
module fifo ( clk, reset, data_in, rd_en, wr_en, empty, full, data_out );
  input [19:0] data_in;
  output [19:0] data_out;
  input clk, reset, rd_en, wr_en;
  output empty, full;
  wire   \buff_mem[19][19] , \buff_mem[19][18] , \buff_mem[19][17] ,
         \buff_mem[19][16] , \buff_mem[19][15] , \buff_mem[19][14] ,
         \buff_mem[19][13] , \buff_mem[19][12] , \buff_mem[19][11] ,
         \buff_mem[19][10] , \buff_mem[19][9] , \buff_mem[19][8] ,
         \buff_mem[19][7] , \buff_mem[19][6] , \buff_mem[19][5] ,
         \buff_mem[19][4] , \buff_mem[19][3] , \buff_mem[19][2] ,
         \buff_mem[19][1] , \buff_mem[19][0] , \buff_mem[18][19] ,
         \buff_mem[18][18] , \buff_mem[18][17] , \buff_mem[18][16] ,
         \buff_mem[18][15] , \buff_mem[18][14] , \buff_mem[18][13] ,
         \buff_mem[18][12] , \buff_mem[18][11] , \buff_mem[18][10] ,
         \buff_mem[18][9] , \buff_mem[18][8] , \buff_mem[18][7] ,
         \buff_mem[18][6] , \buff_mem[18][5] , \buff_mem[18][4] ,
         \buff_mem[18][3] , \buff_mem[18][2] , \buff_mem[18][1] ,
         \buff_mem[18][0] , \buff_mem[17][19] , \buff_mem[17][18] ,
         \buff_mem[17][17] , \buff_mem[17][16] , \buff_mem[17][15] ,
         \buff_mem[17][14] , \buff_mem[17][13] , \buff_mem[17][12] ,
         \buff_mem[17][11] , \buff_mem[17][10] , \buff_mem[17][9] ,
         \buff_mem[17][8] , \buff_mem[17][7] , \buff_mem[17][6] ,
         \buff_mem[17][5] , \buff_mem[17][4] , \buff_mem[17][3] ,
         \buff_mem[17][2] , \buff_mem[17][1] , \buff_mem[17][0] ,
         \buff_mem[16][19] , \buff_mem[16][18] , \buff_mem[16][17] ,
         \buff_mem[16][16] , \buff_mem[16][15] , \buff_mem[16][14] ,
         \buff_mem[16][13] , \buff_mem[16][12] , \buff_mem[16][11] ,
         \buff_mem[16][10] , \buff_mem[16][9] , \buff_mem[16][8] ,
         \buff_mem[16][7] , \buff_mem[16][6] , \buff_mem[16][5] ,
         \buff_mem[16][4] , \buff_mem[16][3] , \buff_mem[16][2] ,
         \buff_mem[16][1] , \buff_mem[16][0] , \buff_mem[15][19] ,
         \buff_mem[15][18] , \buff_mem[15][17] , \buff_mem[15][16] ,
         \buff_mem[15][15] , \buff_mem[15][14] , \buff_mem[15][13] ,
         \buff_mem[15][12] , \buff_mem[15][11] , \buff_mem[15][10] ,
         \buff_mem[15][9] , \buff_mem[15][8] , \buff_mem[15][7] ,
         \buff_mem[15][6] , \buff_mem[15][5] , \buff_mem[15][4] ,
         \buff_mem[15][3] , \buff_mem[15][2] , \buff_mem[15][1] ,
         \buff_mem[15][0] , \buff_mem[14][19] , \buff_mem[14][18] ,
         \buff_mem[14][17] , \buff_mem[14][16] , \buff_mem[14][15] ,
         \buff_mem[14][14] , \buff_mem[14][13] , \buff_mem[14][12] ,
         \buff_mem[14][11] , \buff_mem[14][10] , \buff_mem[14][9] ,
         \buff_mem[14][8] , \buff_mem[14][7] , \buff_mem[14][6] ,
         \buff_mem[14][5] , \buff_mem[14][4] , \buff_mem[14][3] ,
         \buff_mem[14][2] , \buff_mem[14][1] , \buff_mem[14][0] ,
         \buff_mem[13][19] , \buff_mem[13][18] , \buff_mem[13][17] ,
         \buff_mem[13][16] , \buff_mem[13][15] , \buff_mem[13][14] ,
         \buff_mem[13][13] , \buff_mem[13][12] , \buff_mem[13][11] ,
         \buff_mem[13][10] , \buff_mem[13][9] , \buff_mem[13][8] ,
         \buff_mem[13][7] , \buff_mem[13][6] , \buff_mem[13][5] ,
         \buff_mem[13][4] , \buff_mem[13][3] , \buff_mem[13][2] ,
         \buff_mem[13][1] , \buff_mem[13][0] , \buff_mem[12][19] ,
         \buff_mem[12][18] , \buff_mem[12][17] , \buff_mem[12][16] ,
         \buff_mem[12][15] , \buff_mem[12][14] , \buff_mem[12][13] ,
         \buff_mem[12][12] , \buff_mem[12][11] , \buff_mem[12][10] ,
         \buff_mem[12][9] , \buff_mem[12][8] , \buff_mem[12][7] ,
         \buff_mem[12][6] , \buff_mem[12][5] , \buff_mem[12][4] ,
         \buff_mem[12][3] , \buff_mem[12][2] , \buff_mem[12][1] ,
         \buff_mem[12][0] , \buff_mem[11][19] , \buff_mem[11][18] ,
         \buff_mem[11][17] , \buff_mem[11][16] , \buff_mem[11][15] ,
         \buff_mem[11][14] , \buff_mem[11][13] , \buff_mem[11][12] ,
         \buff_mem[11][11] , \buff_mem[11][10] , \buff_mem[11][9] ,
         \buff_mem[11][8] , \buff_mem[11][7] , \buff_mem[11][6] ,
         \buff_mem[11][5] , \buff_mem[11][4] , \buff_mem[11][3] ,
         \buff_mem[11][2] , \buff_mem[11][1] , \buff_mem[11][0] ,
         \buff_mem[10][19] , \buff_mem[10][18] , \buff_mem[10][17] ,
         \buff_mem[10][16] , \buff_mem[10][15] , \buff_mem[10][14] ,
         \buff_mem[10][13] , \buff_mem[10][12] , \buff_mem[10][11] ,
         \buff_mem[10][10] , \buff_mem[10][9] , \buff_mem[10][8] ,
         \buff_mem[10][7] , \buff_mem[10][6] , \buff_mem[10][5] ,
         \buff_mem[10][4] , \buff_mem[10][3] , \buff_mem[10][2] ,
         \buff_mem[10][1] , \buff_mem[10][0] , \buff_mem[9][19] ,
         \buff_mem[9][18] , \buff_mem[9][17] , \buff_mem[9][16] ,
         \buff_mem[9][15] , \buff_mem[9][14] , \buff_mem[9][13] ,
         \buff_mem[9][12] , \buff_mem[9][11] , \buff_mem[9][10] ,
         \buff_mem[9][9] , \buff_mem[9][8] , \buff_mem[9][7] ,
         \buff_mem[9][6] , \buff_mem[9][5] , \buff_mem[9][4] ,
         \buff_mem[9][3] , \buff_mem[9][2] , \buff_mem[9][1] ,
         \buff_mem[9][0] , \buff_mem[8][19] , \buff_mem[8][18] ,
         \buff_mem[8][17] , \buff_mem[8][16] , \buff_mem[8][15] ,
         \buff_mem[8][14] , \buff_mem[8][13] , \buff_mem[8][12] ,
         \buff_mem[8][11] , \buff_mem[8][10] , \buff_mem[8][9] ,
         \buff_mem[8][8] , \buff_mem[8][7] , \buff_mem[8][6] ,
         \buff_mem[8][5] , \buff_mem[8][4] , \buff_mem[8][3] ,
         \buff_mem[8][2] , \buff_mem[8][1] , \buff_mem[8][0] ,
         \buff_mem[7][19] , \buff_mem[7][18] , \buff_mem[7][17] ,
         \buff_mem[7][16] , \buff_mem[7][15] , \buff_mem[7][14] ,
         \buff_mem[7][13] , \buff_mem[7][12] , \buff_mem[7][11] ,
         \buff_mem[7][10] , \buff_mem[7][9] , \buff_mem[7][8] ,
         \buff_mem[7][7] , \buff_mem[7][6] , \buff_mem[7][5] ,
         \buff_mem[7][4] , \buff_mem[7][3] , \buff_mem[7][2] ,
         \buff_mem[7][1] , \buff_mem[7][0] , \buff_mem[6][19] ,
         \buff_mem[6][18] , \buff_mem[6][17] , \buff_mem[6][16] ,
         \buff_mem[6][15] , \buff_mem[6][14] , \buff_mem[6][13] ,
         \buff_mem[6][12] , \buff_mem[6][11] , \buff_mem[6][10] ,
         \buff_mem[6][9] , \buff_mem[6][8] , \buff_mem[6][7] ,
         \buff_mem[6][6] , \buff_mem[6][5] , \buff_mem[6][4] ,
         \buff_mem[6][3] , \buff_mem[6][2] , \buff_mem[6][1] ,
         \buff_mem[6][0] , \buff_mem[5][19] , \buff_mem[5][18] ,
         \buff_mem[5][17] , \buff_mem[5][16] , \buff_mem[5][15] ,
         \buff_mem[5][14] , \buff_mem[5][13] , \buff_mem[5][12] ,
         \buff_mem[5][11] , \buff_mem[5][10] , \buff_mem[5][9] ,
         \buff_mem[5][8] , \buff_mem[5][7] , \buff_mem[5][6] ,
         \buff_mem[5][5] , \buff_mem[5][4] , \buff_mem[5][3] ,
         \buff_mem[5][2] , \buff_mem[5][1] , \buff_mem[5][0] ,
         \buff_mem[4][19] , \buff_mem[4][18] , \buff_mem[4][17] ,
         \buff_mem[4][16] , \buff_mem[4][15] , \buff_mem[4][14] ,
         \buff_mem[4][13] , \buff_mem[4][12] , \buff_mem[4][11] ,
         \buff_mem[4][10] , \buff_mem[4][9] , \buff_mem[4][8] ,
         \buff_mem[4][7] , \buff_mem[4][6] , \buff_mem[4][5] ,
         \buff_mem[4][4] , \buff_mem[4][3] , \buff_mem[4][2] ,
         \buff_mem[4][1] , \buff_mem[4][0] , \buff_mem[3][19] ,
         \buff_mem[3][18] , \buff_mem[3][17] , \buff_mem[3][16] ,
         \buff_mem[3][15] , \buff_mem[3][14] , \buff_mem[3][13] ,
         \buff_mem[3][12] , \buff_mem[3][11] , \buff_mem[3][10] ,
         \buff_mem[3][9] , \buff_mem[3][8] , \buff_mem[3][7] ,
         \buff_mem[3][6] , \buff_mem[3][5] , \buff_mem[3][4] ,
         \buff_mem[3][3] , \buff_mem[3][2] , \buff_mem[3][1] ,
         \buff_mem[3][0] , \buff_mem[2][19] , \buff_mem[2][18] ,
         \buff_mem[2][17] , \buff_mem[2][16] , \buff_mem[2][15] ,
         \buff_mem[2][14] , \buff_mem[2][13] , \buff_mem[2][12] ,
         \buff_mem[2][11] , \buff_mem[2][10] , \buff_mem[2][9] ,
         \buff_mem[2][8] , \buff_mem[2][7] , \buff_mem[2][6] ,
         \buff_mem[2][5] , \buff_mem[2][4] , \buff_mem[2][3] ,
         \buff_mem[2][2] , \buff_mem[2][1] , \buff_mem[2][0] ,
         \buff_mem[1][19] , \buff_mem[1][18] , \buff_mem[1][17] ,
         \buff_mem[1][16] , \buff_mem[1][15] , \buff_mem[1][14] ,
         \buff_mem[1][13] , \buff_mem[1][12] , \buff_mem[1][11] ,
         \buff_mem[1][10] , \buff_mem[1][9] , \buff_mem[1][8] ,
         \buff_mem[1][7] , \buff_mem[1][6] , \buff_mem[1][5] ,
         \buff_mem[1][4] , \buff_mem[1][3] , \buff_mem[1][2] ,
         \buff_mem[1][1] , \buff_mem[1][0] , \buff_mem[0][19] ,
         \buff_mem[0][18] , \buff_mem[0][17] , \buff_mem[0][16] ,
         \buff_mem[0][15] , \buff_mem[0][14] , \buff_mem[0][13] ,
         \buff_mem[0][12] , \buff_mem[0][11] , \buff_mem[0][10] ,
         \buff_mem[0][9] , \buff_mem[0][8] , \buff_mem[0][7] ,
         \buff_mem[0][6] , \buff_mem[0][5] , \buff_mem[0][4] ,
         \buff_mem[0][3] , \buff_mem[0][2] , \buff_mem[0][1] ,
         \buff_mem[0][0] , N142, N143, N144, N145, N146, N147, N148, N149,
         N150, N151, N152, N153, N154, N155, N156, N157, N158, N159, N160,
         N161, n8262, n8263, n4842, n4843, n4852, n4861, n4862, n4863, n4864,
         n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874,
         n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4887, n4888, n4889,
         n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899,
         n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909,
         n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919,
         n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929,
         n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939,
         n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949,
         n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959,
         n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969,
         n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979,
         n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989,
         n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999,
         n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009,
         n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019,
         n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029,
         n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039,
         n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049,
         n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059,
         n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069,
         n5070, n5071, n5072, n5073, n5075, n5076, n5077, n5078, n5079, n5080,
         n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090,
         n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100,
         n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110,
         n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120,
         n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130,
         n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140,
         n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150,
         n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160,
         n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170,
         n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180,
         n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190,
         n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200,
         n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210,
         n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220,
         n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230,
         n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240,
         n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250,
         n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260,
         n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270,
         n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280,
         n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290,
         n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300,
         n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310,
         n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320,
         n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330,
         n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340,
         n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350,
         n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360,
         n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370,
         n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380,
         n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390,
         n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400,
         n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410,
         n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420,
         n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430,
         n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440,
         n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450,
         n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460,
         n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470,
         n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480,
         n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490,
         n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500,
         n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510,
         n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520,
         n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530,
         n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540,
         n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550,
         n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560,
         n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570,
         n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580,
         n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590,
         n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600,
         n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610,
         n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620,
         n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630,
         n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640,
         n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650,
         n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660,
         n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670,
         n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680,
         n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690,
         n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700,
         n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710,
         n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720,
         n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730,
         n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740,
         n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750,
         n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760,
         n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770,
         n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780,
         n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790,
         n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800,
         n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810,
         n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820,
         n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830,
         n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840,
         n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850,
         n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860,
         n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870,
         n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880,
         n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890,
         n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900,
         n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910,
         n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920,
         n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930,
         n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940,
         n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950,
         n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960,
         n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970,
         n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980,
         n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990,
         n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000,
         n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010,
         n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020,
         n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030,
         n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040,
         n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050,
         n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060,
         n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070,
         n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080,
         n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6091,
         n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101,
         n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111,
         n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121,
         n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131,
         n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141,
         n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151,
         n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161,
         n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171,
         n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181,
         n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191,
         n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201,
         n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211,
         n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221,
         n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231,
         n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241,
         n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251,
         n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261,
         n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271,
         n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281,
         n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291,
         n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301,
         n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311,
         n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321,
         n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331,
         n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341,
         n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351,
         n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361,
         n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371,
         n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381,
         n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391,
         n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401,
         n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411,
         n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421,
         n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431,
         n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441,
         n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451,
         n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461,
         n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471,
         n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481,
         n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491,
         n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501,
         n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511,
         n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521,
         n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531,
         n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541,
         n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551,
         n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561,
         n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571,
         n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581,
         n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591,
         n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601,
         n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611,
         n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621,
         n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631,
         n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641,
         n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651,
         n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661,
         n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671,
         n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681,
         n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691,
         n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701,
         n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711,
         n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721,
         n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731,
         n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741,
         n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751,
         n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761,
         n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771,
         n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781,
         n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791,
         n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801,
         n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811,
         n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821,
         n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831,
         n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841,
         n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851,
         n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861,
         n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871,
         n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881,
         n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891,
         n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901,
         n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911,
         n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921,
         n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931,
         n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941,
         n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951,
         n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961,
         n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971,
         n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981,
         n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991,
         n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001,
         n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011,
         n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021,
         n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031,
         n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041,
         n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051,
         n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061,
         n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071,
         n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081,
         n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091,
         n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101,
         n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111,
         n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121,
         n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131,
         n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141,
         n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151,
         n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161,
         n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171,
         n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181,
         n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191,
         n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201,
         n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211,
         n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221,
         n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231,
         n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241,
         n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251,
         n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261,
         n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271,
         n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281,
         n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291,
         n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301,
         n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311,
         n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321,
         n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331,
         n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341,
         n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351,
         n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361,
         n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371,
         n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381,
         n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391,
         n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401,
         n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411,
         n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421,
         n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431,
         n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441,
         n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451,
         n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461,
         n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471,
         n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481,
         n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491,
         n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501,
         n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511,
         n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521,
         n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531,
         n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541,
         n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551,
         n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561,
         n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571,
         n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581,
         n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591,
         n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601,
         n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611,
         n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621,
         n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631,
         n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641,
         n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651,
         n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661,
         n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671,
         n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681,
         n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691,
         n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701,
         n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711,
         n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721,
         n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731,
         n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741,
         n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751,
         n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761,
         n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771,
         n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781,
         n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791,
         n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801,
         n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811,
         n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821,
         n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831,
         n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841,
         n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851,
         n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861,
         n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871,
         n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881,
         n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891,
         n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901,
         n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911,
         n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921,
         n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931,
         n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941,
         n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951,
         n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961,
         n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971,
         n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981,
         n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991,
         n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001,
         n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011,
         n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021,
         n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031,
         n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041,
         n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051,
         n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061,
         n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071,
         n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081,
         n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091,
         n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101,
         n8103, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113,
         n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123,
         n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133,
         n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143,
         n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153,
         n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163,
         n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173,
         n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183,
         n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193,
         n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203,
         n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213,
         n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223,
         n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233,
         n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243,
         n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253,
         n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261;
  wire   [4:0] rd_ptr;
  wire   [4:0] wr_ptr;

  dff_sg \rd_ptr_reg[0]  ( .D(n7257), .CP(clk), .Q(rd_ptr[0]) );
  dff_sg full_reg ( .D(n6888), .CP(clk), .Q(n8263) );
  dff_sg \wr_ptr_reg[0]  ( .D(n7052), .CP(clk), .Q(wr_ptr[0]) );
  dff_sg \wr_ptr_reg[1]  ( .D(n7053), .CP(clk), .Q(wr_ptr[1]) );
  dff_sg \wr_ptr_reg[2]  ( .D(n7054), .CP(clk), .Q(wr_ptr[2]) );
  dff_sg \wr_ptr_reg[3]  ( .D(n7055), .CP(clk), .Q(wr_ptr[3]) );
  dff_sg \wr_ptr_reg[4]  ( .D(n7056), .CP(clk), .Q(wr_ptr[4]) );
  dff_sg \buff_mem_reg[3][12]  ( .D(n7113), .CP(clk), .Q(\buff_mem[3][12] ) );
  dff_sg \buff_mem_reg[2][12]  ( .D(n7076), .CP(clk), .Q(\buff_mem[2][12] ) );
  dff_sg \buff_mem_reg[1][12]  ( .D(n7110), .CP(clk), .Q(\buff_mem[1][12] ) );
  dff_sg \buff_mem_reg[0][12]  ( .D(n7074), .CP(clk), .Q(\buff_mem[0][12] ) );
  dff_sg \buff_mem_reg[19][12]  ( .D(n7137), .CP(clk), .Q(\buff_mem[19][12] )
         );
  dff_sg \buff_mem_reg[18][12]  ( .D(n7156), .CP(clk), .Q(\buff_mem[18][12] )
         );
  dff_sg \buff_mem_reg[17][12]  ( .D(n7179), .CP(clk), .Q(\buff_mem[17][12] )
         );
  dff_sg \buff_mem_reg[16][12]  ( .D(n6876), .CP(clk), .Q(\buff_mem[16][12] )
         );
  dff_sg \buff_mem_reg[15][12]  ( .D(n7048), .CP(clk), .Q(\buff_mem[15][12] )
         );
  dff_sg \buff_mem_reg[14][12]  ( .D(n7024), .CP(clk), .Q(\buff_mem[14][12] )
         );
  dff_sg \buff_mem_reg[13][12]  ( .D(n7014), .CP(clk), .Q(\buff_mem[13][12] )
         );
  dff_sg \buff_mem_reg[12][12]  ( .D(n6859), .CP(clk), .Q(\buff_mem[12][12] )
         );
  dff_sg \buff_mem_reg[11][12]  ( .D(n7220), .CP(clk), .Q(\buff_mem[11][12] )
         );
  dff_sg \buff_mem_reg[10][12]  ( .D(n7216), .CP(clk), .Q(\buff_mem[10][12] )
         );
  dff_sg \buff_mem_reg[9][12]  ( .D(n7242), .CP(clk), .Q(\buff_mem[9][12] ) );
  dff_sg \buff_mem_reg[8][12]  ( .D(n7198), .CP(clk), .Q(\buff_mem[8][12] ) );
  dff_sg \buff_mem_reg[7][12]  ( .D(n6943), .CP(clk), .Q(\buff_mem[7][12] ) );
  dff_sg \buff_mem_reg[6][12]  ( .D(n6997), .CP(clk), .Q(\buff_mem[6][12] ) );
  dff_sg \buff_mem_reg[5][12]  ( .D(n6979), .CP(clk), .Q(\buff_mem[5][12] ) );
  dff_sg \buff_mem_reg[4][12]  ( .D(n6946), .CP(clk), .Q(\buff_mem[4][12] ) );
  dff_sg \buff_mem_reg[3][13]  ( .D(n7125), .CP(clk), .Q(\buff_mem[3][13] ) );
  dff_sg \buff_mem_reg[2][13]  ( .D(n7088), .CP(clk), .Q(\buff_mem[2][13] ) );
  dff_sg \buff_mem_reg[1][13]  ( .D(n7099), .CP(clk), .Q(\buff_mem[1][13] ) );
  dff_sg \buff_mem_reg[0][13]  ( .D(n7066), .CP(clk), .Q(\buff_mem[0][13] ) );
  dff_sg \buff_mem_reg[19][13]  ( .D(n7130), .CP(clk), .Q(\buff_mem[19][13] )
         );
  dff_sg \buff_mem_reg[18][13]  ( .D(n7158), .CP(clk), .Q(\buff_mem[18][13] )
         );
  dff_sg \buff_mem_reg[17][13]  ( .D(n7166), .CP(clk), .Q(\buff_mem[17][13] )
         );
  dff_sg \buff_mem_reg[16][13]  ( .D(n6869), .CP(clk), .Q(\buff_mem[16][13] )
         );
  dff_sg \buff_mem_reg[15][13]  ( .D(n7044), .CP(clk), .Q(\buff_mem[15][13] )
         );
  dff_sg \buff_mem_reg[14][13]  ( .D(n7031), .CP(clk), .Q(\buff_mem[14][13] )
         );
  dff_sg \buff_mem_reg[13][13]  ( .D(n7008), .CP(clk), .Q(\buff_mem[13][13] )
         );
  dff_sg \buff_mem_reg[12][13]  ( .D(n6851), .CP(clk), .Q(\buff_mem[12][13] )
         );
  dff_sg \buff_mem_reg[11][13]  ( .D(n7232), .CP(clk), .Q(\buff_mem[11][13] )
         );
  dff_sg \buff_mem_reg[10][13]  ( .D(n7212), .CP(clk), .Q(\buff_mem[10][13] )
         );
  dff_sg \buff_mem_reg[9][13]  ( .D(n7248), .CP(clk), .Q(\buff_mem[9][13] ) );
  dff_sg \buff_mem_reg[8][13]  ( .D(n7194), .CP(clk), .Q(\buff_mem[8][13] ) );
  dff_sg \buff_mem_reg[7][13]  ( .D(n6937), .CP(clk), .Q(\buff_mem[7][13] ) );
  dff_sg \buff_mem_reg[6][13]  ( .D(n6982), .CP(clk), .Q(\buff_mem[6][13] ) );
  dff_sg \buff_mem_reg[5][13]  ( .D(n6971), .CP(clk), .Q(\buff_mem[5][13] ) );
  dff_sg \buff_mem_reg[4][13]  ( .D(n6958), .CP(clk), .Q(\buff_mem[4][13] ) );
  dff_sg \buff_mem_reg[3][14]  ( .D(n7114), .CP(clk), .Q(\buff_mem[3][14] ) );
  dff_sg \buff_mem_reg[2][14]  ( .D(n7078), .CP(clk), .Q(\buff_mem[2][14] ) );
  dff_sg \buff_mem_reg[1][14]  ( .D(n7093), .CP(clk), .Q(\buff_mem[1][14] ) );
  dff_sg \buff_mem_reg[0][14]  ( .D(n7058), .CP(clk), .Q(\buff_mem[0][14] ) );
  dff_sg \buff_mem_reg[19][14]  ( .D(n7132), .CP(clk), .Q(\buff_mem[19][14] )
         );
  dff_sg \buff_mem_reg[18][14]  ( .D(n7147), .CP(clk), .Q(\buff_mem[18][14] )
         );
  dff_sg \buff_mem_reg[17][14]  ( .D(n7168), .CP(clk), .Q(\buff_mem[17][14] )
         );
  dff_sg \buff_mem_reg[16][14]  ( .D(n6871), .CP(clk), .Q(\buff_mem[16][14] )
         );
  dff_sg \buff_mem_reg[15][14]  ( .D(n7041), .CP(clk), .Q(\buff_mem[15][14] )
         );
  dff_sg \buff_mem_reg[14][14]  ( .D(n7019), .CP(clk), .Q(\buff_mem[14][14] )
         );
  dff_sg \buff_mem_reg[13][14]  ( .D(n7000), .CP(clk), .Q(\buff_mem[13][14] )
         );
  dff_sg \buff_mem_reg[12][14]  ( .D(n6848), .CP(clk), .Q(\buff_mem[12][14] )
         );
  dff_sg \buff_mem_reg[11][14]  ( .D(n7222), .CP(clk), .Q(\buff_mem[11][14] )
         );
  dff_sg \buff_mem_reg[10][14]  ( .D(n7204), .CP(clk), .Q(\buff_mem[10][14] )
         );
  dff_sg \buff_mem_reg[9][14]  ( .D(n7237), .CP(clk), .Q(\buff_mem[9][14] ) );
  dff_sg \buff_mem_reg[8][14]  ( .D(n7186), .CP(clk), .Q(\buff_mem[8][14] ) );
  dff_sg \buff_mem_reg[7][14]  ( .D(n6927), .CP(clk), .Q(\buff_mem[7][14] ) );
  dff_sg \buff_mem_reg[6][14]  ( .D(n6989), .CP(clk), .Q(\buff_mem[6][14] ) );
  dff_sg \buff_mem_reg[5][14]  ( .D(n6964), .CP(clk), .Q(\buff_mem[5][14] ) );
  dff_sg \buff_mem_reg[4][14]  ( .D(n6956), .CP(clk), .Q(\buff_mem[4][14] ) );
  dff_sg \buff_mem_reg[3][15]  ( .D(n7128), .CP(clk), .Q(\buff_mem[3][15] ) );
  dff_sg \buff_mem_reg[2][15]  ( .D(n7092), .CP(clk), .Q(\buff_mem[2][15] ) );
  dff_sg \buff_mem_reg[1][15]  ( .D(n7100), .CP(clk), .Q(\buff_mem[1][15] ) );
  dff_sg \buff_mem_reg[0][15]  ( .D(n7057), .CP(clk), .Q(\buff_mem[0][15] ) );
  dff_sg \buff_mem_reg[19][15]  ( .D(n7146), .CP(clk), .Q(\buff_mem[19][15] )
         );
  dff_sg \buff_mem_reg[18][15]  ( .D(n7159), .CP(clk), .Q(\buff_mem[18][15] )
         );
  dff_sg \buff_mem_reg[17][15]  ( .D(n7182), .CP(clk), .Q(\buff_mem[17][15] )
         );
  dff_sg \buff_mem_reg[16][15]  ( .D(n6886), .CP(clk), .Q(\buff_mem[16][15] )
         );
  dff_sg \buff_mem_reg[15][15]  ( .D(n7035), .CP(clk), .Q(\buff_mem[15][15] )
         );
  dff_sg \buff_mem_reg[14][15]  ( .D(n7033), .CP(clk), .Q(\buff_mem[14][15] )
         );
  dff_sg \buff_mem_reg[13][15]  ( .D(n6999), .CP(clk), .Q(\buff_mem[13][15] )
         );
  dff_sg \buff_mem_reg[12][15]  ( .D(n6854), .CP(clk), .Q(\buff_mem[12][15] )
         );
  dff_sg \buff_mem_reg[11][15]  ( .D(n7236), .CP(clk), .Q(\buff_mem[11][15] )
         );
  dff_sg \buff_mem_reg[10][15]  ( .D(n7217), .CP(clk), .Q(\buff_mem[10][15] )
         );
  dff_sg \buff_mem_reg[9][15]  ( .D(n7243), .CP(clk), .Q(\buff_mem[9][15] ) );
  dff_sg \buff_mem_reg[8][15]  ( .D(n7199), .CP(clk), .Q(\buff_mem[8][15] ) );
  dff_sg \buff_mem_reg[7][15]  ( .D(n6926), .CP(clk), .Q(\buff_mem[7][15] ) );
  dff_sg \buff_mem_reg[6][15]  ( .D(n6985), .CP(clk), .Q(\buff_mem[6][15] ) );
  dff_sg \buff_mem_reg[5][15]  ( .D(n6963), .CP(clk), .Q(\buff_mem[5][15] ) );
  dff_sg \buff_mem_reg[4][15]  ( .D(n6948), .CP(clk), .Q(\buff_mem[4][15] ) );
  dff_sg \buff_mem_reg[3][16]  ( .D(n7120), .CP(clk), .Q(\buff_mem[3][16] ) );
  dff_sg \buff_mem_reg[2][16]  ( .D(n7084), .CP(clk), .Q(\buff_mem[2][16] ) );
  dff_sg \buff_mem_reg[1][16]  ( .D(n7107), .CP(clk), .Q(\buff_mem[1][16] ) );
  dff_sg \buff_mem_reg[0][16]  ( .D(n7069), .CP(clk), .Q(\buff_mem[0][16] ) );
  dff_sg \buff_mem_reg[19][16]  ( .D(n7143), .CP(clk), .Q(\buff_mem[19][16] )
         );
  dff_sg \buff_mem_reg[18][16]  ( .D(n7161), .CP(clk), .Q(\buff_mem[18][16] )
         );
  dff_sg \buff_mem_reg[17][16]  ( .D(n7174), .CP(clk), .Q(\buff_mem[17][16] )
         );
  dff_sg \buff_mem_reg[16][16]  ( .D(n6883), .CP(clk), .Q(\buff_mem[16][16] )
         );
  dff_sg \buff_mem_reg[15][16]  ( .D(n7051), .CP(clk), .Q(\buff_mem[15][16] )
         );
  dff_sg \buff_mem_reg[14][16]  ( .D(n7017), .CP(clk), .Q(\buff_mem[14][16] )
         );
  dff_sg \buff_mem_reg[13][16]  ( .D(n7009), .CP(clk), .Q(\buff_mem[13][16] )
         );
  dff_sg \buff_mem_reg[12][16]  ( .D(n6864), .CP(clk), .Q(\buff_mem[12][16] )
         );
  dff_sg \buff_mem_reg[11][16]  ( .D(n7228), .CP(clk), .Q(\buff_mem[11][16] )
         );
  dff_sg \buff_mem_reg[10][16]  ( .D(n7214), .CP(clk), .Q(\buff_mem[10][16] )
         );
  dff_sg \buff_mem_reg[9][16]  ( .D(n7251), .CP(clk), .Q(\buff_mem[9][16] ) );
  dff_sg \buff_mem_reg[8][16]  ( .D(n7196), .CP(clk), .Q(\buff_mem[8][16] ) );
  dff_sg \buff_mem_reg[7][16]  ( .D(n6938), .CP(clk), .Q(\buff_mem[7][16] ) );
  dff_sg \buff_mem_reg[6][16]  ( .D(n6994), .CP(clk), .Q(\buff_mem[6][16] ) );
  dff_sg \buff_mem_reg[5][16]  ( .D(n6974), .CP(clk), .Q(\buff_mem[5][16] ) );
  dff_sg \buff_mem_reg[4][16]  ( .D(n6955), .CP(clk), .Q(\buff_mem[4][16] ) );
  dff_sg \buff_mem_reg[3][17]  ( .D(n7119), .CP(clk), .Q(\buff_mem[3][17] ) );
  dff_sg \buff_mem_reg[2][17]  ( .D(n7086), .CP(clk), .Q(\buff_mem[2][17] ) );
  dff_sg \buff_mem_reg[1][17]  ( .D(n7097), .CP(clk), .Q(\buff_mem[1][17] ) );
  dff_sg \buff_mem_reg[0][17]  ( .D(n7064), .CP(clk), .Q(\buff_mem[0][17] ) );
  dff_sg \buff_mem_reg[19][17]  ( .D(n7138), .CP(clk), .Q(\buff_mem[19][17] )
         );
  dff_sg \buff_mem_reg[18][17]  ( .D(n7157), .CP(clk), .Q(\buff_mem[18][17] )
         );
  dff_sg \buff_mem_reg[17][17]  ( .D(n7176), .CP(clk), .Q(\buff_mem[17][17] )
         );
  dff_sg \buff_mem_reg[16][17]  ( .D(n6881), .CP(clk), .Q(\buff_mem[16][17] )
         );
  dff_sg \buff_mem_reg[15][17]  ( .D(n7045), .CP(clk), .Q(\buff_mem[15][17] )
         );
  dff_sg \buff_mem_reg[14][17]  ( .D(n7030), .CP(clk), .Q(\buff_mem[14][17] )
         );
  dff_sg \buff_mem_reg[13][17]  ( .D(n7006), .CP(clk), .Q(\buff_mem[13][17] )
         );
  dff_sg \buff_mem_reg[12][17]  ( .D(n6861), .CP(clk), .Q(\buff_mem[12][17] )
         );
  dff_sg \buff_mem_reg[11][17]  ( .D(n7227), .CP(clk), .Q(\buff_mem[11][17] )
         );
  dff_sg \buff_mem_reg[10][17]  ( .D(n7210), .CP(clk), .Q(\buff_mem[10][17] )
         );
  dff_sg \buff_mem_reg[9][17]  ( .D(n7247), .CP(clk), .Q(\buff_mem[9][17] ) );
  dff_sg \buff_mem_reg[8][17]  ( .D(n7191), .CP(clk), .Q(\buff_mem[8][17] ) );
  dff_sg \buff_mem_reg[7][17]  ( .D(n6935), .CP(clk), .Q(\buff_mem[7][17] ) );
  dff_sg \buff_mem_reg[6][17]  ( .D(n6983), .CP(clk), .Q(\buff_mem[6][17] ) );
  dff_sg \buff_mem_reg[5][17]  ( .D(n6969), .CP(clk), .Q(\buff_mem[5][17] ) );
  dff_sg \buff_mem_reg[4][17]  ( .D(n6951), .CP(clk), .Q(\buff_mem[4][17] ) );
  dff_sg \buff_mem_reg[3][18]  ( .D(n7117), .CP(clk), .Q(\buff_mem[3][18] ) );
  dff_sg \buff_mem_reg[2][18]  ( .D(n7081), .CP(clk), .Q(\buff_mem[2][18] ) );
  dff_sg \buff_mem_reg[1][18]  ( .D(n7105), .CP(clk), .Q(\buff_mem[1][18] ) );
  dff_sg \buff_mem_reg[0][18]  ( .D(n7061), .CP(clk), .Q(\buff_mem[0][18] ) );
  dff_sg \buff_mem_reg[19][18]  ( .D(n7144), .CP(clk), .Q(\buff_mem[19][18] )
         );
  dff_sg \buff_mem_reg[18][18]  ( .D(n7150), .CP(clk), .Q(\buff_mem[18][18] )
         );
  dff_sg \buff_mem_reg[17][18]  ( .D(n7165), .CP(clk), .Q(\buff_mem[17][18] )
         );
  dff_sg \buff_mem_reg[16][18]  ( .D(n6868), .CP(clk), .Q(\buff_mem[16][18] )
         );
  dff_sg \buff_mem_reg[15][18]  ( .D(n7042), .CP(clk), .Q(\buff_mem[15][18] )
         );
  dff_sg \buff_mem_reg[14][18]  ( .D(n7022), .CP(clk), .Q(\buff_mem[14][18] )
         );
  dff_sg \buff_mem_reg[13][18]  ( .D(n7003), .CP(clk), .Q(\buff_mem[13][18] )
         );
  dff_sg \buff_mem_reg[12][18]  ( .D(n6860), .CP(clk), .Q(\buff_mem[12][18] )
         );
  dff_sg \buff_mem_reg[11][18]  ( .D(n7225), .CP(clk), .Q(\buff_mem[11][18] )
         );
  dff_sg \buff_mem_reg[10][18]  ( .D(n7207), .CP(clk), .Q(\buff_mem[10][18] )
         );
  dff_sg \buff_mem_reg[9][18]  ( .D(n7246), .CP(clk), .Q(\buff_mem[9][18] ) );
  dff_sg \buff_mem_reg[8][18]  ( .D(n7189), .CP(clk), .Q(\buff_mem[8][18] ) );
  dff_sg \buff_mem_reg[7][18]  ( .D(n6930), .CP(clk), .Q(\buff_mem[7][18] ) );
  dff_sg \buff_mem_reg[6][18]  ( .D(n6981), .CP(clk), .Q(\buff_mem[6][18] ) );
  dff_sg \buff_mem_reg[5][18]  ( .D(n6967), .CP(clk), .Q(\buff_mem[5][18] ) );
  dff_sg \buff_mem_reg[4][18]  ( .D(n6959), .CP(clk), .Q(\buff_mem[4][18] ) );
  dff_sg \buff_mem_reg[3][19]  ( .D(n7112), .CP(clk), .Q(\buff_mem[3][19] ) );
  dff_sg \buff_mem_reg[2][19]  ( .D(n7075), .CP(clk), .Q(\buff_mem[2][19] ) );
  dff_sg \buff_mem_reg[1][19]  ( .D(n7102), .CP(clk), .Q(\buff_mem[1][19] ) );
  dff_sg \buff_mem_reg[0][19]  ( .D(n7068), .CP(clk), .Q(\buff_mem[0][19] ) );
  dff_sg \buff_mem_reg[19][19]  ( .D(n7133), .CP(clk), .Q(\buff_mem[19][19] )
         );
  dff_sg \buff_mem_reg[18][19]  ( .D(n7155), .CP(clk), .Q(\buff_mem[18][19] )
         );
  dff_sg \buff_mem_reg[17][19]  ( .D(n7169), .CP(clk), .Q(\buff_mem[17][19] )
         );
  dff_sg \buff_mem_reg[16][19]  ( .D(n6872), .CP(clk), .Q(\buff_mem[16][19] )
         );
  dff_sg \buff_mem_reg[15][19]  ( .D(n7047), .CP(clk), .Q(\buff_mem[15][19] )
         );
  dff_sg \buff_mem_reg[14][19]  ( .D(n7028), .CP(clk), .Q(\buff_mem[14][19] )
         );
  dff_sg \buff_mem_reg[13][19]  ( .D(n7005), .CP(clk), .Q(\buff_mem[13][19] )
         );
  dff_sg \buff_mem_reg[12][19]  ( .D(n6858), .CP(clk), .Q(\buff_mem[12][19] )
         );
  dff_sg \buff_mem_reg[11][19]  ( .D(n7219), .CP(clk), .Q(\buff_mem[11][19] )
         );
  dff_sg \buff_mem_reg[10][19]  ( .D(n7202), .CP(clk), .Q(\buff_mem[10][19] )
         );
  dff_sg \buff_mem_reg[9][19]  ( .D(n7241), .CP(clk), .Q(\buff_mem[9][19] ) );
  dff_sg \buff_mem_reg[8][19]  ( .D(n7184), .CP(clk), .Q(\buff_mem[8][19] ) );
  dff_sg \buff_mem_reg[7][19]  ( .D(n6933), .CP(clk), .Q(\buff_mem[7][19] ) );
  dff_sg \buff_mem_reg[6][19]  ( .D(n6991), .CP(clk), .Q(\buff_mem[6][19] ) );
  dff_sg \buff_mem_reg[5][19]  ( .D(n6973), .CP(clk), .Q(\buff_mem[5][19] ) );
  dff_sg \buff_mem_reg[4][19]  ( .D(n6944), .CP(clk), .Q(\buff_mem[4][19] ) );
  dff_sg \buff_mem_reg[4][0]  ( .D(n6898), .CP(clk), .Q(\buff_mem[4][0] ) );
  dff_sg \buff_mem_reg[3][0]  ( .D(n6897), .CP(clk), .Q(\buff_mem[3][0] ) );
  dff_sg \buff_mem_reg[2][0]  ( .D(n6894), .CP(clk), .Q(\buff_mem[2][0] ) );
  dff_sg \buff_mem_reg[1][0]  ( .D(n6896), .CP(clk), .Q(\buff_mem[1][0] ) );
  dff_sg \buff_mem_reg[0][0]  ( .D(n6899), .CP(clk), .Q(\buff_mem[0][0] ) );
  dff_sg \buff_mem_reg[19][0]  ( .D(n6895), .CP(clk), .Q(\buff_mem[19][0] ) );
  dff_sg \buff_mem_reg[18][0]  ( .D(n6892), .CP(clk), .Q(\buff_mem[18][0] ) );
  dff_sg \buff_mem_reg[17][0]  ( .D(n6901), .CP(clk), .Q(\buff_mem[17][0] ) );
  dff_sg \buff_mem_reg[16][0]  ( .D(n6887), .CP(clk), .Q(\buff_mem[16][0] ) );
  dff_sg \buff_mem_reg[15][0]  ( .D(n6889), .CP(clk), .Q(\buff_mem[15][0] ) );
  dff_sg \buff_mem_reg[14][0]  ( .D(n6900), .CP(clk), .Q(\buff_mem[14][0] ) );
  dff_sg \buff_mem_reg[13][0]  ( .D(n6893), .CP(clk), .Q(\buff_mem[13][0] ) );
  dff_sg \buff_mem_reg[12][0]  ( .D(n6852), .CP(clk), .Q(\buff_mem[12][0] ) );
  dff_sg \buff_mem_reg[11][0]  ( .D(n6904), .CP(clk), .Q(\buff_mem[11][0] ) );
  dff_sg \buff_mem_reg[10][0]  ( .D(n6902), .CP(clk), .Q(\buff_mem[10][0] ) );
  dff_sg \buff_mem_reg[9][0]  ( .D(n6905), .CP(clk), .Q(\buff_mem[9][0] ) );
  dff_sg \buff_mem_reg[8][0]  ( .D(n6891), .CP(clk), .Q(\buff_mem[8][0] ) );
  dff_sg \buff_mem_reg[7][0]  ( .D(n6903), .CP(clk), .Q(\buff_mem[7][0] ) );
  dff_sg \buff_mem_reg[6][0]  ( .D(n6906), .CP(clk), .Q(\buff_mem[6][0] ) );
  dff_sg \buff_mem_reg[5][0]  ( .D(n6890), .CP(clk), .Q(\buff_mem[5][0] ) );
  dff_sg \buff_mem_reg[4][1]  ( .D(n6960), .CP(clk), .Q(\buff_mem[4][1] ) );
  dff_sg \buff_mem_reg[3][1]  ( .D(n7124), .CP(clk), .Q(\buff_mem[3][1] ) );
  dff_sg \buff_mem_reg[2][1]  ( .D(n7087), .CP(clk), .Q(\buff_mem[2][1] ) );
  dff_sg \buff_mem_reg[1][1]  ( .D(n7106), .CP(clk), .Q(\buff_mem[1][1] ) );
  dff_sg \buff_mem_reg[0][1]  ( .D(n7065), .CP(clk), .Q(\buff_mem[0][1] ) );
  dff_sg \buff_mem_reg[19][1]  ( .D(n7139), .CP(clk), .Q(\buff_mem[19][1] ) );
  dff_sg \buff_mem_reg[18][1]  ( .D(n7160), .CP(clk), .Q(\buff_mem[18][1] ) );
  dff_sg \buff_mem_reg[17][1]  ( .D(n7177), .CP(clk), .Q(\buff_mem[17][1] ) );
  dff_sg \buff_mem_reg[16][1]  ( .D(n6882), .CP(clk), .Q(\buff_mem[16][1] ) );
  dff_sg \buff_mem_reg[15][1]  ( .D(n7050), .CP(clk), .Q(\buff_mem[15][1] ) );
  dff_sg \buff_mem_reg[14][1]  ( .D(n7016), .CP(clk), .Q(\buff_mem[14][1] ) );
  dff_sg \buff_mem_reg[13][1]  ( .D(n7007), .CP(clk), .Q(\buff_mem[13][1] ) );
  dff_sg \buff_mem_reg[12][1]  ( .D(n6863), .CP(clk), .Q(\buff_mem[12][1] ) );
  dff_sg \buff_mem_reg[11][1]  ( .D(n7231), .CP(clk), .Q(\buff_mem[11][1] ) );
  dff_sg \buff_mem_reg[10][1]  ( .D(n7211), .CP(clk), .Q(\buff_mem[10][1] ) );
  dff_sg \buff_mem_reg[9][1]  ( .D(n7250), .CP(clk), .Q(\buff_mem[9][1] ) );
  dff_sg \buff_mem_reg[8][1]  ( .D(n7193), .CP(clk), .Q(\buff_mem[8][1] ) );
  dff_sg \buff_mem_reg[7][1]  ( .D(n6936), .CP(clk), .Q(\buff_mem[7][1] ) );
  dff_sg \buff_mem_reg[6][1]  ( .D(n6993), .CP(clk), .Q(\buff_mem[6][1] ) );
  dff_sg \buff_mem_reg[5][1]  ( .D(n6970), .CP(clk), .Q(\buff_mem[5][1] ) );
  dff_sg \buff_mem_reg[4][2]  ( .D(n6949), .CP(clk), .Q(\buff_mem[4][2] ) );
  dff_sg \buff_mem_reg[3][2]  ( .D(n7122), .CP(clk), .Q(\buff_mem[3][2] ) );
  dff_sg \buff_mem_reg[2][2]  ( .D(n7089), .CP(clk), .Q(\buff_mem[2][2] ) );
  dff_sg \buff_mem_reg[1][2]  ( .D(n7104), .CP(clk), .Q(\buff_mem[1][2] ) );
  dff_sg \buff_mem_reg[0][2]  ( .D(n7067), .CP(clk), .Q(\buff_mem[0][2] ) );
  dff_sg \buff_mem_reg[19][2]  ( .D(n7141), .CP(clk), .Q(\buff_mem[19][2] ) );
  dff_sg \buff_mem_reg[18][2]  ( .D(n7152), .CP(clk), .Q(\buff_mem[18][2] ) );
  dff_sg \buff_mem_reg[17][2]  ( .D(n7173), .CP(clk), .Q(\buff_mem[17][2] ) );
  dff_sg \buff_mem_reg[16][2]  ( .D(n6877), .CP(clk), .Q(\buff_mem[16][2] ) );
  dff_sg \buff_mem_reg[15][2]  ( .D(n7037), .CP(clk), .Q(\buff_mem[15][2] ) );
  dff_sg \buff_mem_reg[14][2]  ( .D(n7027), .CP(clk), .Q(\buff_mem[14][2] ) );
  dff_sg \buff_mem_reg[13][2]  ( .D(n7012), .CP(clk), .Q(\buff_mem[13][2] ) );
  dff_sg \buff_mem_reg[12][2]  ( .D(n6855), .CP(clk), .Q(\buff_mem[12][2] ) );
  dff_sg \buff_mem_reg[11][2]  ( .D(n7233), .CP(clk), .Q(\buff_mem[11][2] ) );
  dff_sg \buff_mem_reg[10][2]  ( .D(n7209), .CP(clk), .Q(\buff_mem[10][2] ) );
  dff_sg \buff_mem_reg[9][2]  ( .D(n7244), .CP(clk), .Q(\buff_mem[9][2] ) );
  dff_sg \buff_mem_reg[8][2]  ( .D(n7195), .CP(clk), .Q(\buff_mem[8][2] ) );
  dff_sg \buff_mem_reg[7][2]  ( .D(n6934), .CP(clk), .Q(\buff_mem[7][2] ) );
  dff_sg \buff_mem_reg[6][2]  ( .D(n6990), .CP(clk), .Q(\buff_mem[6][2] ) );
  dff_sg \buff_mem_reg[5][2]  ( .D(n6972), .CP(clk), .Q(\buff_mem[5][2] ) );
  dff_sg \buff_mem_reg[4][3]  ( .D(n6953), .CP(clk), .Q(\buff_mem[4][3] ) );
  dff_sg \buff_mem_reg[3][3]  ( .D(n7115), .CP(clk), .Q(\buff_mem[3][3] ) );
  dff_sg \buff_mem_reg[2][3]  ( .D(n7079), .CP(clk), .Q(\buff_mem[2][3] ) );
  dff_sg \buff_mem_reg[1][3]  ( .D(n7094), .CP(clk), .Q(\buff_mem[1][3] ) );
  dff_sg \buff_mem_reg[0][3]  ( .D(n7059), .CP(clk), .Q(\buff_mem[0][3] ) );
  dff_sg \buff_mem_reg[19][3]  ( .D(n7129), .CP(clk), .Q(\buff_mem[19][3] ) );
  dff_sg \buff_mem_reg[18][3]  ( .D(n7148), .CP(clk), .Q(\buff_mem[18][3] ) );
  dff_sg \buff_mem_reg[17][3]  ( .D(n7180), .CP(clk), .Q(\buff_mem[17][3] ) );
  dff_sg \buff_mem_reg[16][3]  ( .D(n6884), .CP(clk), .Q(\buff_mem[16][3] ) );
  dff_sg \buff_mem_reg[15][3]  ( .D(n7043), .CP(clk), .Q(\buff_mem[15][3] ) );
  dff_sg \buff_mem_reg[14][3]  ( .D(n7020), .CP(clk), .Q(\buff_mem[14][3] ) );
  dff_sg \buff_mem_reg[13][3]  ( .D(n7001), .CP(clk), .Q(\buff_mem[13][3] ) );
  dff_sg \buff_mem_reg[12][3]  ( .D(n6849), .CP(clk), .Q(\buff_mem[12][3] ) );
  dff_sg \buff_mem_reg[11][3]  ( .D(n7223), .CP(clk), .Q(\buff_mem[11][3] ) );
  dff_sg \buff_mem_reg[10][3]  ( .D(n7205), .CP(clk), .Q(\buff_mem[10][3] ) );
  dff_sg \buff_mem_reg[9][3]  ( .D(n7238), .CP(clk), .Q(\buff_mem[9][3] ) );
  dff_sg \buff_mem_reg[8][3]  ( .D(n7187), .CP(clk), .Q(\buff_mem[8][3] ) );
  dff_sg \buff_mem_reg[7][3]  ( .D(n6928), .CP(clk), .Q(\buff_mem[7][3] ) );
  dff_sg \buff_mem_reg[6][3]  ( .D(n6987), .CP(clk), .Q(\buff_mem[6][3] ) );
  dff_sg \buff_mem_reg[5][3]  ( .D(n6965), .CP(clk), .Q(\buff_mem[5][3] ) );
  dff_sg \buff_mem_reg[4][4]  ( .D(n6961), .CP(clk), .Q(\buff_mem[4][4] ) );
  dff_sg \buff_mem_reg[3][4]  ( .D(n7111), .CP(clk), .Q(\buff_mem[3][4] ) );
  dff_sg \buff_mem_reg[2][4]  ( .D(n7083), .CP(clk), .Q(\buff_mem[2][4] ) );
  dff_sg \buff_mem_reg[1][4]  ( .D(n7103), .CP(clk), .Q(\buff_mem[1][4] ) );
  dff_sg \buff_mem_reg[0][4]  ( .D(n7070), .CP(clk), .Q(\buff_mem[0][4] ) );
  dff_sg \buff_mem_reg[19][4]  ( .D(n7134), .CP(clk), .Q(\buff_mem[19][4] ) );
  dff_sg \buff_mem_reg[18][4]  ( .D(n7164), .CP(clk), .Q(\buff_mem[18][4] ) );
  dff_sg \buff_mem_reg[17][4]  ( .D(n7170), .CP(clk), .Q(\buff_mem[17][4] ) );
  dff_sg \buff_mem_reg[16][4]  ( .D(n6873), .CP(clk), .Q(\buff_mem[16][4] ) );
  dff_sg \buff_mem_reg[15][4]  ( .D(n7040), .CP(clk), .Q(\buff_mem[15][4] ) );
  dff_sg \buff_mem_reg[14][4]  ( .D(n7025), .CP(clk), .Q(\buff_mem[14][4] ) );
  dff_sg \buff_mem_reg[13][4]  ( .D(n7010), .CP(clk), .Q(\buff_mem[13][4] ) );
  dff_sg \buff_mem_reg[12][4]  ( .D(n6867), .CP(clk), .Q(\buff_mem[12][4] ) );
  dff_sg \buff_mem_reg[11][4]  ( .D(n7229), .CP(clk), .Q(\buff_mem[11][4] ) );
  dff_sg \buff_mem_reg[10][4]  ( .D(n7201), .CP(clk), .Q(\buff_mem[10][4] ) );
  dff_sg \buff_mem_reg[9][4]  ( .D(n7254), .CP(clk), .Q(\buff_mem[9][4] ) );
  dff_sg \buff_mem_reg[8][4]  ( .D(n7183), .CP(clk), .Q(\buff_mem[8][4] ) );
  dff_sg \buff_mem_reg[7][4]  ( .D(n6939), .CP(clk), .Q(\buff_mem[7][4] ) );
  dff_sg \buff_mem_reg[6][4]  ( .D(n6996), .CP(clk), .Q(\buff_mem[6][4] ) );
  dff_sg \buff_mem_reg[5][4]  ( .D(n6975), .CP(clk), .Q(\buff_mem[5][4] ) );
  dff_sg \buff_mem_reg[4][5]  ( .D(n6952), .CP(clk), .Q(\buff_mem[4][5] ) );
  dff_sg \buff_mem_reg[3][5]  ( .D(n7118), .CP(clk), .Q(\buff_mem[3][5] ) );
  dff_sg \buff_mem_reg[2][5]  ( .D(n7082), .CP(clk), .Q(\buff_mem[2][5] ) );
  dff_sg \buff_mem_reg[1][5]  ( .D(n7108), .CP(clk), .Q(\buff_mem[1][5] ) );
  dff_sg \buff_mem_reg[0][5]  ( .D(n7062), .CP(clk), .Q(\buff_mem[0][5] ) );
  dff_sg \buff_mem_reg[19][5]  ( .D(n7136), .CP(clk), .Q(\buff_mem[19][5] ) );
  dff_sg \buff_mem_reg[18][5]  ( .D(n7162), .CP(clk), .Q(\buff_mem[18][5] ) );
  dff_sg \buff_mem_reg[17][5]  ( .D(n7172), .CP(clk), .Q(\buff_mem[17][5] ) );
  dff_sg \buff_mem_reg[16][5]  ( .D(n6875), .CP(clk), .Q(\buff_mem[16][5] ) );
  dff_sg \buff_mem_reg[15][5]  ( .D(n7034), .CP(clk), .Q(\buff_mem[15][5] ) );
  dff_sg \buff_mem_reg[14][5]  ( .D(n7023), .CP(clk), .Q(\buff_mem[14][5] ) );
  dff_sg \buff_mem_reg[13][5]  ( .D(n7004), .CP(clk), .Q(\buff_mem[13][5] ) );
  dff_sg \buff_mem_reg[12][5]  ( .D(n6865), .CP(clk), .Q(\buff_mem[12][5] ) );
  dff_sg \buff_mem_reg[11][5]  ( .D(n7226), .CP(clk), .Q(\buff_mem[11][5] ) );
  dff_sg \buff_mem_reg[10][5]  ( .D(n7208), .CP(clk), .Q(\buff_mem[10][5] ) );
  dff_sg \buff_mem_reg[9][5]  ( .D(n7252), .CP(clk), .Q(\buff_mem[9][5] ) );
  dff_sg \buff_mem_reg[8][5]  ( .D(n7190), .CP(clk), .Q(\buff_mem[8][5] ) );
  dff_sg \buff_mem_reg[7][5]  ( .D(n6931), .CP(clk), .Q(\buff_mem[7][5] ) );
  dff_sg \buff_mem_reg[6][5]  ( .D(n6995), .CP(clk), .Q(\buff_mem[6][5] ) );
  dff_sg \buff_mem_reg[5][5]  ( .D(n6968), .CP(clk), .Q(\buff_mem[5][5] ) );
  dff_sg \buff_mem_reg[4][6]  ( .D(n6947), .CP(clk), .Q(\buff_mem[4][6] ) );
  dff_sg \buff_mem_reg[3][6]  ( .D(n7126), .CP(clk), .Q(\buff_mem[3][6] ) );
  dff_sg \buff_mem_reg[2][6]  ( .D(n7091), .CP(clk), .Q(\buff_mem[2][6] ) );
  dff_sg \buff_mem_reg[1][6]  ( .D(n7098), .CP(clk), .Q(\buff_mem[1][6] ) );
  dff_sg \buff_mem_reg[0][6]  ( .D(n7073), .CP(clk), .Q(\buff_mem[0][6] ) );
  dff_sg \buff_mem_reg[19][6]  ( .D(n7145), .CP(clk), .Q(\buff_mem[19][6] ) );
  dff_sg \buff_mem_reg[18][6]  ( .D(n7153), .CP(clk), .Q(\buff_mem[18][6] ) );
  dff_sg \buff_mem_reg[17][6]  ( .D(n7181), .CP(clk), .Q(\buff_mem[17][6] ) );
  dff_sg \buff_mem_reg[16][6]  ( .D(n6885), .CP(clk), .Q(\buff_mem[16][6] ) );
  dff_sg \buff_mem_reg[15][6]  ( .D(n7046), .CP(clk), .Q(\buff_mem[15][6] ) );
  dff_sg \buff_mem_reg[14][6]  ( .D(n7032), .CP(clk), .Q(\buff_mem[14][6] ) );
  dff_sg \buff_mem_reg[13][6]  ( .D(n7013), .CP(clk), .Q(\buff_mem[13][6] ) );
  dff_sg \buff_mem_reg[12][6]  ( .D(n6856), .CP(clk), .Q(\buff_mem[12][6] ) );
  dff_sg \buff_mem_reg[11][6]  ( .D(n7234), .CP(clk), .Q(\buff_mem[11][6] ) );
  dff_sg \buff_mem_reg[10][6]  ( .D(n7215), .CP(clk), .Q(\buff_mem[10][6] ) );
  dff_sg \buff_mem_reg[9][6]  ( .D(n7245), .CP(clk), .Q(\buff_mem[9][6] ) );
  dff_sg \buff_mem_reg[8][6]  ( .D(n7197), .CP(clk), .Q(\buff_mem[8][6] ) );
  dff_sg \buff_mem_reg[7][6]  ( .D(n6942), .CP(clk), .Q(\buff_mem[7][6] ) );
  dff_sg \buff_mem_reg[6][6]  ( .D(n6984), .CP(clk), .Q(\buff_mem[6][6] ) );
  dff_sg \buff_mem_reg[5][6]  ( .D(n6978), .CP(clk), .Q(\buff_mem[5][6] ) );
  dff_sg \buff_mem_reg[4][7]  ( .D(n6945), .CP(clk), .Q(\buff_mem[4][7] ) );
  dff_sg \buff_mem_reg[3][7]  ( .D(n7123), .CP(clk), .Q(\buff_mem[3][7] ) );
  dff_sg \buff_mem_reg[2][7]  ( .D(n7085), .CP(clk), .Q(\buff_mem[2][7] ) );
  dff_sg \buff_mem_reg[1][7]  ( .D(n7096), .CP(clk), .Q(\buff_mem[1][7] ) );
  dff_sg \buff_mem_reg[0][7]  ( .D(n7063), .CP(clk), .Q(\buff_mem[0][7] ) );
  dff_sg \buff_mem_reg[19][7]  ( .D(n7140), .CP(clk), .Q(\buff_mem[19][7] ) );
  dff_sg \buff_mem_reg[18][7]  ( .D(n7151), .CP(clk), .Q(\buff_mem[18][7] ) );
  dff_sg \buff_mem_reg[17][7]  ( .D(n7175), .CP(clk), .Q(\buff_mem[17][7] ) );
  dff_sg \buff_mem_reg[16][7]  ( .D(n6880), .CP(clk), .Q(\buff_mem[16][7] ) );
  dff_sg \buff_mem_reg[15][7]  ( .D(n7038), .CP(clk), .Q(\buff_mem[15][7] ) );
  dff_sg \buff_mem_reg[14][7]  ( .D(n7029), .CP(clk), .Q(\buff_mem[14][7] ) );
  dff_sg \buff_mem_reg[13][7]  ( .D(n6998), .CP(clk), .Q(\buff_mem[13][7] ) );
  dff_sg \buff_mem_reg[12][7]  ( .D(n6862), .CP(clk), .Q(\buff_mem[12][7] ) );
  dff_sg \buff_mem_reg[11][7]  ( .D(n7230), .CP(clk), .Q(\buff_mem[11][7] ) );
  dff_sg \buff_mem_reg[10][7]  ( .D(n7213), .CP(clk), .Q(\buff_mem[10][7] ) );
  dff_sg \buff_mem_reg[9][7]  ( .D(n7249), .CP(clk), .Q(\buff_mem[9][7] ) );
  dff_sg \buff_mem_reg[8][7]  ( .D(n7192), .CP(clk), .Q(\buff_mem[8][7] ) );
  dff_sg \buff_mem_reg[7][7]  ( .D(n6932), .CP(clk), .Q(\buff_mem[7][7] ) );
  dff_sg \buff_mem_reg[6][7]  ( .D(n6986), .CP(clk), .Q(\buff_mem[6][7] ) );
  dff_sg \buff_mem_reg[5][7]  ( .D(n6962), .CP(clk), .Q(\buff_mem[5][7] ) );
  dff_sg \buff_mem_reg[4][8]  ( .D(n6954), .CP(clk), .Q(\buff_mem[4][8] ) );
  dff_sg \buff_mem_reg[3][8]  ( .D(n7121), .CP(clk), .Q(\buff_mem[3][8] ) );
  dff_sg \buff_mem_reg[2][8]  ( .D(n7077), .CP(clk), .Q(\buff_mem[2][8] ) );
  dff_sg \buff_mem_reg[1][8]  ( .D(n7101), .CP(clk), .Q(\buff_mem[1][8] ) );
  dff_sg \buff_mem_reg[0][8]  ( .D(n7071), .CP(clk), .Q(\buff_mem[0][8] ) );
  dff_sg \buff_mem_reg[19][8]  ( .D(n7131), .CP(clk), .Q(\buff_mem[19][8] ) );
  dff_sg \buff_mem_reg[18][8]  ( .D(n7154), .CP(clk), .Q(\buff_mem[18][8] ) );
  dff_sg \buff_mem_reg[17][8]  ( .D(n7167), .CP(clk), .Q(\buff_mem[17][8] ) );
  dff_sg \buff_mem_reg[16][8]  ( .D(n6870), .CP(clk), .Q(\buff_mem[16][8] ) );
  dff_sg \buff_mem_reg[15][8]  ( .D(n7039), .CP(clk), .Q(\buff_mem[15][8] ) );
  dff_sg \buff_mem_reg[14][8]  ( .D(n7026), .CP(clk), .Q(\buff_mem[14][8] ) );
  dff_sg \buff_mem_reg[13][8]  ( .D(n7011), .CP(clk), .Q(\buff_mem[13][8] ) );
  dff_sg \buff_mem_reg[12][8]  ( .D(n6857), .CP(clk), .Q(\buff_mem[12][8] ) );
  dff_sg \buff_mem_reg[11][8]  ( .D(n7221), .CP(clk), .Q(\buff_mem[11][8] ) );
  dff_sg \buff_mem_reg[10][8]  ( .D(n7203), .CP(clk), .Q(\buff_mem[10][8] ) );
  dff_sg \buff_mem_reg[9][8]  ( .D(n7240), .CP(clk), .Q(\buff_mem[9][8] ) );
  dff_sg \buff_mem_reg[8][8]  ( .D(n7185), .CP(clk), .Q(\buff_mem[8][8] ) );
  dff_sg \buff_mem_reg[7][8]  ( .D(n6940), .CP(clk), .Q(\buff_mem[7][8] ) );
  dff_sg \buff_mem_reg[6][8]  ( .D(n6980), .CP(clk), .Q(\buff_mem[6][8] ) );
  dff_sg \buff_mem_reg[5][8]  ( .D(n6976), .CP(clk), .Q(\buff_mem[5][8] ) );
  dff_sg \buff_mem_reg[4][9]  ( .D(n6957), .CP(clk), .Q(\buff_mem[4][9] ) );
  dff_sg \buff_mem_reg[3][9]  ( .D(n7127), .CP(clk), .Q(\buff_mem[3][9] ) );
  dff_sg \buff_mem_reg[2][9]  ( .D(n7090), .CP(clk), .Q(\buff_mem[2][9] ) );
  dff_sg \buff_mem_reg[1][9]  ( .D(n7109), .CP(clk), .Q(\buff_mem[1][9] ) );
  dff_sg \buff_mem_reg[0][9]  ( .D(n7072), .CP(clk), .Q(\buff_mem[0][9] ) );
  dff_sg \buff_mem_reg[19][9]  ( .D(n7135), .CP(clk), .Q(\buff_mem[19][9] ) );
  dff_sg \buff_mem_reg[18][9]  ( .D(n7163), .CP(clk), .Q(\buff_mem[18][9] ) );
  dff_sg \buff_mem_reg[17][9]  ( .D(n7171), .CP(clk), .Q(\buff_mem[17][9] ) );
  dff_sg \buff_mem_reg[16][9]  ( .D(n6874), .CP(clk), .Q(\buff_mem[16][9] ) );
  dff_sg \buff_mem_reg[15][9]  ( .D(n7049), .CP(clk), .Q(\buff_mem[15][9] ) );
  dff_sg \buff_mem_reg[14][9]  ( .D(n7018), .CP(clk), .Q(\buff_mem[14][9] ) );
  dff_sg \buff_mem_reg[13][9]  ( .D(n7015), .CP(clk), .Q(\buff_mem[13][9] ) );
  dff_sg \buff_mem_reg[12][9]  ( .D(n6866), .CP(clk), .Q(\buff_mem[12][9] ) );
  dff_sg \buff_mem_reg[11][9]  ( .D(n7235), .CP(clk), .Q(\buff_mem[11][9] ) );
  dff_sg \buff_mem_reg[10][9]  ( .D(n7218), .CP(clk), .Q(\buff_mem[10][9] ) );
  dff_sg \buff_mem_reg[9][9]  ( .D(n7253), .CP(clk), .Q(\buff_mem[9][9] ) );
  dff_sg \buff_mem_reg[8][9]  ( .D(n7200), .CP(clk), .Q(\buff_mem[8][9] ) );
  dff_sg \buff_mem_reg[7][9]  ( .D(n6941), .CP(clk), .Q(\buff_mem[7][9] ) );
  dff_sg \buff_mem_reg[6][9]  ( .D(n6992), .CP(clk), .Q(\buff_mem[6][9] ) );
  dff_sg \buff_mem_reg[5][9]  ( .D(n6977), .CP(clk), .Q(\buff_mem[5][9] ) );
  dff_sg \buff_mem_reg[4][10]  ( .D(n6950), .CP(clk), .Q(\buff_mem[4][10] ) );
  dff_sg \buff_mem_reg[3][10]  ( .D(n7116), .CP(clk), .Q(\buff_mem[3][10] ) );
  dff_sg \buff_mem_reg[2][10]  ( .D(n7080), .CP(clk), .Q(\buff_mem[2][10] ) );
  dff_sg \buff_mem_reg[1][10]  ( .D(n7095), .CP(clk), .Q(\buff_mem[1][10] ) );
  dff_sg \buff_mem_reg[0][10]  ( .D(n7060), .CP(clk), .Q(\buff_mem[0][10] ) );
  dff_sg \buff_mem_reg[19][10]  ( .D(n7142), .CP(clk), .Q(\buff_mem[19][10] )
         );
  dff_sg \buff_mem_reg[18][10]  ( .D(n7149), .CP(clk), .Q(\buff_mem[18][10] )
         );
  dff_sg \buff_mem_reg[17][10]  ( .D(n7178), .CP(clk), .Q(\buff_mem[17][10] )
         );
  dff_sg \buff_mem_reg[16][10]  ( .D(n6878), .CP(clk), .Q(\buff_mem[16][10] )
         );
  dff_sg \buff_mem_reg[15][10]  ( .D(n7036), .CP(clk), .Q(\buff_mem[15][10] )
         );
  dff_sg \buff_mem_reg[14][10]  ( .D(n7021), .CP(clk), .Q(\buff_mem[14][10] )
         );
  dff_sg \buff_mem_reg[13][10]  ( .D(n7002), .CP(clk), .Q(\buff_mem[13][10] )
         );
  dff_sg \buff_mem_reg[12][10]  ( .D(n6850), .CP(clk), .Q(\buff_mem[12][10] )
         );
  dff_sg \buff_mem_reg[11][10]  ( .D(n7224), .CP(clk), .Q(\buff_mem[11][10] )
         );
  dff_sg \buff_mem_reg[10][10]  ( .D(n7206), .CP(clk), .Q(\buff_mem[10][10] )
         );
  dff_sg \buff_mem_reg[9][10]  ( .D(n7239), .CP(clk), .Q(\buff_mem[9][10] ) );
  dff_sg \buff_mem_reg[8][10]  ( .D(n7188), .CP(clk), .Q(\buff_mem[8][10] ) );
  dff_sg \buff_mem_reg[7][10]  ( .D(n6929), .CP(clk), .Q(\buff_mem[7][10] ) );
  dff_sg \buff_mem_reg[6][10]  ( .D(n6988), .CP(clk), .Q(\buff_mem[6][10] ) );
  dff_sg \buff_mem_reg[5][10]  ( .D(n6966), .CP(clk), .Q(\buff_mem[5][10] ) );
  dff_sg \buff_mem_reg[4][11]  ( .D(n6925), .CP(clk), .Q(\buff_mem[4][11] ) );
  dff_sg \buff_mem_reg[3][11]  ( .D(n6920), .CP(clk), .Q(\buff_mem[3][11] ) );
  dff_sg \buff_mem_reg[2][11]  ( .D(n6912), .CP(clk), .Q(\buff_mem[2][11] ) );
  dff_sg \buff_mem_reg[1][11]  ( .D(n6917), .CP(clk), .Q(\buff_mem[1][11] ) );
  dff_sg \buff_mem_reg[0][11]  ( .D(n6924), .CP(clk), .Q(\buff_mem[0][11] ) );
  dff_sg \buff_mem_reg[19][11]  ( .D(n6913), .CP(clk), .Q(\buff_mem[19][11] )
         );
  dff_sg \buff_mem_reg[18][11]  ( .D(n6908), .CP(clk), .Q(\buff_mem[18][11] )
         );
  dff_sg \buff_mem_reg[17][11]  ( .D(n6911), .CP(clk), .Q(\buff_mem[17][11] )
         );
  dff_sg \buff_mem_reg[16][11]  ( .D(n6879), .CP(clk), .Q(\buff_mem[16][11] )
         );
  dff_sg \buff_mem_reg[15][11]  ( .D(n6914), .CP(clk), .Q(\buff_mem[15][11] )
         );
  dff_sg \buff_mem_reg[14][11]  ( .D(n6909), .CP(clk), .Q(\buff_mem[14][11] )
         );
  dff_sg \buff_mem_reg[13][11]  ( .D(n6916), .CP(clk), .Q(\buff_mem[13][11] )
         );
  dff_sg \buff_mem_reg[12][11]  ( .D(n6853), .CP(clk), .Q(\buff_mem[12][11] )
         );
  dff_sg \buff_mem_reg[11][11]  ( .D(n6915), .CP(clk), .Q(\buff_mem[11][11] )
         );
  dff_sg \buff_mem_reg[10][11]  ( .D(n6919), .CP(clk), .Q(\buff_mem[10][11] )
         );
  dff_sg \buff_mem_reg[9][11]  ( .D(n6922), .CP(clk), .Q(\buff_mem[9][11] ) );
  dff_sg \buff_mem_reg[8][11]  ( .D(n6921), .CP(clk), .Q(\buff_mem[8][11] ) );
  dff_sg \buff_mem_reg[7][11]  ( .D(n6918), .CP(clk), .Q(\buff_mem[7][11] ) );
  dff_sg \buff_mem_reg[6][11]  ( .D(n6910), .CP(clk), .Q(\buff_mem[6][11] ) );
  dff_sg \buff_mem_reg[5][11]  ( .D(n6923), .CP(clk), .Q(\buff_mem[5][11] ) );
  dff_sg empty_reg ( .D(n6907), .CP(clk), .Q(n8262) );
  dff_sg \rd_ptr_reg[4]  ( .D(n7255), .CP(clk), .Q(rd_ptr[4]) );
  dff_sg \rd_ptr_reg[1]  ( .D(n7256), .CP(clk), .Q(rd_ptr[1]) );
  dff_sg \rd_ptr_reg[2]  ( .D(n7259), .CP(clk), .Q(rd_ptr[2]) );
  dff_sg \rd_ptr_reg[3]  ( .D(n7258), .CP(clk), .Q(rd_ptr[3]) );
  dff_sg \data_out_reg[19]  ( .D(N161), .CP(clk), .Q(data_out[19]) );
  dff_sg \data_out_reg[18]  ( .D(N160), .CP(clk), .Q(data_out[18]) );
  dff_sg \data_out_reg[17]  ( .D(N159), .CP(clk), .Q(data_out[17]) );
  dff_sg \data_out_reg[16]  ( .D(N158), .CP(clk), .Q(data_out[16]) );
  dff_sg \data_out_reg[15]  ( .D(N157), .CP(clk), .Q(data_out[15]) );
  dff_sg \data_out_reg[14]  ( .D(N156), .CP(clk), .Q(data_out[14]) );
  dff_sg \data_out_reg[13]  ( .D(N155), .CP(clk), .Q(data_out[13]) );
  dff_sg \data_out_reg[12]  ( .D(N154), .CP(clk), .Q(data_out[12]) );
  dff_sg \data_out_reg[11]  ( .D(N153), .CP(clk), .Q(data_out[11]) );
  dff_sg \data_out_reg[10]  ( .D(N152), .CP(clk), .Q(data_out[10]) );
  dff_sg \data_out_reg[9]  ( .D(N151), .CP(clk), .Q(data_out[9]) );
  dff_sg \data_out_reg[8]  ( .D(N150), .CP(clk), .Q(data_out[8]) );
  dff_sg \data_out_reg[7]  ( .D(N149), .CP(clk), .Q(data_out[7]) );
  dff_sg \data_out_reg[6]  ( .D(N148), .CP(clk), .Q(data_out[6]) );
  dff_sg \data_out_reg[5]  ( .D(N147), .CP(clk), .Q(data_out[5]) );
  dff_sg \data_out_reg[4]  ( .D(N146), .CP(clk), .Q(data_out[4]) );
  dff_sg \data_out_reg[3]  ( .D(N145), .CP(clk), .Q(data_out[3]) );
  dff_sg \data_out_reg[2]  ( .D(N144), .CP(clk), .Q(data_out[2]) );
  dff_sg \data_out_reg[1]  ( .D(N143), .CP(clk), .Q(data_out[1]) );
  dff_sg \data_out_reg[0]  ( .D(N142), .CP(clk), .Q(data_out[0]) );
  nand_x8_sg U3223 ( .A(n5120), .B(n5121), .X(n5081) );
  nand_x8_sg U3284 ( .A(n5120), .B(n5163), .X(n5124) );
  nand_x8_sg U3498 ( .A(n5350), .B(n5351), .X(n5236) );
  nand_x8_sg U3553 ( .A(n5120), .B(n5351), .X(n5221) );
  nand_x8_sg U3608 ( .A(n5424), .B(n5351), .X(n5197) );
  nand_x8_sg U3663 ( .A(n5461), .B(n5351), .X(n5246) );
  nand_x8_sg U3664 ( .A(n5462), .B(n4887), .X(n5351) );
  nand_x8_sg U3721 ( .A(n5424), .B(n5121), .X(n5206) );
  nand_x8_sg U3776 ( .A(n5461), .B(n5121), .X(n5227) );
  nand_x8_sg U3831 ( .A(n5350), .B(n5121), .X(n5194) );
  nand_x8_sg U3832 ( .A(n5573), .B(n4887), .X(n5121) );
  nand_x8_sg U3915 ( .A(n5120), .B(n5629), .X(n5224) );
  nand_x8_sg U3970 ( .A(n5461), .B(n5629), .X(n5209) );
  nand_x8_sg U4025 ( .A(n5424), .B(n5629), .X(n5215) );
  nand_x8_sg U4080 ( .A(n5350), .B(n5629), .X(n5218) );
  nand_x8_sg U4081 ( .A(n5738), .B(n4887), .X(n5629) );
  nand_x8_sg U4137 ( .A(n5350), .B(n5163), .X(n5212) );
  nand_x8_sg U4192 ( .A(n5461), .B(n5163), .X(n5203) );
  nand_x8_sg U4247 ( .A(n5424), .B(n5163), .X(n5230) );
  nand_x8_sg U4248 ( .A(n5848), .B(n4887), .X(n5163) );
  nand_x8_sg U4306 ( .A(n5120), .B(n5887), .X(n5200) );
  nand_x8_sg U4307 ( .A(n5580), .B(n4887), .X(n5120) );
  nand_x8_sg U4363 ( .A(n5461), .B(n5887), .X(n5233) );
  nand_x8_sg U4364 ( .A(n5924), .B(n4887), .X(n5461) );
  nand_x8_sg U4420 ( .A(n5350), .B(n5887), .X(n5239) );
  nand_x8_sg U4421 ( .A(n5579), .B(n4887), .X(n5350) );
  nand_x8_sg U4422 ( .A(n7282), .B(n7331), .X(n5579) );
  nand_x8_sg U4495 ( .A(n5424), .B(n5887), .X(n5242) );
  nand_x8_sg U4496 ( .A(n6015), .B(n4887), .X(n5887) );
  nand_x8_sg U4499 ( .A(n8259), .B(n4911), .X(n5464) );
  nand_x8_sg U4504 ( .A(n6020), .B(n4887), .X(n5424) );
  nor_x2_sg U4534 ( .A(n6040), .B(n6041), .X(n6039) );
  nor_x2_sg U4543 ( .A(n4968), .B(n8210), .X(n6054) );
  nor_x2_sg U4544 ( .A(n4969), .B(n8208), .X(n6053) );
  nor_x2_sg U4552 ( .A(n4974), .B(n8201), .X(n6067) );
  nor_x2_sg U4553 ( .A(n4975), .B(n8199), .X(n6066) );
  nor_x2_sg U4562 ( .A(n4973), .B(n6083), .X(n6082) );
  nor_x2_sg U4563 ( .A(n4971), .B(n8190), .X(n6081) );
  nor_x2_sg U4571 ( .A(n4972), .B(n6096), .X(n6095) );
  nor_x2_sg U4572 ( .A(n4970), .B(n8168), .X(n6094) );
  nor_x2_sg U4574 ( .A(n6099), .B(n6100), .X(n6098) );
  nor_x2_sg U4583 ( .A(n4960), .B(n8209), .X(n6110) );
  nor_x2_sg U4584 ( .A(n4961), .B(n8207), .X(n6109) );
  nor_x2_sg U4592 ( .A(n4966), .B(n8200), .X(n6118) );
  nor_x2_sg U4593 ( .A(n4967), .B(n8198), .X(n6117) );
  nor_x2_sg U4602 ( .A(n4965), .B(n8191), .X(n6128) );
  nor_x2_sg U4603 ( .A(n4963), .B(n8189), .X(n6127) );
  nor_x2_sg U4611 ( .A(n4964), .B(n8169), .X(n6136) );
  nor_x2_sg U4612 ( .A(n4962), .B(n8167), .X(n6135) );
  nor_x2_sg U4614 ( .A(n6138), .B(n6139), .X(n6137) );
  nor_x2_sg U4623 ( .A(n4952), .B(n6055), .X(n6149) );
  nor_x2_sg U4624 ( .A(n4953), .B(n6056), .X(n6148) );
  nor_x2_sg U4632 ( .A(n4958), .B(n6068), .X(n6157) );
  nor_x2_sg U4633 ( .A(n4959), .B(n6069), .X(n6156) );
  nor_x2_sg U4642 ( .A(n4957), .B(n6083), .X(n6167) );
  nor_x2_sg U4643 ( .A(n4955), .B(n6084), .X(n6166) );
  nor_x2_sg U4651 ( .A(n4956), .B(n6096), .X(n6175) );
  nor_x2_sg U4652 ( .A(n4954), .B(n6097), .X(n6174) );
  nor_x2_sg U4654 ( .A(n6177), .B(n6178), .X(n6176) );
  nor_x2_sg U4663 ( .A(n4944), .B(n8210), .X(n6188) );
  nor_x2_sg U4664 ( .A(n4945), .B(n8208), .X(n6187) );
  nor_x2_sg U4672 ( .A(n4950), .B(n8201), .X(n6196) );
  nor_x2_sg U4673 ( .A(n4951), .B(n8199), .X(n6195) );
  nor_x2_sg U4682 ( .A(n4949), .B(n8191), .X(n6206) );
  nor_x2_sg U4683 ( .A(n4947), .B(n8190), .X(n6205) );
  nor_x2_sg U4691 ( .A(n4948), .B(n8169), .X(n6214) );
  nor_x2_sg U4692 ( .A(n4946), .B(n8168), .X(n6213) );
  nor_x2_sg U4694 ( .A(n6216), .B(n6217), .X(n6215) );
  nor_x2_sg U4703 ( .A(n4936), .B(n8209), .X(n6227) );
  nor_x2_sg U4704 ( .A(n4937), .B(n8207), .X(n6226) );
  nor_x2_sg U4712 ( .A(n4942), .B(n8200), .X(n6235) );
  nor_x2_sg U4713 ( .A(n4943), .B(n8198), .X(n6234) );
  nor_x2_sg U4722 ( .A(n4941), .B(n6083), .X(n6245) );
  nor_x2_sg U4723 ( .A(n4939), .B(n8189), .X(n6244) );
  nor_x2_sg U4731 ( .A(n4940), .B(n6096), .X(n6253) );
  nor_x2_sg U4732 ( .A(n4938), .B(n8167), .X(n6252) );
  nor_x2_sg U4734 ( .A(n6255), .B(n6256), .X(n6254) );
  nor_x2_sg U4743 ( .A(n4928), .B(n6055), .X(n6266) );
  nor_x2_sg U4744 ( .A(n4929), .B(n6056), .X(n6265) );
  nor_x2_sg U4752 ( .A(n4934), .B(n6068), .X(n6274) );
  nor_x2_sg U4753 ( .A(n4935), .B(n6069), .X(n6273) );
  nor_x2_sg U4762 ( .A(n4933), .B(n8191), .X(n6284) );
  nor_x2_sg U4763 ( .A(n4931), .B(n6084), .X(n6283) );
  nor_x2_sg U4771 ( .A(n4932), .B(n8169), .X(n6292) );
  nor_x2_sg U4772 ( .A(n4930), .B(n6097), .X(n6291) );
  nor_x2_sg U4774 ( .A(n6294), .B(n6295), .X(n6293) );
  nor_x2_sg U4783 ( .A(n4920), .B(n8210), .X(n6305) );
  nor_x2_sg U4784 ( .A(n4921), .B(n8208), .X(n6304) );
  nor_x2_sg U4792 ( .A(n4926), .B(n8201), .X(n6313) );
  nor_x2_sg U4793 ( .A(n4927), .B(n8199), .X(n6312) );
  nor_x2_sg U4802 ( .A(n4925), .B(n6083), .X(n6323) );
  nor_x2_sg U4803 ( .A(n4923), .B(n8190), .X(n6322) );
  nor_x2_sg U4811 ( .A(n4924), .B(n6096), .X(n6331) );
  nor_x2_sg U4812 ( .A(n4922), .B(n8168), .X(n6330) );
  nor_x2_sg U4814 ( .A(n6333), .B(n6334), .X(n6332) );
  nor_x2_sg U4823 ( .A(n4912), .B(n8209), .X(n6344) );
  nor_x2_sg U4824 ( .A(n4913), .B(n8207), .X(n6343) );
  nor_x2_sg U4832 ( .A(n4918), .B(n8200), .X(n6352) );
  nor_x2_sg U4833 ( .A(n4919), .B(n8198), .X(n6351) );
  nor_x2_sg U4842 ( .A(n4917), .B(n8191), .X(n6362) );
  nor_x2_sg U4843 ( .A(n4915), .B(n8189), .X(n6361) );
  nor_x2_sg U4851 ( .A(n4916), .B(n8169), .X(n6370) );
  nor_x2_sg U4852 ( .A(n4914), .B(n8167), .X(n6369) );
  nor_x2_sg U4854 ( .A(n6372), .B(n6373), .X(n6371) );
  nor_x2_sg U4863 ( .A(n5064), .B(n6055), .X(n6383) );
  nor_x2_sg U4864 ( .A(n5065), .B(n6056), .X(n6382) );
  nor_x2_sg U4872 ( .A(n5070), .B(n6068), .X(n6391) );
  nor_x2_sg U4873 ( .A(n5071), .B(n6069), .X(n6390) );
  nor_x2_sg U4882 ( .A(n5069), .B(n6083), .X(n6401) );
  nor_x2_sg U4883 ( .A(n5067), .B(n6084), .X(n6400) );
  nor_x2_sg U4891 ( .A(n5068), .B(n6096), .X(n6409) );
  nor_x2_sg U4892 ( .A(n5066), .B(n6097), .X(n6408) );
  nor_x2_sg U4894 ( .A(n6411), .B(n6412), .X(n6410) );
  nor_x2_sg U4903 ( .A(n5056), .B(n8210), .X(n6422) );
  nor_x2_sg U4904 ( .A(n5057), .B(n8208), .X(n6421) );
  nor_x2_sg U4912 ( .A(n5062), .B(n8201), .X(n6430) );
  nor_x2_sg U4913 ( .A(n5063), .B(n8199), .X(n6429) );
  nor_x2_sg U4922 ( .A(n5061), .B(n8191), .X(n6440) );
  nor_x2_sg U4923 ( .A(n5059), .B(n8190), .X(n6439) );
  nor_x2_sg U4931 ( .A(n5060), .B(n8169), .X(n6448) );
  nor_x2_sg U4932 ( .A(n5058), .B(n8168), .X(n6447) );
  nor_x2_sg U4934 ( .A(n6450), .B(n6451), .X(n6449) );
  nor_x2_sg U4943 ( .A(n5048), .B(n8209), .X(n6461) );
  nor_x2_sg U4944 ( .A(n5049), .B(n8207), .X(n6460) );
  nor_x2_sg U4952 ( .A(n5054), .B(n8200), .X(n6469) );
  nor_x2_sg U4953 ( .A(n5055), .B(n8198), .X(n6468) );
  nor_x2_sg U4962 ( .A(n5053), .B(n6083), .X(n6479) );
  nor_x2_sg U4963 ( .A(n5051), .B(n8189), .X(n6478) );
  nor_x2_sg U4971 ( .A(n5052), .B(n6096), .X(n6487) );
  nor_x2_sg U4972 ( .A(n5050), .B(n8167), .X(n6486) );
  nor_x2_sg U4974 ( .A(n6489), .B(n6490), .X(n6488) );
  nor_x2_sg U4983 ( .A(n5040), .B(n6055), .X(n6500) );
  nor_x2_sg U4984 ( .A(n5041), .B(n6056), .X(n6499) );
  nor_x2_sg U4992 ( .A(n5046), .B(n6068), .X(n6508) );
  nor_x2_sg U4993 ( .A(n5047), .B(n6069), .X(n6507) );
  nor_x2_sg U5002 ( .A(n5045), .B(n8191), .X(n6518) );
  nor_x2_sg U5003 ( .A(n5043), .B(n6084), .X(n6517) );
  nor_x2_sg U5011 ( .A(n5044), .B(n8169), .X(n6526) );
  nor_x2_sg U5012 ( .A(n5042), .B(n6097), .X(n6525) );
  nor_x2_sg U5014 ( .A(n6528), .B(n6529), .X(n6527) );
  nor_x2_sg U5023 ( .A(n5032), .B(n8210), .X(n6539) );
  nor_x2_sg U5024 ( .A(n5033), .B(n8208), .X(n6538) );
  nor_x2_sg U5032 ( .A(n5038), .B(n8201), .X(n6547) );
  nor_x2_sg U5033 ( .A(n5039), .B(n8199), .X(n6546) );
  nor_x2_sg U5042 ( .A(n5037), .B(n6083), .X(n6557) );
  nor_x2_sg U5043 ( .A(n5035), .B(n8190), .X(n6556) );
  nor_x2_sg U5051 ( .A(n5036), .B(n6096), .X(n6565) );
  nor_x2_sg U5052 ( .A(n5034), .B(n8168), .X(n6564) );
  nor_x2_sg U5054 ( .A(n6567), .B(n6568), .X(n6566) );
  nor_x2_sg U5063 ( .A(n5024), .B(n8209), .X(n6578) );
  nor_x2_sg U5064 ( .A(n5025), .B(n8207), .X(n6577) );
  nor_x2_sg U5072 ( .A(n5030), .B(n8200), .X(n6586) );
  nor_x2_sg U5073 ( .A(n5031), .B(n8198), .X(n6585) );
  nor_x2_sg U5082 ( .A(n5029), .B(n8191), .X(n6596) );
  nor_x2_sg U5083 ( .A(n5027), .B(n8189), .X(n6595) );
  nor_x2_sg U5091 ( .A(n5028), .B(n8169), .X(n6604) );
  nor_x2_sg U5092 ( .A(n5026), .B(n8167), .X(n6603) );
  nor_x2_sg U5094 ( .A(n6606), .B(n6607), .X(n6605) );
  nor_x2_sg U5103 ( .A(n5016), .B(n6055), .X(n6617) );
  nor_x2_sg U5104 ( .A(n5017), .B(n6056), .X(n6616) );
  nor_x2_sg U5112 ( .A(n5022), .B(n6068), .X(n6625) );
  nor_x2_sg U5113 ( .A(n5023), .B(n6069), .X(n6624) );
  nor_x2_sg U5122 ( .A(n5021), .B(n6083), .X(n6635) );
  nor_x2_sg U5123 ( .A(n5019), .B(n6084), .X(n6634) );
  nor_x2_sg U5131 ( .A(n5020), .B(n6096), .X(n6643) );
  nor_x2_sg U5132 ( .A(n5018), .B(n6097), .X(n6642) );
  nor_x2_sg U5134 ( .A(n6645), .B(n6646), .X(n6644) );
  nor_x2_sg U5143 ( .A(n5008), .B(n8210), .X(n6656) );
  nor_x2_sg U5144 ( .A(n5009), .B(n8208), .X(n6655) );
  nor_x2_sg U5152 ( .A(n5014), .B(n8201), .X(n6664) );
  nor_x2_sg U5153 ( .A(n5015), .B(n8199), .X(n6663) );
  nor_x2_sg U5162 ( .A(n5013), .B(n8191), .X(n6674) );
  nor_x2_sg U5163 ( .A(n5011), .B(n8190), .X(n6673) );
  nor_x2_sg U5171 ( .A(n5012), .B(n8169), .X(n6682) );
  nor_x2_sg U5172 ( .A(n5010), .B(n8168), .X(n6681) );
  nor_x2_sg U5174 ( .A(n6684), .B(n6685), .X(n6683) );
  nor_x2_sg U5183 ( .A(n5000), .B(n8209), .X(n6695) );
  nor_x2_sg U5184 ( .A(n5001), .B(n8207), .X(n6694) );
  nor_x2_sg U5192 ( .A(n5006), .B(n8200), .X(n6703) );
  nor_x2_sg U5193 ( .A(n5007), .B(n8198), .X(n6702) );
  nor_x2_sg U5202 ( .A(n5005), .B(n6083), .X(n6713) );
  nor_x2_sg U5203 ( .A(n5003), .B(n8189), .X(n6712) );
  nor_x2_sg U5211 ( .A(n5004), .B(n6096), .X(n6721) );
  nor_x2_sg U5212 ( .A(n5002), .B(n8167), .X(n6720) );
  nor_x2_sg U5214 ( .A(n6723), .B(n6724), .X(n6722) );
  nor_x2_sg U5223 ( .A(n4992), .B(n6055), .X(n6734) );
  nor_x2_sg U5224 ( .A(n4993), .B(n6056), .X(n6733) );
  nor_x2_sg U5232 ( .A(n4998), .B(n6068), .X(n6742) );
  nor_x2_sg U5233 ( .A(n4999), .B(n6069), .X(n6741) );
  nor_x2_sg U5242 ( .A(n4997), .B(n8191), .X(n6752) );
  nor_x2_sg U5243 ( .A(n4995), .B(n6084), .X(n6751) );
  nor_x2_sg U5251 ( .A(n4996), .B(n8169), .X(n6760) );
  nor_x2_sg U5252 ( .A(n4994), .B(n6097), .X(n6759) );
  nor_x2_sg U5254 ( .A(n6762), .B(n6763), .X(n6761) );
  nor_x2_sg U5263 ( .A(n4984), .B(n8210), .X(n6773) );
  nor_x2_sg U5264 ( .A(n4985), .B(n8208), .X(n6772) );
  nor_x2_sg U5272 ( .A(n4990), .B(n8201), .X(n6781) );
  nor_x2_sg U5273 ( .A(n4991), .B(n8199), .X(n6780) );
  nor_x2_sg U5282 ( .A(n4989), .B(n6083), .X(n6791) );
  nor_x2_sg U5283 ( .A(n4987), .B(n8190), .X(n6790) );
  nor_x2_sg U5291 ( .A(n4988), .B(n6096), .X(n6799) );
  nor_x2_sg U5292 ( .A(n4986), .B(n8168), .X(n6798) );
  nand_x8_sg U5294 ( .A(n6801), .B(rd_en), .X(n6038) );
  nor_x2_sg U5296 ( .A(n6802), .B(n6803), .X(n6800) );
  nor_x2_sg U5308 ( .A(n4976), .B(n8209), .X(n6817) );
  nand_x8_sg U5309 ( .A(n6815), .B(n4897), .X(n6055) );
  nor_x2_sg U5312 ( .A(n4977), .B(n8207), .X(n6816) );
  nand_x8_sg U5313 ( .A(n4899), .B(n7340), .X(n6056) );
  nor_x2_sg U5324 ( .A(n4982), .B(n8200), .X(n6827) );
  nand_x8_sg U5325 ( .A(n6828), .B(n4891), .X(n6068) );
  nor_x2_sg U5326 ( .A(n4983), .B(n8198), .X(n6826) );
  nand_x8_sg U5327 ( .A(n4899), .B(n6828), .X(n6069) );
  nand_x8_sg U5335 ( .A(n7334), .B(n5078), .X(n6823) );
  nor_x2_sg U5340 ( .A(n4981), .B(n8191), .X(n6838) );
  nand_x8_sg U5341 ( .A(n4898), .B(n6828), .X(n6083) );
  nor_x2_sg U5342 ( .A(n4979), .B(n8189), .X(n6837) );
  nand_x8_sg U5343 ( .A(n4891), .B(n6839), .X(n6084) );
  nand_x8_sg U5348 ( .A(n7284), .B(n7327), .X(n6811) );
  nand_x8_sg U5354 ( .A(n7284), .B(n7300), .X(n6037) );
  nor_x2_sg U5357 ( .A(n4980), .B(n8169), .X(n6847) );
  nand_x8_sg U5358 ( .A(n4899), .B(n6839), .X(n6096) );
  nand_x8_sg U5359 ( .A(n7327), .B(n4900), .X(n6810) );
  nor_x2_sg U5360 ( .A(n4978), .B(n8167), .X(n6846) );
  nand_x8_sg U5361 ( .A(n4898), .B(n6839), .X(n6097) );
  nand_x8_sg U5363 ( .A(n7300), .B(n4900), .X(n6814) );
  inv_x2_sg U5365 ( .A(n5249), .X(n4843) );
  inv_x2_sg U5411 ( .A(rd_en), .X(n4889) );
  inv_x2_sg U5412 ( .A(wr_en), .X(n4890) );
  inv_x2_sg U5414 ( .A(n5273), .X(n4892) );
  inv_x2_sg U5415 ( .A(n5276), .X(n4893) );
  inv_x2_sg U5416 ( .A(n5270), .X(n4894) );
  inv_x2_sg U5417 ( .A(n5261), .X(n4895) );
  inv_x2_sg U5418 ( .A(n5258), .X(n4896) );
  inv_x2_sg U5425 ( .A(n5188), .X(n4903) );
  inv_x2_sg U5426 ( .A(n5586), .X(n4904) );
  inv_x2_sg U5428 ( .A(n5191), .X(n4906) );
  inv_x2_sg U5429 ( .A(n5588), .X(n4907) );
  inv_x2_sg U5432 ( .A(n8106), .X(n4910) );
  inv_x2_sg U5434 ( .A(n8022), .X(n4912) );
  inv_x2_sg U5435 ( .A(n7942), .X(n4913) );
  inv_x2_sg U5436 ( .A(n7944), .X(n4914) );
  inv_x2_sg U5437 ( .A(n7862), .X(n4915) );
  inv_x2_sg U5438 ( .A(n8024), .X(n4916) );
  inv_x2_sg U5439 ( .A(n7782), .X(n4917) );
  inv_x2_sg U5440 ( .A(n7864), .X(n4918) );
  inv_x2_sg U5441 ( .A(n7784), .X(n4919) );
  inv_x2_sg U5442 ( .A(n8026), .X(n4920) );
  inv_x2_sg U5443 ( .A(n7946), .X(n4921) );
  inv_x2_sg U5444 ( .A(n7948), .X(n4922) );
  inv_x2_sg U5445 ( .A(n7866), .X(n4923) );
  inv_x2_sg U5446 ( .A(n8028), .X(n4924) );
  inv_x2_sg U5447 ( .A(n7786), .X(n4925) );
  inv_x2_sg U5448 ( .A(n7868), .X(n4926) );
  inv_x2_sg U5449 ( .A(n7788), .X(n4927) );
  inv_x2_sg U5450 ( .A(n8030), .X(n4928) );
  inv_x2_sg U5451 ( .A(n7950), .X(n4929) );
  inv_x2_sg U5452 ( .A(n7952), .X(n4930) );
  inv_x2_sg U5453 ( .A(n7870), .X(n4931) );
  inv_x2_sg U5454 ( .A(n8032), .X(n4932) );
  inv_x2_sg U5455 ( .A(n7790), .X(n4933) );
  inv_x2_sg U5456 ( .A(n7872), .X(n4934) );
  inv_x2_sg U5457 ( .A(n7792), .X(n4935) );
  inv_x2_sg U5458 ( .A(n8034), .X(n4936) );
  inv_x2_sg U5459 ( .A(n7954), .X(n4937) );
  inv_x2_sg U5460 ( .A(n7956), .X(n4938) );
  inv_x2_sg U5461 ( .A(n7874), .X(n4939) );
  inv_x2_sg U5462 ( .A(n8036), .X(n4940) );
  inv_x2_sg U5463 ( .A(n7794), .X(n4941) );
  inv_x2_sg U5464 ( .A(n7876), .X(n4942) );
  inv_x2_sg U5465 ( .A(n7796), .X(n4943) );
  inv_x2_sg U5466 ( .A(n8038), .X(n4944) );
  inv_x2_sg U5467 ( .A(n7958), .X(n4945) );
  inv_x2_sg U5468 ( .A(n7960), .X(n4946) );
  inv_x2_sg U5469 ( .A(n7878), .X(n4947) );
  inv_x2_sg U5470 ( .A(n8040), .X(n4948) );
  inv_x2_sg U5471 ( .A(n7798), .X(n4949) );
  inv_x2_sg U5472 ( .A(n7880), .X(n4950) );
  inv_x2_sg U5473 ( .A(n7800), .X(n4951) );
  inv_x2_sg U5474 ( .A(n8042), .X(n4952) );
  inv_x2_sg U5475 ( .A(n7962), .X(n4953) );
  inv_x2_sg U5476 ( .A(n7964), .X(n4954) );
  inv_x2_sg U5477 ( .A(n7882), .X(n4955) );
  inv_x2_sg U5478 ( .A(n8044), .X(n4956) );
  inv_x2_sg U5479 ( .A(n7802), .X(n4957) );
  inv_x2_sg U5480 ( .A(n7884), .X(n4958) );
  inv_x2_sg U5481 ( .A(n7804), .X(n4959) );
  inv_x2_sg U5482 ( .A(n8046), .X(n4960) );
  inv_x2_sg U5483 ( .A(n7966), .X(n4961) );
  inv_x2_sg U5484 ( .A(n7968), .X(n4962) );
  inv_x2_sg U5485 ( .A(n7886), .X(n4963) );
  inv_x2_sg U5486 ( .A(n8048), .X(n4964) );
  inv_x2_sg U5487 ( .A(n7806), .X(n4965) );
  inv_x2_sg U5488 ( .A(n7888), .X(n4966) );
  inv_x2_sg U5489 ( .A(n7808), .X(n4967) );
  inv_x2_sg U5490 ( .A(n8050), .X(n4968) );
  inv_x2_sg U5491 ( .A(n7970), .X(n4969) );
  inv_x2_sg U5492 ( .A(n7972), .X(n4970) );
  inv_x2_sg U5493 ( .A(n7890), .X(n4971) );
  inv_x2_sg U5494 ( .A(n8052), .X(n4972) );
  inv_x2_sg U5495 ( .A(n7810), .X(n4973) );
  inv_x2_sg U5496 ( .A(n7892), .X(n4974) );
  inv_x2_sg U5497 ( .A(n7812), .X(n4975) );
  inv_x2_sg U5498 ( .A(n8054), .X(n4976) );
  inv_x2_sg U5499 ( .A(n7974), .X(n4977) );
  inv_x2_sg U5500 ( .A(n7976), .X(n4978) );
  inv_x2_sg U5501 ( .A(n7894), .X(n4979) );
  inv_x2_sg U5502 ( .A(n8056), .X(n4980) );
  inv_x2_sg U5503 ( .A(n7814), .X(n4981) );
  inv_x2_sg U5504 ( .A(n7896), .X(n4982) );
  inv_x2_sg U5505 ( .A(n7816), .X(n4983) );
  inv_x2_sg U5506 ( .A(n8058), .X(n4984) );
  inv_x2_sg U5507 ( .A(n7978), .X(n4985) );
  inv_x2_sg U5508 ( .A(n7980), .X(n4986) );
  inv_x2_sg U5509 ( .A(n7898), .X(n4987) );
  inv_x2_sg U5510 ( .A(n8060), .X(n4988) );
  inv_x2_sg U5511 ( .A(n7818), .X(n4989) );
  inv_x2_sg U5512 ( .A(n7900), .X(n4990) );
  inv_x2_sg U5513 ( .A(n7820), .X(n4991) );
  inv_x2_sg U5514 ( .A(n8062), .X(n4992) );
  inv_x2_sg U5515 ( .A(n7982), .X(n4993) );
  inv_x2_sg U5516 ( .A(n7984), .X(n4994) );
  inv_x2_sg U5517 ( .A(n7902), .X(n4995) );
  inv_x2_sg U5518 ( .A(n8064), .X(n4996) );
  inv_x2_sg U5519 ( .A(n7822), .X(n4997) );
  inv_x2_sg U5520 ( .A(n7904), .X(n4998) );
  inv_x2_sg U5521 ( .A(n7824), .X(n4999) );
  inv_x2_sg U5522 ( .A(n8066), .X(n5000) );
  inv_x2_sg U5523 ( .A(n7986), .X(n5001) );
  inv_x2_sg U5524 ( .A(n7988), .X(n5002) );
  inv_x2_sg U5525 ( .A(n7906), .X(n5003) );
  inv_x2_sg U5526 ( .A(n8068), .X(n5004) );
  inv_x2_sg U5527 ( .A(n7826), .X(n5005) );
  inv_x2_sg U5528 ( .A(n7908), .X(n5006) );
  inv_x2_sg U5529 ( .A(n7828), .X(n5007) );
  inv_x2_sg U5530 ( .A(n8070), .X(n5008) );
  inv_x2_sg U5531 ( .A(n7990), .X(n5009) );
  inv_x2_sg U5532 ( .A(n7992), .X(n5010) );
  inv_x2_sg U5533 ( .A(n7910), .X(n5011) );
  inv_x2_sg U5534 ( .A(n8072), .X(n5012) );
  inv_x2_sg U5535 ( .A(n7830), .X(n5013) );
  inv_x2_sg U5536 ( .A(n7912), .X(n5014) );
  inv_x2_sg U5537 ( .A(n7832), .X(n5015) );
  inv_x2_sg U5538 ( .A(n8074), .X(n5016) );
  inv_x2_sg U5539 ( .A(n7994), .X(n5017) );
  inv_x2_sg U5540 ( .A(n7996), .X(n5018) );
  inv_x2_sg U5541 ( .A(n7914), .X(n5019) );
  inv_x2_sg U5542 ( .A(n8076), .X(n5020) );
  inv_x2_sg U5543 ( .A(n7834), .X(n5021) );
  inv_x2_sg U5544 ( .A(n7916), .X(n5022) );
  inv_x2_sg U5545 ( .A(n7836), .X(n5023) );
  inv_x2_sg U5546 ( .A(n8078), .X(n5024) );
  inv_x2_sg U5547 ( .A(n7998), .X(n5025) );
  inv_x2_sg U5548 ( .A(n8000), .X(n5026) );
  inv_x2_sg U5549 ( .A(n7918), .X(n5027) );
  inv_x2_sg U5550 ( .A(n8080), .X(n5028) );
  inv_x2_sg U5551 ( .A(n7838), .X(n5029) );
  inv_x2_sg U5552 ( .A(n7920), .X(n5030) );
  inv_x2_sg U5553 ( .A(n7840), .X(n5031) );
  inv_x2_sg U5554 ( .A(n8082), .X(n5032) );
  inv_x2_sg U5555 ( .A(n8002), .X(n5033) );
  inv_x2_sg U5556 ( .A(n8004), .X(n5034) );
  inv_x2_sg U5557 ( .A(n7922), .X(n5035) );
  inv_x2_sg U5558 ( .A(n8084), .X(n5036) );
  inv_x2_sg U5559 ( .A(n7842), .X(n5037) );
  inv_x2_sg U5560 ( .A(n7924), .X(n5038) );
  inv_x2_sg U5561 ( .A(n7844), .X(n5039) );
  inv_x2_sg U5562 ( .A(n8086), .X(n5040) );
  inv_x2_sg U5563 ( .A(n8006), .X(n5041) );
  inv_x2_sg U5564 ( .A(n8008), .X(n5042) );
  inv_x2_sg U5565 ( .A(n7926), .X(n5043) );
  inv_x2_sg U5566 ( .A(n8088), .X(n5044) );
  inv_x2_sg U5567 ( .A(n7846), .X(n5045) );
  inv_x2_sg U5568 ( .A(n7928), .X(n5046) );
  inv_x2_sg U5569 ( .A(n7848), .X(n5047) );
  inv_x2_sg U5570 ( .A(n8090), .X(n5048) );
  inv_x2_sg U5571 ( .A(n8010), .X(n5049) );
  inv_x2_sg U5572 ( .A(n8012), .X(n5050) );
  inv_x2_sg U5573 ( .A(n7930), .X(n5051) );
  inv_x2_sg U5574 ( .A(n8092), .X(n5052) );
  inv_x2_sg U5575 ( .A(n7850), .X(n5053) );
  inv_x2_sg U5576 ( .A(n7932), .X(n5054) );
  inv_x2_sg U5577 ( .A(n7852), .X(n5055) );
  inv_x2_sg U5578 ( .A(n8094), .X(n5056) );
  inv_x2_sg U5579 ( .A(n8014), .X(n5057) );
  inv_x2_sg U5580 ( .A(n8016), .X(n5058) );
  inv_x2_sg U5581 ( .A(n7934), .X(n5059) );
  inv_x2_sg U5582 ( .A(n8096), .X(n5060) );
  inv_x2_sg U5583 ( .A(n7854), .X(n5061) );
  inv_x2_sg U5584 ( .A(n7936), .X(n5062) );
  inv_x2_sg U5585 ( .A(n7856), .X(n5063) );
  inv_x2_sg U5586 ( .A(n8098), .X(n5064) );
  inv_x2_sg U5587 ( .A(n8018), .X(n5065) );
  inv_x2_sg U5588 ( .A(n8020), .X(n5066) );
  inv_x2_sg U5589 ( .A(n7938), .X(n5067) );
  inv_x2_sg U5590 ( .A(n8100), .X(n5068) );
  inv_x2_sg U5591 ( .A(n7858), .X(n5069) );
  inv_x2_sg U5592 ( .A(n7940), .X(n5070) );
  inv_x2_sg U5593 ( .A(n7860), .X(n5071) );
  inv_x4_sg U5601 ( .A(n6839), .X(n5076) );
  inv_x4_sg U5602 ( .A(n8261), .X(n8260) );
  inv_x4_sg U5603 ( .A(n6077), .X(n8194) );
  inv_x4_sg U5604 ( .A(n4863), .X(n8145) );
  inv_x4_sg U5605 ( .A(n6052), .X(n8211) );
  inv_x4_sg U5606 ( .A(n6049), .X(n8213) );
  inv_x4_sg U5607 ( .A(n4879), .X(n8113) );
  inv_x4_sg U5608 ( .A(n4880), .X(n8111) );
  inv_x4_sg U5609 ( .A(n6048), .X(n8215) );
  inv_x4_sg U5610 ( .A(n4866), .X(n8139) );
  inv_x4_sg U5611 ( .A(n4870), .X(n8131) );
  inv_x4_sg U5612 ( .A(n4871), .X(n8129) );
  inv_x4_sg U5613 ( .A(n4865), .X(n8141) );
  inv_x4_sg U5614 ( .A(n4869), .X(n8133) );
  inv_x4_sg U5615 ( .A(n4868), .X(n8135) );
  inv_x4_sg U5616 ( .A(n4864), .X(n8143) );
  inv_x4_sg U5617 ( .A(n4867), .X(n8137) );
  inv_x4_sg U5618 ( .A(n4876), .X(n8119) );
  inv_x4_sg U5619 ( .A(n4875), .X(n8121) );
  inv_x4_sg U5620 ( .A(n4877), .X(n8117) );
  inv_x4_sg U5621 ( .A(n4874), .X(n8123) );
  inv_x4_sg U5622 ( .A(n4872), .X(n8127) );
  inv_x4_sg U5623 ( .A(n4878), .X(n8115) );
  inv_x4_sg U5624 ( .A(n4873), .X(n8125) );
  inv_x4_sg U5625 ( .A(n4862), .X(n8147) );
  inv_x4_sg U5626 ( .A(n4861), .X(n8149) );
  inv_x4_sg U5627 ( .A(n6089), .X(n8187) );
  inv_x4_sg U5628 ( .A(n6080), .X(n8192) );
  inv_x4_sg U5629 ( .A(n6076), .X(n8196) );
  inv_x4_sg U5630 ( .A(n5850), .X(n8261) );
  inv_x1_sg U5631 ( .A(rd_ptr[3]), .X(n7260) );
  inv_x2_sg U5632 ( .A(n7260), .X(n7261) );
  inv_x1_sg U5633 ( .A(rd_ptr[1]), .X(n7262) );
  inv_x2_sg U5634 ( .A(n7262), .X(n7263) );
  inv_x1_sg U5635 ( .A(rd_ptr[4]), .X(n7264) );
  inv_x2_sg U5636 ( .A(n7264), .X(n7265) );
  inv_x1_sg U5637 ( .A(n8262), .X(n7266) );
  inv_x2_sg U5638 ( .A(n7266), .X(n7267) );
  inv_x1_sg U5639 ( .A(wr_ptr[4]), .X(n7268) );
  inv_x2_sg U5640 ( .A(n7268), .X(n7269) );
  inv_x1_sg U5641 ( .A(wr_ptr[3]), .X(n7270) );
  inv_x2_sg U5642 ( .A(n7270), .X(n7271) );
  inv_x1_sg U5643 ( .A(wr_ptr[2]), .X(n7272) );
  inv_x2_sg U5644 ( .A(n7272), .X(n7273) );
  inv_x1_sg U5645 ( .A(wr_ptr[1]), .X(n7274) );
  inv_x2_sg U5646 ( .A(n7274), .X(n7275) );
  inv_x1_sg U5647 ( .A(wr_ptr[0]), .X(n7276) );
  inv_x2_sg U5648 ( .A(n7276), .X(n7277) );
  inv_x1_sg U5649 ( .A(rd_ptr[0]), .X(n7278) );
  inv_x2_sg U5650 ( .A(n7278), .X(n7279) );
  nor_x4_sg U5651 ( .A(n5072), .B(n6814), .X(n6052) );
  nor_x4_sg U5652 ( .A(n6037), .B(n5073), .X(n6076) );
  nor_x4_sg U5653 ( .A(n5072), .B(n6811), .X(n6049) );
  nor_x4_sg U5654 ( .A(n6814), .B(n5073), .X(n6080) );
  nand_x4_sg U5655 ( .A(n4907), .B(n5583), .X(n5191) );
  nand_x4_sg U5656 ( .A(n4895), .B(n6031), .X(n5276) );
  nand_x2_sg U5657 ( .A(n7282), .B(n4902), .X(n5924) );
  nor_x4_sg U5658 ( .A(n5075), .B(n6037), .X(n6093) );
  inv_x4_sg U5659 ( .A(n6828), .X(n5075) );
  nor_x4_sg U5660 ( .A(n6811), .B(n5073), .X(n6089) );
  nor_x8_sg U5661 ( .A(n6823), .B(n6814), .X(n6062) );
  nor_x2_sg U5662 ( .A(n7300), .B(n5176), .X(n5175) );
  nor_x2_sg U5663 ( .A(n4901), .B(n7327), .X(n5174) );
  inv_x4_sg U5664 ( .A(n5176), .X(n4901) );
  inv_x1_sg U5665 ( .A(n5249), .X(n7280) );
  nand_x4_sg U5666 ( .A(n5250), .B(n5251), .X(n5249) );
  inv_x2_sg U5667 ( .A(rd_ptr[2]), .X(n7335) );
  inv_x1_sg U5668 ( .A(\buff_mem[6][12] ), .X(n7285) );
  inv_x1_sg U5669 ( .A(\buff_mem[6][15] ), .X(n7287) );
  inv_x1_sg U5670 ( .A(\buff_mem[6][18] ), .X(n7289) );
  inv_x1_sg U5671 ( .A(\buff_mem[6][0] ), .X(n7291) );
  inv_x1_sg U5672 ( .A(\buff_mem[6][3] ), .X(n7293) );
  inv_x1_sg U5673 ( .A(\buff_mem[6][6] ), .X(n7295) );
  inv_x1_sg U5674 ( .A(\buff_mem[6][9] ), .X(n7297) );
  nor_x4_sg U5675 ( .A(n5072), .B(n6810), .X(n6048) );
  nor_x8_sg U5676 ( .A(n6823), .B(n6814), .X(n8204) );
  inv_x4_sg U5677 ( .A(n7275), .X(n7281) );
  inv_x8_sg U5678 ( .A(n7281), .X(n7282) );
  inv_x4_sg U5679 ( .A(n7279), .X(n7283) );
  inv_x8_sg U5680 ( .A(n7283), .X(n7284) );
  inv_x8_sg U5681 ( .A(n7284), .X(n4900) );
  nor_x2_sg U5682 ( .A(n4911), .B(n5270), .X(n5268) );
  nor_x2_sg U5683 ( .A(n7329), .B(n4894), .X(n5269) );
  inv_x1_sg U5684 ( .A(\buff_mem[6][13] ), .X(n7301) );
  inv_x1_sg U5685 ( .A(\buff_mem[6][14] ), .X(n7303) );
  inv_x1_sg U5686 ( .A(\buff_mem[6][16] ), .X(n7305) );
  inv_x1_sg U5687 ( .A(\buff_mem[6][17] ), .X(n7307) );
  inv_x1_sg U5688 ( .A(\buff_mem[6][19] ), .X(n7309) );
  inv_x1_sg U5689 ( .A(\buff_mem[6][1] ), .X(n7311) );
  inv_x1_sg U5690 ( .A(\buff_mem[6][2] ), .X(n7313) );
  inv_x1_sg U5691 ( .A(\buff_mem[6][4] ), .X(n7315) );
  inv_x1_sg U5692 ( .A(\buff_mem[6][5] ), .X(n7317) );
  inv_x1_sg U5693 ( .A(\buff_mem[6][7] ), .X(n7319) );
  inv_x1_sg U5694 ( .A(\buff_mem[6][8] ), .X(n7321) );
  inv_x1_sg U5695 ( .A(\buff_mem[6][10] ), .X(n7323) );
  inv_x1_sg U5696 ( .A(\buff_mem[6][11] ), .X(n7325) );
  nor_x4_sg U5697 ( .A(n5579), .B(n4909), .X(n5588) );
  inv_x2_sg U5698 ( .A(n7285), .X(n7286) );
  inv_x2_sg U5699 ( .A(n7287), .X(n7288) );
  inv_x2_sg U5700 ( .A(n7289), .X(n7290) );
  inv_x2_sg U5701 ( .A(n7291), .X(n7292) );
  inv_x2_sg U5702 ( .A(n7293), .X(n7294) );
  inv_x2_sg U5703 ( .A(n7295), .X(n7296) );
  inv_x2_sg U5704 ( .A(n7297), .X(n7298) );
  nand_x8_sg U5705 ( .A(n5073), .B(n5078), .X(n6818) );
  nand_x2_sg U5706 ( .A(n7331), .B(n4908), .X(n6020) );
  nand_x4_sg U5707 ( .A(n4908), .B(n4902), .X(n5580) );
  nor_x2_sg U5708 ( .A(n5259), .B(n4908), .X(n5257) );
  inv_x8_sg U5709 ( .A(n7282), .X(n4908) );
  nor_x8_sg U5710 ( .A(reset), .B(n8259), .X(n5250) );
  inv_x4_sg U5711 ( .A(n7263), .X(n7299) );
  inv_x8_sg U5712 ( .A(n7299), .X(n7300) );
  nor_x4_sg U5713 ( .A(n5076), .B(n6037), .X(n8178) );
  inv_x2_sg U5714 ( .A(n7301), .X(n7302) );
  inv_x2_sg U5715 ( .A(n7303), .X(n7304) );
  inv_x2_sg U5716 ( .A(n7305), .X(n7306) );
  inv_x2_sg U5717 ( .A(n7307), .X(n7308) );
  inv_x2_sg U5718 ( .A(n7309), .X(n7310) );
  inv_x2_sg U5719 ( .A(n7311), .X(n7312) );
  inv_x2_sg U5720 ( .A(n7313), .X(n7314) );
  inv_x2_sg U5721 ( .A(n7315), .X(n7316) );
  inv_x2_sg U5722 ( .A(n7317), .X(n7318) );
  inv_x2_sg U5723 ( .A(n7319), .X(n7320) );
  inv_x2_sg U5724 ( .A(n7321), .X(n7322) );
  inv_x2_sg U5725 ( .A(n7323), .X(n7324) );
  inv_x2_sg U5726 ( .A(n7325), .X(n7326) );
  nor_x4_sg U5727 ( .A(n6032), .B(n5078), .X(n5261) );
  inv_x8_sg U5728 ( .A(n7300), .X(n7327) );
  inv_x8_sg U5729 ( .A(n6815), .X(n5072) );
  nor_x8_sg U5730 ( .A(n6818), .B(n7334), .X(n6815) );
  nor_x8_sg U5731 ( .A(n6823), .B(n6814), .X(n8203) );
  inv_x4_sg U5732 ( .A(n7269), .X(n7328) );
  inv_x8_sg U5733 ( .A(n7328), .X(n7329) );
  inv_x8_sg U5734 ( .A(n7329), .X(n4911) );
  inv_x4_sg U5735 ( .A(n7277), .X(n7330) );
  inv_x8_sg U5736 ( .A(n7330), .X(n7331) );
  inv_x8_sg U5737 ( .A(n6037), .X(n4897) );
  nor_x4_sg U5738 ( .A(n4897), .B(n4899), .X(n5259) );
  nand_x4_sg U5739 ( .A(n4897), .B(n7334), .X(n6032) );
  nand_x1_sg U5740 ( .A(n4893), .B(n4910), .X(n5274) );
  nor_x1_sg U5741 ( .A(n5264), .B(n5265), .X(n5252) );
  inv_x1_sg U5742 ( .A(n5464), .X(n4852) );
  nor_x1_sg U5743 ( .A(n6806), .B(n6807), .X(n6805) );
  nor_x1_sg U5744 ( .A(n6816), .B(n6817), .X(n6812) );
  nor_x1_sg U5745 ( .A(n6819), .B(n6820), .X(n6804) );
  nor_x1_sg U5746 ( .A(n6840), .B(n6841), .X(n6829) );
  nor_x1_sg U5747 ( .A(n6846), .B(n6847), .X(n6844) );
  nor_x1_sg U5748 ( .A(n6831), .B(n6832), .X(n6830) );
  nor_x1_sg U5749 ( .A(n6766), .B(n6767), .X(n6765) );
  nor_x1_sg U5750 ( .A(n6772), .B(n6773), .X(n6770) );
  nor_x1_sg U5751 ( .A(n6774), .B(n6775), .X(n6764) );
  nor_x1_sg U5752 ( .A(n6792), .B(n6793), .X(n6782) );
  nor_x1_sg U5753 ( .A(n6798), .B(n6799), .X(n6796) );
  nor_x1_sg U5754 ( .A(n6784), .B(n6785), .X(n6783) );
  nor_x1_sg U5755 ( .A(n6727), .B(n6728), .X(n6726) );
  nor_x1_sg U5756 ( .A(n6733), .B(n6734), .X(n6731) );
  nor_x1_sg U5757 ( .A(n6735), .B(n6736), .X(n6725) );
  nor_x1_sg U5758 ( .A(n6753), .B(n6754), .X(n6743) );
  nor_x1_sg U5759 ( .A(n6759), .B(n6760), .X(n6757) );
  nor_x1_sg U5760 ( .A(n6745), .B(n6746), .X(n6744) );
  nor_x1_sg U5761 ( .A(n6688), .B(n6689), .X(n6687) );
  nor_x1_sg U5762 ( .A(n6694), .B(n6695), .X(n6692) );
  nor_x1_sg U5763 ( .A(n6696), .B(n6697), .X(n6686) );
  nor_x1_sg U5764 ( .A(n6714), .B(n6715), .X(n6704) );
  nor_x1_sg U5765 ( .A(n6720), .B(n6721), .X(n6718) );
  nor_x1_sg U5766 ( .A(n6706), .B(n6707), .X(n6705) );
  nor_x1_sg U5767 ( .A(n6649), .B(n6650), .X(n6648) );
  nor_x1_sg U5768 ( .A(n6655), .B(n6656), .X(n6653) );
  nor_x1_sg U5769 ( .A(n6657), .B(n6658), .X(n6647) );
  nor_x1_sg U5770 ( .A(n6675), .B(n6676), .X(n6665) );
  nor_x1_sg U5771 ( .A(n6681), .B(n6682), .X(n6679) );
  nor_x1_sg U5772 ( .A(n6667), .B(n6668), .X(n6666) );
  nor_x1_sg U5773 ( .A(n6610), .B(n6611), .X(n6609) );
  nor_x1_sg U5774 ( .A(n6616), .B(n6617), .X(n6614) );
  nor_x1_sg U5775 ( .A(n6618), .B(n6619), .X(n6608) );
  nor_x1_sg U5776 ( .A(n6636), .B(n6637), .X(n6626) );
  nor_x1_sg U5777 ( .A(n6642), .B(n6643), .X(n6640) );
  nor_x1_sg U5778 ( .A(n6628), .B(n6629), .X(n6627) );
  nor_x1_sg U5779 ( .A(n6571), .B(n6572), .X(n6570) );
  nor_x1_sg U5780 ( .A(n6577), .B(n6578), .X(n6575) );
  nor_x1_sg U5781 ( .A(n6579), .B(n6580), .X(n6569) );
  nor_x1_sg U5782 ( .A(n6597), .B(n6598), .X(n6587) );
  nor_x1_sg U5783 ( .A(n6603), .B(n6604), .X(n6601) );
  nor_x1_sg U5784 ( .A(n6589), .B(n6590), .X(n6588) );
  nor_x1_sg U5785 ( .A(n6532), .B(n6533), .X(n6531) );
  nor_x1_sg U5786 ( .A(n6538), .B(n6539), .X(n6536) );
  nor_x1_sg U5787 ( .A(n6540), .B(n6541), .X(n6530) );
  nor_x1_sg U5788 ( .A(n6558), .B(n6559), .X(n6548) );
  nor_x1_sg U5789 ( .A(n6564), .B(n6565), .X(n6562) );
  nor_x1_sg U5790 ( .A(n6550), .B(n6551), .X(n6549) );
  nor_x1_sg U5791 ( .A(n6493), .B(n6494), .X(n6492) );
  nor_x1_sg U5792 ( .A(n6499), .B(n6500), .X(n6497) );
  nor_x1_sg U5793 ( .A(n6501), .B(n6502), .X(n6491) );
  nor_x1_sg U5794 ( .A(n6519), .B(n6520), .X(n6509) );
  nor_x1_sg U5795 ( .A(n6525), .B(n6526), .X(n6523) );
  nor_x1_sg U5796 ( .A(n6511), .B(n6512), .X(n6510) );
  nor_x1_sg U5797 ( .A(n6454), .B(n6455), .X(n6453) );
  nor_x1_sg U5798 ( .A(n6460), .B(n6461), .X(n6458) );
  nor_x1_sg U5799 ( .A(n6462), .B(n6463), .X(n6452) );
  nor_x1_sg U5800 ( .A(n6480), .B(n6481), .X(n6470) );
  nor_x1_sg U5801 ( .A(n6486), .B(n6487), .X(n6484) );
  nor_x1_sg U5802 ( .A(n6472), .B(n6473), .X(n6471) );
  nor_x1_sg U5803 ( .A(n6415), .B(n6416), .X(n6414) );
  nor_x1_sg U5804 ( .A(n6421), .B(n6422), .X(n6419) );
  nor_x1_sg U5805 ( .A(n6423), .B(n6424), .X(n6413) );
  nor_x1_sg U5806 ( .A(n6441), .B(n6442), .X(n6431) );
  nor_x1_sg U5807 ( .A(n6447), .B(n6448), .X(n6445) );
  nor_x1_sg U5808 ( .A(n6433), .B(n6434), .X(n6432) );
  nor_x1_sg U5809 ( .A(n6376), .B(n6377), .X(n6375) );
  nor_x1_sg U5810 ( .A(n6382), .B(n6383), .X(n6380) );
  nor_x1_sg U5811 ( .A(n6384), .B(n6385), .X(n6374) );
  nor_x1_sg U5812 ( .A(n6402), .B(n6403), .X(n6392) );
  nor_x1_sg U5813 ( .A(n6408), .B(n6409), .X(n6406) );
  nor_x1_sg U5814 ( .A(n6394), .B(n6395), .X(n6393) );
  nor_x1_sg U5815 ( .A(n6337), .B(n6338), .X(n6336) );
  nor_x1_sg U5816 ( .A(n6343), .B(n6344), .X(n6341) );
  nor_x1_sg U5817 ( .A(n6345), .B(n6346), .X(n6335) );
  nor_x1_sg U5818 ( .A(n6363), .B(n6364), .X(n6353) );
  nor_x1_sg U5819 ( .A(n6369), .B(n6370), .X(n6367) );
  nor_x1_sg U5820 ( .A(n6355), .B(n6356), .X(n6354) );
  nor_x1_sg U5821 ( .A(n6298), .B(n6299), .X(n6297) );
  nor_x1_sg U5822 ( .A(n6304), .B(n6305), .X(n6302) );
  nor_x1_sg U5823 ( .A(n6306), .B(n6307), .X(n6296) );
  nor_x1_sg U5824 ( .A(n6324), .B(n6325), .X(n6314) );
  nor_x1_sg U5825 ( .A(n6330), .B(n6331), .X(n6328) );
  nor_x1_sg U5826 ( .A(n6316), .B(n6317), .X(n6315) );
  nor_x1_sg U5827 ( .A(n6259), .B(n6260), .X(n6258) );
  nor_x1_sg U5828 ( .A(n6265), .B(n6266), .X(n6263) );
  nor_x1_sg U5829 ( .A(n6267), .B(n6268), .X(n6257) );
  nor_x1_sg U5830 ( .A(n6285), .B(n6286), .X(n6275) );
  nor_x1_sg U5831 ( .A(n6291), .B(n6292), .X(n6289) );
  nor_x1_sg U5832 ( .A(n6277), .B(n6278), .X(n6276) );
  nor_x1_sg U5833 ( .A(n6220), .B(n6221), .X(n6219) );
  nor_x1_sg U5834 ( .A(n6226), .B(n6227), .X(n6224) );
  nor_x1_sg U5835 ( .A(n6228), .B(n6229), .X(n6218) );
  nor_x1_sg U5836 ( .A(n6246), .B(n6247), .X(n6236) );
  nor_x1_sg U5837 ( .A(n6252), .B(n6253), .X(n6250) );
  nor_x1_sg U5838 ( .A(n6238), .B(n6239), .X(n6237) );
  nor_x1_sg U5839 ( .A(n6181), .B(n6182), .X(n6180) );
  nor_x1_sg U5840 ( .A(n6187), .B(n6188), .X(n6185) );
  nor_x1_sg U5841 ( .A(n6189), .B(n6190), .X(n6179) );
  nor_x1_sg U5842 ( .A(n6207), .B(n6208), .X(n6197) );
  nor_x1_sg U5843 ( .A(n6213), .B(n6214), .X(n6211) );
  nor_x1_sg U5844 ( .A(n6199), .B(n6200), .X(n6198) );
  nor_x1_sg U5845 ( .A(n6142), .B(n6143), .X(n6141) );
  nor_x1_sg U5846 ( .A(n6148), .B(n6149), .X(n6146) );
  nor_x1_sg U5847 ( .A(n6150), .B(n6151), .X(n6140) );
  nor_x1_sg U5848 ( .A(n6168), .B(n6169), .X(n6158) );
  nor_x1_sg U5849 ( .A(n6174), .B(n6175), .X(n6172) );
  nor_x1_sg U5850 ( .A(n6160), .B(n6161), .X(n6159) );
  nor_x1_sg U5851 ( .A(n6103), .B(n6104), .X(n6102) );
  nor_x1_sg U5852 ( .A(n6109), .B(n6110), .X(n6107) );
  nor_x1_sg U5853 ( .A(n6111), .B(n6112), .X(n6101) );
  nor_x1_sg U5854 ( .A(n6129), .B(n6130), .X(n6119) );
  nor_x1_sg U5855 ( .A(n6135), .B(n6136), .X(n6133) );
  nor_x1_sg U5856 ( .A(n6121), .B(n6122), .X(n6120) );
  nor_x1_sg U5857 ( .A(n6044), .B(n6045), .X(n6043) );
  nor_x1_sg U5858 ( .A(n6053), .B(n6054), .X(n6050) );
  nor_x1_sg U5859 ( .A(n6057), .B(n6058), .X(n6042) );
  nor_x1_sg U5860 ( .A(n6085), .B(n6086), .X(n6070) );
  nor_x1_sg U5861 ( .A(n6094), .B(n6095), .X(n6091) );
  nor_x1_sg U5862 ( .A(n6072), .B(n6073), .X(n6071) );
  nand_x1_sg U5863 ( .A(n5252), .B(n5253), .X(n5251) );
  inv_x1_sg U5864 ( .A(\buff_mem[5][11] ), .X(n7779) );
  inv_x1_sg U5865 ( .A(\buff_mem[7][11] ), .X(n7619) );
  inv_x1_sg U5866 ( .A(\buff_mem[11][11] ), .X(n7777) );
  inv_x1_sg U5867 ( .A(\buff_mem[15][11] ), .X(n7617) );
  inv_x1_sg U5868 ( .A(\buff_mem[17][11] ), .X(n7615) );
  inv_x1_sg U5869 ( .A(\buff_mem[18][11] ), .X(n7613) );
  inv_x1_sg U5870 ( .A(\buff_mem[19][11] ), .X(n7611) );
  inv_x1_sg U5871 ( .A(\buff_mem[0][11] ), .X(n7609) );
  inv_x1_sg U5872 ( .A(\buff_mem[1][11] ), .X(n7775) );
  inv_x1_sg U5873 ( .A(\buff_mem[2][11] ), .X(n7607) );
  inv_x1_sg U5874 ( .A(\buff_mem[4][11] ), .X(n7773) );
  inv_x1_sg U5875 ( .A(\buff_mem[5][10] ), .X(n7771) );
  inv_x1_sg U5876 ( .A(\buff_mem[7][10] ), .X(n7605) );
  inv_x1_sg U5877 ( .A(\buff_mem[11][10] ), .X(n7769) );
  inv_x1_sg U5878 ( .A(\buff_mem[15][10] ), .X(n7603) );
  inv_x1_sg U5879 ( .A(\buff_mem[17][10] ), .X(n7601) );
  inv_x1_sg U5880 ( .A(\buff_mem[18][10] ), .X(n7599) );
  inv_x1_sg U5881 ( .A(\buff_mem[19][10] ), .X(n7597) );
  inv_x1_sg U5882 ( .A(\buff_mem[0][10] ), .X(n7595) );
  inv_x1_sg U5883 ( .A(\buff_mem[1][10] ), .X(n7767) );
  inv_x1_sg U5884 ( .A(\buff_mem[2][10] ), .X(n7593) );
  inv_x1_sg U5885 ( .A(\buff_mem[4][10] ), .X(n7765) );
  inv_x1_sg U5886 ( .A(\buff_mem[5][9] ), .X(n7763) );
  inv_x1_sg U5887 ( .A(\buff_mem[7][9] ), .X(n7591) );
  inv_x1_sg U5888 ( .A(\buff_mem[11][9] ), .X(n7761) );
  inv_x1_sg U5889 ( .A(\buff_mem[15][9] ), .X(n7589) );
  inv_x1_sg U5890 ( .A(\buff_mem[17][9] ), .X(n7587) );
  inv_x1_sg U5891 ( .A(\buff_mem[18][9] ), .X(n7585) );
  inv_x1_sg U5892 ( .A(\buff_mem[19][9] ), .X(n7583) );
  inv_x1_sg U5893 ( .A(\buff_mem[0][9] ), .X(n7581) );
  inv_x1_sg U5894 ( .A(\buff_mem[1][9] ), .X(n7759) );
  inv_x1_sg U5895 ( .A(\buff_mem[2][9] ), .X(n7579) );
  inv_x1_sg U5896 ( .A(\buff_mem[4][9] ), .X(n7757) );
  inv_x1_sg U5897 ( .A(\buff_mem[5][8] ), .X(n7755) );
  inv_x1_sg U5898 ( .A(\buff_mem[7][8] ), .X(n7577) );
  inv_x1_sg U5899 ( .A(\buff_mem[11][8] ), .X(n7753) );
  inv_x1_sg U5900 ( .A(\buff_mem[15][8] ), .X(n7575) );
  inv_x1_sg U5901 ( .A(\buff_mem[17][8] ), .X(n7573) );
  inv_x1_sg U5902 ( .A(\buff_mem[18][8] ), .X(n7571) );
  inv_x1_sg U5903 ( .A(\buff_mem[19][8] ), .X(n7569) );
  inv_x1_sg U5904 ( .A(\buff_mem[0][8] ), .X(n7567) );
  inv_x1_sg U5905 ( .A(\buff_mem[1][8] ), .X(n7751) );
  inv_x1_sg U5906 ( .A(\buff_mem[2][8] ), .X(n7565) );
  inv_x1_sg U5907 ( .A(\buff_mem[4][8] ), .X(n7749) );
  inv_x1_sg U5908 ( .A(\buff_mem[5][7] ), .X(n7747) );
  inv_x1_sg U5909 ( .A(\buff_mem[7][7] ), .X(n7563) );
  inv_x1_sg U5910 ( .A(\buff_mem[11][7] ), .X(n7745) );
  inv_x1_sg U5911 ( .A(\buff_mem[15][7] ), .X(n7561) );
  inv_x1_sg U5912 ( .A(\buff_mem[17][7] ), .X(n7559) );
  inv_x1_sg U5913 ( .A(\buff_mem[18][7] ), .X(n7557) );
  inv_x1_sg U5914 ( .A(\buff_mem[19][7] ), .X(n7555) );
  inv_x1_sg U5915 ( .A(\buff_mem[0][7] ), .X(n7553) );
  inv_x1_sg U5916 ( .A(\buff_mem[1][7] ), .X(n7743) );
  inv_x1_sg U5917 ( .A(\buff_mem[2][7] ), .X(n7551) );
  inv_x1_sg U5918 ( .A(\buff_mem[4][7] ), .X(n7741) );
  inv_x1_sg U5919 ( .A(\buff_mem[5][6] ), .X(n7739) );
  inv_x1_sg U5920 ( .A(\buff_mem[7][6] ), .X(n7549) );
  inv_x1_sg U5921 ( .A(\buff_mem[11][6] ), .X(n7737) );
  inv_x1_sg U5922 ( .A(\buff_mem[15][6] ), .X(n7547) );
  inv_x1_sg U5923 ( .A(\buff_mem[17][6] ), .X(n7545) );
  inv_x1_sg U5924 ( .A(\buff_mem[18][6] ), .X(n7543) );
  inv_x1_sg U5925 ( .A(\buff_mem[19][6] ), .X(n7541) );
  inv_x1_sg U5926 ( .A(\buff_mem[0][6] ), .X(n7539) );
  inv_x1_sg U5927 ( .A(\buff_mem[1][6] ), .X(n7735) );
  inv_x1_sg U5928 ( .A(\buff_mem[2][6] ), .X(n7537) );
  inv_x1_sg U5929 ( .A(\buff_mem[4][6] ), .X(n7733) );
  inv_x1_sg U5930 ( .A(\buff_mem[5][5] ), .X(n7731) );
  inv_x1_sg U5931 ( .A(\buff_mem[7][5] ), .X(n7535) );
  inv_x1_sg U5932 ( .A(\buff_mem[11][5] ), .X(n7729) );
  inv_x1_sg U5933 ( .A(\buff_mem[15][5] ), .X(n7533) );
  inv_x1_sg U5934 ( .A(\buff_mem[17][5] ), .X(n7531) );
  inv_x1_sg U5935 ( .A(\buff_mem[18][5] ), .X(n7529) );
  inv_x1_sg U5936 ( .A(\buff_mem[19][5] ), .X(n7527) );
  inv_x1_sg U5937 ( .A(\buff_mem[0][5] ), .X(n7525) );
  inv_x1_sg U5938 ( .A(\buff_mem[1][5] ), .X(n7727) );
  inv_x1_sg U5939 ( .A(\buff_mem[2][5] ), .X(n7523) );
  inv_x1_sg U5940 ( .A(\buff_mem[4][5] ), .X(n7725) );
  inv_x1_sg U5941 ( .A(\buff_mem[5][4] ), .X(n7723) );
  inv_x1_sg U5942 ( .A(\buff_mem[7][4] ), .X(n7521) );
  inv_x1_sg U5943 ( .A(\buff_mem[11][4] ), .X(n7721) );
  inv_x1_sg U5944 ( .A(\buff_mem[15][4] ), .X(n7519) );
  inv_x1_sg U5945 ( .A(\buff_mem[17][4] ), .X(n7517) );
  inv_x1_sg U5946 ( .A(\buff_mem[18][4] ), .X(n7515) );
  inv_x1_sg U5947 ( .A(\buff_mem[19][4] ), .X(n7513) );
  inv_x1_sg U5948 ( .A(\buff_mem[0][4] ), .X(n7511) );
  inv_x1_sg U5949 ( .A(\buff_mem[1][4] ), .X(n7719) );
  inv_x1_sg U5950 ( .A(\buff_mem[2][4] ), .X(n7509) );
  inv_x1_sg U5951 ( .A(\buff_mem[4][4] ), .X(n7717) );
  inv_x1_sg U5952 ( .A(\buff_mem[5][3] ), .X(n7715) );
  inv_x1_sg U5953 ( .A(\buff_mem[7][3] ), .X(n7507) );
  inv_x1_sg U5954 ( .A(\buff_mem[11][3] ), .X(n7713) );
  inv_x1_sg U5955 ( .A(\buff_mem[15][3] ), .X(n7505) );
  inv_x1_sg U5956 ( .A(\buff_mem[17][3] ), .X(n7503) );
  inv_x1_sg U5957 ( .A(\buff_mem[18][3] ), .X(n7501) );
  inv_x1_sg U5958 ( .A(\buff_mem[19][3] ), .X(n7499) );
  inv_x1_sg U5959 ( .A(\buff_mem[0][3] ), .X(n7497) );
  inv_x1_sg U5960 ( .A(\buff_mem[1][3] ), .X(n7711) );
  inv_x1_sg U5961 ( .A(\buff_mem[2][3] ), .X(n7495) );
  inv_x1_sg U5962 ( .A(\buff_mem[4][3] ), .X(n7709) );
  inv_x1_sg U5963 ( .A(\buff_mem[5][2] ), .X(n7707) );
  inv_x1_sg U5964 ( .A(\buff_mem[7][2] ), .X(n7493) );
  inv_x1_sg U5965 ( .A(\buff_mem[11][2] ), .X(n7705) );
  inv_x1_sg U5966 ( .A(\buff_mem[15][2] ), .X(n7491) );
  inv_x1_sg U5967 ( .A(\buff_mem[17][2] ), .X(n7489) );
  inv_x1_sg U5968 ( .A(\buff_mem[18][2] ), .X(n7487) );
  inv_x1_sg U5969 ( .A(\buff_mem[19][2] ), .X(n7485) );
  inv_x1_sg U5970 ( .A(\buff_mem[0][2] ), .X(n7483) );
  inv_x1_sg U5971 ( .A(\buff_mem[1][2] ), .X(n7703) );
  inv_x1_sg U5972 ( .A(\buff_mem[2][2] ), .X(n7481) );
  inv_x1_sg U5973 ( .A(\buff_mem[4][2] ), .X(n7701) );
  inv_x1_sg U5974 ( .A(\buff_mem[5][1] ), .X(n7699) );
  inv_x1_sg U5975 ( .A(\buff_mem[7][1] ), .X(n7479) );
  inv_x1_sg U5976 ( .A(\buff_mem[11][1] ), .X(n7697) );
  inv_x1_sg U5977 ( .A(\buff_mem[15][1] ), .X(n7477) );
  inv_x1_sg U5978 ( .A(\buff_mem[17][1] ), .X(n7475) );
  inv_x1_sg U5979 ( .A(\buff_mem[18][1] ), .X(n7473) );
  inv_x1_sg U5980 ( .A(\buff_mem[19][1] ), .X(n7471) );
  inv_x1_sg U5981 ( .A(\buff_mem[0][1] ), .X(n7469) );
  inv_x1_sg U5982 ( .A(\buff_mem[1][1] ), .X(n7695) );
  inv_x1_sg U5983 ( .A(\buff_mem[2][1] ), .X(n7467) );
  inv_x1_sg U5984 ( .A(\buff_mem[4][1] ), .X(n7693) );
  inv_x1_sg U5985 ( .A(\buff_mem[5][0] ), .X(n7691) );
  inv_x1_sg U5986 ( .A(\buff_mem[7][0] ), .X(n7465) );
  inv_x1_sg U5987 ( .A(\buff_mem[11][0] ), .X(n7689) );
  inv_x1_sg U5988 ( .A(\buff_mem[15][0] ), .X(n7463) );
  inv_x1_sg U5989 ( .A(\buff_mem[17][0] ), .X(n7461) );
  inv_x1_sg U5990 ( .A(\buff_mem[18][0] ), .X(n7459) );
  inv_x1_sg U5991 ( .A(\buff_mem[19][0] ), .X(n7457) );
  inv_x1_sg U5992 ( .A(\buff_mem[0][0] ), .X(n7455) );
  inv_x1_sg U5993 ( .A(\buff_mem[1][0] ), .X(n7687) );
  inv_x1_sg U5994 ( .A(\buff_mem[2][0] ), .X(n7453) );
  inv_x1_sg U5995 ( .A(\buff_mem[4][0] ), .X(n7685) );
  inv_x1_sg U5996 ( .A(\buff_mem[4][19] ), .X(n7683) );
  inv_x1_sg U5997 ( .A(\buff_mem[5][19] ), .X(n7681) );
  inv_x1_sg U5998 ( .A(\buff_mem[7][19] ), .X(n7451) );
  inv_x1_sg U5999 ( .A(\buff_mem[11][19] ), .X(n7679) );
  inv_x1_sg U6000 ( .A(\buff_mem[15][19] ), .X(n7449) );
  inv_x1_sg U6001 ( .A(\buff_mem[17][19] ), .X(n7447) );
  inv_x1_sg U6002 ( .A(\buff_mem[18][19] ), .X(n7445) );
  inv_x1_sg U6003 ( .A(\buff_mem[19][19] ), .X(n7443) );
  inv_x1_sg U6004 ( .A(\buff_mem[0][19] ), .X(n7441) );
  inv_x1_sg U6005 ( .A(\buff_mem[1][19] ), .X(n7677) );
  inv_x1_sg U6006 ( .A(\buff_mem[2][19] ), .X(n7439) );
  inv_x1_sg U6007 ( .A(\buff_mem[4][18] ), .X(n7675) );
  inv_x1_sg U6008 ( .A(\buff_mem[5][18] ), .X(n7673) );
  inv_x1_sg U6009 ( .A(\buff_mem[7][18] ), .X(n7437) );
  inv_x1_sg U6010 ( .A(\buff_mem[11][18] ), .X(n7671) );
  inv_x1_sg U6011 ( .A(\buff_mem[15][18] ), .X(n7435) );
  inv_x1_sg U6012 ( .A(\buff_mem[17][18] ), .X(n7433) );
  inv_x1_sg U6013 ( .A(\buff_mem[18][18] ), .X(n7431) );
  inv_x1_sg U6014 ( .A(\buff_mem[19][18] ), .X(n7429) );
  inv_x1_sg U6015 ( .A(\buff_mem[0][18] ), .X(n7427) );
  inv_x1_sg U6016 ( .A(\buff_mem[1][18] ), .X(n7669) );
  inv_x1_sg U6017 ( .A(\buff_mem[2][18] ), .X(n7425) );
  inv_x1_sg U6018 ( .A(\buff_mem[4][17] ), .X(n7667) );
  inv_x1_sg U6019 ( .A(\buff_mem[5][17] ), .X(n7665) );
  inv_x1_sg U6020 ( .A(\buff_mem[7][17] ), .X(n7423) );
  inv_x1_sg U6021 ( .A(\buff_mem[11][17] ), .X(n7663) );
  inv_x1_sg U6022 ( .A(\buff_mem[15][17] ), .X(n7421) );
  inv_x1_sg U6023 ( .A(\buff_mem[17][17] ), .X(n7419) );
  inv_x1_sg U6024 ( .A(\buff_mem[18][17] ), .X(n7417) );
  inv_x1_sg U6025 ( .A(\buff_mem[19][17] ), .X(n7415) );
  inv_x1_sg U6026 ( .A(\buff_mem[0][17] ), .X(n7413) );
  inv_x1_sg U6027 ( .A(\buff_mem[1][17] ), .X(n7661) );
  inv_x1_sg U6028 ( .A(\buff_mem[2][17] ), .X(n7411) );
  inv_x1_sg U6029 ( .A(\buff_mem[4][16] ), .X(n7659) );
  inv_x1_sg U6030 ( .A(\buff_mem[5][16] ), .X(n7657) );
  inv_x1_sg U6031 ( .A(\buff_mem[7][16] ), .X(n7409) );
  inv_x1_sg U6032 ( .A(\buff_mem[11][16] ), .X(n7655) );
  inv_x1_sg U6033 ( .A(\buff_mem[15][16] ), .X(n7407) );
  inv_x1_sg U6034 ( .A(\buff_mem[17][16] ), .X(n7405) );
  inv_x1_sg U6035 ( .A(\buff_mem[18][16] ), .X(n7403) );
  inv_x1_sg U6036 ( .A(\buff_mem[19][16] ), .X(n7401) );
  inv_x1_sg U6037 ( .A(\buff_mem[0][16] ), .X(n7399) );
  inv_x1_sg U6038 ( .A(\buff_mem[1][16] ), .X(n7653) );
  inv_x1_sg U6039 ( .A(\buff_mem[2][16] ), .X(n7397) );
  inv_x1_sg U6040 ( .A(\buff_mem[4][15] ), .X(n7651) );
  inv_x1_sg U6041 ( .A(\buff_mem[5][15] ), .X(n7649) );
  inv_x1_sg U6042 ( .A(\buff_mem[7][15] ), .X(n7395) );
  inv_x1_sg U6043 ( .A(\buff_mem[11][15] ), .X(n7647) );
  inv_x1_sg U6044 ( .A(\buff_mem[15][15] ), .X(n7393) );
  inv_x1_sg U6045 ( .A(\buff_mem[17][15] ), .X(n7391) );
  inv_x1_sg U6046 ( .A(\buff_mem[18][15] ), .X(n7389) );
  inv_x1_sg U6047 ( .A(\buff_mem[19][15] ), .X(n7387) );
  inv_x1_sg U6048 ( .A(\buff_mem[0][15] ), .X(n7385) );
  inv_x1_sg U6049 ( .A(\buff_mem[1][15] ), .X(n7645) );
  inv_x1_sg U6050 ( .A(\buff_mem[2][15] ), .X(n7383) );
  inv_x1_sg U6051 ( .A(\buff_mem[4][14] ), .X(n7643) );
  inv_x1_sg U6052 ( .A(\buff_mem[5][14] ), .X(n7641) );
  inv_x1_sg U6053 ( .A(\buff_mem[7][14] ), .X(n7381) );
  inv_x1_sg U6054 ( .A(\buff_mem[11][14] ), .X(n7639) );
  inv_x1_sg U6055 ( .A(\buff_mem[15][14] ), .X(n7379) );
  inv_x1_sg U6056 ( .A(\buff_mem[17][14] ), .X(n7377) );
  inv_x1_sg U6057 ( .A(\buff_mem[18][14] ), .X(n7375) );
  inv_x1_sg U6058 ( .A(\buff_mem[19][14] ), .X(n7373) );
  inv_x1_sg U6059 ( .A(\buff_mem[0][14] ), .X(n7371) );
  inv_x1_sg U6060 ( .A(\buff_mem[1][14] ), .X(n7637) );
  inv_x1_sg U6061 ( .A(\buff_mem[2][14] ), .X(n7369) );
  inv_x1_sg U6062 ( .A(\buff_mem[4][13] ), .X(n7635) );
  inv_x1_sg U6063 ( .A(\buff_mem[5][13] ), .X(n7633) );
  inv_x1_sg U6064 ( .A(\buff_mem[7][13] ), .X(n7367) );
  inv_x1_sg U6065 ( .A(\buff_mem[11][13] ), .X(n7631) );
  inv_x1_sg U6066 ( .A(\buff_mem[15][13] ), .X(n7365) );
  inv_x1_sg U6067 ( .A(\buff_mem[17][13] ), .X(n7363) );
  inv_x1_sg U6068 ( .A(\buff_mem[18][13] ), .X(n7361) );
  inv_x1_sg U6069 ( .A(\buff_mem[19][13] ), .X(n7359) );
  inv_x1_sg U6070 ( .A(\buff_mem[0][13] ), .X(n7357) );
  inv_x1_sg U6071 ( .A(\buff_mem[1][13] ), .X(n7629) );
  inv_x1_sg U6072 ( .A(\buff_mem[2][13] ), .X(n7355) );
  inv_x1_sg U6073 ( .A(\buff_mem[4][12] ), .X(n7627) );
  inv_x1_sg U6074 ( .A(\buff_mem[5][12] ), .X(n7625) );
  inv_x1_sg U6075 ( .A(\buff_mem[7][12] ), .X(n7353) );
  inv_x1_sg U6076 ( .A(\buff_mem[11][12] ), .X(n7623) );
  inv_x1_sg U6077 ( .A(\buff_mem[15][12] ), .X(n7351) );
  inv_x1_sg U6078 ( .A(\buff_mem[17][12] ), .X(n7349) );
  inv_x1_sg U6079 ( .A(\buff_mem[18][12] ), .X(n7347) );
  inv_x1_sg U6080 ( .A(\buff_mem[19][12] ), .X(n7345) );
  inv_x1_sg U6081 ( .A(\buff_mem[0][12] ), .X(n7343) );
  inv_x1_sg U6082 ( .A(\buff_mem[1][12] ), .X(n7621) );
  inv_x1_sg U6083 ( .A(\buff_mem[2][12] ), .X(n7341) );
  nand_x1_sg U6084 ( .A(n5169), .B(n5170), .X(n5168) );
  nand_x1_sg U6085 ( .A(n6029), .B(n6030), .X(n7258) );
  nand_x1_sg U6086 ( .A(n6033), .B(n6034), .X(n7259) );
  nand_x1_sg U6087 ( .A(n6025), .B(n6026), .X(n7256) );
  nand_x1_sg U6088 ( .A(n6021), .B(n6022), .X(n7255) );
  nand_x1_sg U6089 ( .A(n4842), .B(n5247), .X(n6907) );
  inv_x1_sg U6090 ( .A(n5248), .X(n4842) );
  nand_x1_sg U6091 ( .A(n5307), .B(n5308), .X(n6923) );
  nand_x1_sg U6092 ( .A(n8153), .B(n8114), .X(n5308) );
  nand_x1_sg U6093 ( .A(n5281), .B(n5282), .X(n6910) );
  nand_x1_sg U6094 ( .A(n8154), .B(n8114), .X(n5282) );
  nand_x1_sg U6095 ( .A(n5297), .B(n5298), .X(n6918) );
  nand_x1_sg U6096 ( .A(n8151), .B(n8114), .X(n5298) );
  nand_x1_sg U6097 ( .A(n5303), .B(n5304), .X(n6921) );
  nand_x1_sg U6098 ( .A(n8163), .B(n8114), .X(n5304) );
  nand_x1_sg U6099 ( .A(n5305), .B(n5306), .X(n6922) );
  nand_x1_sg U6100 ( .A(n8166), .B(n8114), .X(n5306) );
  nand_x1_sg U6101 ( .A(n5299), .B(n5300), .X(n6919) );
  nand_x1_sg U6102 ( .A(n8164), .B(n8114), .X(n5300) );
  nand_x1_sg U6103 ( .A(n5291), .B(n5292), .X(n6915) );
  nand_x1_sg U6104 ( .A(n8165), .B(n8114), .X(n5292) );
  nand_x1_sg U6105 ( .A(n5090), .B(n5091), .X(n6853) );
  nand_x1_sg U6106 ( .A(n8114), .B(n8155), .X(n5091) );
  nand_x1_sg U6107 ( .A(n5293), .B(n5294), .X(n6916) );
  nand_x1_sg U6108 ( .A(n8156), .B(n8114), .X(n5294) );
  nand_x1_sg U6109 ( .A(n5279), .B(n5280), .X(n6909) );
  nand_x1_sg U6110 ( .A(n8157), .B(n8114), .X(n5280) );
  nand_x1_sg U6111 ( .A(n5289), .B(n5290), .X(n6914) );
  nand_x1_sg U6112 ( .A(n8158), .B(n4879), .X(n5290) );
  nand_x1_sg U6113 ( .A(n5145), .B(n5146), .X(n6879) );
  nand_x1_sg U6114 ( .A(n8107), .B(n8114), .X(n5146) );
  nand_x1_sg U6115 ( .A(n5283), .B(n5284), .X(n6911) );
  nand_x1_sg U6116 ( .A(n8110), .B(n8114), .X(n5284) );
  nand_x1_sg U6117 ( .A(n5277), .B(n5278), .X(n6908) );
  nand_x1_sg U6118 ( .A(n8109), .B(n8114), .X(n5278) );
  nand_x1_sg U6119 ( .A(n5287), .B(n5288), .X(n6913) );
  nand_x1_sg U6120 ( .A(n8108), .B(n8114), .X(n5288) );
  nand_x1_sg U6121 ( .A(n5309), .B(n5310), .X(n6924) );
  nand_x1_sg U6122 ( .A(n8159), .B(n8114), .X(n5310) );
  nand_x1_sg U6123 ( .A(n5295), .B(n5296), .X(n6917) );
  nand_x1_sg U6124 ( .A(n8161), .B(n8114), .X(n5296) );
  nand_x1_sg U6125 ( .A(n5285), .B(n5286), .X(n6912) );
  nand_x1_sg U6126 ( .A(n8160), .B(n8114), .X(n5286) );
  nand_x1_sg U6127 ( .A(n5301), .B(n5302), .X(n6920) );
  nand_x1_sg U6128 ( .A(n8162), .B(n8114), .X(n5302) );
  nand_x1_sg U6129 ( .A(n5311), .B(n5312), .X(n6925) );
  nand_x1_sg U6130 ( .A(n8152), .B(n8114), .X(n5312) );
  nand_x1_sg U6131 ( .A(n5396), .B(n5397), .X(n6966) );
  nand_x1_sg U6132 ( .A(n8153), .B(n8120), .X(n5397) );
  nand_x1_sg U6133 ( .A(n5441), .B(n5442), .X(n6988) );
  nand_x1_sg U6134 ( .A(n8154), .B(n8120), .X(n5442) );
  nand_x1_sg U6135 ( .A(n5320), .B(n5321), .X(n6929) );
  nand_x1_sg U6136 ( .A(n8151), .B(n8120), .X(n5321) );
  nand_x1_sg U6137 ( .A(n5861), .B(n5862), .X(n7188) );
  nand_x1_sg U6138 ( .A(n8163), .B(n8120), .X(n5862) );
  nand_x1_sg U6139 ( .A(n5967), .B(n5968), .X(n7239) );
  nand_x1_sg U6140 ( .A(n8166), .B(n8120), .X(n5968) );
  nand_x1_sg U6141 ( .A(n5898), .B(n5899), .X(n7206) );
  nand_x1_sg U6142 ( .A(n8164), .B(n8120), .X(n5899) );
  nand_x1_sg U6143 ( .A(n5935), .B(n5936), .X(n7224) );
  nand_x1_sg U6144 ( .A(n8165), .B(n8120), .X(n5936) );
  nand_x1_sg U6145 ( .A(n5084), .B(n5085), .X(n6850) );
  nand_x1_sg U6146 ( .A(n8120), .B(n8155), .X(n5085) );
  nand_x1_sg U6147 ( .A(n5473), .B(n5474), .X(n7002) );
  nand_x1_sg U6148 ( .A(n8156), .B(n8120), .X(n5474) );
  nand_x1_sg U6149 ( .A(n5511), .B(n5512), .X(n7021) );
  nand_x1_sg U6150 ( .A(n8157), .B(n8120), .X(n5512) );
  nand_x1_sg U6151 ( .A(n5541), .B(n5542), .X(n7036) );
  nand_x1_sg U6152 ( .A(n8158), .B(n4876), .X(n5542) );
  nand_x1_sg U6153 ( .A(n5143), .B(n5144), .X(n6878) );
  nand_x1_sg U6154 ( .A(n8107), .B(n8120), .X(n5144) );
  nand_x1_sg U6155 ( .A(n5838), .B(n5839), .X(n7178) );
  nand_x1_sg U6156 ( .A(n8110), .B(n8120), .X(n5839) );
  nand_x1_sg U6157 ( .A(n5780), .B(n5781), .X(n7149) );
  nand_x1_sg U6158 ( .A(n8109), .B(n8120), .X(n5781) );
  nand_x1_sg U6159 ( .A(n5766), .B(n5767), .X(n7142) );
  nand_x1_sg U6160 ( .A(n8108), .B(n8120), .X(n5767) );
  nand_x1_sg U6161 ( .A(n5599), .B(n5600), .X(n7060) );
  nand_x1_sg U6162 ( .A(n8159), .B(n8120), .X(n5600) );
  nand_x1_sg U6163 ( .A(n5670), .B(n5671), .X(n7095) );
  nand_x1_sg U6164 ( .A(n8161), .B(n8120), .X(n5671) );
  nand_x1_sg U6165 ( .A(n5640), .B(n5641), .X(n7080) );
  nand_x1_sg U6166 ( .A(n8160), .B(n8120), .X(n5641) );
  nand_x1_sg U6167 ( .A(n5712), .B(n5713), .X(n7116) );
  nand_x1_sg U6168 ( .A(n8162), .B(n8120), .X(n5713) );
  nand_x1_sg U6169 ( .A(n5364), .B(n5365), .X(n6950) );
  nand_x1_sg U6170 ( .A(n8152), .B(n8120), .X(n5365) );
  nand_x1_sg U6171 ( .A(n5418), .B(n5419), .X(n6977) );
  nand_x1_sg U6172 ( .A(n8153), .B(n8148), .X(n5419) );
  nand_x1_sg U6173 ( .A(n5449), .B(n5450), .X(n6992) );
  nand_x1_sg U6174 ( .A(n8154), .B(n8148), .X(n5450) );
  nand_x1_sg U6175 ( .A(n5344), .B(n5345), .X(n6941) );
  nand_x1_sg U6176 ( .A(n8151), .B(n4862), .X(n5345) );
  nand_x1_sg U6177 ( .A(n5885), .B(n5886), .X(n7200) );
  nand_x1_sg U6178 ( .A(n8163), .B(n8148), .X(n5886) );
  nand_x1_sg U6179 ( .A(n6009), .B(n6010), .X(n7253) );
  nand_x1_sg U6180 ( .A(n8166), .B(n8148), .X(n6010) );
  nand_x1_sg U6181 ( .A(n5922), .B(n5923), .X(n7218) );
  nand_x1_sg U6182 ( .A(n8164), .B(n8148), .X(n5923) );
  nand_x1_sg U6183 ( .A(n5957), .B(n5958), .X(n7235) );
  nand_x1_sg U6184 ( .A(n8165), .B(n8148), .X(n5958) );
  nand_x1_sg U6185 ( .A(n5116), .B(n5117), .X(n6866) );
  nand_x1_sg U6186 ( .A(n8148), .B(n8155), .X(n5117) );
  nand_x1_sg U6187 ( .A(n5499), .B(n5500), .X(n7015) );
  nand_x1_sg U6188 ( .A(n8156), .B(n8148), .X(n5500) );
  nand_x1_sg U6189 ( .A(n5505), .B(n5506), .X(n7018) );
  nand_x1_sg U6190 ( .A(n8157), .B(n8148), .X(n5506) );
  nand_x1_sg U6191 ( .A(n5567), .B(n5568), .X(n7049) );
  nand_x1_sg U6192 ( .A(n8158), .B(n8148), .X(n5568) );
  nand_x1_sg U6193 ( .A(n5135), .B(n5136), .X(n6874) );
  nand_x1_sg U6194 ( .A(n8107), .B(n8148), .X(n5136) );
  nand_x1_sg U6195 ( .A(n5824), .B(n5825), .X(n7171) );
  nand_x1_sg U6196 ( .A(n8110), .B(n8148), .X(n5825) );
  nand_x1_sg U6197 ( .A(n5808), .B(n5809), .X(n7163) );
  nand_x1_sg U6198 ( .A(n8109), .B(n8148), .X(n5809) );
  nand_x1_sg U6199 ( .A(n5752), .B(n5753), .X(n7135) );
  nand_x1_sg U6200 ( .A(n8108), .B(n8148), .X(n5753) );
  nand_x1_sg U6201 ( .A(n5623), .B(n5624), .X(n7072) );
  nand_x1_sg U6202 ( .A(n8159), .B(n8148), .X(n5624) );
  nand_x1_sg U6203 ( .A(n5698), .B(n5699), .X(n7109) );
  nand_x1_sg U6204 ( .A(n8161), .B(n8148), .X(n5699) );
  nand_x1_sg U6205 ( .A(n5660), .B(n5661), .X(n7090) );
  nand_x1_sg U6206 ( .A(n8160), .B(n8148), .X(n5661) );
  nand_x1_sg U6207 ( .A(n5734), .B(n5735), .X(n7127) );
  nand_x1_sg U6208 ( .A(n8162), .B(n8148), .X(n5735) );
  nand_x1_sg U6209 ( .A(n5378), .B(n5379), .X(n6957) );
  nand_x1_sg U6210 ( .A(n8152), .B(n8148), .X(n5379) );
  nand_x1_sg U6211 ( .A(n5416), .B(n5417), .X(n6976) );
  nand_x1_sg U6212 ( .A(n8153), .B(n8122), .X(n5417) );
  nand_x1_sg U6213 ( .A(n5425), .B(n5426), .X(n6980) );
  nand_x1_sg U6214 ( .A(n8154), .B(n8122), .X(n5426) );
  nand_x1_sg U6215 ( .A(n5342), .B(n5343), .X(n6940) );
  nand_x1_sg U6216 ( .A(n8151), .B(n8122), .X(n5343) );
  nand_x1_sg U6217 ( .A(n5855), .B(n5856), .X(n7185) );
  nand_x1_sg U6218 ( .A(n8163), .B(n8122), .X(n5856) );
  nand_x1_sg U6219 ( .A(n5970), .B(n5971), .X(n7240) );
  nand_x1_sg U6220 ( .A(n8166), .B(n8122), .X(n5971) );
  nand_x1_sg U6221 ( .A(n5892), .B(n5893), .X(n7203) );
  nand_x1_sg U6222 ( .A(n8164), .B(n8122), .X(n5893) );
  nand_x1_sg U6223 ( .A(n5929), .B(n5930), .X(n7221) );
  nand_x1_sg U6224 ( .A(n8165), .B(n8122), .X(n5930) );
  nand_x1_sg U6225 ( .A(n5098), .B(n5099), .X(n6857) );
  nand_x1_sg U6226 ( .A(n8122), .B(n8155), .X(n5099) );
  nand_x1_sg U6227 ( .A(n5491), .B(n5492), .X(n7011) );
  nand_x1_sg U6228 ( .A(n8156), .B(n8122), .X(n5492) );
  nand_x1_sg U6229 ( .A(n5521), .B(n5522), .X(n7026) );
  nand_x1_sg U6230 ( .A(n8157), .B(n8122), .X(n5522) );
  nand_x1_sg U6231 ( .A(n5547), .B(n5548), .X(n7039) );
  nand_x1_sg U6232 ( .A(n8158), .B(n4875), .X(n5548) );
  nand_x1_sg U6233 ( .A(n5127), .B(n5128), .X(n6870) );
  nand_x1_sg U6234 ( .A(n8107), .B(n8122), .X(n5128) );
  nand_x1_sg U6235 ( .A(n5816), .B(n5817), .X(n7167) );
  nand_x1_sg U6236 ( .A(n8110), .B(n8122), .X(n5817) );
  nand_x1_sg U6237 ( .A(n5790), .B(n5791), .X(n7154) );
  nand_x1_sg U6238 ( .A(n8109), .B(n8122), .X(n5791) );
  nand_x1_sg U6239 ( .A(n5744), .B(n5745), .X(n7131) );
  nand_x1_sg U6240 ( .A(n8108), .B(n8122), .X(n5745) );
  nand_x1_sg U6241 ( .A(n5621), .B(n5622), .X(n7071) );
  nand_x1_sg U6242 ( .A(n8159), .B(n8122), .X(n5622) );
  nand_x1_sg U6243 ( .A(n5682), .B(n5683), .X(n7101) );
  nand_x1_sg U6244 ( .A(n8161), .B(n8122), .X(n5683) );
  nand_x1_sg U6245 ( .A(n5634), .B(n5635), .X(n7077) );
  nand_x1_sg U6246 ( .A(n8160), .B(n8122), .X(n5635) );
  nand_x1_sg U6247 ( .A(n5722), .B(n5723), .X(n7121) );
  nand_x1_sg U6248 ( .A(n8162), .B(n8122), .X(n5723) );
  nand_x1_sg U6249 ( .A(n5372), .B(n5373), .X(n6954) );
  nand_x1_sg U6250 ( .A(n8152), .B(n8122), .X(n5373) );
  nand_x1_sg U6251 ( .A(n5388), .B(n5389), .X(n6962) );
  nand_x1_sg U6252 ( .A(n8153), .B(n8140), .X(n5389) );
  nand_x1_sg U6253 ( .A(n5437), .B(n5438), .X(n6986) );
  nand_x1_sg U6254 ( .A(n8154), .B(n8140), .X(n5438) );
  nand_x1_sg U6255 ( .A(n5326), .B(n5327), .X(n6932) );
  nand_x1_sg U6256 ( .A(n8151), .B(n8140), .X(n5327) );
  nand_x1_sg U6257 ( .A(n5869), .B(n5870), .X(n7192) );
  nand_x1_sg U6258 ( .A(n8163), .B(n8140), .X(n5870) );
  nand_x1_sg U6259 ( .A(n5997), .B(n5998), .X(n7249) );
  nand_x1_sg U6260 ( .A(n8166), .B(n8140), .X(n5998) );
  nand_x1_sg U6261 ( .A(n5912), .B(n5913), .X(n7213) );
  nand_x1_sg U6262 ( .A(n8164), .B(n8140), .X(n5913) );
  nand_x1_sg U6263 ( .A(n5947), .B(n5948), .X(n7230) );
  nand_x1_sg U6264 ( .A(n8165), .B(n8140), .X(n5948) );
  nand_x1_sg U6265 ( .A(n5108), .B(n5109), .X(n6862) );
  nand_x1_sg U6266 ( .A(n8140), .B(n8155), .X(n5109) );
  nand_x1_sg U6267 ( .A(n5465), .B(n5466), .X(n6998) );
  nand_x1_sg U6268 ( .A(n8156), .B(n8140), .X(n5466) );
  nand_x1_sg U6269 ( .A(n5527), .B(n5528), .X(n7029) );
  nand_x1_sg U6270 ( .A(n8157), .B(n8140), .X(n5528) );
  nand_x1_sg U6271 ( .A(n5545), .B(n5546), .X(n7038) );
  nand_x1_sg U6272 ( .A(n8158), .B(n8140), .X(n5546) );
  nand_x1_sg U6273 ( .A(n5147), .B(n5148), .X(n6880) );
  nand_x1_sg U6274 ( .A(n8107), .B(n8140), .X(n5148) );
  nand_x1_sg U6275 ( .A(n5832), .B(n5833), .X(n7175) );
  nand_x1_sg U6276 ( .A(n8110), .B(n8140), .X(n5833) );
  nand_x1_sg U6277 ( .A(n5784), .B(n5785), .X(n7151) );
  nand_x1_sg U6278 ( .A(n8109), .B(n8140), .X(n5785) );
  nand_x1_sg U6279 ( .A(n5762), .B(n5763), .X(n7140) );
  nand_x1_sg U6280 ( .A(n8108), .B(n8140), .X(n5763) );
  nand_x1_sg U6281 ( .A(n5605), .B(n5606), .X(n7063) );
  nand_x1_sg U6282 ( .A(n8159), .B(n8140), .X(n5606) );
  nand_x1_sg U6283 ( .A(n5672), .B(n5673), .X(n7096) );
  nand_x1_sg U6284 ( .A(n8161), .B(n4866), .X(n5673) );
  nand_x1_sg U6285 ( .A(n5650), .B(n5651), .X(n7085) );
  nand_x1_sg U6286 ( .A(n8160), .B(n8140), .X(n5651) );
  nand_x1_sg U6287 ( .A(n5726), .B(n5727), .X(n7123) );
  nand_x1_sg U6288 ( .A(n8162), .B(n8140), .X(n5727) );
  nand_x1_sg U6289 ( .A(n5354), .B(n5355), .X(n6945) );
  nand_x1_sg U6290 ( .A(n8152), .B(n8140), .X(n5355) );
  nand_x1_sg U6291 ( .A(n5420), .B(n5421), .X(n6978) );
  nand_x1_sg U6292 ( .A(n8153), .B(n8132), .X(n5421) );
  nand_x1_sg U6293 ( .A(n5433), .B(n5434), .X(n6984) );
  nand_x1_sg U6294 ( .A(n8154), .B(n8132), .X(n5434) );
  nand_x1_sg U6295 ( .A(n5346), .B(n5347), .X(n6942) );
  nand_x1_sg U6296 ( .A(n8151), .B(n8132), .X(n5347) );
  nand_x1_sg U6297 ( .A(n5879), .B(n5880), .X(n7197) );
  nand_x1_sg U6298 ( .A(n8163), .B(n8132), .X(n5880) );
  nand_x1_sg U6299 ( .A(n5985), .B(n5986), .X(n7245) );
  nand_x1_sg U6300 ( .A(n8166), .B(n8132), .X(n5986) );
  nand_x1_sg U6301 ( .A(n5916), .B(n5917), .X(n7215) );
  nand_x1_sg U6302 ( .A(n8164), .B(n8132), .X(n5917) );
  nand_x1_sg U6303 ( .A(n5955), .B(n5956), .X(n7234) );
  nand_x1_sg U6304 ( .A(n8165), .B(n8132), .X(n5956) );
  nand_x1_sg U6305 ( .A(n5096), .B(n5097), .X(n6856) );
  nand_x1_sg U6306 ( .A(n8132), .B(n8155), .X(n5097) );
  nand_x1_sg U6307 ( .A(n5495), .B(n5496), .X(n7013) );
  nand_x1_sg U6308 ( .A(n8156), .B(n8132), .X(n5496) );
  nand_x1_sg U6309 ( .A(n5533), .B(n5534), .X(n7032) );
  nand_x1_sg U6310 ( .A(n8157), .B(n8132), .X(n5534) );
  nand_x1_sg U6311 ( .A(n5561), .B(n5562), .X(n7046) );
  nand_x1_sg U6312 ( .A(n8158), .B(n8132), .X(n5562) );
  nand_x1_sg U6313 ( .A(n5157), .B(n5158), .X(n6885) );
  nand_x1_sg U6314 ( .A(n8107), .B(n8132), .X(n5158) );
  nand_x1_sg U6315 ( .A(n5844), .B(n5845), .X(n7181) );
  nand_x1_sg U6316 ( .A(n8110), .B(n8132), .X(n5845) );
  nand_x1_sg U6317 ( .A(n5788), .B(n5789), .X(n7153) );
  nand_x1_sg U6318 ( .A(n8109), .B(n4870), .X(n5789) );
  nand_x1_sg U6319 ( .A(n5772), .B(n5773), .X(n7145) );
  nand_x1_sg U6320 ( .A(n8108), .B(n8132), .X(n5773) );
  nand_x1_sg U6321 ( .A(n5625), .B(n5626), .X(n7073) );
  nand_x1_sg U6322 ( .A(n8159), .B(n8132), .X(n5626) );
  nand_x1_sg U6323 ( .A(n5676), .B(n5677), .X(n7098) );
  nand_x1_sg U6324 ( .A(n8161), .B(n8132), .X(n5677) );
  nand_x1_sg U6325 ( .A(n5662), .B(n5663), .X(n7091) );
  nand_x1_sg U6326 ( .A(n8160), .B(n8132), .X(n5663) );
  nand_x1_sg U6327 ( .A(n5732), .B(n5733), .X(n7126) );
  nand_x1_sg U6328 ( .A(n8162), .B(n8132), .X(n5733) );
  nand_x1_sg U6329 ( .A(n5358), .B(n5359), .X(n6947) );
  nand_x1_sg U6330 ( .A(n8152), .B(n8132), .X(n5359) );
  nand_x1_sg U6331 ( .A(n5400), .B(n5401), .X(n6968) );
  nand_x1_sg U6332 ( .A(n8153), .B(n8146), .X(n5401) );
  nand_x1_sg U6333 ( .A(n5455), .B(n5456), .X(n6995) );
  nand_x1_sg U6334 ( .A(n8154), .B(n8146), .X(n5456) );
  nand_x1_sg U6335 ( .A(n5324), .B(n5325), .X(n6931) );
  nand_x1_sg U6336 ( .A(n8151), .B(n8146), .X(n5325) );
  nand_x1_sg U6337 ( .A(n5865), .B(n5866), .X(n7190) );
  nand_x1_sg U6338 ( .A(n8163), .B(n8146), .X(n5866) );
  nand_x1_sg U6339 ( .A(n6006), .B(n6007), .X(n7252) );
  nand_x1_sg U6340 ( .A(n8166), .B(n8146), .X(n6007) );
  nand_x1_sg U6341 ( .A(n5902), .B(n5903), .X(n7208) );
  nand_x1_sg U6342 ( .A(n8164), .B(n8146), .X(n5903) );
  nand_x1_sg U6343 ( .A(n5939), .B(n5940), .X(n7226) );
  nand_x1_sg U6344 ( .A(n8165), .B(n8146), .X(n5940) );
  nand_x1_sg U6345 ( .A(n5114), .B(n5115), .X(n6865) );
  nand_x1_sg U6346 ( .A(n8146), .B(n8155), .X(n5115) );
  nand_x1_sg U6347 ( .A(n5477), .B(n5478), .X(n7004) );
  nand_x1_sg U6348 ( .A(n8156), .B(n8146), .X(n5478) );
  nand_x1_sg U6349 ( .A(n5515), .B(n5516), .X(n7023) );
  nand_x1_sg U6350 ( .A(n8157), .B(n8146), .X(n5516) );
  nand_x1_sg U6351 ( .A(n5537), .B(n5538), .X(n7034) );
  nand_x1_sg U6352 ( .A(n8158), .B(n8146), .X(n5538) );
  nand_x1_sg U6353 ( .A(n5137), .B(n5138), .X(n6875) );
  nand_x1_sg U6354 ( .A(n8107), .B(n8146), .X(n5138) );
  nand_x1_sg U6355 ( .A(n5826), .B(n5827), .X(n7172) );
  nand_x1_sg U6356 ( .A(n8110), .B(n8146), .X(n5827) );
  nand_x1_sg U6357 ( .A(n5806), .B(n5807), .X(n7162) );
  nand_x1_sg U6358 ( .A(n8109), .B(n8146), .X(n5807) );
  nand_x1_sg U6359 ( .A(n5754), .B(n5755), .X(n7136) );
  nand_x1_sg U6360 ( .A(n8108), .B(n8146), .X(n5755) );
  nand_x1_sg U6361 ( .A(n5603), .B(n5604), .X(n7062) );
  nand_x1_sg U6362 ( .A(n8159), .B(n8146), .X(n5604) );
  nand_x1_sg U6363 ( .A(n5696), .B(n5697), .X(n7108) );
  nand_x1_sg U6364 ( .A(n8161), .B(n4863), .X(n5697) );
  nand_x1_sg U6365 ( .A(n5644), .B(n5645), .X(n7082) );
  nand_x1_sg U6366 ( .A(n8160), .B(n8146), .X(n5645) );
  nand_x1_sg U6367 ( .A(n5716), .B(n5717), .X(n7118) );
  nand_x1_sg U6368 ( .A(n8162), .B(n8146), .X(n5717) );
  nand_x1_sg U6369 ( .A(n5368), .B(n5369), .X(n6952) );
  nand_x1_sg U6370 ( .A(n8152), .B(n8146), .X(n5369) );
  nand_x1_sg U6371 ( .A(n5414), .B(n5415), .X(n6975) );
  nand_x1_sg U6372 ( .A(n8153), .B(n8150), .X(n5415) );
  nand_x1_sg U6373 ( .A(n5457), .B(n5458), .X(n6996) );
  nand_x1_sg U6374 ( .A(n8154), .B(n8150), .X(n5458) );
  nand_x1_sg U6375 ( .A(n5340), .B(n5341), .X(n6939) );
  nand_x1_sg U6376 ( .A(n8151), .B(n8150), .X(n5341) );
  nand_x1_sg U6377 ( .A(n5851), .B(n5852), .X(n7183) );
  nand_x1_sg U6378 ( .A(n8163), .B(n8150), .X(n5852) );
  nand_x1_sg U6379 ( .A(n6012), .B(n6013), .X(n7254) );
  nand_x1_sg U6380 ( .A(n8166), .B(n8150), .X(n6013) );
  nand_x1_sg U6381 ( .A(n5888), .B(n5889), .X(n7201) );
  nand_x1_sg U6382 ( .A(n8164), .B(n4861), .X(n5889) );
  nand_x1_sg U6383 ( .A(n5945), .B(n5946), .X(n7229) );
  nand_x1_sg U6384 ( .A(n8165), .B(n8150), .X(n5946) );
  nand_x1_sg U6385 ( .A(n5118), .B(n5119), .X(n6867) );
  nand_x1_sg U6386 ( .A(n8150), .B(n8155), .X(n5119) );
  nand_x1_sg U6387 ( .A(n5489), .B(n5490), .X(n7010) );
  nand_x1_sg U6388 ( .A(n8156), .B(n8150), .X(n5490) );
  nand_x1_sg U6389 ( .A(n5519), .B(n5520), .X(n7025) );
  nand_x1_sg U6390 ( .A(n8157), .B(n8150), .X(n5520) );
  nand_x1_sg U6391 ( .A(n5549), .B(n5550), .X(n7040) );
  nand_x1_sg U6392 ( .A(n8158), .B(n8150), .X(n5550) );
  nand_x1_sg U6393 ( .A(n5133), .B(n5134), .X(n6873) );
  nand_x1_sg U6394 ( .A(n8107), .B(n8150), .X(n5134) );
  nand_x1_sg U6395 ( .A(n5822), .B(n5823), .X(n7170) );
  nand_x1_sg U6396 ( .A(n8110), .B(n8150), .X(n5823) );
  nand_x1_sg U6397 ( .A(n5810), .B(n5811), .X(n7164) );
  nand_x1_sg U6398 ( .A(n8109), .B(n8150), .X(n5811) );
  nand_x1_sg U6399 ( .A(n5750), .B(n5751), .X(n7134) );
  nand_x1_sg U6400 ( .A(n8108), .B(n8150), .X(n5751) );
  nand_x1_sg U6401 ( .A(n5619), .B(n5620), .X(n7070) );
  nand_x1_sg U6402 ( .A(n8159), .B(n8150), .X(n5620) );
  nand_x1_sg U6403 ( .A(n5686), .B(n5687), .X(n7103) );
  nand_x1_sg U6404 ( .A(n8161), .B(n8150), .X(n5687) );
  nand_x1_sg U6405 ( .A(n5646), .B(n5647), .X(n7083) );
  nand_x1_sg U6406 ( .A(n8160), .B(n8150), .X(n5647) );
  nand_x1_sg U6407 ( .A(n5702), .B(n5703), .X(n7111) );
  nand_x1_sg U6408 ( .A(n8162), .B(n8150), .X(n5703) );
  nand_x1_sg U6409 ( .A(n5386), .B(n5387), .X(n6961) );
  nand_x1_sg U6410 ( .A(n8152), .B(n8150), .X(n5387) );
  nand_x1_sg U6411 ( .A(n5394), .B(n5395), .X(n6965) );
  nand_x1_sg U6412 ( .A(n8153), .B(n8118), .X(n5395) );
  nand_x1_sg U6413 ( .A(n5439), .B(n5440), .X(n6987) );
  nand_x1_sg U6414 ( .A(n8154), .B(n8118), .X(n5440) );
  nand_x1_sg U6415 ( .A(n5318), .B(n5319), .X(n6928) );
  nand_x1_sg U6416 ( .A(n8151), .B(n4877), .X(n5319) );
  nand_x1_sg U6417 ( .A(n5859), .B(n5860), .X(n7187) );
  nand_x1_sg U6418 ( .A(n8163), .B(n8118), .X(n5860) );
  nand_x1_sg U6419 ( .A(n5964), .B(n5965), .X(n7238) );
  nand_x1_sg U6420 ( .A(n8166), .B(n8118), .X(n5965) );
  nand_x1_sg U6421 ( .A(n5896), .B(n5897), .X(n7205) );
  nand_x1_sg U6422 ( .A(n8164), .B(n8118), .X(n5897) );
  nand_x1_sg U6423 ( .A(n5933), .B(n5934), .X(n7223) );
  nand_x1_sg U6424 ( .A(n8165), .B(n8118), .X(n5934) );
  nand_x1_sg U6425 ( .A(n5082), .B(n5083), .X(n6849) );
  nand_x1_sg U6426 ( .A(n8118), .B(n8155), .X(n5083) );
  nand_x1_sg U6427 ( .A(n5471), .B(n5472), .X(n7001) );
  nand_x1_sg U6428 ( .A(n8156), .B(n8118), .X(n5472) );
  nand_x1_sg U6429 ( .A(n5509), .B(n5510), .X(n7020) );
  nand_x1_sg U6430 ( .A(n8157), .B(n8118), .X(n5510) );
  nand_x1_sg U6431 ( .A(n5555), .B(n5556), .X(n7043) );
  nand_x1_sg U6432 ( .A(n8158), .B(n8118), .X(n5556) );
  nand_x1_sg U6433 ( .A(n5155), .B(n5156), .X(n6884) );
  nand_x1_sg U6434 ( .A(n8107), .B(n8118), .X(n5156) );
  nand_x1_sg U6435 ( .A(n5842), .B(n5843), .X(n7180) );
  nand_x1_sg U6436 ( .A(n8110), .B(n8118), .X(n5843) );
  nand_x1_sg U6437 ( .A(n5778), .B(n5779), .X(n7148) );
  nand_x1_sg U6438 ( .A(n8109), .B(n8118), .X(n5779) );
  nand_x1_sg U6439 ( .A(n5740), .B(n5741), .X(n7129) );
  nand_x1_sg U6440 ( .A(n8108), .B(n8118), .X(n5741) );
  nand_x1_sg U6441 ( .A(n5597), .B(n5598), .X(n7059) );
  nand_x1_sg U6442 ( .A(n8159), .B(n8118), .X(n5598) );
  nand_x1_sg U6443 ( .A(n5668), .B(n5669), .X(n7094) );
  nand_x1_sg U6444 ( .A(n8161), .B(n8118), .X(n5669) );
  nand_x1_sg U6445 ( .A(n5638), .B(n5639), .X(n7079) );
  nand_x1_sg U6446 ( .A(n8160), .B(n8118), .X(n5639) );
  nand_x1_sg U6447 ( .A(n5710), .B(n5711), .X(n7115) );
  nand_x1_sg U6448 ( .A(n8162), .B(n8118), .X(n5711) );
  nand_x1_sg U6449 ( .A(n5370), .B(n5371), .X(n6953) );
  nand_x1_sg U6450 ( .A(n8152), .B(n8118), .X(n5371) );
  nand_x1_sg U6451 ( .A(n5408), .B(n5409), .X(n6972) );
  nand_x1_sg U6452 ( .A(n8153), .B(n8130), .X(n5409) );
  nand_x1_sg U6453 ( .A(n5445), .B(n5446), .X(n6990) );
  nand_x1_sg U6454 ( .A(n8154), .B(n8130), .X(n5446) );
  nand_x1_sg U6455 ( .A(n5330), .B(n5331), .X(n6934) );
  nand_x1_sg U6456 ( .A(n8151), .B(n4871), .X(n5331) );
  nand_x1_sg U6457 ( .A(n5875), .B(n5876), .X(n7195) );
  nand_x1_sg U6458 ( .A(n8163), .B(n8130), .X(n5876) );
  nand_x1_sg U6459 ( .A(n5982), .B(n5983), .X(n7244) );
  nand_x1_sg U6460 ( .A(n8166), .B(n8130), .X(n5983) );
  nand_x1_sg U6461 ( .A(n5904), .B(n5905), .X(n7209) );
  nand_x1_sg U6462 ( .A(n8164), .B(n8130), .X(n5905) );
  nand_x1_sg U6463 ( .A(n5953), .B(n5954), .X(n7233) );
  nand_x1_sg U6464 ( .A(n8165), .B(n8130), .X(n5954) );
  nand_x1_sg U6465 ( .A(n5094), .B(n5095), .X(n6855) );
  nand_x1_sg U6466 ( .A(n8130), .B(n8155), .X(n5095) );
  nand_x1_sg U6467 ( .A(n5493), .B(n5494), .X(n7012) );
  nand_x1_sg U6468 ( .A(n8156), .B(n8130), .X(n5494) );
  nand_x1_sg U6469 ( .A(n5523), .B(n5524), .X(n7027) );
  nand_x1_sg U6470 ( .A(n8157), .B(n8130), .X(n5524) );
  nand_x1_sg U6471 ( .A(n5543), .B(n5544), .X(n7037) );
  nand_x1_sg U6472 ( .A(n8158), .B(n8130), .X(n5544) );
  nand_x1_sg U6473 ( .A(n5141), .B(n5142), .X(n6877) );
  nand_x1_sg U6474 ( .A(n8107), .B(n8130), .X(n5142) );
  nand_x1_sg U6475 ( .A(n5828), .B(n5829), .X(n7173) );
  nand_x1_sg U6476 ( .A(n8110), .B(n8130), .X(n5829) );
  nand_x1_sg U6477 ( .A(n5786), .B(n5787), .X(n7152) );
  nand_x1_sg U6478 ( .A(n8109), .B(n8130), .X(n5787) );
  nand_x1_sg U6479 ( .A(n5764), .B(n5765), .X(n7141) );
  nand_x1_sg U6480 ( .A(n8108), .B(n8130), .X(n5765) );
  nand_x1_sg U6481 ( .A(n5613), .B(n5614), .X(n7067) );
  nand_x1_sg U6482 ( .A(n8159), .B(n8130), .X(n5614) );
  nand_x1_sg U6483 ( .A(n5688), .B(n5689), .X(n7104) );
  nand_x1_sg U6484 ( .A(n8161), .B(n8130), .X(n5689) );
  nand_x1_sg U6485 ( .A(n5658), .B(n5659), .X(n7089) );
  nand_x1_sg U6486 ( .A(n8160), .B(n8130), .X(n5659) );
  nand_x1_sg U6487 ( .A(n5724), .B(n5725), .X(n7122) );
  nand_x1_sg U6488 ( .A(n8162), .B(n8130), .X(n5725) );
  nand_x1_sg U6489 ( .A(n5362), .B(n5363), .X(n6949) );
  nand_x1_sg U6490 ( .A(n8152), .B(n8130), .X(n5363) );
  nand_x1_sg U6491 ( .A(n5404), .B(n5405), .X(n6970) );
  nand_x1_sg U6492 ( .A(n8153), .B(n8142), .X(n5405) );
  nand_x1_sg U6493 ( .A(n5451), .B(n5452), .X(n6993) );
  nand_x1_sg U6494 ( .A(n8154), .B(n8142), .X(n5452) );
  nand_x1_sg U6495 ( .A(n5334), .B(n5335), .X(n6936) );
  nand_x1_sg U6496 ( .A(n8151), .B(n4865), .X(n5335) );
  nand_x1_sg U6497 ( .A(n5871), .B(n5872), .X(n7193) );
  nand_x1_sg U6498 ( .A(n8163), .B(n8142), .X(n5872) );
  nand_x1_sg U6499 ( .A(n6000), .B(n6001), .X(n7250) );
  nand_x1_sg U6500 ( .A(n8166), .B(n8142), .X(n6001) );
  nand_x1_sg U6501 ( .A(n5908), .B(n5909), .X(n7211) );
  nand_x1_sg U6502 ( .A(n8164), .B(n8142), .X(n5909) );
  nand_x1_sg U6503 ( .A(n5949), .B(n5950), .X(n7231) );
  nand_x1_sg U6504 ( .A(n8165), .B(n8142), .X(n5950) );
  nand_x1_sg U6505 ( .A(n5110), .B(n5111), .X(n6863) );
  nand_x1_sg U6506 ( .A(n8142), .B(n8155), .X(n5111) );
  nand_x1_sg U6507 ( .A(n5483), .B(n5484), .X(n7007) );
  nand_x1_sg U6508 ( .A(n8156), .B(n8142), .X(n5484) );
  nand_x1_sg U6509 ( .A(n5501), .B(n5502), .X(n7016) );
  nand_x1_sg U6510 ( .A(n8157), .B(n8142), .X(n5502) );
  nand_x1_sg U6511 ( .A(n5569), .B(n5570), .X(n7050) );
  nand_x1_sg U6512 ( .A(n8158), .B(n8142), .X(n5570) );
  nand_x1_sg U6513 ( .A(n5151), .B(n5152), .X(n6882) );
  nand_x1_sg U6514 ( .A(n8107), .B(n8142), .X(n5152) );
  nand_x1_sg U6515 ( .A(n5836), .B(n5837), .X(n7177) );
  nand_x1_sg U6516 ( .A(n8110), .B(n8142), .X(n5837) );
  nand_x1_sg U6517 ( .A(n5802), .B(n5803), .X(n7160) );
  nand_x1_sg U6518 ( .A(n8109), .B(n8142), .X(n5803) );
  nand_x1_sg U6519 ( .A(n5760), .B(n5761), .X(n7139) );
  nand_x1_sg U6520 ( .A(n8108), .B(n8142), .X(n5761) );
  nand_x1_sg U6521 ( .A(n5609), .B(n5610), .X(n7065) );
  nand_x1_sg U6522 ( .A(n8159), .B(n8142), .X(n5610) );
  nand_x1_sg U6523 ( .A(n5692), .B(n5693), .X(n7106) );
  nand_x1_sg U6524 ( .A(n8161), .B(n8142), .X(n5693) );
  nand_x1_sg U6525 ( .A(n5654), .B(n5655), .X(n7087) );
  nand_x1_sg U6526 ( .A(n8160), .B(n8142), .X(n5655) );
  nand_x1_sg U6527 ( .A(n5728), .B(n5729), .X(n7124) );
  nand_x1_sg U6528 ( .A(n8162), .B(n8142), .X(n5729) );
  nand_x1_sg U6529 ( .A(n5384), .B(n5385), .X(n6960) );
  nand_x1_sg U6530 ( .A(n8152), .B(n8142), .X(n5385) );
  nand_x1_sg U6531 ( .A(n5195), .B(n5196), .X(n6890) );
  nand_x1_sg U6532 ( .A(n8153), .B(n8112), .X(n5196) );
  nand_x1_sg U6533 ( .A(n5243), .B(n5244), .X(n6906) );
  nand_x1_sg U6534 ( .A(n8154), .B(n8112), .X(n5244) );
  nand_x1_sg U6535 ( .A(n5234), .B(n5235), .X(n6903) );
  nand_x1_sg U6536 ( .A(n8151), .B(n8112), .X(n5235) );
  nand_x1_sg U6537 ( .A(n5198), .B(n5199), .X(n6891) );
  nand_x1_sg U6538 ( .A(n8163), .B(n8112), .X(n5199) );
  nand_x1_sg U6539 ( .A(n5240), .B(n5241), .X(n6905) );
  nand_x1_sg U6540 ( .A(n8166), .B(n8112), .X(n5241) );
  nand_x1_sg U6541 ( .A(n5231), .B(n5232), .X(n6902) );
  nand_x1_sg U6542 ( .A(n8164), .B(n8112), .X(n5232) );
  nand_x1_sg U6543 ( .A(n5237), .B(n5238), .X(n6904) );
  nand_x1_sg U6544 ( .A(n8165), .B(n8112), .X(n5238) );
  nand_x1_sg U6545 ( .A(n5088), .B(n5089), .X(n6852) );
  nand_x1_sg U6546 ( .A(n8112), .B(n8155), .X(n5089) );
  nand_x1_sg U6547 ( .A(n5204), .B(n5205), .X(n6893) );
  nand_x1_sg U6548 ( .A(n8156), .B(n8112), .X(n5205) );
  nand_x1_sg U6549 ( .A(n5225), .B(n5226), .X(n6900) );
  nand_x1_sg U6550 ( .A(n8157), .B(n8112), .X(n5226) );
  nand_x1_sg U6551 ( .A(n5192), .B(n5193), .X(n6889) );
  nand_x1_sg U6552 ( .A(n8158), .B(n4880), .X(n5193) );
  nand_x1_sg U6553 ( .A(n5161), .B(n5162), .X(n6887) );
  nand_x1_sg U6554 ( .A(n8107), .B(n8112), .X(n5162) );
  nand_x1_sg U6555 ( .A(n5228), .B(n5229), .X(n6901) );
  nand_x1_sg U6556 ( .A(n8110), .B(n8112), .X(n5229) );
  nand_x1_sg U6557 ( .A(n5201), .B(n5202), .X(n6892) );
  nand_x1_sg U6558 ( .A(n8109), .B(n8112), .X(n5202) );
  nand_x1_sg U6559 ( .A(n5210), .B(n5211), .X(n6895) );
  nand_x1_sg U6560 ( .A(n8108), .B(n8112), .X(n5211) );
  nand_x1_sg U6561 ( .A(n5222), .B(n5223), .X(n6899) );
  nand_x1_sg U6562 ( .A(n8159), .B(n8112), .X(n5223) );
  nand_x1_sg U6563 ( .A(n5213), .B(n5214), .X(n6896) );
  nand_x1_sg U6564 ( .A(n8161), .B(n8112), .X(n5214) );
  nand_x1_sg U6565 ( .A(n5207), .B(n5208), .X(n6894) );
  nand_x1_sg U6566 ( .A(n8160), .B(n8112), .X(n5208) );
  nand_x1_sg U6567 ( .A(n5216), .B(n5217), .X(n6897) );
  nand_x1_sg U6568 ( .A(n8162), .B(n8112), .X(n5217) );
  nand_x1_sg U6569 ( .A(n5219), .B(n5220), .X(n6898) );
  nand_x1_sg U6570 ( .A(n8152), .B(n8112), .X(n5220) );
  nand_x1_sg U6571 ( .A(n5352), .B(n5353), .X(n6944) );
  nand_x1_sg U6572 ( .A(n8152), .B(n8124), .X(n5353) );
  nand_x1_sg U6573 ( .A(n5410), .B(n5411), .X(n6973) );
  nand_x1_sg U6574 ( .A(n8153), .B(n8124), .X(n5411) );
  nand_x1_sg U6575 ( .A(n5447), .B(n5448), .X(n6991) );
  nand_x1_sg U6576 ( .A(n8154), .B(n8124), .X(n5448) );
  nand_x1_sg U6577 ( .A(n5328), .B(n5329), .X(n6933) );
  nand_x1_sg U6578 ( .A(n8151), .B(n8124), .X(n5329) );
  nand_x1_sg U6579 ( .A(n5853), .B(n5854), .X(n7184) );
  nand_x1_sg U6580 ( .A(n8163), .B(n8124), .X(n5854) );
  nand_x1_sg U6581 ( .A(n5973), .B(n5974), .X(n7241) );
  nand_x1_sg U6582 ( .A(n8166), .B(n8124), .X(n5974) );
  nand_x1_sg U6583 ( .A(n5890), .B(n5891), .X(n7202) );
  nand_x1_sg U6584 ( .A(n8164), .B(n8124), .X(n5891) );
  nand_x1_sg U6585 ( .A(n5925), .B(n5926), .X(n7219) );
  nand_x1_sg U6586 ( .A(n8165), .B(n8124), .X(n5926) );
  nand_x1_sg U6587 ( .A(n5100), .B(n5101), .X(n6858) );
  nand_x1_sg U6588 ( .A(n8124), .B(n8155), .X(n5101) );
  nand_x1_sg U6589 ( .A(n5479), .B(n5480), .X(n7005) );
  nand_x1_sg U6590 ( .A(n8156), .B(n8124), .X(n5480) );
  nand_x1_sg U6591 ( .A(n5525), .B(n5526), .X(n7028) );
  nand_x1_sg U6592 ( .A(n8157), .B(n8124), .X(n5526) );
  nand_x1_sg U6593 ( .A(n5563), .B(n5564), .X(n7047) );
  nand_x1_sg U6594 ( .A(n8158), .B(n4874), .X(n5564) );
  nand_x1_sg U6595 ( .A(n5131), .B(n5132), .X(n6872) );
  nand_x1_sg U6596 ( .A(n8107), .B(n8124), .X(n5132) );
  nand_x1_sg U6597 ( .A(n5820), .B(n5821), .X(n7169) );
  nand_x1_sg U6598 ( .A(n8110), .B(n8124), .X(n5821) );
  nand_x1_sg U6599 ( .A(n5792), .B(n5793), .X(n7155) );
  nand_x1_sg U6600 ( .A(n8109), .B(n8124), .X(n5793) );
  nand_x1_sg U6601 ( .A(n5748), .B(n5749), .X(n7133) );
  nand_x1_sg U6602 ( .A(n8108), .B(n8124), .X(n5749) );
  nand_x1_sg U6603 ( .A(n5615), .B(n5616), .X(n7068) );
  nand_x1_sg U6604 ( .A(n8159), .B(n8124), .X(n5616) );
  nand_x1_sg U6605 ( .A(n5684), .B(n5685), .X(n7102) );
  nand_x1_sg U6606 ( .A(n8161), .B(n8124), .X(n5685) );
  nand_x1_sg U6607 ( .A(n5630), .B(n5631), .X(n7075) );
  nand_x1_sg U6608 ( .A(n8160), .B(n8124), .X(n5631) );
  nand_x1_sg U6609 ( .A(n5704), .B(n5705), .X(n7112) );
  nand_x1_sg U6610 ( .A(n8162), .B(n8124), .X(n5705) );
  nand_x1_sg U6611 ( .A(n5382), .B(n5383), .X(n6959) );
  nand_x1_sg U6612 ( .A(n8152), .B(n8134), .X(n5383) );
  nand_x1_sg U6613 ( .A(n5398), .B(n5399), .X(n6967) );
  nand_x1_sg U6614 ( .A(n8153), .B(n8134), .X(n5399) );
  nand_x1_sg U6615 ( .A(n5427), .B(n5428), .X(n6981) );
  nand_x1_sg U6616 ( .A(n8154), .B(n8134), .X(n5428) );
  nand_x1_sg U6617 ( .A(n5322), .B(n5323), .X(n6930) );
  nand_x1_sg U6618 ( .A(n8151), .B(n8134), .X(n5323) );
  nand_x1_sg U6619 ( .A(n5863), .B(n5864), .X(n7189) );
  nand_x1_sg U6620 ( .A(n8163), .B(n8134), .X(n5864) );
  nand_x1_sg U6621 ( .A(n5988), .B(n5989), .X(n7246) );
  nand_x1_sg U6622 ( .A(n8166), .B(n8134), .X(n5989) );
  nand_x1_sg U6623 ( .A(n5900), .B(n5901), .X(n7207) );
  nand_x1_sg U6624 ( .A(n8164), .B(n8134), .X(n5901) );
  nand_x1_sg U6625 ( .A(n5937), .B(n5938), .X(n7225) );
  nand_x1_sg U6626 ( .A(n8165), .B(n8134), .X(n5938) );
  nand_x1_sg U6627 ( .A(n5104), .B(n5105), .X(n6860) );
  nand_x1_sg U6628 ( .A(n8134), .B(n8155), .X(n5105) );
  nand_x1_sg U6629 ( .A(n5475), .B(n5476), .X(n7003) );
  nand_x1_sg U6630 ( .A(n8156), .B(n8134), .X(n5476) );
  nand_x1_sg U6631 ( .A(n5513), .B(n5514), .X(n7022) );
  nand_x1_sg U6632 ( .A(n8157), .B(n8134), .X(n5514) );
  nand_x1_sg U6633 ( .A(n5553), .B(n5554), .X(n7042) );
  nand_x1_sg U6634 ( .A(n8158), .B(n8134), .X(n5554) );
  nand_x1_sg U6635 ( .A(n5122), .B(n5123), .X(n6868) );
  nand_x1_sg U6636 ( .A(n8107), .B(n8134), .X(n5123) );
  nand_x1_sg U6637 ( .A(n5812), .B(n5813), .X(n7165) );
  nand_x1_sg U6638 ( .A(n8110), .B(n8134), .X(n5813) );
  nand_x1_sg U6639 ( .A(n5782), .B(n5783), .X(n7150) );
  nand_x1_sg U6640 ( .A(n8109), .B(n4869), .X(n5783) );
  nand_x1_sg U6641 ( .A(n5770), .B(n5771), .X(n7144) );
  nand_x1_sg U6642 ( .A(n8108), .B(n8134), .X(n5771) );
  nand_x1_sg U6643 ( .A(n5601), .B(n5602), .X(n7061) );
  nand_x1_sg U6644 ( .A(n8159), .B(n8134), .X(n5602) );
  nand_x1_sg U6645 ( .A(n5690), .B(n5691), .X(n7105) );
  nand_x1_sg U6646 ( .A(n8161), .B(n8134), .X(n5691) );
  nand_x1_sg U6647 ( .A(n5642), .B(n5643), .X(n7081) );
  nand_x1_sg U6648 ( .A(n8160), .B(n8134), .X(n5643) );
  nand_x1_sg U6649 ( .A(n5714), .B(n5715), .X(n7117) );
  nand_x1_sg U6650 ( .A(n8162), .B(n8134), .X(n5715) );
  nand_x1_sg U6651 ( .A(n5366), .B(n5367), .X(n6951) );
  nand_x1_sg U6652 ( .A(n8152), .B(n8136), .X(n5367) );
  nand_x1_sg U6653 ( .A(n5402), .B(n5403), .X(n6969) );
  nand_x1_sg U6654 ( .A(n8153), .B(n8136), .X(n5403) );
  nand_x1_sg U6655 ( .A(n5431), .B(n5432), .X(n6983) );
  nand_x1_sg U6656 ( .A(n8154), .B(n8136), .X(n5432) );
  nand_x1_sg U6657 ( .A(n5332), .B(n5333), .X(n6935) );
  nand_x1_sg U6658 ( .A(n8151), .B(n8136), .X(n5333) );
  nand_x1_sg U6659 ( .A(n5867), .B(n5868), .X(n7191) );
  nand_x1_sg U6660 ( .A(n8163), .B(n8136), .X(n5868) );
  nand_x1_sg U6661 ( .A(n5991), .B(n5992), .X(n7247) );
  nand_x1_sg U6662 ( .A(n8166), .B(n8136), .X(n5992) );
  nand_x1_sg U6663 ( .A(n5906), .B(n5907), .X(n7210) );
  nand_x1_sg U6664 ( .A(n8164), .B(n4868), .X(n5907) );
  nand_x1_sg U6665 ( .A(n5941), .B(n5942), .X(n7227) );
  nand_x1_sg U6666 ( .A(n8165), .B(n8136), .X(n5942) );
  nand_x1_sg U6667 ( .A(n5106), .B(n5107), .X(n6861) );
  nand_x1_sg U6668 ( .A(n8136), .B(n8155), .X(n5107) );
  nand_x1_sg U6669 ( .A(n5481), .B(n5482), .X(n7006) );
  nand_x1_sg U6670 ( .A(n8156), .B(n8136), .X(n5482) );
  nand_x1_sg U6671 ( .A(n5529), .B(n5530), .X(n7030) );
  nand_x1_sg U6672 ( .A(n8157), .B(n8136), .X(n5530) );
  nand_x1_sg U6673 ( .A(n5559), .B(n5560), .X(n7045) );
  nand_x1_sg U6674 ( .A(n8158), .B(n8136), .X(n5560) );
  nand_x1_sg U6675 ( .A(n5149), .B(n5150), .X(n6881) );
  nand_x1_sg U6676 ( .A(n8107), .B(n8136), .X(n5150) );
  nand_x1_sg U6677 ( .A(n5834), .B(n5835), .X(n7176) );
  nand_x1_sg U6678 ( .A(n8110), .B(n8136), .X(n5835) );
  nand_x1_sg U6679 ( .A(n5796), .B(n5797), .X(n7157) );
  nand_x1_sg U6680 ( .A(n8109), .B(n8136), .X(n5797) );
  nand_x1_sg U6681 ( .A(n5758), .B(n5759), .X(n7138) );
  nand_x1_sg U6682 ( .A(n8108), .B(n8136), .X(n5759) );
  nand_x1_sg U6683 ( .A(n5607), .B(n5608), .X(n7064) );
  nand_x1_sg U6684 ( .A(n8159), .B(n8136), .X(n5608) );
  nand_x1_sg U6685 ( .A(n5674), .B(n5675), .X(n7097) );
  nand_x1_sg U6686 ( .A(n8161), .B(n8136), .X(n5675) );
  nand_x1_sg U6687 ( .A(n5652), .B(n5653), .X(n7086) );
  nand_x1_sg U6688 ( .A(n8160), .B(n8136), .X(n5653) );
  nand_x1_sg U6689 ( .A(n5718), .B(n5719), .X(n7119) );
  nand_x1_sg U6690 ( .A(n8162), .B(n8136), .X(n5719) );
  nand_x1_sg U6691 ( .A(n5374), .B(n5375), .X(n6955) );
  nand_x1_sg U6692 ( .A(n8152), .B(n8144), .X(n5375) );
  nand_x1_sg U6693 ( .A(n5412), .B(n5413), .X(n6974) );
  nand_x1_sg U6694 ( .A(n8153), .B(n8144), .X(n5413) );
  nand_x1_sg U6695 ( .A(n5453), .B(n5454), .X(n6994) );
  nand_x1_sg U6696 ( .A(n8154), .B(n8144), .X(n5454) );
  nand_x1_sg U6697 ( .A(n5338), .B(n5339), .X(n6938) );
  nand_x1_sg U6698 ( .A(n8151), .B(n8144), .X(n5339) );
  nand_x1_sg U6699 ( .A(n5877), .B(n5878), .X(n7196) );
  nand_x1_sg U6700 ( .A(n8163), .B(n8144), .X(n5878) );
  nand_x1_sg U6701 ( .A(n6003), .B(n6004), .X(n7251) );
  nand_x1_sg U6702 ( .A(n8166), .B(n8144), .X(n6004) );
  nand_x1_sg U6703 ( .A(n5914), .B(n5915), .X(n7214) );
  nand_x1_sg U6704 ( .A(n8164), .B(n8144), .X(n5915) );
  nand_x1_sg U6705 ( .A(n5943), .B(n5944), .X(n7228) );
  nand_x1_sg U6706 ( .A(n8165), .B(n8144), .X(n5944) );
  nand_x1_sg U6707 ( .A(n5112), .B(n5113), .X(n6864) );
  nand_x1_sg U6708 ( .A(n8144), .B(n8155), .X(n5113) );
  nand_x1_sg U6709 ( .A(n5487), .B(n5488), .X(n7009) );
  nand_x1_sg U6710 ( .A(n8156), .B(n8144), .X(n5488) );
  nand_x1_sg U6711 ( .A(n5503), .B(n5504), .X(n7017) );
  nand_x1_sg U6712 ( .A(n8157), .B(n8144), .X(n5504) );
  nand_x1_sg U6713 ( .A(n5571), .B(n5572), .X(n7051) );
  nand_x1_sg U6714 ( .A(n8158), .B(n4864), .X(n5572) );
  nand_x1_sg U6715 ( .A(n5153), .B(n5154), .X(n6883) );
  nand_x1_sg U6716 ( .A(n8107), .B(n8144), .X(n5154) );
  nand_x1_sg U6717 ( .A(n5830), .B(n5831), .X(n7174) );
  nand_x1_sg U6718 ( .A(n8110), .B(n8144), .X(n5831) );
  nand_x1_sg U6719 ( .A(n5804), .B(n5805), .X(n7161) );
  nand_x1_sg U6720 ( .A(n8109), .B(n8144), .X(n5805) );
  nand_x1_sg U6721 ( .A(n5768), .B(n5769), .X(n7143) );
  nand_x1_sg U6722 ( .A(n8108), .B(n8144), .X(n5769) );
  nand_x1_sg U6723 ( .A(n5617), .B(n5618), .X(n7069) );
  nand_x1_sg U6724 ( .A(n8159), .B(n8144), .X(n5618) );
  nand_x1_sg U6725 ( .A(n5694), .B(n5695), .X(n7107) );
  nand_x1_sg U6726 ( .A(n8161), .B(n8144), .X(n5695) );
  nand_x1_sg U6727 ( .A(n5648), .B(n5649), .X(n7084) );
  nand_x1_sg U6728 ( .A(n8160), .B(n8144), .X(n5649) );
  nand_x1_sg U6729 ( .A(n5720), .B(n5721), .X(n7120) );
  nand_x1_sg U6730 ( .A(n8162), .B(n8144), .X(n5721) );
  nand_x1_sg U6731 ( .A(n5360), .B(n5361), .X(n6948) );
  nand_x1_sg U6732 ( .A(n8152), .B(n8128), .X(n5361) );
  nand_x1_sg U6733 ( .A(n5390), .B(n5391), .X(n6963) );
  nand_x1_sg U6734 ( .A(n8153), .B(n8128), .X(n5391) );
  nand_x1_sg U6735 ( .A(n5435), .B(n5436), .X(n6985) );
  nand_x1_sg U6736 ( .A(n8154), .B(n8128), .X(n5436) );
  nand_x1_sg U6737 ( .A(n5314), .B(n5315), .X(n6926) );
  nand_x1_sg U6738 ( .A(n8151), .B(n8128), .X(n5315) );
  nand_x1_sg U6739 ( .A(n5883), .B(n5884), .X(n7199) );
  nand_x1_sg U6740 ( .A(n8163), .B(n8128), .X(n5884) );
  nand_x1_sg U6741 ( .A(n5979), .B(n5980), .X(n7243) );
  nand_x1_sg U6742 ( .A(n8166), .B(n8128), .X(n5980) );
  nand_x1_sg U6743 ( .A(n5920), .B(n5921), .X(n7217) );
  nand_x1_sg U6744 ( .A(n8164), .B(n8128), .X(n5921) );
  nand_x1_sg U6745 ( .A(n5959), .B(n5960), .X(n7236) );
  nand_x1_sg U6746 ( .A(n8165), .B(n8128), .X(n5960) );
  nand_x1_sg U6747 ( .A(n5092), .B(n5093), .X(n6854) );
  nand_x1_sg U6748 ( .A(n8128), .B(n8155), .X(n5093) );
  nand_x1_sg U6749 ( .A(n5467), .B(n5468), .X(n6999) );
  nand_x1_sg U6750 ( .A(n8156), .B(n8128), .X(n5468) );
  nand_x1_sg U6751 ( .A(n5535), .B(n5536), .X(n7033) );
  nand_x1_sg U6752 ( .A(n8157), .B(n8128), .X(n5536) );
  nand_x1_sg U6753 ( .A(n5539), .B(n5540), .X(n7035) );
  nand_x1_sg U6754 ( .A(n8158), .B(n8128), .X(n5540) );
  nand_x1_sg U6755 ( .A(n5159), .B(n5160), .X(n6886) );
  nand_x1_sg U6756 ( .A(n8107), .B(n8128), .X(n5160) );
  nand_x1_sg U6757 ( .A(n5846), .B(n5847), .X(n7182) );
  nand_x1_sg U6758 ( .A(n8110), .B(n8128), .X(n5847) );
  nand_x1_sg U6759 ( .A(n5800), .B(n5801), .X(n7159) );
  nand_x1_sg U6760 ( .A(n8109), .B(n4872), .X(n5801) );
  nand_x1_sg U6761 ( .A(n5774), .B(n5775), .X(n7146) );
  nand_x1_sg U6762 ( .A(n8108), .B(n8128), .X(n5775) );
  nand_x1_sg U6763 ( .A(n5593), .B(n5594), .X(n7057) );
  nand_x1_sg U6764 ( .A(n8159), .B(n8128), .X(n5594) );
  nand_x1_sg U6765 ( .A(n5680), .B(n5681), .X(n7100) );
  nand_x1_sg U6766 ( .A(n8161), .B(n8128), .X(n5681) );
  nand_x1_sg U6767 ( .A(n5664), .B(n5665), .X(n7092) );
  nand_x1_sg U6768 ( .A(n8160), .B(n8128), .X(n5665) );
  nand_x1_sg U6769 ( .A(n5736), .B(n5737), .X(n7128) );
  nand_x1_sg U6770 ( .A(n8162), .B(n8128), .X(n5737) );
  nand_x1_sg U6771 ( .A(n5376), .B(n5377), .X(n6956) );
  nand_x1_sg U6772 ( .A(n8152), .B(n8116), .X(n5377) );
  nand_x1_sg U6773 ( .A(n5392), .B(n5393), .X(n6964) );
  nand_x1_sg U6774 ( .A(n8153), .B(n8116), .X(n5393) );
  nand_x1_sg U6775 ( .A(n5443), .B(n5444), .X(n6989) );
  nand_x1_sg U6776 ( .A(n8154), .B(n8116), .X(n5444) );
  nand_x1_sg U6777 ( .A(n5316), .B(n5317), .X(n6927) );
  nand_x1_sg U6778 ( .A(n8151), .B(n8116), .X(n5317) );
  nand_x1_sg U6779 ( .A(n5857), .B(n5858), .X(n7186) );
  nand_x1_sg U6780 ( .A(n8163), .B(n8116), .X(n5858) );
  nand_x1_sg U6781 ( .A(n5961), .B(n5962), .X(n7237) );
  nand_x1_sg U6782 ( .A(n8166), .B(n8116), .X(n5962) );
  nand_x1_sg U6783 ( .A(n5894), .B(n5895), .X(n7204) );
  nand_x1_sg U6784 ( .A(n8164), .B(n8116), .X(n5895) );
  nand_x1_sg U6785 ( .A(n5931), .B(n5932), .X(n7222) );
  nand_x1_sg U6786 ( .A(n8165), .B(n8116), .X(n5932) );
  nand_x1_sg U6787 ( .A(n5079), .B(n5080), .X(n6848) );
  nand_x1_sg U6788 ( .A(n8116), .B(n8155), .X(n5080) );
  nand_x1_sg U6789 ( .A(n5469), .B(n5470), .X(n7000) );
  nand_x1_sg U6790 ( .A(n8156), .B(n8116), .X(n5470) );
  nand_x1_sg U6791 ( .A(n5507), .B(n5508), .X(n7019) );
  nand_x1_sg U6792 ( .A(n8157), .B(n8116), .X(n5508) );
  nand_x1_sg U6793 ( .A(n5551), .B(n5552), .X(n7041) );
  nand_x1_sg U6794 ( .A(n8158), .B(n8116), .X(n5552) );
  nand_x1_sg U6795 ( .A(n5129), .B(n5130), .X(n6871) );
  nand_x1_sg U6796 ( .A(n8107), .B(n8116), .X(n5130) );
  nand_x1_sg U6797 ( .A(n5818), .B(n5819), .X(n7168) );
  nand_x1_sg U6798 ( .A(n8110), .B(n8116), .X(n5819) );
  nand_x1_sg U6799 ( .A(n5776), .B(n5777), .X(n7147) );
  nand_x1_sg U6800 ( .A(n8109), .B(n4878), .X(n5777) );
  nand_x1_sg U6801 ( .A(n5746), .B(n5747), .X(n7132) );
  nand_x1_sg U6802 ( .A(n8108), .B(n8116), .X(n5747) );
  nand_x1_sg U6803 ( .A(n5595), .B(n5596), .X(n7058) );
  nand_x1_sg U6804 ( .A(n8159), .B(n8116), .X(n5596) );
  nand_x1_sg U6805 ( .A(n5666), .B(n5667), .X(n7093) );
  nand_x1_sg U6806 ( .A(n8161), .B(n8116), .X(n5667) );
  nand_x1_sg U6807 ( .A(n5636), .B(n5637), .X(n7078) );
  nand_x1_sg U6808 ( .A(n8160), .B(n8116), .X(n5637) );
  nand_x1_sg U6809 ( .A(n5708), .B(n5709), .X(n7114) );
  nand_x1_sg U6810 ( .A(n8162), .B(n8116), .X(n5709) );
  nand_x1_sg U6811 ( .A(n5380), .B(n5381), .X(n6958) );
  nand_x1_sg U6812 ( .A(n8152), .B(n8138), .X(n5381) );
  nand_x1_sg U6813 ( .A(n5406), .B(n5407), .X(n6971) );
  nand_x1_sg U6814 ( .A(n8153), .B(n8138), .X(n5407) );
  nand_x1_sg U6815 ( .A(n5429), .B(n5430), .X(n6982) );
  nand_x1_sg U6816 ( .A(n8154), .B(n8138), .X(n5430) );
  nand_x1_sg U6817 ( .A(n5336), .B(n5337), .X(n6937) );
  nand_x1_sg U6818 ( .A(n8151), .B(n8138), .X(n5337) );
  nand_x1_sg U6819 ( .A(n5873), .B(n5874), .X(n7194) );
  nand_x1_sg U6820 ( .A(n8163), .B(n8138), .X(n5874) );
  nand_x1_sg U6821 ( .A(n5994), .B(n5995), .X(n7248) );
  nand_x1_sg U6822 ( .A(n8166), .B(n8138), .X(n5995) );
  nand_x1_sg U6823 ( .A(n5910), .B(n5911), .X(n7212) );
  nand_x1_sg U6824 ( .A(n8164), .B(n8138), .X(n5911) );
  nand_x1_sg U6825 ( .A(n5951), .B(n5952), .X(n7232) );
  nand_x1_sg U6826 ( .A(n8165), .B(n8138), .X(n5952) );
  nand_x1_sg U6827 ( .A(n5086), .B(n5087), .X(n6851) );
  nand_x1_sg U6828 ( .A(n8138), .B(n8155), .X(n5087) );
  nand_x1_sg U6829 ( .A(n5485), .B(n5486), .X(n7008) );
  nand_x1_sg U6830 ( .A(n8156), .B(n8138), .X(n5486) );
  nand_x1_sg U6831 ( .A(n5531), .B(n5532), .X(n7031) );
  nand_x1_sg U6832 ( .A(n8157), .B(n8138), .X(n5532) );
  nand_x1_sg U6833 ( .A(n5557), .B(n5558), .X(n7044) );
  nand_x1_sg U6834 ( .A(n8158), .B(n4867), .X(n5558) );
  nand_x1_sg U6835 ( .A(n5125), .B(n5126), .X(n6869) );
  nand_x1_sg U6836 ( .A(n8107), .B(n8138), .X(n5126) );
  nand_x1_sg U6837 ( .A(n5814), .B(n5815), .X(n7166) );
  nand_x1_sg U6838 ( .A(n8110), .B(n8138), .X(n5815) );
  nand_x1_sg U6839 ( .A(n5798), .B(n5799), .X(n7158) );
  nand_x1_sg U6840 ( .A(n8109), .B(n8138), .X(n5799) );
  nand_x1_sg U6841 ( .A(n5742), .B(n5743), .X(n7130) );
  nand_x1_sg U6842 ( .A(n8108), .B(n8138), .X(n5743) );
  nand_x1_sg U6843 ( .A(n5611), .B(n5612), .X(n7066) );
  nand_x1_sg U6844 ( .A(n8159), .B(n8138), .X(n5612) );
  nand_x1_sg U6845 ( .A(n5678), .B(n5679), .X(n7099) );
  nand_x1_sg U6846 ( .A(n8161), .B(n8138), .X(n5679) );
  nand_x1_sg U6847 ( .A(n5656), .B(n5657), .X(n7088) );
  nand_x1_sg U6848 ( .A(n8160), .B(n8138), .X(n5657) );
  nand_x1_sg U6849 ( .A(n5730), .B(n5731), .X(n7125) );
  nand_x1_sg U6850 ( .A(n8162), .B(n8138), .X(n5731) );
  nand_x1_sg U6851 ( .A(n5356), .B(n5357), .X(n6946) );
  nand_x1_sg U6852 ( .A(n8152), .B(n8126), .X(n5357) );
  nand_x1_sg U6853 ( .A(n5422), .B(n5423), .X(n6979) );
  nand_x1_sg U6854 ( .A(n8153), .B(n8126), .X(n5423) );
  nand_x1_sg U6855 ( .A(n5459), .B(n5460), .X(n6997) );
  nand_x1_sg U6856 ( .A(n8154), .B(n8126), .X(n5460) );
  nand_x1_sg U6857 ( .A(n5348), .B(n5349), .X(n6943) );
  nand_x1_sg U6858 ( .A(n8151), .B(n8126), .X(n5349) );
  nand_x1_sg U6859 ( .A(n5881), .B(n5882), .X(n7198) );
  nand_x1_sg U6860 ( .A(n8163), .B(n8126), .X(n5882) );
  nand_x1_sg U6861 ( .A(n5976), .B(n5977), .X(n7242) );
  nand_x1_sg U6862 ( .A(n8166), .B(n8126), .X(n5977) );
  nand_x1_sg U6863 ( .A(n5918), .B(n5919), .X(n7216) );
  nand_x1_sg U6864 ( .A(n8164), .B(n4873), .X(n5919) );
  nand_x1_sg U6865 ( .A(n5927), .B(n5928), .X(n7220) );
  nand_x1_sg U6866 ( .A(n8165), .B(n8126), .X(n5928) );
  nand_x1_sg U6867 ( .A(n5102), .B(n5103), .X(n6859) );
  nand_x1_sg U6868 ( .A(n8126), .B(n8155), .X(n5103) );
  nand_x1_sg U6869 ( .A(n5497), .B(n5498), .X(n7014) );
  nand_x1_sg U6870 ( .A(n8156), .B(n8126), .X(n5498) );
  nand_x1_sg U6871 ( .A(n5517), .B(n5518), .X(n7024) );
  nand_x1_sg U6872 ( .A(n8157), .B(n8126), .X(n5518) );
  nand_x1_sg U6873 ( .A(n5565), .B(n5566), .X(n7048) );
  nand_x1_sg U6874 ( .A(n8158), .B(n8126), .X(n5566) );
  nand_x1_sg U6875 ( .A(n5139), .B(n5140), .X(n6876) );
  nand_x1_sg U6876 ( .A(n8107), .B(n8126), .X(n5140) );
  nand_x1_sg U6877 ( .A(n5840), .B(n5841), .X(n7179) );
  nand_x1_sg U6878 ( .A(n8110), .B(n8126), .X(n5841) );
  nand_x1_sg U6879 ( .A(n5794), .B(n5795), .X(n7156) );
  nand_x1_sg U6880 ( .A(n8109), .B(n8126), .X(n5795) );
  nand_x1_sg U6881 ( .A(n5756), .B(n5757), .X(n7137) );
  nand_x1_sg U6882 ( .A(n8108), .B(n8126), .X(n5757) );
  nand_x1_sg U6883 ( .A(n5627), .B(n5628), .X(n7074) );
  nand_x1_sg U6884 ( .A(n8159), .B(n8126), .X(n5628) );
  nand_x1_sg U6885 ( .A(n5700), .B(n5701), .X(n7110) );
  nand_x1_sg U6886 ( .A(n8161), .B(n8126), .X(n5701) );
  nand_x1_sg U6887 ( .A(n5632), .B(n5633), .X(n7076) );
  nand_x1_sg U6888 ( .A(n8160), .B(n8126), .X(n5633) );
  nand_x1_sg U6889 ( .A(n5706), .B(n5707), .X(n7113) );
  nand_x1_sg U6890 ( .A(n8162), .B(n8126), .X(n5707) );
  nand_x1_sg U6891 ( .A(n5589), .B(n5590), .X(n7056) );
  nand_x1_sg U6892 ( .A(n8259), .B(n5188), .X(n5589) );
  nand_x1_sg U6893 ( .A(n5584), .B(n5585), .X(n7055) );
  nand_x1_sg U6894 ( .A(n5581), .B(n5582), .X(n7054) );
  nand_x1_sg U6895 ( .A(n5577), .B(n5578), .X(n7053) );
  nand_x1_sg U6896 ( .A(n5575), .B(n5576), .X(n7052) );
  nand_x1_sg U6897 ( .A(n5164), .B(n5165), .X(n6888) );
  nand_x1_sg U6898 ( .A(n8259), .B(n5166), .X(n5164) );
  nand_x1_sg U6899 ( .A(n6027), .B(n6028), .X(n7257) );
  inv_x4_sg U6900 ( .A(n5996), .X(n4867) );
  inv_x4_sg U6901 ( .A(n6005), .X(n4864) );
  nor_x2_sg U6902 ( .A(n7333), .B(n5185), .X(n5184) );
  nand_x2_sg U6903 ( .A(n5574), .B(n8106), .X(n5573) );
  inv_x4_sg U6904 ( .A(n5978), .X(n4873) );
  inv_x4_sg U6905 ( .A(n5993), .X(n4868) );
  nor_x2_sg U6906 ( .A(n4905), .B(n5078), .X(n5183) );
  nand_x2_sg U6907 ( .A(n6016), .B(n8106), .X(n6015) );
  inv_x4_sg U6908 ( .A(n5963), .X(n4878) );
  inv_x4_sg U6909 ( .A(n5990), .X(n4869) );
  nor_x2_sg U6910 ( .A(n7340), .B(n4903), .X(n5187) );
  nand_x2_sg U6911 ( .A(n5463), .B(n7338), .X(n5462) );
  inv_x4_sg U6912 ( .A(n5981), .X(n4872) );
  inv_x4_sg U6913 ( .A(n6002), .X(n4865) );
  inv_x1_sg U6914 ( .A(n5166), .X(n4881) );
  nor_x1_sg U6915 ( .A(n5271), .B(n5272), .X(n5266) );
  nor_x2_sg U6916 ( .A(n4909), .B(n5273), .X(n5271) );
  nor_x2_sg U6917 ( .A(n7338), .B(n4892), .X(n5272) );
  inv_x4_sg U6918 ( .A(n5975), .X(n4874) );
  inv_x4_sg U6919 ( .A(n5984), .X(n4871) );
  nor_x2_sg U6920 ( .A(empty), .B(n4889), .X(n6019) );
  inv_x4_sg U6921 ( .A(n5966), .X(n4877) );
  inv_x4_sg U6922 ( .A(n6008), .X(n4863) );
  nor_x2_sg U6923 ( .A(n8106), .B(n7338), .X(n5739) );
  inv_x4_sg U6924 ( .A(n7261), .X(n7332) );
  inv_x8_sg U6925 ( .A(n7332), .X(n7333) );
  inv_x8_sg U6926 ( .A(n6814), .X(n4898) );
  inv_x8_sg U6927 ( .A(n6811), .X(n4891) );
  inv_x8_sg U6928 ( .A(n5077), .X(n7334) );
  inv_x4_sg U6929 ( .A(n7335), .X(n7336) );
  inv_x8_sg U6930 ( .A(n7336), .X(n5077) );
  nor_x2_sg U6931 ( .A(n5073), .B(n5188), .X(n5186) );
  inv_x4_sg U6932 ( .A(n7331), .X(n4902) );
  inv_x4_sg U6933 ( .A(n5185), .X(n4905) );
  nand_x4_sg U6934 ( .A(n5586), .B(n5587), .X(n5185) );
  inv_x2_sg U6935 ( .A(\buff_mem[10][12] ), .X(n7781) );
  inv_x2_sg U6936 ( .A(\buff_mem[8][12] ), .X(n7783) );
  inv_x2_sg U6937 ( .A(\buff_mem[10][13] ), .X(n7785) );
  inv_x2_sg U6938 ( .A(\buff_mem[8][13] ), .X(n7787) );
  inv_x2_sg U6939 ( .A(\buff_mem[10][14] ), .X(n7789) );
  inv_x2_sg U6940 ( .A(\buff_mem[8][14] ), .X(n7791) );
  inv_x2_sg U6941 ( .A(\buff_mem[10][15] ), .X(n7793) );
  inv_x2_sg U6942 ( .A(\buff_mem[8][15] ), .X(n7795) );
  inv_x2_sg U6943 ( .A(\buff_mem[10][16] ), .X(n7797) );
  inv_x2_sg U6944 ( .A(\buff_mem[8][16] ), .X(n7799) );
  inv_x2_sg U6945 ( .A(\buff_mem[10][17] ), .X(n7801) );
  inv_x2_sg U6946 ( .A(\buff_mem[8][17] ), .X(n7803) );
  inv_x2_sg U6947 ( .A(\buff_mem[10][18] ), .X(n7805) );
  inv_x2_sg U6948 ( .A(\buff_mem[8][18] ), .X(n7807) );
  inv_x2_sg U6949 ( .A(\buff_mem[10][19] ), .X(n7809) );
  inv_x2_sg U6950 ( .A(\buff_mem[8][19] ), .X(n7811) );
  inv_x2_sg U6951 ( .A(\buff_mem[10][0] ), .X(n7813) );
  inv_x2_sg U6952 ( .A(\buff_mem[8][0] ), .X(n7815) );
  inv_x2_sg U6953 ( .A(\buff_mem[10][1] ), .X(n7817) );
  inv_x2_sg U6954 ( .A(\buff_mem[8][1] ), .X(n7819) );
  inv_x2_sg U6955 ( .A(\buff_mem[10][2] ), .X(n7821) );
  inv_x2_sg U6956 ( .A(\buff_mem[8][2] ), .X(n7823) );
  inv_x2_sg U6957 ( .A(\buff_mem[10][3] ), .X(n7825) );
  inv_x2_sg U6958 ( .A(\buff_mem[8][3] ), .X(n7827) );
  inv_x2_sg U6959 ( .A(\buff_mem[10][4] ), .X(n7829) );
  inv_x2_sg U6960 ( .A(\buff_mem[8][4] ), .X(n7831) );
  inv_x2_sg U6961 ( .A(\buff_mem[10][5] ), .X(n7833) );
  inv_x2_sg U6962 ( .A(\buff_mem[8][5] ), .X(n7835) );
  inv_x2_sg U6963 ( .A(\buff_mem[10][6] ), .X(n7837) );
  inv_x2_sg U6964 ( .A(\buff_mem[8][6] ), .X(n7839) );
  inv_x2_sg U6965 ( .A(\buff_mem[10][7] ), .X(n7841) );
  inv_x2_sg U6966 ( .A(\buff_mem[8][7] ), .X(n7843) );
  inv_x2_sg U6967 ( .A(\buff_mem[10][8] ), .X(n7845) );
  inv_x2_sg U6968 ( .A(\buff_mem[8][8] ), .X(n7847) );
  inv_x2_sg U6969 ( .A(\buff_mem[10][9] ), .X(n7849) );
  inv_x2_sg U6970 ( .A(\buff_mem[8][9] ), .X(n7851) );
  inv_x2_sg U6971 ( .A(\buff_mem[10][10] ), .X(n7853) );
  inv_x2_sg U6972 ( .A(\buff_mem[8][10] ), .X(n7855) );
  inv_x2_sg U6973 ( .A(\buff_mem[10][11] ), .X(n7857) );
  inv_x2_sg U6974 ( .A(\buff_mem[8][11] ), .X(n7859) );
  inv_x2_sg U6975 ( .A(\buff_mem[13][12] ), .X(n7861) );
  inv_x2_sg U6976 ( .A(\buff_mem[9][12] ), .X(n7863) );
  inv_x2_sg U6977 ( .A(\buff_mem[13][13] ), .X(n7865) );
  inv_x2_sg U6978 ( .A(\buff_mem[9][13] ), .X(n7867) );
  inv_x2_sg U6979 ( .A(\buff_mem[13][14] ), .X(n7869) );
  inv_x2_sg U6980 ( .A(\buff_mem[9][14] ), .X(n7871) );
  inv_x2_sg U6981 ( .A(\buff_mem[13][15] ), .X(n7873) );
  inv_x2_sg U6982 ( .A(\buff_mem[9][15] ), .X(n7875) );
  inv_x2_sg U6983 ( .A(\buff_mem[13][16] ), .X(n7877) );
  inv_x2_sg U6984 ( .A(\buff_mem[9][16] ), .X(n7879) );
  inv_x2_sg U6985 ( .A(\buff_mem[13][17] ), .X(n7881) );
  inv_x2_sg U6986 ( .A(\buff_mem[9][17] ), .X(n7883) );
  inv_x2_sg U6987 ( .A(\buff_mem[13][18] ), .X(n7885) );
  inv_x2_sg U6988 ( .A(\buff_mem[9][18] ), .X(n7887) );
  inv_x2_sg U6989 ( .A(\buff_mem[13][19] ), .X(n7889) );
  inv_x2_sg U6990 ( .A(\buff_mem[9][19] ), .X(n7891) );
  inv_x2_sg U6991 ( .A(\buff_mem[13][0] ), .X(n7893) );
  inv_x2_sg U6992 ( .A(\buff_mem[9][0] ), .X(n7895) );
  inv_x2_sg U6993 ( .A(\buff_mem[13][1] ), .X(n7897) );
  inv_x2_sg U6994 ( .A(\buff_mem[9][1] ), .X(n7899) );
  inv_x2_sg U6995 ( .A(\buff_mem[13][2] ), .X(n7901) );
  inv_x2_sg U6996 ( .A(\buff_mem[9][2] ), .X(n7903) );
  inv_x2_sg U6997 ( .A(\buff_mem[13][3] ), .X(n7905) );
  inv_x2_sg U6998 ( .A(\buff_mem[9][3] ), .X(n7907) );
  inv_x2_sg U6999 ( .A(\buff_mem[13][4] ), .X(n7909) );
  inv_x2_sg U7000 ( .A(\buff_mem[9][4] ), .X(n7911) );
  inv_x2_sg U7001 ( .A(\buff_mem[13][5] ), .X(n7913) );
  inv_x2_sg U7002 ( .A(\buff_mem[9][5] ), .X(n7915) );
  inv_x2_sg U7003 ( .A(\buff_mem[13][6] ), .X(n7917) );
  inv_x2_sg U7004 ( .A(\buff_mem[9][6] ), .X(n7919) );
  inv_x2_sg U7005 ( .A(\buff_mem[13][7] ), .X(n7921) );
  inv_x2_sg U7006 ( .A(\buff_mem[9][7] ), .X(n7923) );
  inv_x2_sg U7007 ( .A(\buff_mem[13][8] ), .X(n7925) );
  inv_x2_sg U7008 ( .A(\buff_mem[9][8] ), .X(n7927) );
  inv_x2_sg U7009 ( .A(\buff_mem[13][9] ), .X(n7929) );
  inv_x2_sg U7010 ( .A(\buff_mem[9][9] ), .X(n7931) );
  inv_x2_sg U7011 ( .A(\buff_mem[13][10] ), .X(n7933) );
  inv_x2_sg U7012 ( .A(\buff_mem[9][10] ), .X(n7935) );
  inv_x2_sg U7013 ( .A(\buff_mem[13][11] ), .X(n7937) );
  inv_x2_sg U7014 ( .A(\buff_mem[9][11] ), .X(n7939) );
  inv_x2_sg U7015 ( .A(\buff_mem[16][12] ), .X(n7941) );
  inv_x2_sg U7016 ( .A(\buff_mem[14][12] ), .X(n7943) );
  inv_x2_sg U7017 ( .A(\buff_mem[16][13] ), .X(n7945) );
  inv_x2_sg U7018 ( .A(\buff_mem[14][13] ), .X(n7947) );
  inv_x2_sg U7019 ( .A(\buff_mem[16][14] ), .X(n7949) );
  inv_x2_sg U7020 ( .A(\buff_mem[14][14] ), .X(n7951) );
  inv_x2_sg U7021 ( .A(\buff_mem[16][15] ), .X(n7953) );
  inv_x2_sg U7022 ( .A(\buff_mem[14][15] ), .X(n7955) );
  inv_x2_sg U7023 ( .A(\buff_mem[16][16] ), .X(n7957) );
  inv_x2_sg U7024 ( .A(\buff_mem[14][16] ), .X(n7959) );
  inv_x2_sg U7025 ( .A(\buff_mem[16][17] ), .X(n7961) );
  inv_x2_sg U7026 ( .A(\buff_mem[14][17] ), .X(n7963) );
  inv_x2_sg U7027 ( .A(\buff_mem[16][18] ), .X(n7965) );
  inv_x2_sg U7028 ( .A(\buff_mem[14][18] ), .X(n7967) );
  inv_x2_sg U7029 ( .A(\buff_mem[16][19] ), .X(n7969) );
  inv_x2_sg U7030 ( .A(\buff_mem[14][19] ), .X(n7971) );
  inv_x2_sg U7031 ( .A(\buff_mem[16][0] ), .X(n7973) );
  inv_x2_sg U7032 ( .A(\buff_mem[14][0] ), .X(n7975) );
  inv_x2_sg U7033 ( .A(\buff_mem[16][1] ), .X(n7977) );
  inv_x2_sg U7034 ( .A(\buff_mem[14][1] ), .X(n7979) );
  inv_x2_sg U7035 ( .A(\buff_mem[16][2] ), .X(n7981) );
  inv_x2_sg U7036 ( .A(\buff_mem[14][2] ), .X(n7983) );
  inv_x2_sg U7037 ( .A(\buff_mem[16][3] ), .X(n7985) );
  inv_x2_sg U7038 ( .A(\buff_mem[14][3] ), .X(n7987) );
  inv_x2_sg U7039 ( .A(\buff_mem[16][4] ), .X(n7989) );
  inv_x2_sg U7040 ( .A(\buff_mem[14][4] ), .X(n7991) );
  inv_x2_sg U7041 ( .A(\buff_mem[16][5] ), .X(n7993) );
  inv_x2_sg U7042 ( .A(\buff_mem[14][5] ), .X(n7995) );
  inv_x2_sg U7043 ( .A(\buff_mem[16][6] ), .X(n7997) );
  inv_x2_sg U7044 ( .A(\buff_mem[14][6] ), .X(n7999) );
  inv_x2_sg U7045 ( .A(\buff_mem[16][7] ), .X(n8001) );
  inv_x2_sg U7046 ( .A(\buff_mem[14][7] ), .X(n8003) );
  inv_x2_sg U7047 ( .A(\buff_mem[16][8] ), .X(n8005) );
  inv_x2_sg U7048 ( .A(\buff_mem[14][8] ), .X(n8007) );
  inv_x2_sg U7049 ( .A(\buff_mem[16][9] ), .X(n8009) );
  inv_x2_sg U7050 ( .A(\buff_mem[14][9] ), .X(n8011) );
  inv_x2_sg U7051 ( .A(\buff_mem[16][10] ), .X(n8013) );
  inv_x2_sg U7052 ( .A(\buff_mem[14][10] ), .X(n8015) );
  inv_x2_sg U7053 ( .A(\buff_mem[16][11] ), .X(n8017) );
  inv_x2_sg U7054 ( .A(\buff_mem[14][11] ), .X(n8019) );
  inv_x2_sg U7055 ( .A(\buff_mem[3][12] ), .X(n8021) );
  inv_x2_sg U7056 ( .A(\buff_mem[12][12] ), .X(n8023) );
  inv_x2_sg U7057 ( .A(\buff_mem[3][13] ), .X(n8025) );
  inv_x2_sg U7058 ( .A(\buff_mem[12][13] ), .X(n8027) );
  inv_x2_sg U7059 ( .A(\buff_mem[3][14] ), .X(n8029) );
  inv_x2_sg U7060 ( .A(\buff_mem[12][14] ), .X(n8031) );
  inv_x2_sg U7061 ( .A(\buff_mem[3][15] ), .X(n8033) );
  inv_x2_sg U7062 ( .A(\buff_mem[12][15] ), .X(n8035) );
  inv_x2_sg U7063 ( .A(\buff_mem[3][16] ), .X(n8037) );
  inv_x2_sg U7064 ( .A(\buff_mem[12][16] ), .X(n8039) );
  inv_x2_sg U7065 ( .A(\buff_mem[3][17] ), .X(n8041) );
  inv_x2_sg U7066 ( .A(\buff_mem[12][17] ), .X(n8043) );
  inv_x2_sg U7067 ( .A(\buff_mem[3][18] ), .X(n8045) );
  inv_x2_sg U7068 ( .A(\buff_mem[12][18] ), .X(n8047) );
  inv_x2_sg U7069 ( .A(\buff_mem[3][19] ), .X(n8049) );
  inv_x2_sg U7070 ( .A(\buff_mem[12][19] ), .X(n8051) );
  inv_x2_sg U7071 ( .A(\buff_mem[3][0] ), .X(n8053) );
  inv_x2_sg U7072 ( .A(\buff_mem[12][0] ), .X(n8055) );
  inv_x2_sg U7073 ( .A(\buff_mem[3][1] ), .X(n8057) );
  inv_x2_sg U7074 ( .A(\buff_mem[12][1] ), .X(n8059) );
  inv_x2_sg U7075 ( .A(\buff_mem[3][2] ), .X(n8061) );
  inv_x2_sg U7076 ( .A(\buff_mem[12][2] ), .X(n8063) );
  inv_x2_sg U7077 ( .A(\buff_mem[3][3] ), .X(n8065) );
  inv_x2_sg U7078 ( .A(\buff_mem[12][3] ), .X(n8067) );
  inv_x2_sg U7079 ( .A(\buff_mem[3][4] ), .X(n8069) );
  inv_x2_sg U7080 ( .A(\buff_mem[12][4] ), .X(n8071) );
  inv_x2_sg U7081 ( .A(\buff_mem[3][5] ), .X(n8073) );
  inv_x2_sg U7082 ( .A(\buff_mem[12][5] ), .X(n8075) );
  inv_x2_sg U7083 ( .A(\buff_mem[3][6] ), .X(n8077) );
  inv_x2_sg U7084 ( .A(\buff_mem[12][6] ), .X(n8079) );
  inv_x2_sg U7085 ( .A(\buff_mem[3][7] ), .X(n8081) );
  inv_x2_sg U7086 ( .A(\buff_mem[12][7] ), .X(n8083) );
  inv_x2_sg U7087 ( .A(\buff_mem[3][8] ), .X(n8085) );
  inv_x2_sg U7088 ( .A(\buff_mem[12][8] ), .X(n8087) );
  inv_x2_sg U7089 ( .A(\buff_mem[3][9] ), .X(n8089) );
  inv_x2_sg U7090 ( .A(\buff_mem[12][9] ), .X(n8091) );
  inv_x2_sg U7091 ( .A(\buff_mem[3][10] ), .X(n8093) );
  inv_x2_sg U7092 ( .A(\buff_mem[12][10] ), .X(n8095) );
  inv_x2_sg U7093 ( .A(\buff_mem[3][11] ), .X(n8097) );
  inv_x2_sg U7094 ( .A(\buff_mem[12][11] ), .X(n8099) );
  inv_x2_sg U7095 ( .A(n8263), .X(n8101) );
  inv_x4_sg U7096 ( .A(n5245), .X(n4880) );
  inv_x4_sg U7097 ( .A(n6014), .X(n4861) );
  inv_x4_sg U7098 ( .A(n5987), .X(n4870) );
  inv_x4_sg U7099 ( .A(n5972), .X(n4875) );
  nor_x8_sg U7100 ( .A(reset), .B(empty), .X(n6801) );
  inv_x4_sg U7101 ( .A(n7273), .X(n7337) );
  inv_x8_sg U7102 ( .A(n7337), .X(n7338) );
  inv_x8_sg U7103 ( .A(n7338), .X(n4909) );
  inv_x4_sg U7104 ( .A(n7265), .X(n7339) );
  inv_x8_sg U7105 ( .A(n7339), .X(n7340) );
  inv_x8_sg U7106 ( .A(n7340), .X(n5073) );
  nor_x8_sg U7107 ( .A(n5077), .B(n5078), .X(n6839) );
  nor_x8_sg U7108 ( .A(n5078), .B(n7334), .X(n6828) );
  inv_x8_sg U7109 ( .A(n7333), .X(n5078) );
  inv_x4_sg U7110 ( .A(n5999), .X(n4866) );
  inv_x4_sg U7111 ( .A(n6011), .X(n4862) );
  inv_x4_sg U7112 ( .A(n5969), .X(n4876) );
  inv_x4_sg U7113 ( .A(n5313), .X(n4879) );
  inv_x2_sg U7114 ( .A(n7341), .X(n7342) );
  inv_x2_sg U7115 ( .A(n7343), .X(n7344) );
  inv_x2_sg U7116 ( .A(n7345), .X(n7346) );
  inv_x2_sg U7117 ( .A(n7347), .X(n7348) );
  inv_x2_sg U7118 ( .A(n7349), .X(n7350) );
  inv_x2_sg U7119 ( .A(n7351), .X(n7352) );
  inv_x2_sg U7120 ( .A(n7353), .X(n7354) );
  inv_x2_sg U7121 ( .A(n7355), .X(n7356) );
  inv_x2_sg U7122 ( .A(n7357), .X(n7358) );
  inv_x2_sg U7123 ( .A(n7359), .X(n7360) );
  inv_x2_sg U7124 ( .A(n7361), .X(n7362) );
  inv_x2_sg U7125 ( .A(n7363), .X(n7364) );
  inv_x2_sg U7126 ( .A(n7365), .X(n7366) );
  inv_x2_sg U7127 ( .A(n7367), .X(n7368) );
  inv_x2_sg U7128 ( .A(n7369), .X(n7370) );
  inv_x2_sg U7129 ( .A(n7371), .X(n7372) );
  inv_x2_sg U7130 ( .A(n7373), .X(n7374) );
  inv_x2_sg U7131 ( .A(n7375), .X(n7376) );
  inv_x2_sg U7132 ( .A(n7377), .X(n7378) );
  inv_x2_sg U7133 ( .A(n7379), .X(n7380) );
  inv_x2_sg U7134 ( .A(n7381), .X(n7382) );
  inv_x2_sg U7135 ( .A(n7383), .X(n7384) );
  inv_x2_sg U7136 ( .A(n7385), .X(n7386) );
  inv_x2_sg U7137 ( .A(n7387), .X(n7388) );
  inv_x2_sg U7138 ( .A(n7389), .X(n7390) );
  inv_x2_sg U7139 ( .A(n7391), .X(n7392) );
  inv_x2_sg U7140 ( .A(n7393), .X(n7394) );
  inv_x2_sg U7141 ( .A(n7395), .X(n7396) );
  inv_x2_sg U7142 ( .A(n7397), .X(n7398) );
  inv_x2_sg U7143 ( .A(n7399), .X(n7400) );
  inv_x2_sg U7144 ( .A(n7401), .X(n7402) );
  inv_x2_sg U7145 ( .A(n7403), .X(n7404) );
  inv_x2_sg U7146 ( .A(n7405), .X(n7406) );
  inv_x2_sg U7147 ( .A(n7407), .X(n7408) );
  inv_x2_sg U7148 ( .A(n7409), .X(n7410) );
  inv_x2_sg U7149 ( .A(n7411), .X(n7412) );
  inv_x2_sg U7150 ( .A(n7413), .X(n7414) );
  inv_x2_sg U7151 ( .A(n7415), .X(n7416) );
  inv_x2_sg U7152 ( .A(n7417), .X(n7418) );
  inv_x2_sg U7153 ( .A(n7419), .X(n7420) );
  inv_x2_sg U7154 ( .A(n7421), .X(n7422) );
  inv_x2_sg U7155 ( .A(n7423), .X(n7424) );
  inv_x2_sg U7156 ( .A(n7425), .X(n7426) );
  inv_x2_sg U7157 ( .A(n7427), .X(n7428) );
  inv_x2_sg U7158 ( .A(n7429), .X(n7430) );
  inv_x2_sg U7159 ( .A(n7431), .X(n7432) );
  inv_x2_sg U7160 ( .A(n7433), .X(n7434) );
  inv_x2_sg U7161 ( .A(n7435), .X(n7436) );
  inv_x2_sg U7162 ( .A(n7437), .X(n7438) );
  inv_x2_sg U7163 ( .A(n7439), .X(n7440) );
  inv_x2_sg U7164 ( .A(n7441), .X(n7442) );
  inv_x2_sg U7165 ( .A(n7443), .X(n7444) );
  inv_x2_sg U7166 ( .A(n7445), .X(n7446) );
  inv_x2_sg U7167 ( .A(n7447), .X(n7448) );
  inv_x2_sg U7168 ( .A(n7449), .X(n7450) );
  inv_x2_sg U7169 ( .A(n7451), .X(n7452) );
  inv_x2_sg U7170 ( .A(n7453), .X(n7454) );
  inv_x2_sg U7171 ( .A(n7455), .X(n7456) );
  inv_x2_sg U7172 ( .A(n7457), .X(n7458) );
  inv_x2_sg U7173 ( .A(n7459), .X(n7460) );
  inv_x2_sg U7174 ( .A(n7461), .X(n7462) );
  inv_x2_sg U7175 ( .A(n7463), .X(n7464) );
  inv_x2_sg U7176 ( .A(n7465), .X(n7466) );
  inv_x2_sg U7177 ( .A(n7467), .X(n7468) );
  inv_x2_sg U7178 ( .A(n7469), .X(n7470) );
  inv_x2_sg U7179 ( .A(n7471), .X(n7472) );
  inv_x2_sg U7180 ( .A(n7473), .X(n7474) );
  inv_x2_sg U7181 ( .A(n7475), .X(n7476) );
  inv_x2_sg U7182 ( .A(n7477), .X(n7478) );
  inv_x2_sg U7183 ( .A(n7479), .X(n7480) );
  inv_x2_sg U7184 ( .A(n7481), .X(n7482) );
  inv_x2_sg U7185 ( .A(n7483), .X(n7484) );
  inv_x2_sg U7186 ( .A(n7485), .X(n7486) );
  inv_x2_sg U7187 ( .A(n7487), .X(n7488) );
  inv_x2_sg U7188 ( .A(n7489), .X(n7490) );
  inv_x2_sg U7189 ( .A(n7491), .X(n7492) );
  inv_x2_sg U7190 ( .A(n7493), .X(n7494) );
  inv_x2_sg U7191 ( .A(n7495), .X(n7496) );
  inv_x2_sg U7192 ( .A(n7497), .X(n7498) );
  inv_x2_sg U7193 ( .A(n7499), .X(n7500) );
  inv_x2_sg U7194 ( .A(n7501), .X(n7502) );
  inv_x2_sg U7195 ( .A(n7503), .X(n7504) );
  inv_x2_sg U7196 ( .A(n7505), .X(n7506) );
  inv_x2_sg U7197 ( .A(n7507), .X(n7508) );
  inv_x2_sg U7198 ( .A(n7509), .X(n7510) );
  inv_x2_sg U7199 ( .A(n7511), .X(n7512) );
  inv_x2_sg U7200 ( .A(n7513), .X(n7514) );
  inv_x2_sg U7201 ( .A(n7515), .X(n7516) );
  inv_x2_sg U7202 ( .A(n7517), .X(n7518) );
  inv_x2_sg U7203 ( .A(n7519), .X(n7520) );
  inv_x2_sg U7204 ( .A(n7521), .X(n7522) );
  inv_x2_sg U7205 ( .A(n7523), .X(n7524) );
  inv_x2_sg U7206 ( .A(n7525), .X(n7526) );
  inv_x2_sg U7207 ( .A(n7527), .X(n7528) );
  inv_x2_sg U7208 ( .A(n7529), .X(n7530) );
  inv_x2_sg U7209 ( .A(n7531), .X(n7532) );
  inv_x2_sg U7210 ( .A(n7533), .X(n7534) );
  inv_x2_sg U7211 ( .A(n7535), .X(n7536) );
  inv_x2_sg U7212 ( .A(n7537), .X(n7538) );
  inv_x2_sg U7213 ( .A(n7539), .X(n7540) );
  inv_x2_sg U7214 ( .A(n7541), .X(n7542) );
  inv_x2_sg U7215 ( .A(n7543), .X(n7544) );
  inv_x2_sg U7216 ( .A(n7545), .X(n7546) );
  inv_x2_sg U7217 ( .A(n7547), .X(n7548) );
  inv_x2_sg U7218 ( .A(n7549), .X(n7550) );
  inv_x2_sg U7219 ( .A(n7551), .X(n7552) );
  inv_x2_sg U7220 ( .A(n7553), .X(n7554) );
  inv_x2_sg U7221 ( .A(n7555), .X(n7556) );
  inv_x2_sg U7222 ( .A(n7557), .X(n7558) );
  inv_x2_sg U7223 ( .A(n7559), .X(n7560) );
  inv_x2_sg U7224 ( .A(n7561), .X(n7562) );
  inv_x2_sg U7225 ( .A(n7563), .X(n7564) );
  inv_x2_sg U7226 ( .A(n7565), .X(n7566) );
  inv_x2_sg U7227 ( .A(n7567), .X(n7568) );
  inv_x2_sg U7228 ( .A(n7569), .X(n7570) );
  inv_x2_sg U7229 ( .A(n7571), .X(n7572) );
  inv_x2_sg U7230 ( .A(n7573), .X(n7574) );
  inv_x2_sg U7231 ( .A(n7575), .X(n7576) );
  inv_x2_sg U7232 ( .A(n7577), .X(n7578) );
  inv_x2_sg U7233 ( .A(n7579), .X(n7580) );
  inv_x2_sg U7234 ( .A(n7581), .X(n7582) );
  inv_x2_sg U7235 ( .A(n7583), .X(n7584) );
  inv_x2_sg U7236 ( .A(n7585), .X(n7586) );
  inv_x2_sg U7237 ( .A(n7587), .X(n7588) );
  inv_x2_sg U7238 ( .A(n7589), .X(n7590) );
  inv_x2_sg U7239 ( .A(n7591), .X(n7592) );
  inv_x2_sg U7240 ( .A(n7593), .X(n7594) );
  inv_x2_sg U7241 ( .A(n7595), .X(n7596) );
  inv_x2_sg U7242 ( .A(n7597), .X(n7598) );
  inv_x2_sg U7243 ( .A(n7599), .X(n7600) );
  inv_x2_sg U7244 ( .A(n7601), .X(n7602) );
  inv_x2_sg U7245 ( .A(n7603), .X(n7604) );
  inv_x2_sg U7246 ( .A(n7605), .X(n7606) );
  inv_x2_sg U7247 ( .A(n7607), .X(n7608) );
  inv_x2_sg U7248 ( .A(n7609), .X(n7610) );
  inv_x2_sg U7249 ( .A(n7611), .X(n7612) );
  inv_x2_sg U7250 ( .A(n7613), .X(n7614) );
  inv_x2_sg U7251 ( .A(n7615), .X(n7616) );
  inv_x2_sg U7252 ( .A(n7617), .X(n7618) );
  inv_x2_sg U7253 ( .A(n7619), .X(n7620) );
  inv_x2_sg U7254 ( .A(n7621), .X(n7622) );
  inv_x2_sg U7255 ( .A(n7623), .X(n7624) );
  inv_x2_sg U7256 ( .A(n7625), .X(n7626) );
  inv_x2_sg U7257 ( .A(n7627), .X(n7628) );
  inv_x2_sg U7258 ( .A(n7629), .X(n7630) );
  inv_x2_sg U7259 ( .A(n7631), .X(n7632) );
  inv_x2_sg U7260 ( .A(n7633), .X(n7634) );
  inv_x2_sg U7261 ( .A(n7635), .X(n7636) );
  inv_x2_sg U7262 ( .A(n7637), .X(n7638) );
  inv_x2_sg U7263 ( .A(n7639), .X(n7640) );
  inv_x2_sg U7264 ( .A(n7641), .X(n7642) );
  inv_x2_sg U7265 ( .A(n7643), .X(n7644) );
  inv_x2_sg U7266 ( .A(n7645), .X(n7646) );
  inv_x2_sg U7267 ( .A(n7647), .X(n7648) );
  inv_x2_sg U7268 ( .A(n7649), .X(n7650) );
  inv_x2_sg U7269 ( .A(n7651), .X(n7652) );
  inv_x2_sg U7270 ( .A(n7653), .X(n7654) );
  inv_x2_sg U7271 ( .A(n7655), .X(n7656) );
  inv_x2_sg U7272 ( .A(n7657), .X(n7658) );
  inv_x2_sg U7273 ( .A(n7659), .X(n7660) );
  inv_x2_sg U7274 ( .A(n7661), .X(n7662) );
  inv_x2_sg U7275 ( .A(n7663), .X(n7664) );
  inv_x2_sg U7276 ( .A(n7665), .X(n7666) );
  inv_x2_sg U7277 ( .A(n7667), .X(n7668) );
  inv_x2_sg U7278 ( .A(n7669), .X(n7670) );
  inv_x2_sg U7279 ( .A(n7671), .X(n7672) );
  inv_x2_sg U7280 ( .A(n7673), .X(n7674) );
  inv_x2_sg U7281 ( .A(n7675), .X(n7676) );
  inv_x2_sg U7282 ( .A(n7677), .X(n7678) );
  inv_x2_sg U7283 ( .A(n7679), .X(n7680) );
  inv_x2_sg U7284 ( .A(n7681), .X(n7682) );
  inv_x2_sg U7285 ( .A(n7683), .X(n7684) );
  inv_x2_sg U7286 ( .A(n7685), .X(n7686) );
  inv_x2_sg U7287 ( .A(n7687), .X(n7688) );
  inv_x2_sg U7288 ( .A(n7689), .X(n7690) );
  inv_x2_sg U7289 ( .A(n7691), .X(n7692) );
  inv_x2_sg U7290 ( .A(n7693), .X(n7694) );
  inv_x2_sg U7291 ( .A(n7695), .X(n7696) );
  inv_x2_sg U7292 ( .A(n7697), .X(n7698) );
  inv_x2_sg U7293 ( .A(n7699), .X(n7700) );
  inv_x2_sg U7294 ( .A(n7701), .X(n7702) );
  inv_x2_sg U7295 ( .A(n7703), .X(n7704) );
  inv_x2_sg U7296 ( .A(n7705), .X(n7706) );
  inv_x2_sg U7297 ( .A(n7707), .X(n7708) );
  inv_x2_sg U7298 ( .A(n7709), .X(n7710) );
  inv_x2_sg U7299 ( .A(n7711), .X(n7712) );
  inv_x2_sg U7300 ( .A(n7713), .X(n7714) );
  inv_x2_sg U7301 ( .A(n7715), .X(n7716) );
  inv_x2_sg U7302 ( .A(n7717), .X(n7718) );
  inv_x2_sg U7303 ( .A(n7719), .X(n7720) );
  inv_x2_sg U7304 ( .A(n7721), .X(n7722) );
  inv_x2_sg U7305 ( .A(n7723), .X(n7724) );
  inv_x2_sg U7306 ( .A(n7725), .X(n7726) );
  inv_x2_sg U7307 ( .A(n7727), .X(n7728) );
  inv_x2_sg U7308 ( .A(n7729), .X(n7730) );
  inv_x2_sg U7309 ( .A(n7731), .X(n7732) );
  inv_x2_sg U7310 ( .A(n7733), .X(n7734) );
  inv_x2_sg U7311 ( .A(n7735), .X(n7736) );
  inv_x2_sg U7312 ( .A(n7737), .X(n7738) );
  inv_x2_sg U7313 ( .A(n7739), .X(n7740) );
  inv_x2_sg U7314 ( .A(n7741), .X(n7742) );
  inv_x2_sg U7315 ( .A(n7743), .X(n7744) );
  inv_x2_sg U7316 ( .A(n7745), .X(n7746) );
  inv_x2_sg U7317 ( .A(n7747), .X(n7748) );
  inv_x2_sg U7318 ( .A(n7749), .X(n7750) );
  inv_x2_sg U7319 ( .A(n7751), .X(n7752) );
  inv_x2_sg U7320 ( .A(n7753), .X(n7754) );
  inv_x2_sg U7321 ( .A(n7755), .X(n7756) );
  inv_x2_sg U7322 ( .A(n7757), .X(n7758) );
  inv_x2_sg U7323 ( .A(n7759), .X(n7760) );
  inv_x2_sg U7324 ( .A(n7761), .X(n7762) );
  inv_x2_sg U7325 ( .A(n7763), .X(n7764) );
  inv_x2_sg U7326 ( .A(n7765), .X(n7766) );
  inv_x2_sg U7327 ( .A(n7767), .X(n7768) );
  inv_x2_sg U7328 ( .A(n7769), .X(n7770) );
  inv_x2_sg U7329 ( .A(n7771), .X(n7772) );
  inv_x2_sg U7330 ( .A(n7773), .X(n7774) );
  inv_x2_sg U7331 ( .A(n7775), .X(n7776) );
  inv_x2_sg U7332 ( .A(n7777), .X(n7778) );
  inv_x2_sg U7333 ( .A(n7779), .X(n7780) );
  inv_x4_sg U7334 ( .A(n7781), .X(n7782) );
  inv_x4_sg U7335 ( .A(n7783), .X(n7784) );
  inv_x4_sg U7336 ( .A(n7785), .X(n7786) );
  inv_x4_sg U7337 ( .A(n7787), .X(n7788) );
  inv_x4_sg U7338 ( .A(n7789), .X(n7790) );
  inv_x4_sg U7339 ( .A(n7791), .X(n7792) );
  inv_x4_sg U7340 ( .A(n7793), .X(n7794) );
  inv_x4_sg U7341 ( .A(n7795), .X(n7796) );
  inv_x4_sg U7342 ( .A(n7797), .X(n7798) );
  inv_x4_sg U7343 ( .A(n7799), .X(n7800) );
  inv_x4_sg U7344 ( .A(n7801), .X(n7802) );
  inv_x4_sg U7345 ( .A(n7803), .X(n7804) );
  inv_x4_sg U7346 ( .A(n7805), .X(n7806) );
  inv_x4_sg U7347 ( .A(n7807), .X(n7808) );
  inv_x4_sg U7348 ( .A(n7809), .X(n7810) );
  inv_x4_sg U7349 ( .A(n7811), .X(n7812) );
  inv_x4_sg U7350 ( .A(n7813), .X(n7814) );
  inv_x4_sg U7351 ( .A(n7815), .X(n7816) );
  inv_x4_sg U7352 ( .A(n7817), .X(n7818) );
  inv_x4_sg U7353 ( .A(n7819), .X(n7820) );
  inv_x4_sg U7354 ( .A(n7821), .X(n7822) );
  inv_x4_sg U7355 ( .A(n7823), .X(n7824) );
  inv_x4_sg U7356 ( .A(n7825), .X(n7826) );
  inv_x4_sg U7357 ( .A(n7827), .X(n7828) );
  inv_x4_sg U7358 ( .A(n7829), .X(n7830) );
  inv_x4_sg U7359 ( .A(n7831), .X(n7832) );
  inv_x4_sg U7360 ( .A(n7833), .X(n7834) );
  inv_x4_sg U7361 ( .A(n7835), .X(n7836) );
  inv_x4_sg U7362 ( .A(n7837), .X(n7838) );
  inv_x4_sg U7363 ( .A(n7839), .X(n7840) );
  inv_x4_sg U7364 ( .A(n7841), .X(n7842) );
  inv_x4_sg U7365 ( .A(n7843), .X(n7844) );
  inv_x4_sg U7366 ( .A(n7845), .X(n7846) );
  inv_x4_sg U7367 ( .A(n7847), .X(n7848) );
  inv_x4_sg U7368 ( .A(n7849), .X(n7850) );
  inv_x4_sg U7369 ( .A(n7851), .X(n7852) );
  inv_x4_sg U7370 ( .A(n7853), .X(n7854) );
  inv_x4_sg U7371 ( .A(n7855), .X(n7856) );
  inv_x4_sg U7372 ( .A(n7857), .X(n7858) );
  inv_x4_sg U7373 ( .A(n7859), .X(n7860) );
  inv_x4_sg U7374 ( .A(n7861), .X(n7862) );
  inv_x4_sg U7375 ( .A(n7863), .X(n7864) );
  inv_x4_sg U7376 ( .A(n7865), .X(n7866) );
  inv_x4_sg U7377 ( .A(n7867), .X(n7868) );
  inv_x4_sg U7378 ( .A(n7869), .X(n7870) );
  inv_x4_sg U7379 ( .A(n7871), .X(n7872) );
  inv_x4_sg U7380 ( .A(n7873), .X(n7874) );
  inv_x4_sg U7381 ( .A(n7875), .X(n7876) );
  inv_x4_sg U7382 ( .A(n7877), .X(n7878) );
  inv_x4_sg U7383 ( .A(n7879), .X(n7880) );
  inv_x4_sg U7384 ( .A(n7881), .X(n7882) );
  inv_x4_sg U7385 ( .A(n7883), .X(n7884) );
  inv_x4_sg U7386 ( .A(n7885), .X(n7886) );
  inv_x4_sg U7387 ( .A(n7887), .X(n7888) );
  inv_x4_sg U7388 ( .A(n7889), .X(n7890) );
  inv_x4_sg U7389 ( .A(n7891), .X(n7892) );
  inv_x4_sg U7390 ( .A(n7893), .X(n7894) );
  inv_x4_sg U7391 ( .A(n7895), .X(n7896) );
  inv_x4_sg U7392 ( .A(n7897), .X(n7898) );
  inv_x4_sg U7393 ( .A(n7899), .X(n7900) );
  inv_x4_sg U7394 ( .A(n7901), .X(n7902) );
  inv_x4_sg U7395 ( .A(n7903), .X(n7904) );
  inv_x4_sg U7396 ( .A(n7905), .X(n7906) );
  inv_x4_sg U7397 ( .A(n7907), .X(n7908) );
  inv_x4_sg U7398 ( .A(n7909), .X(n7910) );
  inv_x4_sg U7399 ( .A(n7911), .X(n7912) );
  inv_x4_sg U7400 ( .A(n7913), .X(n7914) );
  inv_x4_sg U7401 ( .A(n7915), .X(n7916) );
  inv_x4_sg U7402 ( .A(n7917), .X(n7918) );
  inv_x4_sg U7403 ( .A(n7919), .X(n7920) );
  inv_x4_sg U7404 ( .A(n7921), .X(n7922) );
  inv_x4_sg U7405 ( .A(n7923), .X(n7924) );
  inv_x4_sg U7406 ( .A(n7925), .X(n7926) );
  inv_x4_sg U7407 ( .A(n7927), .X(n7928) );
  inv_x4_sg U7408 ( .A(n7929), .X(n7930) );
  inv_x4_sg U7409 ( .A(n7931), .X(n7932) );
  inv_x4_sg U7410 ( .A(n7933), .X(n7934) );
  inv_x4_sg U7411 ( .A(n7935), .X(n7936) );
  inv_x4_sg U7412 ( .A(n7937), .X(n7938) );
  inv_x4_sg U7413 ( .A(n7939), .X(n7940) );
  inv_x4_sg U7414 ( .A(n7941), .X(n7942) );
  inv_x4_sg U7415 ( .A(n7943), .X(n7944) );
  inv_x4_sg U7416 ( .A(n7945), .X(n7946) );
  inv_x4_sg U7417 ( .A(n7947), .X(n7948) );
  inv_x4_sg U7418 ( .A(n7949), .X(n7950) );
  inv_x4_sg U7419 ( .A(n7951), .X(n7952) );
  inv_x4_sg U7420 ( .A(n7953), .X(n7954) );
  inv_x4_sg U7421 ( .A(n7955), .X(n7956) );
  inv_x4_sg U7422 ( .A(n7957), .X(n7958) );
  inv_x4_sg U7423 ( .A(n7959), .X(n7960) );
  inv_x4_sg U7424 ( .A(n7961), .X(n7962) );
  inv_x4_sg U7425 ( .A(n7963), .X(n7964) );
  inv_x4_sg U7426 ( .A(n7965), .X(n7966) );
  inv_x4_sg U7427 ( .A(n7967), .X(n7968) );
  inv_x4_sg U7428 ( .A(n7969), .X(n7970) );
  inv_x4_sg U7429 ( .A(n7971), .X(n7972) );
  inv_x4_sg U7430 ( .A(n7973), .X(n7974) );
  inv_x4_sg U7431 ( .A(n7975), .X(n7976) );
  inv_x4_sg U7432 ( .A(n7977), .X(n7978) );
  inv_x4_sg U7433 ( .A(n7979), .X(n7980) );
  inv_x4_sg U7434 ( .A(n7981), .X(n7982) );
  inv_x4_sg U7435 ( .A(n7983), .X(n7984) );
  inv_x4_sg U7436 ( .A(n7985), .X(n7986) );
  inv_x4_sg U7437 ( .A(n7987), .X(n7988) );
  inv_x4_sg U7438 ( .A(n7989), .X(n7990) );
  inv_x4_sg U7439 ( .A(n7991), .X(n7992) );
  inv_x4_sg U7440 ( .A(n7993), .X(n7994) );
  inv_x4_sg U7441 ( .A(n7995), .X(n7996) );
  inv_x4_sg U7442 ( .A(n7997), .X(n7998) );
  inv_x4_sg U7443 ( .A(n7999), .X(n8000) );
  inv_x4_sg U7444 ( .A(n8001), .X(n8002) );
  inv_x4_sg U7445 ( .A(n8003), .X(n8004) );
  inv_x4_sg U7446 ( .A(n8005), .X(n8006) );
  inv_x4_sg U7447 ( .A(n8007), .X(n8008) );
  inv_x4_sg U7448 ( .A(n8009), .X(n8010) );
  inv_x4_sg U7449 ( .A(n8011), .X(n8012) );
  inv_x4_sg U7450 ( .A(n8013), .X(n8014) );
  inv_x4_sg U7451 ( .A(n8015), .X(n8016) );
  inv_x4_sg U7452 ( .A(n8017), .X(n8018) );
  inv_x4_sg U7453 ( .A(n8019), .X(n8020) );
  inv_x4_sg U7454 ( .A(n8021), .X(n8022) );
  inv_x4_sg U7455 ( .A(n8023), .X(n8024) );
  inv_x4_sg U7456 ( .A(n8025), .X(n8026) );
  inv_x4_sg U7457 ( .A(n8027), .X(n8028) );
  inv_x4_sg U7458 ( .A(n8029), .X(n8030) );
  inv_x4_sg U7459 ( .A(n8031), .X(n8032) );
  inv_x4_sg U7460 ( .A(n8033), .X(n8034) );
  inv_x4_sg U7461 ( .A(n8035), .X(n8036) );
  inv_x4_sg U7462 ( .A(n8037), .X(n8038) );
  inv_x4_sg U7463 ( .A(n8039), .X(n8040) );
  inv_x4_sg U7464 ( .A(n8041), .X(n8042) );
  inv_x4_sg U7465 ( .A(n8043), .X(n8044) );
  inv_x4_sg U7466 ( .A(n8045), .X(n8046) );
  inv_x4_sg U7467 ( .A(n8047), .X(n8048) );
  inv_x4_sg U7468 ( .A(n8049), .X(n8050) );
  inv_x4_sg U7469 ( .A(n8051), .X(n8052) );
  inv_x4_sg U7470 ( .A(n8053), .X(n8054) );
  inv_x4_sg U7471 ( .A(n8055), .X(n8056) );
  inv_x4_sg U7472 ( .A(n8057), .X(n8058) );
  inv_x4_sg U7473 ( .A(n8059), .X(n8060) );
  inv_x4_sg U7474 ( .A(n8061), .X(n8062) );
  inv_x4_sg U7475 ( .A(n8063), .X(n8064) );
  inv_x4_sg U7476 ( .A(n8065), .X(n8066) );
  inv_x4_sg U7477 ( .A(n8067), .X(n8068) );
  inv_x4_sg U7478 ( .A(n8069), .X(n8070) );
  inv_x4_sg U7479 ( .A(n8071), .X(n8072) );
  inv_x4_sg U7480 ( .A(n8073), .X(n8074) );
  inv_x4_sg U7481 ( .A(n8075), .X(n8076) );
  inv_x4_sg U7482 ( .A(n8077), .X(n8078) );
  inv_x4_sg U7483 ( .A(n8079), .X(n8080) );
  inv_x4_sg U7484 ( .A(n8081), .X(n8082) );
  inv_x4_sg U7485 ( .A(n8083), .X(n8084) );
  inv_x4_sg U7486 ( .A(n8085), .X(n8086) );
  inv_x4_sg U7487 ( .A(n8087), .X(n8088) );
  inv_x4_sg U7488 ( .A(n8089), .X(n8090) );
  inv_x4_sg U7489 ( .A(n8091), .X(n8092) );
  inv_x4_sg U7490 ( .A(n8093), .X(n8094) );
  inv_x4_sg U7491 ( .A(n8095), .X(n8096) );
  inv_x4_sg U7492 ( .A(n8097), .X(n8098) );
  inv_x4_sg U7493 ( .A(n8099), .X(n8100) );
  inv_x4_sg U7494 ( .A(n8101), .X(full) );
  inv_x4_sg U7495 ( .A(n7267), .X(n8103) );
  inv_x8_sg U7496 ( .A(n8103), .X(empty) );
  nand_x2_sg U7497 ( .A(n5256), .B(n4888), .X(n5255) );
  nor_x8_sg U7498 ( .A(n4888), .B(reset), .X(n5167) );
  inv_x8_sg U7499 ( .A(n6038), .X(n4888) );
  inv_x4_sg U7500 ( .A(n7271), .X(n8105) );
  inv_x8_sg U7501 ( .A(n8105), .X(n8106) );
  nand_x4_sg U7502 ( .A(n5588), .B(n8106), .X(n5586) );
  inv_x8_sg U7503 ( .A(n6810), .X(n4899) );
  nand_x1_sg U7504 ( .A(n8216), .B(n7456), .X(n6809) );
  nand_x1_sg U7505 ( .A(n8216), .B(n7470), .X(n6769) );
  nand_x1_sg U7506 ( .A(n8216), .B(n7498), .X(n6691) );
  nand_x1_sg U7507 ( .A(n8216), .B(n7512), .X(n6652) );
  nand_x1_sg U7508 ( .A(n8216), .B(n7540), .X(n6574) );
  nand_x1_sg U7509 ( .A(n8216), .B(n7554), .X(n6535) );
  nand_x1_sg U7510 ( .A(n8216), .B(n7582), .X(n6457) );
  nand_x1_sg U7511 ( .A(n8216), .B(n7596), .X(n6418) );
  nand_x1_sg U7512 ( .A(n8216), .B(n7344), .X(n6340) );
  nand_x1_sg U7513 ( .A(n8216), .B(n7358), .X(n6301) );
  nand_x1_sg U7514 ( .A(n8216), .B(n7386), .X(n6223) );
  nand_x1_sg U7515 ( .A(n8216), .B(n7400), .X(n6184) );
  nand_x1_sg U7516 ( .A(n8216), .B(n7428), .X(n6106) );
  nand_x1_sg U7517 ( .A(n8216), .B(n7442), .X(n6047) );
  nand_x1_sg U7518 ( .A(n8216), .B(n7484), .X(n6730) );
  nand_x1_sg U7519 ( .A(n8216), .B(n7526), .X(n6613) );
  nand_x1_sg U7520 ( .A(n8216), .B(n7568), .X(n6496) );
  nand_x1_sg U7521 ( .A(n8216), .B(n7610), .X(n6379) );
  nand_x1_sg U7522 ( .A(n6048), .B(n7372), .X(n6262) );
  nand_x1_sg U7523 ( .A(n8216), .B(n7414), .X(n6145) );
  nand_x1_sg U7524 ( .A(n8188), .B(n7462), .X(n6843) );
  nand_x1_sg U7525 ( .A(n8197), .B(n7458), .X(n6834) );
  nand_x1_sg U7526 ( .A(n8188), .B(n7476), .X(n6795) );
  nand_x1_sg U7527 ( .A(n8197), .B(n7472), .X(n6787) );
  nand_x1_sg U7528 ( .A(n8188), .B(n7518), .X(n6678) );
  nand_x1_sg U7529 ( .A(n8197), .B(n7514), .X(n6670) );
  nand_x1_sg U7530 ( .A(n8188), .B(n7532), .X(n6639) );
  nand_x1_sg U7531 ( .A(n8197), .B(n7528), .X(n6631) );
  nand_x1_sg U7532 ( .A(n8188), .B(n7546), .X(n6600) );
  nand_x1_sg U7533 ( .A(n8197), .B(n7542), .X(n6592) );
  nand_x1_sg U7534 ( .A(n8188), .B(n7574), .X(n6522) );
  nand_x1_sg U7535 ( .A(n8197), .B(n7570), .X(n6514) );
  nand_x1_sg U7536 ( .A(n8188), .B(n7588), .X(n6483) );
  nand_x1_sg U7537 ( .A(n8197), .B(n7584), .X(n6475) );
  nand_x1_sg U7538 ( .A(n8188), .B(n7602), .X(n6444) );
  nand_x1_sg U7539 ( .A(n8197), .B(n7598), .X(n6436) );
  nand_x1_sg U7540 ( .A(n8188), .B(n7364), .X(n6327) );
  nand_x1_sg U7541 ( .A(n8197), .B(n7360), .X(n6319) );
  nand_x1_sg U7542 ( .A(n8188), .B(n7378), .X(n6288) );
  nand_x1_sg U7543 ( .A(n8197), .B(n7374), .X(n6280) );
  nand_x1_sg U7544 ( .A(n8188), .B(n7392), .X(n6249) );
  nand_x1_sg U7545 ( .A(n8197), .B(n7388), .X(n6241) );
  nand_x1_sg U7546 ( .A(n8188), .B(n7420), .X(n6171) );
  nand_x1_sg U7547 ( .A(n8197), .B(n7416), .X(n6163) );
  nand_x1_sg U7548 ( .A(n8188), .B(n7434), .X(n6132) );
  nand_x1_sg U7549 ( .A(n8197), .B(n7430), .X(n6124) );
  nand_x1_sg U7550 ( .A(n8188), .B(n7448), .X(n6088) );
  nand_x1_sg U7551 ( .A(n8197), .B(n7444), .X(n6075) );
  nand_x1_sg U7552 ( .A(n8193), .B(n7460), .X(n6836) );
  nand_x1_sg U7553 ( .A(n8193), .B(n7474), .X(n6789) );
  nand_x1_sg U7554 ( .A(n8193), .B(n7516), .X(n6672) );
  nand_x1_sg U7555 ( .A(n8193), .B(n7530), .X(n6633) );
  nand_x1_sg U7556 ( .A(n8193), .B(n7544), .X(n6594) );
  nand_x1_sg U7557 ( .A(n8193), .B(n7572), .X(n6516) );
  nand_x1_sg U7558 ( .A(n8193), .B(n7586), .X(n6477) );
  nand_x1_sg U7559 ( .A(n8193), .B(n7600), .X(n6438) );
  nand_x1_sg U7560 ( .A(n8193), .B(n7362), .X(n6321) );
  nand_x1_sg U7561 ( .A(n8193), .B(n7376), .X(n6282) );
  nand_x1_sg U7562 ( .A(n8193), .B(n7390), .X(n6243) );
  nand_x1_sg U7563 ( .A(n8193), .B(n7418), .X(n6165) );
  nand_x1_sg U7564 ( .A(n8193), .B(n7432), .X(n6126) );
  nand_x1_sg U7565 ( .A(n8193), .B(n7446), .X(n6079) );
  nand_x1_sg U7566 ( .A(n8188), .B(n7490), .X(n6756) );
  nand_x1_sg U7567 ( .A(n8193), .B(n7488), .X(n6750) );
  nand_x1_sg U7568 ( .A(n8197), .B(n7486), .X(n6748) );
  nand_x1_sg U7569 ( .A(n8188), .B(n7504), .X(n6717) );
  nand_x1_sg U7570 ( .A(n8193), .B(n7502), .X(n6711) );
  nand_x1_sg U7571 ( .A(n8197), .B(n7500), .X(n6709) );
  nand_x1_sg U7572 ( .A(n8188), .B(n7560), .X(n6561) );
  nand_x1_sg U7573 ( .A(n8193), .B(n7558), .X(n6555) );
  nand_x1_sg U7574 ( .A(n8197), .B(n7556), .X(n6553) );
  nand_x1_sg U7575 ( .A(n6089), .B(n7616), .X(n6405) );
  nand_x1_sg U7576 ( .A(n6080), .B(n7614), .X(n6399) );
  nand_x1_sg U7577 ( .A(n6076), .B(n7612), .X(n6397) );
  nand_x1_sg U7578 ( .A(n8188), .B(n7350), .X(n6366) );
  nand_x1_sg U7579 ( .A(n8193), .B(n7348), .X(n6360) );
  nand_x1_sg U7580 ( .A(n8197), .B(n7346), .X(n6358) );
  nand_x1_sg U7581 ( .A(n8188), .B(n7406), .X(n6210) );
  nand_x1_sg U7582 ( .A(n8193), .B(n7404), .X(n6204) );
  nand_x1_sg U7583 ( .A(n8197), .B(n7402), .X(n6202) );
  nand_x1_sg U7584 ( .A(n8202), .B(n7466), .X(n6825) );
  nand_x1_sg U7585 ( .A(n6065), .B(n7480), .X(n6779) );
  nand_x1_sg U7586 ( .A(n8202), .B(n7494), .X(n6740) );
  nand_x1_sg U7587 ( .A(n6065), .B(n7508), .X(n6701) );
  nand_x1_sg U7588 ( .A(n8202), .B(n7522), .X(n6662) );
  nand_x1_sg U7589 ( .A(n6065), .B(n7536), .X(n6623) );
  nand_x1_sg U7590 ( .A(n8202), .B(n7550), .X(n6584) );
  nand_x1_sg U7591 ( .A(n6065), .B(n7564), .X(n6545) );
  nand_x1_sg U7592 ( .A(n8202), .B(n7578), .X(n6506) );
  nand_x1_sg U7593 ( .A(n6065), .B(n7592), .X(n6467) );
  nand_x1_sg U7594 ( .A(n8202), .B(n7606), .X(n6428) );
  nand_x1_sg U7595 ( .A(n6065), .B(n7620), .X(n6389) );
  nand_x1_sg U7596 ( .A(n8202), .B(n7354), .X(n6350) );
  nand_x1_sg U7597 ( .A(n6065), .B(n7368), .X(n6311) );
  nand_x1_sg U7598 ( .A(n8202), .B(n7382), .X(n6272) );
  nand_x1_sg U7599 ( .A(n6065), .B(n7396), .X(n6233) );
  nand_x1_sg U7600 ( .A(n8202), .B(n7410), .X(n6194) );
  nand_x1_sg U7601 ( .A(n6065), .B(n7424), .X(n6155) );
  nand_x1_sg U7602 ( .A(n8202), .B(n7438), .X(n6116) );
  nand_x1_sg U7603 ( .A(n6065), .B(n7452), .X(n6064) );
  nand_x2_sg U7604 ( .A(n5262), .B(n5263), .X(n5177) );
  inv_x2_sg U7605 ( .A(n8179), .X(n8183) );
  inv_x2_sg U7606 ( .A(n8179), .X(n8184) );
  inv_x2_sg U7607 ( .A(n8179), .X(n8185) );
  inv_x2_sg U7608 ( .A(n8179), .X(n8186) );
  inv_x2_sg U7609 ( .A(n8173), .X(n8174) );
  inv_x2_sg U7610 ( .A(n8173), .X(n8175) );
  inv_x2_sg U7611 ( .A(n8173), .X(n8177) );
  inv_x2_sg U7612 ( .A(n8173), .X(n8176) );
  nor_x1_sg U7613 ( .A(n5254), .B(n5255), .X(n5253) );
  nor_x1_sg U7614 ( .A(n6800), .B(n8217), .X(N142) );
  nand_x2_sg U7615 ( .A(n6829), .B(n6830), .X(n6802) );
  nand_x2_sg U7616 ( .A(n6804), .B(n6805), .X(n6803) );
  nor_x1_sg U7617 ( .A(n6761), .B(n8218), .X(N143) );
  nand_x2_sg U7618 ( .A(n6782), .B(n6783), .X(n6762) );
  nand_x2_sg U7619 ( .A(n6764), .B(n6765), .X(n6763) );
  nor_x1_sg U7620 ( .A(n6683), .B(n8217), .X(N145) );
  nand_x2_sg U7621 ( .A(n6704), .B(n6705), .X(n6684) );
  nand_x2_sg U7622 ( .A(n6686), .B(n6687), .X(n6685) );
  nor_x1_sg U7623 ( .A(n6644), .B(n8218), .X(N146) );
  nand_x2_sg U7624 ( .A(n6665), .B(n6666), .X(n6645) );
  nand_x2_sg U7625 ( .A(n6647), .B(n6648), .X(n6646) );
  nor_x1_sg U7626 ( .A(n6566), .B(n8217), .X(N148) );
  nand_x2_sg U7627 ( .A(n6587), .B(n6588), .X(n6567) );
  nand_x2_sg U7628 ( .A(n6569), .B(n6570), .X(n6568) );
  nor_x1_sg U7629 ( .A(n6527), .B(n8218), .X(N149) );
  nand_x2_sg U7630 ( .A(n6548), .B(n6549), .X(n6528) );
  nand_x2_sg U7631 ( .A(n6530), .B(n6531), .X(n6529) );
  nor_x1_sg U7632 ( .A(n6449), .B(n8217), .X(N151) );
  nand_x2_sg U7633 ( .A(n6470), .B(n6471), .X(n6450) );
  nand_x2_sg U7634 ( .A(n6452), .B(n6453), .X(n6451) );
  nor_x1_sg U7635 ( .A(n6410), .B(n8218), .X(N152) );
  nand_x2_sg U7636 ( .A(n6431), .B(n6432), .X(n6411) );
  nand_x2_sg U7637 ( .A(n6413), .B(n6414), .X(n6412) );
  nor_x1_sg U7638 ( .A(n6332), .B(n8217), .X(N154) );
  nand_x2_sg U7639 ( .A(n6353), .B(n6354), .X(n6333) );
  nand_x2_sg U7640 ( .A(n6335), .B(n6336), .X(n6334) );
  nor_x1_sg U7641 ( .A(n6293), .B(n8218), .X(N155) );
  nand_x2_sg U7642 ( .A(n6314), .B(n6315), .X(n6294) );
  nand_x2_sg U7643 ( .A(n6296), .B(n6297), .X(n6295) );
  nor_x1_sg U7644 ( .A(n6215), .B(n8217), .X(N157) );
  nand_x2_sg U7645 ( .A(n6236), .B(n6237), .X(n6216) );
  nand_x2_sg U7646 ( .A(n6218), .B(n6219), .X(n6217) );
  nor_x1_sg U7647 ( .A(n6176), .B(n8218), .X(N158) );
  nand_x2_sg U7648 ( .A(n6197), .B(n6198), .X(n6177) );
  nand_x2_sg U7649 ( .A(n6179), .B(n6180), .X(n6178) );
  nor_x1_sg U7650 ( .A(n6098), .B(n8217), .X(N160) );
  nand_x2_sg U7651 ( .A(n6119), .B(n6120), .X(n6099) );
  nand_x2_sg U7652 ( .A(n6101), .B(n6102), .X(n6100) );
  nor_x1_sg U7653 ( .A(n6039), .B(n8218), .X(N161) );
  nand_x2_sg U7654 ( .A(n6070), .B(n6071), .X(n6040) );
  nand_x2_sg U7655 ( .A(n6042), .B(n6043), .X(n6041) );
  nor_x1_sg U7656 ( .A(n6722), .B(n6038), .X(N144) );
  nand_x2_sg U7657 ( .A(n6743), .B(n6744), .X(n6723) );
  nand_x2_sg U7658 ( .A(n6725), .B(n6726), .X(n6724) );
  nor_x1_sg U7659 ( .A(n6605), .B(n6038), .X(N147) );
  nand_x2_sg U7660 ( .A(n6626), .B(n6627), .X(n6606) );
  nand_x2_sg U7661 ( .A(n6608), .B(n6609), .X(n6607) );
  nor_x1_sg U7662 ( .A(n6488), .B(n6038), .X(N150) );
  nand_x2_sg U7663 ( .A(n6509), .B(n6510), .X(n6489) );
  nand_x2_sg U7664 ( .A(n6491), .B(n6492), .X(n6490) );
  nor_x1_sg U7665 ( .A(n6371), .B(n6038), .X(N153) );
  nand_x2_sg U7666 ( .A(n6392), .B(n6393), .X(n6372) );
  nand_x2_sg U7667 ( .A(n6374), .B(n6375), .X(n6373) );
  nor_x1_sg U7668 ( .A(n6254), .B(n6038), .X(N156) );
  nand_x2_sg U7669 ( .A(n6275), .B(n6276), .X(n6255) );
  nand_x2_sg U7670 ( .A(n6257), .B(n6258), .X(n6256) );
  nor_x1_sg U7671 ( .A(n6137), .B(n6038), .X(N159) );
  nand_x2_sg U7672 ( .A(n6158), .B(n6159), .X(n6138) );
  nand_x2_sg U7673 ( .A(n6140), .B(n6141), .X(n6139) );
  nand_x1_sg U7674 ( .A(n6032), .B(n5078), .X(n6031) );
  nand_x1_sg U7675 ( .A(n4908), .B(n5259), .X(n5258) );
  nor_x1_sg U7676 ( .A(n5257), .B(n4896), .X(n5256) );
  nand_x2_sg U7677 ( .A(n5739), .B(n4852), .X(n5738) );
  nand_x2_sg U7678 ( .A(n5167), .B(n5168), .X(n5166) );
  nor_x1_sg U7679 ( .A(n5171), .B(n5172), .X(n5170) );
  nor_x1_sg U7680 ( .A(n5179), .B(n5180), .X(n5169) );
  nand_x1_sg U7681 ( .A(n4907), .B(n4910), .X(n5587) );
  nand_x2_sg U7682 ( .A(n5849), .B(n5739), .X(n5848) );
  nor_x1_sg U7683 ( .A(n5850), .B(n4911), .X(n5849) );
  nand_x1_sg U7684 ( .A(n5579), .B(n4909), .X(n5583) );
  nand_x4_sg U7685 ( .A(n5579), .B(n5580), .X(n5176) );
  nand_x4_sg U7686 ( .A(n6023), .B(n6024), .X(n5270) );
  nand_x1_sg U7687 ( .A(n5261), .B(n5073), .X(n6023) );
  nand_x1_sg U7688 ( .A(n7340), .B(n4895), .X(n6024) );
  nor_x1_sg U7689 ( .A(n5268), .B(n5269), .X(n5267) );
  nand_x2_sg U7690 ( .A(n5274), .B(n5275), .X(n5264) );
  nand_x2_sg U7691 ( .A(n5266), .B(n5267), .X(n5265) );
  nand_x1_sg U7692 ( .A(n8106), .B(n5276), .X(n5275) );
  nand_x1_sg U7693 ( .A(empty), .B(n7280), .X(n5247) );
  nor_x1_sg U7694 ( .A(n4843), .B(n5167), .X(n5248) );
  nand_x1_sg U7695 ( .A(n8212), .B(n7454), .X(n6813) );
  nand_x1_sg U7696 ( .A(n8212), .B(n7468), .X(n6771) );
  nand_x1_sg U7697 ( .A(n8212), .B(n7496), .X(n6693) );
  nand_x1_sg U7698 ( .A(n8212), .B(n7510), .X(n6654) );
  nand_x1_sg U7699 ( .A(n8212), .B(n7538), .X(n6576) );
  nand_x1_sg U7700 ( .A(n8212), .B(n7552), .X(n6537) );
  nand_x1_sg U7701 ( .A(n8212), .B(n7580), .X(n6459) );
  nand_x1_sg U7702 ( .A(n8212), .B(n7594), .X(n6420) );
  nand_x1_sg U7703 ( .A(n8212), .B(n7342), .X(n6342) );
  nand_x1_sg U7704 ( .A(n8212), .B(n7356), .X(n6303) );
  nand_x1_sg U7705 ( .A(n8212), .B(n7384), .X(n6225) );
  nand_x1_sg U7706 ( .A(n8212), .B(n7398), .X(n6186) );
  nand_x1_sg U7707 ( .A(n8212), .B(n7426), .X(n6108) );
  nand_x1_sg U7708 ( .A(n8212), .B(n7440), .X(n6051) );
  nand_x2_sg U7709 ( .A(n6808), .B(n6809), .X(n6807) );
  nand_x2_sg U7710 ( .A(n6812), .B(n6813), .X(n6806) );
  nand_x1_sg U7711 ( .A(n8214), .B(n7688), .X(n6808) );
  nand_x2_sg U7712 ( .A(n6768), .B(n6769), .X(n6767) );
  nand_x2_sg U7713 ( .A(n6770), .B(n6771), .X(n6766) );
  nand_x1_sg U7714 ( .A(n8214), .B(n7696), .X(n6768) );
  nand_x2_sg U7715 ( .A(n6690), .B(n6691), .X(n6689) );
  nand_x2_sg U7716 ( .A(n6692), .B(n6693), .X(n6688) );
  nand_x1_sg U7717 ( .A(n8214), .B(n7712), .X(n6690) );
  nand_x2_sg U7718 ( .A(n6651), .B(n6652), .X(n6650) );
  nand_x2_sg U7719 ( .A(n6653), .B(n6654), .X(n6649) );
  nand_x1_sg U7720 ( .A(n8214), .B(n7720), .X(n6651) );
  nand_x2_sg U7721 ( .A(n6573), .B(n6574), .X(n6572) );
  nand_x2_sg U7722 ( .A(n6575), .B(n6576), .X(n6571) );
  nand_x1_sg U7723 ( .A(n8214), .B(n7736), .X(n6573) );
  nand_x2_sg U7724 ( .A(n6534), .B(n6535), .X(n6533) );
  nand_x2_sg U7725 ( .A(n6536), .B(n6537), .X(n6532) );
  nand_x1_sg U7726 ( .A(n8214), .B(n7744), .X(n6534) );
  nand_x2_sg U7727 ( .A(n6456), .B(n6457), .X(n6455) );
  nand_x2_sg U7728 ( .A(n6458), .B(n6459), .X(n6454) );
  nand_x1_sg U7729 ( .A(n8214), .B(n7760), .X(n6456) );
  nand_x2_sg U7730 ( .A(n6417), .B(n6418), .X(n6416) );
  nand_x2_sg U7731 ( .A(n6419), .B(n6420), .X(n6415) );
  nand_x1_sg U7732 ( .A(n8214), .B(n7768), .X(n6417) );
  nand_x2_sg U7733 ( .A(n6339), .B(n6340), .X(n6338) );
  nand_x2_sg U7734 ( .A(n6341), .B(n6342), .X(n6337) );
  nand_x1_sg U7735 ( .A(n8214), .B(n7622), .X(n6339) );
  nand_x2_sg U7736 ( .A(n6300), .B(n6301), .X(n6299) );
  nand_x2_sg U7737 ( .A(n6302), .B(n6303), .X(n6298) );
  nand_x1_sg U7738 ( .A(n8214), .B(n7630), .X(n6300) );
  nand_x2_sg U7739 ( .A(n6222), .B(n6223), .X(n6221) );
  nand_x2_sg U7740 ( .A(n6224), .B(n6225), .X(n6220) );
  nand_x1_sg U7741 ( .A(n8214), .B(n7646), .X(n6222) );
  nand_x2_sg U7742 ( .A(n6183), .B(n6184), .X(n6182) );
  nand_x2_sg U7743 ( .A(n6185), .B(n6186), .X(n6181) );
  nand_x1_sg U7744 ( .A(n8214), .B(n7654), .X(n6183) );
  nand_x2_sg U7745 ( .A(n6105), .B(n6106), .X(n6104) );
  nand_x2_sg U7746 ( .A(n6107), .B(n6108), .X(n6103) );
  nand_x1_sg U7747 ( .A(n8214), .B(n7670), .X(n6105) );
  nand_x2_sg U7748 ( .A(n6046), .B(n6047), .X(n6045) );
  nand_x2_sg U7749 ( .A(n6050), .B(n6051), .X(n6044) );
  nand_x1_sg U7750 ( .A(n8214), .B(n7678), .X(n6046) );
  nand_x1_sg U7751 ( .A(n8212), .B(n7482), .X(n6732) );
  nand_x1_sg U7752 ( .A(n8212), .B(n7524), .X(n6615) );
  nand_x1_sg U7753 ( .A(n8212), .B(n7566), .X(n6498) );
  nand_x1_sg U7754 ( .A(n8212), .B(n7608), .X(n6381) );
  nand_x1_sg U7755 ( .A(n6052), .B(n7370), .X(n6264) );
  nand_x1_sg U7756 ( .A(n8212), .B(n7412), .X(n6147) );
  nand_x2_sg U7757 ( .A(n6729), .B(n6730), .X(n6728) );
  nand_x2_sg U7758 ( .A(n6731), .B(n6732), .X(n6727) );
  nand_x1_sg U7759 ( .A(n8214), .B(n7704), .X(n6729) );
  nand_x2_sg U7760 ( .A(n6612), .B(n6613), .X(n6611) );
  nand_x2_sg U7761 ( .A(n6614), .B(n6615), .X(n6610) );
  nand_x1_sg U7762 ( .A(n8214), .B(n7728), .X(n6612) );
  nand_x2_sg U7763 ( .A(n6495), .B(n6496), .X(n6494) );
  nand_x2_sg U7764 ( .A(n6497), .B(n6498), .X(n6493) );
  nand_x1_sg U7765 ( .A(n8214), .B(n7752), .X(n6495) );
  nand_x2_sg U7766 ( .A(n6378), .B(n6379), .X(n6377) );
  nand_x2_sg U7767 ( .A(n6380), .B(n6381), .X(n6376) );
  nand_x1_sg U7768 ( .A(n8214), .B(n7776), .X(n6378) );
  nand_x2_sg U7769 ( .A(n6261), .B(n6262), .X(n6260) );
  nand_x2_sg U7770 ( .A(n6263), .B(n6264), .X(n6259) );
  nand_x1_sg U7771 ( .A(n6049), .B(n7638), .X(n6261) );
  nand_x2_sg U7772 ( .A(n6144), .B(n6145), .X(n6143) );
  nand_x2_sg U7773 ( .A(n6146), .B(n6147), .X(n6142) );
  nand_x1_sg U7774 ( .A(n8214), .B(n7662), .X(n6144) );
  nand_x1_sg U7775 ( .A(n8180), .B(n7464), .X(n6842) );
  nand_x1_sg U7776 ( .A(n8181), .B(n7478), .X(n6794) );
  nand_x1_sg U7777 ( .A(n8182), .B(n7492), .X(n6755) );
  nand_x1_sg U7778 ( .A(n8182), .B(n7506), .X(n6716) );
  nand_x1_sg U7779 ( .A(n8180), .B(n7352), .X(n6365) );
  nand_x1_sg U7780 ( .A(n8181), .B(n7366), .X(n6326) );
  nand_x1_sg U7781 ( .A(n8182), .B(n7380), .X(n6287) );
  nand_x1_sg U7782 ( .A(n8181), .B(n7394), .X(n6248) );
  nand_x1_sg U7783 ( .A(n8180), .B(n7408), .X(n6209) );
  nand_x1_sg U7784 ( .A(n8181), .B(n7422), .X(n6170) );
  nand_x1_sg U7785 ( .A(n8182), .B(n7436), .X(n6131) );
  nand_x1_sg U7786 ( .A(n8180), .B(n7450), .X(n6087) );
  nand_x2_sg U7787 ( .A(n6844), .B(n6845), .X(n6840) );
  nand_x2_sg U7788 ( .A(n6842), .B(n6843), .X(n6841) );
  nand_x1_sg U7789 ( .A(n8170), .B(n7690), .X(n6845) );
  nand_x2_sg U7790 ( .A(n6796), .B(n6797), .X(n6792) );
  nand_x2_sg U7791 ( .A(n6794), .B(n6795), .X(n6793) );
  nand_x1_sg U7792 ( .A(n8171), .B(n7698), .X(n6797) );
  nand_x2_sg U7793 ( .A(n6757), .B(n6758), .X(n6753) );
  nand_x2_sg U7794 ( .A(n6755), .B(n6756), .X(n6754) );
  nand_x1_sg U7795 ( .A(n8172), .B(n7706), .X(n6758) );
  nand_x2_sg U7796 ( .A(n6718), .B(n6719), .X(n6714) );
  nand_x2_sg U7797 ( .A(n6716), .B(n6717), .X(n6715) );
  nand_x1_sg U7798 ( .A(n8172), .B(n7714), .X(n6719) );
  nand_x2_sg U7799 ( .A(n6367), .B(n6368), .X(n6363) );
  nand_x2_sg U7800 ( .A(n6365), .B(n6366), .X(n6364) );
  nand_x1_sg U7801 ( .A(n8170), .B(n7624), .X(n6368) );
  nand_x2_sg U7802 ( .A(n6328), .B(n6329), .X(n6324) );
  nand_x2_sg U7803 ( .A(n6326), .B(n6327), .X(n6325) );
  nand_x1_sg U7804 ( .A(n8171), .B(n7632), .X(n6329) );
  nand_x2_sg U7805 ( .A(n6289), .B(n6290), .X(n6285) );
  nand_x2_sg U7806 ( .A(n6287), .B(n6288), .X(n6286) );
  nand_x1_sg U7807 ( .A(n8172), .B(n7640), .X(n6290) );
  nand_x2_sg U7808 ( .A(n6250), .B(n6251), .X(n6246) );
  nand_x2_sg U7809 ( .A(n6248), .B(n6249), .X(n6247) );
  nand_x1_sg U7810 ( .A(n8170), .B(n7648), .X(n6251) );
  nand_x2_sg U7811 ( .A(n6211), .B(n6212), .X(n6207) );
  nand_x2_sg U7812 ( .A(n6209), .B(n6210), .X(n6208) );
  nand_x1_sg U7813 ( .A(n8170), .B(n7656), .X(n6212) );
  nand_x2_sg U7814 ( .A(n6172), .B(n6173), .X(n6168) );
  nand_x2_sg U7815 ( .A(n6170), .B(n6171), .X(n6169) );
  nand_x1_sg U7816 ( .A(n8171), .B(n7664), .X(n6173) );
  nand_x2_sg U7817 ( .A(n6133), .B(n6134), .X(n6129) );
  nand_x2_sg U7818 ( .A(n6131), .B(n6132), .X(n6130) );
  nand_x1_sg U7819 ( .A(n8172), .B(n7672), .X(n6134) );
  nand_x2_sg U7820 ( .A(n6091), .B(n6092), .X(n6085) );
  nand_x2_sg U7821 ( .A(n6087), .B(n6088), .X(n6086) );
  nand_x1_sg U7822 ( .A(n8171), .B(n7680), .X(n6092) );
  nand_x1_sg U7823 ( .A(n8183), .B(n7520), .X(n6677) );
  nand_x1_sg U7824 ( .A(n8184), .B(n7534), .X(n6638) );
  nand_x1_sg U7825 ( .A(n8185), .B(n7548), .X(n6599) );
  nand_x1_sg U7826 ( .A(n8186), .B(n7562), .X(n6560) );
  nand_x1_sg U7827 ( .A(n8183), .B(n7576), .X(n6521) );
  nand_x1_sg U7828 ( .A(n8184), .B(n7590), .X(n6482) );
  nand_x1_sg U7829 ( .A(n8185), .B(n7604), .X(n6443) );
  nand_x1_sg U7830 ( .A(n8186), .B(n7618), .X(n6404) );
  nand_x2_sg U7831 ( .A(n6679), .B(n6680), .X(n6675) );
  nand_x2_sg U7832 ( .A(n6677), .B(n6678), .X(n6676) );
  nand_x1_sg U7833 ( .A(n8174), .B(n7722), .X(n6680) );
  nand_x2_sg U7834 ( .A(n6640), .B(n6641), .X(n6636) );
  nand_x2_sg U7835 ( .A(n6638), .B(n6639), .X(n6637) );
  nand_x1_sg U7836 ( .A(n8175), .B(n7730), .X(n6641) );
  nand_x2_sg U7837 ( .A(n6601), .B(n6602), .X(n6597) );
  nand_x2_sg U7838 ( .A(n6599), .B(n6600), .X(n6598) );
  nand_x1_sg U7839 ( .A(n8176), .B(n7738), .X(n6602) );
  nand_x2_sg U7840 ( .A(n6562), .B(n6563), .X(n6558) );
  nand_x2_sg U7841 ( .A(n6560), .B(n6561), .X(n6559) );
  nand_x1_sg U7842 ( .A(n8177), .B(n7746), .X(n6563) );
  nand_x2_sg U7843 ( .A(n6523), .B(n6524), .X(n6519) );
  nand_x2_sg U7844 ( .A(n6521), .B(n6522), .X(n6520) );
  nand_x1_sg U7845 ( .A(n8174), .B(n7754), .X(n6524) );
  nand_x2_sg U7846 ( .A(n6484), .B(n6485), .X(n6480) );
  nand_x2_sg U7847 ( .A(n6482), .B(n6483), .X(n6481) );
  nand_x1_sg U7848 ( .A(n8175), .B(n7762), .X(n6485) );
  nand_x2_sg U7849 ( .A(n6445), .B(n6446), .X(n6441) );
  nand_x2_sg U7850 ( .A(n6443), .B(n6444), .X(n6442) );
  nand_x1_sg U7851 ( .A(n8176), .B(n7770), .X(n6446) );
  nand_x2_sg U7852 ( .A(n6406), .B(n6407), .X(n6402) );
  nand_x2_sg U7853 ( .A(n6404), .B(n6405), .X(n6403) );
  nand_x1_sg U7854 ( .A(n8177), .B(n7778), .X(n6407) );
  nor_x1_sg U7855 ( .A(n7338), .B(n5464), .X(n6016) );
  nor_x1_sg U7856 ( .A(n5464), .B(n4909), .X(n5574) );
  nor_x1_sg U7857 ( .A(n8106), .B(n5464), .X(n5463) );
  nand_x4_sg U7858 ( .A(n6017), .B(n6018), .X(n5850) );
  nor_x1_sg U7859 ( .A(reset), .B(full), .X(n6018) );
  nor_x1_sg U7860 ( .A(n6019), .B(n4890), .X(n6017) );
  nand_x1_sg U7861 ( .A(n7620), .B(n8253), .X(n5297) );
  nand_x1_sg U7862 ( .A(n7778), .B(n8221), .X(n5291) );
  nand_x1_sg U7863 ( .A(n7618), .B(n8241), .X(n5289) );
  nand_x1_sg U7864 ( .A(n7770), .B(n8221), .X(n5935) );
  nand_x1_sg U7865 ( .A(n7604), .B(n8241), .X(n5541) );
  nand_x1_sg U7866 ( .A(n7762), .B(n8222), .X(n5957) );
  nand_x1_sg U7867 ( .A(n7578), .B(n8253), .X(n5342) );
  nand_x1_sg U7868 ( .A(n7754), .B(n8221), .X(n5929) );
  nand_x1_sg U7869 ( .A(n7576), .B(n8241), .X(n5547) );
  nand_x1_sg U7870 ( .A(n7746), .B(n8221), .X(n5947) );
  nand_x1_sg U7871 ( .A(n7562), .B(n8242), .X(n5545) );
  nand_x1_sg U7872 ( .A(n7550), .B(n8254), .X(n5346) );
  nand_x1_sg U7873 ( .A(n7536), .B(n8253), .X(n5324) );
  nand_x1_sg U7874 ( .A(n7730), .B(n8222), .X(n5939) );
  nand_x1_sg U7875 ( .A(n7522), .B(n8254), .X(n5340) );
  nand_x1_sg U7876 ( .A(n7722), .B(n8222), .X(n5945) );
  nand_x1_sg U7877 ( .A(n7508), .B(n8253), .X(n5318) );
  nand_x1_sg U7878 ( .A(n7714), .B(n8222), .X(n5933) );
  nand_x1_sg U7879 ( .A(n7494), .B(n8253), .X(n5330) );
  nand_x1_sg U7880 ( .A(n7706), .B(n8221), .X(n5953) );
  nand_x1_sg U7881 ( .A(n7480), .B(n8254), .X(n5334) );
  nand_x1_sg U7882 ( .A(n7478), .B(n8242), .X(n5569) );
  nand_x1_sg U7883 ( .A(n7466), .B(n8254), .X(n5234) );
  nand_x1_sg U7884 ( .A(n7690), .B(n8222), .X(n5237) );
  nand_x1_sg U7885 ( .A(n7464), .B(n8242), .X(n5192) );
  nand_x1_sg U7886 ( .A(n7452), .B(n8254), .X(n5328) );
  nand_x1_sg U7887 ( .A(n7450), .B(n8242), .X(n5563) );
  nand_x1_sg U7888 ( .A(n7438), .B(n8254), .X(n5322) );
  nand_x1_sg U7889 ( .A(n7436), .B(n8241), .X(n5553) );
  nand_x1_sg U7890 ( .A(n7664), .B(n8221), .X(n5941) );
  nand_x1_sg U7891 ( .A(n7422), .B(n8241), .X(n5559) );
  nand_x1_sg U7892 ( .A(n7408), .B(n8241), .X(n5571) );
  nand_x1_sg U7893 ( .A(n7648), .B(n8221), .X(n5959) );
  nand_x1_sg U7894 ( .A(n7394), .B(n8242), .X(n5539) );
  nand_x1_sg U7895 ( .A(n7382), .B(n8254), .X(n5316) );
  nand_x1_sg U7896 ( .A(n7380), .B(n8242), .X(n5551) );
  nand_x1_sg U7897 ( .A(n7368), .B(n8253), .X(n5336) );
  nand_x1_sg U7898 ( .A(n7632), .B(n8222), .X(n5951) );
  nand_x1_sg U7899 ( .A(n7366), .B(n8242), .X(n5557) );
  nand_x1_sg U7900 ( .A(n7354), .B(n8253), .X(n5348) );
  nand_x1_sg U7901 ( .A(n7624), .B(n8222), .X(n5927) );
  nand_x1_sg U7902 ( .A(n7352), .B(n8241), .X(n5565) );
  nand_x1_sg U7903 ( .A(n7780), .B(n8249), .X(n5307) );
  nand_x1_sg U7904 ( .A(n7940), .B(n8219), .X(n5305) );
  nand_x1_sg U7905 ( .A(n7938), .B(n8245), .X(n5293) );
  nand_x1_sg U7906 ( .A(n7772), .B(n8250), .X(n5396) );
  nand_x1_sg U7907 ( .A(n7936), .B(n8219), .X(n5967) );
  nand_x1_sg U7908 ( .A(n7934), .B(n8246), .X(n5473) );
  nand_x1_sg U7909 ( .A(n7932), .B(n8220), .X(n6009) );
  nand_x1_sg U7910 ( .A(n7930), .B(n8245), .X(n5499) );
  nand_x1_sg U7911 ( .A(n7756), .B(n8249), .X(n5416) );
  nand_x1_sg U7912 ( .A(n7926), .B(n8246), .X(n5491) );
  nand_x1_sg U7913 ( .A(n7740), .B(n8250), .X(n5420) );
  nand_x1_sg U7914 ( .A(n7920), .B(n8219), .X(n5985) );
  nand_x1_sg U7915 ( .A(n7724), .B(n8250), .X(n5414) );
  nand_x1_sg U7916 ( .A(n7912), .B(n8219), .X(n6012) );
  nand_x1_sg U7917 ( .A(n7908), .B(n8220), .X(n5964) );
  nand_x1_sg U7918 ( .A(n7708), .B(n8250), .X(n5408) );
  nand_x1_sg U7919 ( .A(n7904), .B(n8220), .X(n5982) );
  nand_x1_sg U7920 ( .A(n7902), .B(n8245), .X(n5493) );
  nand_x1_sg U7921 ( .A(n7700), .B(n8249), .X(n5404) );
  nand_x1_sg U7922 ( .A(n7900), .B(n8220), .X(n6000) );
  nand_x1_sg U7923 ( .A(n7692), .B(n8250), .X(n5195) );
  nand_x1_sg U7924 ( .A(n7896), .B(n8220), .X(n5240) );
  nand_x1_sg U7925 ( .A(n7894), .B(n8246), .X(n5204) );
  nand_x1_sg U7926 ( .A(n7682), .B(n8249), .X(n5410) );
  nand_x1_sg U7927 ( .A(n7892), .B(n8220), .X(n5973) );
  nand_x1_sg U7928 ( .A(n7890), .B(n8246), .X(n5479) );
  nand_x1_sg U7929 ( .A(n7674), .B(n8249), .X(n5398) );
  nand_x1_sg U7930 ( .A(n7886), .B(n8245), .X(n5475) );
  nand_x1_sg U7931 ( .A(n7666), .B(n8250), .X(n5402) );
  nand_x1_sg U7932 ( .A(n7884), .B(n8220), .X(n5991) );
  nand_x1_sg U7933 ( .A(n7882), .B(n8245), .X(n5481) );
  nand_x1_sg U7934 ( .A(n7880), .B(n8219), .X(n6003) );
  nand_x1_sg U7935 ( .A(n7878), .B(n8245), .X(n5487) );
  nand_x1_sg U7936 ( .A(n7650), .B(n8250), .X(n5390) );
  nand_x1_sg U7937 ( .A(n7874), .B(n8246), .X(n5467) );
  nand_x1_sg U7938 ( .A(n7642), .B(n8249), .X(n5392) );
  nand_x1_sg U7939 ( .A(n7870), .B(n8245), .X(n5469) );
  nand_x1_sg U7940 ( .A(n7868), .B(n8219), .X(n5994) );
  nand_x1_sg U7941 ( .A(n7866), .B(n8246), .X(n5485) );
  nand_x1_sg U7942 ( .A(n7626), .B(n8249), .X(n5422) );
  nand_x1_sg U7943 ( .A(n7864), .B(n8219), .X(n5976) );
  nand_x1_sg U7944 ( .A(n7862), .B(n8246), .X(n5497) );
  nand_x1_sg U7945 ( .A(n7326), .B(n8247), .X(n5281) );
  nand_x1_sg U7946 ( .A(n7858), .B(n8223), .X(n5299) );
  nand_x1_sg U7947 ( .A(n7324), .B(n8247), .X(n5441) );
  nand_x1_sg U7948 ( .A(n7854), .B(n8223), .X(n5898) );
  nand_x1_sg U7949 ( .A(n7850), .B(n8223), .X(n5922) );
  nand_x1_sg U7950 ( .A(n7846), .B(n8223), .X(n5892) );
  nand_x1_sg U7951 ( .A(n7296), .B(n8248), .X(n5433) );
  nand_x1_sg U7952 ( .A(n7838), .B(n8223), .X(n5916) );
  nand_x1_sg U7953 ( .A(n7834), .B(n8224), .X(n5902) );
  nand_x1_sg U7954 ( .A(n7316), .B(n8248), .X(n5457) );
  nand_x1_sg U7955 ( .A(n7294), .B(n8248), .X(n5439) );
  nand_x1_sg U7956 ( .A(n7826), .B(n8224), .X(n5896) );
  nand_x1_sg U7957 ( .A(n7314), .B(n8248), .X(n5445) );
  nand_x1_sg U7958 ( .A(n7822), .B(n8223), .X(n5904) );
  nand_x1_sg U7959 ( .A(n7312), .B(n8248), .X(n5451) );
  nand_x1_sg U7960 ( .A(n7818), .B(n8224), .X(n5908) );
  nand_x1_sg U7961 ( .A(n7292), .B(n8248), .X(n5243) );
  nand_x1_sg U7962 ( .A(n7814), .B(n8224), .X(n5231) );
  nand_x1_sg U7963 ( .A(n7310), .B(n8247), .X(n5447) );
  nand_x1_sg U7964 ( .A(n7810), .B(n8224), .X(n5890) );
  nand_x1_sg U7965 ( .A(n7290), .B(n8248), .X(n5427) );
  nand_x1_sg U7966 ( .A(n7306), .B(n8247), .X(n5453) );
  nand_x1_sg U7967 ( .A(n7798), .B(n8224), .X(n5914) );
  nand_x1_sg U7968 ( .A(n7288), .B(n8247), .X(n5435) );
  nand_x1_sg U7969 ( .A(n7794), .B(n8224), .X(n5920) );
  nand_x1_sg U7970 ( .A(n7302), .B(n8247), .X(n5429) );
  nand_x1_sg U7971 ( .A(n7786), .B(n8223), .X(n5910) );
  nand_x1_sg U7972 ( .A(n7286), .B(n8247), .X(n5459) );
  nand_x1_sg U7973 ( .A(n7860), .B(n8225), .X(n5303) );
  nand_x1_sg U7974 ( .A(n7774), .B(n8251), .X(n5311) );
  nand_x1_sg U7975 ( .A(n7856), .B(n8225), .X(n5861) );
  nand_x1_sg U7976 ( .A(n7852), .B(n8225), .X(n5885) );
  nand_x1_sg U7977 ( .A(n7758), .B(n8252), .X(n5378) );
  nand_x1_sg U7978 ( .A(n7848), .B(n8225), .X(n5855) );
  nand_x1_sg U7979 ( .A(n7750), .B(n8252), .X(n5372) );
  nand_x1_sg U7980 ( .A(n7742), .B(n8252), .X(n5354) );
  nand_x1_sg U7981 ( .A(n7840), .B(n8225), .X(n5879) );
  nand_x1_sg U7982 ( .A(n7836), .B(n8226), .X(n5865) );
  nand_x1_sg U7983 ( .A(n7726), .B(n8251), .X(n5368) );
  nand_x1_sg U7984 ( .A(n7718), .B(n8251), .X(n5386) );
  nand_x1_sg U7985 ( .A(n7828), .B(n8226), .X(n5859) );
  nand_x1_sg U7986 ( .A(n7702), .B(n8251), .X(n5362) );
  nand_x1_sg U7987 ( .A(n7820), .B(n8226), .X(n5871) );
  nand_x1_sg U7988 ( .A(n7694), .B(n8252), .X(n5384) );
  nand_x1_sg U7989 ( .A(n7816), .B(n8226), .X(n5198) );
  nand_x1_sg U7990 ( .A(n7686), .B(n8252), .X(n5219) );
  nand_x1_sg U7991 ( .A(n7812), .B(n8226), .X(n5853) );
  nand_x1_sg U7992 ( .A(n7668), .B(n8252), .X(n5366) );
  nand_x1_sg U7993 ( .A(n7804), .B(n8225), .X(n5867) );
  nand_x1_sg U7994 ( .A(n7660), .B(n8251), .X(n5374) );
  nand_x1_sg U7995 ( .A(n7800), .B(n8226), .X(n5877) );
  nand_x1_sg U7996 ( .A(n7652), .B(n8252), .X(n5360) );
  nand_x1_sg U7997 ( .A(n7796), .B(n8226), .X(n5883) );
  nand_x1_sg U7998 ( .A(n7636), .B(n8251), .X(n5380) );
  nand_x1_sg U7999 ( .A(n7788), .B(n8225), .X(n5873) );
  nand_x1_sg U8000 ( .A(n7628), .B(n8251), .X(n5356) );
  nand_x1_sg U8001 ( .A(n8020), .B(n8243), .X(n5279) );
  nand_x1_sg U8002 ( .A(n8016), .B(n8243), .X(n5511) );
  nand_x1_sg U8003 ( .A(n8012), .B(n8243), .X(n5505) );
  nand_x1_sg U8004 ( .A(n8008), .B(n8244), .X(n5521) );
  nand_x1_sg U8005 ( .A(n8004), .B(n8244), .X(n5527) );
  nand_x1_sg U8006 ( .A(n8000), .B(n8244), .X(n5533) );
  nand_x1_sg U8007 ( .A(n7996), .B(n8244), .X(n5515) );
  nand_x1_sg U8008 ( .A(n7988), .B(n8244), .X(n5509) );
  nand_x1_sg U8009 ( .A(n7984), .B(n8243), .X(n5523) );
  nand_x1_sg U8010 ( .A(n7976), .B(n8244), .X(n5225) );
  nand_x1_sg U8011 ( .A(n7964), .B(n8243), .X(n5529) );
  nand_x1_sg U8012 ( .A(n7960), .B(n8244), .X(n5503) );
  nand_x1_sg U8013 ( .A(n7956), .B(n8243), .X(n5535) );
  nand_x1_sg U8014 ( .A(n7944), .B(n8243), .X(n5517) );
  nand_x1_sg U8015 ( .A(n8092), .B(n8258), .X(n5116) );
  nand_x1_sg U8016 ( .A(n8088), .B(n8258), .X(n5098) );
  nand_x1_sg U8017 ( .A(n8072), .B(n8257), .X(n5118) );
  nand_x1_sg U8018 ( .A(n8068), .B(n8257), .X(n5082) );
  nand_x1_sg U8019 ( .A(n8064), .B(n8257), .X(n5094) );
  nand_x1_sg U8020 ( .A(n8060), .B(n8258), .X(n5110) );
  nand_x1_sg U8021 ( .A(n8056), .B(n8257), .X(n5088) );
  nand_x1_sg U8022 ( .A(n8052), .B(n8257), .X(n5100) );
  nand_x1_sg U8023 ( .A(n8048), .B(n8258), .X(n5104) );
  nand_x1_sg U8024 ( .A(n8044), .B(n8257), .X(n5106) );
  nand_x1_sg U8025 ( .A(n8040), .B(n8257), .X(n5112) );
  nand_x1_sg U8026 ( .A(n8036), .B(n8258), .X(n5092) );
  nand_x1_sg U8027 ( .A(n8032), .B(n8258), .X(n5079) );
  nand_x1_sg U8028 ( .A(n8028), .B(n8258), .X(n5086) );
  nand_x1_sg U8029 ( .A(n7606), .B(n5236), .X(n5320) );
  nand_x1_sg U8030 ( .A(n7592), .B(n5236), .X(n5344) );
  nand_x1_sg U8031 ( .A(n7564), .B(n5236), .X(n5326) );
  nand_x1_sg U8032 ( .A(n7738), .B(n5239), .X(n5955) );
  nand_x1_sg U8033 ( .A(n7698), .B(n5239), .X(n5949) );
  nand_x1_sg U8034 ( .A(n7680), .B(n5239), .X(n5925) );
  nand_x1_sg U8035 ( .A(n7672), .B(n5239), .X(n5937) );
  nand_x1_sg U8036 ( .A(n7424), .B(n5236), .X(n5332) );
  nand_x1_sg U8037 ( .A(n7410), .B(n5236), .X(n5338) );
  nand_x1_sg U8038 ( .A(n7656), .B(n5239), .X(n5943) );
  nand_x1_sg U8039 ( .A(n7396), .B(n5236), .X(n5314) );
  nand_x1_sg U8040 ( .A(n7640), .B(n5239), .X(n5931) );
  nand_x1_sg U8041 ( .A(n7764), .B(n5197), .X(n5418) );
  nand_x1_sg U8042 ( .A(n7928), .B(n5242), .X(n5970) );
  nand_x1_sg U8043 ( .A(n7748), .B(n5197), .X(n5388) );
  nand_x1_sg U8044 ( .A(n7924), .B(n5242), .X(n5997) );
  nand_x1_sg U8045 ( .A(n7732), .B(n5197), .X(n5400) );
  nand_x1_sg U8046 ( .A(n7916), .B(n5242), .X(n6006) );
  nand_x1_sg U8047 ( .A(n7716), .B(n5197), .X(n5394) );
  nand_x1_sg U8048 ( .A(n7888), .B(n5242), .X(n5988) );
  nand_x1_sg U8049 ( .A(n7658), .B(n5197), .X(n5412) );
  nand_x1_sg U8050 ( .A(n7876), .B(n5242), .X(n5979) );
  nand_x1_sg U8051 ( .A(n7872), .B(n5242), .X(n5961) );
  nand_x1_sg U8052 ( .A(n7634), .B(n5197), .X(n5406) );
  nand_x1_sg U8053 ( .A(n7298), .B(n5246), .X(n5449) );
  nand_x1_sg U8054 ( .A(n7322), .B(n5246), .X(n5425) );
  nand_x1_sg U8055 ( .A(n7320), .B(n5246), .X(n5437) );
  nand_x1_sg U8056 ( .A(n7842), .B(n5233), .X(n5912) );
  nand_x1_sg U8057 ( .A(n7318), .B(n5246), .X(n5455) );
  nand_x1_sg U8058 ( .A(n7830), .B(n5233), .X(n5888) );
  nand_x1_sg U8059 ( .A(n7806), .B(n5233), .X(n5900) );
  nand_x1_sg U8060 ( .A(n7308), .B(n5246), .X(n5431) );
  nand_x1_sg U8061 ( .A(n7802), .B(n5233), .X(n5906) );
  nand_x1_sg U8062 ( .A(n7304), .B(n5246), .X(n5443) );
  nand_x1_sg U8063 ( .A(n7790), .B(n5233), .X(n5894) );
  nand_x1_sg U8064 ( .A(n7782), .B(n5233), .X(n5918) );
  nand_x1_sg U8065 ( .A(n7766), .B(n5221), .X(n5364) );
  nand_x1_sg U8066 ( .A(n7844), .B(n5200), .X(n5869) );
  nand_x1_sg U8067 ( .A(n7734), .B(n5221), .X(n5358) );
  nand_x1_sg U8068 ( .A(n7832), .B(n5200), .X(n5851) );
  nand_x1_sg U8069 ( .A(n7710), .B(n5221), .X(n5370) );
  nand_x1_sg U8070 ( .A(n7824), .B(n5200), .X(n5875) );
  nand_x1_sg U8071 ( .A(n7684), .B(n5221), .X(n5352) );
  nand_x1_sg U8072 ( .A(n7676), .B(n5221), .X(n5382) );
  nand_x1_sg U8073 ( .A(n7808), .B(n5200), .X(n5863) );
  nand_x1_sg U8074 ( .A(n7644), .B(n5221), .X(n5376) );
  nand_x1_sg U8075 ( .A(n7792), .B(n5200), .X(n5857) );
  nand_x1_sg U8076 ( .A(n7784), .B(n5200), .X(n5881) );
  nand_x1_sg U8077 ( .A(n8100), .B(n5081), .X(n5090) );
  nand_x1_sg U8078 ( .A(n7590), .B(n5194), .X(n5567) );
  nand_x1_sg U8079 ( .A(n7548), .B(n5194), .X(n5561) );
  nand_x1_sg U8080 ( .A(n7534), .B(n5194), .X(n5537) );
  nand_x1_sg U8081 ( .A(n7520), .B(n5194), .X(n5549) );
  nand_x1_sg U8082 ( .A(n7506), .B(n5194), .X(n5555) );
  nand_x1_sg U8083 ( .A(n7492), .B(n5194), .X(n5543) );
  nand_x1_sg U8084 ( .A(n7922), .B(n5206), .X(n5465) );
  nand_x1_sg U8085 ( .A(n7918), .B(n5206), .X(n5495) );
  nand_x1_sg U8086 ( .A(n7914), .B(n5206), .X(n5477) );
  nand_x1_sg U8087 ( .A(n7910), .B(n5206), .X(n5489) );
  nand_x1_sg U8088 ( .A(n7906), .B(n5206), .X(n5471) );
  nand_x1_sg U8089 ( .A(n7898), .B(n5206), .X(n5483) );
  nand_x1_sg U8090 ( .A(n7992), .B(n5227), .X(n5519) );
  nand_x1_sg U8091 ( .A(n7980), .B(n5227), .X(n5501) );
  nand_x1_sg U8092 ( .A(n7972), .B(n5227), .X(n5525) );
  nand_x1_sg U8093 ( .A(n7968), .B(n5227), .X(n5513) );
  nand_x1_sg U8094 ( .A(n7952), .B(n5227), .X(n5507) );
  nand_x1_sg U8095 ( .A(n7948), .B(n5227), .X(n5531) );
  nand_x1_sg U8096 ( .A(n8096), .B(n5081), .X(n5084) );
  nand_x1_sg U8097 ( .A(n8084), .B(n5081), .X(n5108) );
  nand_x1_sg U8098 ( .A(n8080), .B(n5081), .X(n5096) );
  nand_x1_sg U8099 ( .A(n8076), .B(n5081), .X(n5114) );
  nand_x1_sg U8100 ( .A(n8024), .B(n5081), .X(n5102) );
  nand_x1_sg U8101 ( .A(n8098), .B(n8233), .X(n5301) );
  nand_x1_sg U8102 ( .A(n8094), .B(n8233), .X(n5712) );
  nand_x1_sg U8103 ( .A(n8090), .B(n8234), .X(n5734) );
  nand_x1_sg U8104 ( .A(n8086), .B(n8234), .X(n5722) );
  nand_x1_sg U8105 ( .A(n8074), .B(n8234), .X(n5716) );
  nand_x1_sg U8106 ( .A(n8066), .B(n8234), .X(n5710) );
  nand_x1_sg U8107 ( .A(n8062), .B(n8233), .X(n5724) );
  nand_x1_sg U8108 ( .A(n8058), .B(n8234), .X(n5728) );
  nand_x1_sg U8109 ( .A(n8054), .B(n8234), .X(n5216) );
  nand_x1_sg U8110 ( .A(n8050), .B(n8234), .X(n5704) );
  nand_x1_sg U8111 ( .A(n8042), .B(n8233), .X(n5718) );
  nand_x1_sg U8112 ( .A(n8034), .B(n8233), .X(n5736) );
  nand_x1_sg U8113 ( .A(n8026), .B(n8233), .X(n5730) );
  nand_x1_sg U8114 ( .A(n8022), .B(n8233), .X(n5706) );
  nand_x1_sg U8115 ( .A(n7776), .B(n8235), .X(n5295) );
  nand_x1_sg U8116 ( .A(n7768), .B(n8235), .X(n5670) );
  nand_x1_sg U8117 ( .A(n7760), .B(n8236), .X(n5698) );
  nand_x1_sg U8118 ( .A(n7752), .B(n8235), .X(n5682) );
  nand_x1_sg U8119 ( .A(n7736), .B(n8235), .X(n5676) );
  nand_x1_sg U8120 ( .A(n7720), .B(n8236), .X(n5686) );
  nand_x1_sg U8121 ( .A(n7712), .B(n8236), .X(n5668) );
  nand_x1_sg U8122 ( .A(n7704), .B(n8235), .X(n5688) );
  nand_x1_sg U8123 ( .A(n7696), .B(n8236), .X(n5692) );
  nand_x1_sg U8124 ( .A(n7688), .B(n8236), .X(n5213) );
  nand_x1_sg U8125 ( .A(n7662), .B(n8236), .X(n5674) );
  nand_x1_sg U8126 ( .A(n7654), .B(n8235), .X(n5694) );
  nand_x1_sg U8127 ( .A(n7646), .B(n8236), .X(n5680) );
  nand_x1_sg U8128 ( .A(n7622), .B(n8235), .X(n5700) );
  nand_x1_sg U8129 ( .A(n7608), .B(n8237), .X(n5285) );
  nand_x1_sg U8130 ( .A(n7594), .B(n8237), .X(n5640) );
  nand_x1_sg U8131 ( .A(n7566), .B(n8237), .X(n5634) );
  nand_x1_sg U8132 ( .A(n7552), .B(n8238), .X(n5650) );
  nand_x1_sg U8133 ( .A(n7538), .B(n8238), .X(n5662) );
  nand_x1_sg U8134 ( .A(n7524), .B(n8238), .X(n5644) );
  nand_x1_sg U8135 ( .A(n7510), .B(n8237), .X(n5646) );
  nand_x1_sg U8136 ( .A(n7496), .B(n8238), .X(n5638) );
  nand_x1_sg U8137 ( .A(n7482), .B(n8237), .X(n5658) );
  nand_x1_sg U8138 ( .A(n7454), .B(n8238), .X(n5207) );
  nand_x1_sg U8139 ( .A(n7412), .B(n8237), .X(n5652) );
  nand_x1_sg U8140 ( .A(n7384), .B(n8237), .X(n5664) );
  nand_x1_sg U8141 ( .A(n7356), .B(n8238), .X(n5656) );
  nand_x1_sg U8142 ( .A(n7342), .B(n8238), .X(n5632) );
  nand_x1_sg U8143 ( .A(n7610), .B(n8239), .X(n5309) );
  nand_x1_sg U8144 ( .A(n7568), .B(n8239), .X(n5621) );
  nand_x1_sg U8145 ( .A(n7540), .B(n8240), .X(n5625) );
  nand_x1_sg U8146 ( .A(n7526), .B(n8239), .X(n5603) );
  nand_x1_sg U8147 ( .A(n7512), .B(n8240), .X(n5619) );
  nand_x1_sg U8148 ( .A(n7498), .B(n8239), .X(n5597) );
  nand_x1_sg U8149 ( .A(n7484), .B(n8240), .X(n5613) );
  nand_x1_sg U8150 ( .A(n7470), .B(n8239), .X(n5609) );
  nand_x1_sg U8151 ( .A(n7456), .B(n8240), .X(n5222) );
  nand_x1_sg U8152 ( .A(n7442), .B(n8239), .X(n5615) );
  nand_x1_sg U8153 ( .A(n7428), .B(n8240), .X(n5601) );
  nand_x1_sg U8154 ( .A(n7414), .B(n8240), .X(n5607) );
  nand_x1_sg U8155 ( .A(n7372), .B(n8240), .X(n5595) );
  nand_x1_sg U8156 ( .A(n7344), .B(n8239), .X(n5627) );
  nand_x1_sg U8157 ( .A(n8082), .B(n5218), .X(n5726) );
  nand_x1_sg U8158 ( .A(n8078), .B(n5218), .X(n5732) );
  nand_x1_sg U8159 ( .A(n8070), .B(n5218), .X(n5702) );
  nand_x1_sg U8160 ( .A(n8046), .B(n5218), .X(n5714) );
  nand_x1_sg U8161 ( .A(n8038), .B(n5218), .X(n5720) );
  nand_x1_sg U8162 ( .A(n8030), .B(n5218), .X(n5708) );
  nand_x1_sg U8163 ( .A(n7744), .B(n5215), .X(n5672) );
  nand_x1_sg U8164 ( .A(n7728), .B(n5215), .X(n5696) );
  nand_x1_sg U8165 ( .A(n7678), .B(n5215), .X(n5684) );
  nand_x1_sg U8166 ( .A(n7670), .B(n5215), .X(n5690) );
  nand_x1_sg U8167 ( .A(n7638), .B(n5215), .X(n5666) );
  nand_x1_sg U8168 ( .A(n7630), .B(n5215), .X(n5678) );
  nand_x1_sg U8169 ( .A(n7580), .B(n5209), .X(n5660) );
  nand_x1_sg U8170 ( .A(n7468), .B(n5209), .X(n5654) );
  nand_x1_sg U8171 ( .A(n7440), .B(n5209), .X(n5630) );
  nand_x1_sg U8172 ( .A(n7426), .B(n5209), .X(n5642) );
  nand_x1_sg U8173 ( .A(n7398), .B(n5209), .X(n5648) );
  nand_x1_sg U8174 ( .A(n7370), .B(n5209), .X(n5636) );
  nand_x1_sg U8175 ( .A(n7596), .B(n5224), .X(n5599) );
  nand_x1_sg U8176 ( .A(n7582), .B(n5224), .X(n5623) );
  nand_x1_sg U8177 ( .A(n7554), .B(n5224), .X(n5605) );
  nand_x1_sg U8178 ( .A(n7400), .B(n5224), .X(n5617) );
  nand_x1_sg U8179 ( .A(n7386), .B(n5224), .X(n5593) );
  nand_x1_sg U8180 ( .A(n7358), .B(n5224), .X(n5611) );
  nor_x1_sg U8181 ( .A(n6837), .B(n6838), .X(n6835) );
  nor_x1_sg U8182 ( .A(n6790), .B(n6791), .X(n6788) );
  nor_x1_sg U8183 ( .A(n6712), .B(n6713), .X(n6710) );
  nor_x1_sg U8184 ( .A(n6673), .B(n6674), .X(n6671) );
  nor_x1_sg U8185 ( .A(n6595), .B(n6596), .X(n6593) );
  nor_x1_sg U8186 ( .A(n6556), .B(n6557), .X(n6554) );
  nor_x1_sg U8187 ( .A(n6478), .B(n6479), .X(n6476) );
  nor_x1_sg U8188 ( .A(n6439), .B(n6440), .X(n6437) );
  nor_x1_sg U8189 ( .A(n6361), .B(n6362), .X(n6359) );
  nor_x1_sg U8190 ( .A(n6322), .B(n6323), .X(n6320) );
  nor_x1_sg U8191 ( .A(n6244), .B(n6245), .X(n6242) );
  nor_x1_sg U8192 ( .A(n6205), .B(n6206), .X(n6203) );
  nor_x1_sg U8193 ( .A(n6127), .B(n6128), .X(n6125) );
  nor_x1_sg U8194 ( .A(n6081), .B(n6082), .X(n6078) );
  nand_x2_sg U8195 ( .A(n6833), .B(n6834), .X(n6832) );
  nand_x2_sg U8196 ( .A(n6835), .B(n6836), .X(n6831) );
  nand_x1_sg U8197 ( .A(n8195), .B(n7686), .X(n6833) );
  nand_x2_sg U8198 ( .A(n6786), .B(n6787), .X(n6785) );
  nand_x2_sg U8199 ( .A(n6788), .B(n6789), .X(n6784) );
  nand_x1_sg U8200 ( .A(n8195), .B(n7694), .X(n6786) );
  nand_x2_sg U8201 ( .A(n6708), .B(n6709), .X(n6707) );
  nand_x2_sg U8202 ( .A(n6710), .B(n6711), .X(n6706) );
  nand_x1_sg U8203 ( .A(n8195), .B(n7710), .X(n6708) );
  nand_x2_sg U8204 ( .A(n6669), .B(n6670), .X(n6668) );
  nand_x2_sg U8205 ( .A(n6671), .B(n6672), .X(n6667) );
  nand_x1_sg U8206 ( .A(n8195), .B(n7718), .X(n6669) );
  nand_x2_sg U8207 ( .A(n6591), .B(n6592), .X(n6590) );
  nand_x2_sg U8208 ( .A(n6593), .B(n6594), .X(n6589) );
  nand_x1_sg U8209 ( .A(n8195), .B(n7734), .X(n6591) );
  nand_x2_sg U8210 ( .A(n6552), .B(n6553), .X(n6551) );
  nand_x2_sg U8211 ( .A(n6554), .B(n6555), .X(n6550) );
  nand_x1_sg U8212 ( .A(n8195), .B(n7742), .X(n6552) );
  nand_x2_sg U8213 ( .A(n6474), .B(n6475), .X(n6473) );
  nand_x2_sg U8214 ( .A(n6476), .B(n6477), .X(n6472) );
  nand_x1_sg U8215 ( .A(n8195), .B(n7758), .X(n6474) );
  nand_x2_sg U8216 ( .A(n6435), .B(n6436), .X(n6434) );
  nand_x2_sg U8217 ( .A(n6437), .B(n6438), .X(n6433) );
  nand_x1_sg U8218 ( .A(n8195), .B(n7766), .X(n6435) );
  nand_x2_sg U8219 ( .A(n6357), .B(n6358), .X(n6356) );
  nand_x2_sg U8220 ( .A(n6359), .B(n6360), .X(n6355) );
  nand_x1_sg U8221 ( .A(n8195), .B(n7628), .X(n6357) );
  nand_x2_sg U8222 ( .A(n6318), .B(n6319), .X(n6317) );
  nand_x2_sg U8223 ( .A(n6320), .B(n6321), .X(n6316) );
  nand_x1_sg U8224 ( .A(n8195), .B(n7636), .X(n6318) );
  nand_x2_sg U8225 ( .A(n6240), .B(n6241), .X(n6239) );
  nand_x2_sg U8226 ( .A(n6242), .B(n6243), .X(n6238) );
  nand_x1_sg U8227 ( .A(n8195), .B(n7652), .X(n6240) );
  nand_x2_sg U8228 ( .A(n6201), .B(n6202), .X(n6200) );
  nand_x2_sg U8229 ( .A(n6203), .B(n6204), .X(n6199) );
  nand_x1_sg U8230 ( .A(n8195), .B(n7660), .X(n6201) );
  nand_x2_sg U8231 ( .A(n6123), .B(n6124), .X(n6122) );
  nand_x2_sg U8232 ( .A(n6125), .B(n6126), .X(n6121) );
  nand_x1_sg U8233 ( .A(n8195), .B(n7676), .X(n6123) );
  nand_x2_sg U8234 ( .A(n6074), .B(n6075), .X(n6073) );
  nand_x2_sg U8235 ( .A(n6078), .B(n6079), .X(n6072) );
  nand_x1_sg U8236 ( .A(n8195), .B(n7684), .X(n6074) );
  nand_x2_sg U8237 ( .A(n5177), .B(n5260), .X(n5254) );
  nand_x1_sg U8238 ( .A(n5261), .B(n7340), .X(n5260) );
  nor_x1_sg U8239 ( .A(n6751), .B(n6752), .X(n6749) );
  nor_x1_sg U8240 ( .A(n6634), .B(n6635), .X(n6632) );
  nor_x1_sg U8241 ( .A(n6517), .B(n6518), .X(n6515) );
  nor_x1_sg U8242 ( .A(n6400), .B(n6401), .X(n6398) );
  nor_x1_sg U8243 ( .A(n6283), .B(n6284), .X(n6281) );
  nor_x1_sg U8244 ( .A(n6166), .B(n6167), .X(n6164) );
  nand_x2_sg U8245 ( .A(n6747), .B(n6748), .X(n6746) );
  nand_x2_sg U8246 ( .A(n6749), .B(n6750), .X(n6745) );
  nand_x1_sg U8247 ( .A(n8195), .B(n7702), .X(n6747) );
  nand_x2_sg U8248 ( .A(n6630), .B(n6631), .X(n6629) );
  nand_x2_sg U8249 ( .A(n6632), .B(n6633), .X(n6628) );
  nand_x1_sg U8250 ( .A(n8195), .B(n7726), .X(n6630) );
  nand_x2_sg U8251 ( .A(n6513), .B(n6514), .X(n6512) );
  nand_x2_sg U8252 ( .A(n6515), .B(n6516), .X(n6511) );
  nand_x1_sg U8253 ( .A(n8195), .B(n7750), .X(n6513) );
  nand_x2_sg U8254 ( .A(n6396), .B(n6397), .X(n6395) );
  nand_x2_sg U8255 ( .A(n6398), .B(n6399), .X(n6394) );
  nand_x1_sg U8256 ( .A(n6077), .B(n7774), .X(n6396) );
  nand_x2_sg U8257 ( .A(n6279), .B(n6280), .X(n6278) );
  nand_x2_sg U8258 ( .A(n6281), .B(n6282), .X(n6277) );
  nand_x1_sg U8259 ( .A(n8195), .B(n7644), .X(n6279) );
  nand_x2_sg U8260 ( .A(n6162), .B(n6163), .X(n6161) );
  nand_x2_sg U8261 ( .A(n6164), .B(n6165), .X(n6160) );
  nand_x1_sg U8262 ( .A(n8195), .B(n7668), .X(n6162) );
  nand_x4_sg U8263 ( .A(n6035), .B(n6036), .X(n5273) );
  nand_x1_sg U8264 ( .A(n7334), .B(n6037), .X(n6036) );
  nand_x1_sg U8265 ( .A(n4897), .B(n5077), .X(n6035) );
  nand_x1_sg U8266 ( .A(full), .B(n4881), .X(n5165) );
  nand_x2_sg U8267 ( .A(n5181), .B(n5182), .X(n5180) );
  nor_x1_sg U8268 ( .A(n5183), .B(n5184), .X(n5182) );
  nor_x1_sg U8269 ( .A(n5186), .B(n5187), .X(n5181) );
  nand_x4_sg U8270 ( .A(n5591), .B(n5592), .X(n5188) );
  nand_x1_sg U8271 ( .A(n7329), .B(n5586), .X(n5592) );
  nand_x1_sg U8272 ( .A(n4904), .B(n4911), .X(n5591) );
  nor_x1_sg U8273 ( .A(n6826), .B(n6827), .X(n6824) );
  nor_x1_sg U8274 ( .A(n6780), .B(n6781), .X(n6778) );
  nor_x1_sg U8275 ( .A(n6702), .B(n6703), .X(n6700) );
  nor_x1_sg U8276 ( .A(n6663), .B(n6664), .X(n6661) );
  nor_x1_sg U8277 ( .A(n6585), .B(n6586), .X(n6583) );
  nor_x1_sg U8278 ( .A(n6546), .B(n6547), .X(n6544) );
  nor_x1_sg U8279 ( .A(n6468), .B(n6469), .X(n6466) );
  nor_x1_sg U8280 ( .A(n6429), .B(n6430), .X(n6427) );
  nor_x1_sg U8281 ( .A(n6351), .B(n6352), .X(n6349) );
  nor_x1_sg U8282 ( .A(n6312), .B(n6313), .X(n6310) );
  nor_x1_sg U8283 ( .A(n6234), .B(n6235), .X(n6232) );
  nor_x1_sg U8284 ( .A(n6195), .B(n6196), .X(n6193) );
  nor_x1_sg U8285 ( .A(n6117), .B(n6118), .X(n6115) );
  nor_x1_sg U8286 ( .A(n6066), .B(n6067), .X(n6063) );
  nand_x2_sg U8287 ( .A(n6821), .B(n6822), .X(n6820) );
  nand_x2_sg U8288 ( .A(n6824), .B(n6825), .X(n6819) );
  nand_x1_sg U8289 ( .A(n8205), .B(n7692), .X(n6822) );
  nand_x2_sg U8290 ( .A(n6776), .B(n6777), .X(n6775) );
  nand_x2_sg U8291 ( .A(n6778), .B(n6779), .X(n6774) );
  nand_x1_sg U8292 ( .A(n8206), .B(n7700), .X(n6777) );
  nand_x2_sg U8293 ( .A(n6698), .B(n6699), .X(n6697) );
  nand_x2_sg U8294 ( .A(n6700), .B(n6701), .X(n6696) );
  nand_x1_sg U8295 ( .A(n8205), .B(n7716), .X(n6699) );
  nand_x2_sg U8296 ( .A(n6659), .B(n6660), .X(n6658) );
  nand_x2_sg U8297 ( .A(n6661), .B(n6662), .X(n6657) );
  nand_x1_sg U8298 ( .A(n8206), .B(n7724), .X(n6660) );
  nand_x2_sg U8299 ( .A(n6581), .B(n6582), .X(n6580) );
  nand_x2_sg U8300 ( .A(n6583), .B(n6584), .X(n6579) );
  nand_x1_sg U8301 ( .A(n8205), .B(n7740), .X(n6582) );
  nand_x2_sg U8302 ( .A(n6542), .B(n6543), .X(n6541) );
  nand_x2_sg U8303 ( .A(n6544), .B(n6545), .X(n6540) );
  nand_x1_sg U8304 ( .A(n8206), .B(n7748), .X(n6543) );
  nand_x2_sg U8305 ( .A(n6464), .B(n6465), .X(n6463) );
  nand_x2_sg U8306 ( .A(n6466), .B(n6467), .X(n6462) );
  nand_x1_sg U8307 ( .A(n8205), .B(n7764), .X(n6465) );
  nand_x2_sg U8308 ( .A(n6425), .B(n6426), .X(n6424) );
  nand_x2_sg U8309 ( .A(n6427), .B(n6428), .X(n6423) );
  nand_x1_sg U8310 ( .A(n8206), .B(n7772), .X(n6426) );
  nand_x2_sg U8311 ( .A(n6347), .B(n6348), .X(n6346) );
  nand_x2_sg U8312 ( .A(n6349), .B(n6350), .X(n6345) );
  nand_x1_sg U8313 ( .A(n8205), .B(n7626), .X(n6348) );
  nand_x2_sg U8314 ( .A(n6308), .B(n6309), .X(n6307) );
  nand_x2_sg U8315 ( .A(n6310), .B(n6311), .X(n6306) );
  nand_x1_sg U8316 ( .A(n8206), .B(n7634), .X(n6309) );
  nand_x2_sg U8317 ( .A(n6230), .B(n6231), .X(n6229) );
  nand_x2_sg U8318 ( .A(n6232), .B(n6233), .X(n6228) );
  nand_x1_sg U8319 ( .A(n8205), .B(n7650), .X(n6231) );
  nand_x2_sg U8320 ( .A(n6191), .B(n6192), .X(n6190) );
  nand_x2_sg U8321 ( .A(n6193), .B(n6194), .X(n6189) );
  nand_x1_sg U8322 ( .A(n8206), .B(n7658), .X(n6192) );
  nand_x2_sg U8323 ( .A(n6113), .B(n6114), .X(n6112) );
  nand_x2_sg U8324 ( .A(n6115), .B(n6116), .X(n6111) );
  nand_x1_sg U8325 ( .A(n8205), .B(n7674), .X(n6114) );
  nand_x2_sg U8326 ( .A(n6059), .B(n6060), .X(n6058) );
  nand_x2_sg U8327 ( .A(n6063), .B(n6064), .X(n6057) );
  nand_x1_sg U8328 ( .A(n8206), .B(n7682), .X(n6060) );
  nor_x1_sg U8329 ( .A(n6741), .B(n6742), .X(n6739) );
  nor_x1_sg U8330 ( .A(n6624), .B(n6625), .X(n6622) );
  nor_x1_sg U8331 ( .A(n6507), .B(n6508), .X(n6505) );
  nor_x1_sg U8332 ( .A(n6390), .B(n6391), .X(n6388) );
  nor_x1_sg U8333 ( .A(n6273), .B(n6274), .X(n6271) );
  nor_x1_sg U8334 ( .A(n6156), .B(n6157), .X(n6154) );
  nand_x2_sg U8335 ( .A(n6737), .B(n6738), .X(n6736) );
  nand_x2_sg U8336 ( .A(n6739), .B(n6740), .X(n6735) );
  nand_x1_sg U8337 ( .A(n6061), .B(n7708), .X(n6738) );
  nand_x2_sg U8338 ( .A(n6620), .B(n6621), .X(n6619) );
  nand_x2_sg U8339 ( .A(n6622), .B(n6623), .X(n6618) );
  nand_x1_sg U8340 ( .A(n6061), .B(n7732), .X(n6621) );
  nand_x2_sg U8341 ( .A(n6503), .B(n6504), .X(n6502) );
  nand_x2_sg U8342 ( .A(n6505), .B(n6506), .X(n6501) );
  nand_x1_sg U8343 ( .A(n6061), .B(n7756), .X(n6504) );
  nand_x2_sg U8344 ( .A(n6386), .B(n6387), .X(n6385) );
  nand_x2_sg U8345 ( .A(n6388), .B(n6389), .X(n6384) );
  nand_x1_sg U8346 ( .A(n6061), .B(n7780), .X(n6387) );
  nand_x2_sg U8347 ( .A(n6269), .B(n6270), .X(n6268) );
  nand_x2_sg U8348 ( .A(n6271), .B(n6272), .X(n6267) );
  nand_x1_sg U8349 ( .A(n6061), .B(n7642), .X(n6270) );
  nand_x2_sg U8350 ( .A(n6152), .B(n6153), .X(n6151) );
  nand_x2_sg U8351 ( .A(n6154), .B(n6155), .X(n6150) );
  nand_x1_sg U8352 ( .A(n6061), .B(n7666), .X(n6153) );
  nand_x1_sg U8353 ( .A(n5167), .B(n7333), .X(n6029) );
  nand_x1_sg U8354 ( .A(n4888), .B(n4893), .X(n6030) );
  nand_x1_sg U8355 ( .A(n5167), .B(n7340), .X(n6021) );
  nand_x1_sg U8356 ( .A(n4888), .B(n5270), .X(n6022) );
  nand_x1_sg U8357 ( .A(n8014), .B(n8255), .X(n5143) );
  nand_x1_sg U8358 ( .A(n8010), .B(n8256), .X(n5135) );
  nand_x1_sg U8359 ( .A(n8002), .B(n8256), .X(n5147) );
  nand_x1_sg U8360 ( .A(n7994), .B(n8255), .X(n5137) );
  nand_x1_sg U8361 ( .A(n7986), .B(n8255), .X(n5155) );
  nand_x1_sg U8362 ( .A(n7982), .B(n8256), .X(n5141) );
  nand_x1_sg U8363 ( .A(n7974), .B(n8255), .X(n5161) );
  nand_x1_sg U8364 ( .A(n7970), .B(n8255), .X(n5131) );
  nand_x1_sg U8365 ( .A(n7966), .B(n8256), .X(n5122) );
  nand_x1_sg U8366 ( .A(n7962), .B(n8255), .X(n5149) );
  nand_x1_sg U8367 ( .A(n7958), .B(n8256), .X(n5153) );
  nand_x1_sg U8368 ( .A(n7954), .B(n8256), .X(n5159) );
  nand_x1_sg U8369 ( .A(n7950), .B(n8256), .X(n5129) );
  nand_x1_sg U8370 ( .A(n7946), .B(n8255), .X(n5125) );
  nand_x1_sg U8371 ( .A(n7614), .B(n8229), .X(n5277) );
  nand_x1_sg U8372 ( .A(n7600), .B(n8229), .X(n5780) );
  nand_x1_sg U8373 ( .A(n7586), .B(n8230), .X(n5808) );
  nand_x1_sg U8374 ( .A(n7572), .B(n8230), .X(n5790) );
  nand_x1_sg U8375 ( .A(n7558), .B(n8230), .X(n5784) );
  nand_x1_sg U8376 ( .A(n7516), .B(n8229), .X(n5810) );
  nand_x1_sg U8377 ( .A(n7502), .B(n8230), .X(n5778) );
  nand_x1_sg U8378 ( .A(n7488), .B(n8229), .X(n5786) );
  nand_x1_sg U8379 ( .A(n7474), .B(n8230), .X(n5802) );
  nand_x1_sg U8380 ( .A(n7460), .B(n8230), .X(n5201) );
  nand_x1_sg U8381 ( .A(n7446), .B(n8229), .X(n5792) );
  nand_x1_sg U8382 ( .A(n7418), .B(n8230), .X(n5796) );
  nand_x1_sg U8383 ( .A(n7404), .B(n8229), .X(n5804) );
  nand_x1_sg U8384 ( .A(n7362), .B(n8229), .X(n5798) );
  nand_x1_sg U8385 ( .A(n8018), .B(n5124), .X(n5145) );
  nand_x1_sg U8386 ( .A(n8006), .B(n5124), .X(n5127) );
  nand_x1_sg U8387 ( .A(n7998), .B(n5124), .X(n5157) );
  nand_x1_sg U8388 ( .A(n7990), .B(n5124), .X(n5133) );
  nand_x1_sg U8389 ( .A(n7978), .B(n5124), .X(n5151) );
  nand_x1_sg U8390 ( .A(n7942), .B(n5124), .X(n5139) );
  nand_x1_sg U8391 ( .A(n7544), .B(n5203), .X(n5788) );
  nand_x1_sg U8392 ( .A(n7530), .B(n5203), .X(n5806) );
  nand_x1_sg U8393 ( .A(n7432), .B(n5203), .X(n5782) );
  nand_x1_sg U8394 ( .A(n7390), .B(n5203), .X(n5800) );
  nand_x1_sg U8395 ( .A(n7376), .B(n5203), .X(n5776) );
  nand_x1_sg U8396 ( .A(n7348), .B(n5203), .X(n5794) );
  nand_x1_sg U8397 ( .A(n7612), .B(n8231), .X(n5287) );
  nand_x1_sg U8398 ( .A(n7598), .B(n8232), .X(n5766) );
  nand_x1_sg U8399 ( .A(n7570), .B(n8231), .X(n5744) );
  nand_x1_sg U8400 ( .A(n7556), .B(n8231), .X(n5762) );
  nand_x1_sg U8401 ( .A(n7542), .B(n8232), .X(n5772) );
  nand_x1_sg U8402 ( .A(n7528), .B(n8232), .X(n5754) );
  nand_x1_sg U8403 ( .A(n7514), .B(n8231), .X(n5750) );
  nand_x1_sg U8404 ( .A(n7472), .B(n8232), .X(n5760) );
  nand_x1_sg U8405 ( .A(n7458), .B(n8232), .X(n5210) );
  nand_x1_sg U8406 ( .A(n7444), .B(n8232), .X(n5748) );
  nand_x1_sg U8407 ( .A(n7402), .B(n8231), .X(n5768) );
  nand_x1_sg U8408 ( .A(n7388), .B(n8231), .X(n5774) );
  nand_x1_sg U8409 ( .A(n7360), .B(n8232), .X(n5742) );
  nand_x1_sg U8410 ( .A(n7346), .B(n8231), .X(n5756) );
  nand_x1_sg U8411 ( .A(n7616), .B(n8227), .X(n5283) );
  nand_x1_sg U8412 ( .A(n7602), .B(n8228), .X(n5838) );
  nand_x1_sg U8413 ( .A(n7574), .B(n8227), .X(n5816) );
  nand_x1_sg U8414 ( .A(n7560), .B(n8228), .X(n5832) );
  nand_x1_sg U8415 ( .A(n7546), .B(n8228), .X(n5844) );
  nand_x1_sg U8416 ( .A(n7532), .B(n8228), .X(n5826) );
  nand_x1_sg U8417 ( .A(n7518), .B(n8227), .X(n5822) );
  nand_x1_sg U8418 ( .A(n7490), .B(n8227), .X(n5828) );
  nand_x1_sg U8419 ( .A(n7462), .B(n8228), .X(n5228) );
  nand_x1_sg U8420 ( .A(n7448), .B(n8228), .X(n5820) );
  nand_x1_sg U8421 ( .A(n7420), .B(n8227), .X(n5834) );
  nand_x1_sg U8422 ( .A(n7392), .B(n8227), .X(n5846) );
  nand_x1_sg U8423 ( .A(n7364), .B(n8228), .X(n5814) );
  nand_x1_sg U8424 ( .A(n7350), .B(n8227), .X(n5840) );
  nand_x1_sg U8425 ( .A(n7584), .B(n5212), .X(n5752) );
  nand_x1_sg U8426 ( .A(n7500), .B(n5212), .X(n5740) );
  nand_x1_sg U8427 ( .A(n7486), .B(n5212), .X(n5764) );
  nand_x1_sg U8428 ( .A(n7430), .B(n5212), .X(n5770) );
  nand_x1_sg U8429 ( .A(n7416), .B(n5212), .X(n5758) );
  nand_x1_sg U8430 ( .A(n7374), .B(n5212), .X(n5746) );
  nand_x1_sg U8431 ( .A(n7588), .B(n5230), .X(n5824) );
  nand_x1_sg U8432 ( .A(n7504), .B(n5230), .X(n5842) );
  nand_x1_sg U8433 ( .A(n7476), .B(n5230), .X(n5836) );
  nand_x1_sg U8434 ( .A(n7434), .B(n5230), .X(n5812) );
  nand_x1_sg U8435 ( .A(n7406), .B(n5230), .X(n5830) );
  nand_x1_sg U8436 ( .A(n7378), .B(n5230), .X(n5818) );
  nand_x2_sg U8437 ( .A(n5189), .B(n5190), .X(n5179) );
  nand_x1_sg U8438 ( .A(n7334), .B(n5191), .X(n5190) );
  nand_x1_sg U8439 ( .A(n4906), .B(n5077), .X(n5189) );
  nand_x2_sg U8440 ( .A(n5177), .B(n5178), .X(n5171) );
  nand_x1_sg U8441 ( .A(n4904), .B(n7329), .X(n5178) );
  nand_x1_sg U8442 ( .A(n4888), .B(n5273), .X(n6033) );
  nand_x1_sg U8443 ( .A(n5167), .B(n7334), .X(n6034) );
  nand_x1_sg U8444 ( .A(n4888), .B(n5259), .X(n6026) );
  nand_x1_sg U8445 ( .A(n5167), .B(n7300), .X(n6025) );
  nand_x1_sg U8446 ( .A(n4888), .B(n4900), .X(n6027) );
  nand_x1_sg U8447 ( .A(n5167), .B(n7284), .X(n6028) );
  nand_x1_sg U8448 ( .A(n8203), .B(n7292), .X(n6821) );
  nand_x1_sg U8449 ( .A(n8204), .B(n7312), .X(n6776) );
  nand_x1_sg U8450 ( .A(n8203), .B(n7294), .X(n6698) );
  nand_x1_sg U8451 ( .A(n8204), .B(n7316), .X(n6659) );
  nand_x1_sg U8452 ( .A(n8203), .B(n7296), .X(n6581) );
  nand_x1_sg U8453 ( .A(n8204), .B(n7320), .X(n6542) );
  nand_x1_sg U8454 ( .A(n8203), .B(n7298), .X(n6464) );
  nand_x1_sg U8455 ( .A(n8204), .B(n7324), .X(n6425) );
  nand_x1_sg U8456 ( .A(n8203), .B(n7286), .X(n6347) );
  nand_x1_sg U8457 ( .A(n8204), .B(n7302), .X(n6308) );
  nand_x1_sg U8458 ( .A(n8203), .B(n7288), .X(n6230) );
  nand_x1_sg U8459 ( .A(n8204), .B(n7306), .X(n6191) );
  nand_x1_sg U8460 ( .A(n8203), .B(n7290), .X(n6113) );
  nand_x1_sg U8461 ( .A(n8204), .B(n7310), .X(n6059) );
  nand_x1_sg U8462 ( .A(n6062), .B(n7314), .X(n6737) );
  nand_x1_sg U8463 ( .A(n6062), .B(n7318), .X(n6620) );
  nand_x1_sg U8464 ( .A(n6062), .B(n7322), .X(n6503) );
  nand_x1_sg U8465 ( .A(n6062), .B(n7326), .X(n6386) );
  nand_x1_sg U8466 ( .A(n6062), .B(n7304), .X(n6269) );
  nand_x1_sg U8467 ( .A(n6062), .B(n7308), .X(n6152) );
  nand_x1_sg U8468 ( .A(n5250), .B(n7329), .X(n5590) );
  nand_x1_sg U8469 ( .A(n5250), .B(n8106), .X(n5584) );
  nand_x1_sg U8470 ( .A(n4905), .B(n8259), .X(n5585) );
  nand_x2_sg U8471 ( .A(n5173), .B(n8259), .X(n5172) );
  nor_x1_sg U8472 ( .A(n5174), .B(n5175), .X(n5173) );
  nand_x2_sg U8473 ( .A(data_in[11]), .B(n8261), .X(n5313) );
  nand_x2_sg U8474 ( .A(data_in[0]), .B(n8259), .X(n5245) );
  nand_x2_sg U8475 ( .A(data_in[10]), .B(n8259), .X(n5969) );
  nand_x2_sg U8476 ( .A(data_in[8]), .B(n8259), .X(n5972) );
  nand_x2_sg U8477 ( .A(data_in[7]), .B(n8259), .X(n5999) );
  nand_x2_sg U8478 ( .A(data_in[6]), .B(n8259), .X(n5987) );
  nand_x2_sg U8479 ( .A(data_in[5]), .B(n8259), .X(n6008) );
  nand_x2_sg U8480 ( .A(data_in[3]), .B(n8259), .X(n5966) );
  nand_x2_sg U8481 ( .A(data_in[2]), .B(n8259), .X(n5984) );
  nand_x2_sg U8482 ( .A(data_in[1]), .B(n8259), .X(n6002) );
  nand_x2_sg U8483 ( .A(data_in[19]), .B(n8259), .X(n5975) );
  nand_x2_sg U8484 ( .A(data_in[18]), .B(n8259), .X(n5990) );
  nand_x2_sg U8485 ( .A(data_in[17]), .B(n8259), .X(n5993) );
  nand_x2_sg U8486 ( .A(data_in[16]), .B(n8259), .X(n6005) );
  nand_x2_sg U8487 ( .A(data_in[15]), .B(n8259), .X(n5981) );
  nand_x2_sg U8488 ( .A(data_in[14]), .B(n8259), .X(n5963) );
  nand_x2_sg U8489 ( .A(data_in[13]), .B(n8259), .X(n5996) );
  nand_x2_sg U8490 ( .A(data_in[12]), .B(n8259), .X(n5978) );
  nand_x1_sg U8491 ( .A(n4906), .B(n8259), .X(n5582) );
  nand_x1_sg U8492 ( .A(n5250), .B(n7338), .X(n5581) );
  nand_x1_sg U8493 ( .A(n8259), .B(n4902), .X(n5575) );
  nand_x1_sg U8494 ( .A(n5250), .B(n7331), .X(n5576) );
  nand_x1_sg U8495 ( .A(n4901), .B(n8259), .X(n5578) );
  nand_x1_sg U8496 ( .A(n5250), .B(n7282), .X(n5577) );
  nand_x2_sg U8497 ( .A(data_in[9]), .B(n8259), .X(n6011) );
  nand_x2_sg U8498 ( .A(data_in[4]), .B(n8259), .X(n6014) );
  nand_x1_sg U8499 ( .A(n7284), .B(n4902), .X(n5262) );
  nand_x1_sg U8500 ( .A(n7331), .B(n4900), .X(n5263) );
  inv_x8_sg U8501 ( .A(reset), .X(n4887) );
  inv_x8_sg U8502 ( .A(n8256), .X(n8107) );
  inv_x8_sg U8503 ( .A(n8232), .X(n8108) );
  inv_x8_sg U8504 ( .A(n8230), .X(n8109) );
  inv_x8_sg U8505 ( .A(n8228), .X(n8110) );
  inv_x8_sg U8506 ( .A(n8111), .X(n8112) );
  inv_x8_sg U8507 ( .A(n8113), .X(n8114) );
  inv_x8_sg U8508 ( .A(n8115), .X(n8116) );
  inv_x8_sg U8509 ( .A(n8117), .X(n8118) );
  inv_x8_sg U8510 ( .A(n8119), .X(n8120) );
  inv_x8_sg U8511 ( .A(n8121), .X(n8122) );
  inv_x8_sg U8512 ( .A(n8123), .X(n8124) );
  inv_x8_sg U8513 ( .A(n8125), .X(n8126) );
  inv_x8_sg U8514 ( .A(n8127), .X(n8128) );
  inv_x8_sg U8515 ( .A(n8129), .X(n8130) );
  inv_x8_sg U8516 ( .A(n8131), .X(n8132) );
  inv_x8_sg U8517 ( .A(n8133), .X(n8134) );
  inv_x8_sg U8518 ( .A(n8135), .X(n8136) );
  inv_x8_sg U8519 ( .A(n8137), .X(n8138) );
  inv_x8_sg U8520 ( .A(n8139), .X(n8140) );
  inv_x8_sg U8521 ( .A(n8141), .X(n8142) );
  inv_x8_sg U8522 ( .A(n8143), .X(n8144) );
  inv_x8_sg U8523 ( .A(n8145), .X(n8146) );
  inv_x8_sg U8524 ( .A(n8147), .X(n8148) );
  inv_x8_sg U8525 ( .A(n8149), .X(n8150) );
  inv_x8_sg U8526 ( .A(n8254), .X(n8151) );
  inv_x8_sg U8527 ( .A(n8252), .X(n8152) );
  inv_x8_sg U8528 ( .A(n8250), .X(n8153) );
  inv_x8_sg U8529 ( .A(n8248), .X(n8154) );
  inv_x8_sg U8530 ( .A(n8257), .X(n8155) );
  inv_x8_sg U8531 ( .A(n8245), .X(n8156) );
  inv_x8_sg U8532 ( .A(n8244), .X(n8157) );
  inv_x8_sg U8533 ( .A(n8242), .X(n8158) );
  inv_x8_sg U8534 ( .A(n8240), .X(n8159) );
  inv_x8_sg U8535 ( .A(n8237), .X(n8160) );
  inv_x8_sg U8536 ( .A(n8236), .X(n8161) );
  inv_x8_sg U8537 ( .A(n8234), .X(n8162) );
  inv_x8_sg U8538 ( .A(n8226), .X(n8163) );
  inv_x8_sg U8539 ( .A(n8224), .X(n8164) );
  inv_x8_sg U8540 ( .A(n8222), .X(n8165) );
  inv_x8_sg U8541 ( .A(n8220), .X(n8166) );
  nand_x8_sg U8542 ( .A(n4898), .B(n6839), .X(n8167) );
  nand_x8_sg U8543 ( .A(n4898), .B(n6839), .X(n8168) );
  nand_x8_sg U8544 ( .A(n4899), .B(n6839), .X(n8169) );
  inv_x4_sg U8545 ( .A(n8173), .X(n8170) );
  inv_x4_sg U8546 ( .A(n8173), .X(n8171) );
  inv_x4_sg U8547 ( .A(n8173), .X(n8172) );
  inv_x8_sg U8548 ( .A(n6093), .X(n8173) );
  inv_x8_sg U8549 ( .A(n8178), .X(n8179) );
  inv_x4_sg U8550 ( .A(n8179), .X(n8180) );
  inv_x4_sg U8551 ( .A(n8179), .X(n8181) );
  inv_x4_sg U8552 ( .A(n8179), .X(n8182) );
  inv_x8_sg U8553 ( .A(n8187), .X(n8188) );
  nand_x8_sg U8554 ( .A(n4891), .B(n6839), .X(n8189) );
  nand_x8_sg U8555 ( .A(n4891), .B(n6839), .X(n8190) );
  nand_x8_sg U8556 ( .A(n4898), .B(n6828), .X(n8191) );
  inv_x8_sg U8557 ( .A(n8192), .X(n8193) );
  inv_x8_sg U8558 ( .A(n8194), .X(n8195) );
  nor_x4_sg U8559 ( .A(n6823), .B(n6810), .X(n6077) );
  inv_x8_sg U8560 ( .A(n8196), .X(n8197) );
  nand_x8_sg U8561 ( .A(n4899), .B(n6828), .X(n8198) );
  nand_x8_sg U8562 ( .A(n4899), .B(n6828), .X(n8199) );
  nand_x8_sg U8563 ( .A(n6828), .B(n4891), .X(n8200) );
  nand_x8_sg U8564 ( .A(n6828), .B(n4891), .X(n8201) );
  nor_x8_sg U8565 ( .A(n6823), .B(n6037), .X(n8202) );
  nor_x8_sg U8566 ( .A(n6823), .B(n6037), .X(n6065) );
  nor_x8_sg U8567 ( .A(n6823), .B(n6811), .X(n8205) );
  nor_x8_sg U8568 ( .A(n6823), .B(n6811), .X(n8206) );
  nor_x8_sg U8569 ( .A(n6823), .B(n6811), .X(n6061) );
  nand_x8_sg U8570 ( .A(n4899), .B(n7340), .X(n8207) );
  nand_x8_sg U8571 ( .A(n4899), .B(n7340), .X(n8208) );
  nand_x8_sg U8572 ( .A(n6815), .B(n4897), .X(n8209) );
  nand_x8_sg U8573 ( .A(n6815), .B(n4897), .X(n8210) );
  inv_x8_sg U8574 ( .A(n8211), .X(n8212) );
  inv_x8_sg U8575 ( .A(n8213), .X(n8214) );
  inv_x8_sg U8576 ( .A(n8215), .X(n8216) );
  nand_x8_sg U8577 ( .A(n6801), .B(rd_en), .X(n8217) );
  nand_x8_sg U8578 ( .A(n6801), .B(rd_en), .X(n8218) );
  nand_x8_sg U8579 ( .A(n5424), .B(n5887), .X(n8219) );
  nand_x8_sg U8580 ( .A(n5424), .B(n5887), .X(n8220) );
  nand_x8_sg U8581 ( .A(n5350), .B(n5887), .X(n8221) );
  nand_x8_sg U8582 ( .A(n5350), .B(n5887), .X(n8222) );
  nand_x8_sg U8583 ( .A(n5461), .B(n5887), .X(n8223) );
  nand_x8_sg U8584 ( .A(n5461), .B(n5887), .X(n8224) );
  nand_x8_sg U8585 ( .A(n5120), .B(n5887), .X(n8225) );
  nand_x8_sg U8586 ( .A(n5120), .B(n5887), .X(n8226) );
  nand_x8_sg U8587 ( .A(n5424), .B(n5163), .X(n8227) );
  nand_x8_sg U8588 ( .A(n5424), .B(n5163), .X(n8228) );
  nand_x8_sg U8589 ( .A(n5461), .B(n5163), .X(n8229) );
  nand_x8_sg U8590 ( .A(n5461), .B(n5163), .X(n8230) );
  nand_x8_sg U8591 ( .A(n5350), .B(n5163), .X(n8231) );
  nand_x8_sg U8592 ( .A(n5350), .B(n5163), .X(n8232) );
  nand_x8_sg U8593 ( .A(n5350), .B(n5629), .X(n8233) );
  nand_x8_sg U8594 ( .A(n5350), .B(n5629), .X(n8234) );
  nand_x8_sg U8595 ( .A(n5424), .B(n5629), .X(n8235) );
  nand_x8_sg U8596 ( .A(n5424), .B(n5629), .X(n8236) );
  nand_x8_sg U8597 ( .A(n5461), .B(n5629), .X(n8237) );
  nand_x8_sg U8598 ( .A(n5461), .B(n5629), .X(n8238) );
  nand_x8_sg U8599 ( .A(n5120), .B(n5629), .X(n8239) );
  nand_x8_sg U8600 ( .A(n5120), .B(n5629), .X(n8240) );
  nand_x8_sg U8601 ( .A(n5350), .B(n5121), .X(n8241) );
  nand_x8_sg U8602 ( .A(n5350), .B(n5121), .X(n8242) );
  nand_x8_sg U8603 ( .A(n5461), .B(n5121), .X(n8243) );
  nand_x8_sg U8604 ( .A(n5461), .B(n5121), .X(n8244) );
  nand_x8_sg U8605 ( .A(n5424), .B(n5121), .X(n8245) );
  nand_x8_sg U8606 ( .A(n5424), .B(n5121), .X(n8246) );
  nand_x8_sg U8607 ( .A(n5461), .B(n5351), .X(n8247) );
  nand_x8_sg U8608 ( .A(n5461), .B(n5351), .X(n8248) );
  nand_x8_sg U8609 ( .A(n5424), .B(n5351), .X(n8249) );
  nand_x8_sg U8610 ( .A(n5424), .B(n5351), .X(n8250) );
  nand_x8_sg U8611 ( .A(n5120), .B(n5351), .X(n8251) );
  nand_x8_sg U8612 ( .A(n5120), .B(n5351), .X(n8252) );
  nand_x8_sg U8613 ( .A(n5350), .B(n5351), .X(n8253) );
  nand_x8_sg U8614 ( .A(n5350), .B(n5351), .X(n8254) );
  nand_x8_sg U8615 ( .A(n5120), .B(n5163), .X(n8255) );
  nand_x8_sg U8616 ( .A(n5120), .B(n5163), .X(n8256) );
  nand_x8_sg U8617 ( .A(n5120), .B(n5121), .X(n8257) );
  nand_x8_sg U8618 ( .A(n5120), .B(n5121), .X(n8258) );
  inv_x8_sg U8619 ( .A(n8260), .X(n8259) );
endmodule

