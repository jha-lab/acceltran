
module pooling ( clk, reset, .im({\im[3][19] , \im[3][18] , \im[3][17] , 
        \im[3][16] , \im[3][15] , \im[3][14] , \im[3][13] , \im[3][12] , 
        \im[3][11] , \im[3][10] , \im[3][9] , \im[3][8] , \im[3][7] , 
        \im[3][6] , \im[3][5] , \im[3][4] , \im[3][3] , \im[3][2] , \im[3][1] , 
        \im[3][0] , \im[2][19] , \im[2][18] , \im[2][17] , \im[2][16] , 
        \im[2][15] , \im[2][14] , \im[2][13] , \im[2][12] , \im[2][11] , 
        \im[2][10] , \im[2][9] , \im[2][8] , \im[2][7] , \im[2][6] , 
        \im[2][5] , \im[2][4] , \im[2][3] , \im[2][2] , \im[2][1] , \im[2][0] , 
        \im[1][19] , \im[1][18] , \im[1][17] , \im[1][16] , \im[1][15] , 
        \im[1][14] , \im[1][13] , \im[1][12] , \im[1][11] , \im[1][10] , 
        \im[1][9] , \im[1][8] , \im[1][7] , \im[1][6] , \im[1][5] , \im[1][4] , 
        \im[1][3] , \im[1][2] , \im[1][1] , \im[1][0] , \im[0][19] , 
        \im[0][18] , \im[0][17] , \im[0][16] , \im[0][15] , \im[0][14] , 
        \im[0][13] , \im[0][12] , \im[0][11] , \im[0][10] , \im[0][9] , 
        \im[0][8] , \im[0][7] , \im[0][6] , \im[0][5] , \im[0][4] , \im[0][3] , 
        \im[0][2] , \im[0][1] , \im[0][0] }), input_ready, output_taken, mode, 
        om, state );
  input [1:0] mode;
  output [19:0] om;
  output [1:0] state;
  input clk, reset, \im[3][19] , \im[3][18] , \im[3][17] , \im[3][16] ,
         \im[3][15] , \im[3][14] , \im[3][13] , \im[3][12] , \im[3][11] ,
         \im[3][10] , \im[3][9] , \im[3][8] , \im[3][7] , \im[3][6] ,
         \im[3][5] , \im[3][4] , \im[3][3] , \im[3][2] , \im[3][1] ,
         \im[3][0] , \im[2][19] , \im[2][18] , \im[2][17] , \im[2][16] ,
         \im[2][15] , \im[2][14] , \im[2][13] , \im[2][12] , \im[2][11] ,
         \im[2][10] , \im[2][9] , \im[2][8] , \im[2][7] , \im[2][6] ,
         \im[2][5] , \im[2][4] , \im[2][3] , \im[2][2] , \im[2][1] ,
         \im[2][0] , \im[1][19] , \im[1][18] , \im[1][17] , \im[1][16] ,
         \im[1][15] , \im[1][14] , \im[1][13] , \im[1][12] , \im[1][11] ,
         \im[1][10] , \im[1][9] , \im[1][8] , \im[1][7] , \im[1][6] ,
         \im[1][5] , \im[1][4] , \im[1][3] , \im[1][2] , \im[1][1] ,
         \im[1][0] , \im[0][19] , \im[0][18] , \im[0][17] , \im[0][16] ,
         \im[0][15] , \im[0][14] , \im[0][13] , \im[0][12] , \im[0][11] ,
         \im[0][10] , \im[0][9] , \im[0][8] , \im[0][7] , \im[0][6] ,
         \im[0][5] , \im[0][4] , \im[0][3] , \im[0][2] , \im[0][1] ,
         \im[0][0] , input_ready, output_taken;
  wire   \reg_im[3][19] , \reg_im[3][18] , \reg_im[3][17] , \reg_im[3][16] ,
         \reg_im[3][15] , \reg_im[3][14] , \reg_im[3][13] , \reg_im[3][12] ,
         \reg_im[3][11] , \reg_im[3][10] , \reg_im[3][9] , \reg_im[3][8] ,
         \reg_im[3][7] , \reg_im[3][6] , \reg_im[3][5] , \reg_im[3][4] ,
         \reg_im[3][3] , \reg_im[3][2] , \reg_im[3][1] , \reg_im[3][0] ,
         \reg_im[2][19] , \reg_im[2][18] , \reg_im[2][17] , \reg_im[2][16] ,
         \reg_im[2][15] , \reg_im[2][14] , \reg_im[2][13] , \reg_im[2][12] ,
         \reg_im[2][11] , \reg_im[2][10] , \reg_im[2][9] , \reg_im[2][8] ,
         \reg_im[2][7] , \reg_im[2][6] , \reg_im[2][5] , \reg_im[2][4] ,
         \reg_im[2][3] , \reg_im[2][2] , \reg_im[2][1] , \reg_im[2][0] ,
         \reg_im[1][19] , \reg_im[1][18] , \reg_im[1][17] , \reg_im[1][16] ,
         \reg_im[1][15] , \reg_im[1][14] , \reg_im[1][13] , \reg_im[1][12] ,
         \reg_im[1][11] , \reg_im[1][10] , \reg_im[1][9] , \reg_im[1][8] ,
         \reg_im[1][7] , \reg_im[1][6] , \reg_im[1][5] , \reg_im[1][4] ,
         \reg_im[1][3] , \reg_im[1][2] , \reg_im[1][1] , \reg_im[1][0] ,
         \reg_im[0][19] , \reg_im[0][18] , \reg_im[0][17] , \reg_im[0][16] ,
         \reg_im[0][15] , \reg_im[0][14] , \reg_im[0][13] , \reg_im[0][12] ,
         \reg_im[0][11] , \reg_im[0][10] , \reg_im[0][9] , \reg_im[0][8] ,
         \reg_im[0][7] , \reg_im[0][6] , \reg_im[0][5] , \reg_im[0][4] ,
         \reg_im[0][3] , \reg_im[0][2] , \reg_im[0][1] , \reg_im[0][0] , N112,
         reg_input_ready, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, \max_pooling_0/n352 ,
         \max_pooling_0/n351 , \max_pooling_0/n350 , \max_pooling_0/n349 ,
         \max_pooling_0/n348 , \max_pooling_0/n347 , \max_pooling_0/n346 ,
         \max_pooling_0/n345 , \max_pooling_0/n344 , \max_pooling_0/n343 ,
         \max_pooling_0/n342 , \max_pooling_0/n341 , \max_pooling_0/n340 ,
         \max_pooling_0/n339 , \max_pooling_0/n338 , \max_pooling_0/n337 ,
         \max_pooling_0/n336 , \max_pooling_0/n335 , \max_pooling_0/n334 ,
         \max_pooling_0/n333 , \max_pooling_0/n332 , \max_pooling_0/n331 ,
         \max_pooling_0/n330 , \max_pooling_0/n329 , \max_pooling_0/n328 ,
         \max_pooling_0/n327 , \max_pooling_0/n326 , \max_pooling_0/n325 ,
         \max_pooling_0/n324 , \max_pooling_0/n323 , \max_pooling_0/n322 ,
         \max_pooling_0/n321 , \max_pooling_0/n320 , \max_pooling_0/n319 ,
         \max_pooling_0/n318 , \max_pooling_0/n317 , \max_pooling_0/n316 ,
         \max_pooling_0/n315 , \max_pooling_0/n314 , \max_pooling_0/n313 ,
         \max_pooling_0/n312 , \max_pooling_0/n311 , \max_pooling_0/n643 ,
         \max_pooling_0/n642 , \max_pooling_0/n641 , \max_pooling_0/n640 ,
         \max_pooling_0/n639 , \max_pooling_0/N4 , \max_pooling_0/N3 ,
         \mean_pooling_0/n265 , \mean_pooling_0/n264 , \mean_pooling_0/n263 ,
         \mean_pooling_0/n262 , \mean_pooling_0/n261 , \mean_pooling_0/n260 ,
         \mean_pooling_0/n259 , \mean_pooling_0/n258 , \mean_pooling_0/n257 ,
         \mean_pooling_0/n256 , \mean_pooling_0/n255 , \mean_pooling_0/n254 ,
         \mean_pooling_0/n253 , \mean_pooling_0/n252 , \mean_pooling_0/n251 ,
         \mean_pooling_0/n250 , \mean_pooling_0/n249 , \mean_pooling_0/n248 ,
         \mean_pooling_0/n247 , \mean_pooling_0/n246 , \mean_pooling_0/N5 ,
         \mean_pooling_0/N4 , \min_pooling_0/n413 , \min_pooling_0/n412 ,
         \min_pooling_0/n411 , \min_pooling_0/n410 , \min_pooling_0/n409 ,
         \min_pooling_0/n408 , \min_pooling_0/n407 , \min_pooling_0/n406 ,
         \min_pooling_0/n405 , \min_pooling_0/n404 , \min_pooling_0/n403 ,
         \min_pooling_0/n402 , \min_pooling_0/n401 , \min_pooling_0/n400 ,
         \min_pooling_0/n399 , \min_pooling_0/n398 , \min_pooling_0/n397 ,
         \min_pooling_0/n396 , \min_pooling_0/n395 , \min_pooling_0/n394 ,
         \min_pooling_0/n393 , \min_pooling_0/n392 , \min_pooling_0/n265 ,
         \min_pooling_0/n264 , \min_pooling_0/n263 , \min_pooling_0/n262 ,
         \min_pooling_0/n261 , \min_pooling_0/n260 , \min_pooling_0/n259 ,
         \min_pooling_0/n258 , \min_pooling_0/n257 , \min_pooling_0/n256 ,
         \min_pooling_0/n255 , \min_pooling_0/n254 , \min_pooling_0/n253 ,
         \min_pooling_0/n252 , \min_pooling_0/n251 , \min_pooling_0/n250 ,
         \min_pooling_0/n249 , \min_pooling_0/n248 , \min_pooling_0/n247 ,
         \min_pooling_0/n246 , \min_pooling_0/n724 , \min_pooling_0/n723 ,
         \min_pooling_0/n722 , \min_pooling_0/N4 , \min_pooling_0/N3 , n2454,
         n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
         n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474,
         n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
         n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
         n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
         n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
         n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524,
         n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534,
         n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544,
         n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554,
         n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564,
         n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574,
         n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584,
         n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594,
         n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604,
         n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614,
         n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624,
         n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634,
         n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2643, n2644, n2645,
         n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655,
         n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665,
         n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675,
         n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685,
         n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695,
         n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705,
         n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715,
         n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725,
         n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735,
         n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745,
         n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755,
         n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765,
         n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775,
         n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785,
         n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795,
         n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805,
         n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815,
         n2816, n2817, n2818, n2819, n2820, n441, n437, n433, n429, n425, n422,
         n421, n418, n417, n414, n413, n410, n406, n405, n401, n397, n393,
         n389, n385, n381, n377, n373, n369, n365, n361, n357, n353, n349,
         n2179, n2178, n2177, n2176, n2175, n2174, n2173, n2172, n2171, n2170,
         n2169, n2168, n2167, n2166, n2165, n2164, n2163, n2162, n2161, n2160,
         n2159, n2158, n2157, n2156, n2155, n2154, n2153, n2152, n2151, n2150,
         n2149, n2148, n2147, n2146, n2145, n2144, n2143, n2142, n2141, n2140,
         n2139, n2138, n2137, n2136, n2135, n2134, n2133, n2132, n2131, n2130,
         n2129, n2128, n2127, n2126, n2125, n2124, n2123, n2122, n2121, n2120,
         n2119, n2118, n2117, n2116, n2115, n2114, n2113, n2112, n2111, n2110,
         n2109, n2108, n2107, n2106, n2105, n2104, n2103, n2102, n2101, n2100,
         n2099, n2098, n2097, n2096, n2095, n2094, n2093, n2092, n2091, n2090,
         n2089, n2088, n2087, n2086, n2085, n2084, n2083, n2082, n2081, n2080,
         n2079, n2078, n2077, n2076, n2075, n2074, n2073, n2072, n2071, n2070,
         n2069, n2068, n2067, n2066, n2065, n2064, n2063, n2062, n2061, n2060,
         n2059, n2058, n2057, n2056, n2055, n2054, n2053, n2052, n2051, n2050,
         n2049, n2048, n2047, n2046, n2045, n2044, n2043, n2042, n2041, n2040,
         n2039, n2038, n2037, n2036, n2035, n2034, n2033, n2032, n2031, n2030,
         n2029, n2028, n2027, n2026, n2025, n2024, n2023, n2022, n2021, n2020,
         n2019, n2018, n2017, n2016, n2015, n2014, n2013, n2012, n2011, n2010,
         n2009, n2008, n2007, n2006, n2005, n2004, n2003, n2002, n2001, n2000,
         n1999, n1998, n1997, n1996, n1995, n1994, n1993, n1992, n1991, n1989,
         n1988, n1987, n1986, n1985, n1984, n1983, n1982, n1981, n1980, n1979,
         n1978, n1977, n1976, n1975, n1974, n1973, n1972, n1971, n1970, n1969,
         n1968, n1967, n1966, n1965, n1964, n1963, n1962, n1961, n1960, n1959,
         n1958, n1957, n1956, n1955, n1954, n1953, n1952, n1951, n1950, n1949,
         n1948, n1947, n1946, n1945, n1944, n1943, n1942, n1941, n1940, n1939,
         n1938, n1937, n1936, n1935, n1934, n1933, n1932, n1931, n1930, n1929,
         n1928, n1927, n1926, n1925, n1924, n1923, n1922, n1921, n1920, n1919,
         n1918, n1917, n1916, n1915, n1914, n1913, n1912, n1911, n1910, n1909,
         n1908, n1907, n1906, n1905, n1904, n1903, n1902, n1901, n1900, n1899,
         n1898, n1897, n1896, n1895, n1894, n1893, n1892, n1891, n1890, n1889,
         n1888, n1887, n1886, n1885, n1884, n1883, n1882, n1881, n1880, n1879,
         n1878, n1877, n1876, n1875, n1874, n1873, n1872, n1870, n1869, n1868,
         n1867, n1866, n1865, n1864, n1863, n1862, n1861, n1860, n1859, n1858,
         n1857, n1856, n1855, n1854, n1853, n1852, n1851, n1850, n1849, n1848,
         n1847, n1846, n1845, n1844, n1843, n1842, n1841, n1840, n1839, n1838,
         n1837, n1836, n1835, n1834, n1833, n1832, n1831, n1830, n1829, n1828,
         n1827, n1826, n1825, n1824, n1823, n1822, n1821, n1820, n1819, n1818,
         n1817, n1816, n1815, n1814, n1813, n1812, n1811, n1810, n1809, n1808,
         n1807, n1806, n1805, n1804, n1803, n1802, n1801, n1800, n1799, n1798,
         n1797, n1796, n1795, n1794, n1793, n1792, n1791, n1790, n1789, n1788,
         n1787, n1786, n1785, n1784, n1783, n1782, n1781, n1780, n1779, n1778,
         n1777, n1776, n1775, n1774, n1773, n1772, n1771, n1770, n1769, n1768,
         n1767, n1766, n1765, n1764, n1763, n1762, n1761, n1760, n1759, n1758,
         n1757, n1756, n1755, n1754, n1753, n1752, n1751, n1750, n1749, n1748,
         n1747, n1746, n1745, n1744, n1743, n1742, n1741, n1740, n1739, n1738,
         n1737, n1736, n1735, n1734, n1733, n1732, n1731, n1730, n1729, n1728,
         n1727, n1726, n1725, n1724, n1723, n1722, n1721, n1720, n1719, n1718,
         n1717, n1716, n1715, n1714, n1713, n1712, n1711, n1710, n1709, n1708,
         n1707, n1706, n1705, n1704, n1703, n1702, n1701, n1700, n1699, n1698,
         n1697, n1696, n1695, n1694, n1693, n1692, n1691, n1690, n1689, n1688,
         n1687, n1686, n1685, n1684, n1683, n1682, n1681, n1680, n1679, n1678,
         n1677, n1676, n1675, n1674, n1673, n1672, n1671, n1670, n1669, n1668,
         n1667, n1666, n1665, n1664, n1663, n1662, n1661, n1660, n1659, n1658,
         n1657, n1656, n1655, n1654, n1653, n1652, n1651, n1650, n1649, n1648,
         n1647, n1646, n1645, n1644, n1643, n1642, n1641, n1640, n1639, n1638,
         n1637, n1636, n1635, n1634, n1633, n1632, n1631, n1630, n1629, n1628,
         n1627, n1626, n1625, n1624, n1623, n1622, n1621, n1620, n1619, n1618,
         n1617, n1616, n1615, n1614, n1613, n1612, n1611, n1610, n1609, n1608,
         n1607, n1606, n1605, n1604, n1603, n1602, n1601, n1600, n1599, n1598,
         n1597, n1596, n1595, n1594, n1593, n1592, n1591, n1590, n1589, n1588,
         n1587, n1586, n1585, n1584, n1583, n1582, n1581, n1580, n1579, n1578,
         n1577, n1576, n1575, n1574, n1573, n1572, n1571, n1570, n1569, n1568,
         n1567, n1566, n1565, n1564, n1563, n1562, n1561, n1560, n1559, n1558,
         n1557, n1556, n1555, n1554, n1553, n1552, n1551, n1550, n1549, n1548,
         n1547, n1546, n1545, n1544, n1543, n1542, n1541, n1540, n1539, n1538,
         n1537, n1536, n1535, n1534, n1533, n1532, n1531, n1530, n1529, n1528,
         n1527, n1526, n1525, n1524, n1523, n1522, n1521, n1520, n1519, n1518,
         n1517, n1516, n1515, n1514, n1513, n1512, n1511, n1510, n1509, n1508,
         n1507, n1506, n1505, n1504, n1503, n1502, n1501, n1500, n1499, n1498,
         n1497, n1496, n1495, n1494, n1493, n1492, n1491, n1490, n1489, n1488,
         n1487, n1486, n1485, n1484, n1483, n1482, n1481, n1480, n1479, n1478,
         n1477, n1476, n1475, n1474, n1473, n1472, n1471, n1470, n1469, n1468,
         n1467, n1466, n1465, n1464, n1463, n1462, n1461, n1460, n1459, n1458,
         n1457, n1456, n1455, n1454, n1453, n1452, n1451, n1450, n1449, n1448,
         n1447, n1446, n1445, n1444, n1443, n1442, n1441, n1440, n1439, n1438,
         n1437, n1436, n1435, n1434, n1433, n1432, n1431, n1430, n1429, n1428,
         n1427, n1426, n1425, n1424, n1423, n1422, n1421, n1420, n1419, n1418,
         n1417, n1416, n1415, n1414, n1413, n1412, n1411, n1410, n1409, n1408,
         n1407, n1406, n1405, n1404, n1403, n1402, n1401, n1400, n1399, n1398,
         n1397, n1396, n1395, n1394, n1393, n1392, n1391, n1390, n1389, n1388,
         n1387, n1386, n1385, n1384, n1383, n1382, n1381, n1380, n1379, n1378,
         n1377, n1376, n1375, n1374, n1373, n1372, n1371, n1370, n1369, n1368,
         n1367, n1366, n1365, n1364, n1363, n1362, n1361, n1360, n1359, n1358,
         n1357, n1356, n1355, n1354, n1353, n1352, n1351, n1350, n1349, n1348,
         n1347, n1346, n1345, n1344, n1343, n1342, n1341, n1340, n1339, n1338,
         n1337, n1336, n1335, n1334, n1333, n1332, n1331, n1330, n1329, n1328,
         n1326, n1325, n1324, n1323, n1322, n1321, n1320, n1319, n1318, n1317,
         n1316, n1315, n1314, n1313, n1312, n1311, n1310, n1309, n1308, n1307,
         n1306, n1305, n1304, n1303, n1302, n1301, n1300, n1299, n1298, n1297,
         n1296, n1295, n1294, n1293, n1292, n1291, n1290, n1289, n1288, n1287,
         n1286, n1285, n1284, n1283, n1282, n1281, n1280, n1279, n1278, n1277,
         n1276, n1275, n1274, n1273, n1272, n1271, n1270, n1269, n1268, n1267,
         n1266, n1265, n1264, n1263, n1262, n1261, n1260, n1259, n1258, n1257,
         n1256, n1255, n1254, n1253, n1252, n1251, n1250, n1249, n1248, n1247,
         n1246, n1245, n1244, n1243, n1242, n1241, n1240, n1239, n1238, n1237,
         n1236, n1235, n1234, n1233, n1232, n1231, n1230, n1229, n1228, n1227,
         n1226, n1225, n1224, n1223, n1222, n1221, n1220, n1219, n1218, n1217,
         n1216, n1215, n1214, n1213, n1212, n1211, n1210, n1209, n1208, n1207,
         n1206, n1205, n1204, n1203, n1202, n1201, n1200, n1199, n1198, n1197,
         n1196, n1195, n1194, n1193, n1192, n1191, n1190, n1189, n1188, n1187,
         n1186, n1185, n1184, n1183, n1182, n1181, n1180, n1179, n1178, n1177,
         n1176, n1175, n1174, n1173, n1172, n1171, n1170, n1169, n1168, n1167,
         n1166, n1165, n1164, n1163, n1162, n1161, n1160, n1159, n1158, n1157,
         n1156, n1155, n1154, n1153, n1152, n1151, n1150, n1149, n1148, n1147,
         n1146, n1145, n1144, n1143, n1142, n1141, n1140, n1139, n1138, n1137,
         n1136, n1135, n1134, n1133, n1132, n1131, n1130, n1129, n1128, n1127,
         n1126, n1125, n1124, n1123, n1122, n1121, n1120, n1119, n1118, n1117,
         n1116, n1115, n1113, n1112, n1111, n1110, n1109, n1108, n1107, n1106,
         n1105, n1104, n1103, n1102, n1101, n1100, n1099, n1098, n1097, n1096,
         n1095, n1094, n1093, \min_pooling_0/n390 , \min_pooling_0/n389 ,
         \min_pooling_0/n386 , \min_pooling_0/n385 , \min_pooling_0/n382 ,
         \min_pooling_0/n381 , \min_pooling_0/n378 , \min_pooling_0/n377 ,
         \min_pooling_0/n374 , \min_pooling_0/n373 , \min_pooling_0/n370 ,
         \min_pooling_0/n369 , \min_pooling_0/n366 , \min_pooling_0/n365 ,
         \min_pooling_0/n362 , \min_pooling_0/n361 , \min_pooling_0/n358 ,
         \min_pooling_0/n357 , \min_pooling_0/n354 , \min_pooling_0/n353 ,
         \min_pooling_0/n350 , \min_pooling_0/n349 , \min_pooling_0/n346 ,
         \min_pooling_0/n345 , \min_pooling_0/n342 , \min_pooling_0/n341 ,
         \min_pooling_0/n338 , \min_pooling_0/n337 , \min_pooling_0/n334 ,
         \min_pooling_0/n333 , \min_pooling_0/n330 , \min_pooling_0/n329 ,
         \min_pooling_0/n326 , \min_pooling_0/n325 , \min_pooling_0/n322 ,
         \min_pooling_0/n321 , \min_pooling_0/n318 , \min_pooling_0/n317 ,
         \min_pooling_0/n314 , \min_pooling_0/n313 , \min_pooling_0/n310 ,
         \min_pooling_0/n309 , \mean_pooling_0/n244 , \mean_pooling_0/n243 ,
         \mean_pooling_0/n240 , \mean_pooling_0/n239 , \mean_pooling_0/n236 ,
         \mean_pooling_0/n235 , \mean_pooling_0/n232 , \mean_pooling_0/n231 ,
         \mean_pooling_0/n228 , \mean_pooling_0/n227 , \mean_pooling_0/n224 ,
         \mean_pooling_0/n223 , \mean_pooling_0/n220 , \mean_pooling_0/n219 ,
         \mean_pooling_0/n216 , \mean_pooling_0/n215 , \mean_pooling_0/n212 ,
         \mean_pooling_0/n211 , \mean_pooling_0/n208 , \mean_pooling_0/n207 ,
         \mean_pooling_0/n204 , \mean_pooling_0/n203 , \mean_pooling_0/n200 ,
         \mean_pooling_0/n199 , \mean_pooling_0/n196 , \mean_pooling_0/n195 ,
         \mean_pooling_0/n192 , \mean_pooling_0/n191 , \mean_pooling_0/n188 ,
         \mean_pooling_0/n187 , \mean_pooling_0/n184 , \mean_pooling_0/n183 ,
         \mean_pooling_0/n180 , \mean_pooling_0/n179 , \mean_pooling_0/n176 ,
         \mean_pooling_0/n175 , \mean_pooling_0/n172 , \mean_pooling_0/n171 ,
         \mean_pooling_0/n168 , \mean_pooling_0/n167 , \mean_pooling_0/n164 ,
         \mean_pooling_0/n163 , \max_pooling_0/n309 , \max_pooling_0/n308 ,
         \max_pooling_0/n305 , \max_pooling_0/n304 , \max_pooling_0/n301 ,
         \max_pooling_0/n300 , \max_pooling_0/n297 , \max_pooling_0/n296 ,
         \max_pooling_0/n293 , \max_pooling_0/n292 , \max_pooling_0/n289 ,
         \max_pooling_0/n288 , \max_pooling_0/n285 , \max_pooling_0/n284 ,
         \max_pooling_0/n281 , \max_pooling_0/n280 , \max_pooling_0/n277 ,
         \max_pooling_0/n276 , \max_pooling_0/n273 , \max_pooling_0/n272 ,
         \max_pooling_0/n269 , \max_pooling_0/n268 , \max_pooling_0/n265 ,
         \max_pooling_0/n264 , \max_pooling_0/n261 , \max_pooling_0/n260 ,
         \max_pooling_0/n257 , \max_pooling_0/n256 , \max_pooling_0/n253 ,
         \max_pooling_0/n252 , \max_pooling_0/n249 , \max_pooling_0/n248 ,
         \max_pooling_0/n245 , \max_pooling_0/n244 , \max_pooling_0/n241 ,
         \max_pooling_0/n240 , \max_pooling_0/n237 , \max_pooling_0/n236 ,
         \max_pooling_0/n233 , \max_pooling_0/n232 , \max_pooling_0/n229 ,
         \max_pooling_0/n228 , n2821, n2822, n2823, n2824, n2825, n2826, n2827,
         n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837,
         n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847,
         n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857,
         n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867,
         n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877,
         n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887,
         n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897,
         n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907,
         n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917,
         n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927,
         n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937,
         n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947,
         n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957,
         n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967,
         n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977,
         n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987,
         n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997,
         n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007,
         n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017,
         n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027,
         n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037,
         n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047,
         n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057,
         n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067,
         n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077,
         n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087,
         n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097,
         n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107,
         n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117,
         n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127,
         n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137,
         n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147,
         n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157,
         n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167,
         n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177,
         n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187,
         n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197,
         n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207,
         n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217,
         n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227,
         n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237,
         n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247,
         n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3603, n3604, n3605,
         n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615,
         n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625,
         n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635,
         n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645,
         n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655,
         n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665,
         n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675,
         n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685,
         n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695,
         n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705,
         n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715,
         n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725,
         n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735,
         n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745,
         n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753;
  wire   [19:0] om_max;
  wire   [19:0] om_mean;
  wire   [19:0] om_min;

  dff_sg \state_reg[1]  ( .D(n526), .CP(clk), .Q(state[1]) );
  dff_sg \state_reg[0]  ( .D(n525), .CP(clk), .Q(state[0]) );
  dff_sg \reg_im_reg[3][19]  ( .D(n445), .CP(clk), .Q(\reg_im[3][19] ) );
  dff_sg \reg_im_reg[3][18]  ( .D(n446), .CP(clk), .Q(\reg_im[3][18] ) );
  dff_sg \reg_im_reg[3][17]  ( .D(n447), .CP(clk), .Q(\reg_im[3][17] ) );
  dff_sg \reg_im_reg[3][16]  ( .D(n448), .CP(clk), .Q(\reg_im[3][16] ) );
  dff_sg \reg_im_reg[3][15]  ( .D(n449), .CP(clk), .Q(\reg_im[3][15] ) );
  dff_sg \reg_im_reg[3][14]  ( .D(n450), .CP(clk), .Q(\reg_im[3][14] ) );
  dff_sg \reg_im_reg[3][13]  ( .D(n451), .CP(clk), .Q(\reg_im[3][13] ) );
  dff_sg \reg_im_reg[3][12]  ( .D(n452), .CP(clk), .Q(\reg_im[3][12] ) );
  dff_sg \reg_im_reg[3][11]  ( .D(n453), .CP(clk), .Q(\reg_im[3][11] ) );
  dff_sg \reg_im_reg[3][10]  ( .D(n454), .CP(clk), .Q(\reg_im[3][10] ) );
  dff_sg \reg_im_reg[3][9]  ( .D(n455), .CP(clk), .Q(\reg_im[3][9] ) );
  dff_sg \reg_im_reg[3][8]  ( .D(n456), .CP(clk), .Q(\reg_im[3][8] ) );
  dff_sg \reg_im_reg[3][7]  ( .D(n457), .CP(clk), .Q(\reg_im[3][7] ) );
  dff_sg \reg_im_reg[3][6]  ( .D(n458), .CP(clk), .Q(\reg_im[3][6] ) );
  dff_sg \reg_im_reg[3][5]  ( .D(n459), .CP(clk), .Q(\reg_im[3][5] ) );
  dff_sg \reg_im_reg[3][4]  ( .D(n460), .CP(clk), .Q(\reg_im[3][4] ) );
  dff_sg \reg_im_reg[3][3]  ( .D(n461), .CP(clk), .Q(\reg_im[3][3] ) );
  dff_sg \reg_im_reg[3][2]  ( .D(n462), .CP(clk), .Q(\reg_im[3][2] ) );
  dff_sg \reg_im_reg[3][1]  ( .D(n463), .CP(clk), .Q(\reg_im[3][1] ) );
  dff_sg \reg_im_reg[3][0]  ( .D(n464), .CP(clk), .Q(\reg_im[3][0] ) );
  dff_sg \reg_im_reg[2][19]  ( .D(n465), .CP(clk), .Q(\reg_im[2][19] ) );
  dff_sg \reg_im_reg[2][18]  ( .D(n466), .CP(clk), .Q(\reg_im[2][18] ) );
  dff_sg \reg_im_reg[2][17]  ( .D(n467), .CP(clk), .Q(\reg_im[2][17] ) );
  dff_sg \reg_im_reg[2][16]  ( .D(n468), .CP(clk), .Q(\reg_im[2][16] ) );
  dff_sg \reg_im_reg[2][15]  ( .D(n469), .CP(clk), .Q(\reg_im[2][15] ) );
  dff_sg \reg_im_reg[2][14]  ( .D(n470), .CP(clk), .Q(\reg_im[2][14] ) );
  dff_sg \reg_im_reg[2][13]  ( .D(n471), .CP(clk), .Q(\reg_im[2][13] ) );
  dff_sg \reg_im_reg[2][12]  ( .D(n472), .CP(clk), .Q(\reg_im[2][12] ) );
  dff_sg \reg_im_reg[2][11]  ( .D(n473), .CP(clk), .Q(\reg_im[2][11] ) );
  dff_sg \reg_im_reg[2][10]  ( .D(n474), .CP(clk), .Q(\reg_im[2][10] ) );
  dff_sg \reg_im_reg[2][9]  ( .D(n475), .CP(clk), .Q(\reg_im[2][9] ) );
  dff_sg \reg_im_reg[2][8]  ( .D(n476), .CP(clk), .Q(\reg_im[2][8] ) );
  dff_sg \reg_im_reg[2][7]  ( .D(n477), .CP(clk), .Q(\reg_im[2][7] ) );
  dff_sg \reg_im_reg[2][6]  ( .D(n478), .CP(clk), .Q(\reg_im[2][6] ) );
  dff_sg \reg_im_reg[2][5]  ( .D(n479), .CP(clk), .Q(\reg_im[2][5] ) );
  dff_sg \reg_im_reg[2][4]  ( .D(n480), .CP(clk), .Q(\reg_im[2][4] ) );
  dff_sg \reg_im_reg[2][3]  ( .D(n481), .CP(clk), .Q(\reg_im[2][3] ) );
  dff_sg \reg_im_reg[2][2]  ( .D(n482), .CP(clk), .Q(\reg_im[2][2] ) );
  dff_sg \reg_im_reg[2][1]  ( .D(n483), .CP(clk), .Q(\reg_im[2][1] ) );
  dff_sg \reg_im_reg[2][0]  ( .D(n484), .CP(clk), .Q(\reg_im[2][0] ) );
  dff_sg \reg_im_reg[1][19]  ( .D(n485), .CP(clk), .Q(\reg_im[1][19] ) );
  dff_sg \reg_im_reg[1][18]  ( .D(n486), .CP(clk), .Q(\reg_im[1][18] ) );
  dff_sg \reg_im_reg[1][17]  ( .D(n487), .CP(clk), .Q(\reg_im[1][17] ) );
  dff_sg \reg_im_reg[1][16]  ( .D(n488), .CP(clk), .Q(\reg_im[1][16] ) );
  dff_sg \reg_im_reg[1][15]  ( .D(n489), .CP(clk), .Q(\reg_im[1][15] ) );
  dff_sg \reg_im_reg[1][14]  ( .D(n490), .CP(clk), .Q(\reg_im[1][14] ) );
  dff_sg \reg_im_reg[1][13]  ( .D(n491), .CP(clk), .Q(\reg_im[1][13] ) );
  dff_sg \reg_im_reg[1][12]  ( .D(n492), .CP(clk), .Q(\reg_im[1][12] ) );
  dff_sg \reg_im_reg[1][11]  ( .D(n493), .CP(clk), .Q(\reg_im[1][11] ) );
  dff_sg \reg_im_reg[1][10]  ( .D(n494), .CP(clk), .Q(\reg_im[1][10] ) );
  dff_sg \reg_im_reg[1][9]  ( .D(n495), .CP(clk), .Q(\reg_im[1][9] ) );
  dff_sg \reg_im_reg[1][8]  ( .D(n496), .CP(clk), .Q(\reg_im[1][8] ) );
  dff_sg \reg_im_reg[1][7]  ( .D(n497), .CP(clk), .Q(\reg_im[1][7] ) );
  dff_sg \reg_im_reg[1][6]  ( .D(n498), .CP(clk), .Q(\reg_im[1][6] ) );
  dff_sg \reg_im_reg[1][5]  ( .D(n499), .CP(clk), .Q(\reg_im[1][5] ) );
  dff_sg \reg_im_reg[1][4]  ( .D(n500), .CP(clk), .Q(\reg_im[1][4] ) );
  dff_sg \reg_im_reg[1][3]  ( .D(n501), .CP(clk), .Q(\reg_im[1][3] ) );
  dff_sg \reg_im_reg[1][2]  ( .D(n502), .CP(clk), .Q(\reg_im[1][2] ) );
  dff_sg \reg_im_reg[1][1]  ( .D(n503), .CP(clk), .Q(\reg_im[1][1] ) );
  dff_sg \reg_im_reg[1][0]  ( .D(n504), .CP(clk), .Q(\reg_im[1][0] ) );
  dff_sg \reg_im_reg[0][19]  ( .D(n505), .CP(clk), .Q(\reg_im[0][19] ) );
  dff_sg \reg_im_reg[0][18]  ( .D(n506), .CP(clk), .Q(\reg_im[0][18] ) );
  dff_sg \reg_im_reg[0][17]  ( .D(n507), .CP(clk), .Q(\reg_im[0][17] ) );
  dff_sg \reg_im_reg[0][16]  ( .D(n508), .CP(clk), .Q(\reg_im[0][16] ) );
  dff_sg \reg_im_reg[0][15]  ( .D(n509), .CP(clk), .Q(\reg_im[0][15] ) );
  dff_sg \reg_im_reg[0][14]  ( .D(n510), .CP(clk), .Q(\reg_im[0][14] ) );
  dff_sg \reg_im_reg[0][13]  ( .D(n511), .CP(clk), .Q(\reg_im[0][13] ) );
  dff_sg \reg_im_reg[0][12]  ( .D(n512), .CP(clk), .Q(\reg_im[0][12] ) );
  dff_sg \reg_im_reg[0][11]  ( .D(n513), .CP(clk), .Q(\reg_im[0][11] ) );
  dff_sg \reg_im_reg[0][10]  ( .D(n514), .CP(clk), .Q(\reg_im[0][10] ) );
  dff_sg \reg_im_reg[0][9]  ( .D(n515), .CP(clk), .Q(\reg_im[0][9] ) );
  dff_sg \reg_im_reg[0][8]  ( .D(n516), .CP(clk), .Q(\reg_im[0][8] ) );
  dff_sg \reg_im_reg[0][7]  ( .D(n517), .CP(clk), .Q(\reg_im[0][7] ) );
  dff_sg \reg_im_reg[0][6]  ( .D(n518), .CP(clk), .Q(\reg_im[0][6] ) );
  dff_sg \reg_im_reg[0][5]  ( .D(n519), .CP(clk), .Q(\reg_im[0][5] ) );
  dff_sg \reg_im_reg[0][4]  ( .D(n520), .CP(clk), .Q(\reg_im[0][4] ) );
  dff_sg \reg_im_reg[0][3]  ( .D(n521), .CP(clk), .Q(\reg_im[0][3] ) );
  dff_sg \reg_im_reg[0][2]  ( .D(n522), .CP(clk), .Q(\reg_im[0][2] ) );
  dff_sg \reg_im_reg[0][1]  ( .D(n523), .CP(clk), .Q(\reg_im[0][1] ) );
  dff_sg \reg_im_reg[0][0]  ( .D(n524), .CP(clk), .Q(\reg_im[0][0] ) );
  dff_sg reg_input_ready_reg ( .D(N112), .CP(clk), .Q(reg_input_ready) );
  dff_sg \max_pooling_0/om_reg[1]  ( .D(\max_pooling_0/n331 ), .CP(clk), .Q(
        om_max[1]) );
  dff_sg \max_pooling_0/om_reg[2]  ( .D(\max_pooling_0/n332 ), .CP(clk), .Q(
        om_max[2]) );
  dff_sg \max_pooling_0/om_reg[3]  ( .D(\max_pooling_0/n333 ), .CP(clk), .Q(
        om_max[3]) );
  dff_sg \max_pooling_0/om_reg[4]  ( .D(\max_pooling_0/n334 ), .CP(clk), .Q(
        \max_pooling_0/n643 ) );
  dff_sg \max_pooling_0/om_reg[5]  ( .D(\max_pooling_0/n335 ), .CP(clk), .Q(
        om_max[5]) );
  dff_sg \max_pooling_0/om_reg[6]  ( .D(\max_pooling_0/n336 ), .CP(clk), .Q(
        \max_pooling_0/n642 ) );
  dff_sg \max_pooling_0/om_reg[7]  ( .D(\max_pooling_0/n337 ), .CP(clk), .Q(
        om_max[7]) );
  dff_sg \max_pooling_0/om_reg[8]  ( .D(\max_pooling_0/n338 ), .CP(clk), .Q(
        \max_pooling_0/n641 ) );
  dff_sg \max_pooling_0/om_reg[9]  ( .D(\max_pooling_0/n339 ), .CP(clk), .Q(
        om_max[9]) );
  dff_sg \max_pooling_0/om_reg[10]  ( .D(\max_pooling_0/n340 ), .CP(clk), .Q(
        \max_pooling_0/n640 ) );
  dff_sg \max_pooling_0/om_reg[11]  ( .D(\max_pooling_0/n341 ), .CP(clk), .Q(
        om_max[11]) );
  dff_sg \max_pooling_0/om_reg[12]  ( .D(\max_pooling_0/n342 ), .CP(clk), .Q(
        \max_pooling_0/n639 ) );
  dff_sg \max_pooling_0/om_reg[13]  ( .D(\max_pooling_0/n343 ), .CP(clk), .Q(
        om_max[13]) );
  dff_sg \max_pooling_0/om_reg[14]  ( .D(\max_pooling_0/n344 ), .CP(clk), .Q(
        om_max[14]) );
  dff_sg \max_pooling_0/om_reg[15]  ( .D(\max_pooling_0/n345 ), .CP(clk), .Q(
        om_max[15]) );
  dff_sg \max_pooling_0/om_reg[16]  ( .D(\max_pooling_0/n346 ), .CP(clk), .Q(
        om_max[16]) );
  dff_sg \max_pooling_0/om_reg[17]  ( .D(\max_pooling_0/n347 ), .CP(clk), .Q(
        om_max[17]) );
  dff_sg \max_pooling_0/om_reg[18]  ( .D(\max_pooling_0/n348 ), .CP(clk), .Q(
        om_max[18]) );
  dff_sg \max_pooling_0/om_reg[19]  ( .D(\max_pooling_0/n349 ), .CP(clk), .Q(
        om_max[19]) );
  dff_sg \max_pooling_0/om_reg[0]  ( .D(\max_pooling_0/n350 ), .CP(clk), .Q(
        om_max[0]) );
  dff_sg \max_pooling_0/pointer_reg[1]  ( .D(\max_pooling_0/n351 ), .CP(clk), 
        .Q(\max_pooling_0/N4 ) );
  dff_sg \max_pooling_0/pointer_reg[0]  ( .D(\max_pooling_0/n352 ), .CP(clk), 
        .Q(\max_pooling_0/N3 ) );
  dff_sg \mean_pooling_0/om_reg[17]  ( .D(\mean_pooling_0/n248 ), .CP(clk), 
        .Q(om_mean[17]) );
  dff_sg \mean_pooling_0/om_reg[16]  ( .D(\mean_pooling_0/n249 ), .CP(clk), 
        .Q(om_mean[16]) );
  dff_sg \mean_pooling_0/om_reg[15]  ( .D(\mean_pooling_0/n250 ), .CP(clk), 
        .Q(om_mean[15]) );
  dff_sg \mean_pooling_0/om_reg[14]  ( .D(\mean_pooling_0/n251 ), .CP(clk), 
        .Q(om_mean[14]) );
  dff_sg \mean_pooling_0/om_reg[13]  ( .D(\mean_pooling_0/n252 ), .CP(clk), 
        .Q(om_mean[13]) );
  dff_sg \mean_pooling_0/om_reg[12]  ( .D(\mean_pooling_0/n253 ), .CP(clk), 
        .Q(om_mean[12]) );
  dff_sg \mean_pooling_0/om_reg[11]  ( .D(\mean_pooling_0/n254 ), .CP(clk), 
        .Q(om_mean[11]) );
  dff_sg \mean_pooling_0/om_reg[10]  ( .D(\mean_pooling_0/n255 ), .CP(clk), 
        .Q(om_mean[10]) );
  dff_sg \mean_pooling_0/om_reg[9]  ( .D(\mean_pooling_0/n256 ), .CP(clk), .Q(
        om_mean[9]) );
  dff_sg \mean_pooling_0/om_reg[8]  ( .D(\mean_pooling_0/n257 ), .CP(clk), .Q(
        om_mean[8]) );
  dff_sg \mean_pooling_0/om_reg[7]  ( .D(\mean_pooling_0/n258 ), .CP(clk), .Q(
        om_mean[7]) );
  dff_sg \mean_pooling_0/om_reg[6]  ( .D(\mean_pooling_0/n259 ), .CP(clk), .Q(
        om_mean[6]) );
  dff_sg \mean_pooling_0/om_reg[5]  ( .D(\mean_pooling_0/n260 ), .CP(clk), .Q(
        om_mean[5]) );
  dff_sg \mean_pooling_0/om_reg[4]  ( .D(\mean_pooling_0/n261 ), .CP(clk), .Q(
        om_mean[4]) );
  dff_sg \mean_pooling_0/om_reg[3]  ( .D(\mean_pooling_0/n262 ), .CP(clk), .Q(
        om_mean[3]) );
  dff_sg \mean_pooling_0/om_reg[2]  ( .D(\mean_pooling_0/n263 ), .CP(clk), .Q(
        om_mean[2]) );
  dff_sg \mean_pooling_0/om_reg[1]  ( .D(\mean_pooling_0/n264 ), .CP(clk), .Q(
        om_mean[1]) );
  dff_sg \mean_pooling_0/om_reg[0]  ( .D(\mean_pooling_0/n265 ), .CP(clk), .Q(
        om_mean[0]) );
  dff_sg \mean_pooling_0/pointer_reg[1]  ( .D(\mean_pooling_0/n246 ), .CP(clk), 
        .Q(\mean_pooling_0/N5 ) );
  dff_sg \mean_pooling_0/pointer_reg[0]  ( .D(\mean_pooling_0/n247 ), .CP(clk), 
        .Q(\mean_pooling_0/N4 ) );
  dff_sg \min_pooling_0/om_reg[1]  ( .D(\min_pooling_0/n392 ), .CP(clk), .Q(
        om_min[1]) );
  dff_sg \min_pooling_0/om_reg[2]  ( .D(\min_pooling_0/n393 ), .CP(clk), .Q(
        \min_pooling_0/n724 ) );
  dff_sg \min_pooling_0/om_reg[3]  ( .D(\min_pooling_0/n394 ), .CP(clk), .Q(
        om_min[3]) );
  dff_sg \min_pooling_0/om_reg[4]  ( .D(\min_pooling_0/n395 ), .CP(clk), .Q(
        om_min[4]) );
  dff_sg \min_pooling_0/om_reg[5]  ( .D(\min_pooling_0/n396 ), .CP(clk), .Q(
        om_min[5]) );
  dff_sg \min_pooling_0/om_reg[6]  ( .D(\min_pooling_0/n397 ), .CP(clk), .Q(
        om_min[6]) );
  dff_sg \min_pooling_0/om_reg[7]  ( .D(\min_pooling_0/n398 ), .CP(clk), .Q(
        om_min[7]) );
  dff_sg \min_pooling_0/om_reg[8]  ( .D(\min_pooling_0/n399 ), .CP(clk), .Q(
        om_min[8]) );
  dff_sg \min_pooling_0/om_reg[9]  ( .D(\min_pooling_0/n400 ), .CP(clk), .Q(
        om_min[9]) );
  dff_sg \min_pooling_0/om_reg[10]  ( .D(\min_pooling_0/n401 ), .CP(clk), .Q(
        om_min[10]) );
  dff_sg \min_pooling_0/om_reg[11]  ( .D(\min_pooling_0/n402 ), .CP(clk), .Q(
        om_min[11]) );
  dff_sg \min_pooling_0/om_reg[12]  ( .D(\min_pooling_0/n403 ), .CP(clk), .Q(
        om_min[12]) );
  dff_sg \min_pooling_0/om_reg[13]  ( .D(\min_pooling_0/n404 ), .CP(clk), .Q(
        om_min[13]) );
  dff_sg \min_pooling_0/om_reg[14]  ( .D(\min_pooling_0/n405 ), .CP(clk), .Q(
        \min_pooling_0/n723 ) );
  dff_sg \min_pooling_0/om_reg[15]  ( .D(\min_pooling_0/n406 ), .CP(clk), .Q(
        om_min[15]) );
  dff_sg \min_pooling_0/om_reg[16]  ( .D(\min_pooling_0/n407 ), .CP(clk), .Q(
        \min_pooling_0/n722 ) );
  dff_sg \min_pooling_0/om_reg[17]  ( .D(\min_pooling_0/n408 ), .CP(clk), .Q(
        om_min[17]) );
  dff_sg \min_pooling_0/om_reg[18]  ( .D(\min_pooling_0/n409 ), .CP(clk), .Q(
        om_min[18]) );
  dff_sg \min_pooling_0/om_reg[19]  ( .D(\min_pooling_0/n410 ), .CP(clk), .Q(
        om_min[19]) );
  dff_sg \min_pooling_0/om_reg[0]  ( .D(\min_pooling_0/n411 ), .CP(clk), .Q(
        om_min[0]) );
  dff_sg \min_pooling_0/pointer_reg[1]  ( .D(\min_pooling_0/n412 ), .CP(clk), 
        .Q(\min_pooling_0/N4 ) );
  dff_sg \min_pooling_0/pointer_reg[0]  ( .D(\min_pooling_0/n413 ), .CP(clk), 
        .Q(\min_pooling_0/N3 ) );
  \**FFGEN**  \om_reg[0]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(
        1'b0), .force_01(n349), .force_10(n3141), .force_11(1'b0), .Q(om[0])
         );
  \**FFGEN**  \om_reg[1]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(
        1'b0), .force_01(n397), .force_10(n3140), .force_11(1'b0), .Q(om[1])
         );
  \**FFGEN**  \om_reg[2]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(
        1'b0), .force_01(n393), .force_10(n3159), .force_11(1'b0), .Q(om[2])
         );
  \**FFGEN**  \om_reg[3]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(
        1'b0), .force_01(n389), .force_10(n3154), .force_11(1'b0), .Q(om[3])
         );
  \**FFGEN**  \om_reg[4]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(
        1'b0), .force_01(n385), .force_10(n3143), .force_11(1'b0), .Q(om[4])
         );
  \**FFGEN**  \om_reg[5]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(
        1'b0), .force_01(n381), .force_10(n3155), .force_11(1'b0), .Q(om[5])
         );
  \**FFGEN**  \om_reg[6]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(
        1'b0), .force_01(n377), .force_10(n3156), .force_11(1'b0), .Q(om[6])
         );
  \**FFGEN**  \om_reg[7]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(
        1'b0), .force_01(n373), .force_10(n3168), .force_11(1'b0), .Q(om[7])
         );
  \**FFGEN**  \om_reg[8]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(
        1'b0), .force_01(n369), .force_10(n3142), .force_11(1'b0), .Q(om[8])
         );
  \**FFGEN**  \om_reg[9]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(
        1'b0), .force_01(n365), .force_10(n3160), .force_11(1'b0), .Q(om[9])
         );
  \**FFGEN**  \om_reg[10]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(
        1'b0), .force_01(n361), .force_10(n3157), .force_11(1'b0), .Q(om[10])
         );
  \**FFGEN**  \om_reg[11]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(
        1'b0), .force_01(n357), .force_10(n3144), .force_11(1'b0), .Q(om[11])
         );
  \**FFGEN**  \om_reg[12]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(
        1'b0), .force_01(n353), .force_10(n3161), .force_11(1'b0), .Q(om[12])
         );
  \**FFGEN**  \om_reg[13]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(
        1'b0), .force_01(n441), .force_10(n3162), .force_11(1'b0), .Q(om[13])
         );
  \**FFGEN**  \om_reg[14]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(
        1'b0), .force_01(n437), .force_10(n3169), .force_11(1'b0), .Q(om[14])
         );
  \**FFGEN**  \om_reg[15]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(
        1'b0), .force_01(n433), .force_10(n3163), .force_11(1'b0), .Q(om[15])
         );
  \**FFGEN**  \om_reg[16]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(
        1'b0), .force_01(n429), .force_10(n3170), .force_11(1'b0), .Q(om[16])
         );
  \**FFGEN**  \om_reg[17]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(
        1'b0), .force_01(n425), .force_10(n3171), .force_11(1'b0), .Q(om[17])
         );
  \**FFGEN**  \om_reg[18]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(
        1'b0), .force_01(n421), .force_10(n422), .force_11(1'b0), .Q(om[18])
         );
  \**FFGEN**  \om_reg[19]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(
        1'b0), .force_01(n417), .force_10(n418), .force_11(1'b0), .Q(om[19])
         );
  \**FFGEN**  en_mean_reg ( .next_state(1'b0), .clocked_on(1'b0), .force_00(
        1'b0), .force_01(n413), .force_10(n414), .force_11(1'b0), .Q(n3252), 
        .QN(n2820) );
  \**FFGEN**  en_max_reg ( .next_state(1'b0), .clocked_on(1'b0), .force_00(
        1'b0), .force_01(n1093), .force_10(n410), .force_11(1'b0), .QN(n2819)
         );
  \**FFGEN**  en_min_reg ( .next_state(1'b0), .clocked_on(1'b0), .force_00(
        1'b0), .force_01(n405), .force_10(n406), .force_11(1'b0), .Q(n2824), 
        .QN(n2818) );
  \**FFGEN**  done_reg ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), 
        .force_01(n401), .force_10(n3172), .force_11(1'b0), .Q(n444) );
  \**FFGEN**  \max_pooling_0/done_reg  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\max_pooling_0/n232 ), .force_10(
        \max_pooling_0/n233 ), .force_11(1'b0), .QN(n1116) );
  \**FFGEN**  \max_pooling_0/max_num_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\max_pooling_0/n236 ), .force_10(
        \max_pooling_0/n237 ), .force_11(1'b0), .Q(\max_pooling_0/n330 ) );
  \**FFGEN**  \max_pooling_0/max_num_reg[19]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\max_pooling_0/n240 ), 
        .force_10(\max_pooling_0/n241 ), .force_11(1'b0), .Q(
        \max_pooling_0/n329 ) );
  \**FFGEN**  \max_pooling_0/max_num_reg[18]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\max_pooling_0/n244 ), 
        .force_10(\max_pooling_0/n245 ), .force_11(1'b0), .Q(
        \max_pooling_0/n328 ) );
  \**FFGEN**  \max_pooling_0/max_num_reg[17]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\max_pooling_0/n248 ), 
        .force_10(\max_pooling_0/n249 ), .force_11(1'b0), .Q(
        \max_pooling_0/n327 ) );
  \**FFGEN**  \max_pooling_0/max_num_reg[16]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\max_pooling_0/n252 ), 
        .force_10(\max_pooling_0/n253 ), .force_11(1'b0), .Q(
        \max_pooling_0/n326 ) );
  \**FFGEN**  \max_pooling_0/max_num_reg[15]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\max_pooling_0/n256 ), 
        .force_10(\max_pooling_0/n257 ), .force_11(1'b0), .Q(
        \max_pooling_0/n325 ) );
  \**FFGEN**  \max_pooling_0/max_num_reg[14]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\max_pooling_0/n260 ), 
        .force_10(\max_pooling_0/n261 ), .force_11(1'b0), .Q(
        \max_pooling_0/n324 ) );
  \**FFGEN**  \max_pooling_0/max_num_reg[13]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\max_pooling_0/n264 ), 
        .force_10(\max_pooling_0/n265 ), .force_11(1'b0), .Q(
        \max_pooling_0/n323 ) );
  \**FFGEN**  \max_pooling_0/max_num_reg[12]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\max_pooling_0/n268 ), 
        .force_10(\max_pooling_0/n269 ), .force_11(1'b0), .Q(
        \max_pooling_0/n322 ) );
  \**FFGEN**  \max_pooling_0/max_num_reg[11]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\max_pooling_0/n272 ), 
        .force_10(\max_pooling_0/n273 ), .force_11(1'b0), .Q(
        \max_pooling_0/n321 ) );
  \**FFGEN**  \max_pooling_0/max_num_reg[10]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\max_pooling_0/n276 ), 
        .force_10(\max_pooling_0/n277 ), .force_11(1'b0), .Q(
        \max_pooling_0/n320 ) );
  \**FFGEN**  \max_pooling_0/max_num_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\max_pooling_0/n280 ), .force_10(
        \max_pooling_0/n281 ), .force_11(1'b0), .Q(\max_pooling_0/n319 ) );
  \**FFGEN**  \max_pooling_0/max_num_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\max_pooling_0/n284 ), .force_10(
        \max_pooling_0/n285 ), .force_11(1'b0), .Q(\max_pooling_0/n318 ) );
  \**FFGEN**  \max_pooling_0/max_num_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\max_pooling_0/n288 ), .force_10(
        \max_pooling_0/n289 ), .force_11(1'b0), .Q(\max_pooling_0/n317 ) );
  \**FFGEN**  \max_pooling_0/max_num_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\max_pooling_0/n292 ), .force_10(
        \max_pooling_0/n293 ), .force_11(1'b0), .Q(\max_pooling_0/n316 ) );
  \**FFGEN**  \max_pooling_0/max_num_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\max_pooling_0/n296 ), .force_10(
        \max_pooling_0/n297 ), .force_11(1'b0), .Q(\max_pooling_0/n315 ) );
  \**FFGEN**  \max_pooling_0/max_num_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\max_pooling_0/n300 ), .force_10(
        \max_pooling_0/n301 ), .force_11(1'b0), .Q(\max_pooling_0/n314 ) );
  \**FFGEN**  \max_pooling_0/max_num_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\max_pooling_0/n304 ), .force_10(
        \max_pooling_0/n305 ), .force_11(1'b0), .Q(\max_pooling_0/n313 ) );
  \**FFGEN**  \max_pooling_0/max_num_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\max_pooling_0/n308 ), .force_10(
        \max_pooling_0/n309 ), .force_11(1'b0), .Q(\max_pooling_0/n312 ) );
  \**FFGEN**  \max_pooling_0/max_num_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\max_pooling_0/n228 ), .force_10(
        \max_pooling_0/n229 ), .force_11(1'b0), .Q(\max_pooling_0/n311 ) );
  \**FFGEN**  \mean_pooling_0/done_reg  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\mean_pooling_0/n167 ), .force_10(
        \mean_pooling_0/n168 ), .force_11(1'b0), .Q(n2841) );
  \**FFGEN**  \mean_pooling_0/sum_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\mean_pooling_0/n171 ), .force_10(
        \mean_pooling_0/n172 ), .force_11(1'b0), .Q(n2825), .QN(n1094) );
  \**FFGEN**  \mean_pooling_0/sum_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\mean_pooling_0/n175 ), .force_10(
        \mean_pooling_0/n176 ), .force_11(1'b0), .Q(n2842), .QN(n1095) );
  \**FFGEN**  \mean_pooling_0/sum_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\mean_pooling_0/n179 ), .force_10(
        \mean_pooling_0/n180 ), .force_11(1'b0), .Q(n2822), .QN(n1096) );
  \**FFGEN**  \mean_pooling_0/sum_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\mean_pooling_0/n183 ), .force_10(
        \mean_pooling_0/n184 ), .force_11(1'b0), .Q(n2826), .QN(n1097) );
  \**FFGEN**  \mean_pooling_0/sum_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\mean_pooling_0/n187 ), .force_10(
        \mean_pooling_0/n188 ), .force_11(1'b0), .Q(n2840), .QN(n1098) );
  \**FFGEN**  \mean_pooling_0/sum_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\mean_pooling_0/n191 ), .force_10(
        \mean_pooling_0/n192 ), .force_11(1'b0), .Q(n2839), .QN(n1099) );
  \**FFGEN**  \mean_pooling_0/sum_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\mean_pooling_0/n195 ), .force_10(
        \mean_pooling_0/n196 ), .force_11(1'b0), .Q(n2838), .QN(n1100) );
  \**FFGEN**  \mean_pooling_0/sum_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\mean_pooling_0/n199 ), .force_10(
        \mean_pooling_0/n200 ), .force_11(1'b0), .Q(n2837), .QN(n1101) );
  \**FFGEN**  \mean_pooling_0/sum_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\mean_pooling_0/n203 ), .force_10(
        \mean_pooling_0/n204 ), .force_11(1'b0), .Q(n2836), .QN(n1102) );
  \**FFGEN**  \mean_pooling_0/sum_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\mean_pooling_0/n207 ), .force_10(
        \mean_pooling_0/n208 ), .force_11(1'b0), .Q(n2835), .QN(n1103) );
  \**FFGEN**  \mean_pooling_0/sum_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\mean_pooling_0/n211 ), .force_10(
        \mean_pooling_0/n212 ), .force_11(1'b0), .Q(n2834), .QN(n1104) );
  \**FFGEN**  \mean_pooling_0/sum_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\mean_pooling_0/n215 ), .force_10(
        \mean_pooling_0/n216 ), .force_11(1'b0), .Q(n2833), .QN(n1105) );
  \**FFGEN**  \mean_pooling_0/sum_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\mean_pooling_0/n219 ), .force_10(
        \mean_pooling_0/n220 ), .force_11(1'b0), .Q(n2832), .QN(n1106) );
  \**FFGEN**  \mean_pooling_0/sum_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\mean_pooling_0/n223 ), .force_10(
        \mean_pooling_0/n224 ), .force_11(1'b0), .Q(n2831), .QN(n1107) );
  \**FFGEN**  \mean_pooling_0/sum_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\mean_pooling_0/n227 ), .force_10(
        \mean_pooling_0/n228 ), .force_11(1'b0), .Q(n2830), .QN(n1108) );
  \**FFGEN**  \mean_pooling_0/sum_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\mean_pooling_0/n231 ), .force_10(
        \mean_pooling_0/n232 ), .force_11(1'b0), .Q(n2829), .QN(n1109) );
  \**FFGEN**  \mean_pooling_0/sum_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\mean_pooling_0/n235 ), .force_10(
        \mean_pooling_0/n236 ), .force_11(1'b0), .Q(n2828), .QN(n1110) );
  \**FFGEN**  \mean_pooling_0/sum_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\mean_pooling_0/n239 ), .force_10(
        \mean_pooling_0/n240 ), .force_11(1'b0), .Q(n2827), .QN(n1111) );
  \**FFGEN**  \mean_pooling_0/sum_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\mean_pooling_0/n243 ), .force_10(
        \mean_pooling_0/n244 ), .force_11(1'b0), .Q(n2823), .QN(n1112) );
  \**FFGEN**  \mean_pooling_0/sum_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\mean_pooling_0/n163 ), .force_10(
        \mean_pooling_0/n164 ), .force_11(1'b0), .Q(n2821), .QN(n1113) );
  \**FFGEN**  \min_pooling_0/done_reg  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\min_pooling_0/n313 ), .force_10(
        \min_pooling_0/n314 ), .force_11(1'b0), .QN(n1115) );
  \**FFGEN**  \min_pooling_0/min_num_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\min_pooling_0/n317 ), .force_10(
        \min_pooling_0/n318 ), .force_11(1'b0), .QN(\min_pooling_0/n265 ) );
  \**FFGEN**  \min_pooling_0/min_num_reg[19]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\min_pooling_0/n321 ), 
        .force_10(\min_pooling_0/n322 ), .force_11(1'b0), .QN(
        \min_pooling_0/n264 ) );
  \**FFGEN**  \min_pooling_0/min_num_reg[18]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\min_pooling_0/n325 ), 
        .force_10(\min_pooling_0/n326 ), .force_11(1'b0), .QN(
        \min_pooling_0/n263 ) );
  \**FFGEN**  \min_pooling_0/min_num_reg[17]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\min_pooling_0/n329 ), 
        .force_10(\min_pooling_0/n330 ), .force_11(1'b0), .QN(
        \min_pooling_0/n262 ) );
  \**FFGEN**  \min_pooling_0/min_num_reg[16]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\min_pooling_0/n333 ), 
        .force_10(\min_pooling_0/n334 ), .force_11(1'b0), .QN(
        \min_pooling_0/n261 ) );
  \**FFGEN**  \min_pooling_0/min_num_reg[15]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\min_pooling_0/n337 ), 
        .force_10(\min_pooling_0/n338 ), .force_11(1'b0), .QN(
        \min_pooling_0/n260 ) );
  \**FFGEN**  \min_pooling_0/min_num_reg[14]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\min_pooling_0/n341 ), 
        .force_10(\min_pooling_0/n342 ), .force_11(1'b0), .QN(
        \min_pooling_0/n259 ) );
  \**FFGEN**  \min_pooling_0/min_num_reg[13]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\min_pooling_0/n345 ), 
        .force_10(\min_pooling_0/n346 ), .force_11(1'b0), .QN(
        \min_pooling_0/n258 ) );
  \**FFGEN**  \min_pooling_0/min_num_reg[12]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\min_pooling_0/n349 ), 
        .force_10(\min_pooling_0/n350 ), .force_11(1'b0), .QN(
        \min_pooling_0/n257 ) );
  \**FFGEN**  \min_pooling_0/min_num_reg[11]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\min_pooling_0/n353 ), 
        .force_10(\min_pooling_0/n354 ), .force_11(1'b0), .QN(
        \min_pooling_0/n256 ) );
  \**FFGEN**  \min_pooling_0/min_num_reg[10]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\min_pooling_0/n357 ), 
        .force_10(\min_pooling_0/n358 ), .force_11(1'b0), .QN(
        \min_pooling_0/n255 ) );
  \**FFGEN**  \min_pooling_0/min_num_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\min_pooling_0/n361 ), .force_10(
        \min_pooling_0/n362 ), .force_11(1'b0), .QN(\min_pooling_0/n254 ) );
  \**FFGEN**  \min_pooling_0/min_num_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\min_pooling_0/n365 ), .force_10(
        \min_pooling_0/n366 ), .force_11(1'b0), .QN(\min_pooling_0/n253 ) );
  \**FFGEN**  \min_pooling_0/min_num_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\min_pooling_0/n369 ), .force_10(
        \min_pooling_0/n370 ), .force_11(1'b0), .QN(\min_pooling_0/n252 ) );
  \**FFGEN**  \min_pooling_0/min_num_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\min_pooling_0/n373 ), .force_10(
        \min_pooling_0/n374 ), .force_11(1'b0), .QN(\min_pooling_0/n251 ) );
  \**FFGEN**  \min_pooling_0/min_num_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\min_pooling_0/n377 ), .force_10(
        \min_pooling_0/n378 ), .force_11(1'b0), .QN(\min_pooling_0/n250 ) );
  \**FFGEN**  \min_pooling_0/min_num_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\min_pooling_0/n381 ), .force_10(
        \min_pooling_0/n382 ), .force_11(1'b0), .QN(\min_pooling_0/n249 ) );
  \**FFGEN**  \min_pooling_0/min_num_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\min_pooling_0/n385 ), .force_10(
        \min_pooling_0/n386 ), .force_11(1'b0), .QN(\min_pooling_0/n248 ) );
  \**FFGEN**  \min_pooling_0/min_num_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\min_pooling_0/n389 ), .force_10(
        \min_pooling_0/n390 ), .force_11(1'b0), .QN(\min_pooling_0/n247 ) );
  \**FFGEN**  \min_pooling_0/min_num_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\min_pooling_0/n309 ), .force_10(
        \min_pooling_0/n310 ), .force_11(1'b0), .QN(\min_pooling_0/n246 ) );
  nand_x8_sg U2221 ( .A(mode[0]), .B(mode[1]), .X(n1147) );
  nand_x1_sg U2897 ( .A(n1678), .B(n1742), .X(n1670) );
  nand_x1_sg U2898 ( .A(n1743), .B(n2842), .X(n1678) );
  inv_x1_sg U2899 ( .A(n1208), .X(n3634) );
  inv_x1_sg U2900 ( .A(n1223), .X(n3647) );
  inv_x1_sg U2901 ( .A(n1243), .X(n3670) );
  inv_x1_sg U2902 ( .A(n1293), .X(n3724) );
  inv_x1_sg U2903 ( .A(n1957), .X(n3727) );
  inv_x1_sg U2904 ( .A(n1218), .X(n3643) );
  nand_x1_sg U2905 ( .A(n2027), .B(n2028), .X(n2024) );
  nand_x1_sg U2906 ( .A(n1365), .B(n1366), .X(n1362) );
  nand_x1_sg U2907 ( .A(n2114), .B(n3687), .X(n2113) );
  nand_x1_sg U2908 ( .A(n2014), .B(n2015), .X(n2013) );
  nand_x1_sg U2909 ( .A(n2112), .B(n2113), .X(n2111) );
  nand_x1_sg U2910 ( .A(n1694), .B(n1695), .X(n1526) );
  nand_x1_sg U2911 ( .A(n1697), .B(n1698), .X(n1535) );
  nand_x1_sg U2912 ( .A(n1700), .B(n1701), .X(n1544) );
  nand_x1_sg U2913 ( .A(n1703), .B(n1704), .X(n1553) );
  nand_x1_sg U2914 ( .A(n1706), .B(n1707), .X(n1562) );
  nand_x1_sg U2915 ( .A(n1709), .B(n1710), .X(n1571) );
  nand_x1_sg U2916 ( .A(n1712), .B(n1713), .X(n1580) );
  nand_x1_sg U2917 ( .A(n1715), .B(n1716), .X(n1589) );
  nand_x1_sg U2918 ( .A(n1718), .B(n1719), .X(n1598) );
  nand_x1_sg U2919 ( .A(n1721), .B(n1722), .X(n1607) );
  nand_x1_sg U2920 ( .A(n1724), .B(n1725), .X(n1616) );
  nand_x1_sg U2921 ( .A(n1727), .B(n1728), .X(n1625) );
  nand_x1_sg U2922 ( .A(n1730), .B(n1731), .X(n1634) );
  nand_x1_sg U2923 ( .A(n1733), .B(n1734), .X(n1643) );
  nand_x1_sg U2924 ( .A(n1736), .B(n1737), .X(n1652) );
  inv_x1_sg U2925 ( .A(n1661), .X(n3636) );
  nand_x1_sg U2926 ( .A(n1853), .B(n1854), .X(n1523) );
  nand_x2_sg U2927 ( .A(n1847), .B(n1848), .X(n1532) );
  nand_x2_sg U2928 ( .A(n1841), .B(n1842), .X(n1541) );
  nand_x2_sg U2929 ( .A(n1835), .B(n1836), .X(n1550) );
  nand_x2_sg U2930 ( .A(n1829), .B(n1830), .X(n1559) );
  nand_x2_sg U2931 ( .A(n1823), .B(n1824), .X(n1568) );
  nand_x2_sg U2932 ( .A(n1817), .B(n1818), .X(n1577) );
  nand_x2_sg U2933 ( .A(n1811), .B(n1812), .X(n1586) );
  nand_x2_sg U2934 ( .A(n1805), .B(n1806), .X(n1595) );
  nand_x2_sg U2935 ( .A(n1799), .B(n1800), .X(n1604) );
  nand_x2_sg U2936 ( .A(n1793), .B(n1794), .X(n1613) );
  nand_x2_sg U2937 ( .A(n1787), .B(n1788), .X(n1622) );
  nand_x2_sg U2938 ( .A(n1781), .B(n1782), .X(n1631) );
  nand_x2_sg U2939 ( .A(n1775), .B(n1776), .X(n1640) );
  nand_x2_sg U2940 ( .A(n1769), .B(n1770), .X(n1649) );
  nand_x2_sg U2941 ( .A(n1763), .B(n1764), .X(n1658) );
  nand_x2_sg U2942 ( .A(n1757), .B(n1758), .X(n1667) );
  nor_x1_sg U2943 ( .A(n1094), .B(n3625), .X(n1675) );
  nand_x2_sg U2944 ( .A(n1387), .B(n1388), .X(n1304) );
  nand_x1_sg U2945 ( .A(n1377), .B(n1378), .X(n1208) );
  nand_x2_sg U2946 ( .A(n1399), .B(n1400), .X(n1213) );
  nand_x1_sg U2947 ( .A(n1406), .B(n1407), .X(n1218) );
  nand_x1_sg U2948 ( .A(n1412), .B(n1413), .X(n1223) );
  inv_x1_sg U2949 ( .A(n1228), .X(n3654) );
  nand_x2_sg U2950 ( .A(n1425), .B(n1426), .X(n1233) );
  nand_x2_sg U2951 ( .A(n1466), .B(n1467), .X(n1238) );
  nand_x1_sg U2952 ( .A(n1460), .B(n1461), .X(n1243) );
  inv_x1_sg U2953 ( .A(n1248), .X(n3677) );
  nand_x2_sg U2954 ( .A(n1479), .B(n1480), .X(n1253) );
  nand_x2_sg U2955 ( .A(n1437), .B(n1438), .X(n1258) );
  nand_x2_sg U2956 ( .A(n1443), .B(n1444), .X(n1263) );
  inv_x1_sg U2957 ( .A(n1268), .X(n3699) );
  nand_x2_sg U2958 ( .A(n1492), .B(n1493), .X(n1273) );
  nand_x2_sg U2959 ( .A(n1323), .B(n1324), .X(n1278) );
  inv_x1_sg U2960 ( .A(n1283), .X(n3715) );
  inv_x1_sg U2961 ( .A(n1288), .X(n3720) );
  nand_x1_sg U2962 ( .A(n1512), .B(n1513), .X(n1293) );
  inv_x1_sg U2963 ( .A(n1298), .X(n3624) );
  inv_x1_sg U2964 ( .A(n1666), .X(n3631) );
  nand_x2_sg U2965 ( .A(n2054), .B(n2055), .X(n1968) );
  inv_x1_sg U2966 ( .A(n1872), .X(n3637) );
  inv_x1_sg U2967 ( .A(n1877), .X(n3642) );
  nand_x2_sg U2968 ( .A(n2067), .B(n2068), .X(n1887) );
  nand_x2_sg U2969 ( .A(n2080), .B(n2081), .X(n1892) );
  inv_x1_sg U2970 ( .A(n1897), .X(n3663) );
  nand_x2_sg U2971 ( .A(n2122), .B(n2123), .X(n1902) );
  nand_x2_sg U2972 ( .A(n2128), .B(n2129), .X(n1907) );
  inv_x1_sg U2973 ( .A(n1912), .X(n3681) );
  inv_x1_sg U2974 ( .A(n1917), .X(n3686) );
  nand_x2_sg U2975 ( .A(n2098), .B(n2099), .X(n1922) );
  nand_x2_sg U2976 ( .A(n2104), .B(n2105), .X(n1927) );
  nand_x2_sg U2977 ( .A(n2148), .B(n2149), .X(n1932) );
  inv_x1_sg U2978 ( .A(n1937), .X(n3708) );
  nand_x2_sg U2979 ( .A(n1986), .B(n1987), .X(n1942) );
  nand_x2_sg U2980 ( .A(n2162), .B(n2163), .X(n1947) );
  nand_x2_sg U2981 ( .A(n2168), .B(n2169), .X(n1952) );
  nand_x1_sg U2982 ( .A(n2174), .B(n2175), .X(n1957) );
  nand_x1_sg U2983 ( .A(n1685), .B(n3252), .X(n1686) );
  nand_x1_sg U2984 ( .A(n1518), .B(n3252), .X(n1519) );
  nand_x1_sg U2985 ( .A(n1527), .B(n3252), .X(n1528) );
  nand_x1_sg U2986 ( .A(n1536), .B(n3252), .X(n1537) );
  nand_x1_sg U2987 ( .A(n1545), .B(n3252), .X(n1546) );
  nand_x1_sg U2988 ( .A(n1554), .B(n3252), .X(n1555) );
  nand_x1_sg U2989 ( .A(n1563), .B(n3252), .X(n1564) );
  nand_x1_sg U2990 ( .A(n1572), .B(n3252), .X(n1573) );
  nand_x1_sg U2991 ( .A(n1581), .B(n3252), .X(n1582) );
  nand_x1_sg U2992 ( .A(n1590), .B(n3252), .X(n1591) );
  nand_x1_sg U2993 ( .A(n1599), .B(n3252), .X(n1600) );
  nand_x1_sg U2994 ( .A(n1608), .B(n3252), .X(n1609) );
  nand_x1_sg U2995 ( .A(n1617), .B(n3252), .X(n1618) );
  nand_x1_sg U2996 ( .A(n1626), .B(n3252), .X(n1627) );
  nand_x1_sg U2997 ( .A(n1635), .B(n3252), .X(n1636) );
  nand_x1_sg U2998 ( .A(n1644), .B(n3252), .X(n1645) );
  nand_x1_sg U2999 ( .A(n1653), .B(n3252), .X(n1654) );
  nand_x1_sg U3000 ( .A(n1662), .B(n3252), .X(n1663) );
  nand_x1_sg U3001 ( .A(n2460), .B(n2456), .X(n2459) );
  nand_x1_sg U3002 ( .A(n2464), .B(n444), .X(n2461) );
  inv_x1_sg U3003 ( .A(n1141), .X(n2843) );
  nor_x4_sg U3004 ( .A(n2844), .B(mode[0]), .X(n1141) );
  inv_x16_sg U3005 ( .A(mode[1]), .X(n2844) );
  inv_x8_sg U3006 ( .A(mode[1]), .X(n3165) );
  inv_x1_sg U3007 ( .A(n2973), .X(n2845) );
  inv_x2_sg U3008 ( .A(n1145), .X(n2846) );
  nand_x16_sg U3009 ( .A(n2817), .B(input_ready), .X(n2463) );
  nor_x1_sg U3010 ( .A(n3165), .B(mode[0]), .X(n2847) );
  inv_x1_sg U3011 ( .A(n3116), .X(n2848) );
  inv_x1_sg U3012 ( .A(n3117), .X(n2849) );
  inv_x1_sg U3013 ( .A(n3118), .X(n2850) );
  inv_x1_sg U3014 ( .A(n3119), .X(n2851) );
  inv_x1_sg U3015 ( .A(n3120), .X(n2852) );
  inv_x1_sg U3016 ( .A(n3121), .X(n2853) );
  inv_x1_sg U3017 ( .A(n3122), .X(n2854) );
  inv_x1_sg U3018 ( .A(n3123), .X(n2855) );
  inv_x1_sg U3019 ( .A(n3124), .X(n2856) );
  inv_x1_sg U3020 ( .A(n3125), .X(n2857) );
  inv_x1_sg U3021 ( .A(n3126), .X(n2858) );
  inv_x1_sg U3022 ( .A(n2963), .X(n2859) );
  inv_x1_sg U3023 ( .A(n2757), .X(n2860) );
  inv_x4_sg U3024 ( .A(n2757), .X(n2968) );
  inv_x1_sg U3025 ( .A(n2968), .X(n2861) );
  inv_x1_sg U3026 ( .A(n1748), .X(n2862) );
  inv_x1_sg U3027 ( .A(n2980), .X(n2863) );
  inv_x1_sg U3028 ( .A(n3250), .X(n2864) );
  inv_x1_sg U3029 ( .A(n2985), .X(n2865) );
  inv_x1_sg U3030 ( .A(n3251), .X(n2866) );
  inv_x1_sg U3031 ( .A(n2990), .X(n2867) );
  inv_x1_sg U3032 ( .A(n2997), .X(n2868) );
  inv_x1_sg U3033 ( .A(n3002), .X(n2869) );
  inv_x1_sg U3034 ( .A(n3007), .X(n2870) );
  inv_x1_sg U3035 ( .A(n3013), .X(n2871) );
  inv_x1_sg U3036 ( .A(n2871), .X(n2872) );
  inv_x1_sg U3037 ( .A(n3017), .X(n2873) );
  inv_x1_sg U3038 ( .A(n2873), .X(n2874) );
  inv_x1_sg U3039 ( .A(n3022), .X(n2875) );
  inv_x1_sg U3040 ( .A(n2875), .X(n2876) );
  inv_x1_sg U3041 ( .A(n3027), .X(n2877) );
  inv_x1_sg U3042 ( .A(n2877), .X(n2878) );
  inv_x1_sg U3043 ( .A(n3032), .X(n2879) );
  inv_x1_sg U3044 ( .A(n2879), .X(n2880) );
  inv_x1_sg U3045 ( .A(n3037), .X(n2881) );
  inv_x1_sg U3046 ( .A(n2881), .X(n2882) );
  inv_x1_sg U3047 ( .A(n3042), .X(n2883) );
  inv_x1_sg U3048 ( .A(n2883), .X(n2884) );
  inv_x1_sg U3049 ( .A(n3254), .X(n2885) );
  inv_x1_sg U3050 ( .A(n2885), .X(n2886) );
  inv_x1_sg U3051 ( .A(n3075), .X(n2887) );
  inv_x1_sg U3052 ( .A(n1870), .X(n2888) );
  inv_x1_sg U3053 ( .A(n2888), .X(n2889) );
  inv_x1_sg U3054 ( .A(n3080), .X(n2890) );
  inv_x1_sg U3055 ( .A(n1207), .X(n2891) );
  inv_x1_sg U3056 ( .A(n2891), .X(n2892) );
  inv_x1_sg U3057 ( .A(n3085), .X(n2893) );
  inv_x1_sg U3058 ( .A(n3129), .X(n2894) );
  inv_x1_sg U3059 ( .A(n2894), .X(n2895) );
  inv_x1_sg U3060 ( .A(n1308), .X(n2896) );
  inv_x1_sg U3061 ( .A(n2467), .X(n2897) );
  inv_x1_sg U3062 ( .A(n3098), .X(n2898) );
  inv_x1_sg U3063 ( .A(n2898), .X(n2899) );
  inv_x1_sg U3064 ( .A(n3100), .X(n2900) );
  inv_x1_sg U3065 ( .A(n2923), .X(n2901) );
  inv_x1_sg U3066 ( .A(n3127), .X(n2902) );
  inv_x1_sg U3067 ( .A(n3012), .X(n2903) );
  inv_x1_sg U3068 ( .A(n3016), .X(n2904) );
  inv_x1_sg U3069 ( .A(n3021), .X(n2905) );
  inv_x1_sg U3070 ( .A(n3026), .X(n2906) );
  inv_x1_sg U3071 ( .A(n3031), .X(n2907) );
  inv_x1_sg U3072 ( .A(n3036), .X(n2908) );
  inv_x1_sg U3073 ( .A(n3041), .X(n2909) );
  inv_x1_sg U3074 ( .A(n2761), .X(n2910) );
  inv_x1_sg U3075 ( .A(n3051), .X(n2911) );
  inv_x1_sg U3076 ( .A(n1965), .X(n2912) );
  inv_x1_sg U3077 ( .A(n2912), .X(n2913) );
  inv_x1_sg U3078 ( .A(n3063), .X(n2914) );
  inv_x1_sg U3079 ( .A(n1301), .X(n2915) );
  inv_x1_sg U3080 ( .A(n2915), .X(n2916) );
  inv_x1_sg U3081 ( .A(n3067), .X(n2917) );
  inv_x1_sg U3082 ( .A(n1684), .X(n2918) );
  inv_x1_sg U3083 ( .A(n2918), .X(n2919) );
  inv_x1_sg U3084 ( .A(n3071), .X(n2920) );
  inv_x1_sg U3085 ( .A(n3094), .X(n2921) );
  inv_x1_sg U3086 ( .A(n3094), .X(n2922) );
  inv_x1_sg U3087 ( .A(n2468), .X(n2923) );
  inv_x1_sg U3088 ( .A(n3099), .X(n2924) );
  inv_x1_sg U3089 ( .A(n3254), .X(n2925) );
  inv_x1_sg U3090 ( .A(n3075), .X(n2926) );
  inv_x1_sg U3091 ( .A(n2925), .X(n2927) );
  inv_x1_sg U3092 ( .A(n1870), .X(n2928) );
  inv_x1_sg U3093 ( .A(n3080), .X(n2929) );
  inv_x1_sg U3094 ( .A(n2928), .X(n2930) );
  inv_x1_sg U3095 ( .A(n1207), .X(n2931) );
  inv_x1_sg U3096 ( .A(n3085), .X(n2932) );
  inv_x1_sg U3097 ( .A(n2931), .X(n2933) );
  inv_x1_sg U3098 ( .A(n3129), .X(n2934) );
  inv_x1_sg U3099 ( .A(n1308), .X(n2935) );
  inv_x1_sg U3100 ( .A(n2934), .X(n2936) );
  inv_x1_sg U3101 ( .A(n2467), .X(n2937) );
  inv_x1_sg U3102 ( .A(n2897), .X(n2938) );
  inv_x1_sg U3103 ( .A(n2937), .X(n2939) );
  inv_x1_sg U3104 ( .A(n2923), .X(n2940) );
  inv_x1_sg U3105 ( .A(n2923), .X(n2941) );
  inv_x1_sg U3106 ( .A(n2924), .X(n2942) );
  inv_x1_sg U3107 ( .A(n3105), .X(n2943) );
  inv_x1_sg U3108 ( .A(n3110), .X(n2944) );
  inv_x1_sg U3109 ( .A(n3110), .X(n2945) );
  inv_x1_sg U3110 ( .A(n1145), .X(n2946) );
  inv_x1_sg U3111 ( .A(n2885), .X(n2947) );
  inv_x1_sg U3112 ( .A(n2885), .X(n2948) );
  inv_x1_sg U3113 ( .A(n2888), .X(n2949) );
  inv_x1_sg U3114 ( .A(n2888), .X(n2950) );
  inv_x1_sg U3115 ( .A(n2891), .X(n2951) );
  inv_x1_sg U3116 ( .A(n2891), .X(n2952) );
  inv_x1_sg U3117 ( .A(n2894), .X(n2953) );
  inv_x1_sg U3118 ( .A(n2894), .X(n2954) );
  inv_x1_sg U3119 ( .A(reg_input_ready), .X(n2955) );
  inv_x1_sg U3120 ( .A(n2955), .X(n2956) );
  inv_x1_sg U3121 ( .A(n2955), .X(n2957) );
  inv_x1_sg U3122 ( .A(n2721), .X(n2958) );
  inv_x1_sg U3123 ( .A(n2958), .X(n2959) );
  inv_x1_sg U3124 ( .A(n2958), .X(n2960) );
  inv_x1_sg U3125 ( .A(n2958), .X(n2961) );
  inv_x1_sg U3126 ( .A(n2958), .X(n2962) );
  inv_x1_sg U3127 ( .A(n3131), .X(n2963) );
  inv_x1_sg U3128 ( .A(n2756), .X(n2964) );
  inv_x1_sg U3129 ( .A(n2963), .X(n2965) );
  inv_x1_sg U3130 ( .A(n2963), .X(n2966) );
  inv_x1_sg U3131 ( .A(n2963), .X(n2967) );
  inv_x1_sg U3132 ( .A(n2860), .X(n2969) );
  inv_x1_sg U3133 ( .A(n2860), .X(n2970) );
  inv_x1_sg U3134 ( .A(n2860), .X(n2971) );
  inv_x1_sg U3135 ( .A(n2968), .X(n2972) );
  nand_x1_sg U3136 ( .A(n2956), .B(n2824), .X(n2973) );
  inv_x1_sg U3137 ( .A(n2973), .X(n2974) );
  inv_x1_sg U3138 ( .A(n2974), .X(n2975) );
  inv_x1_sg U3139 ( .A(n2974), .X(n2976) );
  inv_x1_sg U3140 ( .A(n2974), .X(n2977) );
  inv_x1_sg U3141 ( .A(n2974), .X(n2978) );
  inv_x1_sg U3142 ( .A(n2845), .X(n2979) );
  inv_x1_sg U3143 ( .A(n1748), .X(n2980) );
  inv_x1_sg U3144 ( .A(n2980), .X(n2981) );
  inv_x1_sg U3145 ( .A(n2980), .X(n2982) );
  inv_x1_sg U3146 ( .A(n2980), .X(n2983) );
  inv_x1_sg U3147 ( .A(n2862), .X(n2984) );
  inv_x1_sg U3148 ( .A(n3250), .X(n2985) );
  inv_x1_sg U3149 ( .A(n2985), .X(n2986) );
  inv_x1_sg U3150 ( .A(n2985), .X(n2987) );
  inv_x1_sg U3151 ( .A(n2985), .X(n2988) );
  inv_x1_sg U3152 ( .A(n2864), .X(n2989) );
  inv_x1_sg U3153 ( .A(n3251), .X(n2990) );
  inv_x1_sg U3154 ( .A(n2990), .X(n2991) );
  inv_x1_sg U3155 ( .A(n2990), .X(n2992) );
  inv_x1_sg U3156 ( .A(n2990), .X(n2993) );
  inv_x1_sg U3157 ( .A(n2866), .X(n2994) );
  inv_x1_sg U3158 ( .A(n2897), .X(n2995) );
  inv_x1_sg U3159 ( .A(n2937), .X(n2996) );
  inv_x1_sg U3160 ( .A(n2899), .X(n2997) );
  inv_x1_sg U3161 ( .A(n2997), .X(n2998) );
  inv_x1_sg U3162 ( .A(n2997), .X(n2999) );
  inv_x1_sg U3163 ( .A(n2997), .X(n3000) );
  inv_x1_sg U3164 ( .A(n2897), .X(n3001) );
  inv_x1_sg U3165 ( .A(n3098), .X(n3002) );
  inv_x1_sg U3166 ( .A(n3002), .X(n3003) );
  inv_x1_sg U3167 ( .A(n3002), .X(n3004) );
  inv_x1_sg U3168 ( .A(n3002), .X(n3005) );
  inv_x1_sg U3169 ( .A(n2937), .X(n3006) );
  inv_x1_sg U3170 ( .A(n2843), .X(n3007) );
  inv_x1_sg U3171 ( .A(n3007), .X(n3008) );
  inv_x1_sg U3172 ( .A(n3007), .X(n3009) );
  inv_x1_sg U3173 ( .A(n3007), .X(n3010) );
  inv_x1_sg U3174 ( .A(n2847), .X(n3011) );
  inv_x1_sg U3175 ( .A(n1117), .X(n3012) );
  inv_x1_sg U3176 ( .A(n3012), .X(n3013) );
  inv_x1_sg U3177 ( .A(n3012), .X(n3014) );
  inv_x1_sg U3178 ( .A(n3012), .X(n3015) );
  inv_x1_sg U3179 ( .A(n2776), .X(n3016) );
  inv_x1_sg U3180 ( .A(n3016), .X(n3017) );
  inv_x1_sg U3181 ( .A(n2873), .X(n3018) );
  inv_x1_sg U3182 ( .A(n3016), .X(n3019) );
  inv_x1_sg U3183 ( .A(n3016), .X(n3020) );
  inv_x1_sg U3184 ( .A(n2637), .X(n3021) );
  inv_x1_sg U3185 ( .A(n3021), .X(n3022) );
  inv_x1_sg U3186 ( .A(n2875), .X(n3023) );
  inv_x1_sg U3187 ( .A(n3021), .X(n3024) );
  inv_x1_sg U3188 ( .A(n3021), .X(n3025) );
  inv_x1_sg U3189 ( .A(n2767), .X(n3026) );
  inv_x1_sg U3190 ( .A(n3026), .X(n3027) );
  inv_x1_sg U3191 ( .A(n2877), .X(n3028) );
  inv_x1_sg U3192 ( .A(n3026), .X(n3029) );
  inv_x1_sg U3193 ( .A(n3026), .X(n3030) );
  inv_x1_sg U3194 ( .A(n2775), .X(n3031) );
  inv_x1_sg U3195 ( .A(n3031), .X(n3032) );
  inv_x1_sg U3196 ( .A(n2879), .X(n3033) );
  inv_x1_sg U3197 ( .A(n3031), .X(n3034) );
  inv_x1_sg U3198 ( .A(n3031), .X(n3035) );
  inv_x1_sg U3199 ( .A(n2766), .X(n3036) );
  inv_x1_sg U3200 ( .A(n3036), .X(n3037) );
  inv_x1_sg U3201 ( .A(n2881), .X(n3038) );
  inv_x1_sg U3202 ( .A(n3036), .X(n3039) );
  inv_x1_sg U3203 ( .A(n3036), .X(n3040) );
  inv_x1_sg U3204 ( .A(n2636), .X(n3041) );
  inv_x1_sg U3205 ( .A(n3041), .X(n3042) );
  inv_x1_sg U3206 ( .A(n2883), .X(n3043) );
  inv_x1_sg U3207 ( .A(n3041), .X(n3044) );
  inv_x1_sg U3208 ( .A(n3041), .X(n3045) );
  inv_x1_sg U3209 ( .A(n3128), .X(n3046) );
  inv_x1_sg U3210 ( .A(n3046), .X(n3047) );
  inv_x1_sg U3211 ( .A(n3046), .X(n3048) );
  inv_x1_sg U3212 ( .A(n3046), .X(n3049) );
  inv_x1_sg U3213 ( .A(n3046), .X(n3050) );
  inv_x1_sg U3214 ( .A(n3132), .X(n3051) );
  inv_x1_sg U3215 ( .A(n2631), .X(n3052) );
  inv_x1_sg U3216 ( .A(n3051), .X(n3053) );
  inv_x1_sg U3217 ( .A(n3051), .X(n3054) );
  inv_x1_sg U3218 ( .A(n3051), .X(n3055) );
  inv_x1_sg U3219 ( .A(n3060), .X(n3056) );
  inv_x1_sg U3220 ( .A(n3752), .X(n3057) );
  inv_x1_sg U3221 ( .A(n3060), .X(n3058) );
  inv_x1_sg U3222 ( .A(n3752), .X(n3059) );
  inv_x1_sg U3223 ( .A(n2770), .X(n3060) );
  inv_x1_sg U3224 ( .A(n3060), .X(n3061) );
  inv_x1_sg U3225 ( .A(n3060), .X(n3062) );
  inv_x1_sg U3226 ( .A(n1965), .X(n3063) );
  inv_x1_sg U3227 ( .A(n2912), .X(n3064) );
  inv_x1_sg U3228 ( .A(n2912), .X(n3065) );
  inv_x1_sg U3229 ( .A(n3063), .X(n3066) );
  inv_x1_sg U3230 ( .A(n1301), .X(n3067) );
  inv_x1_sg U3231 ( .A(n2915), .X(n3068) );
  inv_x1_sg U3232 ( .A(n2915), .X(n3069) );
  inv_x1_sg U3233 ( .A(n3067), .X(n3070) );
  inv_x1_sg U3234 ( .A(n1684), .X(n3071) );
  inv_x1_sg U3235 ( .A(n2918), .X(n3072) );
  inv_x1_sg U3236 ( .A(n2918), .X(n3073) );
  inv_x1_sg U3237 ( .A(n3071), .X(n3074) );
  inv_x1_sg U3238 ( .A(n3254), .X(n3075) );
  inv_x1_sg U3239 ( .A(n3075), .X(n3076) );
  inv_x1_sg U3240 ( .A(n2925), .X(n3077) );
  inv_x1_sg U3241 ( .A(n2925), .X(n3078) );
  inv_x1_sg U3242 ( .A(n3075), .X(n3079) );
  inv_x1_sg U3243 ( .A(n1870), .X(n3080) );
  inv_x1_sg U3244 ( .A(n3080), .X(n3081) );
  inv_x1_sg U3245 ( .A(n2928), .X(n3082) );
  inv_x1_sg U3246 ( .A(n2928), .X(n3083) );
  inv_x1_sg U3247 ( .A(n3080), .X(n3084) );
  inv_x1_sg U3248 ( .A(n1207), .X(n3085) );
  inv_x1_sg U3249 ( .A(n3085), .X(n3086) );
  inv_x1_sg U3250 ( .A(n2931), .X(n3087) );
  inv_x1_sg U3251 ( .A(n2931), .X(n3088) );
  inv_x1_sg U3252 ( .A(n3085), .X(n3089) );
  inv_x1_sg U3253 ( .A(n1308), .X(n3090) );
  inv_x1_sg U3254 ( .A(n2934), .X(n3091) );
  inv_x1_sg U3255 ( .A(n2934), .X(n3092) );
  inv_x1_sg U3256 ( .A(n2894), .X(n3093) );
  inv_x1_sg U3257 ( .A(n2467), .X(n3094) );
  inv_x1_sg U3258 ( .A(n2937), .X(n3095) );
  inv_x1_sg U3259 ( .A(n2897), .X(n3096) );
  inv_x1_sg U3260 ( .A(n3094), .X(n3097) );
  inv_x1_sg U3261 ( .A(n3094), .X(n3098) );
  nor_x1_sg U3262 ( .A(n2463), .B(n3148), .X(n3099) );
  inv_x1_sg U3263 ( .A(n3099), .X(n3100) );
  inv_x1_sg U3264 ( .A(n2923), .X(n3101) );
  inv_x1_sg U3265 ( .A(n3100), .X(n3102) );
  inv_x1_sg U3266 ( .A(n3100), .X(n3103) );
  inv_x1_sg U3267 ( .A(n3100), .X(n3104) );
  inv_x1_sg U3268 ( .A(n3099), .X(n3105) );
  inv_x1_sg U3269 ( .A(n2924), .X(n3106) );
  inv_x1_sg U3270 ( .A(n3105), .X(n3107) );
  inv_x1_sg U3271 ( .A(n2924), .X(n3108) );
  inv_x1_sg U3272 ( .A(n3105), .X(n3109) );
  inv_x1_sg U3273 ( .A(n2468), .X(n3110) );
  inv_x1_sg U3274 ( .A(n3110), .X(n3111) );
  inv_x1_sg U3275 ( .A(n2924), .X(n3112) );
  inv_x1_sg U3276 ( .A(n3105), .X(n3113) );
  inv_x1_sg U3277 ( .A(n3110), .X(n3114) );
  inv_x2_sg U3278 ( .A(n3133), .X(n3115) );
  inv_x16_sg U3279 ( .A(n3166), .X(n3134) );
  nor_x1_sg U3280 ( .A(n2627), .B(reset), .X(n2456) );
  nor_x1_sg U3281 ( .A(n2819), .B(n2957), .X(n2770) );
  nor_x16_sg U3282 ( .A(mode[0]), .B(mode[1]), .X(n3133) );
  inv_x1_sg U3283 ( .A(om_min[19]), .X(n3116) );
  inv_x1_sg U3284 ( .A(om_min[17]), .X(n3117) );
  inv_x1_sg U3285 ( .A(om_min[5]), .X(n3118) );
  inv_x1_sg U3286 ( .A(om_max[19]), .X(n3119) );
  inv_x1_sg U3287 ( .A(om_max[15]), .X(n3120) );
  inv_x1_sg U3288 ( .A(om_max[11]), .X(n3121) );
  inv_x1_sg U3289 ( .A(\max_pooling_0/n640 ), .X(n3122) );
  inv_x1_sg U3290 ( .A(om_max[9]), .X(n3123) );
  inv_x1_sg U3291 ( .A(om_max[7]), .X(n3124) );
  inv_x1_sg U3292 ( .A(om_max[3]), .X(n3125) );
  inv_x1_sg U3293 ( .A(om_max[2]), .X(n3126) );
  inv_x1_sg U3294 ( .A(om_min[18]), .X(n3127) );
  inv_x1_sg U3295 ( .A(n2761), .X(n3128) );
  inv_x1_sg U3296 ( .A(n1308), .X(n3129) );
  inv_x1_sg U3297 ( .A(n3138), .X(n3130) );
  inv_x1_sg U3298 ( .A(n2756), .X(n3131) );
  inv_x1_sg U3299 ( .A(n2631), .X(n3132) );
  inv_x4_sg U3300 ( .A(n3138), .X(n3245) );
  nand_x16_sg U3301 ( .A(n2956), .B(n3252), .X(n2757) );
  inv_x1_sg U3302 ( .A(n1140), .X(n3135) );
  nor_x1_sg U3303 ( .A(n2819), .B(n3728), .X(n3254) );
  inv_x1_sg U3304 ( .A(n1145), .X(n3136) );
  inv_x16_sg U3305 ( .A(mode[1]), .X(n3137) );
  nand_x16_sg U3306 ( .A(mode[0]), .B(n3137), .X(n3138) );
  nand_x1_sg U3307 ( .A(n1309), .B(n1310), .X(n1307) );
  nand_x4_sg U3308 ( .A(n2824), .B(n1307), .X(n1308) );
  nand_x2_sg U3309 ( .A(n1972), .B(n1973), .X(n1971) );
  inv_x1_sg U3310 ( .A(n3133), .X(n3139) );
  nand_x1_sg U3311 ( .A(n1152), .B(n1153), .X(n3140) );
  nand_x1_sg U3312 ( .A(n1201), .B(n1202), .X(n3141) );
  nand_x1_sg U3313 ( .A(n1180), .B(n1181), .X(n3142) );
  nand_x1_sg U3314 ( .A(n1164), .B(n1165), .X(n3143) );
  nand_x1_sg U3315 ( .A(n1192), .B(n1193), .X(n3144) );
  inv_x1_sg U3316 ( .A(n1962), .X(n3145) );
  inv_x1_sg U3317 ( .A(n2461), .X(n3146) );
  inv_x1_sg U3318 ( .A(n3133), .X(n3147) );
  inv_x1_sg U3319 ( .A(n2456), .X(n3148) );
  inv_x1_sg U3320 ( .A(n1140), .X(n3149) );
  inv_x1_sg U3321 ( .A(\max_pooling_0/n643 ), .X(n3150) );
  inv_x1_sg U3322 ( .A(om_max[0]), .X(n3151) );
  inv_x1_sg U3323 ( .A(n1882), .X(n3152) );
  inv_x1_sg U3324 ( .A(om_max[5]), .X(n3153) );
  nand_x1_sg U3325 ( .A(n1160), .B(n1161), .X(n3154) );
  nand_x1_sg U3326 ( .A(n1168), .B(n1169), .X(n3155) );
  nand_x1_sg U3327 ( .A(n1172), .B(n1173), .X(n3156) );
  nand_x1_sg U3328 ( .A(n1188), .B(n1189), .X(n3157) );
  inv_x16_sg U3329 ( .A(n3133), .X(n3158) );
  nor_x16_sg U3330 ( .A(mode[0]), .B(mode[1]), .X(n3167) );
  nand_x1_sg U3331 ( .A(n1156), .B(n1157), .X(n3159) );
  nand_x1_sg U3332 ( .A(n1184), .B(n1185), .X(n3160) );
  nand_x1_sg U3333 ( .A(n1196), .B(n1197), .X(n3161) );
  nand_x1_sg U3334 ( .A(n1118), .B(n1119), .X(n3162) );
  nand_x1_sg U3335 ( .A(n1126), .B(n1127), .X(n3163) );
  inv_x16_sg U3336 ( .A(n3167), .X(n3164) );
  nor_x16_sg U3337 ( .A(mode[0]), .B(mode[1]), .X(n3166) );
  nand_x1_sg U3338 ( .A(n1176), .B(n1177), .X(n3168) );
  nand_x1_sg U3339 ( .A(n1122), .B(n1123), .X(n3169) );
  nand_x1_sg U3340 ( .A(n1130), .B(n1131), .X(n3170) );
  nand_x1_sg U3341 ( .A(n1134), .B(n1135), .X(n3171) );
  nand_x1_sg U3342 ( .A(n1148), .B(n1149), .X(n3172) );
  inv_x1_sg U3343 ( .A(n3138), .X(n3244) );
  inv_x1_sg U3344 ( .A(\reg_im[3][19] ), .X(n3173) );
  inv_x1_sg U3345 ( .A(\reg_im[3][17] ), .X(n3174) );
  inv_x1_sg U3346 ( .A(\reg_im[3][15] ), .X(n3175) );
  inv_x1_sg U3347 ( .A(om_max[17]), .X(n3176) );
  inv_x1_sg U3348 ( .A(n3167), .X(n3177) );
  inv_x1_sg U3349 ( .A(n3167), .X(n3178) );
  nand_x2_sg U3350 ( .A(n1336), .B(n1337), .X(n1332) );
  nand_x2_sg U3351 ( .A(n1338), .B(n1339), .X(n1337) );
  inv_x1_sg U3352 ( .A(om_min[9]), .X(n3179) );
  inv_x1_sg U3353 ( .A(n2464), .X(n3180) );
  inv_x1_sg U3354 ( .A(\reg_im[1][12] ), .X(n3181) );
  inv_x1_sg U3355 ( .A(\reg_im[2][2] ), .X(n3182) );
  inv_x1_sg U3356 ( .A(\reg_im[2][5] ), .X(n3183) );
  inv_x1_sg U3357 ( .A(\reg_im[2][8] ), .X(n3184) );
  inv_x1_sg U3358 ( .A(\reg_im[3][1] ), .X(n3185) );
  inv_x1_sg U3359 ( .A(\reg_im[3][14] ), .X(n3186) );
  inv_x1_sg U3360 ( .A(\reg_im[1][6] ), .X(n3187) );
  inv_x1_sg U3361 ( .A(\reg_im[3][10] ), .X(n3188) );
  inv_x1_sg U3362 ( .A(\reg_im[1][9] ), .X(n3189) );
  inv_x1_sg U3363 ( .A(\reg_im[3][5] ), .X(n3190) );
  inv_x1_sg U3364 ( .A(\reg_im[3][2] ), .X(n3191) );
  inv_x1_sg U3365 ( .A(\reg_im[3][0] ), .X(n3192) );
  inv_x1_sg U3366 ( .A(\max_pooling_0/n639 ), .X(n3193) );
  inv_x1_sg U3367 ( .A(\min_pooling_0/n724 ), .X(n3194) );
  inv_x16_sg U3368 ( .A(mode[1]), .X(n3729) );
  nand_x1_sg U3369 ( .A(n3061), .B(\max_pooling_0/n325 ), .X(n2788) );
  inv_x1_sg U3370 ( .A(\max_pooling_0/N3 ), .X(n3195) );
  inv_x1_sg U3371 ( .A(n1140), .X(n3196) );
  nand_x1_sg U3372 ( .A(n1677), .B(n1678), .X(n3197) );
  nand_x4_sg U3373 ( .A(n1095), .B(n3628), .X(n1677) );
  inv_x1_sg U3374 ( .A(\reg_im[2][18] ), .X(n3198) );
  inv_x1_sg U3375 ( .A(\reg_im[2][17] ), .X(n3199) );
  inv_x1_sg U3376 ( .A(\reg_im[2][12] ), .X(n3200) );
  inv_x1_sg U3377 ( .A(\reg_im[3][12] ), .X(n3201) );
  inv_x1_sg U3378 ( .A(\reg_im[2][1] ), .X(n3202) );
  inv_x1_sg U3379 ( .A(\reg_im[2][0] ), .X(n3203) );
  inv_x1_sg U3380 ( .A(\reg_im[2][3] ), .X(n3204) );
  inv_x1_sg U3381 ( .A(\reg_im[2][4] ), .X(n3205) );
  inv_x1_sg U3382 ( .A(\reg_im[2][6] ), .X(n3206) );
  inv_x1_sg U3383 ( .A(\reg_im[2][7] ), .X(n3207) );
  inv_x1_sg U3384 ( .A(\reg_im[2][9] ), .X(n3208) );
  inv_x1_sg U3385 ( .A(\reg_im[2][10] ), .X(n3209) );
  inv_x1_sg U3386 ( .A(\reg_im[2][11] ), .X(n3210) );
  inv_x1_sg U3387 ( .A(\reg_im[2][13] ), .X(n3211) );
  inv_x1_sg U3388 ( .A(\reg_im[2][14] ), .X(n3212) );
  inv_x1_sg U3389 ( .A(\reg_im[2][15] ), .X(n3213) );
  inv_x1_sg U3390 ( .A(\reg_im[2][16] ), .X(n3214) );
  inv_x1_sg U3391 ( .A(\reg_im[2][19] ), .X(n3215) );
  inv_x1_sg U3392 ( .A(\reg_im[1][19] ), .X(n3216) );
  inv_x1_sg U3393 ( .A(\reg_im[1][17] ), .X(n3217) );
  inv_x1_sg U3394 ( .A(\reg_im[3][18] ), .X(n3218) );
  inv_x1_sg U3395 ( .A(\reg_im[1][18] ), .X(n3219) );
  inv_x1_sg U3396 ( .A(\reg_im[3][16] ), .X(n3220) );
  inv_x1_sg U3397 ( .A(\reg_im[1][16] ), .X(n3221) );
  inv_x1_sg U3398 ( .A(\reg_im[1][1] ), .X(n3222) );
  inv_x1_sg U3399 ( .A(\reg_im[1][15] ), .X(n3223) );
  inv_x1_sg U3400 ( .A(\reg_im[1][14] ), .X(n3224) );
  inv_x1_sg U3401 ( .A(\reg_im[3][13] ), .X(n3225) );
  inv_x1_sg U3402 ( .A(\reg_im[1][13] ), .X(n3226) );
  inv_x1_sg U3403 ( .A(\reg_im[3][6] ), .X(n3227) );
  inv_x1_sg U3404 ( .A(\reg_im[3][11] ), .X(n3228) );
  inv_x1_sg U3405 ( .A(\reg_im[1][11] ), .X(n3229) );
  inv_x1_sg U3406 ( .A(\reg_im[1][10] ), .X(n3230) );
  inv_x1_sg U3407 ( .A(\reg_im[3][9] ), .X(n3231) );
  inv_x1_sg U3408 ( .A(\reg_im[3][7] ), .X(n3232) );
  inv_x1_sg U3409 ( .A(\reg_im[1][7] ), .X(n3233) );
  inv_x1_sg U3410 ( .A(\reg_im[3][8] ), .X(n3234) );
  inv_x1_sg U3411 ( .A(\reg_im[1][8] ), .X(n3235) );
  inv_x1_sg U3412 ( .A(\reg_im[3][4] ), .X(n3236) );
  inv_x1_sg U3413 ( .A(\reg_im[1][4] ), .X(n3237) );
  inv_x1_sg U3414 ( .A(\reg_im[1][5] ), .X(n3238) );
  inv_x1_sg U3415 ( .A(\reg_im[3][3] ), .X(n3239) );
  inv_x1_sg U3416 ( .A(\reg_im[1][3] ), .X(n3240) );
  inv_x1_sg U3417 ( .A(\reg_im[1][2] ), .X(n3241) );
  inv_x1_sg U3418 ( .A(\reg_im[1][0] ), .X(n3242) );
  inv_x1_sg U3419 ( .A(om_min[13]), .X(n3243) );
  nor_x16_sg U3420 ( .A(mode[0]), .B(mode[1]), .X(n1140) );
  nand_x16_sg U3421 ( .A(mode[0]), .B(n3729), .X(n1145) );
  inv_x1_sg U3422 ( .A(n1385), .X(n3627) );
  nor_x1_sg U3423 ( .A(n1373), .B(n1374), .X(n1372) );
  nand_x1_sg U3424 ( .A(n1375), .B(n1376), .X(n1374) );
  nand_x1_sg U3425 ( .A(n2029), .B(n2030), .X(n2028) );
  nand_x1_sg U3426 ( .A(n1367), .B(n1368), .X(n1366) );
  nand_x1_sg U3427 ( .A(n1358), .B(n1359), .X(n1357) );
  inv_x1_sg U3428 ( .A(n1458), .X(n3671) );
  nand_x2_sg U3429 ( .A(n2018), .B(n2019), .X(n2014) );
  inv_x1_sg U3430 ( .A(n2115), .X(n3687) );
  nand_x1_sg U3431 ( .A(n1352), .B(n1353), .X(n1351) );
  nand_x1_sg U3432 ( .A(n1356), .B(n1357), .X(n1352) );
  inv_x1_sg U3433 ( .A(n1345), .X(n3249) );
  nand_x1_sg U3434 ( .A(n2134), .B(n2116), .X(n2112) );
  nor_x1_sg U3435 ( .A(n2005), .B(n2006), .X(n2004) );
  nand_x1_sg U3436 ( .A(n2008), .B(n2009), .X(n2005) );
  nand_x1_sg U3437 ( .A(n1332), .B(n1333), .X(n1331) );
  nand_x4_sg U3438 ( .A(n1751), .B(n1752), .X(n1743) );
  nand_x4_sg U3439 ( .A(n1862), .B(n1863), .X(n1861) );
  nor_x1_sg U3440 ( .A(n1739), .B(n1740), .X(n1661) );
  nor_x1_sg U3441 ( .A(n1741), .B(n1096), .X(n1740) );
  nand_x1_sg U3442 ( .A(n1311), .B(n1312), .X(n1310) );
  nand_x1_sg U3443 ( .A(n1313), .B(n1314), .X(n1311) );
  nor_x1_sg U3444 ( .A(n1691), .B(n1692), .X(n1688) );
  nor_x1_sg U3445 ( .A(n1693), .B(n1112), .X(n1692) );
  nor_x1_sg U3446 ( .A(n1859), .B(n1860), .X(n1689) );
  nand_x1_sg U3447 ( .A(n1524), .B(n1525), .X(n1522) );
  nand_x1_sg U3448 ( .A(n1533), .B(n1534), .X(n1531) );
  nand_x1_sg U3449 ( .A(n1542), .B(n1543), .X(n1540) );
  nand_x1_sg U3450 ( .A(n1551), .B(n1552), .X(n1549) );
  nand_x1_sg U3451 ( .A(n1560), .B(n1561), .X(n1558) );
  nand_x1_sg U3452 ( .A(n1569), .B(n1570), .X(n1567) );
  nand_x1_sg U3453 ( .A(n1578), .B(n1579), .X(n1576) );
  nand_x1_sg U3454 ( .A(n1587), .B(n1588), .X(n1585) );
  nand_x1_sg U3455 ( .A(n1596), .B(n1597), .X(n1594) );
  nand_x1_sg U3456 ( .A(n1605), .B(n1606), .X(n1603) );
  nand_x1_sg U3457 ( .A(n1614), .B(n1615), .X(n1612) );
  nand_x1_sg U3458 ( .A(n1623), .B(n1624), .X(n1621) );
  nand_x1_sg U3459 ( .A(n1632), .B(n1633), .X(n1630) );
  nand_x1_sg U3460 ( .A(n1641), .B(n1642), .X(n1639) );
  nand_x1_sg U3461 ( .A(n1650), .B(n1651), .X(n1648) );
  nand_x1_sg U3462 ( .A(n1659), .B(n1660), .X(n1657) );
  nand_x1_sg U3463 ( .A(n1668), .B(n1669), .X(n1666) );
  nand_x4_sg U3464 ( .A(n1744), .B(n1745), .X(n1683) );
  nand_x2_sg U3465 ( .A(n1419), .B(n1420), .X(n1228) );
  nand_x2_sg U3466 ( .A(n1473), .B(n1474), .X(n1248) );
  nand_x2_sg U3467 ( .A(n1486), .B(n1487), .X(n1268) );
  nand_x2_sg U3468 ( .A(n1500), .B(n1501), .X(n1283) );
  nand_x2_sg U3469 ( .A(n1506), .B(n1507), .X(n1288) );
  nand_x2_sg U3470 ( .A(n1393), .B(n1394), .X(n1298) );
  nand_x1_sg U3471 ( .A(n3726), .B(n1687), .X(n1685) );
  nand_x1_sg U3472 ( .A(n1520), .B(n3722), .X(n1518) );
  nand_x1_sg U3473 ( .A(n1529), .B(n3716), .X(n1527) );
  nand_x1_sg U3474 ( .A(n1538), .B(n3711), .X(n1536) );
  nand_x1_sg U3475 ( .A(n1547), .B(n3705), .X(n1545) );
  nand_x1_sg U3476 ( .A(n1556), .B(n3700), .X(n1554) );
  nand_x1_sg U3477 ( .A(n1565), .B(n3694), .X(n1563) );
  nand_x1_sg U3478 ( .A(n1574), .B(n3689), .X(n1572) );
  nand_x1_sg U3479 ( .A(n1583), .B(n3683), .X(n1581) );
  nand_x1_sg U3480 ( .A(n1592), .B(n3678), .X(n1590) );
  nand_x1_sg U3481 ( .A(n1601), .B(n3672), .X(n1599) );
  nand_x1_sg U3482 ( .A(n1610), .B(n3666), .X(n1608) );
  nand_x1_sg U3483 ( .A(n1619), .B(n3660), .X(n1617) );
  nand_x1_sg U3484 ( .A(n1628), .B(n3655), .X(n1626) );
  nand_x1_sg U3485 ( .A(n1637), .B(n3649), .X(n1635) );
  nand_x1_sg U3486 ( .A(n1646), .B(n3644), .X(n1644) );
  nand_x1_sg U3487 ( .A(n1655), .B(n3639), .X(n1653) );
  nand_x1_sg U3488 ( .A(n1664), .B(n1665), .X(n1662) );
  inv_x1_sg U3489 ( .A(n1676), .X(n3629) );
  nor_x1_sg U3490 ( .A(n1681), .B(n1682), .X(n1679) );
  nand_x2_sg U3491 ( .A(n2038), .B(n2039), .X(n1872) );
  nand_x2_sg U3492 ( .A(n2060), .B(n2061), .X(n1877) );
  nand_x2_sg U3493 ( .A(n2073), .B(n2074), .X(n1882) );
  nand_x2_sg U3494 ( .A(n2086), .B(n2087), .X(n1897) );
  nand_x2_sg U3495 ( .A(n2135), .B(n2136), .X(n1912) );
  nand_x2_sg U3496 ( .A(n2141), .B(n2142), .X(n1917) );
  nand_x2_sg U3497 ( .A(n2154), .B(n2155), .X(n1937) );
  nand_x2_sg U3498 ( .A(n2048), .B(n2049), .X(n1962) );
  nand_x1_sg U3499 ( .A(n1969), .B(n1970), .X(\max_pooling_0/n228 ) );
  nand_x1_sg U3500 ( .A(n1893), .B(n1894), .X(\max_pooling_0/n292 ) );
  nand_x1_sg U3501 ( .A(n1898), .B(n1899), .X(\max_pooling_0/n288 ) );
  nand_x1_sg U3502 ( .A(n1903), .B(n1904), .X(\max_pooling_0/n284 ) );
  nand_x1_sg U3503 ( .A(n1908), .B(n1909), .X(\max_pooling_0/n280 ) );
  nand_x1_sg U3504 ( .A(n1923), .B(n1924), .X(\max_pooling_0/n268 ) );
  nand_x1_sg U3505 ( .A(n1948), .B(n1949), .X(\max_pooling_0/n248 ) );
  nand_x1_sg U3506 ( .A(n1953), .B(n1954), .X(\max_pooling_0/n244 ) );
  nand_x1_sg U3507 ( .A(n1142), .B(n1143), .X(n418) );
  nand_x1_sg U3508 ( .A(n1138), .B(n1139), .X(n422) );
  nand_x2_sg U3509 ( .A(n2757), .B(n2758), .X(n2756) );
  nand_x2_sg U3510 ( .A(n3252), .B(n2841), .X(n2758) );
  inv_x1_sg U3511 ( .A(\mean_pooling_0/N5 ), .X(n3246) );
  inv_x1_sg U3512 ( .A(\max_pooling_0/N4 ), .X(n3247) );
  inv_x1_sg U3513 ( .A(\min_pooling_0/N3 ), .X(n3248) );
  nand_x1_sg U3514 ( .A(n1432), .B(n1436), .X(n1345) );
  nand_x2_sg U3515 ( .A(n1978), .B(n1979), .X(n1977) );
  nand_x2_sg U3516 ( .A(n1980), .B(n1981), .X(n1979) );
  nand_x1_sg U3517 ( .A(n3753), .B(n3246), .X(n1748) );
  nand_x1_sg U3518 ( .A(n3248), .B(n3603), .X(n3250) );
  nand_x1_sg U3519 ( .A(n3195), .B(n3247), .X(n3251) );
  inv_x1_sg U3520 ( .A(n2007), .X(n3698) );
  nand_x2_sg U3521 ( .A(n1974), .B(n1975), .X(n1973) );
  nand_x1_sg U3522 ( .A(n3249), .B(n1344), .X(n1343) );
  inv_x1_sg U3523 ( .A(n1738), .X(n3640) );
  inv_x1_sg U3524 ( .A(n1735), .X(n3645) );
  inv_x1_sg U3525 ( .A(n1732), .X(n3650) );
  inv_x1_sg U3526 ( .A(n1729), .X(n3656) );
  inv_x1_sg U3527 ( .A(n1726), .X(n3661) );
  inv_x1_sg U3528 ( .A(n1723), .X(n3667) );
  inv_x1_sg U3529 ( .A(n1720), .X(n3673) );
  inv_x1_sg U3530 ( .A(n1717), .X(n3679) );
  inv_x1_sg U3531 ( .A(n1714), .X(n3684) );
  inv_x1_sg U3532 ( .A(n1711), .X(n3690) );
  inv_x1_sg U3533 ( .A(n1708), .X(n3695) );
  inv_x1_sg U3534 ( .A(n1705), .X(n3701) );
  inv_x1_sg U3535 ( .A(n1702), .X(n3706) );
  inv_x1_sg U3536 ( .A(n1699), .X(n3712) );
  inv_x1_sg U3537 ( .A(n1696), .X(n3717) );
  nand_x1_sg U3538 ( .A(n1369), .B(n3634), .X(n1368) );
  inv_x1_sg U3539 ( .A(n1521), .X(n3722) );
  inv_x1_sg U3540 ( .A(n1656), .X(n3639) );
  inv_x1_sg U3541 ( .A(n1530), .X(n3716) );
  inv_x1_sg U3542 ( .A(n1539), .X(n3711) );
  inv_x1_sg U3543 ( .A(n1548), .X(n3705) );
  inv_x1_sg U3544 ( .A(n1557), .X(n3700) );
  inv_x1_sg U3545 ( .A(n1566), .X(n3694) );
  inv_x1_sg U3546 ( .A(n1575), .X(n3689) );
  inv_x1_sg U3547 ( .A(n1584), .X(n3683) );
  inv_x1_sg U3548 ( .A(n1593), .X(n3678) );
  inv_x1_sg U3549 ( .A(n1602), .X(n3672) );
  inv_x1_sg U3550 ( .A(n1611), .X(n3666) );
  inv_x1_sg U3551 ( .A(n1620), .X(n3660) );
  inv_x1_sg U3552 ( .A(n1629), .X(n3655) );
  inv_x1_sg U3553 ( .A(n1638), .X(n3649) );
  inv_x1_sg U3554 ( .A(n1647), .X(n3644) );
  nand_x1_sg U3555 ( .A(n2971), .B(n1686), .X(\mean_pooling_0/n163 ) );
  nand_x1_sg U3556 ( .A(n2970), .B(n1519), .X(\mean_pooling_0/n243 ) );
  nand_x1_sg U3557 ( .A(n2970), .B(n1528), .X(\mean_pooling_0/n239 ) );
  nand_x1_sg U3558 ( .A(n2971), .B(n1546), .X(\mean_pooling_0/n231 ) );
  nand_x1_sg U3559 ( .A(n2969), .B(n1537), .X(\mean_pooling_0/n235 ) );
  inv_x1_sg U3560 ( .A(n1690), .X(n3726) );
  nand_x2_sg U3561 ( .A(n1315), .B(n1316), .X(n1314) );
  nand_x2_sg U3562 ( .A(n2020), .B(n2021), .X(n2019) );
  inv_x1_sg U3563 ( .A(n2047), .X(n3633) );
  nand_x1_sg U3564 ( .A(n1209), .B(n1210), .X(\min_pooling_0/n389 ) );
  nand_x1_sg U3565 ( .A(n1214), .B(n1215), .X(\min_pooling_0/n385 ) );
  nand_x1_sg U3566 ( .A(n1224), .B(n1225), .X(\min_pooling_0/n377 ) );
  nand_x1_sg U3567 ( .A(n1249), .B(n1250), .X(\min_pooling_0/n357 ) );
  nand_x1_sg U3568 ( .A(n1254), .B(n1255), .X(\min_pooling_0/n353 ) );
  nand_x1_sg U3569 ( .A(n1269), .B(n1270), .X(\min_pooling_0/n341 ) );
  nand_x1_sg U3570 ( .A(n1274), .B(n1275), .X(\min_pooling_0/n337 ) );
  nand_x1_sg U3571 ( .A(n1279), .B(n1280), .X(\min_pooling_0/n333 ) );
  nand_x1_sg U3572 ( .A(n1284), .B(n1285), .X(\min_pooling_0/n329 ) );
  nand_x1_sg U3573 ( .A(n1294), .B(n1295), .X(\min_pooling_0/n321 ) );
  nand_x1_sg U3574 ( .A(n1299), .B(n1300), .X(\min_pooling_0/n317 ) );
  nand_x1_sg U3575 ( .A(n1305), .B(n1306), .X(\min_pooling_0/n309 ) );
  nand_x1_sg U3576 ( .A(n1219), .B(n1220), .X(\min_pooling_0/n381 ) );
  nand_x1_sg U3577 ( .A(n1259), .B(n1260), .X(\min_pooling_0/n349 ) );
  nand_x1_sg U3578 ( .A(n1264), .B(n1265), .X(\min_pooling_0/n345 ) );
  nand_x1_sg U3579 ( .A(n1928), .B(n1929), .X(\max_pooling_0/n264 ) );
  nand_x1_sg U3580 ( .A(n1933), .B(n1934), .X(\max_pooling_0/n260 ) );
  nand_x1_sg U3581 ( .A(n1943), .B(n1944), .X(\max_pooling_0/n252 ) );
  nand_x1_sg U3582 ( .A(n1883), .B(n1884), .X(\max_pooling_0/n300 ) );
  nand_x1_sg U3583 ( .A(n1873), .B(n1874), .X(\max_pooling_0/n308 ) );
  nand_x1_sg U3584 ( .A(n1878), .B(n1879), .X(\max_pooling_0/n304 ) );
  nand_x1_sg U3585 ( .A(n1888), .B(n1889), .X(\max_pooling_0/n296 ) );
  nand_x1_sg U3586 ( .A(n1913), .B(n1914), .X(\max_pooling_0/n276 ) );
  nand_x1_sg U3587 ( .A(n1918), .B(n1919), .X(\max_pooling_0/n272 ) );
  nand_x1_sg U3588 ( .A(n1938), .B(n1939), .X(\max_pooling_0/n256 ) );
  nand_x1_sg U3589 ( .A(n1958), .B(n1959), .X(\max_pooling_0/n240 ) );
  nand_x1_sg U3590 ( .A(n1963), .B(n1964), .X(\max_pooling_0/n236 ) );
  nand_x1_sg U3591 ( .A(n1229), .B(n1230), .X(\min_pooling_0/n373 ) );
  nand_x1_sg U3592 ( .A(n1234), .B(n1235), .X(\min_pooling_0/n369 ) );
  nand_x1_sg U3593 ( .A(n1239), .B(n1240), .X(\min_pooling_0/n365 ) );
  nand_x1_sg U3594 ( .A(n1244), .B(n1245), .X(\min_pooling_0/n361 ) );
  nand_x1_sg U3595 ( .A(n2722), .B(n2723), .X(\mean_pooling_0/n264 ) );
  nand_x1_sg U3596 ( .A(n2724), .B(n2725), .X(\mean_pooling_0/n263 ) );
  nand_x1_sg U3597 ( .A(n2726), .B(n2727), .X(\mean_pooling_0/n262 ) );
  nand_x1_sg U3598 ( .A(n2728), .B(n2729), .X(\mean_pooling_0/n261 ) );
  nand_x1_sg U3599 ( .A(n2730), .B(n2731), .X(\mean_pooling_0/n260 ) );
  nand_x1_sg U3600 ( .A(n2732), .B(n2733), .X(\mean_pooling_0/n259 ) );
  nand_x1_sg U3601 ( .A(n2734), .B(n2735), .X(\mean_pooling_0/n258 ) );
  nand_x1_sg U3602 ( .A(n2736), .B(n2737), .X(\mean_pooling_0/n257 ) );
  nand_x1_sg U3603 ( .A(n2738), .B(n2739), .X(\mean_pooling_0/n256 ) );
  nand_x1_sg U3604 ( .A(n2740), .B(n2741), .X(\mean_pooling_0/n255 ) );
  nand_x1_sg U3605 ( .A(n2742), .B(n2743), .X(\mean_pooling_0/n254 ) );
  nand_x1_sg U3606 ( .A(n2744), .B(n2745), .X(\mean_pooling_0/n253 ) );
  nand_x1_sg U3607 ( .A(n2746), .B(n2747), .X(\mean_pooling_0/n252 ) );
  nand_x1_sg U3608 ( .A(n2748), .B(n2749), .X(\mean_pooling_0/n251 ) );
  nand_x1_sg U3609 ( .A(n2750), .B(n2751), .X(\mean_pooling_0/n250 ) );
  nand_x1_sg U3610 ( .A(n2752), .B(n2753), .X(\mean_pooling_0/n249 ) );
  nand_x1_sg U3611 ( .A(n2754), .B(n2755), .X(\mean_pooling_0/n248 ) );
  nand_x1_sg U3612 ( .A(n2719), .B(n2720), .X(\mean_pooling_0/n265 ) );
  nand_x1_sg U3613 ( .A(n2960), .B(n2822), .X(n2720) );
  nand_x1_sg U3614 ( .A(n2511), .B(n2512), .X(n502) );
  nand_x1_sg U3615 ( .A(n2513), .B(n2514), .X(n501) );
  nand_x1_sg U3616 ( .A(n2583), .B(n2584), .X(n466) );
  nand_x1_sg U3617 ( .A(n2585), .B(n2586), .X(n465) );
  nand_x1_sg U3618 ( .A(n2587), .B(n2588), .X(n464) );
  nand_x1_sg U3619 ( .A(n2589), .B(n2590), .X(n463) );
  nand_x1_sg U3620 ( .A(n2465), .B(n2466), .X(n524) );
  nand_x1_sg U3621 ( .A(n2469), .B(n2470), .X(n523) );
  nand_x1_sg U3622 ( .A(n2471), .B(n2472), .X(n522) );
  nand_x1_sg U3623 ( .A(n2473), .B(n2474), .X(n521) );
  nand_x1_sg U3624 ( .A(n2475), .B(n2476), .X(n520) );
  nand_x1_sg U3625 ( .A(n2477), .B(n2478), .X(n519) );
  nand_x1_sg U3626 ( .A(n2479), .B(n2480), .X(n518) );
  nand_x1_sg U3627 ( .A(n2481), .B(n2482), .X(n517) );
  nand_x1_sg U3628 ( .A(n2483), .B(n2484), .X(n516) );
  nand_x1_sg U3629 ( .A(n2485), .B(n2486), .X(n515) );
  nand_x1_sg U3630 ( .A(n2487), .B(n2488), .X(n514) );
  nand_x1_sg U3631 ( .A(n2489), .B(n2490), .X(n513) );
  nand_x1_sg U3632 ( .A(n2491), .B(n2492), .X(n512) );
  nand_x1_sg U3633 ( .A(n2493), .B(n2494), .X(n511) );
  nand_x1_sg U3634 ( .A(n2495), .B(n2496), .X(n510) );
  nand_x1_sg U3635 ( .A(n2497), .B(n2498), .X(n509) );
  nand_x1_sg U3636 ( .A(n2499), .B(n2500), .X(n508) );
  nand_x1_sg U3637 ( .A(n2501), .B(n2502), .X(n507) );
  nand_x1_sg U3638 ( .A(n2503), .B(n2504), .X(n506) );
  nand_x1_sg U3639 ( .A(n2505), .B(n2506), .X(n505) );
  nand_x1_sg U3640 ( .A(n2507), .B(n2508), .X(n504) );
  nand_x1_sg U3641 ( .A(n2509), .B(n2510), .X(n503) );
  nand_x1_sg U3642 ( .A(n2515), .B(n2516), .X(n500) );
  nand_x1_sg U3643 ( .A(n2537), .B(n2538), .X(n489) );
  nand_x1_sg U3644 ( .A(n2539), .B(n2540), .X(n488) );
  nand_x1_sg U3645 ( .A(n2541), .B(n2542), .X(n487) );
  nand_x1_sg U3646 ( .A(n2543), .B(n2544), .X(n486) );
  nand_x1_sg U3647 ( .A(n2545), .B(n2546), .X(n485) );
  nand_x1_sg U3648 ( .A(n2547), .B(n2548), .X(n484) );
  nand_x1_sg U3649 ( .A(n2549), .B(n2550), .X(n483) );
  nand_x1_sg U3650 ( .A(n2551), .B(n2552), .X(n482) );
  nand_x1_sg U3651 ( .A(n2553), .B(n2554), .X(n481) );
  nand_x1_sg U3652 ( .A(n2555), .B(n2556), .X(n480) );
  nand_x1_sg U3653 ( .A(n2557), .B(n2558), .X(n479) );
  nand_x1_sg U3654 ( .A(n2559), .B(n2560), .X(n478) );
  nand_x1_sg U3655 ( .A(n2561), .B(n2562), .X(n477) );
  nand_x1_sg U3656 ( .A(n2563), .B(n2564), .X(n476) );
  nand_x1_sg U3657 ( .A(n2565), .B(n2566), .X(n475) );
  nand_x1_sg U3658 ( .A(n2567), .B(n2568), .X(n474) );
  nand_x1_sg U3659 ( .A(n2569), .B(n2570), .X(n473) );
  nand_x1_sg U3660 ( .A(n2571), .B(n2572), .X(n472) );
  nand_x1_sg U3661 ( .A(n2573), .B(n2574), .X(n471) );
  nand_x1_sg U3662 ( .A(n2575), .B(n2576), .X(n470) );
  nand_x1_sg U3663 ( .A(n2577), .B(n2578), .X(n469) );
  nand_x1_sg U3664 ( .A(n2579), .B(n2580), .X(n468) );
  nand_x1_sg U3665 ( .A(n2581), .B(n2582), .X(n467) );
  nand_x1_sg U3666 ( .A(n2591), .B(n2592), .X(n462) );
  nand_x1_sg U3667 ( .A(n2593), .B(n2594), .X(n461) );
  nand_x1_sg U3668 ( .A(n2595), .B(n2596), .X(n460) );
  nand_x1_sg U3669 ( .A(n2597), .B(n2598), .X(n459) );
  nand_x1_sg U3670 ( .A(n2599), .B(n2600), .X(n458) );
  nand_x1_sg U3671 ( .A(n2601), .B(n2602), .X(n457) );
  nand_x1_sg U3672 ( .A(n2603), .B(n2604), .X(n456) );
  nand_x1_sg U3673 ( .A(n2605), .B(n2606), .X(n455) );
  nand_x1_sg U3674 ( .A(n2607), .B(n2608), .X(n454) );
  nand_x1_sg U3675 ( .A(n2609), .B(n2610), .X(n453) );
  nand_x1_sg U3676 ( .A(n2611), .B(n2612), .X(n452) );
  nand_x1_sg U3677 ( .A(n2613), .B(n2614), .X(n451) );
  nand_x1_sg U3678 ( .A(n2615), .B(n2616), .X(n450) );
  nand_x1_sg U3679 ( .A(n2617), .B(n2618), .X(n449) );
  nand_x1_sg U3680 ( .A(n2619), .B(n2620), .X(n448) );
  nand_x1_sg U3681 ( .A(n2621), .B(n2622), .X(n447) );
  nand_x1_sg U3682 ( .A(n2623), .B(n2624), .X(n446) );
  nand_x1_sg U3683 ( .A(n2625), .B(n2626), .X(n445) );
  nand_x1_sg U3684 ( .A(n2523), .B(n2524), .X(n496) );
  nand_x1_sg U3685 ( .A(n2525), .B(n2526), .X(n495) );
  nand_x1_sg U3686 ( .A(n2517), .B(n2518), .X(n499) );
  nand_x1_sg U3687 ( .A(n2519), .B(n2520), .X(n498) );
  nand_x1_sg U3688 ( .A(n2521), .B(n2522), .X(n497) );
  nand_x1_sg U3689 ( .A(n2527), .B(n2528), .X(n494) );
  nand_x1_sg U3690 ( .A(n2529), .B(n2530), .X(n493) );
  nand_x1_sg U3691 ( .A(n2531), .B(n2532), .X(n492) );
  nand_x1_sg U3692 ( .A(n2533), .B(n2534), .X(n491) );
  nand_x1_sg U3693 ( .A(n2535), .B(n2536), .X(n490) );
  nand_x1_sg U3694 ( .A(n2651), .B(n2652), .X(\min_pooling_0/n408 ) );
  nand_x1_sg U3695 ( .A(n2699), .B(n2700), .X(\min_pooling_0/n396 ) );
  nand_x1_sg U3696 ( .A(n2632), .B(n2633), .X(\min_pooling_0/n412 ) );
  nand_x1_sg U3697 ( .A(n2643), .B(n2644), .X(\min_pooling_0/n410 ) );
  nand_x1_sg U3698 ( .A(n2659), .B(n2660), .X(\min_pooling_0/n406 ) );
  nand_x1_sg U3699 ( .A(n2667), .B(n2668), .X(\min_pooling_0/n404 ) );
  nand_x1_sg U3700 ( .A(n2675), .B(n2676), .X(\min_pooling_0/n402 ) );
  nand_x1_sg U3701 ( .A(n2683), .B(n2684), .X(\min_pooling_0/n400 ) );
  nand_x1_sg U3702 ( .A(n2691), .B(n2692), .X(\min_pooling_0/n398 ) );
  nand_x1_sg U3703 ( .A(n2707), .B(n2708), .X(\min_pooling_0/n394 ) );
  nand_x1_sg U3704 ( .A(n2715), .B(n2716), .X(\min_pooling_0/n392 ) );
  nand_x1_sg U3705 ( .A(n2762), .B(n2763), .X(\mean_pooling_0/n246 ) );
  nand_x1_sg U3706 ( .A(n2638), .B(n2639), .X(\min_pooling_0/n411 ) );
  nand_x1_sg U3707 ( .A(n2655), .B(n2656), .X(\min_pooling_0/n407 ) );
  nand_x1_sg U3708 ( .A(n2663), .B(n2664), .X(\min_pooling_0/n405 ) );
  nand_x1_sg U3709 ( .A(n2671), .B(n2672), .X(\min_pooling_0/n403 ) );
  nand_x1_sg U3710 ( .A(n2679), .B(n2680), .X(\min_pooling_0/n401 ) );
  nand_x1_sg U3711 ( .A(n2687), .B(n2688), .X(\min_pooling_0/n399 ) );
  nand_x1_sg U3712 ( .A(n2695), .B(n2696), .X(\min_pooling_0/n397 ) );
  nand_x1_sg U3713 ( .A(n2703), .B(n2704), .X(\min_pooling_0/n395 ) );
  nand_x1_sg U3714 ( .A(n2711), .B(n2712), .X(\min_pooling_0/n393 ) );
  nand_x1_sg U3715 ( .A(n2647), .B(n2648), .X(\min_pooling_0/n409 ) );
  nand_x1_sg U3716 ( .A(n2771), .B(n2772), .X(\max_pooling_0/n351 ) );
  nand_x1_sg U3717 ( .A(n2458), .B(n2459), .X(n525) );
  nand_x1_sg U3718 ( .A(n2454), .B(n2455), .X(n526) );
  nand_x1_sg U3719 ( .A(n2811), .B(n2812), .X(\max_pooling_0/n333 ) );
  nand_x1_sg U3720 ( .A(n2813), .B(n2814), .X(\max_pooling_0/n332 ) );
  nand_x1_sg U3721 ( .A(n2777), .B(n2778), .X(\max_pooling_0/n350 ) );
  nand_x1_sg U3722 ( .A(n2785), .B(n2786), .X(\max_pooling_0/n346 ) );
  nand_x1_sg U3723 ( .A(n2789), .B(n2790), .X(\max_pooling_0/n344 ) );
  nand_x1_sg U3724 ( .A(n2791), .B(n2792), .X(\max_pooling_0/n343 ) );
  nand_x1_sg U3725 ( .A(n2801), .B(n2802), .X(\max_pooling_0/n338 ) );
  nand_x1_sg U3726 ( .A(n2805), .B(n2806), .X(\max_pooling_0/n336 ) );
  nand_x1_sg U3727 ( .A(n2809), .B(n2810), .X(\max_pooling_0/n334 ) );
  nand_x1_sg U3728 ( .A(n2779), .B(n2780), .X(\max_pooling_0/n349 ) );
  nand_x1_sg U3729 ( .A(n2799), .B(n2800), .X(\max_pooling_0/n339 ) );
  nand_x1_sg U3730 ( .A(n2781), .B(n2782), .X(\max_pooling_0/n348 ) );
  nand_x1_sg U3731 ( .A(n2807), .B(n2808), .X(\max_pooling_0/n335 ) );
  nand_x1_sg U3732 ( .A(n2815), .B(n2816), .X(\max_pooling_0/n331 ) );
  nand_x1_sg U3733 ( .A(n2783), .B(n2784), .X(\max_pooling_0/n347 ) );
  nand_x1_sg U3734 ( .A(n2793), .B(n2794), .X(\max_pooling_0/n342 ) );
  nand_x1_sg U3735 ( .A(n2629), .B(n2630), .X(\min_pooling_0/n413 ) );
  nand_x1_sg U3736 ( .A(n2759), .B(n2760), .X(\mean_pooling_0/n247 ) );
  nand_x1_sg U3737 ( .A(n2768), .B(n2769), .X(\max_pooling_0/n352 ) );
  nand_x1_sg U3738 ( .A(n2787), .B(n2788), .X(\max_pooling_0/n345 ) );
  nand_x1_sg U3739 ( .A(n2795), .B(n2796), .X(\max_pooling_0/n341 ) );
  nand_x1_sg U3740 ( .A(n3057), .B(\max_pooling_0/n321 ), .X(n2796) );
  nand_x1_sg U3741 ( .A(n2797), .B(n2798), .X(\max_pooling_0/n340 ) );
  nand_x1_sg U3742 ( .A(n3056), .B(\max_pooling_0/n320 ), .X(n2798) );
  nand_x1_sg U3743 ( .A(n2803), .B(n2804), .X(\max_pooling_0/n337 ) );
  nand_x1_sg U3744 ( .A(n3057), .B(\max_pooling_0/n317 ), .X(n2804) );
  nand_x1_sg U3745 ( .A(n3633), .B(n2044), .X(n2035) );
  nand_x1_sg U3746 ( .A(n1302), .B(n1303), .X(\min_pooling_0/n310 ) );
  nand_x1_sg U3747 ( .A(n1205), .B(n1206), .X(\min_pooling_0/n390 ) );
  nand_x1_sg U3748 ( .A(n1211), .B(n1212), .X(\min_pooling_0/n386 ) );
  nand_x1_sg U3749 ( .A(n1216), .B(n1217), .X(\min_pooling_0/n382 ) );
  nand_x1_sg U3750 ( .A(n1221), .B(n1222), .X(\min_pooling_0/n378 ) );
  nand_x1_sg U3751 ( .A(n1246), .B(n1247), .X(\min_pooling_0/n358 ) );
  nand_x1_sg U3752 ( .A(n1251), .B(n1252), .X(\min_pooling_0/n354 ) );
  nand_x1_sg U3753 ( .A(n1256), .B(n1257), .X(\min_pooling_0/n350 ) );
  nand_x1_sg U3754 ( .A(n1261), .B(n1262), .X(\min_pooling_0/n346 ) );
  nand_x1_sg U3755 ( .A(n1266), .B(n1267), .X(\min_pooling_0/n342 ) );
  nand_x1_sg U3756 ( .A(n1271), .B(n1272), .X(\min_pooling_0/n338 ) );
  nand_x1_sg U3757 ( .A(n1276), .B(n1277), .X(\min_pooling_0/n334 ) );
  nand_x1_sg U3758 ( .A(n1281), .B(n1282), .X(\min_pooling_0/n330 ) );
  nand_x1_sg U3759 ( .A(n1286), .B(n1287), .X(\min_pooling_0/n326 ) );
  nand_x1_sg U3760 ( .A(n1291), .B(n1292), .X(\min_pooling_0/n322 ) );
  nand_x1_sg U3761 ( .A(n1296), .B(n1297), .X(\min_pooling_0/n318 ) );
  nand_x1_sg U3762 ( .A(n1289), .B(n1290), .X(\min_pooling_0/n325 ) );
  nand_x1_sg U3763 ( .A(n1966), .B(n1967), .X(\max_pooling_0/n229 ) );
  nand_x1_sg U3764 ( .A(n1885), .B(n1886), .X(\max_pooling_0/n297 ) );
  nand_x1_sg U3765 ( .A(n1920), .B(n1921), .X(\max_pooling_0/n269 ) );
  nand_x1_sg U3766 ( .A(n1945), .B(n1946), .X(\max_pooling_0/n249 ) );
  nand_x1_sg U3767 ( .A(n1950), .B(n1951), .X(\max_pooling_0/n245 ) );
  nand_x1_sg U3768 ( .A(n1925), .B(n1926), .X(\max_pooling_0/n265 ) );
  nand_x1_sg U3769 ( .A(n1930), .B(n1931), .X(\max_pooling_0/n261 ) );
  nand_x1_sg U3770 ( .A(n1940), .B(n1941), .X(\max_pooling_0/n253 ) );
  nand_x1_sg U3771 ( .A(n1955), .B(n1956), .X(\max_pooling_0/n241 ) );
  nand_x1_sg U3772 ( .A(n1868), .B(n1869), .X(\max_pooling_0/n309 ) );
  nand_x1_sg U3773 ( .A(n1875), .B(n1876), .X(\max_pooling_0/n305 ) );
  nand_x1_sg U3774 ( .A(n1880), .B(n1881), .X(\max_pooling_0/n301 ) );
  nand_x1_sg U3775 ( .A(n1910), .B(n1911), .X(\max_pooling_0/n277 ) );
  nand_x1_sg U3776 ( .A(n1915), .B(n1916), .X(\max_pooling_0/n273 ) );
  nand_x1_sg U3777 ( .A(n1935), .B(n1936), .X(\max_pooling_0/n257 ) );
  nand_x1_sg U3778 ( .A(n1960), .B(n1961), .X(\max_pooling_0/n237 ) );
  nand_x1_sg U3779 ( .A(n1890), .B(n1891), .X(\max_pooling_0/n293 ) );
  nand_x1_sg U3780 ( .A(n1895), .B(n1896), .X(\max_pooling_0/n289 ) );
  nand_x1_sg U3781 ( .A(n1900), .B(n1901), .X(\max_pooling_0/n285 ) );
  nand_x1_sg U3782 ( .A(n1905), .B(n1906), .X(\max_pooling_0/n281 ) );
  nand_x1_sg U3783 ( .A(n1226), .B(n1227), .X(\min_pooling_0/n374 ) );
  nand_x1_sg U3784 ( .A(n1231), .B(n1232), .X(\min_pooling_0/n370 ) );
  nand_x1_sg U3785 ( .A(n1236), .B(n1237), .X(\min_pooling_0/n366 ) );
  nand_x1_sg U3786 ( .A(n1241), .B(n1242), .X(\min_pooling_0/n362 ) );
  nand_x1_sg U3787 ( .A(n2031), .B(n2032), .X(n2030) );
  nor_x1_sg U3788 ( .A(n3052), .B(n3022), .X(n2634) );
  nor_x1_sg U3789 ( .A(n3128), .B(n3027), .X(n2764) );
  nor_x1_sg U3790 ( .A(n3148), .B(n3101), .X(n2467) );
  nor_x1_sg U3791 ( .A(n1535), .B(n1532), .X(n1696) );
  nor_x1_sg U3792 ( .A(n1544), .B(n1541), .X(n1699) );
  nor_x1_sg U3793 ( .A(n1553), .B(n1550), .X(n1702) );
  nor_x1_sg U3794 ( .A(n1562), .B(n1559), .X(n1705) );
  nor_x1_sg U3795 ( .A(n1571), .B(n1568), .X(n1708) );
  nor_x1_sg U3796 ( .A(n1580), .B(n1577), .X(n1711) );
  nor_x1_sg U3797 ( .A(n1589), .B(n1586), .X(n1714) );
  nor_x1_sg U3798 ( .A(n1598), .B(n1595), .X(n1717) );
  nor_x1_sg U3799 ( .A(n1607), .B(n1604), .X(n1720) );
  nor_x1_sg U3800 ( .A(n1616), .B(n1613), .X(n1723) );
  nor_x1_sg U3801 ( .A(n1625), .B(n1622), .X(n1726) );
  nor_x1_sg U3802 ( .A(n1634), .B(n1631), .X(n1729) );
  nor_x1_sg U3803 ( .A(n1643), .B(n1640), .X(n1732) );
  nor_x1_sg U3804 ( .A(n1652), .B(n1649), .X(n1735) );
  nor_x1_sg U3805 ( .A(n3636), .B(n1658), .X(n1738) );
  inv_x1_sg U3806 ( .A(n1971), .X(n3728) );
  nor_x1_sg U3807 ( .A(n1523), .B(n1526), .X(n1693) );
  nor_x1_sg U3808 ( .A(n1218), .B(n1362), .X(n1361) );
  nor_x1_sg U3809 ( .A(n3009), .B(n3180), .X(n406) );
  inv_x1_sg U3810 ( .A(n1213), .X(n3638) );
  inv_x1_sg U3811 ( .A(n1683), .X(n3625) );
  inv_x1_sg U3812 ( .A(n1253), .X(n3682) );
  inv_x1_sg U3813 ( .A(n1927), .X(n3697) );
  inv_x1_sg U3814 ( .A(n1273), .X(n3704) );
  inv_x1_sg U3815 ( .A(n1932), .X(n3703) );
  inv_x1_sg U3816 ( .A(n1278), .X(n3710) );
  inv_x1_sg U3817 ( .A(n1942), .X(n3714) );
  inv_x1_sg U3818 ( .A(n1667), .X(n3635) );
  inv_x1_sg U3819 ( .A(n1238), .X(n3665) );
  inv_x1_sg U3820 ( .A(n1902), .X(n3669) );
  inv_x1_sg U3821 ( .A(n1892), .X(n3658) );
  inv_x1_sg U3822 ( .A(n1233), .X(n3659) );
  inv_x1_sg U3823 ( .A(n1670), .X(n3630) );
  inv_x1_sg U3824 ( .A(n1526), .X(n3718) );
  inv_x1_sg U3825 ( .A(n1907), .X(n3675) );
  inv_x1_sg U3826 ( .A(n1887), .X(n3652) );
  nor_x1_sg U3827 ( .A(n1671), .B(n3050), .X(\mean_pooling_0/n176 ) );
  nor_x1_sg U3828 ( .A(n3049), .B(n1518), .X(\mean_pooling_0/n244 ) );
  nor_x1_sg U3829 ( .A(n3050), .B(n1536), .X(\mean_pooling_0/n236 ) );
  nor_x1_sg U3830 ( .A(n2910), .B(n1554), .X(\mean_pooling_0/n228 ) );
  nor_x1_sg U3831 ( .A(n3048), .B(n1572), .X(\mean_pooling_0/n220 ) );
  nor_x1_sg U3832 ( .A(n3047), .B(n1590), .X(\mean_pooling_0/n212 ) );
  nor_x1_sg U3833 ( .A(n3047), .B(n1608), .X(\mean_pooling_0/n204 ) );
  nor_x1_sg U3834 ( .A(n2910), .B(n1626), .X(\mean_pooling_0/n196 ) );
  nor_x1_sg U3835 ( .A(n3050), .B(n1644), .X(\mean_pooling_0/n188 ) );
  nor_x1_sg U3836 ( .A(n3050), .B(n1662), .X(\mean_pooling_0/n180 ) );
  nor_x1_sg U3837 ( .A(n2910), .B(n1685), .X(\mean_pooling_0/n164 ) );
  nor_x1_sg U3838 ( .A(n3049), .B(n1527), .X(\mean_pooling_0/n240 ) );
  nor_x1_sg U3839 ( .A(n3049), .B(n1545), .X(\mean_pooling_0/n232 ) );
  nor_x1_sg U3840 ( .A(n2910), .B(n1563), .X(\mean_pooling_0/n224 ) );
  nor_x1_sg U3841 ( .A(n3048), .B(n1581), .X(\mean_pooling_0/n216 ) );
  nor_x1_sg U3842 ( .A(n3048), .B(n1599), .X(\mean_pooling_0/n208 ) );
  nor_x1_sg U3843 ( .A(n3047), .B(n1617), .X(\mean_pooling_0/n200 ) );
  nor_x1_sg U3844 ( .A(n3049), .B(n1635), .X(\mean_pooling_0/n192 ) );
  nor_x1_sg U3845 ( .A(n3047), .B(n1653), .X(\mean_pooling_0/n184 ) );
  nor_x1_sg U3846 ( .A(n2463), .B(n3148), .X(n2468) );
  nor_x1_sg U3847 ( .A(n2964), .B(n2956), .X(n2721) );
  nor_x1_sg U3848 ( .A(n2462), .B(n3148), .X(n2457) );
  nand_x1_sg U3849 ( .A(n2463), .B(n2461), .X(n2462) );
  nor_x1_sg U3850 ( .A(n3752), .B(n3017), .X(n2773) );
  inv_x1_sg U3851 ( .A(n2770), .X(n3752) );
  nor_x1_sg U3852 ( .A(n2092), .B(n2097), .X(n2007) );
  nor_x1_sg U3853 ( .A(n1922), .B(n3193), .X(n2097) );
  nor_x1_sg U3854 ( .A(n1927), .B(n3620), .X(n2092) );
  nor_x1_sg U3855 ( .A(n1200), .B(n1141), .X(n1117) );
  nand_x1_sg U3856 ( .A(n3138), .B(n3115), .X(n1200) );
  nor_x1_sg U3857 ( .A(n1238), .B(n3611), .X(n1457) );
  nor_x1_sg U3858 ( .A(n3629), .B(n1673), .X(n1671) );
  nor_x1_sg U3859 ( .A(n3197), .B(n1675), .X(n1673) );
  nand_x1_sg U3860 ( .A(n1675), .B(n1674), .X(n1676) );
  nand_x1_sg U3861 ( .A(n1957), .B(n3119), .X(n1972) );
  nand_x2_sg U3862 ( .A(n1976), .B(n1977), .X(n1974) );
  nor_x1_sg U3863 ( .A(n1857), .B(n1858), .X(n1853) );
  nor_x1_sg U3864 ( .A(n1855), .B(n1856), .X(n1854) );
  nor_x1_sg U3865 ( .A(n3198), .B(n2882), .X(n1857) );
  nor_x1_sg U3866 ( .A(n1410), .B(n1411), .X(n1406) );
  nor_x1_sg U3867 ( .A(n1408), .B(n1409), .X(n1407) );
  nor_x1_sg U3868 ( .A(n3205), .B(n3044), .X(n1410) );
  nor_x1_sg U3869 ( .A(n1403), .B(n1404), .X(n1399) );
  nor_x1_sg U3870 ( .A(n1401), .B(n1402), .X(n1400) );
  nor_x1_sg U3871 ( .A(n3204), .B(n3045), .X(n1403) );
  nor_x1_sg U3872 ( .A(n1391), .B(n1392), .X(n1387) );
  nor_x1_sg U3873 ( .A(n1389), .B(n1390), .X(n1388) );
  nor_x1_sg U3874 ( .A(n3202), .B(n3042), .X(n1391) );
  nor_x1_sg U3875 ( .A(n1441), .B(n1442), .X(n1437) );
  nor_x1_sg U3876 ( .A(n1439), .B(n1440), .X(n1438) );
  nor_x1_sg U3877 ( .A(n3200), .B(n2884), .X(n1441) );
  nor_x1_sg U3878 ( .A(n1447), .B(n1448), .X(n1443) );
  nor_x1_sg U3879 ( .A(n1445), .B(n1446), .X(n1444) );
  nor_x1_sg U3880 ( .A(n3211), .B(n3045), .X(n1447) );
  nor_x1_sg U3881 ( .A(n2058), .B(n2059), .X(n2054) );
  nor_x1_sg U3882 ( .A(n2056), .B(n2057), .X(n2055) );
  nor_x1_sg U3883 ( .A(n3202), .B(n3033), .X(n2058) );
  nor_x1_sg U3884 ( .A(n2132), .B(n2133), .X(n2128) );
  nor_x1_sg U3885 ( .A(n2130), .B(n2131), .X(n2129) );
  nor_x1_sg U3886 ( .A(n3208), .B(n2907), .X(n2132) );
  nor_x1_sg U3887 ( .A(n2102), .B(n2103), .X(n2098) );
  nor_x1_sg U3888 ( .A(n2100), .B(n2101), .X(n2099) );
  nor_x1_sg U3889 ( .A(n3200), .B(n3035), .X(n2102) );
  nor_x1_sg U3890 ( .A(n2166), .B(n2167), .X(n2162) );
  nor_x1_sg U3891 ( .A(n2164), .B(n2165), .X(n2163) );
  nor_x1_sg U3892 ( .A(n3199), .B(n3033), .X(n2166) );
  nor_x1_sg U3893 ( .A(n2172), .B(n2173), .X(n2168) );
  nor_x1_sg U3894 ( .A(n2170), .B(n2171), .X(n2169) );
  nor_x1_sg U3895 ( .A(n3198), .B(n2880), .X(n2172) );
  nor_x1_sg U3896 ( .A(n2071), .B(n2072), .X(n2067) );
  nor_x1_sg U3897 ( .A(n2069), .B(n2070), .X(n2068) );
  nor_x1_sg U3898 ( .A(n3183), .B(n2907), .X(n2071) );
  nand_x1_sg U3899 ( .A(n3712), .B(n2828), .X(n1698) );
  nand_x1_sg U3900 ( .A(n1541), .B(n1544), .X(n1697) );
  nand_x1_sg U3901 ( .A(n3706), .B(n2829), .X(n1701) );
  nand_x1_sg U3902 ( .A(n1550), .B(n1553), .X(n1700) );
  nand_x1_sg U3903 ( .A(n3701), .B(n2830), .X(n1704) );
  nand_x1_sg U3904 ( .A(n1559), .B(n1562), .X(n1703) );
  nand_x1_sg U3905 ( .A(n3695), .B(n2831), .X(n1707) );
  nand_x1_sg U3906 ( .A(n1568), .B(n1571), .X(n1706) );
  nand_x1_sg U3907 ( .A(n3690), .B(n2832), .X(n1710) );
  nand_x1_sg U3908 ( .A(n1577), .B(n1580), .X(n1709) );
  nand_x1_sg U3909 ( .A(n3684), .B(n2833), .X(n1713) );
  nand_x1_sg U3910 ( .A(n1586), .B(n1589), .X(n1712) );
  nand_x1_sg U3911 ( .A(n3679), .B(n2834), .X(n1716) );
  nand_x1_sg U3912 ( .A(n1595), .B(n1598), .X(n1715) );
  nand_x1_sg U3913 ( .A(n3673), .B(n2835), .X(n1719) );
  nand_x1_sg U3914 ( .A(n1604), .B(n1607), .X(n1718) );
  nand_x1_sg U3915 ( .A(n3667), .B(n2836), .X(n1722) );
  nand_x1_sg U3916 ( .A(n1613), .B(n1616), .X(n1721) );
  nand_x1_sg U3917 ( .A(n3661), .B(n2837), .X(n1725) );
  nand_x1_sg U3918 ( .A(n1622), .B(n1625), .X(n1724) );
  nand_x1_sg U3919 ( .A(n3656), .B(n2838), .X(n1728) );
  nand_x1_sg U3920 ( .A(n1631), .B(n1634), .X(n1727) );
  nand_x1_sg U3921 ( .A(n3650), .B(n2839), .X(n1731) );
  nand_x1_sg U3922 ( .A(n1640), .B(n1643), .X(n1730) );
  nand_x1_sg U3923 ( .A(n3645), .B(n2840), .X(n1734) );
  nand_x1_sg U3924 ( .A(n1649), .B(n1652), .X(n1733) );
  nand_x1_sg U3925 ( .A(n3640), .B(n2826), .X(n1737) );
  nand_x1_sg U3926 ( .A(n1658), .B(n3636), .X(n1736) );
  nor_x1_sg U3927 ( .A(n1851), .B(n1852), .X(n1847) );
  nor_x1_sg U3928 ( .A(n1849), .B(n1850), .X(n1848) );
  nor_x1_sg U3929 ( .A(n3199), .B(n3038), .X(n1851) );
  nor_x1_sg U3930 ( .A(n1845), .B(n1846), .X(n1841) );
  nor_x1_sg U3931 ( .A(n1843), .B(n1844), .X(n1842) );
  nor_x1_sg U3932 ( .A(n3214), .B(n3040), .X(n1845) );
  nor_x1_sg U3933 ( .A(n1839), .B(n1840), .X(n1835) );
  nor_x1_sg U3934 ( .A(n1837), .B(n1838), .X(n1836) );
  nor_x1_sg U3935 ( .A(n3213), .B(n3039), .X(n1839) );
  nor_x1_sg U3936 ( .A(n1833), .B(n1834), .X(n1829) );
  nor_x1_sg U3937 ( .A(n1831), .B(n1832), .X(n1830) );
  nor_x1_sg U3938 ( .A(n3212), .B(n3038), .X(n1833) );
  nor_x1_sg U3939 ( .A(n1827), .B(n1828), .X(n1823) );
  nor_x1_sg U3940 ( .A(n1825), .B(n1826), .X(n1824) );
  nor_x1_sg U3941 ( .A(n3211), .B(n3040), .X(n1827) );
  nor_x1_sg U3942 ( .A(n1821), .B(n1822), .X(n1817) );
  nor_x1_sg U3943 ( .A(n1819), .B(n1820), .X(n1818) );
  nor_x1_sg U3944 ( .A(n3200), .B(n2908), .X(n1821) );
  nor_x1_sg U3945 ( .A(n1809), .B(n1810), .X(n1805) );
  nor_x1_sg U3946 ( .A(n1807), .B(n1808), .X(n1806) );
  nor_x1_sg U3947 ( .A(n3209), .B(n3039), .X(n1809) );
  nor_x1_sg U3948 ( .A(n1803), .B(n1804), .X(n1799) );
  nor_x1_sg U3949 ( .A(n1801), .B(n1802), .X(n1800) );
  nor_x1_sg U3950 ( .A(n3208), .B(n3037), .X(n1803) );
  nor_x1_sg U3951 ( .A(n1773), .B(n1774), .X(n1769) );
  nor_x1_sg U3952 ( .A(n1771), .B(n1772), .X(n1770) );
  nor_x1_sg U3953 ( .A(n3205), .B(n2908), .X(n1773) );
  nor_x1_sg U3954 ( .A(n1767), .B(n1768), .X(n1763) );
  nor_x1_sg U3955 ( .A(n1765), .B(n1766), .X(n1764) );
  nor_x1_sg U3956 ( .A(n3204), .B(n3040), .X(n1767) );
  nor_x1_sg U3957 ( .A(n1815), .B(n1816), .X(n1811) );
  nor_x1_sg U3958 ( .A(n1813), .B(n1814), .X(n1812) );
  nor_x1_sg U3959 ( .A(n3210), .B(n3039), .X(n1815) );
  nor_x1_sg U3960 ( .A(n1797), .B(n1798), .X(n1793) );
  nor_x1_sg U3961 ( .A(n1795), .B(n1796), .X(n1794) );
  nor_x1_sg U3962 ( .A(n3184), .B(n3038), .X(n1797) );
  nor_x1_sg U3963 ( .A(n1791), .B(n1792), .X(n1787) );
  nor_x1_sg U3964 ( .A(n1789), .B(n1790), .X(n1788) );
  nor_x1_sg U3965 ( .A(n3207), .B(n2908), .X(n1791) );
  nor_x1_sg U3966 ( .A(n1785), .B(n1786), .X(n1781) );
  nor_x1_sg U3967 ( .A(n1783), .B(n1784), .X(n1782) );
  nor_x1_sg U3968 ( .A(n3206), .B(n2882), .X(n1785) );
  nor_x1_sg U3969 ( .A(n1779), .B(n1780), .X(n1775) );
  nor_x1_sg U3970 ( .A(n1777), .B(n1778), .X(n1776) );
  nor_x1_sg U3971 ( .A(n3183), .B(n3039), .X(n1779) );
  nor_x1_sg U3972 ( .A(n1145), .B(n3180), .X(n414) );
  nor_x1_sg U3973 ( .A(n1470), .B(n1471), .X(n1466) );
  nor_x1_sg U3974 ( .A(n1468), .B(n1469), .X(n1467) );
  nor_x1_sg U3975 ( .A(n3184), .B(n3042), .X(n1470) );
  nor_x1_sg U3976 ( .A(n2108), .B(n2109), .X(n2104) );
  nor_x1_sg U3977 ( .A(n2106), .B(n2107), .X(n2105) );
  nor_x1_sg U3978 ( .A(n3211), .B(n2907), .X(n2108) );
  nor_x1_sg U3979 ( .A(n1483), .B(n1484), .X(n1479) );
  nor_x1_sg U3980 ( .A(n1481), .B(n1482), .X(n1480) );
  nor_x1_sg U3981 ( .A(n3210), .B(n2909), .X(n1483) );
  nor_x1_sg U3982 ( .A(n1496), .B(n1497), .X(n1492) );
  nor_x1_sg U3983 ( .A(n1494), .B(n1495), .X(n1493) );
  nor_x1_sg U3984 ( .A(n3213), .B(n3045), .X(n1496) );
  nor_x1_sg U3985 ( .A(n2152), .B(n2153), .X(n2148) );
  nor_x1_sg U3986 ( .A(n2150), .B(n2151), .X(n2149) );
  nor_x1_sg U3987 ( .A(n3212), .B(n3034), .X(n2152) );
  nor_x1_sg U3988 ( .A(n1328), .B(n1329), .X(n1323) );
  nor_x1_sg U3989 ( .A(n1325), .B(n1326), .X(n1324) );
  nor_x1_sg U3990 ( .A(n3214), .B(n2909), .X(n1328) );
  nor_x1_sg U3991 ( .A(n1991), .B(n1992), .X(n1986) );
  nor_x1_sg U3992 ( .A(n1988), .B(n1989), .X(n1987) );
  nor_x1_sg U3993 ( .A(n3214), .B(n3035), .X(n1991) );
  nor_x1_sg U3994 ( .A(n1761), .B(n1762), .X(n1757) );
  nor_x1_sg U3995 ( .A(n1759), .B(n1760), .X(n1758) );
  nor_x1_sg U3996 ( .A(n3182), .B(n3038), .X(n1761) );
  nor_x1_sg U3997 ( .A(n1429), .B(n1430), .X(n1425) );
  nor_x1_sg U3998 ( .A(n1427), .B(n1428), .X(n1426) );
  nor_x1_sg U3999 ( .A(n3207), .B(n3044), .X(n1429) );
  nor_x1_sg U4000 ( .A(n2084), .B(n2085), .X(n2080) );
  nor_x1_sg U4001 ( .A(n2082), .B(n2083), .X(n2081) );
  nor_x1_sg U4002 ( .A(n3206), .B(n3034), .X(n2084) );
  nor_x1_sg U4003 ( .A(n2126), .B(n2127), .X(n2122) );
  nor_x1_sg U4004 ( .A(n2124), .B(n2125), .X(n2123) );
  nor_x1_sg U4005 ( .A(n3184), .B(n3035), .X(n2126) );
  nor_x1_sg U4006 ( .A(n3153), .B(n1887), .X(n2066) );
  nand_x1_sg U4007 ( .A(n1675), .B(n1677), .X(n1742) );
  nor_x1_sg U4008 ( .A(n3243), .B(n1263), .X(n1434) );
  nor_x1_sg U4009 ( .A(n3176), .B(n1947), .X(n2161) );
  nor_x1_sg U4010 ( .A(n3612), .B(n1233), .X(n1350) );
  nor_x1_sg U4011 ( .A(n3606), .B(n1273), .X(n1330) );
  nor_x1_sg U4012 ( .A(n3605), .B(n1278), .X(n1320) );
  nand_x1_sg U4013 ( .A(n3717), .B(n2827), .X(n1695) );
  nand_x1_sg U4014 ( .A(n1532), .B(n1535), .X(n1694) );
  nor_x1_sg U4015 ( .A(n3751), .B(n2988), .X(n1395) );
  nor_x1_sg U4016 ( .A(n3751), .B(n2994), .X(n2050) );
  nor_x1_sg U4017 ( .A(n3749), .B(n2989), .X(n1379) );
  nor_x1_sg U4018 ( .A(n3748), .B(n2989), .X(n1401) );
  nor_x1_sg U4019 ( .A(n3749), .B(n2993), .X(n2040) );
  nor_x1_sg U4020 ( .A(n3748), .B(n2991), .X(n2062) );
  nor_x1_sg U4021 ( .A(n3746), .B(n2986), .X(n1414) );
  nor_x1_sg U4022 ( .A(n3746), .B(n2992), .X(n2069) );
  nor_x1_sg U4023 ( .A(n3747), .B(n2991), .X(n2075) );
  nor_x1_sg U4024 ( .A(n3743), .B(n2987), .X(n1468) );
  nor_x1_sg U4025 ( .A(n3741), .B(n2993), .X(n2137) );
  nor_x1_sg U4026 ( .A(n3744), .B(n2991), .X(n2088) );
  nor_x1_sg U4027 ( .A(n3744), .B(n2986), .X(n1427) );
  nor_x1_sg U4028 ( .A(n3741), .B(n2865), .X(n1475) );
  nor_x1_sg U4029 ( .A(n3740), .B(n2867), .X(n2143) );
  nor_x1_sg U4030 ( .A(n3738), .B(n2991), .X(n2106) );
  nor_x1_sg U4031 ( .A(n3740), .B(n2865), .X(n1481) );
  nor_x1_sg U4032 ( .A(n3736), .B(n2987), .X(n1494) );
  nor_x1_sg U4033 ( .A(n3737), .B(n2992), .X(n2150) );
  nor_x1_sg U4034 ( .A(n3737), .B(n2865), .X(n1488) );
  nor_x1_sg U4035 ( .A(n3750), .B(n2983), .X(n1753) );
  nor_x1_sg U4036 ( .A(n3736), .B(n2867), .X(n2156) );
  nor_x1_sg U4037 ( .A(n3735), .B(n2989), .X(n1325) );
  nor_x1_sg U4038 ( .A(n3735), .B(n2994), .X(n1988) );
  nor_x1_sg U4039 ( .A(n3734), .B(n2987), .X(n1502) );
  nor_x1_sg U4040 ( .A(n3732), .B(n2986), .X(n1514) );
  nor_x1_sg U4041 ( .A(n3732), .B(n2994), .X(n2176) );
  nor_x1_sg U4042 ( .A(n3732), .B(n2982), .X(n1864) );
  nor_x1_sg U4043 ( .A(n3745), .B(n2988), .X(n1421) );
  nor_x1_sg U4044 ( .A(n3733), .B(n2986), .X(n1508) );
  nor_x1_sg U4045 ( .A(n3733), .B(n2982), .X(n1855) );
  nor_x1_sg U4046 ( .A(n3734), .B(n2863), .X(n1849) );
  nor_x1_sg U4047 ( .A(n3735), .B(n2863), .X(n1843) );
  nor_x1_sg U4048 ( .A(n3736), .B(n2981), .X(n1837) );
  nor_x1_sg U4049 ( .A(n3737), .B(n2863), .X(n1831) );
  nor_x1_sg U4050 ( .A(n3738), .B(n2982), .X(n1825) );
  nor_x1_sg U4051 ( .A(n3739), .B(n2983), .X(n1819) );
  nor_x1_sg U4052 ( .A(n3740), .B(n2982), .X(n1813) );
  nor_x1_sg U4053 ( .A(n3741), .B(n2981), .X(n1807) );
  nor_x1_sg U4054 ( .A(n3742), .B(n2984), .X(n1801) );
  nor_x1_sg U4055 ( .A(n3743), .B(n2983), .X(n1795) );
  nor_x1_sg U4056 ( .A(n3744), .B(n2984), .X(n1789) );
  nor_x1_sg U4057 ( .A(n3745), .B(n2984), .X(n1783) );
  nor_x1_sg U4058 ( .A(n3746), .B(n2863), .X(n1777) );
  nor_x1_sg U4059 ( .A(n3747), .B(n2981), .X(n1771) );
  nor_x1_sg U4060 ( .A(n3748), .B(n2981), .X(n1765) );
  nor_x1_sg U4061 ( .A(n3749), .B(n2984), .X(n1759) );
  nor_x1_sg U4062 ( .A(n3751), .B(n2983), .X(n1746) );
  nor_x1_sg U4063 ( .A(n3750), .B(n2989), .X(n1389) );
  nor_x1_sg U4064 ( .A(n3747), .B(n2987), .X(n1408) );
  nor_x1_sg U4065 ( .A(n3742), .B(n2865), .X(n1462) );
  nor_x1_sg U4066 ( .A(n3739), .B(n2988), .X(n1439) );
  nor_x1_sg U4067 ( .A(n3738), .B(n2988), .X(n1445) );
  nor_x1_sg U4068 ( .A(n3750), .B(n2993), .X(n2056) );
  nor_x1_sg U4069 ( .A(n3745), .B(n2992), .X(n2082) );
  nor_x1_sg U4070 ( .A(n3743), .B(n2992), .X(n2124) );
  nor_x1_sg U4071 ( .A(n3742), .B(n2994), .X(n2130) );
  nor_x1_sg U4072 ( .A(n3739), .B(n2867), .X(n2100) );
  nor_x1_sg U4073 ( .A(n3734), .B(n2867), .X(n2164) );
  nor_x1_sg U4074 ( .A(n3733), .B(n2993), .X(n2170) );
  nor_x1_sg U4075 ( .A(n3617), .B(n1952), .X(n2160) );
  nor_x1_sg U4076 ( .A(n2092), .B(n2093), .X(n2003) );
  nand_x1_sg U4077 ( .A(n1922), .B(n3193), .X(n2093) );
  nor_x1_sg U4078 ( .A(n1381), .B(n1382), .X(n1377) );
  nor_x1_sg U4079 ( .A(n1379), .B(n1380), .X(n1378) );
  nor_x1_sg U4080 ( .A(n3182), .B(n2884), .X(n1381) );
  nor_x1_sg U4081 ( .A(n1516), .B(n1517), .X(n1512) );
  nor_x1_sg U4082 ( .A(n1514), .B(n1515), .X(n1513) );
  nor_x1_sg U4083 ( .A(n3215), .B(n3045), .X(n1516) );
  nor_x1_sg U4084 ( .A(n2178), .B(n2179), .X(n2174) );
  nor_x1_sg U4085 ( .A(n2176), .B(n2177), .X(n2175) );
  nor_x1_sg U4086 ( .A(n3215), .B(n3034), .X(n2178) );
  nor_x1_sg U4087 ( .A(n1416), .B(n1417), .X(n1412) );
  nor_x1_sg U4088 ( .A(n1414), .B(n1415), .X(n1413) );
  nor_x1_sg U4089 ( .A(n3183), .B(n3043), .X(n1416) );
  nor_x1_sg U4090 ( .A(n1464), .B(n1465), .X(n1460) );
  nor_x1_sg U4091 ( .A(n1462), .B(n1463), .X(n1461) );
  nor_x1_sg U4092 ( .A(n3208), .B(n3043), .X(n1464) );
  nor_x1_sg U4093 ( .A(n3242), .B(n3022), .X(n1396) );
  nor_x1_sg U4094 ( .A(n3192), .B(n2916), .X(n1398) );
  nor_x1_sg U4095 ( .A(n3242), .B(n2874), .X(n2051) );
  nor_x1_sg U4096 ( .A(n3192), .B(n3064), .X(n2053) );
  nor_x1_sg U4097 ( .A(n3241), .B(n2905), .X(n1380) );
  nor_x1_sg U4098 ( .A(n3191), .B(n2917), .X(n1382) );
  nor_x1_sg U4099 ( .A(n3240), .B(n3023), .X(n1402) );
  nor_x1_sg U4100 ( .A(n3239), .B(n3068), .X(n1404) );
  nor_x1_sg U4101 ( .A(n3241), .B(n3020), .X(n2041) );
  nor_x1_sg U4102 ( .A(n3191), .B(n3065), .X(n2043) );
  nor_x1_sg U4103 ( .A(n3240), .B(n2904), .X(n2063) );
  nor_x1_sg U4104 ( .A(n3239), .B(n2913), .X(n2065) );
  nor_x1_sg U4105 ( .A(n3238), .B(n3024), .X(n1415) );
  nor_x1_sg U4106 ( .A(n3190), .B(n2917), .X(n1417) );
  nor_x1_sg U4107 ( .A(n3238), .B(n3018), .X(n2070) );
  nor_x1_sg U4108 ( .A(n3190), .B(n2914), .X(n2072) );
  nor_x1_sg U4109 ( .A(n3237), .B(n3019), .X(n2076) );
  nor_x1_sg U4110 ( .A(n3236), .B(n3066), .X(n2078) );
  nor_x1_sg U4111 ( .A(n3235), .B(n3024), .X(n1469) );
  nor_x1_sg U4112 ( .A(n3234), .B(n3070), .X(n1471) );
  nor_x1_sg U4113 ( .A(n3230), .B(n2874), .X(n2138) );
  nor_x1_sg U4114 ( .A(n3188), .B(n3066), .X(n2140) );
  nor_x1_sg U4115 ( .A(n3233), .B(n3020), .X(n2089) );
  nor_x1_sg U4116 ( .A(n3232), .B(n1965), .X(n2091) );
  nor_x1_sg U4117 ( .A(n3233), .B(n3025), .X(n1428) );
  nor_x1_sg U4118 ( .A(n3232), .B(n3068), .X(n1430) );
  nor_x1_sg U4119 ( .A(n3230), .B(n2905), .X(n1476) );
  nor_x1_sg U4120 ( .A(n3188), .B(n2917), .X(n1478) );
  nor_x1_sg U4121 ( .A(n3229), .B(n2904), .X(n2144) );
  nor_x1_sg U4122 ( .A(n3228), .B(n3066), .X(n2146) );
  nor_x1_sg U4123 ( .A(n3226), .B(n3019), .X(n2107) );
  nor_x1_sg U4124 ( .A(n3225), .B(n3064), .X(n2109) );
  nor_x1_sg U4125 ( .A(n3229), .B(n3023), .X(n1482) );
  nor_x1_sg U4126 ( .A(n3228), .B(n3070), .X(n1484) );
  nor_x1_sg U4127 ( .A(n3223), .B(n3025), .X(n1495) );
  nor_x1_sg U4128 ( .A(n3175), .B(n2916), .X(n1497) );
  nor_x1_sg U4129 ( .A(n3224), .B(n3020), .X(n2151) );
  nor_x1_sg U4130 ( .A(n3186), .B(n2913), .X(n2153) );
  nor_x1_sg U4131 ( .A(n3224), .B(n2876), .X(n1489) );
  nor_x1_sg U4132 ( .A(n3186), .B(n3069), .X(n1491) );
  nor_x1_sg U4133 ( .A(n3222), .B(n3029), .X(n1754) );
  nor_x1_sg U4134 ( .A(n3185), .B(n3073), .X(n1756) );
  nor_x1_sg U4135 ( .A(n3223), .B(n3018), .X(n2157) );
  nor_x1_sg U4136 ( .A(n3175), .B(n3065), .X(n2159) );
  nor_x1_sg U4137 ( .A(n3221), .B(n3023), .X(n1326) );
  nor_x1_sg U4138 ( .A(n3220), .B(n3068), .X(n1329) );
  nor_x1_sg U4139 ( .A(n3221), .B(n3019), .X(n1989) );
  nor_x1_sg U4140 ( .A(n3220), .B(n2913), .X(n1992) );
  nor_x1_sg U4141 ( .A(n3217), .B(n2905), .X(n1503) );
  nor_x1_sg U4142 ( .A(n3174), .B(n1301), .X(n1505) );
  nor_x1_sg U4143 ( .A(n3216), .B(n3025), .X(n1515) );
  nor_x1_sg U4144 ( .A(n3173), .B(n2917), .X(n1517) );
  nor_x1_sg U4145 ( .A(n3216), .B(n3019), .X(n2177) );
  nor_x1_sg U4146 ( .A(n3173), .B(n2914), .X(n2179) );
  nor_x1_sg U4147 ( .A(n3216), .B(n3030), .X(n1865) );
  nor_x1_sg U4148 ( .A(n3173), .B(n3073), .X(n1867) );
  nor_x1_sg U4149 ( .A(n3187), .B(n3024), .X(n1422) );
  nor_x1_sg U4150 ( .A(n3227), .B(n2916), .X(n1424) );
  nor_x1_sg U4151 ( .A(n3219), .B(n3025), .X(n1509) );
  nor_x1_sg U4152 ( .A(n3218), .B(n3069), .X(n1511) );
  nor_x1_sg U4153 ( .A(n3219), .B(n3028), .X(n1856) );
  nor_x1_sg U4154 ( .A(n3218), .B(n3072), .X(n1858) );
  nor_x1_sg U4155 ( .A(n3217), .B(n2906), .X(n1850) );
  nor_x1_sg U4156 ( .A(n3174), .B(n2920), .X(n1852) );
  nor_x1_sg U4157 ( .A(n3221), .B(n3028), .X(n1844) );
  nor_x1_sg U4158 ( .A(n3220), .B(n2920), .X(n1846) );
  nor_x1_sg U4159 ( .A(n3223), .B(n3028), .X(n1838) );
  nor_x1_sg U4160 ( .A(n3175), .B(n3074), .X(n1840) );
  nor_x1_sg U4161 ( .A(n3224), .B(n3029), .X(n1832) );
  nor_x1_sg U4162 ( .A(n3186), .B(n3074), .X(n1834) );
  nor_x1_sg U4163 ( .A(n3226), .B(n3028), .X(n1826) );
  nor_x1_sg U4164 ( .A(n3225), .B(n2919), .X(n1828) );
  nor_x1_sg U4165 ( .A(n3181), .B(n2878), .X(n1820) );
  nor_x1_sg U4166 ( .A(n3201), .B(n2920), .X(n1822) );
  nor_x1_sg U4167 ( .A(n3229), .B(n3030), .X(n1814) );
  nor_x1_sg U4168 ( .A(n3228), .B(n2919), .X(n1816) );
  nor_x1_sg U4169 ( .A(n3230), .B(n3030), .X(n1808) );
  nor_x1_sg U4170 ( .A(n3188), .B(n3074), .X(n1810) );
  nor_x1_sg U4171 ( .A(n3189), .B(n2906), .X(n1802) );
  nor_x1_sg U4172 ( .A(n3231), .B(n3072), .X(n1804) );
  nor_x1_sg U4173 ( .A(n3235), .B(n3030), .X(n1796) );
  nor_x1_sg U4174 ( .A(n3234), .B(n2919), .X(n1798) );
  nor_x1_sg U4175 ( .A(n3233), .B(n3029), .X(n1790) );
  nor_x1_sg U4176 ( .A(n3232), .B(n1684), .X(n1792) );
  nor_x1_sg U4177 ( .A(n3187), .B(n2878), .X(n1784) );
  nor_x1_sg U4178 ( .A(n3227), .B(n3072), .X(n1786) );
  nor_x1_sg U4179 ( .A(n3238), .B(n3027), .X(n1778) );
  nor_x1_sg U4180 ( .A(n3190), .B(n3074), .X(n1780) );
  nor_x1_sg U4181 ( .A(n3237), .B(n2906), .X(n1772) );
  nor_x1_sg U4182 ( .A(n3236), .B(n1684), .X(n1774) );
  nor_x1_sg U4183 ( .A(n3240), .B(n3027), .X(n1766) );
  nor_x1_sg U4184 ( .A(n3239), .B(n2919), .X(n1768) );
  nor_x1_sg U4185 ( .A(n3241), .B(n3029), .X(n1760) );
  nor_x1_sg U4186 ( .A(n3191), .B(n3073), .X(n1762) );
  nor_x1_sg U4187 ( .A(n3242), .B(n2906), .X(n1747) );
  nor_x1_sg U4188 ( .A(n3192), .B(n2920), .X(n1750) );
  nor_x1_sg U4189 ( .A(n3222), .B(n3022), .X(n1390) );
  nor_x1_sg U4190 ( .A(n3185), .B(n3070), .X(n1392) );
  nor_x1_sg U4191 ( .A(n3237), .B(n2876), .X(n1409) );
  nor_x1_sg U4192 ( .A(n3236), .B(n1301), .X(n1411) );
  nor_x1_sg U4193 ( .A(n3189), .B(n3023), .X(n1463) );
  nor_x1_sg U4194 ( .A(n3231), .B(n3070), .X(n1465) );
  nor_x1_sg U4195 ( .A(n3181), .B(n2905), .X(n1440) );
  nor_x1_sg U4196 ( .A(n3201), .B(n2916), .X(n1442) );
  nor_x1_sg U4197 ( .A(n3226), .B(n3024), .X(n1446) );
  nor_x1_sg U4198 ( .A(n3225), .B(n3069), .X(n1448) );
  nor_x1_sg U4199 ( .A(n3222), .B(n2904), .X(n2057) );
  nor_x1_sg U4200 ( .A(n3185), .B(n2914), .X(n2059) );
  nor_x1_sg U4201 ( .A(n3187), .B(n3018), .X(n2083) );
  nor_x1_sg U4202 ( .A(n3227), .B(n2913), .X(n2085) );
  nor_x1_sg U4203 ( .A(n3235), .B(n3018), .X(n2125) );
  nor_x1_sg U4204 ( .A(n3234), .B(n3066), .X(n2127) );
  nor_x1_sg U4205 ( .A(n3189), .B(n3017), .X(n2131) );
  nor_x1_sg U4206 ( .A(n3231), .B(n3065), .X(n2133) );
  nor_x1_sg U4207 ( .A(n3181), .B(n3020), .X(n2101) );
  nor_x1_sg U4208 ( .A(n3201), .B(n3064), .X(n2103) );
  nor_x1_sg U4209 ( .A(n3217), .B(n3017), .X(n2165) );
  nor_x1_sg U4210 ( .A(n3174), .B(n3065), .X(n2167) );
  nor_x1_sg U4211 ( .A(n3219), .B(n2904), .X(n2171) );
  nor_x1_sg U4212 ( .A(n3218), .B(n1965), .X(n2173) );
  nor_x1_sg U4213 ( .A(n3008), .B(n3615), .X(n1163) );
  nor_x1_sg U4214 ( .A(n3178), .B(n3153), .X(n1170) );
  nor_x1_sg U4215 ( .A(n2096), .B(n3698), .X(n2094) );
  nor_x1_sg U4216 ( .A(n2110), .B(n2111), .X(n2096) );
  nor_x1_sg U4217 ( .A(n3134), .B(n3176), .X(n1136) );
  nor_x1_sg U4218 ( .A(n2843), .B(n3243), .X(n1121) );
  nor_x1_sg U4219 ( .A(n3253), .B(n3193), .X(n1198) );
  nor_x1_sg U4220 ( .A(n3008), .B(n3194), .X(n1159) );
  nor_x1_sg U4221 ( .A(n1363), .B(n3614), .X(n1360) );
  nor_x1_sg U4222 ( .A(n1364), .B(n3648), .X(n1363) );
  inv_x1_sg U4223 ( .A(n1362), .X(n3648) );
  nor_x1_sg U4224 ( .A(n1405), .B(n1218), .X(n1364) );
  nor_x1_sg U4225 ( .A(n1435), .B(n1345), .X(n1433) );
  nor_x1_sg U4226 ( .A(n1449), .B(n1450), .X(n1435) );
  nand_x1_sg U4227 ( .A(n1451), .B(n1452), .X(n1450) );
  nor_x1_sg U4228 ( .A(n3609), .B(n1253), .X(n1449) );
  nor_x1_sg U4229 ( .A(n3010), .B(n3605), .X(n1133) );
  nor_x1_sg U4230 ( .A(n3010), .B(n3606), .X(n1129) );
  nor_x1_sg U4231 ( .A(n3008), .B(n3607), .X(n1125) );
  nor_x1_sg U4232 ( .A(n3009), .B(n3609), .X(n1195) );
  nor_x1_sg U4233 ( .A(n2870), .B(n3610), .X(n1191) );
  nor_x1_sg U4234 ( .A(n3010), .B(n3179), .X(n1187) );
  nor_x1_sg U4235 ( .A(n3008), .B(n3611), .X(n1183) );
  nor_x1_sg U4236 ( .A(n3011), .B(n3612), .X(n1179) );
  nor_x1_sg U4237 ( .A(n2870), .B(n3613), .X(n1175) );
  nor_x1_sg U4238 ( .A(n3011), .B(n3614), .X(n1167) );
  nor_x1_sg U4239 ( .A(n3011), .B(n3616), .X(n1155) );
  nor_x1_sg U4240 ( .A(n3009), .B(n3604), .X(n1204) );
  nor_x1_sg U4241 ( .A(n1371), .B(n1372), .X(n1367) );
  nor_x1_sg U4242 ( .A(n3615), .B(n1213), .X(n1371) );
  nand_x1_sg U4243 ( .A(n1383), .B(n1384), .X(n1373) );
  nor_x1_sg U4244 ( .A(n1866), .B(n1867), .X(n1862) );
  nor_x1_sg U4245 ( .A(n1864), .B(n1865), .X(n1863) );
  nor_x1_sg U4246 ( .A(n3215), .B(n2908), .X(n1866) );
  nor_x1_sg U4247 ( .A(n1749), .B(n1750), .X(n1744) );
  nor_x1_sg U4248 ( .A(n1746), .B(n1747), .X(n1745) );
  nor_x1_sg U4249 ( .A(n3203), .B(n3040), .X(n1749) );
  nor_x1_sg U4250 ( .A(n1340), .B(n1341), .X(n1339) );
  nor_x1_sg U4251 ( .A(n1342), .B(n1343), .X(n1341) );
  nor_x1_sg U4252 ( .A(n1258), .B(n1431), .X(n1340) );
  nand_x4_sg U4253 ( .A(n1346), .B(n1347), .X(n1342) );
  nand_x1_sg U4254 ( .A(n1258), .B(n3608), .X(n1436) );
  nand_x1_sg U4255 ( .A(n3243), .B(n1263), .X(n1432) );
  nor_x1_sg U4256 ( .A(n3664), .B(n2079), .X(n2018) );
  inv_x1_sg U4257 ( .A(n2017), .X(n3664) );
  nor_x1_sg U4258 ( .A(n3622), .B(n1892), .X(n2079) );
  nor_x1_sg U4259 ( .A(n3709), .B(n2147), .X(n1999) );
  inv_x1_sg U4260 ( .A(n1998), .X(n3709) );
  nor_x1_sg U4261 ( .A(n3619), .B(n1932), .X(n2147) );
  nand_x1_sg U4262 ( .A(n1223), .B(n3118), .X(n1365) );
  nor_x1_sg U4263 ( .A(n1397), .B(n1398), .X(n1393) );
  nor_x1_sg U4264 ( .A(n1395), .B(n1396), .X(n1394) );
  nor_x1_sg U4265 ( .A(n3203), .B(n3044), .X(n1397) );
  nor_x1_sg U4266 ( .A(n2052), .B(n2053), .X(n2048) );
  nor_x1_sg U4267 ( .A(n2050), .B(n2051), .X(n2049) );
  nor_x1_sg U4268 ( .A(n3203), .B(n3032), .X(n2052) );
  nor_x1_sg U4269 ( .A(n2042), .B(n2043), .X(n2038) );
  nor_x1_sg U4270 ( .A(n2040), .B(n2041), .X(n2039) );
  nor_x1_sg U4271 ( .A(n3182), .B(n3034), .X(n2042) );
  nor_x1_sg U4272 ( .A(n2064), .B(n2065), .X(n2060) );
  nor_x1_sg U4273 ( .A(n2062), .B(n2063), .X(n2061) );
  nor_x1_sg U4274 ( .A(n3204), .B(n3035), .X(n2064) );
  nor_x1_sg U4275 ( .A(n2139), .B(n2140), .X(n2135) );
  nor_x1_sg U4276 ( .A(n2137), .B(n2138), .X(n2136) );
  nor_x1_sg U4277 ( .A(n3209), .B(n2907), .X(n2139) );
  nor_x1_sg U4278 ( .A(n1477), .B(n1478), .X(n1473) );
  nor_x1_sg U4279 ( .A(n1475), .B(n1476), .X(n1474) );
  nor_x1_sg U4280 ( .A(n3209), .B(n3043), .X(n1477) );
  nor_x1_sg U4281 ( .A(n2145), .B(n2146), .X(n2141) );
  nor_x1_sg U4282 ( .A(n2143), .B(n2144), .X(n2142) );
  nor_x1_sg U4283 ( .A(n3210), .B(n2880), .X(n2145) );
  nor_x1_sg U4284 ( .A(n1490), .B(n1491), .X(n1486) );
  nor_x1_sg U4285 ( .A(n1488), .B(n1489), .X(n1487) );
  nor_x1_sg U4286 ( .A(n3212), .B(n2909), .X(n1490) );
  nor_x1_sg U4287 ( .A(n1755), .B(n1756), .X(n1751) );
  nor_x1_sg U4288 ( .A(n1753), .B(n1754), .X(n1752) );
  nor_x1_sg U4289 ( .A(n3202), .B(n3037), .X(n1755) );
  nor_x1_sg U4290 ( .A(n2158), .B(n2159), .X(n2154) );
  nor_x1_sg U4291 ( .A(n2156), .B(n2157), .X(n2155) );
  nor_x1_sg U4292 ( .A(n3213), .B(n3032), .X(n2158) );
  nor_x1_sg U4293 ( .A(n1504), .B(n1505), .X(n1500) );
  nor_x1_sg U4294 ( .A(n1502), .B(n1503), .X(n1501) );
  nor_x1_sg U4295 ( .A(n3199), .B(n3044), .X(n1504) );
  nor_x1_sg U4296 ( .A(n1510), .B(n1511), .X(n1506) );
  nor_x1_sg U4297 ( .A(n1508), .B(n1509), .X(n1507) );
  nor_x1_sg U4298 ( .A(n3198), .B(n3043), .X(n1510) );
  nor_x1_sg U4299 ( .A(n2077), .B(n2078), .X(n2073) );
  nor_x1_sg U4300 ( .A(n2075), .B(n2076), .X(n2074) );
  nor_x1_sg U4301 ( .A(n3205), .B(n3033), .X(n2077) );
  nor_x1_sg U4302 ( .A(n2090), .B(n2091), .X(n2086) );
  nor_x1_sg U4303 ( .A(n2088), .B(n2089), .X(n2087) );
  nor_x1_sg U4304 ( .A(n3207), .B(n3033), .X(n2090) );
  nor_x1_sg U4305 ( .A(n1423), .B(n1424), .X(n1419) );
  nor_x1_sg U4306 ( .A(n1421), .B(n1422), .X(n1420) );
  nor_x1_sg U4307 ( .A(n3206), .B(n2909), .X(n1423) );
  nand_x1_sg U4308 ( .A(n1677), .B(n1678), .X(n1674) );
  nand_x1_sg U4309 ( .A(n1146), .B(n2464), .X(n1093) );
  nor_x1_sg U4310 ( .A(n3245), .B(n1141), .X(n1146) );
  nand_x1_sg U4311 ( .A(n1522), .B(n1523), .X(n1520) );
  nor_x1_sg U4312 ( .A(n1522), .B(n1523), .X(n1521) );
  nand_x1_sg U4313 ( .A(n1531), .B(n1532), .X(n1529) );
  nor_x1_sg U4314 ( .A(n1531), .B(n1532), .X(n1530) );
  nand_x1_sg U4315 ( .A(n1540), .B(n1541), .X(n1538) );
  nor_x1_sg U4316 ( .A(n1540), .B(n1541), .X(n1539) );
  nand_x1_sg U4317 ( .A(n1549), .B(n1550), .X(n1547) );
  nor_x1_sg U4318 ( .A(n1549), .B(n1550), .X(n1548) );
  nand_x1_sg U4319 ( .A(n1558), .B(n1559), .X(n1556) );
  nor_x1_sg U4320 ( .A(n1558), .B(n1559), .X(n1557) );
  nand_x1_sg U4321 ( .A(n1567), .B(n1568), .X(n1565) );
  nor_x1_sg U4322 ( .A(n1567), .B(n1568), .X(n1566) );
  nand_x1_sg U4323 ( .A(n1576), .B(n1577), .X(n1574) );
  nor_x1_sg U4324 ( .A(n1576), .B(n1577), .X(n1575) );
  nand_x1_sg U4325 ( .A(n1585), .B(n1586), .X(n1583) );
  nor_x1_sg U4326 ( .A(n1585), .B(n1586), .X(n1584) );
  nand_x1_sg U4327 ( .A(n1594), .B(n1595), .X(n1592) );
  nor_x1_sg U4328 ( .A(n1594), .B(n1595), .X(n1593) );
  nand_x1_sg U4329 ( .A(n1603), .B(n1604), .X(n1601) );
  nor_x1_sg U4330 ( .A(n1603), .B(n1604), .X(n1602) );
  nand_x1_sg U4331 ( .A(n1612), .B(n1613), .X(n1610) );
  nor_x1_sg U4332 ( .A(n1612), .B(n1613), .X(n1611) );
  nand_x1_sg U4333 ( .A(n1621), .B(n1622), .X(n1619) );
  nor_x1_sg U4334 ( .A(n1621), .B(n1622), .X(n1620) );
  nand_x1_sg U4335 ( .A(n1630), .B(n1631), .X(n1628) );
  nor_x1_sg U4336 ( .A(n1630), .B(n1631), .X(n1629) );
  nand_x1_sg U4337 ( .A(n1639), .B(n1640), .X(n1637) );
  nor_x1_sg U4338 ( .A(n1639), .B(n1640), .X(n1638) );
  nand_x1_sg U4339 ( .A(n1648), .B(n1649), .X(n1646) );
  nor_x1_sg U4340 ( .A(n1648), .B(n1649), .X(n1647) );
  nand_x1_sg U4341 ( .A(n1657), .B(n1658), .X(n1655) );
  nor_x1_sg U4342 ( .A(n1657), .B(n1658), .X(n1656) );
  nand_x1_sg U4343 ( .A(n3631), .B(n3635), .X(n1665) );
  nand_x1_sg U4344 ( .A(n1666), .B(n1667), .X(n1664) );
  nand_x1_sg U4345 ( .A(n1688), .B(n1689), .X(n1687) );
  nor_x1_sg U4346 ( .A(n1689), .B(n1688), .X(n1690) );
  nand_x1_sg U4347 ( .A(n3179), .B(n1459), .X(n1458) );
  nand_x1_sg U4348 ( .A(n1457), .B(n3670), .X(n1459) );
  nand_x1_sg U4349 ( .A(n2007), .B(n3687), .X(n2006) );
  nand_x1_sg U4350 ( .A(n1952), .B(n3617), .X(n1976) );
  nand_x1_sg U4351 ( .A(n1386), .B(n1304), .X(n1383) );
  nand_x1_sg U4352 ( .A(n3116), .B(n1293), .X(n1312) );
  nand_x1_sg U4353 ( .A(n1243), .B(n3179), .X(n1347) );
  nand_x1_sg U4354 ( .A(n1354), .B(n3654), .X(n1353) );
  nor_x1_sg U4355 ( .A(n1355), .B(n3613), .X(n1354) );
  nor_x1_sg U4356 ( .A(n1355), .B(n1418), .X(n1356) );
  nor_x1_sg U4357 ( .A(n1360), .B(n1361), .X(n1358) );
  nand_x1_sg U4358 ( .A(n1472), .B(n3677), .X(n1451) );
  nor_x1_sg U4359 ( .A(n1454), .B(n3610), .X(n1472) );
  nand_x1_sg U4360 ( .A(n1334), .B(n3699), .X(n1333) );
  nor_x1_sg U4361 ( .A(n1335), .B(n3607), .X(n1334) );
  nor_x1_sg U4362 ( .A(n1335), .B(n1485), .X(n1336) );
  nor_x1_sg U4363 ( .A(n1433), .B(n1434), .X(n1338) );
  nand_x2_sg U4364 ( .A(n1317), .B(n1318), .X(n1316) );
  nor_x1_sg U4365 ( .A(n1498), .B(n1499), .X(n1315) );
  nor_x1_sg U4366 ( .A(n1319), .B(n1320), .X(n1317) );
  nand_x1_sg U4367 ( .A(n1887), .B(n3153), .X(n2021) );
  nor_x1_sg U4368 ( .A(n2022), .B(n2023), .X(n2020) );
  nor_x1_sg U4369 ( .A(n3152), .B(n2024), .X(n2023) );
  nand_x1_sg U4370 ( .A(n1208), .B(n3194), .X(n1376) );
  nand_x1_sg U4371 ( .A(n1213), .B(n3615), .X(n1375) );
  nand_x1_sg U4372 ( .A(n1453), .B(n1344), .X(n1452) );
  nor_x1_sg U4373 ( .A(n3671), .B(n1456), .X(n1453) );
  nor_x1_sg U4374 ( .A(n3670), .B(n1457), .X(n1456) );
  nand_x1_sg U4375 ( .A(n3627), .B(n3616), .X(n1384) );
  nor_x1_sg U4376 ( .A(n1304), .B(n1386), .X(n1385) );
  nor_x1_sg U4377 ( .A(n1679), .B(n3048), .X(\mean_pooling_0/n172 ) );
  nor_x1_sg U4378 ( .A(n2160), .B(n2161), .X(n1978) );
  nand_x1_sg U4379 ( .A(n1947), .B(n3176), .X(n1981) );
  nand_x4_sg U4380 ( .A(n2001), .B(n2002), .X(n2000) );
  nor_x1_sg U4381 ( .A(n2003), .B(n2004), .X(n2002) );
  nor_x1_sg U4382 ( .A(n2094), .B(n2095), .X(n2001) );
  nor_x1_sg U4383 ( .A(n3676), .B(n2118), .X(n2114) );
  inv_x1_sg U4384 ( .A(n2120), .X(n3676) );
  nor_x1_sg U4385 ( .A(n2119), .B(n1907), .X(n2118) );
  nor_x1_sg U4386 ( .A(n414), .B(n1144), .X(n413) );
  nor_x1_sg U4387 ( .A(n406), .B(n1144), .X(n405) );
  nor_x1_sg U4388 ( .A(n1093), .B(n1144), .X(n410) );
  nor_x1_sg U4389 ( .A(n3172), .B(n2872), .X(n401) );
  nor_x1_sg U4390 ( .A(n418), .B(n3014), .X(n417) );
  nor_x1_sg U4391 ( .A(n422), .B(n3013), .X(n421) );
  nor_x1_sg U4392 ( .A(n3171), .B(n2872), .X(n425) );
  nor_x1_sg U4393 ( .A(n3170), .B(n1117), .X(n429) );
  nor_x1_sg U4394 ( .A(n3163), .B(n1117), .X(n433) );
  nor_x1_sg U4395 ( .A(n3169), .B(n1117), .X(n437) );
  nor_x1_sg U4396 ( .A(n3162), .B(n2903), .X(n441) );
  nor_x1_sg U4397 ( .A(n3161), .B(n2872), .X(n353) );
  nor_x1_sg U4398 ( .A(n3144), .B(n2903), .X(n357) );
  nor_x1_sg U4399 ( .A(n3157), .B(n3014), .X(n361) );
  nor_x1_sg U4400 ( .A(n3160), .B(n3015), .X(n365) );
  nor_x1_sg U4401 ( .A(n3142), .B(n2903), .X(n369) );
  nor_x1_sg U4402 ( .A(n3168), .B(n2903), .X(n373) );
  nor_x1_sg U4403 ( .A(n3156), .B(n3015), .X(n377) );
  nor_x1_sg U4404 ( .A(n3155), .B(n3015), .X(n381) );
  nor_x1_sg U4405 ( .A(n3143), .B(n3013), .X(n385) );
  nor_x1_sg U4406 ( .A(n3154), .B(n3014), .X(n389) );
  nor_x1_sg U4407 ( .A(n3159), .B(n3015), .X(n393) );
  nor_x1_sg U4408 ( .A(n3140), .B(n3013), .X(n397) );
  nor_x1_sg U4409 ( .A(n3141), .B(n3014), .X(n349) );
  nor_x1_sg U4410 ( .A(n1968), .B(n2046), .X(n2047) );
  nand_x1_sg U4411 ( .A(n2861), .B(n1555), .X(\mean_pooling_0/n227 ) );
  nand_x1_sg U4412 ( .A(n2970), .B(n1564), .X(\mean_pooling_0/n223 ) );
  nand_x1_sg U4413 ( .A(n2861), .B(n1573), .X(\mean_pooling_0/n219 ) );
  nand_x1_sg U4414 ( .A(n2972), .B(n1582), .X(\mean_pooling_0/n215 ) );
  nand_x1_sg U4415 ( .A(n2969), .B(n1591), .X(\mean_pooling_0/n211 ) );
  nand_x1_sg U4416 ( .A(n2972), .B(n1600), .X(\mean_pooling_0/n207 ) );
  nand_x1_sg U4417 ( .A(n2972), .B(n1609), .X(\mean_pooling_0/n203 ) );
  nand_x1_sg U4418 ( .A(n2861), .B(n1618), .X(\mean_pooling_0/n199 ) );
  nand_x1_sg U4419 ( .A(n2971), .B(n1627), .X(\mean_pooling_0/n195 ) );
  nand_x1_sg U4420 ( .A(n2970), .B(n1636), .X(\mean_pooling_0/n191 ) );
  nand_x1_sg U4421 ( .A(n2971), .B(n1645), .X(\mean_pooling_0/n187 ) );
  nand_x1_sg U4422 ( .A(n2969), .B(n1654), .X(\mean_pooling_0/n183 ) );
  nand_x1_sg U4423 ( .A(n2861), .B(n1663), .X(\mean_pooling_0/n179 ) );
  nand_x1_sg U4424 ( .A(n2972), .B(n1672), .X(\mean_pooling_0/n175 ) );
  nand_x1_sg U4425 ( .A(n1671), .B(n3252), .X(n1672) );
  nand_x1_sg U4426 ( .A(n2969), .B(n1680), .X(\mean_pooling_0/n171 ) );
  nand_x1_sg U4427 ( .A(n1679), .B(n3252), .X(n1680) );
  nand_x1_sg U4428 ( .A(n3088), .B(n3616), .X(n1306) );
  nand_x1_sg U4429 ( .A(n2935), .B(n3626), .X(n1305) );
  inv_x1_sg U4430 ( .A(n1304), .X(n3626) );
  nand_x1_sg U4431 ( .A(n3086), .B(n3194), .X(n1210) );
  nand_x1_sg U4432 ( .A(n3092), .B(n3634), .X(n1209) );
  nand_x1_sg U4433 ( .A(n2893), .B(n3615), .X(n1215) );
  nand_x1_sg U4434 ( .A(n3091), .B(n3638), .X(n1214) );
  nand_x1_sg U4435 ( .A(n2933), .B(n3614), .X(n1220) );
  nand_x1_sg U4436 ( .A(n2936), .B(n3643), .X(n1219) );
  nand_x1_sg U4437 ( .A(n3089), .B(n3118), .X(n1225) );
  nand_x1_sg U4438 ( .A(n2895), .B(n3647), .X(n1224) );
  nand_x1_sg U4439 ( .A(n3087), .B(n3613), .X(n1230) );
  nand_x1_sg U4440 ( .A(n3093), .B(n3654), .X(n1229) );
  nand_x1_sg U4441 ( .A(n3087), .B(n3612), .X(n1235) );
  nand_x1_sg U4442 ( .A(n2953), .B(n3659), .X(n1234) );
  nand_x1_sg U4443 ( .A(n2952), .B(n3611), .X(n1240) );
  nand_x1_sg U4444 ( .A(n2954), .B(n3665), .X(n1239) );
  nand_x1_sg U4445 ( .A(n2932), .B(n3179), .X(n1245) );
  nand_x1_sg U4446 ( .A(n2896), .B(n3670), .X(n1244) );
  nand_x1_sg U4447 ( .A(n2933), .B(n3610), .X(n1250) );
  nand_x1_sg U4448 ( .A(n3091), .B(n3677), .X(n1249) );
  nand_x1_sg U4449 ( .A(n2893), .B(n3609), .X(n1255) );
  nand_x1_sg U4450 ( .A(n3093), .B(n3682), .X(n1254) );
  nand_x1_sg U4451 ( .A(n2952), .B(n3608), .X(n1260) );
  nand_x1_sg U4452 ( .A(n2953), .B(n3688), .X(n1259) );
  inv_x1_sg U4453 ( .A(n1258), .X(n3688) );
  nand_x1_sg U4454 ( .A(n2951), .B(n3243), .X(n1265) );
  nand_x1_sg U4455 ( .A(n2895), .B(n3693), .X(n1264) );
  inv_x1_sg U4456 ( .A(n1263), .X(n3693) );
  nand_x1_sg U4457 ( .A(n2951), .B(n3607), .X(n1270) );
  nand_x1_sg U4458 ( .A(n3090), .B(n3699), .X(n1269) );
  nand_x1_sg U4459 ( .A(n2892), .B(n3606), .X(n1275) );
  nand_x1_sg U4460 ( .A(n2936), .B(n3704), .X(n1274) );
  nand_x1_sg U4461 ( .A(n2932), .B(n3605), .X(n1280) );
  nand_x1_sg U4462 ( .A(n3090), .B(n3710), .X(n1279) );
  nand_x1_sg U4463 ( .A(n2933), .B(n3117), .X(n1285) );
  nand_x1_sg U4464 ( .A(n3090), .B(n3715), .X(n1284) );
  nand_x1_sg U4465 ( .A(n3086), .B(n3116), .X(n1295) );
  nand_x1_sg U4466 ( .A(n2954), .B(n3724), .X(n1294) );
  nand_x1_sg U4467 ( .A(n2952), .B(n3604), .X(n1300) );
  nand_x1_sg U4468 ( .A(n2936), .B(n3624), .X(n1299) );
  nand_x1_sg U4469 ( .A(n3152), .B(n2926), .X(n1883) );
  nand_x1_sg U4470 ( .A(n3082), .B(n3150), .X(n1884) );
  nand_x1_sg U4471 ( .A(n3145), .B(n2927), .X(n1963) );
  nand_x1_sg U4472 ( .A(n3084), .B(n3151), .X(n1964) );
  nand_x1_sg U4473 ( .A(n2886), .B(n3632), .X(n1969) );
  nand_x1_sg U4474 ( .A(n2930), .B(n3623), .X(n1970) );
  inv_x1_sg U4475 ( .A(n1968), .X(n3632) );
  nand_x1_sg U4476 ( .A(n3076), .B(n3637), .X(n1873) );
  nand_x1_sg U4477 ( .A(n3082), .B(n3126), .X(n1874) );
  nand_x1_sg U4478 ( .A(n2887), .B(n3642), .X(n1878) );
  nand_x1_sg U4479 ( .A(n2949), .B(n3125), .X(n1879) );
  nand_x1_sg U4480 ( .A(n3076), .B(n3652), .X(n1888) );
  nand_x1_sg U4481 ( .A(n2950), .B(n3153), .X(n1889) );
  nand_x1_sg U4482 ( .A(n2948), .B(n3681), .X(n1913) );
  nand_x1_sg U4483 ( .A(n2890), .B(n3122), .X(n1914) );
  nand_x1_sg U4484 ( .A(n2926), .B(n3686), .X(n1918) );
  nand_x1_sg U4485 ( .A(n2929), .B(n3121), .X(n1919) );
  nand_x1_sg U4486 ( .A(n2947), .B(n3692), .X(n1923) );
  nand_x1_sg U4487 ( .A(n2949), .B(n3193), .X(n1924) );
  inv_x1_sg U4488 ( .A(n1922), .X(n3692) );
  nand_x1_sg U4489 ( .A(n2947), .B(n3697), .X(n1928) );
  nand_x1_sg U4490 ( .A(n3081), .B(n3620), .X(n1929) );
  nand_x1_sg U4491 ( .A(n2948), .B(n3703), .X(n1933) );
  nand_x1_sg U4492 ( .A(n2889), .B(n3619), .X(n1934) );
  nand_x1_sg U4493 ( .A(n2926), .B(n3708), .X(n1938) );
  nand_x1_sg U4494 ( .A(n3081), .B(n3120), .X(n1939) );
  nand_x1_sg U4495 ( .A(n2948), .B(n3714), .X(n1943) );
  nand_x1_sg U4496 ( .A(n2930), .B(n3618), .X(n1944) );
  nand_x1_sg U4497 ( .A(n3079), .B(n3719), .X(n1948) );
  nand_x1_sg U4498 ( .A(n2949), .B(n3176), .X(n1949) );
  inv_x1_sg U4499 ( .A(n1947), .X(n3719) );
  nand_x1_sg U4500 ( .A(n2886), .B(n3723), .X(n1953) );
  nand_x1_sg U4501 ( .A(n2950), .B(n3617), .X(n1954) );
  inv_x1_sg U4502 ( .A(n1952), .X(n3723) );
  nand_x1_sg U4503 ( .A(n3078), .B(n3727), .X(n1958) );
  nand_x1_sg U4504 ( .A(n3084), .B(n3119), .X(n1959) );
  nand_x1_sg U4505 ( .A(n2926), .B(n3658), .X(n1893) );
  nand_x1_sg U4506 ( .A(n3084), .B(n3622), .X(n1894) );
  nand_x1_sg U4507 ( .A(n2947), .B(n3663), .X(n1898) );
  nand_x1_sg U4508 ( .A(n3083), .B(n3124), .X(n1899) );
  nand_x1_sg U4509 ( .A(n3079), .B(n3669), .X(n1903) );
  nand_x1_sg U4510 ( .A(n3081), .B(n3621), .X(n1904) );
  nand_x1_sg U4511 ( .A(n2927), .B(n3675), .X(n1908) );
  nand_x1_sg U4512 ( .A(n2930), .B(n3123), .X(n1909) );
  nor_x1_sg U4513 ( .A(n2628), .B(n3730), .X(n2627) );
  nand_x1_sg U4514 ( .A(n3731), .B(output_taken), .X(n2628) );
  inv_x1_sg U4515 ( .A(state[1]), .X(n3730) );
  nand_x1_sg U4516 ( .A(\im[0][0] ), .B(n3101), .X(n2465) );
  nand_x1_sg U4517 ( .A(\reg_im[0][0] ), .B(n3003), .X(n2466) );
  nand_x1_sg U4518 ( .A(\im[0][1] ), .B(n2945), .X(n2469) );
  nand_x1_sg U4519 ( .A(\reg_im[0][1] ), .B(n3097), .X(n2470) );
  nand_x1_sg U4520 ( .A(\im[0][2] ), .B(n3107), .X(n2471) );
  nand_x1_sg U4521 ( .A(\reg_im[0][2] ), .B(n2998), .X(n2472) );
  nand_x1_sg U4522 ( .A(\im[0][3] ), .B(n2901), .X(n2473) );
  nand_x1_sg U4523 ( .A(\reg_im[0][3] ), .B(n2995), .X(n2474) );
  nand_x1_sg U4524 ( .A(\im[0][4] ), .B(n2940), .X(n2475) );
  nand_x1_sg U4525 ( .A(\reg_im[0][4] ), .B(n3001), .X(n2476) );
  nand_x1_sg U4526 ( .A(\im[0][5] ), .B(n3103), .X(n2477) );
  nand_x1_sg U4527 ( .A(\reg_im[0][5] ), .B(n2939), .X(n2478) );
  nand_x1_sg U4528 ( .A(\im[0][6] ), .B(n3103), .X(n2479) );
  nand_x1_sg U4529 ( .A(\reg_im[0][6] ), .B(n3095), .X(n2480) );
  nand_x1_sg U4530 ( .A(\im[0][7] ), .B(n2940), .X(n2481) );
  nand_x1_sg U4531 ( .A(\reg_im[0][7] ), .B(n2922), .X(n2482) );
  nand_x1_sg U4532 ( .A(\im[0][8] ), .B(n2940), .X(n2483) );
  nand_x1_sg U4533 ( .A(\reg_im[0][8] ), .B(n2922), .X(n2484) );
  nand_x1_sg U4534 ( .A(\im[0][9] ), .B(n2941), .X(n2485) );
  nand_x1_sg U4535 ( .A(\reg_im[0][9] ), .B(n2996), .X(n2486) );
  nand_x1_sg U4536 ( .A(\im[0][10] ), .B(n3106), .X(n2487) );
  nand_x1_sg U4537 ( .A(\reg_im[0][10] ), .B(n2899), .X(n2488) );
  nand_x1_sg U4538 ( .A(\im[0][11] ), .B(n3107), .X(n2489) );
  nand_x1_sg U4539 ( .A(\reg_im[0][11] ), .B(n3003), .X(n2490) );
  nand_x1_sg U4540 ( .A(\im[0][12] ), .B(n3109), .X(n2491) );
  nand_x1_sg U4541 ( .A(\reg_im[0][12] ), .B(n2868), .X(n2492) );
  nand_x1_sg U4542 ( .A(\im[0][13] ), .B(n3111), .X(n2493) );
  nand_x1_sg U4543 ( .A(\reg_im[0][13] ), .B(n3095), .X(n2494) );
  nand_x1_sg U4544 ( .A(\im[0][14] ), .B(n2468), .X(n2495) );
  nand_x1_sg U4545 ( .A(\reg_im[0][14] ), .B(n2995), .X(n2496) );
  nand_x1_sg U4546 ( .A(\im[0][15] ), .B(n3114), .X(n2497) );
  nand_x1_sg U4547 ( .A(\reg_im[0][15] ), .B(n2922), .X(n2498) );
  nand_x1_sg U4548 ( .A(\im[0][16] ), .B(n3104), .X(n2499) );
  nand_x1_sg U4549 ( .A(\reg_im[0][16] ), .B(n3004), .X(n2500) );
  nand_x1_sg U4550 ( .A(\im[0][17] ), .B(n3107), .X(n2501) );
  nand_x1_sg U4551 ( .A(\reg_im[0][17] ), .B(n2999), .X(n2502) );
  nand_x1_sg U4552 ( .A(\im[0][18] ), .B(n3106), .X(n2503) );
  nand_x1_sg U4553 ( .A(\reg_im[0][18] ), .B(n3001), .X(n2504) );
  nand_x1_sg U4554 ( .A(\im[0][19] ), .B(n3108), .X(n2505) );
  nand_x1_sg U4555 ( .A(\reg_im[0][19] ), .B(n3004), .X(n2506) );
  nand_x1_sg U4556 ( .A(\im[1][0] ), .B(n3104), .X(n2507) );
  nand_x1_sg U4557 ( .A(\reg_im[1][0] ), .B(n3000), .X(n2508) );
  nand_x1_sg U4558 ( .A(\im[1][1] ), .B(n2900), .X(n2509) );
  nand_x1_sg U4559 ( .A(\reg_im[1][1] ), .B(n3006), .X(n2510) );
  nand_x1_sg U4560 ( .A(\im[1][2] ), .B(n2941), .X(n2511) );
  nand_x1_sg U4561 ( .A(\reg_im[1][2] ), .B(n2996), .X(n2512) );
  nand_x1_sg U4562 ( .A(\im[1][3] ), .B(n3104), .X(n2513) );
  nand_x1_sg U4563 ( .A(\reg_im[1][3] ), .B(n2938), .X(n2514) );
  nand_x1_sg U4564 ( .A(\im[1][4] ), .B(n2942), .X(n2515) );
  nand_x1_sg U4565 ( .A(\reg_im[1][4] ), .B(n2869), .X(n2516) );
  nand_x1_sg U4566 ( .A(\im[1][15] ), .B(n3113), .X(n2537) );
  nand_x1_sg U4567 ( .A(\reg_im[1][15] ), .B(n2922), .X(n2538) );
  nand_x1_sg U4568 ( .A(\im[1][16] ), .B(n2945), .X(n2539) );
  nand_x1_sg U4569 ( .A(\reg_im[1][16] ), .B(n2939), .X(n2540) );
  nand_x1_sg U4570 ( .A(\im[1][17] ), .B(n3113), .X(n2541) );
  nand_x1_sg U4571 ( .A(\reg_im[1][17] ), .B(n2999), .X(n2542) );
  nand_x1_sg U4572 ( .A(\im[1][18] ), .B(n3112), .X(n2543) );
  nand_x1_sg U4573 ( .A(\reg_im[1][18] ), .B(n3000), .X(n2544) );
  nand_x1_sg U4574 ( .A(\im[1][19] ), .B(n3113), .X(n2545) );
  nand_x1_sg U4575 ( .A(\reg_im[1][19] ), .B(n2996), .X(n2546) );
  nand_x1_sg U4576 ( .A(\im[2][0] ), .B(n3108), .X(n2547) );
  nand_x1_sg U4577 ( .A(\reg_im[2][0] ), .B(n3005), .X(n2548) );
  nand_x1_sg U4578 ( .A(\im[2][1] ), .B(n3108), .X(n2549) );
  nand_x1_sg U4579 ( .A(\reg_im[2][1] ), .B(n3001), .X(n2550) );
  nand_x1_sg U4580 ( .A(\im[2][2] ), .B(n3104), .X(n2551) );
  nand_x1_sg U4581 ( .A(\reg_im[2][2] ), .B(n3000), .X(n2552) );
  nand_x1_sg U4582 ( .A(\im[2][3] ), .B(n3113), .X(n2553) );
  nand_x1_sg U4583 ( .A(\reg_im[2][3] ), .B(n3004), .X(n2554) );
  nand_x1_sg U4584 ( .A(\im[2][4] ), .B(n2944), .X(n2555) );
  nand_x1_sg U4585 ( .A(\reg_im[2][4] ), .B(n2938), .X(n2556) );
  nand_x1_sg U4586 ( .A(\im[2][5] ), .B(n2942), .X(n2557) );
  nand_x1_sg U4587 ( .A(\reg_im[2][5] ), .B(n2921), .X(n2558) );
  nand_x1_sg U4588 ( .A(\im[2][6] ), .B(n3108), .X(n2559) );
  nand_x1_sg U4589 ( .A(\reg_im[2][6] ), .B(n2921), .X(n2560) );
  nand_x1_sg U4590 ( .A(\im[2][7] ), .B(n3101), .X(n2561) );
  nand_x1_sg U4591 ( .A(\reg_im[2][7] ), .B(n3003), .X(n2562) );
  nand_x1_sg U4592 ( .A(\im[2][8] ), .B(n2944), .X(n2563) );
  nand_x1_sg U4593 ( .A(\reg_im[2][8] ), .B(n3096), .X(n2564) );
  nand_x1_sg U4594 ( .A(\im[2][9] ), .B(n3102), .X(n2565) );
  nand_x1_sg U4595 ( .A(\reg_im[2][9] ), .B(n3095), .X(n2566) );
  nand_x1_sg U4596 ( .A(\im[2][10] ), .B(n2900), .X(n2567) );
  nand_x1_sg U4597 ( .A(\reg_im[2][10] ), .B(n2999), .X(n2568) );
  nand_x1_sg U4598 ( .A(\im[2][11] ), .B(n3111), .X(n2569) );
  nand_x1_sg U4599 ( .A(\reg_im[2][11] ), .B(n3098), .X(n2570) );
  nand_x1_sg U4600 ( .A(\im[2][12] ), .B(n2942), .X(n2571) );
  nand_x1_sg U4601 ( .A(\reg_im[2][12] ), .B(n2998), .X(n2572) );
  nand_x1_sg U4602 ( .A(\im[2][13] ), .B(n2945), .X(n2573) );
  nand_x1_sg U4603 ( .A(\reg_im[2][13] ), .B(n2999), .X(n2574) );
  nand_x1_sg U4604 ( .A(\im[2][14] ), .B(n2942), .X(n2575) );
  nand_x1_sg U4605 ( .A(\reg_im[2][14] ), .B(n2868), .X(n2576) );
  nand_x1_sg U4606 ( .A(\im[2][15] ), .B(n3112), .X(n2577) );
  nand_x1_sg U4607 ( .A(\reg_im[2][15] ), .B(n2938), .X(n2578) );
  nand_x1_sg U4608 ( .A(\im[2][16] ), .B(n3103), .X(n2579) );
  nand_x1_sg U4609 ( .A(\reg_im[2][16] ), .B(n2939), .X(n2580) );
  nand_x1_sg U4610 ( .A(\im[2][17] ), .B(n3111), .X(n2581) );
  nand_x1_sg U4611 ( .A(\reg_im[2][17] ), .B(n2998), .X(n2582) );
  nand_x1_sg U4612 ( .A(\im[2][18] ), .B(n3102), .X(n2583) );
  nand_x1_sg U4613 ( .A(\reg_im[2][18] ), .B(n2868), .X(n2584) );
  nand_x1_sg U4614 ( .A(\im[2][19] ), .B(n3107), .X(n2585) );
  nand_x1_sg U4615 ( .A(\reg_im[2][19] ), .B(n2921), .X(n2586) );
  nand_x1_sg U4616 ( .A(\im[3][0] ), .B(n3112), .X(n2587) );
  nand_x1_sg U4617 ( .A(\reg_im[3][0] ), .B(n3097), .X(n2588) );
  nand_x1_sg U4618 ( .A(\im[3][1] ), .B(n3109), .X(n2589) );
  nand_x1_sg U4619 ( .A(\reg_im[3][1] ), .B(n2996), .X(n2590) );
  nand_x1_sg U4620 ( .A(\im[3][2] ), .B(n3114), .X(n2591) );
  nand_x1_sg U4621 ( .A(\reg_im[3][2] ), .B(n2938), .X(n2592) );
  nand_x1_sg U4622 ( .A(\im[3][3] ), .B(n3109), .X(n2593) );
  nand_x1_sg U4623 ( .A(\reg_im[3][3] ), .B(n3096), .X(n2594) );
  nand_x1_sg U4624 ( .A(\im[3][4] ), .B(n2943), .X(n2595) );
  nand_x1_sg U4625 ( .A(\reg_im[3][4] ), .B(n3006), .X(n2596) );
  nand_x1_sg U4626 ( .A(\im[3][5] ), .B(n3109), .X(n2597) );
  nand_x1_sg U4627 ( .A(\reg_im[3][5] ), .B(n3001), .X(n2598) );
  nand_x1_sg U4628 ( .A(\im[3][6] ), .B(n2468), .X(n2599) );
  nand_x1_sg U4629 ( .A(\reg_im[3][6] ), .B(n2995), .X(n2600) );
  nand_x1_sg U4630 ( .A(\im[3][7] ), .B(n3114), .X(n2601) );
  nand_x1_sg U4631 ( .A(\reg_im[3][7] ), .B(n3004), .X(n2602) );
  nand_x1_sg U4632 ( .A(\im[3][8] ), .B(n2945), .X(n2603) );
  nand_x1_sg U4633 ( .A(\reg_im[3][8] ), .B(n3097), .X(n2604) );
  nand_x1_sg U4634 ( .A(\im[3][9] ), .B(n2943), .X(n2605) );
  nand_x1_sg U4635 ( .A(\reg_im[3][9] ), .B(n3005), .X(n2606) );
  nand_x1_sg U4636 ( .A(\im[3][10] ), .B(n2944), .X(n2607) );
  nand_x1_sg U4637 ( .A(\reg_im[3][10] ), .B(n2869), .X(n2608) );
  nand_x1_sg U4638 ( .A(\im[3][11] ), .B(n2900), .X(n2609) );
  nand_x1_sg U4639 ( .A(\reg_im[3][11] ), .B(n2921), .X(n2610) );
  nand_x1_sg U4640 ( .A(\im[3][12] ), .B(n3111), .X(n2611) );
  nand_x1_sg U4641 ( .A(\reg_im[3][12] ), .B(n3096), .X(n2612) );
  nand_x1_sg U4642 ( .A(\im[3][13] ), .B(n2940), .X(n2613) );
  nand_x1_sg U4643 ( .A(\reg_im[3][13] ), .B(n2868), .X(n2614) );
  nand_x1_sg U4644 ( .A(\im[3][14] ), .B(n3106), .X(n2615) );
  nand_x1_sg U4645 ( .A(\reg_im[3][14] ), .B(n2869), .X(n2616) );
  nand_x1_sg U4646 ( .A(\im[3][15] ), .B(n3106), .X(n2617) );
  nand_x1_sg U4647 ( .A(\reg_im[3][15] ), .B(n3096), .X(n2618) );
  nand_x1_sg U4648 ( .A(\im[3][16] ), .B(n2901), .X(n2619) );
  nand_x1_sg U4649 ( .A(\reg_im[3][16] ), .B(n3098), .X(n2620) );
  nand_x1_sg U4650 ( .A(\im[3][17] ), .B(n3103), .X(n2621) );
  nand_x1_sg U4651 ( .A(\reg_im[3][17] ), .B(n3006), .X(n2622) );
  nand_x1_sg U4652 ( .A(\im[3][18] ), .B(n2941), .X(n2623) );
  nand_x1_sg U4653 ( .A(\reg_im[3][18] ), .B(n3006), .X(n2624) );
  nand_x1_sg U4654 ( .A(\im[3][19] ), .B(n3102), .X(n2625) );
  nand_x1_sg U4655 ( .A(\reg_im[3][19] ), .B(n3000), .X(n2626) );
  inv_x1_sg U4656 ( .A(state[0]), .X(n3731) );
  nand_x1_sg U4657 ( .A(\im[1][5] ), .B(n2943), .X(n2517) );
  nand_x1_sg U4658 ( .A(\reg_im[1][5] ), .B(n3095), .X(n2518) );
  nand_x1_sg U4659 ( .A(\im[1][6] ), .B(n2944), .X(n2519) );
  nand_x1_sg U4660 ( .A(\reg_im[1][6] ), .B(n2869), .X(n2520) );
  nand_x1_sg U4661 ( .A(\im[1][7] ), .B(n2901), .X(n2521) );
  nand_x1_sg U4662 ( .A(\reg_im[1][7] ), .B(n2899), .X(n2522) );
  nand_x1_sg U4663 ( .A(\im[1][8] ), .B(n3101), .X(n2523) );
  nand_x1_sg U4664 ( .A(\reg_im[1][8] ), .B(n2939), .X(n2524) );
  nand_x1_sg U4665 ( .A(\im[1][9] ), .B(n2900), .X(n2525) );
  nand_x1_sg U4666 ( .A(\reg_im[1][9] ), .B(n3005), .X(n2526) );
  nand_x1_sg U4667 ( .A(\im[1][10] ), .B(n2943), .X(n2527) );
  nand_x1_sg U4668 ( .A(\reg_im[1][10] ), .B(n3097), .X(n2528) );
  nand_x1_sg U4669 ( .A(\im[1][11] ), .B(n3112), .X(n2529) );
  nand_x1_sg U4670 ( .A(\reg_im[1][11] ), .B(n3003), .X(n2530) );
  nand_x1_sg U4671 ( .A(\im[1][12] ), .B(n2941), .X(n2531) );
  nand_x1_sg U4672 ( .A(\reg_im[1][12] ), .B(n2995), .X(n2532) );
  nand_x1_sg U4673 ( .A(\im[1][13] ), .B(n3114), .X(n2533) );
  nand_x1_sg U4674 ( .A(\reg_im[1][13] ), .B(n2998), .X(n2534) );
  nand_x1_sg U4675 ( .A(\im[1][14] ), .B(n3102), .X(n2535) );
  nand_x1_sg U4676 ( .A(\reg_im[1][14] ), .B(n3005), .X(n2536) );
  nor_x1_sg U4677 ( .A(state[1]), .B(state[0]), .X(n2817) );
  nand_x1_sg U4678 ( .A(n2966), .B(om_mean[0]), .X(n2719) );
  nand_x1_sg U4679 ( .A(n2966), .B(om_mean[1]), .X(n2722) );
  nand_x1_sg U4680 ( .A(n2962), .B(n2826), .X(n2723) );
  nand_x1_sg U4681 ( .A(n2965), .B(om_mean[2]), .X(n2724) );
  nand_x1_sg U4682 ( .A(n2959), .B(n2840), .X(n2725) );
  nand_x1_sg U4683 ( .A(n2964), .B(om_mean[3]), .X(n2726) );
  nand_x1_sg U4684 ( .A(n2959), .B(n2839), .X(n2727) );
  nand_x1_sg U4685 ( .A(n2965), .B(om_mean[4]), .X(n2728) );
  nand_x1_sg U4686 ( .A(n2960), .B(n2838), .X(n2729) );
  nand_x1_sg U4687 ( .A(n2966), .B(om_mean[5]), .X(n2730) );
  nand_x1_sg U4688 ( .A(n2959), .B(n2837), .X(n2731) );
  nand_x1_sg U4689 ( .A(n2859), .B(om_mean[6]), .X(n2732) );
  nand_x1_sg U4690 ( .A(n2960), .B(n2836), .X(n2733) );
  nand_x1_sg U4691 ( .A(n2964), .B(om_mean[7]), .X(n2734) );
  nand_x1_sg U4692 ( .A(n2959), .B(n2835), .X(n2735) );
  nand_x1_sg U4693 ( .A(n2964), .B(om_mean[8]), .X(n2736) );
  nand_x1_sg U4694 ( .A(n2961), .B(n2834), .X(n2737) );
  nand_x1_sg U4695 ( .A(n2967), .B(om_mean[9]), .X(n2738) );
  nand_x1_sg U4696 ( .A(n2962), .B(n2833), .X(n2739) );
  nand_x1_sg U4697 ( .A(n2967), .B(om_mean[10]), .X(n2740) );
  nand_x1_sg U4698 ( .A(n2961), .B(n2832), .X(n2741) );
  nand_x1_sg U4699 ( .A(n2965), .B(om_mean[11]), .X(n2742) );
  nand_x1_sg U4700 ( .A(n2961), .B(n2831), .X(n2743) );
  nand_x1_sg U4701 ( .A(n2859), .B(om_mean[12]), .X(n2744) );
  nand_x1_sg U4702 ( .A(n2962), .B(n2830), .X(n2745) );
  nand_x1_sg U4703 ( .A(n2859), .B(om_mean[13]), .X(n2746) );
  nand_x1_sg U4704 ( .A(n2962), .B(n2829), .X(n2747) );
  nand_x1_sg U4705 ( .A(n2966), .B(om_mean[14]), .X(n2748) );
  nand_x1_sg U4706 ( .A(n2961), .B(n2828), .X(n2749) );
  nand_x1_sg U4707 ( .A(n2967), .B(om_mean[15]), .X(n2750) );
  nand_x1_sg U4708 ( .A(n2721), .B(n2827), .X(n2751) );
  nand_x1_sg U4709 ( .A(n2967), .B(om_mean[16]), .X(n2752) );
  nand_x1_sg U4710 ( .A(n2721), .B(n2823), .X(n2753) );
  nand_x1_sg U4711 ( .A(n2965), .B(om_mean[17]), .X(n2754) );
  nand_x1_sg U4712 ( .A(n2960), .B(n2821), .X(n2755) );
  nor_x1_sg U4713 ( .A(n2818), .B(n2957), .X(n2631) );
  nor_x1_sg U4714 ( .A(n2820), .B(n2957), .X(n2761) );
  nor_x1_sg U4715 ( .A(n3052), .B(\min_pooling_0/n264 ), .X(n2645) );
  nor_x1_sg U4716 ( .A(n3052), .B(\min_pooling_0/n262 ), .X(n2653) );
  nor_x1_sg U4717 ( .A(n2911), .B(\min_pooling_0/n260 ), .X(n2661) );
  nor_x1_sg U4718 ( .A(n3055), .B(\min_pooling_0/n258 ), .X(n2669) );
  nor_x1_sg U4719 ( .A(n3055), .B(\min_pooling_0/n256 ), .X(n2677) );
  nor_x1_sg U4720 ( .A(n3054), .B(\min_pooling_0/n254 ), .X(n2685) );
  nor_x1_sg U4721 ( .A(n3055), .B(\min_pooling_0/n252 ), .X(n2693) );
  nor_x1_sg U4722 ( .A(n3053), .B(\min_pooling_0/n250 ), .X(n2701) );
  nor_x1_sg U4723 ( .A(n2911), .B(\min_pooling_0/n248 ), .X(n2709) );
  nor_x1_sg U4724 ( .A(n3054), .B(\min_pooling_0/n246 ), .X(n2717) );
  nand_x1_sg U4725 ( .A(n2818), .B(om_min[15]), .X(n2660) );
  nor_x1_sg U4726 ( .A(n2661), .B(n2662), .X(n2659) );
  nor_x1_sg U4727 ( .A(n3736), .B(n2979), .X(n2662) );
  nand_x1_sg U4728 ( .A(n2818), .B(om_min[11]), .X(n2676) );
  nor_x1_sg U4729 ( .A(n2677), .B(n2678), .X(n2675) );
  nor_x1_sg U4730 ( .A(n3740), .B(n2976), .X(n2678) );
  nand_x1_sg U4731 ( .A(n2818), .B(om_min[7]), .X(n2692) );
  nor_x1_sg U4732 ( .A(n2693), .B(n2694), .X(n2691) );
  nor_x1_sg U4733 ( .A(n3744), .B(n2976), .X(n2694) );
  nand_x1_sg U4734 ( .A(n2818), .B(om_min[3]), .X(n2708) );
  nor_x1_sg U4735 ( .A(n2709), .B(n2710), .X(n2707) );
  nor_x1_sg U4736 ( .A(n3748), .B(n2978), .X(n2710) );
  nand_x1_sg U4737 ( .A(n2818), .B(n2848), .X(n2644) );
  nor_x1_sg U4738 ( .A(n2645), .B(n2646), .X(n2643) );
  nor_x1_sg U4739 ( .A(n3732), .B(n2978), .X(n2646) );
  nand_x1_sg U4740 ( .A(n2818), .B(n2849), .X(n2652) );
  nor_x1_sg U4741 ( .A(n2653), .B(n2654), .X(n2651) );
  nor_x1_sg U4742 ( .A(n3734), .B(n2977), .X(n2654) );
  nand_x1_sg U4743 ( .A(n2818), .B(n2850), .X(n2700) );
  nor_x1_sg U4744 ( .A(n2701), .B(n2702), .X(n2699) );
  nor_x1_sg U4745 ( .A(n3746), .B(n2978), .X(n2702) );
  nand_x1_sg U4746 ( .A(\min_pooling_0/N4 ), .B(n2818), .X(n2633) );
  nor_x1_sg U4747 ( .A(n2634), .B(n2635), .X(n2632) );
  nor_x1_sg U4748 ( .A(n2957), .B(n3042), .X(n2635) );
  nand_x1_sg U4749 ( .A(\mean_pooling_0/N5 ), .B(n2820), .X(n2763) );
  nor_x1_sg U4750 ( .A(n2764), .B(n2765), .X(n2762) );
  nor_x1_sg U4751 ( .A(n2956), .B(n3037), .X(n2765) );
  nand_x1_sg U4752 ( .A(n2818), .B(om_min[13]), .X(n2668) );
  nor_x1_sg U4753 ( .A(n2669), .B(n2670), .X(n2667) );
  nor_x1_sg U4754 ( .A(n3738), .B(n2978), .X(n2670) );
  nand_x1_sg U4755 ( .A(n2818), .B(om_min[9]), .X(n2684) );
  nor_x1_sg U4756 ( .A(n2685), .B(n2686), .X(n2683) );
  nor_x1_sg U4757 ( .A(n3742), .B(n2979), .X(n2686) );
  nand_x1_sg U4758 ( .A(n2818), .B(om_min[1]), .X(n2716) );
  nor_x1_sg U4759 ( .A(n2717), .B(n2718), .X(n2715) );
  nor_x1_sg U4760 ( .A(n3750), .B(n2976), .X(n2718) );
  nor_x1_sg U4761 ( .A(n3053), .B(\min_pooling_0/n265 ), .X(n2640) );
  nor_x1_sg U4762 ( .A(n3055), .B(\min_pooling_0/n263 ), .X(n2649) );
  nor_x1_sg U4763 ( .A(n3054), .B(\min_pooling_0/n261 ), .X(n2657) );
  nor_x1_sg U4764 ( .A(n2911), .B(\min_pooling_0/n259 ), .X(n2665) );
  nor_x1_sg U4765 ( .A(n2911), .B(\min_pooling_0/n257 ), .X(n2673) );
  nor_x1_sg U4766 ( .A(n3053), .B(\min_pooling_0/n255 ), .X(n2681) );
  nor_x1_sg U4767 ( .A(n3053), .B(\min_pooling_0/n253 ), .X(n2689) );
  nor_x1_sg U4768 ( .A(n3054), .B(\min_pooling_0/n251 ), .X(n2697) );
  nor_x1_sg U4769 ( .A(n3132), .B(\min_pooling_0/n249 ), .X(n2705) );
  nor_x1_sg U4770 ( .A(n3052), .B(\min_pooling_0/n247 ), .X(n2713) );
  nand_x1_sg U4771 ( .A(n2818), .B(om_min[0]), .X(n2639) );
  nor_x1_sg U4772 ( .A(n2640), .B(n2641), .X(n2638) );
  nor_x1_sg U4773 ( .A(n3751), .B(n2975), .X(n2641) );
  nand_x1_sg U4774 ( .A(n2818), .B(om_min[12]), .X(n2672) );
  nor_x1_sg U4775 ( .A(n2673), .B(n2674), .X(n2671) );
  nor_x1_sg U4776 ( .A(n3739), .B(n2976), .X(n2674) );
  nand_x1_sg U4777 ( .A(n2818), .B(\min_pooling_0/n722 ), .X(n2656) );
  nor_x1_sg U4778 ( .A(n2657), .B(n2658), .X(n2655) );
  nor_x1_sg U4779 ( .A(n3735), .B(n2975), .X(n2658) );
  nand_x1_sg U4780 ( .A(n2818), .B(\min_pooling_0/n723 ), .X(n2664) );
  nor_x1_sg U4781 ( .A(n2665), .B(n2666), .X(n2663) );
  nor_x1_sg U4782 ( .A(n3737), .B(n2977), .X(n2666) );
  nand_x1_sg U4783 ( .A(n2818), .B(om_min[10]), .X(n2680) );
  nor_x1_sg U4784 ( .A(n2681), .B(n2682), .X(n2679) );
  nor_x1_sg U4785 ( .A(n3741), .B(n2977), .X(n2682) );
  nand_x1_sg U4786 ( .A(n2818), .B(om_min[8]), .X(n2688) );
  nor_x1_sg U4787 ( .A(n2689), .B(n2690), .X(n2687) );
  nor_x1_sg U4788 ( .A(n3743), .B(n2977), .X(n2690) );
  nand_x1_sg U4789 ( .A(n2818), .B(om_min[6]), .X(n2696) );
  nor_x1_sg U4790 ( .A(n2697), .B(n2698), .X(n2695) );
  nor_x1_sg U4791 ( .A(n3745), .B(n2979), .X(n2698) );
  nand_x1_sg U4792 ( .A(n2818), .B(om_min[18]), .X(n2648) );
  nor_x1_sg U4793 ( .A(n2649), .B(n2650), .X(n2647) );
  nor_x1_sg U4794 ( .A(n3733), .B(n2975), .X(n2650) );
  nand_x1_sg U4795 ( .A(n2818), .B(om_min[4]), .X(n2704) );
  nor_x1_sg U4796 ( .A(n2705), .B(n2706), .X(n2703) );
  nor_x1_sg U4797 ( .A(n3747), .B(n2975), .X(n2706) );
  nand_x1_sg U4798 ( .A(n2818), .B(\min_pooling_0/n724 ), .X(n2712) );
  nor_x1_sg U4799 ( .A(n2713), .B(n2714), .X(n2711) );
  nor_x1_sg U4800 ( .A(n3749), .B(n2979), .X(n2714) );
  nand_x1_sg U4801 ( .A(n2457), .B(state[0]), .X(n2458) );
  nor_x1_sg U4802 ( .A(n2457), .B(n3146), .X(n2460) );
  nand_x1_sg U4803 ( .A(n2456), .B(n3146), .X(n2455) );
  nand_x1_sg U4804 ( .A(n2457), .B(state[1]), .X(n2454) );
  nand_x1_sg U4805 ( .A(\max_pooling_0/N4 ), .B(n2819), .X(n2772) );
  nor_x1_sg U4806 ( .A(n2773), .B(n2774), .X(n2771) );
  nor_x1_sg U4807 ( .A(reg_input_ready), .B(n3032), .X(n2774) );
  nor_x1_sg U4808 ( .A(n3731), .B(state[1]), .X(n2464) );
  nand_x1_sg U4809 ( .A(\max_pooling_0/N3 ), .B(n3247), .X(n2776) );
  nand_x1_sg U4810 ( .A(\min_pooling_0/N3 ), .B(n3603), .X(n2637) );
  nand_x1_sg U4811 ( .A(\mean_pooling_0/N4 ), .B(n3246), .X(n2767) );
  inv_x1_sg U4812 ( .A(\min_pooling_0/N4 ), .X(n3603) );
  inv_x1_sg U4813 ( .A(\mean_pooling_0/N4 ), .X(n3753) );
  nand_x1_sg U4814 ( .A(\max_pooling_0/N4 ), .B(n3195), .X(n2775) );
  nand_x1_sg U4815 ( .A(\mean_pooling_0/N5 ), .B(n3753), .X(n2766) );
  nand_x1_sg U4816 ( .A(\min_pooling_0/N4 ), .B(n3248), .X(n2636) );
  nand_x1_sg U4817 ( .A(n2819), .B(n2852), .X(n2787) );
  nand_x1_sg U4818 ( .A(n2819), .B(n2853), .X(n2795) );
  nand_x1_sg U4819 ( .A(n2819), .B(n2854), .X(n2797) );
  nand_x1_sg U4820 ( .A(n2819), .B(n2856), .X(n2803) );
  nand_x1_sg U4821 ( .A(n2819), .B(n2857), .X(n2811) );
  nand_x1_sg U4822 ( .A(n3058), .B(\max_pooling_0/n313 ), .X(n2812) );
  nand_x1_sg U4823 ( .A(n2819), .B(n2858), .X(n2813) );
  nand_x1_sg U4824 ( .A(n3058), .B(\max_pooling_0/n312 ), .X(n2814) );
  nand_x1_sg U4825 ( .A(n2819), .B(n2851), .X(n2779) );
  nand_x1_sg U4826 ( .A(n3061), .B(\max_pooling_0/n329 ), .X(n2780) );
  nand_x1_sg U4827 ( .A(n2819), .B(n2855), .X(n2799) );
  nand_x1_sg U4828 ( .A(n3062), .B(\max_pooling_0/n319 ), .X(n2800) );
  nand_x1_sg U4829 ( .A(n2819), .B(om_max[0]), .X(n2777) );
  nand_x1_sg U4830 ( .A(n3057), .B(\max_pooling_0/n330 ), .X(n2778) );
  nand_x1_sg U4831 ( .A(n2819), .B(om_max[16]), .X(n2785) );
  nand_x1_sg U4832 ( .A(n3056), .B(\max_pooling_0/n326 ), .X(n2786) );
  nand_x1_sg U4833 ( .A(n2819), .B(om_max[14]), .X(n2789) );
  nand_x1_sg U4834 ( .A(n3058), .B(\max_pooling_0/n324 ), .X(n2790) );
  nand_x1_sg U4835 ( .A(n2819), .B(om_max[13]), .X(n2791) );
  nand_x1_sg U4836 ( .A(n3057), .B(\max_pooling_0/n323 ), .X(n2792) );
  nand_x1_sg U4837 ( .A(n2819), .B(\max_pooling_0/n641 ), .X(n2801) );
  nand_x1_sg U4838 ( .A(n3062), .B(\max_pooling_0/n318 ), .X(n2802) );
  nand_x1_sg U4839 ( .A(n2819), .B(\max_pooling_0/n642 ), .X(n2805) );
  nand_x1_sg U4840 ( .A(n3059), .B(\max_pooling_0/n316 ), .X(n2806) );
  nand_x1_sg U4841 ( .A(n2819), .B(\max_pooling_0/n643 ), .X(n2809) );
  nand_x1_sg U4842 ( .A(n3058), .B(\max_pooling_0/n314 ), .X(n2810) );
  nand_x1_sg U4843 ( .A(n2818), .B(\min_pooling_0/N3 ), .X(n2629) );
  nand_x1_sg U4844 ( .A(n2631), .B(n3248), .X(n2630) );
  nand_x1_sg U4845 ( .A(n2820), .B(\mean_pooling_0/N4 ), .X(n2759) );
  nand_x1_sg U4846 ( .A(n2761), .B(n3753), .X(n2760) );
  nand_x1_sg U4847 ( .A(n2819), .B(\max_pooling_0/N3 ), .X(n2768) );
  nand_x1_sg U4848 ( .A(n3059), .B(n3195), .X(n2769) );
  nand_x1_sg U4849 ( .A(n2819), .B(om_max[18]), .X(n2781) );
  nand_x1_sg U4850 ( .A(n3059), .B(\max_pooling_0/n328 ), .X(n2782) );
  nand_x1_sg U4851 ( .A(n2819), .B(om_max[5]), .X(n2807) );
  nand_x1_sg U4852 ( .A(n3061), .B(\max_pooling_0/n315 ), .X(n2808) );
  nand_x1_sg U4853 ( .A(n2819), .B(om_max[1]), .X(n2815) );
  nand_x1_sg U4854 ( .A(n3056), .B(\max_pooling_0/n311 ), .X(n2816) );
  nand_x1_sg U4855 ( .A(n2819), .B(om_max[17]), .X(n2783) );
  nand_x1_sg U4856 ( .A(n3056), .B(\max_pooling_0/n327 ), .X(n2784) );
  nand_x1_sg U4857 ( .A(n2819), .B(\max_pooling_0/n639 ), .X(n2793) );
  nand_x1_sg U4858 ( .A(n3062), .B(\max_pooling_0/n322 ), .X(n2794) );
  nor_x1_sg U4859 ( .A(reset), .B(n2463), .X(N112) );
  inv_x1_sg U4860 ( .A(\reg_im[0][0] ), .X(n3751) );
  inv_x1_sg U4861 ( .A(\reg_im[0][19] ), .X(n3732) );
  inv_x1_sg U4862 ( .A(\reg_im[0][18] ), .X(n3733) );
  inv_x1_sg U4863 ( .A(\reg_im[0][17] ), .X(n3734) );
  inv_x1_sg U4864 ( .A(\reg_im[0][16] ), .X(n3735) );
  inv_x1_sg U4865 ( .A(\reg_im[0][15] ), .X(n3736) );
  inv_x1_sg U4866 ( .A(\reg_im[0][14] ), .X(n3737) );
  inv_x1_sg U4867 ( .A(\reg_im[0][13] ), .X(n3738) );
  inv_x1_sg U4868 ( .A(\reg_im[0][12] ), .X(n3739) );
  inv_x1_sg U4869 ( .A(\reg_im[0][11] ), .X(n3740) );
  inv_x1_sg U4870 ( .A(\reg_im[0][10] ), .X(n3741) );
  inv_x1_sg U4871 ( .A(\reg_im[0][9] ), .X(n3742) );
  inv_x1_sg U4872 ( .A(\reg_im[0][8] ), .X(n3743) );
  inv_x1_sg U4873 ( .A(\reg_im[0][7] ), .X(n3744) );
  inv_x1_sg U4874 ( .A(\reg_im[0][6] ), .X(n3745) );
  inv_x1_sg U4875 ( .A(\reg_im[0][5] ), .X(n3746) );
  inv_x1_sg U4876 ( .A(\reg_im[0][4] ), .X(n3747) );
  inv_x1_sg U4877 ( .A(\reg_im[0][3] ), .X(n3748) );
  inv_x1_sg U4878 ( .A(\reg_im[0][2] ), .X(n3749) );
  inv_x1_sg U4879 ( .A(\reg_im[0][1] ), .X(n3750) );
  nor_x1_sg U4880 ( .A(n1147), .B(n3180), .X(n1144) );
  nor_x1_sg U4881 ( .A(om_min[7]), .B(n3659), .X(n1355) );
  nor_x1_sg U4882 ( .A(om_min[11]), .B(n3682), .X(n1454) );
  nor_x1_sg U4883 ( .A(om_min[15]), .B(n3704), .X(n1335) );
  nor_x1_sg U4884 ( .A(om_max[0]), .B(n3145), .X(n2046) );
  nor_x1_sg U4885 ( .A(\max_pooling_0/n641 ), .B(n3669), .X(n2119) );
  nor_x1_sg U4886 ( .A(om_min[18]), .B(n3720), .X(n1498) );
  inv_x1_sg U4887 ( .A(om_min[3]), .X(n3615) );
  nor_x1_sg U4888 ( .A(om_max[11]), .B(n3686), .X(n2110) );
  nor_x1_sg U4889 ( .A(om_min[17]), .B(n3715), .X(n1499) );
  nor_x1_sg U4890 ( .A(n3647), .B(om_min[5]), .X(n1405) );
  nor_x1_sg U4891 ( .A(n3635), .B(n3630), .X(n1739) );
  nor_x1_sg U4892 ( .A(n1670), .B(n1667), .X(n1741) );
  inv_x1_sg U4893 ( .A(\min_pooling_0/n722 ), .X(n3605) );
  inv_x1_sg U4894 ( .A(om_min[15]), .X(n3606) );
  inv_x1_sg U4895 ( .A(\min_pooling_0/n723 ), .X(n3607) );
  inv_x1_sg U4896 ( .A(om_min[11]), .X(n3609) );
  inv_x1_sg U4897 ( .A(om_min[10]), .X(n3610) );
  inv_x1_sg U4898 ( .A(om_min[6]), .X(n3613) );
  inv_x1_sg U4899 ( .A(om_min[7]), .X(n3612) );
  inv_x1_sg U4900 ( .A(om_min[8]), .X(n3611) );
  inv_x1_sg U4901 ( .A(\max_pooling_0/n642 ), .X(n3622) );
  inv_x1_sg U4902 ( .A(\max_pooling_0/n641 ), .X(n3621) );
  inv_x1_sg U4903 ( .A(om_max[13]), .X(n3620) );
  inv_x1_sg U4904 ( .A(om_max[14]), .X(n3619) );
  inv_x1_sg U4905 ( .A(om_max[16]), .X(n3618) );
  nor_x1_sg U4906 ( .A(om_max[2]), .B(n3637), .X(n2031) );
  nor_x1_sg U4907 ( .A(\max_pooling_0/n643 ), .B(n2025), .X(n2022) );
  nor_x1_sg U4908 ( .A(n2026), .B(n3653), .X(n2025) );
  inv_x1_sg U4909 ( .A(n2024), .X(n3653) );
  nor_x1_sg U4910 ( .A(n3152), .B(n2066), .X(n2026) );
  nor_x1_sg U4911 ( .A(om_min[6]), .B(n3654), .X(n1418) );
  nor_x1_sg U4912 ( .A(om_max[13]), .B(n3697), .X(n2095) );
  nor_x1_sg U4913 ( .A(\min_pooling_0/n723 ), .B(n3699), .X(n1485) );
  nor_x1_sg U4914 ( .A(n1454), .B(n1455), .X(n1344) );
  nor_x1_sg U4915 ( .A(n3677), .B(om_min[10]), .X(n1455) );
  nor_x1_sg U4916 ( .A(n2821), .B(n3725), .X(n1860) );
  nor_x1_sg U4917 ( .A(n1861), .B(n1113), .X(n1859) );
  inv_x1_sg U4918 ( .A(n1861), .X(n3725) );
  nor_x1_sg U4919 ( .A(n2825), .B(n3625), .X(n1682) );
  nor_x1_sg U4920 ( .A(n1683), .B(n1094), .X(n1681) );
  nor_x1_sg U4921 ( .A(n3721), .B(n3718), .X(n1691) );
  inv_x1_sg U4922 ( .A(n1523), .X(n3721) );
  inv_x1_sg U4923 ( .A(om_min[12]), .X(n3608) );
  inv_x1_sg U4924 ( .A(om_max[18]), .X(n3617) );
  nand_x1_sg U4925 ( .A(n3663), .B(om_max[7]), .X(n2017) );
  nand_x1_sg U4926 ( .A(n3708), .B(om_max[15]), .X(n1998) );
  inv_x1_sg U4927 ( .A(om_min[4]), .X(n3614) );
  nand_x1_sg U4928 ( .A(n3724), .B(om_min[19]), .X(n1309) );
  nand_x1_sg U4929 ( .A(n3642), .B(om_max[3]), .X(n2032) );
  nand_x1_sg U4930 ( .A(n3686), .B(om_max[11]), .X(n2116) );
  inv_x1_sg U4931 ( .A(om_min[1]), .X(n3616) );
  nand_x1_sg U4932 ( .A(n3624), .B(om_min[0]), .X(n1386) );
  inv_x1_sg U4933 ( .A(om_min[0]), .X(n3604) );
  inv_x1_sg U4934 ( .A(om_max[1]), .X(n3623) );
  nor_x1_sg U4935 ( .A(n1971), .B(n2819), .X(n1870) );
  nor_x1_sg U4936 ( .A(n1307), .B(n2818), .X(n1207) );
  nand_x1_sg U4937 ( .A(n3720), .B(om_min[18]), .X(n1313) );
  nand_x1_sg U4938 ( .A(om_min[12]), .B(n1432), .X(n1431) );
  nand_x1_sg U4939 ( .A(n2121), .B(om_max[9]), .X(n2120) );
  nand_x1_sg U4940 ( .A(n1907), .B(n2119), .X(n2121) );
  nand_x1_sg U4941 ( .A(om_max[1]), .B(n2045), .X(n2044) );
  nand_x1_sg U4942 ( .A(n2046), .B(n1968), .X(n2045) );
  nor_x1_sg U4943 ( .A(n2012), .B(n2013), .X(n2010) );
  nor_x1_sg U4944 ( .A(om_max[7]), .B(n3663), .X(n2012) );
  nor_x1_sg U4945 ( .A(n1993), .B(n1994), .X(n1984) );
  nand_x4_sg U4946 ( .A(n1995), .B(n1996), .X(n1994) );
  nor_x1_sg U4947 ( .A(om_max[15]), .B(n3708), .X(n1993) );
  nand_x4_sg U4948 ( .A(n1999), .B(n2000), .X(n1995) );
  nand_x1_sg U4949 ( .A(n3647), .B(om_min[5]), .X(n1359) );
  nand_x1_sg U4950 ( .A(n3715), .B(om_min[17]), .X(n1318) );
  nand_x1_sg U4951 ( .A(\max_pooling_0/N4 ), .B(\max_pooling_0/N3 ), .X(n1965)
         );
  nand_x1_sg U4952 ( .A(\min_pooling_0/N4 ), .B(\min_pooling_0/N3 ), .X(n1301)
         );
  nand_x1_sg U4953 ( .A(\mean_pooling_0/N5 ), .B(\mean_pooling_0/N4 ), .X(
        n1684) );
  nand_x1_sg U4954 ( .A(n3727), .B(om_max[19]), .X(n1975) );
  nor_x1_sg U4955 ( .A(n1321), .B(n1322), .X(n1319) );
  nor_x1_sg U4956 ( .A(n1330), .B(n1331), .X(n1321) );
  nor_x1_sg U4957 ( .A(n3710), .B(\min_pooling_0/n722 ), .X(n1322) );
  nor_x1_sg U4958 ( .A(n2033), .B(n2034), .X(n2029) );
  nor_x1_sg U4959 ( .A(n2035), .B(n2036), .X(n2034) );
  nor_x1_sg U4960 ( .A(om_max[3]), .B(n3642), .X(n2033) );
  nor_x1_sg U4961 ( .A(n1115), .B(n3011), .X(n1151) );
  nor_x1_sg U4962 ( .A(n1370), .B(n3194), .X(n1369) );
  nor_x1_sg U4963 ( .A(om_min[3]), .B(n3638), .X(n1370) );
  nor_x1_sg U4964 ( .A(n1348), .B(n1349), .X(n1346) );
  nor_x1_sg U4965 ( .A(n1350), .B(n1351), .X(n1348) );
  nor_x1_sg U4966 ( .A(om_min[8]), .B(n3665), .X(n1349) );
  nor_x1_sg U4967 ( .A(n1982), .B(n1983), .X(n1980) );
  nor_x1_sg U4968 ( .A(n1984), .B(n1985), .X(n1982) );
  nor_x1_sg U4969 ( .A(om_max[16]), .B(n3714), .X(n1983) );
  nor_x1_sg U4970 ( .A(n3618), .B(n1942), .X(n1985) );
  nand_x1_sg U4971 ( .A(n3652), .B(om_max[5]), .X(n2027) );
  nand_x1_sg U4972 ( .A(n3630), .B(n2822), .X(n1668) );
  nand_x1_sg U4973 ( .A(n1096), .B(n1670), .X(n1669) );
  nand_x1_sg U4974 ( .A(n1097), .B(n3636), .X(n1660) );
  nand_x1_sg U4975 ( .A(n1661), .B(n2826), .X(n1659) );
  nand_x1_sg U4976 ( .A(n3713), .B(n2827), .X(n1533) );
  nand_x1_sg U4977 ( .A(n1111), .B(n1535), .X(n1534) );
  inv_x1_sg U4978 ( .A(n1535), .X(n3713) );
  nand_x1_sg U4979 ( .A(n3707), .B(n2828), .X(n1542) );
  nand_x1_sg U4980 ( .A(n1110), .B(n1544), .X(n1543) );
  inv_x1_sg U4981 ( .A(n1544), .X(n3707) );
  nand_x1_sg U4982 ( .A(n3702), .B(n2829), .X(n1551) );
  nand_x1_sg U4983 ( .A(n1109), .B(n1553), .X(n1552) );
  inv_x1_sg U4984 ( .A(n1553), .X(n3702) );
  nand_x1_sg U4985 ( .A(n3696), .B(n2830), .X(n1560) );
  nand_x1_sg U4986 ( .A(n1108), .B(n1562), .X(n1561) );
  inv_x1_sg U4987 ( .A(n1562), .X(n3696) );
  nand_x1_sg U4988 ( .A(n3691), .B(n2831), .X(n1569) );
  nand_x1_sg U4989 ( .A(n1107), .B(n1571), .X(n1570) );
  inv_x1_sg U4990 ( .A(n1571), .X(n3691) );
  nand_x1_sg U4991 ( .A(n3685), .B(n2832), .X(n1578) );
  nand_x1_sg U4992 ( .A(n1106), .B(n1580), .X(n1579) );
  inv_x1_sg U4993 ( .A(n1580), .X(n3685) );
  nand_x1_sg U4994 ( .A(n3680), .B(n2833), .X(n1587) );
  nand_x1_sg U4995 ( .A(n1105), .B(n1589), .X(n1588) );
  inv_x1_sg U4996 ( .A(n1589), .X(n3680) );
  nand_x1_sg U4997 ( .A(n3674), .B(n2834), .X(n1596) );
  nand_x1_sg U4998 ( .A(n1104), .B(n1598), .X(n1597) );
  inv_x1_sg U4999 ( .A(n1598), .X(n3674) );
  nand_x1_sg U5000 ( .A(n3668), .B(n2835), .X(n1605) );
  nand_x1_sg U5001 ( .A(n1103), .B(n1607), .X(n1606) );
  inv_x1_sg U5002 ( .A(n1607), .X(n3668) );
  nand_x1_sg U5003 ( .A(n3662), .B(n2836), .X(n1614) );
  nand_x1_sg U5004 ( .A(n1102), .B(n1616), .X(n1615) );
  inv_x1_sg U5005 ( .A(n1616), .X(n3662) );
  nand_x1_sg U5006 ( .A(n3657), .B(n2837), .X(n1623) );
  nand_x1_sg U5007 ( .A(n1101), .B(n1625), .X(n1624) );
  inv_x1_sg U5008 ( .A(n1625), .X(n3657) );
  nand_x1_sg U5009 ( .A(n3651), .B(n2838), .X(n1632) );
  nand_x1_sg U5010 ( .A(n1100), .B(n1634), .X(n1633) );
  inv_x1_sg U5011 ( .A(n1634), .X(n3651) );
  nand_x1_sg U5012 ( .A(n3646), .B(n2839), .X(n1641) );
  nand_x1_sg U5013 ( .A(n1099), .B(n1643), .X(n1642) );
  inv_x1_sg U5014 ( .A(n1643), .X(n3646) );
  nand_x1_sg U5015 ( .A(n3641), .B(n2840), .X(n1650) );
  nand_x1_sg U5016 ( .A(n1098), .B(n1652), .X(n1651) );
  inv_x1_sg U5017 ( .A(n1652), .X(n3641) );
  nand_x1_sg U5018 ( .A(n3718), .B(n2823), .X(n1524) );
  nand_x1_sg U5019 ( .A(n1112), .B(n1526), .X(n1525) );
  inv_x1_sg U5020 ( .A(n1743), .X(n3628) );
  nand_x1_sg U5021 ( .A(om_max[18]), .B(n3166), .X(n1139) );
  nand_x1_sg U5022 ( .A(n2902), .B(n2847), .X(n1138) );
  nor_x1_sg U5023 ( .A(\max_pooling_0/n640 ), .B(n3681), .X(n2134) );
  nand_x1_sg U5024 ( .A(om_min[19]), .B(n2847), .X(n1142) );
  nand_x1_sg U5025 ( .A(om_max[19]), .B(n3167), .X(n1143) );
  nand_x1_sg U5026 ( .A(n2016), .B(n2017), .X(n2015) );
  nor_x1_sg U5027 ( .A(\max_pooling_0/n642 ), .B(n3658), .X(n2016) );
  nand_x1_sg U5028 ( .A(n1997), .B(n1998), .X(n1996) );
  nor_x1_sg U5029 ( .A(om_max[14]), .B(n3703), .X(n1997) );
  nand_x1_sg U5030 ( .A(om_mean[5]), .B(n3245), .X(n1169) );
  nor_x1_sg U5031 ( .A(n1170), .B(n1171), .X(n1168) );
  nor_x1_sg U5032 ( .A(n3010), .B(n3118), .X(n1171) );
  nand_x1_sg U5033 ( .A(om_mean[17]), .B(n3130), .X(n1135) );
  nor_x1_sg U5034 ( .A(n1136), .B(n1137), .X(n1134) );
  nor_x1_sg U5035 ( .A(n2870), .B(n3117), .X(n1137) );
  nand_x1_sg U5036 ( .A(om_mean[12]), .B(n3130), .X(n1197) );
  nor_x1_sg U5037 ( .A(n1198), .B(n1199), .X(n1196) );
  nor_x1_sg U5038 ( .A(n3009), .B(n3608), .X(n1199) );
  nand_x1_sg U5039 ( .A(n2037), .B(n2032), .X(n2036) );
  nand_x1_sg U5040 ( .A(n3637), .B(om_max[2]), .X(n2037) );
  nand_x1_sg U5041 ( .A(om_mean[16]), .B(n3130), .X(n1131) );
  nor_x1_sg U5042 ( .A(n1132), .B(n1133), .X(n1130) );
  nor_x1_sg U5043 ( .A(n3177), .B(n3618), .X(n1132) );
  nand_x1_sg U5044 ( .A(om_mean[14]), .B(n2946), .X(n1123) );
  nor_x1_sg U5045 ( .A(n1124), .B(n1125), .X(n1122) );
  nor_x1_sg U5046 ( .A(n3134), .B(n3619), .X(n1124) );
  nand_x1_sg U5047 ( .A(om_mean[13]), .B(n2846), .X(n1119) );
  nor_x1_sg U5048 ( .A(n1120), .B(n1121), .X(n1118) );
  nor_x1_sg U5049 ( .A(n3139), .B(n3620), .X(n1120) );
  nand_x1_sg U5050 ( .A(om_mean[8]), .B(n2946), .X(n1181) );
  nor_x1_sg U5051 ( .A(n1182), .B(n1183), .X(n1180) );
  nor_x1_sg U5052 ( .A(n3147), .B(n3621), .X(n1182) );
  nand_x1_sg U5053 ( .A(om_mean[6]), .B(n3136), .X(n1173) );
  nor_x1_sg U5054 ( .A(n1174), .B(n1175), .X(n1172) );
  nor_x1_sg U5055 ( .A(n3158), .B(n3622), .X(n1174) );
  nand_x1_sg U5056 ( .A(om_mean[15]), .B(n3136), .X(n1127) );
  nor_x1_sg U5057 ( .A(n1128), .B(n1129), .X(n1126) );
  nor_x1_sg U5058 ( .A(n3134), .B(n3120), .X(n1128) );
  nand_x1_sg U5059 ( .A(om_mean[11]), .B(n2946), .X(n1193) );
  nor_x1_sg U5060 ( .A(n1194), .B(n1195), .X(n1192) );
  nor_x1_sg U5061 ( .A(n3196), .B(n3121), .X(n1194) );
  nand_x1_sg U5062 ( .A(om_mean[10]), .B(n3245), .X(n1189) );
  nor_x1_sg U5063 ( .A(n1190), .B(n1191), .X(n1188) );
  nor_x1_sg U5064 ( .A(n3164), .B(n3122), .X(n1190) );
  nand_x1_sg U5065 ( .A(om_mean[7]), .B(n3136), .X(n1177) );
  nor_x1_sg U5066 ( .A(n1178), .B(n1179), .X(n1176) );
  nor_x1_sg U5067 ( .A(n3135), .B(n3124), .X(n1178) );
  nand_x1_sg U5068 ( .A(om_mean[3]), .B(n3244), .X(n1161) );
  nor_x1_sg U5069 ( .A(n1162), .B(n1163), .X(n1160) );
  nor_x1_sg U5070 ( .A(n3149), .B(n3125), .X(n1162) );
  nand_x1_sg U5071 ( .A(om_mean[2]), .B(n3244), .X(n1157) );
  nor_x1_sg U5072 ( .A(n1158), .B(n1159), .X(n1156) );
  nor_x1_sg U5073 ( .A(n3164), .B(n3126), .X(n1158) );
  nand_x1_sg U5074 ( .A(om_mean[9]), .B(n3244), .X(n1185) );
  nor_x1_sg U5075 ( .A(n1186), .B(n1187), .X(n1184) );
  nor_x1_sg U5076 ( .A(n3253), .B(n3123), .X(n1186) );
  nand_x1_sg U5077 ( .A(om_mean[4]), .B(n3136), .X(n1165) );
  nor_x1_sg U5078 ( .A(n1166), .B(n1167), .X(n1164) );
  nor_x1_sg U5079 ( .A(n3158), .B(n3150), .X(n1166) );
  nand_x1_sg U5080 ( .A(om_mean[0]), .B(n3244), .X(n1202) );
  nor_x1_sg U5081 ( .A(n1203), .B(n1204), .X(n1201) );
  nor_x1_sg U5082 ( .A(n3253), .B(n3151), .X(n1203) );
  nand_x1_sg U5083 ( .A(om_mean[1]), .B(n2946), .X(n1153) );
  nor_x1_sg U5084 ( .A(n1154), .B(n1155), .X(n1152) );
  nor_x1_sg U5085 ( .A(n3164), .B(n3623), .X(n1154) );
  nand_x1_sg U5086 ( .A(n3130), .B(n2841), .X(n1149) );
  nor_x1_sg U5087 ( .A(n1150), .B(n1151), .X(n1148) );
  nor_x1_sg U5088 ( .A(n1116), .B(n3158), .X(n1150) );
  nor_x1_sg U5089 ( .A(n2010), .B(n2011), .X(n2008) );
  nand_x1_sg U5090 ( .A(n3675), .B(om_max[9]), .X(n2009) );
  nor_x1_sg U5091 ( .A(n3621), .B(n1902), .X(n2011) );
  nand_x1_sg U5092 ( .A(n2116), .B(n2117), .X(n2115) );
  nand_x1_sg U5093 ( .A(n3681), .B(\max_pooling_0/n640 ), .X(n2117) );
  nor_x1_sg U5094 ( .A(n2818), .B(n3069), .X(\min_pooling_0/n314 ) );
  nor_x1_sg U5095 ( .A(n2820), .B(n3073), .X(\mean_pooling_0/n168 ) );
  nor_x1_sg U5096 ( .A(n2819), .B(n2914), .X(\max_pooling_0/n233 ) );
  nor_x1_sg U5097 ( .A(n2818), .B(n3067), .X(\min_pooling_0/n313 ) );
  nor_x1_sg U5098 ( .A(n2820), .B(n3071), .X(\mean_pooling_0/n167 ) );
  nor_x1_sg U5099 ( .A(n2819), .B(n3063), .X(\max_pooling_0/n232 ) );
  nand_x1_sg U5100 ( .A(n3091), .B(n1258), .X(n1256) );
  nand_x1_sg U5101 ( .A(n3089), .B(om_min[12]), .X(n1257) );
  nand_x1_sg U5102 ( .A(n2953), .B(n1298), .X(n1296) );
  nand_x1_sg U5103 ( .A(n2932), .B(om_min[0]), .X(n1297) );
  nand_x1_sg U5104 ( .A(n3079), .B(n1968), .X(n1966) );
  nand_x1_sg U5105 ( .A(n2890), .B(om_max[1]), .X(n1967) );
  nand_x1_sg U5106 ( .A(n3078), .B(n1887), .X(n1885) );
  nand_x1_sg U5107 ( .A(n3083), .B(om_max[5]), .X(n1886) );
  nand_x1_sg U5108 ( .A(n2887), .B(n1952), .X(n1950) );
  nand_x1_sg U5109 ( .A(n3082), .B(om_max[18]), .X(n1951) );
  nand_x1_sg U5110 ( .A(n3091), .B(n1213), .X(n1211) );
  nand_x1_sg U5111 ( .A(n3087), .B(om_min[3]), .X(n1212) );
  nand_x1_sg U5112 ( .A(n2953), .B(n1228), .X(n1226) );
  nand_x1_sg U5113 ( .A(n3086), .B(om_min[6]), .X(n1227) );
  nand_x1_sg U5114 ( .A(n3092), .B(n1233), .X(n1231) );
  nand_x1_sg U5115 ( .A(n3086), .B(om_min[7]), .X(n1232) );
  nand_x1_sg U5116 ( .A(n2935), .B(n1238), .X(n1236) );
  nand_x1_sg U5117 ( .A(n2892), .B(om_min[8]), .X(n1237) );
  nand_x1_sg U5118 ( .A(n3093), .B(n1248), .X(n1246) );
  nand_x1_sg U5119 ( .A(n2893), .B(om_min[10]), .X(n1247) );
  nand_x1_sg U5120 ( .A(n2954), .B(n1253), .X(n1251) );
  nand_x1_sg U5121 ( .A(n3087), .B(om_min[11]), .X(n1252) );
  nand_x1_sg U5122 ( .A(n2896), .B(n1268), .X(n1266) );
  nand_x1_sg U5123 ( .A(n2892), .B(\min_pooling_0/n723 ), .X(n1267) );
  nand_x1_sg U5124 ( .A(n2935), .B(n1273), .X(n1271) );
  nand_x1_sg U5125 ( .A(n2892), .B(om_min[15]), .X(n1272) );
  nand_x1_sg U5126 ( .A(n2895), .B(n1278), .X(n1276) );
  nand_x1_sg U5127 ( .A(n3088), .B(\min_pooling_0/n722 ), .X(n1277) );
  nand_x1_sg U5128 ( .A(n3076), .B(n1882), .X(n1880) );
  nand_x1_sg U5129 ( .A(n2929), .B(\max_pooling_0/n643 ), .X(n1881) );
  nand_x1_sg U5130 ( .A(n3077), .B(n1892), .X(n1890) );
  nand_x1_sg U5131 ( .A(n2929), .B(\max_pooling_0/n642 ), .X(n1891) );
  nand_x1_sg U5132 ( .A(n2927), .B(n1902), .X(n1900) );
  nand_x1_sg U5133 ( .A(n2889), .B(\max_pooling_0/n641 ), .X(n1901) );
  nand_x1_sg U5134 ( .A(n3078), .B(n1927), .X(n1925) );
  nand_x1_sg U5135 ( .A(n2950), .B(om_max[13]), .X(n1926) );
  nand_x1_sg U5136 ( .A(n3076), .B(n1932), .X(n1930) );
  nand_x1_sg U5137 ( .A(n3082), .B(om_max[14]), .X(n1931) );
  nand_x1_sg U5138 ( .A(n2886), .B(n1942), .X(n1940) );
  nand_x1_sg U5139 ( .A(n3084), .B(om_max[16]), .X(n1941) );
  nand_x1_sg U5140 ( .A(n3078), .B(n1962), .X(n1960) );
  nand_x1_sg U5141 ( .A(n2929), .B(om_max[0]), .X(n1961) );
  nand_x1_sg U5142 ( .A(n2954), .B(n1293), .X(n1291) );
  nand_x1_sg U5143 ( .A(n2952), .B(om_min[19]), .X(n1292) );
  nand_x1_sg U5144 ( .A(n3077), .B(n1907), .X(n1905) );
  nand_x1_sg U5145 ( .A(n2950), .B(om_max[9]), .X(n1906) );
  nand_x1_sg U5146 ( .A(n2948), .B(n1957), .X(n1955) );
  nand_x1_sg U5147 ( .A(n2890), .B(om_max[19]), .X(n1956) );
  nand_x1_sg U5148 ( .A(n3092), .B(n1223), .X(n1221) );
  nand_x1_sg U5149 ( .A(n3088), .B(om_min[5]), .X(n1222) );
  nand_x1_sg U5150 ( .A(n3090), .B(n1283), .X(n1281) );
  nand_x1_sg U5151 ( .A(n2932), .B(om_min[17]), .X(n1282) );
  nand_x1_sg U5152 ( .A(n3079), .B(n1872), .X(n1868) );
  nand_x1_sg U5153 ( .A(n2890), .B(om_max[2]), .X(n1869) );
  nand_x1_sg U5154 ( .A(n3077), .B(n1877), .X(n1875) );
  nand_x1_sg U5155 ( .A(n3083), .B(om_max[3]), .X(n1876) );
  nand_x1_sg U5156 ( .A(n2887), .B(n1897), .X(n1895) );
  nand_x1_sg U5157 ( .A(n2930), .B(om_max[7]), .X(n1896) );
  nand_x1_sg U5158 ( .A(n2886), .B(n1912), .X(n1910) );
  nand_x1_sg U5159 ( .A(n2889), .B(\max_pooling_0/n640 ), .X(n1911) );
  nand_x1_sg U5160 ( .A(n2887), .B(n1917), .X(n1915) );
  nand_x1_sg U5161 ( .A(n2949), .B(om_max[11]), .X(n1916) );
  nand_x1_sg U5162 ( .A(n2947), .B(n1937), .X(n1935) );
  nand_x1_sg U5163 ( .A(n2889), .B(om_max[15]), .X(n1936) );
  nand_x1_sg U5164 ( .A(n2896), .B(n1288), .X(n1286) );
  nand_x1_sg U5165 ( .A(n3088), .B(n2902), .X(n1287) );
  nand_x1_sg U5166 ( .A(n3089), .B(om_min[1]), .X(n1303) );
  nand_x1_sg U5167 ( .A(n2936), .B(n1304), .X(n1302) );
  nand_x1_sg U5168 ( .A(n2893), .B(\min_pooling_0/n724 ), .X(n1206) );
  nand_x1_sg U5169 ( .A(n2896), .B(n1208), .X(n1205) );
  nand_x1_sg U5170 ( .A(n2951), .B(om_min[4]), .X(n1217) );
  nand_x1_sg U5171 ( .A(n2895), .B(n1218), .X(n1216) );
  nand_x1_sg U5172 ( .A(n2951), .B(om_min[9]), .X(n1242) );
  nand_x1_sg U5173 ( .A(n3093), .B(n1243), .X(n1241) );
  nand_x1_sg U5174 ( .A(n3089), .B(om_min[13]), .X(n1262) );
  nand_x1_sg U5175 ( .A(n3092), .B(n1263), .X(n1261) );
  nand_x1_sg U5176 ( .A(n2927), .B(n1922), .X(n1920) );
  nand_x1_sg U5177 ( .A(n3083), .B(\max_pooling_0/n639 ), .X(n1921) );
  nand_x1_sg U5178 ( .A(n3077), .B(n1947), .X(n1945) );
  nand_x1_sg U5179 ( .A(n3081), .B(om_max[17]), .X(n1946) );
  nand_x1_sg U5180 ( .A(n2933), .B(n3127), .X(n1290) );
  nand_x1_sg U5181 ( .A(n2935), .B(n3720), .X(n1289) );
  inv_x16_sg U5182 ( .A(n1140), .X(n3253) );
endmodule

