
module transposer ( clk, reset, input_ready, output_taken, state, .in({
        \in[3][3][19] , \in[3][3][18] , \in[3][3][17] , \in[3][3][16] , 
        \in[3][3][15] , \in[3][3][14] , \in[3][3][13] , \in[3][3][12] , 
        \in[3][3][11] , \in[3][3][10] , \in[3][3][9] , \in[3][3][8] , 
        \in[3][3][7] , \in[3][3][6] , \in[3][3][5] , \in[3][3][4] , 
        \in[3][3][3] , \in[3][3][2] , \in[3][3][1] , \in[3][3][0] , 
        \in[3][2][19] , \in[3][2][18] , \in[3][2][17] , \in[3][2][16] , 
        \in[3][2][15] , \in[3][2][14] , \in[3][2][13] , \in[3][2][12] , 
        \in[3][2][11] , \in[3][2][10] , \in[3][2][9] , \in[3][2][8] , 
        \in[3][2][7] , \in[3][2][6] , \in[3][2][5] , \in[3][2][4] , 
        \in[3][2][3] , \in[3][2][2] , \in[3][2][1] , \in[3][2][0] , 
        \in[3][1][19] , \in[3][1][18] , \in[3][1][17] , \in[3][1][16] , 
        \in[3][1][15] , \in[3][1][14] , \in[3][1][13] , \in[3][1][12] , 
        \in[3][1][11] , \in[3][1][10] , \in[3][1][9] , \in[3][1][8] , 
        \in[3][1][7] , \in[3][1][6] , \in[3][1][5] , \in[3][1][4] , 
        \in[3][1][3] , \in[3][1][2] , \in[3][1][1] , \in[3][1][0] , 
        \in[3][0][19] , \in[3][0][18] , \in[3][0][17] , \in[3][0][16] , 
        \in[3][0][15] , \in[3][0][14] , \in[3][0][13] , \in[3][0][12] , 
        \in[3][0][11] , \in[3][0][10] , \in[3][0][9] , \in[3][0][8] , 
        \in[3][0][7] , \in[3][0][6] , \in[3][0][5] , \in[3][0][4] , 
        \in[3][0][3] , \in[3][0][2] , \in[3][0][1] , \in[3][0][0] , 
        \in[2][3][19] , \in[2][3][18] , \in[2][3][17] , \in[2][3][16] , 
        \in[2][3][15] , \in[2][3][14] , \in[2][3][13] , \in[2][3][12] , 
        \in[2][3][11] , \in[2][3][10] , \in[2][3][9] , \in[2][3][8] , 
        \in[2][3][7] , \in[2][3][6] , \in[2][3][5] , \in[2][3][4] , 
        \in[2][3][3] , \in[2][3][2] , \in[2][3][1] , \in[2][3][0] , 
        \in[2][2][19] , \in[2][2][18] , \in[2][2][17] , \in[2][2][16] , 
        \in[2][2][15] , \in[2][2][14] , \in[2][2][13] , \in[2][2][12] , 
        \in[2][2][11] , \in[2][2][10] , \in[2][2][9] , \in[2][2][8] , 
        \in[2][2][7] , \in[2][2][6] , \in[2][2][5] , \in[2][2][4] , 
        \in[2][2][3] , \in[2][2][2] , \in[2][2][1] , \in[2][2][0] , 
        \in[2][1][19] , \in[2][1][18] , \in[2][1][17] , \in[2][1][16] , 
        \in[2][1][15] , \in[2][1][14] , \in[2][1][13] , \in[2][1][12] , 
        \in[2][1][11] , \in[2][1][10] , \in[2][1][9] , \in[2][1][8] , 
        \in[2][1][7] , \in[2][1][6] , \in[2][1][5] , \in[2][1][4] , 
        \in[2][1][3] , \in[2][1][2] , \in[2][1][1] , \in[2][1][0] , 
        \in[2][0][19] , \in[2][0][18] , \in[2][0][17] , \in[2][0][16] , 
        \in[2][0][15] , \in[2][0][14] , \in[2][0][13] , \in[2][0][12] , 
        \in[2][0][11] , \in[2][0][10] , \in[2][0][9] , \in[2][0][8] , 
        \in[2][0][7] , \in[2][0][6] , \in[2][0][5] , \in[2][0][4] , 
        \in[2][0][3] , \in[2][0][2] , \in[2][0][1] , \in[2][0][0] , 
        \in[1][3][19] , \in[1][3][18] , \in[1][3][17] , \in[1][3][16] , 
        \in[1][3][15] , \in[1][3][14] , \in[1][3][13] , \in[1][3][12] , 
        \in[1][3][11] , \in[1][3][10] , \in[1][3][9] , \in[1][3][8] , 
        \in[1][3][7] , \in[1][3][6] , \in[1][3][5] , \in[1][3][4] , 
        \in[1][3][3] , \in[1][3][2] , \in[1][3][1] , \in[1][3][0] , 
        \in[1][2][19] , \in[1][2][18] , \in[1][2][17] , \in[1][2][16] , 
        \in[1][2][15] , \in[1][2][14] , \in[1][2][13] , \in[1][2][12] , 
        \in[1][2][11] , \in[1][2][10] , \in[1][2][9] , \in[1][2][8] , 
        \in[1][2][7] , \in[1][2][6] , \in[1][2][5] , \in[1][2][4] , 
        \in[1][2][3] , \in[1][2][2] , \in[1][2][1] , \in[1][2][0] , 
        \in[1][1][19] , \in[1][1][18] , \in[1][1][17] , \in[1][1][16] , 
        \in[1][1][15] , \in[1][1][14] , \in[1][1][13] , \in[1][1][12] , 
        \in[1][1][11] , \in[1][1][10] , \in[1][1][9] , \in[1][1][8] , 
        \in[1][1][7] , \in[1][1][6] , \in[1][1][5] , \in[1][1][4] , 
        \in[1][1][3] , \in[1][1][2] , \in[1][1][1] , \in[1][1][0] , 
        \in[1][0][19] , \in[1][0][18] , \in[1][0][17] , \in[1][0][16] , 
        \in[1][0][15] , \in[1][0][14] , \in[1][0][13] , \in[1][0][12] , 
        \in[1][0][11] , \in[1][0][10] , \in[1][0][9] , \in[1][0][8] , 
        \in[1][0][7] , \in[1][0][6] , \in[1][0][5] , \in[1][0][4] , 
        \in[1][0][3] , \in[1][0][2] , \in[1][0][1] , \in[1][0][0] , 
        \in[0][3][19] , \in[0][3][18] , \in[0][3][17] , \in[0][3][16] , 
        \in[0][3][15] , \in[0][3][14] , \in[0][3][13] , \in[0][3][12] , 
        \in[0][3][11] , \in[0][3][10] , \in[0][3][9] , \in[0][3][8] , 
        \in[0][3][7] , \in[0][3][6] , \in[0][3][5] , \in[0][3][4] , 
        \in[0][3][3] , \in[0][3][2] , \in[0][3][1] , \in[0][3][0] , 
        \in[0][2][19] , \in[0][2][18] , \in[0][2][17] , \in[0][2][16] , 
        \in[0][2][15] , \in[0][2][14] , \in[0][2][13] , \in[0][2][12] , 
        \in[0][2][11] , \in[0][2][10] , \in[0][2][9] , \in[0][2][8] , 
        \in[0][2][7] , \in[0][2][6] , \in[0][2][5] , \in[0][2][4] , 
        \in[0][2][3] , \in[0][2][2] , \in[0][2][1] , \in[0][2][0] , 
        \in[0][1][19] , \in[0][1][18] , \in[0][1][17] , \in[0][1][16] , 
        \in[0][1][15] , \in[0][1][14] , \in[0][1][13] , \in[0][1][12] , 
        \in[0][1][11] , \in[0][1][10] , \in[0][1][9] , \in[0][1][8] , 
        \in[0][1][7] , \in[0][1][6] , \in[0][1][5] , \in[0][1][4] , 
        \in[0][1][3] , \in[0][1][2] , \in[0][1][1] , \in[0][1][0] , 
        \in[0][0][19] , \in[0][0][18] , \in[0][0][17] , \in[0][0][16] , 
        \in[0][0][15] , \in[0][0][14] , \in[0][0][13] , \in[0][0][12] , 
        \in[0][0][11] , \in[0][0][10] , \in[0][0][9] , \in[0][0][8] , 
        \in[0][0][7] , \in[0][0][6] , \in[0][0][5] , \in[0][0][4] , 
        \in[0][0][3] , \in[0][0][2] , \in[0][0][1] , \in[0][0][0] }), .out({
        \out[3][3][19] , \out[3][3][18] , \out[3][3][17] , \out[3][3][16] , 
        \out[3][3][15] , \out[3][3][14] , \out[3][3][13] , \out[3][3][12] , 
        \out[3][3][11] , \out[3][3][10] , \out[3][3][9] , \out[3][3][8] , 
        \out[3][3][7] , \out[3][3][6] , \out[3][3][5] , \out[3][3][4] , 
        \out[3][3][3] , \out[3][3][2] , \out[3][3][1] , \out[3][3][0] , 
        \out[3][2][19] , \out[3][2][18] , \out[3][2][17] , \out[3][2][16] , 
        \out[3][2][15] , \out[3][2][14] , \out[3][2][13] , \out[3][2][12] , 
        \out[3][2][11] , \out[3][2][10] , \out[3][2][9] , \out[3][2][8] , 
        \out[3][2][7] , \out[3][2][6] , \out[3][2][5] , \out[3][2][4] , 
        \out[3][2][3] , \out[3][2][2] , \out[3][2][1] , \out[3][2][0] , 
        \out[3][1][19] , \out[3][1][18] , \out[3][1][17] , \out[3][1][16] , 
        \out[3][1][15] , \out[3][1][14] , \out[3][1][13] , \out[3][1][12] , 
        \out[3][1][11] , \out[3][1][10] , \out[3][1][9] , \out[3][1][8] , 
        \out[3][1][7] , \out[3][1][6] , \out[3][1][5] , \out[3][1][4] , 
        \out[3][1][3] , \out[3][1][2] , \out[3][1][1] , \out[3][1][0] , 
        \out[3][0][19] , \out[3][0][18] , \out[3][0][17] , \out[3][0][16] , 
        \out[3][0][15] , \out[3][0][14] , \out[3][0][13] , \out[3][0][12] , 
        \out[3][0][11] , \out[3][0][10] , \out[3][0][9] , \out[3][0][8] , 
        \out[3][0][7] , \out[3][0][6] , \out[3][0][5] , \out[3][0][4] , 
        \out[3][0][3] , \out[3][0][2] , \out[3][0][1] , \out[3][0][0] , 
        \out[2][3][19] , \out[2][3][18] , \out[2][3][17] , \out[2][3][16] , 
        \out[2][3][15] , \out[2][3][14] , \out[2][3][13] , \out[2][3][12] , 
        \out[2][3][11] , \out[2][3][10] , \out[2][3][9] , \out[2][3][8] , 
        \out[2][3][7] , \out[2][3][6] , \out[2][3][5] , \out[2][3][4] , 
        \out[2][3][3] , \out[2][3][2] , \out[2][3][1] , \out[2][3][0] , 
        \out[2][2][19] , \out[2][2][18] , \out[2][2][17] , \out[2][2][16] , 
        \out[2][2][15] , \out[2][2][14] , \out[2][2][13] , \out[2][2][12] , 
        \out[2][2][11] , \out[2][2][10] , \out[2][2][9] , \out[2][2][8] , 
        \out[2][2][7] , \out[2][2][6] , \out[2][2][5] , \out[2][2][4] , 
        \out[2][2][3] , \out[2][2][2] , \out[2][2][1] , \out[2][2][0] , 
        \out[2][1][19] , \out[2][1][18] , \out[2][1][17] , \out[2][1][16] , 
        \out[2][1][15] , \out[2][1][14] , \out[2][1][13] , \out[2][1][12] , 
        \out[2][1][11] , \out[2][1][10] , \out[2][1][9] , \out[2][1][8] , 
        \out[2][1][7] , \out[2][1][6] , \out[2][1][5] , \out[2][1][4] , 
        \out[2][1][3] , \out[2][1][2] , \out[2][1][1] , \out[2][1][0] , 
        \out[2][0][19] , \out[2][0][18] , \out[2][0][17] , \out[2][0][16] , 
        \out[2][0][15] , \out[2][0][14] , \out[2][0][13] , \out[2][0][12] , 
        \out[2][0][11] , \out[2][0][10] , \out[2][0][9] , \out[2][0][8] , 
        \out[2][0][7] , \out[2][0][6] , \out[2][0][5] , \out[2][0][4] , 
        \out[2][0][3] , \out[2][0][2] , \out[2][0][1] , \out[2][0][0] , 
        \out[1][3][19] , \out[1][3][18] , \out[1][3][17] , \out[1][3][16] , 
        \out[1][3][15] , \out[1][3][14] , \out[1][3][13] , \out[1][3][12] , 
        \out[1][3][11] , \out[1][3][10] , \out[1][3][9] , \out[1][3][8] , 
        \out[1][3][7] , \out[1][3][6] , \out[1][3][5] , \out[1][3][4] , 
        \out[1][3][3] , \out[1][3][2] , \out[1][3][1] , \out[1][3][0] , 
        \out[1][2][19] , \out[1][2][18] , \out[1][2][17] , \out[1][2][16] , 
        \out[1][2][15] , \out[1][2][14] , \out[1][2][13] , \out[1][2][12] , 
        \out[1][2][11] , \out[1][2][10] , \out[1][2][9] , \out[1][2][8] , 
        \out[1][2][7] , \out[1][2][6] , \out[1][2][5] , \out[1][2][4] , 
        \out[1][2][3] , \out[1][2][2] , \out[1][2][1] , \out[1][2][0] , 
        \out[1][1][19] , \out[1][1][18] , \out[1][1][17] , \out[1][1][16] , 
        \out[1][1][15] , \out[1][1][14] , \out[1][1][13] , \out[1][1][12] , 
        \out[1][1][11] , \out[1][1][10] , \out[1][1][9] , \out[1][1][8] , 
        \out[1][1][7] , \out[1][1][6] , \out[1][1][5] , \out[1][1][4] , 
        \out[1][1][3] , \out[1][1][2] , \out[1][1][1] , \out[1][1][0] , 
        \out[1][0][19] , \out[1][0][18] , \out[1][0][17] , \out[1][0][16] , 
        \out[1][0][15] , \out[1][0][14] , \out[1][0][13] , \out[1][0][12] , 
        \out[1][0][11] , \out[1][0][10] , \out[1][0][9] , \out[1][0][8] , 
        \out[1][0][7] , \out[1][0][6] , \out[1][0][5] , \out[1][0][4] , 
        \out[1][0][3] , \out[1][0][2] , \out[1][0][1] , \out[1][0][0] , 
        \out[0][3][19] , \out[0][3][18] , \out[0][3][17] , \out[0][3][16] , 
        \out[0][3][15] , \out[0][3][14] , \out[0][3][13] , \out[0][3][12] , 
        \out[0][3][11] , \out[0][3][10] , \out[0][3][9] , \out[0][3][8] , 
        \out[0][3][7] , \out[0][3][6] , \out[0][3][5] , \out[0][3][4] , 
        \out[0][3][3] , \out[0][3][2] , \out[0][3][1] , \out[0][3][0] , 
        \out[0][2][19] , \out[0][2][18] , \out[0][2][17] , \out[0][2][16] , 
        \out[0][2][15] , \out[0][2][14] , \out[0][2][13] , \out[0][2][12] , 
        \out[0][2][11] , \out[0][2][10] , \out[0][2][9] , \out[0][2][8] , 
        \out[0][2][7] , \out[0][2][6] , \out[0][2][5] , \out[0][2][4] , 
        \out[0][2][3] , \out[0][2][2] , \out[0][2][1] , \out[0][2][0] , 
        \out[0][1][19] , \out[0][1][18] , \out[0][1][17] , \out[0][1][16] , 
        \out[0][1][15] , \out[0][1][14] , \out[0][1][13] , \out[0][1][12] , 
        \out[0][1][11] , \out[0][1][10] , \out[0][1][9] , \out[0][1][8] , 
        \out[0][1][7] , \out[0][1][6] , \out[0][1][5] , \out[0][1][4] , 
        \out[0][1][3] , \out[0][1][2] , \out[0][1][1] , \out[0][1][0] , 
        \out[0][0][19] , \out[0][0][18] , \out[0][0][17] , \out[0][0][16] , 
        \out[0][0][15] , \out[0][0][14] , \out[0][0][13] , \out[0][0][12] , 
        \out[0][0][11] , \out[0][0][10] , \out[0][0][9] , \out[0][0][8] , 
        \out[0][0][7] , \out[0][0][6] , \out[0][0][5] , \out[0][0][4] , 
        \out[0][0][3] , \out[0][0][2] , \out[0][0][1] , \out[0][0][0] }) );
  output [1:0] state;
  input clk, reset, input_ready, output_taken, \in[3][3][19] , \in[3][3][18] ,
         \in[3][3][17] , \in[3][3][16] , \in[3][3][15] , \in[3][3][14] ,
         \in[3][3][13] , \in[3][3][12] , \in[3][3][11] , \in[3][3][10] ,
         \in[3][3][9] , \in[3][3][8] , \in[3][3][7] , \in[3][3][6] ,
         \in[3][3][5] , \in[3][3][4] , \in[3][3][3] , \in[3][3][2] ,
         \in[3][3][1] , \in[3][3][0] , \in[3][2][19] , \in[3][2][18] ,
         \in[3][2][17] , \in[3][2][16] , \in[3][2][15] , \in[3][2][14] ,
         \in[3][2][13] , \in[3][2][12] , \in[3][2][11] , \in[3][2][10] ,
         \in[3][2][9] , \in[3][2][8] , \in[3][2][7] , \in[3][2][6] ,
         \in[3][2][5] , \in[3][2][4] , \in[3][2][3] , \in[3][2][2] ,
         \in[3][2][1] , \in[3][2][0] , \in[3][1][19] , \in[3][1][18] ,
         \in[3][1][17] , \in[3][1][16] , \in[3][1][15] , \in[3][1][14] ,
         \in[3][1][13] , \in[3][1][12] , \in[3][1][11] , \in[3][1][10] ,
         \in[3][1][9] , \in[3][1][8] , \in[3][1][7] , \in[3][1][6] ,
         \in[3][1][5] , \in[3][1][4] , \in[3][1][3] , \in[3][1][2] ,
         \in[3][1][1] , \in[3][1][0] , \in[3][0][19] , \in[3][0][18] ,
         \in[3][0][17] , \in[3][0][16] , \in[3][0][15] , \in[3][0][14] ,
         \in[3][0][13] , \in[3][0][12] , \in[3][0][11] , \in[3][0][10] ,
         \in[3][0][9] , \in[3][0][8] , \in[3][0][7] , \in[3][0][6] ,
         \in[3][0][5] , \in[3][0][4] , \in[3][0][3] , \in[3][0][2] ,
         \in[3][0][1] , \in[3][0][0] , \in[2][3][19] , \in[2][3][18] ,
         \in[2][3][17] , \in[2][3][16] , \in[2][3][15] , \in[2][3][14] ,
         \in[2][3][13] , \in[2][3][12] , \in[2][3][11] , \in[2][3][10] ,
         \in[2][3][9] , \in[2][3][8] , \in[2][3][7] , \in[2][3][6] ,
         \in[2][3][5] , \in[2][3][4] , \in[2][3][3] , \in[2][3][2] ,
         \in[2][3][1] , \in[2][3][0] , \in[2][2][19] , \in[2][2][18] ,
         \in[2][2][17] , \in[2][2][16] , \in[2][2][15] , \in[2][2][14] ,
         \in[2][2][13] , \in[2][2][12] , \in[2][2][11] , \in[2][2][10] ,
         \in[2][2][9] , \in[2][2][8] , \in[2][2][7] , \in[2][2][6] ,
         \in[2][2][5] , \in[2][2][4] , \in[2][2][3] , \in[2][2][2] ,
         \in[2][2][1] , \in[2][2][0] , \in[2][1][19] , \in[2][1][18] ,
         \in[2][1][17] , \in[2][1][16] , \in[2][1][15] , \in[2][1][14] ,
         \in[2][1][13] , \in[2][1][12] , \in[2][1][11] , \in[2][1][10] ,
         \in[2][1][9] , \in[2][1][8] , \in[2][1][7] , \in[2][1][6] ,
         \in[2][1][5] , \in[2][1][4] , \in[2][1][3] , \in[2][1][2] ,
         \in[2][1][1] , \in[2][1][0] , \in[2][0][19] , \in[2][0][18] ,
         \in[2][0][17] , \in[2][0][16] , \in[2][0][15] , \in[2][0][14] ,
         \in[2][0][13] , \in[2][0][12] , \in[2][0][11] , \in[2][0][10] ,
         \in[2][0][9] , \in[2][0][8] , \in[2][0][7] , \in[2][0][6] ,
         \in[2][0][5] , \in[2][0][4] , \in[2][0][3] , \in[2][0][2] ,
         \in[2][0][1] , \in[2][0][0] , \in[1][3][19] , \in[1][3][18] ,
         \in[1][3][17] , \in[1][3][16] , \in[1][3][15] , \in[1][3][14] ,
         \in[1][3][13] , \in[1][3][12] , \in[1][3][11] , \in[1][3][10] ,
         \in[1][3][9] , \in[1][3][8] , \in[1][3][7] , \in[1][3][6] ,
         \in[1][3][5] , \in[1][3][4] , \in[1][3][3] , \in[1][3][2] ,
         \in[1][3][1] , \in[1][3][0] , \in[1][2][19] , \in[1][2][18] ,
         \in[1][2][17] , \in[1][2][16] , \in[1][2][15] , \in[1][2][14] ,
         \in[1][2][13] , \in[1][2][12] , \in[1][2][11] , \in[1][2][10] ,
         \in[1][2][9] , \in[1][2][8] , \in[1][2][7] , \in[1][2][6] ,
         \in[1][2][5] , \in[1][2][4] , \in[1][2][3] , \in[1][2][2] ,
         \in[1][2][1] , \in[1][2][0] , \in[1][1][19] , \in[1][1][18] ,
         \in[1][1][17] , \in[1][1][16] , \in[1][1][15] , \in[1][1][14] ,
         \in[1][1][13] , \in[1][1][12] , \in[1][1][11] , \in[1][1][10] ,
         \in[1][1][9] , \in[1][1][8] , \in[1][1][7] , \in[1][1][6] ,
         \in[1][1][5] , \in[1][1][4] , \in[1][1][3] , \in[1][1][2] ,
         \in[1][1][1] , \in[1][1][0] , \in[1][0][19] , \in[1][0][18] ,
         \in[1][0][17] , \in[1][0][16] , \in[1][0][15] , \in[1][0][14] ,
         \in[1][0][13] , \in[1][0][12] , \in[1][0][11] , \in[1][0][10] ,
         \in[1][0][9] , \in[1][0][8] , \in[1][0][7] , \in[1][0][6] ,
         \in[1][0][5] , \in[1][0][4] , \in[1][0][3] , \in[1][0][2] ,
         \in[1][0][1] , \in[1][0][0] , \in[0][3][19] , \in[0][3][18] ,
         \in[0][3][17] , \in[0][3][16] , \in[0][3][15] , \in[0][3][14] ,
         \in[0][3][13] , \in[0][3][12] , \in[0][3][11] , \in[0][3][10] ,
         \in[0][3][9] , \in[0][3][8] , \in[0][3][7] , \in[0][3][6] ,
         \in[0][3][5] , \in[0][3][4] , \in[0][3][3] , \in[0][3][2] ,
         \in[0][3][1] , \in[0][3][0] , \in[0][2][19] , \in[0][2][18] ,
         \in[0][2][17] , \in[0][2][16] , \in[0][2][15] , \in[0][2][14] ,
         \in[0][2][13] , \in[0][2][12] , \in[0][2][11] , \in[0][2][10] ,
         \in[0][2][9] , \in[0][2][8] , \in[0][2][7] , \in[0][2][6] ,
         \in[0][2][5] , \in[0][2][4] , \in[0][2][3] , \in[0][2][2] ,
         \in[0][2][1] , \in[0][2][0] , \in[0][1][19] , \in[0][1][18] ,
         \in[0][1][17] , \in[0][1][16] , \in[0][1][15] , \in[0][1][14] ,
         \in[0][1][13] , \in[0][1][12] , \in[0][1][11] , \in[0][1][10] ,
         \in[0][1][9] , \in[0][1][8] , \in[0][1][7] , \in[0][1][6] ,
         \in[0][1][5] , \in[0][1][4] , \in[0][1][3] , \in[0][1][2] ,
         \in[0][1][1] , \in[0][1][0] , \in[0][0][19] , \in[0][0][18] ,
         \in[0][0][17] , \in[0][0][16] , \in[0][0][15] , \in[0][0][14] ,
         \in[0][0][13] , \in[0][0][12] , \in[0][0][11] , \in[0][0][10] ,
         \in[0][0][9] , \in[0][0][8] , \in[0][0][7] , \in[0][0][6] ,
         \in[0][0][5] , \in[0][0][4] , \in[0][0][3] , \in[0][0][2] ,
         \in[0][0][1] , \in[0][0][0] ;
  output \out[3][3][19] , \out[3][3][18] , \out[3][3][17] , \out[3][3][16] ,
         \out[3][3][15] , \out[3][3][14] , \out[3][3][13] , \out[3][3][12] ,
         \out[3][3][11] , \out[3][3][10] , \out[3][3][9] , \out[3][3][8] ,
         \out[3][3][7] , \out[3][3][6] , \out[3][3][5] , \out[3][3][4] ,
         \out[3][3][3] , \out[3][3][2] , \out[3][3][1] , \out[3][3][0] ,
         \out[3][2][19] , \out[3][2][18] , \out[3][2][17] , \out[3][2][16] ,
         \out[3][2][15] , \out[3][2][14] , \out[3][2][13] , \out[3][2][12] ,
         \out[3][2][11] , \out[3][2][10] , \out[3][2][9] , \out[3][2][8] ,
         \out[3][2][7] , \out[3][2][6] , \out[3][2][5] , \out[3][2][4] ,
         \out[3][2][3] , \out[3][2][2] , \out[3][2][1] , \out[3][2][0] ,
         \out[3][1][19] , \out[3][1][18] , \out[3][1][17] , \out[3][1][16] ,
         \out[3][1][15] , \out[3][1][14] , \out[3][1][13] , \out[3][1][12] ,
         \out[3][1][11] , \out[3][1][10] , \out[3][1][9] , \out[3][1][8] ,
         \out[3][1][7] , \out[3][1][6] , \out[3][1][5] , \out[3][1][4] ,
         \out[3][1][3] , \out[3][1][2] , \out[3][1][1] , \out[3][1][0] ,
         \out[3][0][19] , \out[3][0][18] , \out[3][0][17] , \out[3][0][16] ,
         \out[3][0][15] , \out[3][0][14] , \out[3][0][13] , \out[3][0][12] ,
         \out[3][0][11] , \out[3][0][10] , \out[3][0][9] , \out[3][0][8] ,
         \out[3][0][7] , \out[3][0][6] , \out[3][0][5] , \out[3][0][4] ,
         \out[3][0][3] , \out[3][0][2] , \out[3][0][1] , \out[3][0][0] ,
         \out[2][3][19] , \out[2][3][18] , \out[2][3][17] , \out[2][3][16] ,
         \out[2][3][15] , \out[2][3][14] , \out[2][3][13] , \out[2][3][12] ,
         \out[2][3][11] , \out[2][3][10] , \out[2][3][9] , \out[2][3][8] ,
         \out[2][3][7] , \out[2][3][6] , \out[2][3][5] , \out[2][3][4] ,
         \out[2][3][3] , \out[2][3][2] , \out[2][3][1] , \out[2][3][0] ,
         \out[2][2][19] , \out[2][2][18] , \out[2][2][17] , \out[2][2][16] ,
         \out[2][2][15] , \out[2][2][14] , \out[2][2][13] , \out[2][2][12] ,
         \out[2][2][11] , \out[2][2][10] , \out[2][2][9] , \out[2][2][8] ,
         \out[2][2][7] , \out[2][2][6] , \out[2][2][5] , \out[2][2][4] ,
         \out[2][2][3] , \out[2][2][2] , \out[2][2][1] , \out[2][2][0] ,
         \out[2][1][19] , \out[2][1][18] , \out[2][1][17] , \out[2][1][16] ,
         \out[2][1][15] , \out[2][1][14] , \out[2][1][13] , \out[2][1][12] ,
         \out[2][1][11] , \out[2][1][10] , \out[2][1][9] , \out[2][1][8] ,
         \out[2][1][7] , \out[2][1][6] , \out[2][1][5] , \out[2][1][4] ,
         \out[2][1][3] , \out[2][1][2] , \out[2][1][1] , \out[2][1][0] ,
         \out[2][0][19] , \out[2][0][18] , \out[2][0][17] , \out[2][0][16] ,
         \out[2][0][15] , \out[2][0][14] , \out[2][0][13] , \out[2][0][12] ,
         \out[2][0][11] , \out[2][0][10] , \out[2][0][9] , \out[2][0][8] ,
         \out[2][0][7] , \out[2][0][6] , \out[2][0][5] , \out[2][0][4] ,
         \out[2][0][3] , \out[2][0][2] , \out[2][0][1] , \out[2][0][0] ,
         \out[1][3][19] , \out[1][3][18] , \out[1][3][17] , \out[1][3][16] ,
         \out[1][3][15] , \out[1][3][14] , \out[1][3][13] , \out[1][3][12] ,
         \out[1][3][11] , \out[1][3][10] , \out[1][3][9] , \out[1][3][8] ,
         \out[1][3][7] , \out[1][3][6] , \out[1][3][5] , \out[1][3][4] ,
         \out[1][3][3] , \out[1][3][2] , \out[1][3][1] , \out[1][3][0] ,
         \out[1][2][19] , \out[1][2][18] , \out[1][2][17] , \out[1][2][16] ,
         \out[1][2][15] , \out[1][2][14] , \out[1][2][13] , \out[1][2][12] ,
         \out[1][2][11] , \out[1][2][10] , \out[1][2][9] , \out[1][2][8] ,
         \out[1][2][7] , \out[1][2][6] , \out[1][2][5] , \out[1][2][4] ,
         \out[1][2][3] , \out[1][2][2] , \out[1][2][1] , \out[1][2][0] ,
         \out[1][1][19] , \out[1][1][18] , \out[1][1][17] , \out[1][1][16] ,
         \out[1][1][15] , \out[1][1][14] , \out[1][1][13] , \out[1][1][12] ,
         \out[1][1][11] , \out[1][1][10] , \out[1][1][9] , \out[1][1][8] ,
         \out[1][1][7] , \out[1][1][6] , \out[1][1][5] , \out[1][1][4] ,
         \out[1][1][3] , \out[1][1][2] , \out[1][1][1] , \out[1][1][0] ,
         \out[1][0][19] , \out[1][0][18] , \out[1][0][17] , \out[1][0][16] ,
         \out[1][0][15] , \out[1][0][14] , \out[1][0][13] , \out[1][0][12] ,
         \out[1][0][11] , \out[1][0][10] , \out[1][0][9] , \out[1][0][8] ,
         \out[1][0][7] , \out[1][0][6] , \out[1][0][5] , \out[1][0][4] ,
         \out[1][0][3] , \out[1][0][2] , \out[1][0][1] , \out[1][0][0] ,
         \out[0][3][19] , \out[0][3][18] , \out[0][3][17] , \out[0][3][16] ,
         \out[0][3][15] , \out[0][3][14] , \out[0][3][13] , \out[0][3][12] ,
         \out[0][3][11] , \out[0][3][10] , \out[0][3][9] , \out[0][3][8] ,
         \out[0][3][7] , \out[0][3][6] , \out[0][3][5] , \out[0][3][4] ,
         \out[0][3][3] , \out[0][3][2] , \out[0][3][1] , \out[0][3][0] ,
         \out[0][2][19] , \out[0][2][18] , \out[0][2][17] , \out[0][2][16] ,
         \out[0][2][15] , \out[0][2][14] , \out[0][2][13] , \out[0][2][12] ,
         \out[0][2][11] , \out[0][2][10] , \out[0][2][9] , \out[0][2][8] ,
         \out[0][2][7] , \out[0][2][6] , \out[0][2][5] , \out[0][2][4] ,
         \out[0][2][3] , \out[0][2][2] , \out[0][2][1] , \out[0][2][0] ,
         \out[0][1][19] , \out[0][1][18] , \out[0][1][17] , \out[0][1][16] ,
         \out[0][1][15] , \out[0][1][14] , \out[0][1][13] , \out[0][1][12] ,
         \out[0][1][11] , \out[0][1][10] , \out[0][1][9] , \out[0][1][8] ,
         \out[0][1][7] , \out[0][1][6] , \out[0][1][5] , \out[0][1][4] ,
         \out[0][1][3] , \out[0][1][2] , \out[0][1][1] , \out[0][1][0] ,
         \out[0][0][19] , \out[0][0][18] , \out[0][0][17] , \out[0][0][16] ,
         \out[0][0][15] , \out[0][0][14] , \out[0][0][13] , \out[0][0][12] ,
         \out[0][0][11] , \out[0][0][10] , \out[0][0][9] , \out[0][0][8] ,
         \out[0][0][7] , \out[0][0][6] , \out[0][0][5] , \out[0][0][4] ,
         \out[0][0][3] , \out[0][0][2] , \out[0][0][1] , \out[0][0][0] ;
  wire   \reg_in[3][3][19] , \reg_in[3][3][18] , \reg_in[3][3][17] ,
         \reg_in[3][3][16] , \reg_in[3][3][15] , \reg_in[3][3][14] ,
         \reg_in[3][3][13] , \reg_in[3][3][12] , \reg_in[3][3][11] ,
         \reg_in[3][3][10] , \reg_in[3][3][9] , \reg_in[3][3][8] ,
         \reg_in[3][3][7] , \reg_in[3][3][6] , \reg_in[3][3][5] ,
         \reg_in[3][3][4] , \reg_in[3][3][3] , \reg_in[3][3][2] ,
         \reg_in[3][3][1] , \reg_in[3][3][0] , \reg_in[3][2][19] ,
         \reg_in[3][2][18] , \reg_in[3][2][17] , \reg_in[3][2][16] ,
         \reg_in[3][2][15] , \reg_in[3][2][14] , \reg_in[3][2][13] ,
         \reg_in[3][2][12] , \reg_in[3][2][11] , \reg_in[3][2][10] ,
         \reg_in[3][2][9] , \reg_in[3][2][8] , \reg_in[3][2][7] ,
         \reg_in[3][2][6] , \reg_in[3][2][5] , \reg_in[3][2][4] ,
         \reg_in[3][2][3] , \reg_in[3][2][2] , \reg_in[3][2][1] ,
         \reg_in[3][2][0] , \reg_in[3][1][19] , \reg_in[3][1][18] ,
         \reg_in[3][1][17] , \reg_in[3][1][16] , \reg_in[3][1][15] ,
         \reg_in[3][1][14] , \reg_in[3][1][13] , \reg_in[3][1][12] ,
         \reg_in[3][1][11] , \reg_in[3][1][10] , \reg_in[3][1][9] ,
         \reg_in[3][1][8] , \reg_in[3][1][7] , \reg_in[3][1][6] ,
         \reg_in[3][1][5] , \reg_in[3][1][4] , \reg_in[3][1][3] ,
         \reg_in[3][1][2] , \reg_in[3][1][1] , \reg_in[3][1][0] ,
         \reg_in[3][0][19] , \reg_in[3][0][18] , \reg_in[3][0][17] ,
         \reg_in[3][0][16] , \reg_in[3][0][15] , \reg_in[3][0][14] ,
         \reg_in[3][0][13] , \reg_in[3][0][12] , \reg_in[3][0][11] ,
         \reg_in[3][0][10] , \reg_in[3][0][9] , \reg_in[3][0][8] ,
         \reg_in[3][0][7] , \reg_in[3][0][6] , \reg_in[3][0][5] ,
         \reg_in[3][0][4] , \reg_in[3][0][3] , \reg_in[3][0][2] ,
         \reg_in[3][0][1] , \reg_in[3][0][0] , \reg_in[2][3][19] ,
         \reg_in[2][3][18] , \reg_in[2][3][17] , \reg_in[2][3][16] ,
         \reg_in[2][3][15] , \reg_in[2][3][14] , \reg_in[2][3][13] ,
         \reg_in[2][3][12] , \reg_in[2][3][11] , \reg_in[2][3][10] ,
         \reg_in[2][3][9] , \reg_in[2][3][8] , \reg_in[2][3][7] ,
         \reg_in[2][3][6] , \reg_in[2][3][5] , \reg_in[2][3][4] ,
         \reg_in[2][3][3] , \reg_in[2][3][2] , \reg_in[2][3][1] ,
         \reg_in[2][3][0] , \reg_in[2][2][19] , \reg_in[2][2][18] ,
         \reg_in[2][2][17] , \reg_in[2][2][16] , \reg_in[2][2][15] ,
         \reg_in[2][2][14] , \reg_in[2][2][13] , \reg_in[2][2][12] ,
         \reg_in[2][2][11] , \reg_in[2][2][10] , \reg_in[2][2][9] ,
         \reg_in[2][2][8] , \reg_in[2][2][7] , \reg_in[2][2][6] ,
         \reg_in[2][2][5] , \reg_in[2][2][4] , \reg_in[2][2][3] ,
         \reg_in[2][2][2] , \reg_in[2][2][1] , \reg_in[2][2][0] ,
         \reg_in[2][1][19] , \reg_in[2][1][18] , \reg_in[2][1][17] ,
         \reg_in[2][1][16] , \reg_in[2][1][15] , \reg_in[2][1][14] ,
         \reg_in[2][1][13] , \reg_in[2][1][12] , \reg_in[2][1][11] ,
         \reg_in[2][1][10] , \reg_in[2][1][9] , \reg_in[2][1][8] ,
         \reg_in[2][1][7] , \reg_in[2][1][6] , \reg_in[2][1][5] ,
         \reg_in[2][1][4] , \reg_in[2][1][3] , \reg_in[2][1][2] ,
         \reg_in[2][1][1] , \reg_in[2][1][0] , \reg_in[2][0][19] ,
         \reg_in[2][0][18] , \reg_in[2][0][17] , \reg_in[2][0][16] ,
         \reg_in[2][0][15] , \reg_in[2][0][14] , \reg_in[2][0][13] ,
         \reg_in[2][0][12] , \reg_in[2][0][11] , \reg_in[2][0][10] ,
         \reg_in[2][0][9] , \reg_in[2][0][8] , \reg_in[2][0][7] ,
         \reg_in[2][0][6] , \reg_in[2][0][5] , \reg_in[2][0][4] ,
         \reg_in[2][0][3] , \reg_in[2][0][2] , \reg_in[2][0][1] ,
         \reg_in[2][0][0] , \reg_in[1][3][19] , \reg_in[1][3][18] ,
         \reg_in[1][3][17] , \reg_in[1][3][16] , \reg_in[1][3][15] ,
         \reg_in[1][3][14] , \reg_in[1][3][13] , \reg_in[1][3][12] ,
         \reg_in[1][3][11] , \reg_in[1][3][10] , \reg_in[1][3][9] ,
         \reg_in[1][3][8] , \reg_in[1][3][7] , \reg_in[1][3][6] ,
         \reg_in[1][3][5] , \reg_in[1][3][4] , \reg_in[1][3][3] ,
         \reg_in[1][3][2] , \reg_in[1][3][1] , \reg_in[1][3][0] ,
         \reg_in[1][2][19] , \reg_in[1][2][18] , \reg_in[1][2][17] ,
         \reg_in[1][2][16] , \reg_in[1][2][15] , \reg_in[1][2][14] ,
         \reg_in[1][2][13] , \reg_in[1][2][12] , \reg_in[1][2][11] ,
         \reg_in[1][2][10] , \reg_in[1][2][9] , \reg_in[1][2][8] ,
         \reg_in[1][2][7] , \reg_in[1][2][6] , \reg_in[1][2][5] ,
         \reg_in[1][2][4] , \reg_in[1][2][3] , \reg_in[1][2][2] ,
         \reg_in[1][2][1] , \reg_in[1][2][0] , \reg_in[1][1][19] ,
         \reg_in[1][1][18] , \reg_in[1][1][17] , \reg_in[1][1][16] ,
         \reg_in[1][1][15] , \reg_in[1][1][14] , \reg_in[1][1][13] ,
         \reg_in[1][1][12] , \reg_in[1][1][11] , \reg_in[1][1][10] ,
         \reg_in[1][1][9] , \reg_in[1][1][8] , \reg_in[1][1][7] ,
         \reg_in[1][1][6] , \reg_in[1][1][5] , \reg_in[1][1][4] ,
         \reg_in[1][1][3] , \reg_in[1][1][2] , \reg_in[1][1][1] ,
         \reg_in[1][1][0] , \reg_in[1][0][19] , \reg_in[1][0][18] ,
         \reg_in[1][0][17] , \reg_in[1][0][16] , \reg_in[1][0][15] ,
         \reg_in[1][0][14] , \reg_in[1][0][13] , \reg_in[1][0][12] ,
         \reg_in[1][0][11] , \reg_in[1][0][10] , \reg_in[1][0][9] ,
         \reg_in[1][0][8] , \reg_in[1][0][7] , \reg_in[1][0][6] ,
         \reg_in[1][0][5] , \reg_in[1][0][4] , \reg_in[1][0][3] ,
         \reg_in[1][0][2] , \reg_in[1][0][1] , \reg_in[1][0][0] ,
         \reg_in[0][3][19] , \reg_in[0][3][18] , \reg_in[0][3][17] ,
         \reg_in[0][3][16] , \reg_in[0][3][15] , \reg_in[0][3][14] ,
         \reg_in[0][3][13] , \reg_in[0][3][12] , \reg_in[0][3][11] ,
         \reg_in[0][3][10] , \reg_in[0][3][9] , \reg_in[0][3][8] ,
         \reg_in[0][3][7] , \reg_in[0][3][6] , \reg_in[0][3][5] ,
         \reg_in[0][3][4] , \reg_in[0][3][3] , \reg_in[0][3][2] ,
         \reg_in[0][3][1] , \reg_in[0][3][0] , \reg_in[0][2][19] ,
         \reg_in[0][2][18] , \reg_in[0][2][17] , \reg_in[0][2][16] ,
         \reg_in[0][2][15] , \reg_in[0][2][14] , \reg_in[0][2][13] ,
         \reg_in[0][2][12] , \reg_in[0][2][11] , \reg_in[0][2][10] ,
         \reg_in[0][2][9] , \reg_in[0][2][8] , \reg_in[0][2][7] ,
         \reg_in[0][2][6] , \reg_in[0][2][5] , \reg_in[0][2][4] ,
         \reg_in[0][2][3] , \reg_in[0][2][2] , \reg_in[0][2][1] ,
         \reg_in[0][2][0] , \reg_in[0][1][19] , \reg_in[0][1][18] ,
         \reg_in[0][1][17] , \reg_in[0][1][16] , \reg_in[0][1][15] ,
         \reg_in[0][1][14] , \reg_in[0][1][13] , \reg_in[0][1][12] ,
         \reg_in[0][1][11] , \reg_in[0][1][10] , \reg_in[0][1][9] ,
         \reg_in[0][1][8] , \reg_in[0][1][7] , \reg_in[0][1][6] ,
         \reg_in[0][1][5] , \reg_in[0][1][4] , \reg_in[0][1][3] ,
         \reg_in[0][1][2] , \reg_in[0][1][1] , \reg_in[0][1][0] ,
         \reg_in[0][0][19] , \reg_in[0][0][18] , \reg_in[0][0][17] ,
         \reg_in[0][0][16] , \reg_in[0][0][15] , \reg_in[0][0][14] ,
         \reg_in[0][0][13] , \reg_in[0][0][12] , \reg_in[0][0][11] ,
         \reg_in[0][0][10] , \reg_in[0][0][9] , \reg_in[0][0][8] ,
         \reg_in[0][0][7] , \reg_in[0][0][6] , \reg_in[0][0][5] ,
         \reg_in[0][0][4] , \reg_in[0][0][3] , \reg_in[0][0][2] ,
         \reg_in[0][0][1] , \reg_in[0][0][0] , n3546, n3547, n3548, n3549,
         n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559,
         n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569,
         n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579,
         n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589,
         n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599,
         n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609,
         n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619,
         n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629,
         n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639,
         n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649,
         n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659,
         n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669,
         n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679,
         n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689,
         n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699,
         n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709,
         n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719,
         n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729,
         n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739,
         n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749,
         n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759,
         n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769,
         n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779,
         n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789,
         n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799,
         n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809,
         n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819,
         n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829,
         n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839,
         n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849,
         n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859,
         n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869,
         n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879,
         n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889,
         n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899,
         n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909,
         n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919,
         n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929,
         n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939,
         n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949,
         n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959,
         n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969,
         n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979,
         n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989,
         n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999,
         n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009,
         n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019,
         n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029,
         n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039,
         n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049,
         n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059,
         n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069,
         n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079,
         n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089,
         n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099,
         n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109,
         n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119,
         n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129,
         n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139,
         n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149,
         n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159,
         n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169,
         n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179,
         n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189,
         n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199,
         n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209,
         n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219,
         n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229,
         n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239,
         n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249,
         n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259,
         n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269,
         n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279,
         n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289,
         n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299,
         n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309,
         n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319,
         n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329,
         n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339,
         n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349,
         n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359,
         n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369,
         n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379,
         n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389,
         n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399,
         n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409,
         n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419,
         n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429,
         n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439,
         n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449,
         n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459,
         n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469,
         n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479,
         n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489,
         n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499,
         n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n8707, n8708,
         n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718,
         n8719, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729,
         n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739,
         n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749,
         n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759,
         n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769,
         n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779,
         n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789,
         n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799,
         n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809,
         n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819,
         n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829,
         n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839,
         n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849,
         n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859,
         n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869,
         n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879,
         n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889,
         n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899,
         n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909,
         n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919,
         n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929,
         n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939,
         n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949,
         n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959,
         n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969,
         n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979,
         n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989,
         n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999,
         n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009,
         n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019,
         n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029,
         n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039,
         n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049,
         n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059,
         n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069,
         n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079,
         n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089,
         n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099,
         n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109,
         n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119,
         n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129,
         n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139,
         n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149,
         n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159,
         n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169,
         n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179,
         n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189,
         n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199,
         n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209,
         n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219,
         n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229,
         n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239,
         n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249,
         n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259,
         n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269,
         n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279,
         n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289,
         n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299,
         n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309,
         n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319,
         n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329,
         n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339,
         n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349,
         n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359,
         n9360, n9361, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370,
         n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380,
         n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390,
         n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400,
         n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410,
         n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420,
         n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430,
         n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440,
         n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450,
         n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460,
         n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470,
         n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480,
         n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490,
         n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500,
         n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510,
         n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520,
         n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530,
         n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540,
         n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550,
         n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560,
         n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570,
         n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580,
         n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590,
         n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600,
         n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610,
         n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620,
         n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630,
         n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640,
         n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650,
         n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660,
         n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670,
         n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680,
         n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690,
         n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700,
         n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710,
         n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720,
         n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730,
         n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740,
         n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750,
         n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760,
         n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770,
         n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780,
         n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790,
         n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800,
         n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810,
         n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820,
         n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830,
         n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840,
         n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850,
         n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860,
         n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870,
         n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880,
         n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890,
         n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900,
         n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910,
         n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920,
         n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930,
         n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940,
         n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950,
         n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960,
         n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970,
         n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980,
         n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990,
         n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n8381, n8380, n8379, n8378, n8377, n8376, n8375,
         n8374, n8373, n8372, n8371, n8370, n8369, n8368, n8367, n8366, n8365,
         n8364, n8363, n8362, n8361, n8360, n8359, n8358, n8357, n8356, n8355,
         n8354, n8353, n8352, n8351, n8350, n8349, n8348, n8347, n8346, n8345,
         n8344, n8343, n8342, n8341, n8340, n8339, n8338, n8337, n8336, n8335,
         n8334, n8333, n8332, n8331, n8330, n8329, n8328, n8327, n8326, n8325,
         n8324, n8323, n8322, n8321, n8320, n8319, n8318, n8317, n8316, n8315,
         n8314, n8313, n8312, n8311, n8310, n8309, n8308, n8307, n8306, n8305,
         n8304, n8303, n8302, n8301, n8300, n8299, n8298, n8297, n8296, n8295,
         n8294, n8293, n8292, n8291, n8290, n8289, n8288, n8287, n8286, n8285,
         n8284, n8283, n8282, n8281, n8280, n8279, n8278, n8277, n8276, n8275,
         n8274, n8273, n8272, n8271, n8270, n8269, n8268, n8267, n8266, n8265,
         n8264, n8263, n8262, n8261, n8260, n8259, n8258, n8257, n8256, n8255,
         n8254, n8253, n8252, n8251, n8250, n8249, n8248, n8247, n8246, n8245,
         n8244, n8243, n8242, n8241, n8240, n8239, n8238, n8237, n8236, n8235,
         n8234, n8233, n8232, n8231, n8230, n8229, n8228, n8227, n8226, n8225,
         n8224, n8223, n8222, n8221, n8220, n8219, n8218, n8217, n8216, n8215,
         n8214, n8213, n8212, n8211, n8210, n8209, n8208, n8207, n8206, n8205,
         n8204, n8203, n8202, n8201, n8200, n8199, n8198, n8197, n8196, n8195,
         n8194, n8193, n8192, n8191, n8190, n8189, n8188, n8187, n8186, n8185,
         n8184, n8183, n8182, n8181, n8180, n8179, n8178, n8177, n8176, n8175,
         n8174, n8173, n8172, n8171, n8170, n8169, n8168, n8167, n8166, n8165,
         n8164, n8163, n8162, n8161, n8160, n8159, n8158, n8157, n8156, n8155,
         n8154, n8153, n8152, n8151, n8150, n8149, n8148, n8147, n8146, n8145,
         n8144, n8143, n8142, n8141, n8140, n8139, n8138, n8137, n8136, n8135,
         n8134, n8133, n8132, n8131, n8130, n8129, n8128, n8127, n8126, n8125,
         n8124, n8123, n8122, n8121, n8120, n8119, n8118, n8117, n8116, n8115,
         n8114, n8113, n8112, n8111, n8110, n8109, n8108, n8107, n8106, n8105,
         n8104, n8103, n8102, n8101, n8100, n8099, n8098, n8097, n8096, n8095,
         n8094, n8093, n8092, n8091, n8090, n8089, n8088, n8087, n8086, n8085,
         n8084, n8083, n8082, n8081, n8080, n8079, n8078, n8077, n8076, n8075,
         n8074, n8073, n8072, n8071, n8070, n8069, n8068, n8067, n8066, n8065,
         n8064, n8063, n8062, n3543, n3539, n3535, n3531, n3527, n3523, n3519,
         n3515, n3511, n3507, n3503, n3499, n3495, n3491, n3487, n3483, n3479,
         n3475, n3471, n3467, n3463, n3459, n3455, n3451, n3447, n3443, n3439,
         n3435, n3431, n3427, n3423, n3419, n3415, n3411, n3407, n3403, n3399,
         n3395, n3391, n3387, n3383, n3379, n3375, n3371, n3367, n3363, n3359,
         n3355, n3351, n3347, n3343, n3339, n3335, n3331, n3327, n3323, n3319,
         n3315, n3311, n3307, n3303, n3299, n3295, n3291, n3287, n3283, n3279,
         n3275, n3271, n3267, n3263, n3259, n3255, n3251, n3247, n3243, n3239,
         n3235, n3231, n3227, n3223, n3219, n3215, n3211, n3207, n3203, n3199,
         n3195, n3191, n3187, n3183, n3179, n3175, n3171, n3167, n3163, n3159,
         n3155, n3151, n3147, n3143, n3139, n3135, n3131, n3127, n3123, n3119,
         n3115, n3111, n3107, n3103, n3099, n3095, n3091, n3087, n3083, n3079,
         n3075, n3071, n3067, n3063, n3059, n3055, n3051, n3047, n3043, n3039,
         n3035, n3031, n3027, n3023, n3019, n3015, n3011, n3007, n3003, n2999,
         n2995, n2991, n2987, n2983, n2979, n2975, n2971, n2967, n2963, n2959,
         n2955, n2951, n2947, n2943, n2939, n2935, n2931, n2927, n2923, n2919,
         n2915, n2911, n2907, n2903, n2899, n2895, n2891, n2887, n2883, n2879,
         n2875, n2871, n2867, n2863, n2859, n2855, n2851, n2847, n2843, n2839,
         n2835, n2831, n2827, n2823, n2819, n2815, n2811, n2807, n2803, n2799,
         n2795, n2791, n2787, n2783, n2779, n2775, n2771, n2767, n2763, n2759,
         n2755, n2751, n2747, n2743, n2739, n2735, n2731, n2727, n2723, n2719,
         n2715, n2711, n2707, n2703, n2699, n2695, n2691, n2687, n2683, n2679,
         n2675, n2671, n2667, n2663, n2659, n2655, n2651, n2647, n2643, n2639,
         n2635, n2631, n2627, n2623, n2619, n2615, n2611, n2607, n2603, n2599,
         n2595, n2591, n2587, n2583, n2579, n2575, n2571, n2567, n2563, n2559,
         n2555, n2551, n2547, n2543, n2539, n2535, n2531, n2527, n2523, n2519,
         n2515, n2511, n2507, n2503, n2499, n2495, n2491, n2487, n2483, n2479,
         n2475, n2471, n2467, n2463, n2459, n2455, n2451, n2447, n2443, n2439,
         n2435, n2431, n2427, n2423, n2419, n2415, n2411, n2407, n2403, n2399,
         n2395, n2391, n2387, n2383, n2379, n2375, n2371, n2367, n2363, n2359,
         n2355, n2351, n2347, n2343, n2339, n2335, n2331, n2327, n2323, n2319,
         n2315, n2311, n2307, n2303, n2299, n2295, n2291, n2287, n2283, n2279,
         n2275, n2271, n2267, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
         n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512,
         n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
         n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
         n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536,
         n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
         n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552,
         n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560,
         n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568,
         n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576,
         n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584,
         n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592,
         n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600,
         n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608,
         n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616,
         n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624,
         n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632,
         n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640,
         n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648,
         n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656,
         n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664,
         n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672,
         n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680,
         n10681, n10682, n10683, n10684, n10685, n11966, n11967, n11968,
         n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976,
         n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984,
         n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992,
         n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000,
         n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008,
         n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016,
         n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024,
         n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032,
         n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040,
         n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048,
         n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056,
         n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064,
         n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072,
         n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080,
         n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088,
         n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096,
         n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104,
         n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112,
         n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120,
         n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128,
         n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136,
         n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144,
         n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152,
         n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160,
         n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168,
         n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176,
         n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184,
         n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192,
         n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200,
         n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208,
         n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216,
         n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224,
         n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232,
         n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240,
         n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248,
         n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256,
         n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264,
         n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272,
         n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280,
         n12281, n12282, n12283, n12284, n12285, n12286, n12287;

  dff_sg \state_reg[0]  ( .D(n4507), .CP(clk), .Q(state[0]) );
  dff_sg \state_reg[1]  ( .D(n4506), .CP(clk), .Q(state[1]) );
  dff_sg \reg_in_reg[3][3][19]  ( .D(n4505), .CP(clk), .Q(\reg_in[3][3][19] )
         );
  dff_sg \reg_in_reg[3][3][18]  ( .D(n4504), .CP(clk), .Q(\reg_in[3][3][18] )
         );
  dff_sg \reg_in_reg[3][3][17]  ( .D(n4503), .CP(clk), .Q(\reg_in[3][3][17] )
         );
  dff_sg \reg_in_reg[3][3][16]  ( .D(n4502), .CP(clk), .Q(\reg_in[3][3][16] )
         );
  dff_sg \reg_in_reg[3][3][15]  ( .D(n4501), .CP(clk), .Q(\reg_in[3][3][15] )
         );
  dff_sg \reg_in_reg[3][3][14]  ( .D(n4500), .CP(clk), .Q(\reg_in[3][3][14] )
         );
  dff_sg \reg_in_reg[3][3][13]  ( .D(n4499), .CP(clk), .Q(\reg_in[3][3][13] )
         );
  dff_sg \reg_in_reg[3][3][12]  ( .D(n4498), .CP(clk), .Q(\reg_in[3][3][12] )
         );
  dff_sg \reg_in_reg[3][3][11]  ( .D(n4497), .CP(clk), .Q(\reg_in[3][3][11] )
         );
  dff_sg \reg_in_reg[3][3][10]  ( .D(n4496), .CP(clk), .Q(\reg_in[3][3][10] )
         );
  dff_sg \reg_in_reg[3][3][9]  ( .D(n4495), .CP(clk), .Q(\reg_in[3][3][9] ) );
  dff_sg \reg_in_reg[3][3][8]  ( .D(n4494), .CP(clk), .Q(\reg_in[3][3][8] ) );
  dff_sg \reg_in_reg[3][3][7]  ( .D(n4493), .CP(clk), .Q(\reg_in[3][3][7] ) );
  dff_sg \reg_in_reg[3][3][6]  ( .D(n4492), .CP(clk), .Q(\reg_in[3][3][6] ) );
  dff_sg \reg_in_reg[3][3][5]  ( .D(n4491), .CP(clk), .Q(\reg_in[3][3][5] ) );
  dff_sg \reg_in_reg[3][3][4]  ( .D(n4490), .CP(clk), .Q(\reg_in[3][3][4] ) );
  dff_sg \reg_in_reg[3][3][3]  ( .D(n4489), .CP(clk), .Q(\reg_in[3][3][3] ) );
  dff_sg \reg_in_reg[3][3][2]  ( .D(n4488), .CP(clk), .Q(\reg_in[3][3][2] ) );
  dff_sg \reg_in_reg[3][3][1]  ( .D(n4487), .CP(clk), .Q(\reg_in[3][3][1] ) );
  dff_sg \reg_in_reg[3][3][0]  ( .D(n4486), .CP(clk), .Q(\reg_in[3][3][0] ) );
  dff_sg \reg_in_reg[3][2][19]  ( .D(n4485), .CP(clk), .Q(\reg_in[3][2][19] )
         );
  dff_sg \reg_in_reg[3][2][18]  ( .D(n4484), .CP(clk), .Q(\reg_in[3][2][18] )
         );
  dff_sg \reg_in_reg[3][2][17]  ( .D(n4483), .CP(clk), .Q(\reg_in[3][2][17] )
         );
  dff_sg \reg_in_reg[3][2][16]  ( .D(n4482), .CP(clk), .Q(\reg_in[3][2][16] )
         );
  dff_sg \reg_in_reg[3][2][15]  ( .D(n4481), .CP(clk), .Q(\reg_in[3][2][15] )
         );
  dff_sg \reg_in_reg[3][2][14]  ( .D(n4480), .CP(clk), .Q(\reg_in[3][2][14] )
         );
  dff_sg \reg_in_reg[3][2][13]  ( .D(n4479), .CP(clk), .Q(\reg_in[3][2][13] )
         );
  dff_sg \reg_in_reg[3][2][12]  ( .D(n4478), .CP(clk), .Q(\reg_in[3][2][12] )
         );
  dff_sg \reg_in_reg[3][2][11]  ( .D(n4477), .CP(clk), .Q(\reg_in[3][2][11] )
         );
  dff_sg \reg_in_reg[3][2][10]  ( .D(n4476), .CP(clk), .Q(\reg_in[3][2][10] )
         );
  dff_sg \reg_in_reg[3][2][9]  ( .D(n4475), .CP(clk), .Q(\reg_in[3][2][9] ) );
  dff_sg \reg_in_reg[3][2][8]  ( .D(n4474), .CP(clk), .Q(\reg_in[3][2][8] ) );
  dff_sg \reg_in_reg[3][2][7]  ( .D(n4473), .CP(clk), .Q(\reg_in[3][2][7] ) );
  dff_sg \reg_in_reg[3][2][6]  ( .D(n4472), .CP(clk), .Q(\reg_in[3][2][6] ) );
  dff_sg \reg_in_reg[3][2][5]  ( .D(n4471), .CP(clk), .Q(\reg_in[3][2][5] ) );
  dff_sg \reg_in_reg[3][2][4]  ( .D(n4470), .CP(clk), .Q(\reg_in[3][2][4] ) );
  dff_sg \reg_in_reg[3][2][3]  ( .D(n4469), .CP(clk), .Q(\reg_in[3][2][3] ) );
  dff_sg \reg_in_reg[3][2][2]  ( .D(n4468), .CP(clk), .Q(\reg_in[3][2][2] ) );
  dff_sg \reg_in_reg[3][2][1]  ( .D(n4467), .CP(clk), .Q(\reg_in[3][2][1] ) );
  dff_sg \reg_in_reg[3][2][0]  ( .D(n4466), .CP(clk), .Q(\reg_in[3][2][0] ) );
  dff_sg \reg_in_reg[3][1][19]  ( .D(n4465), .CP(clk), .Q(\reg_in[3][1][19] )
         );
  dff_sg \reg_in_reg[3][1][18]  ( .D(n4464), .CP(clk), .Q(\reg_in[3][1][18] )
         );
  dff_sg \reg_in_reg[3][1][17]  ( .D(n4463), .CP(clk), .Q(\reg_in[3][1][17] )
         );
  dff_sg \reg_in_reg[3][1][16]  ( .D(n4462), .CP(clk), .Q(\reg_in[3][1][16] )
         );
  dff_sg \reg_in_reg[3][1][15]  ( .D(n4461), .CP(clk), .Q(\reg_in[3][1][15] )
         );
  dff_sg \reg_in_reg[3][1][14]  ( .D(n4460), .CP(clk), .Q(\reg_in[3][1][14] )
         );
  dff_sg \reg_in_reg[3][1][13]  ( .D(n4459), .CP(clk), .Q(\reg_in[3][1][13] )
         );
  dff_sg \reg_in_reg[3][1][12]  ( .D(n4458), .CP(clk), .Q(\reg_in[3][1][12] )
         );
  dff_sg \reg_in_reg[3][1][11]  ( .D(n4457), .CP(clk), .Q(\reg_in[3][1][11] )
         );
  dff_sg \reg_in_reg[3][1][10]  ( .D(n4456), .CP(clk), .Q(\reg_in[3][1][10] )
         );
  dff_sg \reg_in_reg[3][1][9]  ( .D(n4455), .CP(clk), .Q(\reg_in[3][1][9] ) );
  dff_sg \reg_in_reg[3][1][8]  ( .D(n4454), .CP(clk), .Q(\reg_in[3][1][8] ) );
  dff_sg \reg_in_reg[3][1][7]  ( .D(n4453), .CP(clk), .Q(\reg_in[3][1][7] ) );
  dff_sg \reg_in_reg[3][1][6]  ( .D(n4452), .CP(clk), .Q(\reg_in[3][1][6] ) );
  dff_sg \reg_in_reg[3][1][5]  ( .D(n4451), .CP(clk), .Q(\reg_in[3][1][5] ) );
  dff_sg \reg_in_reg[3][1][4]  ( .D(n4450), .CP(clk), .Q(\reg_in[3][1][4] ) );
  dff_sg \reg_in_reg[3][1][3]  ( .D(n4449), .CP(clk), .Q(\reg_in[3][1][3] ) );
  dff_sg \reg_in_reg[3][1][2]  ( .D(n4448), .CP(clk), .Q(\reg_in[3][1][2] ) );
  dff_sg \reg_in_reg[3][1][1]  ( .D(n4447), .CP(clk), .Q(\reg_in[3][1][1] ) );
  dff_sg \reg_in_reg[3][1][0]  ( .D(n4446), .CP(clk), .Q(\reg_in[3][1][0] ) );
  dff_sg \reg_in_reg[3][0][19]  ( .D(n4445), .CP(clk), .Q(\reg_in[3][0][19] )
         );
  dff_sg \reg_in_reg[3][0][18]  ( .D(n4444), .CP(clk), .Q(\reg_in[3][0][18] )
         );
  dff_sg \reg_in_reg[3][0][17]  ( .D(n4443), .CP(clk), .Q(\reg_in[3][0][17] )
         );
  dff_sg \reg_in_reg[3][0][16]  ( .D(n4442), .CP(clk), .Q(\reg_in[3][0][16] )
         );
  dff_sg \reg_in_reg[3][0][15]  ( .D(n4441), .CP(clk), .Q(\reg_in[3][0][15] )
         );
  dff_sg \reg_in_reg[3][0][14]  ( .D(n4440), .CP(clk), .Q(\reg_in[3][0][14] )
         );
  dff_sg \reg_in_reg[3][0][13]  ( .D(n4439), .CP(clk), .Q(\reg_in[3][0][13] )
         );
  dff_sg \reg_in_reg[3][0][12]  ( .D(n4438), .CP(clk), .Q(\reg_in[3][0][12] )
         );
  dff_sg \reg_in_reg[3][0][11]  ( .D(n4437), .CP(clk), .Q(\reg_in[3][0][11] )
         );
  dff_sg \reg_in_reg[3][0][10]  ( .D(n4436), .CP(clk), .Q(\reg_in[3][0][10] )
         );
  dff_sg \reg_in_reg[3][0][9]  ( .D(n4435), .CP(clk), .Q(\reg_in[3][0][9] ) );
  dff_sg \reg_in_reg[3][0][8]  ( .D(n4434), .CP(clk), .Q(\reg_in[3][0][8] ) );
  dff_sg \reg_in_reg[3][0][7]  ( .D(n4433), .CP(clk), .Q(\reg_in[3][0][7] ) );
  dff_sg \reg_in_reg[3][0][6]  ( .D(n4432), .CP(clk), .Q(\reg_in[3][0][6] ) );
  dff_sg \reg_in_reg[3][0][5]  ( .D(n4431), .CP(clk), .Q(\reg_in[3][0][5] ) );
  dff_sg \reg_in_reg[3][0][4]  ( .D(n4430), .CP(clk), .Q(\reg_in[3][0][4] ) );
  dff_sg \reg_in_reg[3][0][3]  ( .D(n4429), .CP(clk), .Q(\reg_in[3][0][3] ) );
  dff_sg \reg_in_reg[3][0][2]  ( .D(n4428), .CP(clk), .Q(\reg_in[3][0][2] ) );
  dff_sg \reg_in_reg[3][0][1]  ( .D(n4427), .CP(clk), .Q(\reg_in[3][0][1] ) );
  dff_sg \reg_in_reg[3][0][0]  ( .D(n4426), .CP(clk), .Q(\reg_in[3][0][0] ) );
  dff_sg \reg_in_reg[2][3][19]  ( .D(n4425), .CP(clk), .Q(\reg_in[2][3][19] )
         );
  dff_sg \reg_in_reg[2][3][18]  ( .D(n4424), .CP(clk), .Q(\reg_in[2][3][18] )
         );
  dff_sg \reg_in_reg[2][3][17]  ( .D(n4423), .CP(clk), .Q(\reg_in[2][3][17] )
         );
  dff_sg \reg_in_reg[2][3][16]  ( .D(n4422), .CP(clk), .Q(\reg_in[2][3][16] )
         );
  dff_sg \reg_in_reg[2][3][15]  ( .D(n4421), .CP(clk), .Q(\reg_in[2][3][15] )
         );
  dff_sg \reg_in_reg[2][3][14]  ( .D(n4420), .CP(clk), .Q(\reg_in[2][3][14] )
         );
  dff_sg \reg_in_reg[2][3][13]  ( .D(n4419), .CP(clk), .Q(\reg_in[2][3][13] )
         );
  dff_sg \reg_in_reg[2][3][12]  ( .D(n4418), .CP(clk), .Q(\reg_in[2][3][12] )
         );
  dff_sg \reg_in_reg[2][3][11]  ( .D(n4417), .CP(clk), .Q(\reg_in[2][3][11] )
         );
  dff_sg \reg_in_reg[2][3][10]  ( .D(n4416), .CP(clk), .Q(\reg_in[2][3][10] )
         );
  dff_sg \reg_in_reg[2][3][9]  ( .D(n4415), .CP(clk), .Q(\reg_in[2][3][9] ) );
  dff_sg \reg_in_reg[2][3][8]  ( .D(n4414), .CP(clk), .Q(\reg_in[2][3][8] ) );
  dff_sg \reg_in_reg[2][3][7]  ( .D(n4413), .CP(clk), .Q(\reg_in[2][3][7] ) );
  dff_sg \reg_in_reg[2][3][6]  ( .D(n4412), .CP(clk), .Q(\reg_in[2][3][6] ) );
  dff_sg \reg_in_reg[2][3][5]  ( .D(n4411), .CP(clk), .Q(\reg_in[2][3][5] ) );
  dff_sg \reg_in_reg[2][3][4]  ( .D(n4410), .CP(clk), .Q(\reg_in[2][3][4] ) );
  dff_sg \reg_in_reg[2][3][3]  ( .D(n4409), .CP(clk), .Q(\reg_in[2][3][3] ) );
  dff_sg \reg_in_reg[2][3][2]  ( .D(n4408), .CP(clk), .Q(\reg_in[2][3][2] ) );
  dff_sg \reg_in_reg[2][3][1]  ( .D(n4407), .CP(clk), .Q(\reg_in[2][3][1] ) );
  dff_sg \reg_in_reg[2][3][0]  ( .D(n4406), .CP(clk), .Q(\reg_in[2][3][0] ) );
  dff_sg \reg_in_reg[2][2][19]  ( .D(n4405), .CP(clk), .Q(\reg_in[2][2][19] )
         );
  dff_sg \reg_in_reg[2][2][18]  ( .D(n4404), .CP(clk), .Q(\reg_in[2][2][18] )
         );
  dff_sg \reg_in_reg[2][2][17]  ( .D(n4403), .CP(clk), .Q(\reg_in[2][2][17] )
         );
  dff_sg \reg_in_reg[2][2][16]  ( .D(n4402), .CP(clk), .Q(\reg_in[2][2][16] )
         );
  dff_sg \reg_in_reg[2][2][15]  ( .D(n4401), .CP(clk), .Q(\reg_in[2][2][15] )
         );
  dff_sg \reg_in_reg[2][2][14]  ( .D(n4400), .CP(clk), .Q(\reg_in[2][2][14] )
         );
  dff_sg \reg_in_reg[2][2][13]  ( .D(n4399), .CP(clk), .Q(\reg_in[2][2][13] )
         );
  dff_sg \reg_in_reg[2][2][12]  ( .D(n4398), .CP(clk), .Q(\reg_in[2][2][12] )
         );
  dff_sg \reg_in_reg[2][2][11]  ( .D(n4397), .CP(clk), .Q(\reg_in[2][2][11] )
         );
  dff_sg \reg_in_reg[2][2][10]  ( .D(n4396), .CP(clk), .Q(\reg_in[2][2][10] )
         );
  dff_sg \reg_in_reg[2][2][9]  ( .D(n4395), .CP(clk), .Q(\reg_in[2][2][9] ) );
  dff_sg \reg_in_reg[2][2][8]  ( .D(n4394), .CP(clk), .Q(\reg_in[2][2][8] ) );
  dff_sg \reg_in_reg[2][2][7]  ( .D(n4393), .CP(clk), .Q(\reg_in[2][2][7] ) );
  dff_sg \reg_in_reg[2][2][6]  ( .D(n4392), .CP(clk), .Q(\reg_in[2][2][6] ) );
  dff_sg \reg_in_reg[2][2][5]  ( .D(n4391), .CP(clk), .Q(\reg_in[2][2][5] ) );
  dff_sg \reg_in_reg[2][2][4]  ( .D(n4390), .CP(clk), .Q(\reg_in[2][2][4] ) );
  dff_sg \reg_in_reg[2][2][3]  ( .D(n4389), .CP(clk), .Q(\reg_in[2][2][3] ) );
  dff_sg \reg_in_reg[2][2][2]  ( .D(n4388), .CP(clk), .Q(\reg_in[2][2][2] ) );
  dff_sg \reg_in_reg[2][2][1]  ( .D(n4387), .CP(clk), .Q(\reg_in[2][2][1] ) );
  dff_sg \reg_in_reg[2][2][0]  ( .D(n4386), .CP(clk), .Q(\reg_in[2][2][0] ) );
  dff_sg \reg_in_reg[2][1][19]  ( .D(n4385), .CP(clk), .Q(\reg_in[2][1][19] )
         );
  dff_sg \reg_in_reg[2][1][18]  ( .D(n4384), .CP(clk), .Q(\reg_in[2][1][18] )
         );
  dff_sg \reg_in_reg[2][1][17]  ( .D(n4383), .CP(clk), .Q(\reg_in[2][1][17] )
         );
  dff_sg \reg_in_reg[2][1][16]  ( .D(n4382), .CP(clk), .Q(\reg_in[2][1][16] )
         );
  dff_sg \reg_in_reg[2][1][15]  ( .D(n4381), .CP(clk), .Q(\reg_in[2][1][15] )
         );
  dff_sg \reg_in_reg[2][1][14]  ( .D(n4380), .CP(clk), .Q(\reg_in[2][1][14] )
         );
  dff_sg \reg_in_reg[2][1][13]  ( .D(n4379), .CP(clk), .Q(\reg_in[2][1][13] )
         );
  dff_sg \reg_in_reg[2][1][12]  ( .D(n4378), .CP(clk), .Q(\reg_in[2][1][12] )
         );
  dff_sg \reg_in_reg[2][1][11]  ( .D(n4377), .CP(clk), .Q(\reg_in[2][1][11] )
         );
  dff_sg \reg_in_reg[2][1][10]  ( .D(n4376), .CP(clk), .Q(\reg_in[2][1][10] )
         );
  dff_sg \reg_in_reg[2][1][9]  ( .D(n4375), .CP(clk), .Q(\reg_in[2][1][9] ) );
  dff_sg \reg_in_reg[2][1][8]  ( .D(n4374), .CP(clk), .Q(\reg_in[2][1][8] ) );
  dff_sg \reg_in_reg[2][1][7]  ( .D(n4373), .CP(clk), .Q(\reg_in[2][1][7] ) );
  dff_sg \reg_in_reg[2][1][6]  ( .D(n4372), .CP(clk), .Q(\reg_in[2][1][6] ) );
  dff_sg \reg_in_reg[2][1][5]  ( .D(n4371), .CP(clk), .Q(\reg_in[2][1][5] ) );
  dff_sg \reg_in_reg[2][1][4]  ( .D(n4370), .CP(clk), .Q(\reg_in[2][1][4] ) );
  dff_sg \reg_in_reg[2][1][3]  ( .D(n4369), .CP(clk), .Q(\reg_in[2][1][3] ) );
  dff_sg \reg_in_reg[2][1][2]  ( .D(n4368), .CP(clk), .Q(\reg_in[2][1][2] ) );
  dff_sg \reg_in_reg[2][1][1]  ( .D(n4367), .CP(clk), .Q(\reg_in[2][1][1] ) );
  dff_sg \reg_in_reg[2][1][0]  ( .D(n4366), .CP(clk), .Q(\reg_in[2][1][0] ) );
  dff_sg \reg_in_reg[2][0][19]  ( .D(n4365), .CP(clk), .Q(\reg_in[2][0][19] )
         );
  dff_sg \reg_in_reg[2][0][18]  ( .D(n4364), .CP(clk), .Q(\reg_in[2][0][18] )
         );
  dff_sg \reg_in_reg[2][0][17]  ( .D(n4363), .CP(clk), .Q(\reg_in[2][0][17] )
         );
  dff_sg \reg_in_reg[2][0][16]  ( .D(n4362), .CP(clk), .Q(\reg_in[2][0][16] )
         );
  dff_sg \reg_in_reg[2][0][15]  ( .D(n4361), .CP(clk), .Q(\reg_in[2][0][15] )
         );
  dff_sg \reg_in_reg[2][0][14]  ( .D(n4360), .CP(clk), .Q(\reg_in[2][0][14] )
         );
  dff_sg \reg_in_reg[2][0][13]  ( .D(n4359), .CP(clk), .Q(\reg_in[2][0][13] )
         );
  dff_sg \reg_in_reg[2][0][12]  ( .D(n4358), .CP(clk), .Q(\reg_in[2][0][12] )
         );
  dff_sg \reg_in_reg[2][0][11]  ( .D(n4357), .CP(clk), .Q(\reg_in[2][0][11] )
         );
  dff_sg \reg_in_reg[2][0][10]  ( .D(n4356), .CP(clk), .Q(\reg_in[2][0][10] )
         );
  dff_sg \reg_in_reg[2][0][9]  ( .D(n4355), .CP(clk), .Q(\reg_in[2][0][9] ) );
  dff_sg \reg_in_reg[2][0][8]  ( .D(n4354), .CP(clk), .Q(\reg_in[2][0][8] ) );
  dff_sg \reg_in_reg[2][0][7]  ( .D(n4353), .CP(clk), .Q(\reg_in[2][0][7] ) );
  dff_sg \reg_in_reg[2][0][6]  ( .D(n4352), .CP(clk), .Q(\reg_in[2][0][6] ) );
  dff_sg \reg_in_reg[2][0][5]  ( .D(n4351), .CP(clk), .Q(\reg_in[2][0][5] ) );
  dff_sg \reg_in_reg[2][0][4]  ( .D(n4350), .CP(clk), .Q(\reg_in[2][0][4] ) );
  dff_sg \reg_in_reg[2][0][3]  ( .D(n4349), .CP(clk), .Q(\reg_in[2][0][3] ) );
  dff_sg \reg_in_reg[2][0][2]  ( .D(n4348), .CP(clk), .Q(\reg_in[2][0][2] ) );
  dff_sg \reg_in_reg[2][0][1]  ( .D(n4347), .CP(clk), .Q(\reg_in[2][0][1] ) );
  dff_sg \reg_in_reg[2][0][0]  ( .D(n4346), .CP(clk), .Q(\reg_in[2][0][0] ) );
  dff_sg \reg_in_reg[1][3][19]  ( .D(n4345), .CP(clk), .Q(\reg_in[1][3][19] )
         );
  dff_sg \reg_in_reg[1][3][18]  ( .D(n4344), .CP(clk), .Q(\reg_in[1][3][18] )
         );
  dff_sg \reg_in_reg[1][3][17]  ( .D(n4343), .CP(clk), .Q(\reg_in[1][3][17] )
         );
  dff_sg \reg_in_reg[1][3][16]  ( .D(n4342), .CP(clk), .Q(\reg_in[1][3][16] )
         );
  dff_sg \reg_in_reg[1][3][15]  ( .D(n4341), .CP(clk), .Q(\reg_in[1][3][15] )
         );
  dff_sg \reg_in_reg[1][3][14]  ( .D(n4340), .CP(clk), .Q(\reg_in[1][3][14] )
         );
  dff_sg \reg_in_reg[1][3][13]  ( .D(n4339), .CP(clk), .Q(\reg_in[1][3][13] )
         );
  dff_sg \reg_in_reg[1][3][12]  ( .D(n4338), .CP(clk), .Q(\reg_in[1][3][12] )
         );
  dff_sg \reg_in_reg[1][3][11]  ( .D(n4337), .CP(clk), .Q(\reg_in[1][3][11] )
         );
  dff_sg \reg_in_reg[1][3][10]  ( .D(n4336), .CP(clk), .Q(\reg_in[1][3][10] )
         );
  dff_sg \reg_in_reg[1][3][9]  ( .D(n4335), .CP(clk), .Q(\reg_in[1][3][9] ) );
  dff_sg \reg_in_reg[1][3][8]  ( .D(n4334), .CP(clk), .Q(\reg_in[1][3][8] ) );
  dff_sg \reg_in_reg[1][3][7]  ( .D(n4333), .CP(clk), .Q(\reg_in[1][3][7] ) );
  dff_sg \reg_in_reg[1][3][6]  ( .D(n4332), .CP(clk), .Q(\reg_in[1][3][6] ) );
  dff_sg \reg_in_reg[1][3][5]  ( .D(n4331), .CP(clk), .Q(\reg_in[1][3][5] ) );
  dff_sg \reg_in_reg[1][3][4]  ( .D(n4330), .CP(clk), .Q(\reg_in[1][3][4] ) );
  dff_sg \reg_in_reg[1][3][3]  ( .D(n4329), .CP(clk), .Q(\reg_in[1][3][3] ) );
  dff_sg \reg_in_reg[1][3][2]  ( .D(n4328), .CP(clk), .Q(\reg_in[1][3][2] ) );
  dff_sg \reg_in_reg[1][3][1]  ( .D(n4327), .CP(clk), .Q(\reg_in[1][3][1] ) );
  dff_sg \reg_in_reg[1][3][0]  ( .D(n4326), .CP(clk), .Q(\reg_in[1][3][0] ) );
  dff_sg \reg_in_reg[1][2][19]  ( .D(n4325), .CP(clk), .Q(\reg_in[1][2][19] )
         );
  dff_sg \reg_in_reg[1][2][18]  ( .D(n4324), .CP(clk), .Q(\reg_in[1][2][18] )
         );
  dff_sg \reg_in_reg[1][2][17]  ( .D(n4323), .CP(clk), .Q(\reg_in[1][2][17] )
         );
  dff_sg \reg_in_reg[1][2][16]  ( .D(n4322), .CP(clk), .Q(\reg_in[1][2][16] )
         );
  dff_sg \reg_in_reg[1][2][15]  ( .D(n4321), .CP(clk), .Q(\reg_in[1][2][15] )
         );
  dff_sg \reg_in_reg[1][2][14]  ( .D(n4320), .CP(clk), .Q(\reg_in[1][2][14] )
         );
  dff_sg \reg_in_reg[1][2][13]  ( .D(n4319), .CP(clk), .Q(\reg_in[1][2][13] )
         );
  dff_sg \reg_in_reg[1][2][12]  ( .D(n4318), .CP(clk), .Q(\reg_in[1][2][12] )
         );
  dff_sg \reg_in_reg[1][2][11]  ( .D(n4317), .CP(clk), .Q(\reg_in[1][2][11] )
         );
  dff_sg \reg_in_reg[1][2][10]  ( .D(n4316), .CP(clk), .Q(\reg_in[1][2][10] )
         );
  dff_sg \reg_in_reg[1][2][9]  ( .D(n4315), .CP(clk), .Q(\reg_in[1][2][9] ) );
  dff_sg \reg_in_reg[1][2][8]  ( .D(n4314), .CP(clk), .Q(\reg_in[1][2][8] ) );
  dff_sg \reg_in_reg[1][2][7]  ( .D(n4313), .CP(clk), .Q(\reg_in[1][2][7] ) );
  dff_sg \reg_in_reg[1][2][6]  ( .D(n4312), .CP(clk), .Q(\reg_in[1][2][6] ) );
  dff_sg \reg_in_reg[1][2][5]  ( .D(n4311), .CP(clk), .Q(\reg_in[1][2][5] ) );
  dff_sg \reg_in_reg[1][2][4]  ( .D(n4310), .CP(clk), .Q(\reg_in[1][2][4] ) );
  dff_sg \reg_in_reg[1][2][3]  ( .D(n4309), .CP(clk), .Q(\reg_in[1][2][3] ) );
  dff_sg \reg_in_reg[1][2][2]  ( .D(n4308), .CP(clk), .Q(\reg_in[1][2][2] ) );
  dff_sg \reg_in_reg[1][2][1]  ( .D(n4307), .CP(clk), .Q(\reg_in[1][2][1] ) );
  dff_sg \reg_in_reg[1][2][0]  ( .D(n4306), .CP(clk), .Q(\reg_in[1][2][0] ) );
  dff_sg \reg_in_reg[1][1][19]  ( .D(n4305), .CP(clk), .Q(\reg_in[1][1][19] )
         );
  dff_sg \reg_in_reg[1][1][18]  ( .D(n4304), .CP(clk), .Q(\reg_in[1][1][18] )
         );
  dff_sg \reg_in_reg[1][1][17]  ( .D(n4303), .CP(clk), .Q(\reg_in[1][1][17] )
         );
  dff_sg \reg_in_reg[1][1][16]  ( .D(n4302), .CP(clk), .Q(\reg_in[1][1][16] )
         );
  dff_sg \reg_in_reg[1][1][15]  ( .D(n4301), .CP(clk), .Q(\reg_in[1][1][15] )
         );
  dff_sg \reg_in_reg[1][1][14]  ( .D(n4300), .CP(clk), .Q(\reg_in[1][1][14] )
         );
  dff_sg \reg_in_reg[1][1][13]  ( .D(n4299), .CP(clk), .Q(\reg_in[1][1][13] )
         );
  dff_sg \reg_in_reg[1][1][12]  ( .D(n4298), .CP(clk), .Q(\reg_in[1][1][12] )
         );
  dff_sg \reg_in_reg[1][1][11]  ( .D(n4297), .CP(clk), .Q(\reg_in[1][1][11] )
         );
  dff_sg \reg_in_reg[1][1][10]  ( .D(n4296), .CP(clk), .Q(\reg_in[1][1][10] )
         );
  dff_sg \reg_in_reg[1][1][9]  ( .D(n4295), .CP(clk), .Q(\reg_in[1][1][9] ) );
  dff_sg \reg_in_reg[1][1][8]  ( .D(n4294), .CP(clk), .Q(\reg_in[1][1][8] ) );
  dff_sg \reg_in_reg[1][1][7]  ( .D(n4293), .CP(clk), .Q(\reg_in[1][1][7] ) );
  dff_sg \reg_in_reg[1][1][6]  ( .D(n4292), .CP(clk), .Q(\reg_in[1][1][6] ) );
  dff_sg \reg_in_reg[1][1][5]  ( .D(n4291), .CP(clk), .Q(\reg_in[1][1][5] ) );
  dff_sg \reg_in_reg[1][1][4]  ( .D(n4290), .CP(clk), .Q(\reg_in[1][1][4] ) );
  dff_sg \reg_in_reg[1][1][3]  ( .D(n4289), .CP(clk), .Q(\reg_in[1][1][3] ) );
  dff_sg \reg_in_reg[1][1][2]  ( .D(n4288), .CP(clk), .Q(\reg_in[1][1][2] ) );
  dff_sg \reg_in_reg[1][1][1]  ( .D(n4287), .CP(clk), .Q(\reg_in[1][1][1] ) );
  dff_sg \reg_in_reg[1][1][0]  ( .D(n4286), .CP(clk), .Q(\reg_in[1][1][0] ) );
  dff_sg \reg_in_reg[1][0][19]  ( .D(n4285), .CP(clk), .Q(\reg_in[1][0][19] )
         );
  dff_sg \reg_in_reg[1][0][18]  ( .D(n4284), .CP(clk), .Q(\reg_in[1][0][18] )
         );
  dff_sg \reg_in_reg[1][0][17]  ( .D(n4283), .CP(clk), .Q(\reg_in[1][0][17] )
         );
  dff_sg \reg_in_reg[1][0][16]  ( .D(n4282), .CP(clk), .Q(\reg_in[1][0][16] )
         );
  dff_sg \reg_in_reg[1][0][15]  ( .D(n4281), .CP(clk), .Q(\reg_in[1][0][15] )
         );
  dff_sg \reg_in_reg[1][0][14]  ( .D(n4280), .CP(clk), .Q(\reg_in[1][0][14] )
         );
  dff_sg \reg_in_reg[1][0][13]  ( .D(n4279), .CP(clk), .Q(\reg_in[1][0][13] )
         );
  dff_sg \reg_in_reg[1][0][12]  ( .D(n4278), .CP(clk), .Q(\reg_in[1][0][12] )
         );
  dff_sg \reg_in_reg[1][0][11]  ( .D(n4277), .CP(clk), .Q(\reg_in[1][0][11] )
         );
  dff_sg \reg_in_reg[1][0][10]  ( .D(n4276), .CP(clk), .Q(\reg_in[1][0][10] )
         );
  dff_sg \reg_in_reg[1][0][9]  ( .D(n4275), .CP(clk), .Q(\reg_in[1][0][9] ) );
  dff_sg \reg_in_reg[1][0][8]  ( .D(n4274), .CP(clk), .Q(\reg_in[1][0][8] ) );
  dff_sg \reg_in_reg[1][0][7]  ( .D(n4273), .CP(clk), .Q(\reg_in[1][0][7] ) );
  dff_sg \reg_in_reg[1][0][6]  ( .D(n4272), .CP(clk), .Q(\reg_in[1][0][6] ) );
  dff_sg \reg_in_reg[1][0][5]  ( .D(n4271), .CP(clk), .Q(\reg_in[1][0][5] ) );
  dff_sg \reg_in_reg[1][0][4]  ( .D(n4270), .CP(clk), .Q(\reg_in[1][0][4] ) );
  dff_sg \reg_in_reg[1][0][3]  ( .D(n4269), .CP(clk), .Q(\reg_in[1][0][3] ) );
  dff_sg \reg_in_reg[1][0][2]  ( .D(n4268), .CP(clk), .Q(\reg_in[1][0][2] ) );
  dff_sg \reg_in_reg[1][0][1]  ( .D(n4267), .CP(clk), .Q(\reg_in[1][0][1] ) );
  dff_sg \reg_in_reg[1][0][0]  ( .D(n4266), .CP(clk), .Q(\reg_in[1][0][0] ) );
  dff_sg \reg_in_reg[0][3][19]  ( .D(n4265), .CP(clk), .Q(\reg_in[0][3][19] )
         );
  dff_sg \reg_in_reg[0][3][18]  ( .D(n4264), .CP(clk), .Q(\reg_in[0][3][18] )
         );
  dff_sg \reg_in_reg[0][3][17]  ( .D(n4263), .CP(clk), .Q(\reg_in[0][3][17] )
         );
  dff_sg \reg_in_reg[0][3][16]  ( .D(n4262), .CP(clk), .Q(\reg_in[0][3][16] )
         );
  dff_sg \reg_in_reg[0][3][15]  ( .D(n4261), .CP(clk), .Q(\reg_in[0][3][15] )
         );
  dff_sg \reg_in_reg[0][3][14]  ( .D(n4260), .CP(clk), .Q(\reg_in[0][3][14] )
         );
  dff_sg \reg_in_reg[0][3][13]  ( .D(n4259), .CP(clk), .Q(\reg_in[0][3][13] )
         );
  dff_sg \reg_in_reg[0][3][12]  ( .D(n4258), .CP(clk), .Q(\reg_in[0][3][12] )
         );
  dff_sg \reg_in_reg[0][3][11]  ( .D(n4257), .CP(clk), .Q(\reg_in[0][3][11] )
         );
  dff_sg \reg_in_reg[0][3][10]  ( .D(n4256), .CP(clk), .Q(\reg_in[0][3][10] )
         );
  dff_sg \reg_in_reg[0][3][9]  ( .D(n4255), .CP(clk), .Q(\reg_in[0][3][9] ) );
  dff_sg \reg_in_reg[0][3][8]  ( .D(n4254), .CP(clk), .Q(\reg_in[0][3][8] ) );
  dff_sg \reg_in_reg[0][3][7]  ( .D(n4253), .CP(clk), .Q(\reg_in[0][3][7] ) );
  dff_sg \reg_in_reg[0][3][6]  ( .D(n4252), .CP(clk), .Q(\reg_in[0][3][6] ) );
  dff_sg \reg_in_reg[0][3][5]  ( .D(n4251), .CP(clk), .Q(\reg_in[0][3][5] ) );
  dff_sg \reg_in_reg[0][3][4]  ( .D(n4250), .CP(clk), .Q(\reg_in[0][3][4] ) );
  dff_sg \reg_in_reg[0][3][3]  ( .D(n4249), .CP(clk), .Q(\reg_in[0][3][3] ) );
  dff_sg \reg_in_reg[0][3][2]  ( .D(n4248), .CP(clk), .Q(\reg_in[0][3][2] ) );
  dff_sg \reg_in_reg[0][3][1]  ( .D(n4247), .CP(clk), .Q(\reg_in[0][3][1] ) );
  dff_sg \reg_in_reg[0][3][0]  ( .D(n4246), .CP(clk), .Q(\reg_in[0][3][0] ) );
  dff_sg \reg_in_reg[0][2][19]  ( .D(n4245), .CP(clk), .Q(\reg_in[0][2][19] )
         );
  dff_sg \reg_in_reg[0][2][18]  ( .D(n4244), .CP(clk), .Q(\reg_in[0][2][18] )
         );
  dff_sg \reg_in_reg[0][2][17]  ( .D(n4243), .CP(clk), .Q(\reg_in[0][2][17] )
         );
  dff_sg \reg_in_reg[0][2][16]  ( .D(n4242), .CP(clk), .Q(\reg_in[0][2][16] )
         );
  dff_sg \reg_in_reg[0][2][15]  ( .D(n4241), .CP(clk), .Q(\reg_in[0][2][15] )
         );
  dff_sg \reg_in_reg[0][2][14]  ( .D(n4240), .CP(clk), .Q(\reg_in[0][2][14] )
         );
  dff_sg \reg_in_reg[0][2][13]  ( .D(n4239), .CP(clk), .Q(\reg_in[0][2][13] )
         );
  dff_sg \reg_in_reg[0][2][12]  ( .D(n4238), .CP(clk), .Q(\reg_in[0][2][12] )
         );
  dff_sg \reg_in_reg[0][2][11]  ( .D(n4237), .CP(clk), .Q(\reg_in[0][2][11] )
         );
  dff_sg \reg_in_reg[0][2][10]  ( .D(n4236), .CP(clk), .Q(\reg_in[0][2][10] )
         );
  dff_sg \reg_in_reg[0][2][9]  ( .D(n4235), .CP(clk), .Q(\reg_in[0][2][9] ) );
  dff_sg \reg_in_reg[0][2][8]  ( .D(n4234), .CP(clk), .Q(\reg_in[0][2][8] ) );
  dff_sg \reg_in_reg[0][2][7]  ( .D(n4233), .CP(clk), .Q(\reg_in[0][2][7] ) );
  dff_sg \reg_in_reg[0][2][6]  ( .D(n4232), .CP(clk), .Q(\reg_in[0][2][6] ) );
  dff_sg \reg_in_reg[0][2][5]  ( .D(n4231), .CP(clk), .Q(\reg_in[0][2][5] ) );
  dff_sg \reg_in_reg[0][2][4]  ( .D(n4230), .CP(clk), .Q(\reg_in[0][2][4] ) );
  dff_sg \reg_in_reg[0][2][3]  ( .D(n4229), .CP(clk), .Q(\reg_in[0][2][3] ) );
  dff_sg \reg_in_reg[0][2][2]  ( .D(n4228), .CP(clk), .Q(\reg_in[0][2][2] ) );
  dff_sg \reg_in_reg[0][2][1]  ( .D(n4227), .CP(clk), .Q(\reg_in[0][2][1] ) );
  dff_sg \reg_in_reg[0][2][0]  ( .D(n4226), .CP(clk), .Q(\reg_in[0][2][0] ) );
  dff_sg \reg_in_reg[0][1][19]  ( .D(n4225), .CP(clk), .Q(\reg_in[0][1][19] )
         );
  dff_sg \reg_in_reg[0][1][18]  ( .D(n4224), .CP(clk), .Q(\reg_in[0][1][18] )
         );
  dff_sg \reg_in_reg[0][1][17]  ( .D(n4223), .CP(clk), .Q(\reg_in[0][1][17] )
         );
  dff_sg \reg_in_reg[0][1][16]  ( .D(n4222), .CP(clk), .Q(\reg_in[0][1][16] )
         );
  dff_sg \reg_in_reg[0][1][15]  ( .D(n4221), .CP(clk), .Q(\reg_in[0][1][15] )
         );
  dff_sg \reg_in_reg[0][1][14]  ( .D(n4220), .CP(clk), .Q(\reg_in[0][1][14] )
         );
  dff_sg \reg_in_reg[0][1][13]  ( .D(n4219), .CP(clk), .Q(\reg_in[0][1][13] )
         );
  dff_sg \reg_in_reg[0][1][12]  ( .D(n4218), .CP(clk), .Q(\reg_in[0][1][12] )
         );
  dff_sg \reg_in_reg[0][1][11]  ( .D(n4217), .CP(clk), .Q(\reg_in[0][1][11] )
         );
  dff_sg \reg_in_reg[0][1][10]  ( .D(n4216), .CP(clk), .Q(\reg_in[0][1][10] )
         );
  dff_sg \reg_in_reg[0][1][9]  ( .D(n4215), .CP(clk), .Q(\reg_in[0][1][9] ) );
  dff_sg \reg_in_reg[0][1][8]  ( .D(n4214), .CP(clk), .Q(\reg_in[0][1][8] ) );
  dff_sg \reg_in_reg[0][1][7]  ( .D(n4213), .CP(clk), .Q(\reg_in[0][1][7] ) );
  dff_sg \reg_in_reg[0][1][6]  ( .D(n4212), .CP(clk), .Q(\reg_in[0][1][6] ) );
  dff_sg \reg_in_reg[0][1][5]  ( .D(n4211), .CP(clk), .Q(\reg_in[0][1][5] ) );
  dff_sg \reg_in_reg[0][1][4]  ( .D(n4210), .CP(clk), .Q(\reg_in[0][1][4] ) );
  dff_sg \reg_in_reg[0][1][3]  ( .D(n4209), .CP(clk), .Q(\reg_in[0][1][3] ) );
  dff_sg \reg_in_reg[0][1][2]  ( .D(n4208), .CP(clk), .Q(\reg_in[0][1][2] ) );
  dff_sg \reg_in_reg[0][1][1]  ( .D(n4207), .CP(clk), .Q(\reg_in[0][1][1] ) );
  dff_sg \reg_in_reg[0][1][0]  ( .D(n4206), .CP(clk), .Q(\reg_in[0][1][0] ) );
  dff_sg \reg_in_reg[0][0][19]  ( .D(n4205), .CP(clk), .Q(\reg_in[0][0][19] )
         );
  dff_sg \reg_in_reg[0][0][18]  ( .D(n4204), .CP(clk), .Q(\reg_in[0][0][18] )
         );
  dff_sg \reg_in_reg[0][0][17]  ( .D(n4203), .CP(clk), .Q(\reg_in[0][0][17] )
         );
  dff_sg \reg_in_reg[0][0][16]  ( .D(n4202), .CP(clk), .Q(\reg_in[0][0][16] )
         );
  dff_sg \reg_in_reg[0][0][15]  ( .D(n4201), .CP(clk), .Q(\reg_in[0][0][15] )
         );
  dff_sg \reg_in_reg[0][0][14]  ( .D(n4200), .CP(clk), .Q(\reg_in[0][0][14] )
         );
  dff_sg \reg_in_reg[0][0][13]  ( .D(n4199), .CP(clk), .Q(\reg_in[0][0][13] )
         );
  dff_sg \reg_in_reg[0][0][12]  ( .D(n4198), .CP(clk), .Q(\reg_in[0][0][12] )
         );
  dff_sg \reg_in_reg[0][0][11]  ( .D(n4197), .CP(clk), .Q(\reg_in[0][0][11] )
         );
  dff_sg \reg_in_reg[0][0][10]  ( .D(n4196), .CP(clk), .Q(\reg_in[0][0][10] )
         );
  dff_sg \reg_in_reg[0][0][9]  ( .D(n4195), .CP(clk), .Q(\reg_in[0][0][9] ) );
  dff_sg \reg_in_reg[0][0][8]  ( .D(n4194), .CP(clk), .Q(\reg_in[0][0][8] ) );
  dff_sg \reg_in_reg[0][0][7]  ( .D(n4193), .CP(clk), .Q(\reg_in[0][0][7] ) );
  dff_sg \reg_in_reg[0][0][6]  ( .D(n4192), .CP(clk), .Q(\reg_in[0][0][6] ) );
  dff_sg \reg_in_reg[0][0][5]  ( .D(n4191), .CP(clk), .Q(\reg_in[0][0][5] ) );
  dff_sg \reg_in_reg[0][0][4]  ( .D(n4190), .CP(clk), .Q(\reg_in[0][0][4] ) );
  dff_sg \reg_in_reg[0][0][3]  ( .D(n4189), .CP(clk), .Q(\reg_in[0][0][3] ) );
  dff_sg \reg_in_reg[0][0][2]  ( .D(n4188), .CP(clk), .Q(\reg_in[0][0][2] ) );
  dff_sg \reg_in_reg[0][0][1]  ( .D(n4187), .CP(clk), .Q(\reg_in[0][0][1] ) );
  dff_sg \reg_in_reg[0][0][0]  ( .D(n4186), .CP(clk), .Q(\reg_in[0][0][0] ) );
  dff_sg \out_reg[3][3][19]  ( .D(n4185), .CP(clk), .Q(\out[3][3][19] ) );
  dff_sg \out_reg[3][3][18]  ( .D(n4184), .CP(clk), .Q(\out[3][3][18] ) );
  dff_sg \out_reg[3][3][17]  ( .D(n4183), .CP(clk), .Q(\out[3][3][17] ) );
  dff_sg \out_reg[3][3][16]  ( .D(n4182), .CP(clk), .Q(\out[3][3][16] ) );
  dff_sg \out_reg[3][3][15]  ( .D(n4181), .CP(clk), .Q(\out[3][3][15] ) );
  dff_sg \out_reg[3][3][14]  ( .D(n4180), .CP(clk), .Q(\out[3][3][14] ) );
  dff_sg \out_reg[3][3][13]  ( .D(n4179), .CP(clk), .Q(\out[3][3][13] ) );
  dff_sg \out_reg[3][3][12]  ( .D(n4178), .CP(clk), .Q(\out[3][3][12] ) );
  dff_sg \out_reg[3][3][11]  ( .D(n4177), .CP(clk), .Q(\out[3][3][11] ) );
  dff_sg \out_reg[3][3][10]  ( .D(n4176), .CP(clk), .Q(\out[3][3][10] ) );
  dff_sg \out_reg[3][3][9]  ( .D(n4175), .CP(clk), .Q(\out[3][3][9] ) );
  dff_sg \out_reg[3][3][8]  ( .D(n4174), .CP(clk), .Q(\out[3][3][8] ) );
  dff_sg \out_reg[3][3][7]  ( .D(n4173), .CP(clk), .Q(\out[3][3][7] ) );
  dff_sg \out_reg[3][3][6]  ( .D(n4172), .CP(clk), .Q(\out[3][3][6] ) );
  dff_sg \out_reg[3][3][5]  ( .D(n4171), .CP(clk), .Q(\out[3][3][5] ) );
  dff_sg \out_reg[3][3][4]  ( .D(n4170), .CP(clk), .Q(\out[3][3][4] ) );
  dff_sg \out_reg[3][3][3]  ( .D(n4169), .CP(clk), .Q(\out[3][3][3] ) );
  dff_sg \out_reg[3][3][2]  ( .D(n4168), .CP(clk), .Q(\out[3][3][2] ) );
  dff_sg \out_reg[3][3][1]  ( .D(n4167), .CP(clk), .Q(\out[3][3][1] ) );
  dff_sg \out_reg[3][3][0]  ( .D(n4166), .CP(clk), .Q(\out[3][3][0] ) );
  dff_sg \out_reg[3][2][19]  ( .D(n4165), .CP(clk), .Q(\out[3][2][19] ) );
  dff_sg \out_reg[3][2][18]  ( .D(n4164), .CP(clk), .Q(\out[3][2][18] ) );
  dff_sg \out_reg[3][2][17]  ( .D(n4163), .CP(clk), .Q(\out[3][2][17] ) );
  dff_sg \out_reg[3][2][16]  ( .D(n4162), .CP(clk), .Q(\out[3][2][16] ) );
  dff_sg \out_reg[3][2][15]  ( .D(n4161), .CP(clk), .Q(\out[3][2][15] ) );
  dff_sg \out_reg[3][2][14]  ( .D(n4160), .CP(clk), .Q(\out[3][2][14] ) );
  dff_sg \out_reg[3][2][13]  ( .D(n4159), .CP(clk), .Q(\out[3][2][13] ) );
  dff_sg \out_reg[3][2][12]  ( .D(n4158), .CP(clk), .Q(\out[3][2][12] ) );
  dff_sg \out_reg[3][2][11]  ( .D(n4157), .CP(clk), .Q(\out[3][2][11] ) );
  dff_sg \out_reg[3][2][10]  ( .D(n4156), .CP(clk), .Q(\out[3][2][10] ) );
  dff_sg \out_reg[3][2][9]  ( .D(n4155), .CP(clk), .Q(\out[3][2][9] ) );
  dff_sg \out_reg[3][2][8]  ( .D(n4154), .CP(clk), .Q(\out[3][2][8] ) );
  dff_sg \out_reg[3][2][7]  ( .D(n4153), .CP(clk), .Q(\out[3][2][7] ) );
  dff_sg \out_reg[3][2][6]  ( .D(n4152), .CP(clk), .Q(\out[3][2][6] ) );
  dff_sg \out_reg[3][2][5]  ( .D(n4151), .CP(clk), .Q(\out[3][2][5] ) );
  dff_sg \out_reg[3][2][4]  ( .D(n4150), .CP(clk), .Q(\out[3][2][4] ) );
  dff_sg \out_reg[3][2][3]  ( .D(n4149), .CP(clk), .Q(\out[3][2][3] ) );
  dff_sg \out_reg[3][2][2]  ( .D(n4148), .CP(clk), .Q(\out[3][2][2] ) );
  dff_sg \out_reg[3][2][1]  ( .D(n4147), .CP(clk), .Q(\out[3][2][1] ) );
  dff_sg \out_reg[3][2][0]  ( .D(n4146), .CP(clk), .Q(\out[3][2][0] ) );
  dff_sg \out_reg[3][1][19]  ( .D(n4145), .CP(clk), .Q(\out[3][1][19] ) );
  dff_sg \out_reg[3][1][18]  ( .D(n4144), .CP(clk), .Q(\out[3][1][18] ) );
  dff_sg \out_reg[3][1][17]  ( .D(n4143), .CP(clk), .Q(\out[3][1][17] ) );
  dff_sg \out_reg[3][1][16]  ( .D(n4142), .CP(clk), .Q(\out[3][1][16] ) );
  dff_sg \out_reg[3][1][15]  ( .D(n4141), .CP(clk), .Q(\out[3][1][15] ) );
  dff_sg \out_reg[3][1][14]  ( .D(n4140), .CP(clk), .Q(\out[3][1][14] ) );
  dff_sg \out_reg[3][1][13]  ( .D(n4139), .CP(clk), .Q(\out[3][1][13] ) );
  dff_sg \out_reg[3][1][12]  ( .D(n4138), .CP(clk), .Q(\out[3][1][12] ) );
  dff_sg \out_reg[3][1][11]  ( .D(n4137), .CP(clk), .Q(\out[3][1][11] ) );
  dff_sg \out_reg[3][1][10]  ( .D(n4136), .CP(clk), .Q(\out[3][1][10] ) );
  dff_sg \out_reg[3][1][9]  ( .D(n4135), .CP(clk), .Q(\out[3][1][9] ) );
  dff_sg \out_reg[3][1][8]  ( .D(n4134), .CP(clk), .Q(\out[3][1][8] ) );
  dff_sg \out_reg[3][1][7]  ( .D(n4133), .CP(clk), .Q(\out[3][1][7] ) );
  dff_sg \out_reg[3][1][6]  ( .D(n4132), .CP(clk), .Q(\out[3][1][6] ) );
  dff_sg \out_reg[3][1][5]  ( .D(n4131), .CP(clk), .Q(\out[3][1][5] ) );
  dff_sg \out_reg[3][1][4]  ( .D(n4130), .CP(clk), .Q(\out[3][1][4] ) );
  dff_sg \out_reg[3][1][3]  ( .D(n4129), .CP(clk), .Q(\out[3][1][3] ) );
  dff_sg \out_reg[3][1][2]  ( .D(n4128), .CP(clk), .Q(\out[3][1][2] ) );
  dff_sg \out_reg[3][1][1]  ( .D(n4127), .CP(clk), .Q(\out[3][1][1] ) );
  dff_sg \out_reg[3][1][0]  ( .D(n4126), .CP(clk), .Q(\out[3][1][0] ) );
  dff_sg \out_reg[3][0][19]  ( .D(n4125), .CP(clk), .Q(\out[3][0][19] ) );
  dff_sg \out_reg[3][0][18]  ( .D(n4124), .CP(clk), .Q(\out[3][0][18] ) );
  dff_sg \out_reg[3][0][17]  ( .D(n4123), .CP(clk), .Q(\out[3][0][17] ) );
  dff_sg \out_reg[3][0][16]  ( .D(n4122), .CP(clk), .Q(\out[3][0][16] ) );
  dff_sg \out_reg[3][0][15]  ( .D(n4121), .CP(clk), .Q(\out[3][0][15] ) );
  dff_sg \out_reg[3][0][14]  ( .D(n4120), .CP(clk), .Q(\out[3][0][14] ) );
  dff_sg \out_reg[3][0][13]  ( .D(n4119), .CP(clk), .Q(\out[3][0][13] ) );
  dff_sg \out_reg[3][0][12]  ( .D(n4118), .CP(clk), .Q(\out[3][0][12] ) );
  dff_sg \out_reg[3][0][11]  ( .D(n4117), .CP(clk), .Q(\out[3][0][11] ) );
  dff_sg \out_reg[3][0][10]  ( .D(n4116), .CP(clk), .Q(\out[3][0][10] ) );
  dff_sg \out_reg[3][0][9]  ( .D(n4115), .CP(clk), .Q(\out[3][0][9] ) );
  dff_sg \out_reg[3][0][8]  ( .D(n4114), .CP(clk), .Q(\out[3][0][8] ) );
  dff_sg \out_reg[3][0][7]  ( .D(n4113), .CP(clk), .Q(\out[3][0][7] ) );
  dff_sg \out_reg[3][0][6]  ( .D(n4112), .CP(clk), .Q(\out[3][0][6] ) );
  dff_sg \out_reg[3][0][5]  ( .D(n4111), .CP(clk), .Q(\out[3][0][5] ) );
  dff_sg \out_reg[3][0][4]  ( .D(n4110), .CP(clk), .Q(\out[3][0][4] ) );
  dff_sg \out_reg[3][0][3]  ( .D(n4109), .CP(clk), .Q(\out[3][0][3] ) );
  dff_sg \out_reg[3][0][2]  ( .D(n4108), .CP(clk), .Q(\out[3][0][2] ) );
  dff_sg \out_reg[3][0][1]  ( .D(n4107), .CP(clk), .Q(\out[3][0][1] ) );
  dff_sg \out_reg[3][0][0]  ( .D(n4106), .CP(clk), .Q(\out[3][0][0] ) );
  dff_sg \out_reg[2][3][19]  ( .D(n4105), .CP(clk), .Q(\out[2][3][19] ) );
  dff_sg \out_reg[2][3][18]  ( .D(n4104), .CP(clk), .Q(\out[2][3][18] ) );
  dff_sg \out_reg[2][3][17]  ( .D(n4103), .CP(clk), .Q(\out[2][3][17] ) );
  dff_sg \out_reg[2][3][16]  ( .D(n4102), .CP(clk), .Q(\out[2][3][16] ) );
  dff_sg \out_reg[2][3][15]  ( .D(n4101), .CP(clk), .Q(\out[2][3][15] ) );
  dff_sg \out_reg[2][3][14]  ( .D(n4100), .CP(clk), .Q(\out[2][3][14] ) );
  dff_sg \out_reg[2][3][13]  ( .D(n4099), .CP(clk), .Q(\out[2][3][13] ) );
  dff_sg \out_reg[2][3][12]  ( .D(n4098), .CP(clk), .Q(\out[2][3][12] ) );
  dff_sg \out_reg[2][3][11]  ( .D(n4097), .CP(clk), .Q(\out[2][3][11] ) );
  dff_sg \out_reg[2][3][10]  ( .D(n4096), .CP(clk), .Q(\out[2][3][10] ) );
  dff_sg \out_reg[2][3][9]  ( .D(n4095), .CP(clk), .Q(\out[2][3][9] ) );
  dff_sg \out_reg[2][3][8]  ( .D(n4094), .CP(clk), .Q(\out[2][3][8] ) );
  dff_sg \out_reg[2][3][7]  ( .D(n4093), .CP(clk), .Q(\out[2][3][7] ) );
  dff_sg \out_reg[2][3][6]  ( .D(n4092), .CP(clk), .Q(\out[2][3][6] ) );
  dff_sg \out_reg[2][3][5]  ( .D(n4091), .CP(clk), .Q(\out[2][3][5] ) );
  dff_sg \out_reg[2][3][4]  ( .D(n4090), .CP(clk), .Q(\out[2][3][4] ) );
  dff_sg \out_reg[2][3][3]  ( .D(n4089), .CP(clk), .Q(\out[2][3][3] ) );
  dff_sg \out_reg[2][3][2]  ( .D(n4088), .CP(clk), .Q(\out[2][3][2] ) );
  dff_sg \out_reg[2][3][1]  ( .D(n4087), .CP(clk), .Q(\out[2][3][1] ) );
  dff_sg \out_reg[2][3][0]  ( .D(n4086), .CP(clk), .Q(\out[2][3][0] ) );
  dff_sg \out_reg[2][2][19]  ( .D(n4085), .CP(clk), .Q(\out[2][2][19] ) );
  dff_sg \out_reg[2][2][18]  ( .D(n4084), .CP(clk), .Q(\out[2][2][18] ) );
  dff_sg \out_reg[2][2][17]  ( .D(n4083), .CP(clk), .Q(\out[2][2][17] ) );
  dff_sg \out_reg[2][2][16]  ( .D(n4082), .CP(clk), .Q(\out[2][2][16] ) );
  dff_sg \out_reg[2][2][15]  ( .D(n4081), .CP(clk), .Q(\out[2][2][15] ) );
  dff_sg \out_reg[2][2][14]  ( .D(n4080), .CP(clk), .Q(\out[2][2][14] ) );
  dff_sg \out_reg[2][2][13]  ( .D(n4079), .CP(clk), .Q(\out[2][2][13] ) );
  dff_sg \out_reg[2][2][12]  ( .D(n4078), .CP(clk), .Q(\out[2][2][12] ) );
  dff_sg \out_reg[2][2][11]  ( .D(n4077), .CP(clk), .Q(\out[2][2][11] ) );
  dff_sg \out_reg[2][2][10]  ( .D(n4076), .CP(clk), .Q(\out[2][2][10] ) );
  dff_sg \out_reg[2][2][9]  ( .D(n4075), .CP(clk), .Q(\out[2][2][9] ) );
  dff_sg \out_reg[2][2][8]  ( .D(n4074), .CP(clk), .Q(\out[2][2][8] ) );
  dff_sg \out_reg[2][2][7]  ( .D(n4073), .CP(clk), .Q(\out[2][2][7] ) );
  dff_sg \out_reg[2][2][6]  ( .D(n4072), .CP(clk), .Q(\out[2][2][6] ) );
  dff_sg \out_reg[2][2][5]  ( .D(n4071), .CP(clk), .Q(\out[2][2][5] ) );
  dff_sg \out_reg[2][2][4]  ( .D(n4070), .CP(clk), .Q(\out[2][2][4] ) );
  dff_sg \out_reg[2][2][3]  ( .D(n4069), .CP(clk), .Q(\out[2][2][3] ) );
  dff_sg \out_reg[2][2][2]  ( .D(n4068), .CP(clk), .Q(\out[2][2][2] ) );
  dff_sg \out_reg[2][2][1]  ( .D(n4067), .CP(clk), .Q(\out[2][2][1] ) );
  dff_sg \out_reg[2][2][0]  ( .D(n4066), .CP(clk), .Q(\out[2][2][0] ) );
  dff_sg \out_reg[2][1][19]  ( .D(n4065), .CP(clk), .Q(\out[2][1][19] ) );
  dff_sg \out_reg[2][1][18]  ( .D(n4064), .CP(clk), .Q(\out[2][1][18] ) );
  dff_sg \out_reg[2][1][17]  ( .D(n4063), .CP(clk), .Q(\out[2][1][17] ) );
  dff_sg \out_reg[2][1][16]  ( .D(n4062), .CP(clk), .Q(\out[2][1][16] ) );
  dff_sg \out_reg[2][1][15]  ( .D(n4061), .CP(clk), .Q(\out[2][1][15] ) );
  dff_sg \out_reg[2][1][14]  ( .D(n4060), .CP(clk), .Q(\out[2][1][14] ) );
  dff_sg \out_reg[2][1][13]  ( .D(n4059), .CP(clk), .Q(\out[2][1][13] ) );
  dff_sg \out_reg[2][1][12]  ( .D(n4058), .CP(clk), .Q(\out[2][1][12] ) );
  dff_sg \out_reg[2][1][11]  ( .D(n4057), .CP(clk), .Q(\out[2][1][11] ) );
  dff_sg \out_reg[2][1][10]  ( .D(n4056), .CP(clk), .Q(\out[2][1][10] ) );
  dff_sg \out_reg[2][1][9]  ( .D(n4055), .CP(clk), .Q(\out[2][1][9] ) );
  dff_sg \out_reg[2][1][8]  ( .D(n4054), .CP(clk), .Q(\out[2][1][8] ) );
  dff_sg \out_reg[2][1][7]  ( .D(n4053), .CP(clk), .Q(\out[2][1][7] ) );
  dff_sg \out_reg[2][1][6]  ( .D(n4052), .CP(clk), .Q(\out[2][1][6] ) );
  dff_sg \out_reg[2][1][5]  ( .D(n4051), .CP(clk), .Q(\out[2][1][5] ) );
  dff_sg \out_reg[2][1][4]  ( .D(n4050), .CP(clk), .Q(\out[2][1][4] ) );
  dff_sg \out_reg[2][1][3]  ( .D(n4049), .CP(clk), .Q(\out[2][1][3] ) );
  dff_sg \out_reg[2][1][2]  ( .D(n4048), .CP(clk), .Q(\out[2][1][2] ) );
  dff_sg \out_reg[2][1][1]  ( .D(n4047), .CP(clk), .Q(\out[2][1][1] ) );
  dff_sg \out_reg[2][1][0]  ( .D(n4046), .CP(clk), .Q(\out[2][1][0] ) );
  dff_sg \out_reg[2][0][19]  ( .D(n4045), .CP(clk), .Q(\out[2][0][19] ) );
  dff_sg \out_reg[2][0][18]  ( .D(n4044), .CP(clk), .Q(\out[2][0][18] ) );
  dff_sg \out_reg[2][0][17]  ( .D(n4043), .CP(clk), .Q(\out[2][0][17] ) );
  dff_sg \out_reg[2][0][16]  ( .D(n4042), .CP(clk), .Q(\out[2][0][16] ) );
  dff_sg \out_reg[2][0][15]  ( .D(n4041), .CP(clk), .Q(\out[2][0][15] ) );
  dff_sg \out_reg[2][0][14]  ( .D(n4040), .CP(clk), .Q(\out[2][0][14] ) );
  dff_sg \out_reg[2][0][13]  ( .D(n4039), .CP(clk), .Q(\out[2][0][13] ) );
  dff_sg \out_reg[2][0][12]  ( .D(n4038), .CP(clk), .Q(\out[2][0][12] ) );
  dff_sg \out_reg[2][0][11]  ( .D(n4037), .CP(clk), .Q(\out[2][0][11] ) );
  dff_sg \out_reg[2][0][10]  ( .D(n4036), .CP(clk), .Q(\out[2][0][10] ) );
  dff_sg \out_reg[2][0][9]  ( .D(n4035), .CP(clk), .Q(\out[2][0][9] ) );
  dff_sg \out_reg[2][0][8]  ( .D(n4034), .CP(clk), .Q(\out[2][0][8] ) );
  dff_sg \out_reg[2][0][7]  ( .D(n4033), .CP(clk), .Q(\out[2][0][7] ) );
  dff_sg \out_reg[2][0][6]  ( .D(n4032), .CP(clk), .Q(\out[2][0][6] ) );
  dff_sg \out_reg[2][0][5]  ( .D(n4031), .CP(clk), .Q(\out[2][0][5] ) );
  dff_sg \out_reg[2][0][4]  ( .D(n4030), .CP(clk), .Q(\out[2][0][4] ) );
  dff_sg \out_reg[2][0][3]  ( .D(n4029), .CP(clk), .Q(\out[2][0][3] ) );
  dff_sg \out_reg[2][0][2]  ( .D(n4028), .CP(clk), .Q(\out[2][0][2] ) );
  dff_sg \out_reg[2][0][1]  ( .D(n4027), .CP(clk), .Q(\out[2][0][1] ) );
  dff_sg \out_reg[2][0][0]  ( .D(n4026), .CP(clk), .Q(\out[2][0][0] ) );
  dff_sg \out_reg[1][3][19]  ( .D(n4025), .CP(clk), .Q(\out[1][3][19] ) );
  dff_sg \out_reg[1][3][18]  ( .D(n4024), .CP(clk), .Q(\out[1][3][18] ) );
  dff_sg \out_reg[1][3][17]  ( .D(n4023), .CP(clk), .Q(\out[1][3][17] ) );
  dff_sg \out_reg[1][3][16]  ( .D(n4022), .CP(clk), .Q(\out[1][3][16] ) );
  dff_sg \out_reg[1][3][15]  ( .D(n4021), .CP(clk), .Q(\out[1][3][15] ) );
  dff_sg \out_reg[1][3][14]  ( .D(n4020), .CP(clk), .Q(\out[1][3][14] ) );
  dff_sg \out_reg[1][3][13]  ( .D(n4019), .CP(clk), .Q(\out[1][3][13] ) );
  dff_sg \out_reg[1][3][12]  ( .D(n4018), .CP(clk), .Q(\out[1][3][12] ) );
  dff_sg \out_reg[1][3][11]  ( .D(n4017), .CP(clk), .Q(\out[1][3][11] ) );
  dff_sg \out_reg[1][3][10]  ( .D(n4016), .CP(clk), .Q(\out[1][3][10] ) );
  dff_sg \out_reg[1][3][9]  ( .D(n4015), .CP(clk), .Q(\out[1][3][9] ) );
  dff_sg \out_reg[1][3][8]  ( .D(n4014), .CP(clk), .Q(\out[1][3][8] ) );
  dff_sg \out_reg[1][3][7]  ( .D(n4013), .CP(clk), .Q(\out[1][3][7] ) );
  dff_sg \out_reg[1][3][6]  ( .D(n4012), .CP(clk), .Q(\out[1][3][6] ) );
  dff_sg \out_reg[1][3][5]  ( .D(n4011), .CP(clk), .Q(\out[1][3][5] ) );
  dff_sg \out_reg[1][3][4]  ( .D(n4010), .CP(clk), .Q(\out[1][3][4] ) );
  dff_sg \out_reg[1][3][3]  ( .D(n4009), .CP(clk), .Q(\out[1][3][3] ) );
  dff_sg \out_reg[1][3][2]  ( .D(n4008), .CP(clk), .Q(\out[1][3][2] ) );
  dff_sg \out_reg[1][3][1]  ( .D(n4007), .CP(clk), .Q(\out[1][3][1] ) );
  dff_sg \out_reg[1][3][0]  ( .D(n4006), .CP(clk), .Q(\out[1][3][0] ) );
  dff_sg \out_reg[1][2][19]  ( .D(n4005), .CP(clk), .Q(\out[1][2][19] ) );
  dff_sg \out_reg[1][2][18]  ( .D(n4004), .CP(clk), .Q(\out[1][2][18] ) );
  dff_sg \out_reg[1][2][17]  ( .D(n4003), .CP(clk), .Q(\out[1][2][17] ) );
  dff_sg \out_reg[1][2][16]  ( .D(n4002), .CP(clk), .Q(\out[1][2][16] ) );
  dff_sg \out_reg[1][2][15]  ( .D(n4001), .CP(clk), .Q(\out[1][2][15] ) );
  dff_sg \out_reg[1][2][14]  ( .D(n4000), .CP(clk), .Q(\out[1][2][14] ) );
  dff_sg \out_reg[1][2][13]  ( .D(n3999), .CP(clk), .Q(\out[1][2][13] ) );
  dff_sg \out_reg[1][2][12]  ( .D(n3998), .CP(clk), .Q(\out[1][2][12] ) );
  dff_sg \out_reg[1][2][11]  ( .D(n3997), .CP(clk), .Q(\out[1][2][11] ) );
  dff_sg \out_reg[1][2][10]  ( .D(n3996), .CP(clk), .Q(\out[1][2][10] ) );
  dff_sg \out_reg[1][2][9]  ( .D(n3995), .CP(clk), .Q(\out[1][2][9] ) );
  dff_sg \out_reg[1][2][8]  ( .D(n3994), .CP(clk), .Q(\out[1][2][8] ) );
  dff_sg \out_reg[1][2][7]  ( .D(n3993), .CP(clk), .Q(\out[1][2][7] ) );
  dff_sg \out_reg[1][2][6]  ( .D(n3992), .CP(clk), .Q(\out[1][2][6] ) );
  dff_sg \out_reg[1][2][5]  ( .D(n3991), .CP(clk), .Q(\out[1][2][5] ) );
  dff_sg \out_reg[1][2][4]  ( .D(n3990), .CP(clk), .Q(\out[1][2][4] ) );
  dff_sg \out_reg[1][2][3]  ( .D(n3989), .CP(clk), .Q(\out[1][2][3] ) );
  dff_sg \out_reg[1][2][2]  ( .D(n3988), .CP(clk), .Q(\out[1][2][2] ) );
  dff_sg \out_reg[1][2][1]  ( .D(n3987), .CP(clk), .Q(\out[1][2][1] ) );
  dff_sg \out_reg[1][2][0]  ( .D(n3986), .CP(clk), .Q(\out[1][2][0] ) );
  dff_sg \out_reg[1][1][19]  ( .D(n3985), .CP(clk), .Q(\out[1][1][19] ) );
  dff_sg \out_reg[1][1][18]  ( .D(n3984), .CP(clk), .Q(\out[1][1][18] ) );
  dff_sg \out_reg[1][1][17]  ( .D(n3983), .CP(clk), .Q(\out[1][1][17] ) );
  dff_sg \out_reg[1][1][16]  ( .D(n3982), .CP(clk), .Q(\out[1][1][16] ) );
  dff_sg \out_reg[1][1][15]  ( .D(n3981), .CP(clk), .Q(\out[1][1][15] ) );
  dff_sg \out_reg[1][1][14]  ( .D(n3980), .CP(clk), .Q(\out[1][1][14] ) );
  dff_sg \out_reg[1][1][13]  ( .D(n3979), .CP(clk), .Q(\out[1][1][13] ) );
  dff_sg \out_reg[1][1][12]  ( .D(n3978), .CP(clk), .Q(\out[1][1][12] ) );
  dff_sg \out_reg[1][1][11]  ( .D(n3977), .CP(clk), .Q(\out[1][1][11] ) );
  dff_sg \out_reg[1][1][10]  ( .D(n3976), .CP(clk), .Q(\out[1][1][10] ) );
  dff_sg \out_reg[1][1][9]  ( .D(n3975), .CP(clk), .Q(\out[1][1][9] ) );
  dff_sg \out_reg[1][1][8]  ( .D(n3974), .CP(clk), .Q(\out[1][1][8] ) );
  dff_sg \out_reg[1][1][7]  ( .D(n3973), .CP(clk), .Q(\out[1][1][7] ) );
  dff_sg \out_reg[1][1][6]  ( .D(n3972), .CP(clk), .Q(\out[1][1][6] ) );
  dff_sg \out_reg[1][1][5]  ( .D(n3971), .CP(clk), .Q(\out[1][1][5] ) );
  dff_sg \out_reg[1][1][4]  ( .D(n3970), .CP(clk), .Q(\out[1][1][4] ) );
  dff_sg \out_reg[1][1][3]  ( .D(n3969), .CP(clk), .Q(\out[1][1][3] ) );
  dff_sg \out_reg[1][1][2]  ( .D(n3968), .CP(clk), .Q(\out[1][1][2] ) );
  dff_sg \out_reg[1][1][1]  ( .D(n3967), .CP(clk), .Q(\out[1][1][1] ) );
  dff_sg \out_reg[1][1][0]  ( .D(n3966), .CP(clk), .Q(\out[1][1][0] ) );
  dff_sg \out_reg[1][0][19]  ( .D(n3965), .CP(clk), .Q(\out[1][0][19] ) );
  dff_sg \out_reg[1][0][18]  ( .D(n3964), .CP(clk), .Q(\out[1][0][18] ) );
  dff_sg \out_reg[1][0][17]  ( .D(n3963), .CP(clk), .Q(\out[1][0][17] ) );
  dff_sg \out_reg[1][0][16]  ( .D(n3962), .CP(clk), .Q(\out[1][0][16] ) );
  dff_sg \out_reg[1][0][15]  ( .D(n3961), .CP(clk), .Q(\out[1][0][15] ) );
  dff_sg \out_reg[1][0][14]  ( .D(n3960), .CP(clk), .Q(\out[1][0][14] ) );
  dff_sg \out_reg[1][0][13]  ( .D(n3959), .CP(clk), .Q(\out[1][0][13] ) );
  dff_sg \out_reg[1][0][12]  ( .D(n3958), .CP(clk), .Q(\out[1][0][12] ) );
  dff_sg \out_reg[1][0][11]  ( .D(n3957), .CP(clk), .Q(\out[1][0][11] ) );
  dff_sg \out_reg[1][0][10]  ( .D(n3956), .CP(clk), .Q(\out[1][0][10] ) );
  dff_sg \out_reg[1][0][9]  ( .D(n3955), .CP(clk), .Q(\out[1][0][9] ) );
  dff_sg \out_reg[1][0][8]  ( .D(n3954), .CP(clk), .Q(\out[1][0][8] ) );
  dff_sg \out_reg[1][0][7]  ( .D(n3953), .CP(clk), .Q(\out[1][0][7] ) );
  dff_sg \out_reg[1][0][6]  ( .D(n3952), .CP(clk), .Q(\out[1][0][6] ) );
  dff_sg \out_reg[1][0][5]  ( .D(n3951), .CP(clk), .Q(\out[1][0][5] ) );
  dff_sg \out_reg[1][0][4]  ( .D(n3950), .CP(clk), .Q(\out[1][0][4] ) );
  dff_sg \out_reg[1][0][3]  ( .D(n3949), .CP(clk), .Q(\out[1][0][3] ) );
  dff_sg \out_reg[1][0][2]  ( .D(n3948), .CP(clk), .Q(\out[1][0][2] ) );
  dff_sg \out_reg[1][0][1]  ( .D(n3947), .CP(clk), .Q(\out[1][0][1] ) );
  dff_sg \out_reg[1][0][0]  ( .D(n3946), .CP(clk), .Q(\out[1][0][0] ) );
  dff_sg \out_reg[0][3][19]  ( .D(n3945), .CP(clk), .Q(\out[0][3][19] ) );
  dff_sg \out_reg[0][3][18]  ( .D(n3944), .CP(clk), .Q(\out[0][3][18] ) );
  dff_sg \out_reg[0][3][17]  ( .D(n3943), .CP(clk), .Q(\out[0][3][17] ) );
  dff_sg \out_reg[0][3][16]  ( .D(n3942), .CP(clk), .Q(\out[0][3][16] ) );
  dff_sg \out_reg[0][3][15]  ( .D(n3941), .CP(clk), .Q(\out[0][3][15] ) );
  dff_sg \out_reg[0][3][14]  ( .D(n3940), .CP(clk), .Q(\out[0][3][14] ) );
  dff_sg \out_reg[0][3][13]  ( .D(n3939), .CP(clk), .Q(\out[0][3][13] ) );
  dff_sg \out_reg[0][3][12]  ( .D(n3938), .CP(clk), .Q(\out[0][3][12] ) );
  dff_sg \out_reg[0][3][11]  ( .D(n3937), .CP(clk), .Q(\out[0][3][11] ) );
  dff_sg \out_reg[0][3][10]  ( .D(n3936), .CP(clk), .Q(\out[0][3][10] ) );
  dff_sg \out_reg[0][3][9]  ( .D(n3935), .CP(clk), .Q(\out[0][3][9] ) );
  dff_sg \out_reg[0][3][8]  ( .D(n3934), .CP(clk), .Q(\out[0][3][8] ) );
  dff_sg \out_reg[0][3][7]  ( .D(n3933), .CP(clk), .Q(\out[0][3][7] ) );
  dff_sg \out_reg[0][3][6]  ( .D(n3932), .CP(clk), .Q(\out[0][3][6] ) );
  dff_sg \out_reg[0][3][5]  ( .D(n3931), .CP(clk), .Q(\out[0][3][5] ) );
  dff_sg \out_reg[0][3][4]  ( .D(n3930), .CP(clk), .Q(\out[0][3][4] ) );
  dff_sg \out_reg[0][3][3]  ( .D(n3929), .CP(clk), .Q(\out[0][3][3] ) );
  dff_sg \out_reg[0][3][2]  ( .D(n3928), .CP(clk), .Q(\out[0][3][2] ) );
  dff_sg \out_reg[0][3][1]  ( .D(n3927), .CP(clk), .Q(\out[0][3][1] ) );
  dff_sg \out_reg[0][3][0]  ( .D(n3926), .CP(clk), .Q(\out[0][3][0] ) );
  dff_sg \out_reg[0][2][19]  ( .D(n3925), .CP(clk), .Q(\out[0][2][19] ) );
  dff_sg \out_reg[0][2][18]  ( .D(n3924), .CP(clk), .Q(\out[0][2][18] ) );
  dff_sg \out_reg[0][2][17]  ( .D(n3923), .CP(clk), .Q(\out[0][2][17] ) );
  dff_sg \out_reg[0][2][16]  ( .D(n3922), .CP(clk), .Q(\out[0][2][16] ) );
  dff_sg \out_reg[0][2][15]  ( .D(n3921), .CP(clk), .Q(\out[0][2][15] ) );
  dff_sg \out_reg[0][2][14]  ( .D(n3920), .CP(clk), .Q(\out[0][2][14] ) );
  dff_sg \out_reg[0][2][13]  ( .D(n3919), .CP(clk), .Q(\out[0][2][13] ) );
  dff_sg \out_reg[0][2][12]  ( .D(n3918), .CP(clk), .Q(\out[0][2][12] ) );
  dff_sg \out_reg[0][2][11]  ( .D(n3917), .CP(clk), .Q(\out[0][2][11] ) );
  dff_sg \out_reg[0][2][10]  ( .D(n3916), .CP(clk), .Q(\out[0][2][10] ) );
  dff_sg \out_reg[0][2][9]  ( .D(n3915), .CP(clk), .Q(\out[0][2][9] ) );
  dff_sg \out_reg[0][2][8]  ( .D(n3914), .CP(clk), .Q(\out[0][2][8] ) );
  dff_sg \out_reg[0][2][7]  ( .D(n3913), .CP(clk), .Q(\out[0][2][7] ) );
  dff_sg \out_reg[0][2][6]  ( .D(n3912), .CP(clk), .Q(\out[0][2][6] ) );
  dff_sg \out_reg[0][2][5]  ( .D(n3911), .CP(clk), .Q(\out[0][2][5] ) );
  dff_sg \out_reg[0][2][4]  ( .D(n3910), .CP(clk), .Q(\out[0][2][4] ) );
  dff_sg \out_reg[0][2][3]  ( .D(n3909), .CP(clk), .Q(\out[0][2][3] ) );
  dff_sg \out_reg[0][2][2]  ( .D(n3908), .CP(clk), .Q(\out[0][2][2] ) );
  dff_sg \out_reg[0][2][1]  ( .D(n3907), .CP(clk), .Q(\out[0][2][1] ) );
  dff_sg \out_reg[0][2][0]  ( .D(n3906), .CP(clk), .Q(\out[0][2][0] ) );
  dff_sg \out_reg[0][1][19]  ( .D(n3905), .CP(clk), .Q(\out[0][1][19] ) );
  dff_sg \out_reg[0][1][18]  ( .D(n3904), .CP(clk), .Q(\out[0][1][18] ) );
  dff_sg \out_reg[0][1][17]  ( .D(n3903), .CP(clk), .Q(\out[0][1][17] ) );
  dff_sg \out_reg[0][1][16]  ( .D(n3902), .CP(clk), .Q(\out[0][1][16] ) );
  dff_sg \out_reg[0][1][15]  ( .D(n3901), .CP(clk), .Q(\out[0][1][15] ) );
  dff_sg \out_reg[0][1][14]  ( .D(n3900), .CP(clk), .Q(\out[0][1][14] ) );
  dff_sg \out_reg[0][1][13]  ( .D(n3899), .CP(clk), .Q(\out[0][1][13] ) );
  dff_sg \out_reg[0][1][12]  ( .D(n3898), .CP(clk), .Q(\out[0][1][12] ) );
  dff_sg \out_reg[0][1][11]  ( .D(n3897), .CP(clk), .Q(\out[0][1][11] ) );
  dff_sg \out_reg[0][1][10]  ( .D(n3896), .CP(clk), .Q(\out[0][1][10] ) );
  dff_sg \out_reg[0][1][9]  ( .D(n3895), .CP(clk), .Q(\out[0][1][9] ) );
  dff_sg \out_reg[0][1][8]  ( .D(n3894), .CP(clk), .Q(\out[0][1][8] ) );
  dff_sg \out_reg[0][1][7]  ( .D(n3893), .CP(clk), .Q(\out[0][1][7] ) );
  dff_sg \out_reg[0][1][6]  ( .D(n3892), .CP(clk), .Q(\out[0][1][6] ) );
  dff_sg \out_reg[0][1][5]  ( .D(n3891), .CP(clk), .Q(\out[0][1][5] ) );
  dff_sg \out_reg[0][1][4]  ( .D(n3890), .CP(clk), .Q(\out[0][1][4] ) );
  dff_sg \out_reg[0][1][3]  ( .D(n3889), .CP(clk), .Q(\out[0][1][3] ) );
  dff_sg \out_reg[0][1][2]  ( .D(n3888), .CP(clk), .Q(\out[0][1][2] ) );
  dff_sg \out_reg[0][1][1]  ( .D(n3887), .CP(clk), .Q(\out[0][1][1] ) );
  dff_sg \out_reg[0][1][0]  ( .D(n3886), .CP(clk), .Q(\out[0][1][0] ) );
  dff_sg \out_reg[0][0][19]  ( .D(n3885), .CP(clk), .Q(\out[0][0][19] ) );
  dff_sg \out_reg[0][0][18]  ( .D(n3884), .CP(clk), .Q(\out[0][0][18] ) );
  dff_sg \out_reg[0][0][17]  ( .D(n3883), .CP(clk), .Q(\out[0][0][17] ) );
  dff_sg \out_reg[0][0][16]  ( .D(n3882), .CP(clk), .Q(\out[0][0][16] ) );
  dff_sg \out_reg[0][0][15]  ( .D(n3881), .CP(clk), .Q(\out[0][0][15] ) );
  dff_sg \out_reg[0][0][14]  ( .D(n3880), .CP(clk), .Q(\out[0][0][14] ) );
  dff_sg \out_reg[0][0][13]  ( .D(n3879), .CP(clk), .Q(\out[0][0][13] ) );
  dff_sg \out_reg[0][0][12]  ( .D(n3878), .CP(clk), .Q(\out[0][0][12] ) );
  dff_sg \out_reg[0][0][11]  ( .D(n3877), .CP(clk), .Q(\out[0][0][11] ) );
  dff_sg \out_reg[0][0][10]  ( .D(n3876), .CP(clk), .Q(\out[0][0][10] ) );
  dff_sg \out_reg[0][0][9]  ( .D(n3875), .CP(clk), .Q(\out[0][0][9] ) );
  dff_sg \out_reg[0][0][8]  ( .D(n3874), .CP(clk), .Q(\out[0][0][8] ) );
  dff_sg \out_reg[0][0][7]  ( .D(n3873), .CP(clk), .Q(\out[0][0][7] ) );
  dff_sg \out_reg[0][0][6]  ( .D(n3872), .CP(clk), .Q(\out[0][0][6] ) );
  dff_sg \out_reg[0][0][5]  ( .D(n3871), .CP(clk), .Q(\out[0][0][5] ) );
  dff_sg \out_reg[0][0][4]  ( .D(n3870), .CP(clk), .Q(\out[0][0][4] ) );
  dff_sg \out_reg[0][0][3]  ( .D(n3869), .CP(clk), .Q(\out[0][0][3] ) );
  dff_sg \out_reg[0][0][2]  ( .D(n3868), .CP(clk), .Q(\out[0][0][2] ) );
  dff_sg \out_reg[0][0][1]  ( .D(n3867), .CP(clk), .Q(\out[0][0][1] ) );
  dff_sg \out_reg[0][0][0]  ( .D(n3866), .CP(clk), .Q(\out[0][0][0] ) );
  \**FFGEN**  \reg_out_reg[3][3][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2271), .force_10(n11967), .force_11(1'b0), 
        .Q(n3865) );
  \**FFGEN**  \reg_out_reg[3][3][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2275), .force_10(n11968), .force_11(1'b0), 
        .Q(n3864) );
  \**FFGEN**  \reg_out_reg[3][3][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2279), .force_10(n11969), .force_11(1'b0), 
        .Q(n3863) );
  \**FFGEN**  \reg_out_reg[3][3][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2283), .force_10(n11970), .force_11(1'b0), 
        .Q(n3862) );
  \**FFGEN**  \reg_out_reg[3][3][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2287), .force_10(n11971), .force_11(1'b0), 
        .Q(n3861) );
  \**FFGEN**  \reg_out_reg[3][3][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2291), .force_10(n11972), .force_11(1'b0), 
        .Q(n3860) );
  \**FFGEN**  \reg_out_reg[3][3][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2295), .force_10(n11973), .force_11(1'b0), 
        .Q(n3859) );
  \**FFGEN**  \reg_out_reg[3][3][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2299), .force_10(n11974), .force_11(1'b0), 
        .Q(n3858) );
  \**FFGEN**  \reg_out_reg[3][3][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2303), .force_10(n11975), .force_11(1'b0), 
        .Q(n3857) );
  \**FFGEN**  \reg_out_reg[3][3][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2307), .force_10(n11976), .force_11(1'b0), 
        .Q(n3856) );
  \**FFGEN**  \reg_out_reg[3][3][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2311), .force_10(n11977), .force_11(1'b0), 
        .Q(n3855) );
  \**FFGEN**  \reg_out_reg[3][3][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2315), .force_10(n11978), .force_11(1'b0), 
        .Q(n3854) );
  \**FFGEN**  \reg_out_reg[3][3][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2319), .force_10(n11979), .force_11(1'b0), 
        .Q(n3853) );
  \**FFGEN**  \reg_out_reg[3][3][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2323), .force_10(n11980), .force_11(1'b0), 
        .Q(n3852) );
  \**FFGEN**  \reg_out_reg[3][3][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2327), .force_10(n11981), .force_11(1'b0), 
        .Q(n3851) );
  \**FFGEN**  \reg_out_reg[3][3][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2331), .force_10(n11982), .force_11(1'b0), 
        .Q(n3850) );
  \**FFGEN**  \reg_out_reg[3][3][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2335), .force_10(n11983), .force_11(1'b0), 
        .Q(n3849) );
  \**FFGEN**  \reg_out_reg[3][3][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2339), .force_10(n11984), .force_11(1'b0), 
        .Q(n3848) );
  \**FFGEN**  \reg_out_reg[3][3][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2343), .force_10(n11985), .force_11(1'b0), 
        .Q(n3847) );
  \**FFGEN**  \reg_out_reg[3][3][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2347), .force_10(n11986), .force_11(1'b0), 
        .Q(n3846) );
  \**FFGEN**  \reg_out_reg[3][2][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2351), .force_10(n11987), .force_11(1'b0), 
        .Q(n3845) );
  \**FFGEN**  \reg_out_reg[3][2][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2355), .force_10(n11988), .force_11(1'b0), 
        .Q(n3844) );
  \**FFGEN**  \reg_out_reg[3][2][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2359), .force_10(n11989), .force_11(1'b0), 
        .Q(n3843) );
  \**FFGEN**  \reg_out_reg[3][2][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2363), .force_10(n11990), .force_11(1'b0), 
        .Q(n3842) );
  \**FFGEN**  \reg_out_reg[3][2][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2367), .force_10(n11991), .force_11(1'b0), 
        .Q(n3841) );
  \**FFGEN**  \reg_out_reg[3][2][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2371), .force_10(n11992), .force_11(1'b0), 
        .Q(n3840) );
  \**FFGEN**  \reg_out_reg[3][2][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2375), .force_10(n11993), .force_11(1'b0), 
        .Q(n3839) );
  \**FFGEN**  \reg_out_reg[3][2][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2379), .force_10(n11994), .force_11(1'b0), 
        .Q(n3838) );
  \**FFGEN**  \reg_out_reg[3][2][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2383), .force_10(n11995), .force_11(1'b0), 
        .Q(n3837) );
  \**FFGEN**  \reg_out_reg[3][2][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2387), .force_10(n11996), .force_11(1'b0), 
        .Q(n3836) );
  \**FFGEN**  \reg_out_reg[3][2][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2391), .force_10(n11997), .force_11(1'b0), 
        .Q(n3835) );
  \**FFGEN**  \reg_out_reg[3][2][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2395), .force_10(n11998), .force_11(1'b0), 
        .Q(n3834) );
  \**FFGEN**  \reg_out_reg[3][2][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2399), .force_10(n11999), .force_11(1'b0), 
        .Q(n3833) );
  \**FFGEN**  \reg_out_reg[3][2][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2403), .force_10(n12000), .force_11(1'b0), 
        .Q(n3832) );
  \**FFGEN**  \reg_out_reg[3][2][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2407), .force_10(n12001), .force_11(1'b0), 
        .Q(n3831) );
  \**FFGEN**  \reg_out_reg[3][2][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2411), .force_10(n12002), .force_11(1'b0), 
        .Q(n3830) );
  \**FFGEN**  \reg_out_reg[3][2][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2415), .force_10(n12003), .force_11(1'b0), 
        .Q(n3829) );
  \**FFGEN**  \reg_out_reg[3][2][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2419), .force_10(n12004), .force_11(1'b0), 
        .Q(n3828) );
  \**FFGEN**  \reg_out_reg[3][2][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2423), .force_10(n12005), .force_11(1'b0), 
        .Q(n3827) );
  \**FFGEN**  \reg_out_reg[3][2][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2427), .force_10(n12006), .force_11(1'b0), 
        .Q(n3826) );
  \**FFGEN**  \reg_out_reg[3][1][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2431), .force_10(n12007), .force_11(1'b0), 
        .Q(n3825) );
  \**FFGEN**  \reg_out_reg[3][1][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2435), .force_10(n12008), .force_11(1'b0), 
        .Q(n3824) );
  \**FFGEN**  \reg_out_reg[3][1][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2439), .force_10(n12009), .force_11(1'b0), 
        .Q(n3823) );
  \**FFGEN**  \reg_out_reg[3][1][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2443), .force_10(n12010), .force_11(1'b0), 
        .Q(n3822) );
  \**FFGEN**  \reg_out_reg[3][1][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2447), .force_10(n12011), .force_11(1'b0), 
        .Q(n3821) );
  \**FFGEN**  \reg_out_reg[3][1][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2451), .force_10(n12012), .force_11(1'b0), 
        .Q(n3820) );
  \**FFGEN**  \reg_out_reg[3][1][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2455), .force_10(n12013), .force_11(1'b0), 
        .Q(n3819) );
  \**FFGEN**  \reg_out_reg[3][1][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2459), .force_10(n12014), .force_11(1'b0), 
        .Q(n3818) );
  \**FFGEN**  \reg_out_reg[3][1][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2463), .force_10(n12015), .force_11(1'b0), 
        .Q(n3817) );
  \**FFGEN**  \reg_out_reg[3][1][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2467), .force_10(n12016), .force_11(1'b0), 
        .Q(n3816) );
  \**FFGEN**  \reg_out_reg[3][1][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2471), .force_10(n12017), .force_11(1'b0), 
        .Q(n3815) );
  \**FFGEN**  \reg_out_reg[3][1][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2475), .force_10(n12018), .force_11(1'b0), 
        .Q(n3814) );
  \**FFGEN**  \reg_out_reg[3][1][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2479), .force_10(n12019), .force_11(1'b0), 
        .Q(n3813) );
  \**FFGEN**  \reg_out_reg[3][1][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2483), .force_10(n12020), .force_11(1'b0), 
        .Q(n3812) );
  \**FFGEN**  \reg_out_reg[3][1][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2487), .force_10(n12021), .force_11(1'b0), 
        .Q(n3811) );
  \**FFGEN**  \reg_out_reg[3][1][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2491), .force_10(n12022), .force_11(1'b0), 
        .Q(n3810) );
  \**FFGEN**  \reg_out_reg[3][1][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2495), .force_10(n12023), .force_11(1'b0), 
        .Q(n3809) );
  \**FFGEN**  \reg_out_reg[3][1][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2499), .force_10(n12024), .force_11(1'b0), 
        .Q(n3808) );
  \**FFGEN**  \reg_out_reg[3][1][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2503), .force_10(n12025), .force_11(1'b0), 
        .Q(n3807) );
  \**FFGEN**  \reg_out_reg[3][1][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2507), .force_10(n12026), .force_11(1'b0), 
        .Q(n3806) );
  \**FFGEN**  \reg_out_reg[3][0][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2511), .force_10(n12027), .force_11(1'b0), 
        .Q(n3805) );
  \**FFGEN**  \reg_out_reg[3][0][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2515), .force_10(n12028), .force_11(1'b0), 
        .Q(n3804) );
  \**FFGEN**  \reg_out_reg[3][0][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2519), .force_10(n12029), .force_11(1'b0), 
        .Q(n3803) );
  \**FFGEN**  \reg_out_reg[3][0][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2523), .force_10(n12030), .force_11(1'b0), 
        .Q(n3802) );
  \**FFGEN**  \reg_out_reg[3][0][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2527), .force_10(n12031), .force_11(1'b0), 
        .Q(n3801) );
  \**FFGEN**  \reg_out_reg[3][0][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2531), .force_10(n12032), .force_11(1'b0), 
        .Q(n3800) );
  \**FFGEN**  \reg_out_reg[3][0][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2535), .force_10(n12033), .force_11(1'b0), 
        .Q(n3799) );
  \**FFGEN**  \reg_out_reg[3][0][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2539), .force_10(n12034), .force_11(1'b0), 
        .Q(n3798) );
  \**FFGEN**  \reg_out_reg[3][0][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2543), .force_10(n12035), .force_11(1'b0), 
        .Q(n3797) );
  \**FFGEN**  \reg_out_reg[3][0][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2547), .force_10(n12036), .force_11(1'b0), 
        .Q(n3796) );
  \**FFGEN**  \reg_out_reg[3][0][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2551), .force_10(n12037), .force_11(1'b0), 
        .Q(n3795) );
  \**FFGEN**  \reg_out_reg[3][0][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2555), .force_10(n12038), .force_11(1'b0), 
        .Q(n3794) );
  \**FFGEN**  \reg_out_reg[3][0][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2559), .force_10(n12039), .force_11(1'b0), 
        .Q(n3793) );
  \**FFGEN**  \reg_out_reg[3][0][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2563), .force_10(n12040), .force_11(1'b0), 
        .Q(n3792) );
  \**FFGEN**  \reg_out_reg[3][0][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2567), .force_10(n12041), .force_11(1'b0), 
        .Q(n3791) );
  \**FFGEN**  \reg_out_reg[3][0][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2571), .force_10(n12042), .force_11(1'b0), 
        .Q(n3790) );
  \**FFGEN**  \reg_out_reg[3][0][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2575), .force_10(n12043), .force_11(1'b0), 
        .Q(n3789) );
  \**FFGEN**  \reg_out_reg[3][0][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2579), .force_10(n12044), .force_11(1'b0), 
        .Q(n3788) );
  \**FFGEN**  \reg_out_reg[3][0][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2583), .force_10(n12045), .force_11(1'b0), 
        .Q(n3787) );
  \**FFGEN**  \reg_out_reg[3][0][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2587), .force_10(n12046), .force_11(1'b0), 
        .Q(n3786) );
  \**FFGEN**  \reg_out_reg[2][3][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2591), .force_10(n12047), .force_11(1'b0), 
        .Q(n3785) );
  \**FFGEN**  \reg_out_reg[2][3][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2595), .force_10(n12048), .force_11(1'b0), 
        .Q(n3784) );
  \**FFGEN**  \reg_out_reg[2][3][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2599), .force_10(n12049), .force_11(1'b0), 
        .Q(n3783) );
  \**FFGEN**  \reg_out_reg[2][3][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2603), .force_10(n12050), .force_11(1'b0), 
        .Q(n3782) );
  \**FFGEN**  \reg_out_reg[2][3][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2607), .force_10(n12051), .force_11(1'b0), 
        .Q(n3781) );
  \**FFGEN**  \reg_out_reg[2][3][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2611), .force_10(n12052), .force_11(1'b0), 
        .Q(n3780) );
  \**FFGEN**  \reg_out_reg[2][3][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2615), .force_10(n12053), .force_11(1'b0), 
        .Q(n3779) );
  \**FFGEN**  \reg_out_reg[2][3][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2619), .force_10(n12054), .force_11(1'b0), 
        .Q(n3778) );
  \**FFGEN**  \reg_out_reg[2][3][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2623), .force_10(n12055), .force_11(1'b0), 
        .Q(n3777) );
  \**FFGEN**  \reg_out_reg[2][3][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2627), .force_10(n12056), .force_11(1'b0), 
        .Q(n3776) );
  \**FFGEN**  \reg_out_reg[2][3][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2631), .force_10(n12057), .force_11(1'b0), 
        .Q(n3775) );
  \**FFGEN**  \reg_out_reg[2][3][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2635), .force_10(n12058), .force_11(1'b0), 
        .Q(n3774) );
  \**FFGEN**  \reg_out_reg[2][3][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2639), .force_10(n12059), .force_11(1'b0), 
        .Q(n3773) );
  \**FFGEN**  \reg_out_reg[2][3][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2643), .force_10(n12060), .force_11(1'b0), 
        .Q(n3772) );
  \**FFGEN**  \reg_out_reg[2][3][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2647), .force_10(n12061), .force_11(1'b0), 
        .Q(n3771) );
  \**FFGEN**  \reg_out_reg[2][3][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2651), .force_10(n12062), .force_11(1'b0), 
        .Q(n3770) );
  \**FFGEN**  \reg_out_reg[2][3][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2655), .force_10(n12063), .force_11(1'b0), 
        .Q(n3769) );
  \**FFGEN**  \reg_out_reg[2][3][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2659), .force_10(n12064), .force_11(1'b0), 
        .Q(n3768) );
  \**FFGEN**  \reg_out_reg[2][3][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2663), .force_10(n12065), .force_11(1'b0), 
        .Q(n3767) );
  \**FFGEN**  \reg_out_reg[2][3][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2667), .force_10(n12066), .force_11(1'b0), 
        .Q(n3766) );
  \**FFGEN**  \reg_out_reg[2][2][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2671), .force_10(n12067), .force_11(1'b0), 
        .Q(n3765) );
  \**FFGEN**  \reg_out_reg[2][2][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2675), .force_10(n12068), .force_11(1'b0), 
        .Q(n3764) );
  \**FFGEN**  \reg_out_reg[2][2][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2679), .force_10(n12069), .force_11(1'b0), 
        .Q(n3763) );
  \**FFGEN**  \reg_out_reg[2][2][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2683), .force_10(n12070), .force_11(1'b0), 
        .Q(n3762) );
  \**FFGEN**  \reg_out_reg[2][2][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2687), .force_10(n12071), .force_11(1'b0), 
        .Q(n3761) );
  \**FFGEN**  \reg_out_reg[2][2][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2691), .force_10(n12072), .force_11(1'b0), 
        .Q(n3760) );
  \**FFGEN**  \reg_out_reg[2][2][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2695), .force_10(n12073), .force_11(1'b0), 
        .Q(n3759) );
  \**FFGEN**  \reg_out_reg[2][2][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2699), .force_10(n12074), .force_11(1'b0), 
        .Q(n3758) );
  \**FFGEN**  \reg_out_reg[2][2][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2703), .force_10(n12075), .force_11(1'b0), 
        .Q(n3757) );
  \**FFGEN**  \reg_out_reg[2][2][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2707), .force_10(n12076), .force_11(1'b0), 
        .Q(n3756) );
  \**FFGEN**  \reg_out_reg[2][2][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2711), .force_10(n12077), .force_11(1'b0), 
        .Q(n3755) );
  \**FFGEN**  \reg_out_reg[2][2][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2715), .force_10(n12078), .force_11(1'b0), 
        .Q(n3754) );
  \**FFGEN**  \reg_out_reg[2][2][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2719), .force_10(n12079), .force_11(1'b0), 
        .Q(n3753) );
  \**FFGEN**  \reg_out_reg[2][2][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2723), .force_10(n12080), .force_11(1'b0), 
        .Q(n3752) );
  \**FFGEN**  \reg_out_reg[2][2][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2727), .force_10(n12081), .force_11(1'b0), 
        .Q(n3751) );
  \**FFGEN**  \reg_out_reg[2][2][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2731), .force_10(n12082), .force_11(1'b0), 
        .Q(n3750) );
  \**FFGEN**  \reg_out_reg[2][2][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2735), .force_10(n12083), .force_11(1'b0), 
        .Q(n3749) );
  \**FFGEN**  \reg_out_reg[2][2][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2739), .force_10(n12084), .force_11(1'b0), 
        .Q(n3748) );
  \**FFGEN**  \reg_out_reg[2][2][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2743), .force_10(n12085), .force_11(1'b0), 
        .Q(n3747) );
  \**FFGEN**  \reg_out_reg[2][2][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2747), .force_10(n12086), .force_11(1'b0), 
        .Q(n3746) );
  \**FFGEN**  \reg_out_reg[2][1][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2751), .force_10(n12087), .force_11(1'b0), 
        .Q(n3745) );
  \**FFGEN**  \reg_out_reg[2][1][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2755), .force_10(n12088), .force_11(1'b0), 
        .Q(n3744) );
  \**FFGEN**  \reg_out_reg[2][1][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2759), .force_10(n12089), .force_11(1'b0), 
        .Q(n3743) );
  \**FFGEN**  \reg_out_reg[2][1][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2763), .force_10(n12090), .force_11(1'b0), 
        .Q(n3742) );
  \**FFGEN**  \reg_out_reg[2][1][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2767), .force_10(n12091), .force_11(1'b0), 
        .Q(n3741) );
  \**FFGEN**  \reg_out_reg[2][1][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2771), .force_10(n12092), .force_11(1'b0), 
        .Q(n3740) );
  \**FFGEN**  \reg_out_reg[2][1][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2775), .force_10(n12093), .force_11(1'b0), 
        .Q(n3739) );
  \**FFGEN**  \reg_out_reg[2][1][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2779), .force_10(n12094), .force_11(1'b0), 
        .Q(n3738) );
  \**FFGEN**  \reg_out_reg[2][1][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2783), .force_10(n12095), .force_11(1'b0), 
        .Q(n3737) );
  \**FFGEN**  \reg_out_reg[2][1][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2787), .force_10(n12096), .force_11(1'b0), 
        .Q(n3736) );
  \**FFGEN**  \reg_out_reg[2][1][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2791), .force_10(n12097), .force_11(1'b0), 
        .Q(n3735) );
  \**FFGEN**  \reg_out_reg[2][1][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2795), .force_10(n12098), .force_11(1'b0), 
        .Q(n3734) );
  \**FFGEN**  \reg_out_reg[2][1][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2799), .force_10(n12099), .force_11(1'b0), 
        .Q(n3733) );
  \**FFGEN**  \reg_out_reg[2][1][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2803), .force_10(n12100), .force_11(1'b0), 
        .Q(n3732) );
  \**FFGEN**  \reg_out_reg[2][1][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2807), .force_10(n12101), .force_11(1'b0), 
        .Q(n3731) );
  \**FFGEN**  \reg_out_reg[2][1][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2811), .force_10(n12102), .force_11(1'b0), 
        .Q(n3730) );
  \**FFGEN**  \reg_out_reg[2][1][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2815), .force_10(n12103), .force_11(1'b0), 
        .Q(n3729) );
  \**FFGEN**  \reg_out_reg[2][1][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2819), .force_10(n12104), .force_11(1'b0), 
        .Q(n3728) );
  \**FFGEN**  \reg_out_reg[2][1][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2823), .force_10(n12105), .force_11(1'b0), 
        .Q(n3727) );
  \**FFGEN**  \reg_out_reg[2][1][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2827), .force_10(n12106), .force_11(1'b0), 
        .Q(n3726) );
  \**FFGEN**  \reg_out_reg[2][0][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2831), .force_10(n12107), .force_11(1'b0), 
        .Q(n3725) );
  \**FFGEN**  \reg_out_reg[2][0][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2835), .force_10(n12108), .force_11(1'b0), 
        .Q(n3724) );
  \**FFGEN**  \reg_out_reg[2][0][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2839), .force_10(n12109), .force_11(1'b0), 
        .Q(n3723) );
  \**FFGEN**  \reg_out_reg[2][0][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2843), .force_10(n12110), .force_11(1'b0), 
        .Q(n3722) );
  \**FFGEN**  \reg_out_reg[2][0][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2847), .force_10(n12111), .force_11(1'b0), 
        .Q(n3721) );
  \**FFGEN**  \reg_out_reg[2][0][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2851), .force_10(n12112), .force_11(1'b0), 
        .Q(n3720) );
  \**FFGEN**  \reg_out_reg[2][0][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2855), .force_10(n12113), .force_11(1'b0), 
        .Q(n3719) );
  \**FFGEN**  \reg_out_reg[2][0][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2859), .force_10(n12114), .force_11(1'b0), 
        .Q(n3718) );
  \**FFGEN**  \reg_out_reg[2][0][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2863), .force_10(n12115), .force_11(1'b0), 
        .Q(n3717) );
  \**FFGEN**  \reg_out_reg[2][0][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2867), .force_10(n12116), .force_11(1'b0), 
        .Q(n3716) );
  \**FFGEN**  \reg_out_reg[2][0][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2871), .force_10(n12117), .force_11(1'b0), 
        .Q(n3715) );
  \**FFGEN**  \reg_out_reg[2][0][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2875), .force_10(n12118), .force_11(1'b0), 
        .Q(n3714) );
  \**FFGEN**  \reg_out_reg[2][0][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2879), .force_10(n12119), .force_11(1'b0), 
        .Q(n3713) );
  \**FFGEN**  \reg_out_reg[2][0][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2883), .force_10(n12120), .force_11(1'b0), 
        .Q(n3712) );
  \**FFGEN**  \reg_out_reg[2][0][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2887), .force_10(n12121), .force_11(1'b0), 
        .Q(n3711) );
  \**FFGEN**  \reg_out_reg[2][0][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2891), .force_10(n12122), .force_11(1'b0), 
        .Q(n3710) );
  \**FFGEN**  \reg_out_reg[2][0][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2895), .force_10(n12123), .force_11(1'b0), 
        .Q(n3709) );
  \**FFGEN**  \reg_out_reg[2][0][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2899), .force_10(n12124), .force_11(1'b0), 
        .Q(n3708) );
  \**FFGEN**  \reg_out_reg[2][0][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2903), .force_10(n12125), .force_11(1'b0), 
        .Q(n3707) );
  \**FFGEN**  \reg_out_reg[2][0][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2907), .force_10(n12126), .force_11(1'b0), 
        .Q(n3706) );
  \**FFGEN**  \reg_out_reg[1][3][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2911), .force_10(n12127), .force_11(1'b0), 
        .Q(n3705) );
  \**FFGEN**  \reg_out_reg[1][3][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2915), .force_10(n12128), .force_11(1'b0), 
        .Q(n3704) );
  \**FFGEN**  \reg_out_reg[1][3][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2919), .force_10(n12129), .force_11(1'b0), 
        .Q(n3703) );
  \**FFGEN**  \reg_out_reg[1][3][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2923), .force_10(n12130), .force_11(1'b0), 
        .Q(n3702) );
  \**FFGEN**  \reg_out_reg[1][3][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2927), .force_10(n12131), .force_11(1'b0), 
        .Q(n3701) );
  \**FFGEN**  \reg_out_reg[1][3][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2931), .force_10(n12132), .force_11(1'b0), 
        .Q(n3700) );
  \**FFGEN**  \reg_out_reg[1][3][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2935), .force_10(n12133), .force_11(1'b0), 
        .Q(n3699) );
  \**FFGEN**  \reg_out_reg[1][3][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2939), .force_10(n12134), .force_11(1'b0), 
        .Q(n3698) );
  \**FFGEN**  \reg_out_reg[1][3][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2943), .force_10(n12135), .force_11(1'b0), 
        .Q(n3697) );
  \**FFGEN**  \reg_out_reg[1][3][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2947), .force_10(n12136), .force_11(1'b0), 
        .Q(n3696) );
  \**FFGEN**  \reg_out_reg[1][3][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2951), .force_10(n12137), .force_11(1'b0), 
        .Q(n3695) );
  \**FFGEN**  \reg_out_reg[1][3][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2955), .force_10(n12138), .force_11(1'b0), 
        .Q(n3694) );
  \**FFGEN**  \reg_out_reg[1][3][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2959), .force_10(n12139), .force_11(1'b0), 
        .Q(n3693) );
  \**FFGEN**  \reg_out_reg[1][3][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2963), .force_10(n12140), .force_11(1'b0), 
        .Q(n3692) );
  \**FFGEN**  \reg_out_reg[1][3][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2967), .force_10(n12141), .force_11(1'b0), 
        .Q(n3691) );
  \**FFGEN**  \reg_out_reg[1][3][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2971), .force_10(n12142), .force_11(1'b0), 
        .Q(n3690) );
  \**FFGEN**  \reg_out_reg[1][3][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2975), .force_10(n12143), .force_11(1'b0), 
        .Q(n3689) );
  \**FFGEN**  \reg_out_reg[1][3][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2979), .force_10(n12144), .force_11(1'b0), 
        .Q(n3688) );
  \**FFGEN**  \reg_out_reg[1][3][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2983), .force_10(n12145), .force_11(1'b0), 
        .Q(n3687) );
  \**FFGEN**  \reg_out_reg[1][3][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2987), .force_10(n12146), .force_11(1'b0), 
        .Q(n3686) );
  \**FFGEN**  \reg_out_reg[1][2][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2991), .force_10(n12147), .force_11(1'b0), 
        .Q(n3685) );
  \**FFGEN**  \reg_out_reg[1][2][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2995), .force_10(n12148), .force_11(1'b0), 
        .Q(n3684) );
  \**FFGEN**  \reg_out_reg[1][2][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2999), .force_10(n12149), .force_11(1'b0), 
        .Q(n3683) );
  \**FFGEN**  \reg_out_reg[1][2][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3003), .force_10(n12150), .force_11(1'b0), 
        .Q(n3682) );
  \**FFGEN**  \reg_out_reg[1][2][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3007), .force_10(n12151), .force_11(1'b0), 
        .Q(n3681) );
  \**FFGEN**  \reg_out_reg[1][2][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3011), .force_10(n12152), .force_11(1'b0), 
        .Q(n3680) );
  \**FFGEN**  \reg_out_reg[1][2][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3015), .force_10(n12153), .force_11(1'b0), 
        .Q(n3679) );
  \**FFGEN**  \reg_out_reg[1][2][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3019), .force_10(n12154), .force_11(1'b0), 
        .Q(n3678) );
  \**FFGEN**  \reg_out_reg[1][2][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3023), .force_10(n12155), .force_11(1'b0), 
        .Q(n3677) );
  \**FFGEN**  \reg_out_reg[1][2][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3027), .force_10(n12156), .force_11(1'b0), 
        .Q(n3676) );
  \**FFGEN**  \reg_out_reg[1][2][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3031), .force_10(n12157), .force_11(1'b0), 
        .Q(n3675) );
  \**FFGEN**  \reg_out_reg[1][2][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3035), .force_10(n12158), .force_11(1'b0), 
        .Q(n3674) );
  \**FFGEN**  \reg_out_reg[1][2][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3039), .force_10(n12159), .force_11(1'b0), 
        .Q(n3673) );
  \**FFGEN**  \reg_out_reg[1][2][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3043), .force_10(n12160), .force_11(1'b0), 
        .Q(n3672) );
  \**FFGEN**  \reg_out_reg[1][2][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3047), .force_10(n12161), .force_11(1'b0), 
        .Q(n3671) );
  \**FFGEN**  \reg_out_reg[1][2][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3051), .force_10(n12162), .force_11(1'b0), 
        .Q(n3670) );
  \**FFGEN**  \reg_out_reg[1][2][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3055), .force_10(n12163), .force_11(1'b0), 
        .Q(n3669) );
  \**FFGEN**  \reg_out_reg[1][2][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3059), .force_10(n12164), .force_11(1'b0), 
        .Q(n3668) );
  \**FFGEN**  \reg_out_reg[1][2][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3063), .force_10(n12165), .force_11(1'b0), 
        .Q(n3667) );
  \**FFGEN**  \reg_out_reg[1][2][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3067), .force_10(n12166), .force_11(1'b0), 
        .Q(n3666) );
  \**FFGEN**  \reg_out_reg[1][1][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3071), .force_10(n12167), .force_11(1'b0), 
        .Q(n3665) );
  \**FFGEN**  \reg_out_reg[1][1][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3075), .force_10(n12168), .force_11(1'b0), 
        .Q(n3664) );
  \**FFGEN**  \reg_out_reg[1][1][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3079), .force_10(n12169), .force_11(1'b0), 
        .Q(n3663) );
  \**FFGEN**  \reg_out_reg[1][1][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3083), .force_10(n12170), .force_11(1'b0), 
        .Q(n3662) );
  \**FFGEN**  \reg_out_reg[1][1][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3087), .force_10(n12171), .force_11(1'b0), 
        .Q(n3661) );
  \**FFGEN**  \reg_out_reg[1][1][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3091), .force_10(n12172), .force_11(1'b0), 
        .Q(n3660) );
  \**FFGEN**  \reg_out_reg[1][1][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3095), .force_10(n12173), .force_11(1'b0), 
        .Q(n3659) );
  \**FFGEN**  \reg_out_reg[1][1][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3099), .force_10(n12174), .force_11(1'b0), 
        .Q(n3658) );
  \**FFGEN**  \reg_out_reg[1][1][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3103), .force_10(n12175), .force_11(1'b0), 
        .Q(n3657) );
  \**FFGEN**  \reg_out_reg[1][1][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3107), .force_10(n12176), .force_11(1'b0), 
        .Q(n3656) );
  \**FFGEN**  \reg_out_reg[1][1][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3111), .force_10(n12177), .force_11(1'b0), 
        .Q(n3655) );
  \**FFGEN**  \reg_out_reg[1][1][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3115), .force_10(n12178), .force_11(1'b0), 
        .Q(n3654) );
  \**FFGEN**  \reg_out_reg[1][1][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3119), .force_10(n12179), .force_11(1'b0), 
        .Q(n3653) );
  \**FFGEN**  \reg_out_reg[1][1][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3123), .force_10(n12180), .force_11(1'b0), 
        .Q(n3652) );
  \**FFGEN**  \reg_out_reg[1][1][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3127), .force_10(n12181), .force_11(1'b0), 
        .Q(n3651) );
  \**FFGEN**  \reg_out_reg[1][1][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3131), .force_10(n12182), .force_11(1'b0), 
        .Q(n3650) );
  \**FFGEN**  \reg_out_reg[1][1][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3135), .force_10(n12183), .force_11(1'b0), 
        .Q(n3649) );
  \**FFGEN**  \reg_out_reg[1][1][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3139), .force_10(n12184), .force_11(1'b0), 
        .Q(n3648) );
  \**FFGEN**  \reg_out_reg[1][1][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3143), .force_10(n12185), .force_11(1'b0), 
        .Q(n3647) );
  \**FFGEN**  \reg_out_reg[1][1][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3147), .force_10(n12186), .force_11(1'b0), 
        .Q(n3646) );
  \**FFGEN**  \reg_out_reg[1][0][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3151), .force_10(n12187), .force_11(1'b0), 
        .Q(n3645) );
  \**FFGEN**  \reg_out_reg[1][0][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3155), .force_10(n12188), .force_11(1'b0), 
        .Q(n3644) );
  \**FFGEN**  \reg_out_reg[1][0][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3159), .force_10(n12189), .force_11(1'b0), 
        .Q(n3643) );
  \**FFGEN**  \reg_out_reg[1][0][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3163), .force_10(n12190), .force_11(1'b0), 
        .Q(n3642) );
  \**FFGEN**  \reg_out_reg[1][0][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3167), .force_10(n12191), .force_11(1'b0), 
        .Q(n3641) );
  \**FFGEN**  \reg_out_reg[1][0][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3171), .force_10(n12192), .force_11(1'b0), 
        .Q(n3640) );
  \**FFGEN**  \reg_out_reg[1][0][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3175), .force_10(n12193), .force_11(1'b0), 
        .Q(n3639) );
  \**FFGEN**  \reg_out_reg[1][0][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3179), .force_10(n12194), .force_11(1'b0), 
        .Q(n3638) );
  \**FFGEN**  \reg_out_reg[1][0][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3183), .force_10(n12195), .force_11(1'b0), 
        .Q(n3637) );
  \**FFGEN**  \reg_out_reg[1][0][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3187), .force_10(n12196), .force_11(1'b0), 
        .Q(n3636) );
  \**FFGEN**  \reg_out_reg[1][0][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3191), .force_10(n12197), .force_11(1'b0), 
        .Q(n3635) );
  \**FFGEN**  \reg_out_reg[1][0][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3195), .force_10(n12198), .force_11(1'b0), 
        .Q(n3634) );
  \**FFGEN**  \reg_out_reg[1][0][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3199), .force_10(n12199), .force_11(1'b0), 
        .Q(n3633) );
  \**FFGEN**  \reg_out_reg[1][0][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3203), .force_10(n12200), .force_11(1'b0), 
        .Q(n3632) );
  \**FFGEN**  \reg_out_reg[1][0][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3207), .force_10(n12201), .force_11(1'b0), 
        .Q(n3631) );
  \**FFGEN**  \reg_out_reg[1][0][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3211), .force_10(n12202), .force_11(1'b0), 
        .Q(n3630) );
  \**FFGEN**  \reg_out_reg[1][0][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3215), .force_10(n12203), .force_11(1'b0), 
        .Q(n3629) );
  \**FFGEN**  \reg_out_reg[1][0][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3219), .force_10(n12204), .force_11(1'b0), 
        .Q(n3628) );
  \**FFGEN**  \reg_out_reg[1][0][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3223), .force_10(n12205), .force_11(1'b0), 
        .Q(n3627) );
  \**FFGEN**  \reg_out_reg[1][0][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3227), .force_10(n12206), .force_11(1'b0), 
        .Q(n3626) );
  \**FFGEN**  \reg_out_reg[0][3][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3231), .force_10(n12207), .force_11(1'b0), 
        .Q(n3625) );
  \**FFGEN**  \reg_out_reg[0][3][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3235), .force_10(n12208), .force_11(1'b0), 
        .Q(n3624) );
  \**FFGEN**  \reg_out_reg[0][3][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3239), .force_10(n12209), .force_11(1'b0), 
        .Q(n3623) );
  \**FFGEN**  \reg_out_reg[0][3][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3243), .force_10(n12210), .force_11(1'b0), 
        .Q(n3622) );
  \**FFGEN**  \reg_out_reg[0][3][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3247), .force_10(n12211), .force_11(1'b0), 
        .Q(n3621) );
  \**FFGEN**  \reg_out_reg[0][3][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3251), .force_10(n12212), .force_11(1'b0), 
        .Q(n3620) );
  \**FFGEN**  \reg_out_reg[0][3][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3255), .force_10(n12213), .force_11(1'b0), 
        .Q(n3619) );
  \**FFGEN**  \reg_out_reg[0][3][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3259), .force_10(n12214), .force_11(1'b0), 
        .Q(n3618) );
  \**FFGEN**  \reg_out_reg[0][3][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3263), .force_10(n12215), .force_11(1'b0), 
        .Q(n3617) );
  \**FFGEN**  \reg_out_reg[0][3][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3267), .force_10(n12216), .force_11(1'b0), 
        .Q(n3616) );
  \**FFGEN**  \reg_out_reg[0][3][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3271), .force_10(n12217), .force_11(1'b0), 
        .Q(n3615) );
  \**FFGEN**  \reg_out_reg[0][3][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3275), .force_10(n12218), .force_11(1'b0), 
        .Q(n3614) );
  \**FFGEN**  \reg_out_reg[0][3][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3279), .force_10(n12219), .force_11(1'b0), 
        .Q(n3613) );
  \**FFGEN**  \reg_out_reg[0][3][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3283), .force_10(n12220), .force_11(1'b0), 
        .Q(n3612) );
  \**FFGEN**  \reg_out_reg[0][3][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3287), .force_10(n12221), .force_11(1'b0), 
        .Q(n3611) );
  \**FFGEN**  \reg_out_reg[0][3][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3291), .force_10(n12222), .force_11(1'b0), 
        .Q(n3610) );
  \**FFGEN**  \reg_out_reg[0][3][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3295), .force_10(n12223), .force_11(1'b0), 
        .Q(n3609) );
  \**FFGEN**  \reg_out_reg[0][3][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3299), .force_10(n12224), .force_11(1'b0), 
        .Q(n3608) );
  \**FFGEN**  \reg_out_reg[0][3][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3303), .force_10(n12225), .force_11(1'b0), 
        .Q(n3607) );
  \**FFGEN**  \reg_out_reg[0][3][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3307), .force_10(n12226), .force_11(1'b0), 
        .Q(n3606) );
  \**FFGEN**  \reg_out_reg[0][2][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3311), .force_10(n12227), .force_11(1'b0), 
        .Q(n3605) );
  \**FFGEN**  \reg_out_reg[0][2][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3315), .force_10(n12228), .force_11(1'b0), 
        .Q(n3604) );
  \**FFGEN**  \reg_out_reg[0][2][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3319), .force_10(n12229), .force_11(1'b0), 
        .Q(n3603) );
  \**FFGEN**  \reg_out_reg[0][2][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3323), .force_10(n12230), .force_11(1'b0), 
        .Q(n3602) );
  \**FFGEN**  \reg_out_reg[0][2][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3327), .force_10(n12231), .force_11(1'b0), 
        .Q(n3601) );
  \**FFGEN**  \reg_out_reg[0][2][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3331), .force_10(n12232), .force_11(1'b0), 
        .Q(n3600) );
  \**FFGEN**  \reg_out_reg[0][2][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3335), .force_10(n12233), .force_11(1'b0), 
        .Q(n3599) );
  \**FFGEN**  \reg_out_reg[0][2][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3339), .force_10(n12234), .force_11(1'b0), 
        .Q(n3598) );
  \**FFGEN**  \reg_out_reg[0][2][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3343), .force_10(n12235), .force_11(1'b0), 
        .Q(n3597) );
  \**FFGEN**  \reg_out_reg[0][2][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3347), .force_10(n12236), .force_11(1'b0), 
        .Q(n3596) );
  \**FFGEN**  \reg_out_reg[0][2][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3351), .force_10(n12237), .force_11(1'b0), 
        .Q(n3595) );
  \**FFGEN**  \reg_out_reg[0][2][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3355), .force_10(n12238), .force_11(1'b0), 
        .Q(n3594) );
  \**FFGEN**  \reg_out_reg[0][2][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3359), .force_10(n12239), .force_11(1'b0), 
        .Q(n3593) );
  \**FFGEN**  \reg_out_reg[0][2][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3363), .force_10(n12240), .force_11(1'b0), 
        .Q(n3592) );
  \**FFGEN**  \reg_out_reg[0][2][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3367), .force_10(n12241), .force_11(1'b0), 
        .Q(n3591) );
  \**FFGEN**  \reg_out_reg[0][2][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3371), .force_10(n12242), .force_11(1'b0), 
        .Q(n3590) );
  \**FFGEN**  \reg_out_reg[0][2][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3375), .force_10(n12243), .force_11(1'b0), 
        .Q(n3589) );
  \**FFGEN**  \reg_out_reg[0][2][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3379), .force_10(n12244), .force_11(1'b0), 
        .Q(n3588) );
  \**FFGEN**  \reg_out_reg[0][2][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3383), .force_10(n12245), .force_11(1'b0), 
        .Q(n3587) );
  \**FFGEN**  \reg_out_reg[0][2][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3387), .force_10(n12246), .force_11(1'b0), 
        .Q(n3586) );
  \**FFGEN**  \reg_out_reg[0][1][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3391), .force_10(n12247), .force_11(1'b0), 
        .Q(n3585) );
  \**FFGEN**  \reg_out_reg[0][1][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3395), .force_10(n12248), .force_11(1'b0), 
        .Q(n3584) );
  \**FFGEN**  \reg_out_reg[0][1][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3399), .force_10(n12249), .force_11(1'b0), 
        .Q(n3583) );
  \**FFGEN**  \reg_out_reg[0][1][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3403), .force_10(n12250), .force_11(1'b0), 
        .Q(n3582) );
  \**FFGEN**  \reg_out_reg[0][1][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3407), .force_10(n12251), .force_11(1'b0), 
        .Q(n3581) );
  \**FFGEN**  \reg_out_reg[0][1][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3411), .force_10(n12252), .force_11(1'b0), 
        .Q(n3580) );
  \**FFGEN**  \reg_out_reg[0][1][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3415), .force_10(n12253), .force_11(1'b0), 
        .Q(n3579) );
  \**FFGEN**  \reg_out_reg[0][1][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3419), .force_10(n12254), .force_11(1'b0), 
        .Q(n3578) );
  \**FFGEN**  \reg_out_reg[0][1][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3423), .force_10(n12255), .force_11(1'b0), 
        .Q(n3577) );
  \**FFGEN**  \reg_out_reg[0][1][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3427), .force_10(n12256), .force_11(1'b0), 
        .Q(n3576) );
  \**FFGEN**  \reg_out_reg[0][1][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3431), .force_10(n12257), .force_11(1'b0), 
        .Q(n3575) );
  \**FFGEN**  \reg_out_reg[0][1][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3435), .force_10(n12258), .force_11(1'b0), 
        .Q(n3574) );
  \**FFGEN**  \reg_out_reg[0][1][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3439), .force_10(n12259), .force_11(1'b0), 
        .Q(n3573) );
  \**FFGEN**  \reg_out_reg[0][1][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3443), .force_10(n12260), .force_11(1'b0), 
        .Q(n3572) );
  \**FFGEN**  \reg_out_reg[0][1][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3447), .force_10(n12261), .force_11(1'b0), 
        .Q(n3571) );
  \**FFGEN**  \reg_out_reg[0][1][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3451), .force_10(n12262), .force_11(1'b0), 
        .Q(n3570) );
  \**FFGEN**  \reg_out_reg[0][1][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3455), .force_10(n12263), .force_11(1'b0), 
        .Q(n3569) );
  \**FFGEN**  \reg_out_reg[0][1][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3459), .force_10(n12264), .force_11(1'b0), 
        .Q(n3568) );
  \**FFGEN**  \reg_out_reg[0][1][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3463), .force_10(n12265), .force_11(1'b0), 
        .Q(n3567) );
  \**FFGEN**  \reg_out_reg[0][1][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3467), .force_10(n12266), .force_11(1'b0), 
        .Q(n3566) );
  \**FFGEN**  \reg_out_reg[0][0][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3471), .force_10(n12267), .force_11(1'b0), 
        .Q(n3565) );
  \**FFGEN**  \reg_out_reg[0][0][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3475), .force_10(n12268), .force_11(1'b0), 
        .Q(n3564) );
  \**FFGEN**  \reg_out_reg[0][0][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3479), .force_10(n12269), .force_11(1'b0), 
        .Q(n3563) );
  \**FFGEN**  \reg_out_reg[0][0][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3483), .force_10(n12270), .force_11(1'b0), 
        .Q(n3562) );
  \**FFGEN**  \reg_out_reg[0][0][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3487), .force_10(n12271), .force_11(1'b0), 
        .Q(n3561) );
  \**FFGEN**  \reg_out_reg[0][0][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3491), .force_10(n12272), .force_11(1'b0), 
        .Q(n3560) );
  \**FFGEN**  \reg_out_reg[0][0][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3495), .force_10(n12273), .force_11(1'b0), 
        .Q(n3559) );
  \**FFGEN**  \reg_out_reg[0][0][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3499), .force_10(n12274), .force_11(1'b0), 
        .Q(n3558) );
  \**FFGEN**  \reg_out_reg[0][0][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3503), .force_10(n12275), .force_11(1'b0), 
        .Q(n3557) );
  \**FFGEN**  \reg_out_reg[0][0][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3507), .force_10(n12276), .force_11(1'b0), 
        .Q(n3556) );
  \**FFGEN**  \reg_out_reg[0][0][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3511), .force_10(n12277), .force_11(1'b0), 
        .Q(n3555) );
  \**FFGEN**  \reg_out_reg[0][0][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3515), .force_10(n12278), .force_11(1'b0), 
        .Q(n3554) );
  \**FFGEN**  \reg_out_reg[0][0][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3519), .force_10(n12279), .force_11(1'b0), 
        .Q(n3553) );
  \**FFGEN**  \reg_out_reg[0][0][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3523), .force_10(n12280), .force_11(1'b0), 
        .Q(n3552) );
  \**FFGEN**  \reg_out_reg[0][0][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3527), .force_10(n12281), .force_11(1'b0), 
        .Q(n3551) );
  \**FFGEN**  \reg_out_reg[0][0][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3531), .force_10(n12282), .force_11(1'b0), 
        .Q(n3550) );
  \**FFGEN**  \reg_out_reg[0][0][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3535), .force_10(n12283), .force_11(1'b0), 
        .Q(n3549) );
  \**FFGEN**  \reg_out_reg[0][0][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3539), .force_10(n12284), .force_11(1'b0), 
        .Q(n3548) );
  \**FFGEN**  \reg_out_reg[0][0][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n3543), .force_10(n12285), .force_11(1'b0), 
        .Q(n3547) );
  \**FFGEN**  \reg_out_reg[0][0][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n2267), .force_10(n11966), .force_11(1'b0), 
        .Q(n3546) );
  nand_x1_sg U8370 ( .A(n8709), .B(n8710), .X(n8708) );
  inv_x1_sg U8371 ( .A(n8710), .X(n10682) );
  nor_x1_sg U8372 ( .A(reset), .B(n10001), .X(n8710) );
  nand_x1_sg U8373 ( .A(n10666), .B(n3573), .X(n9945) );
  nand_x1_sg U8374 ( .A(n10104), .B(n3666), .X(n9759) );
  nand_x1_sg U8375 ( .A(n10667), .B(n3790), .X(n9511) );
  nand_x1_sg U8376 ( .A(n10384), .B(n3856), .X(n9379) );
  nand_x16_sg U8377 ( .A(input_ready), .B(n12287), .X(n8715) );
  inv_x1_sg U8378 ( .A(n10375), .X(n10003) );
  inv_x1_sg U8379 ( .A(n10124), .X(n10004) );
  inv_x1_sg U8380 ( .A(n10004), .X(n10005) );
  inv_x1_sg U8381 ( .A(n10128), .X(n10006) );
  inv_x1_sg U8382 ( .A(n10133), .X(n10007) );
  inv_x1_sg U8383 ( .A(n10137), .X(n10008) );
  inv_x1_sg U8384 ( .A(n10142), .X(n10009) );
  inv_x1_sg U8385 ( .A(n10158), .X(n10010) );
  inv_x1_sg U8386 ( .A(n10220), .X(n10011) );
  inv_x1_sg U8387 ( .A(n10167), .X(n10012) );
  inv_x1_sg U8388 ( .A(n10175), .X(n10013) );
  inv_x1_sg U8389 ( .A(n10180), .X(n10014) );
  inv_x1_sg U8390 ( .A(n10185), .X(n10015) );
  inv_x1_sg U8391 ( .A(n10243), .X(n10016) );
  inv_x1_sg U8392 ( .A(n10290), .X(n10017) );
  inv_x1_sg U8393 ( .A(n10017), .X(n10018) );
  inv_x1_sg U8394 ( .A(n10309), .X(n10019) );
  inv_x1_sg U8395 ( .A(n10019), .X(n10020) );
  inv_x1_sg U8396 ( .A(n10257), .X(n10021) );
  inv_x1_sg U8397 ( .A(n10099), .X(n10022) );
  inv_x1_sg U8398 ( .A(n10078), .X(n10023) );
  inv_x1_sg U8399 ( .A(n10027), .X(n10024) );
  inv_x1_sg U8400 ( .A(n10027), .X(n10025) );
  inv_x1_sg U8401 ( .A(n10500), .X(n10026) );
  inv_x1_sg U8402 ( .A(n10429), .X(n10027) );
  inv_x1_sg U8403 ( .A(n10027), .X(n10028) );
  inv_x1_sg U8404 ( .A(n10030), .X(n10029) );
  inv_x1_sg U8405 ( .A(n10434), .X(n10030) );
  inv_x1_sg U8406 ( .A(n10030), .X(n10031) );
  inv_x1_sg U8407 ( .A(n10458), .X(n10032) );
  inv_x1_sg U8408 ( .A(n10117), .X(n10033) );
  inv_x1_sg U8409 ( .A(n10117), .X(n10034) );
  inv_x1_sg U8410 ( .A(n10456), .X(n10035) );
  inv_x1_sg U8411 ( .A(n10035), .X(n10036) );
  inv_x1_sg U8412 ( .A(n10124), .X(n10037) );
  inv_x1_sg U8413 ( .A(n10006), .X(n10038) );
  inv_x1_sg U8414 ( .A(n10130), .X(n10039) );
  inv_x1_sg U8415 ( .A(n10007), .X(n10040) );
  inv_x1_sg U8416 ( .A(n10008), .X(n10041) );
  inv_x1_sg U8417 ( .A(n10009), .X(n10042) );
  inv_x1_sg U8418 ( .A(n10139), .X(n10043) );
  inv_x1_sg U8419 ( .A(n10495), .X(n10044) );
  inv_x1_sg U8420 ( .A(n10149), .X(n10045) );
  inv_x1_sg U8421 ( .A(n10155), .X(n10046) );
  inv_x1_sg U8422 ( .A(n10160), .X(n10047) );
  inv_x1_sg U8423 ( .A(n10010), .X(n10048) );
  inv_x1_sg U8424 ( .A(n10163), .X(n10049) );
  inv_x1_sg U8425 ( .A(n10011), .X(n10050) );
  inv_x1_sg U8426 ( .A(n10012), .X(n10051) );
  inv_x1_sg U8427 ( .A(n10169), .X(n10052) );
  inv_x1_sg U8428 ( .A(n10517), .X(n10053) );
  inv_x1_sg U8429 ( .A(n10176), .X(n10054) );
  inv_x1_sg U8430 ( .A(n10013), .X(n10055) );
  inv_x1_sg U8431 ( .A(n10182), .X(n10056) );
  inv_x1_sg U8432 ( .A(n10014), .X(n10057) );
  inv_x1_sg U8433 ( .A(n10187), .X(n10058) );
  inv_x1_sg U8434 ( .A(n10015), .X(n10059) );
  inv_x1_sg U8435 ( .A(n10537), .X(n10060) );
  inv_x1_sg U8436 ( .A(n10019), .X(n10061) );
  inv_x1_sg U8437 ( .A(n10203), .X(n10062) );
  inv_x1_sg U8438 ( .A(n10244), .X(n10063) );
  inv_x1_sg U8439 ( .A(n10245), .X(n10064) );
  inv_x1_sg U8440 ( .A(n10557), .X(n10065) );
  inv_x1_sg U8441 ( .A(n10065), .X(n10066) );
  inv_x1_sg U8442 ( .A(n10557), .X(n10067) );
  inv_x1_sg U8443 ( .A(n10677), .X(n10068) );
  inv_x1_sg U8444 ( .A(n10248), .X(n10069) );
  inv_x1_sg U8445 ( .A(n10568), .X(n10070) );
  inv_x1_sg U8446 ( .A(n10582), .X(n10071) );
  inv_x1_sg U8447 ( .A(n10595), .X(n10072) );
  inv_x1_sg U8448 ( .A(n10076), .X(n10073) );
  inv_x1_sg U8449 ( .A(n10598), .X(n10074) );
  inv_x1_sg U8450 ( .A(n10599), .X(n10075) );
  inv_x1_sg U8451 ( .A(n10595), .X(n10076) );
  inv_x1_sg U8452 ( .A(n10597), .X(n10077) );
  inv_x1_sg U8453 ( .A(n10596), .X(n10078) );
  inv_x1_sg U8454 ( .A(n10082), .X(n10079) );
  inv_x1_sg U8455 ( .A(n10609), .X(n10080) );
  inv_x1_sg U8456 ( .A(n10610), .X(n10081) );
  inv_x1_sg U8457 ( .A(n10596), .X(n10082) );
  inv_x1_sg U8458 ( .A(n10611), .X(n10083) );
  inv_x1_sg U8459 ( .A(n10621), .X(n10084) );
  inv_x1_sg U8460 ( .A(n10075), .X(n10085) );
  inv_x1_sg U8461 ( .A(n10622), .X(n10086) );
  inv_x1_sg U8462 ( .A(n10635), .X(n10087) );
  inv_x1_sg U8463 ( .A(n10087), .X(n10088) );
  inv_x1_sg U8464 ( .A(n10639), .X(n10089) );
  inv_x1_sg U8465 ( .A(n10089), .X(n10090) );
  inv_x1_sg U8466 ( .A(n10090), .X(n10091) );
  inv_x1_sg U8467 ( .A(n10345), .X(n10092) );
  inv_x1_sg U8468 ( .A(n10096), .X(n10093) );
  inv_x1_sg U8469 ( .A(n10381), .X(n10094) );
  inv_x1_sg U8470 ( .A(n10101), .X(n10095) );
  inv_x1_sg U8471 ( .A(n8716), .X(n10096) );
  inv_x1_sg U8472 ( .A(n10640), .X(n10097) );
  inv_x1_sg U8473 ( .A(n10369), .X(n10098) );
  inv_x1_sg U8474 ( .A(n10003), .X(n10099) );
  inv_x1_sg U8475 ( .A(n10641), .X(n10100) );
  inv_x1_sg U8476 ( .A(n10108), .X(n10101) );
  inv_x1_sg U8477 ( .A(n10101), .X(n10102) );
  inv_x1_sg U8478 ( .A(n8716), .X(n10103) );
  inv_x1_sg U8479 ( .A(n10640), .X(n10104) );
  inv_x1_sg U8480 ( .A(n10665), .X(n10105) );
  inv_x1_sg U8481 ( .A(n10663), .X(n10106) );
  inv_x1_sg U8482 ( .A(n10260), .X(n10107) );
  inv_x1_sg U8483 ( .A(n10664), .X(n10108) );
  inv_x1_sg U8484 ( .A(n10414), .X(n10109) );
  inv_x1_sg U8485 ( .A(n10561), .X(n10110) );
  inv_x1_sg U8486 ( .A(n10418), .X(n10111) );
  inv_x1_sg U8487 ( .A(n10422), .X(n10112) );
  inv_x1_sg U8488 ( .A(n10423), .X(n10113) );
  inv_x1_sg U8489 ( .A(n10426), .X(n10114) );
  inv_x1_sg U8490 ( .A(n10438), .X(n10115) );
  inv_x1_sg U8491 ( .A(n10115), .X(n10116) );
  inv_x1_sg U8492 ( .A(n10202), .X(n10117) );
  inv_x1_sg U8493 ( .A(n10452), .X(n10118) );
  inv_x1_sg U8494 ( .A(n10118), .X(n10119) );
  inv_x1_sg U8495 ( .A(n10118), .X(n10120) );
  inv_x1_sg U8496 ( .A(n10120), .X(n10121) );
  inv_x1_sg U8497 ( .A(n10119), .X(n10122) );
  inv_x1_sg U8498 ( .A(n10044), .X(n10123) );
  inv_x1_sg U8499 ( .A(n10123), .X(n10124) );
  inv_x1_sg U8500 ( .A(n10123), .X(n10125) );
  inv_x1_sg U8501 ( .A(n10125), .X(n10126) );
  inv_x1_sg U8502 ( .A(n10124), .X(n10127) );
  inv_x1_sg U8503 ( .A(n10255), .X(n10128) );
  inv_x1_sg U8504 ( .A(n10128), .X(n10129) );
  inv_x1_sg U8505 ( .A(n10128), .X(n10130) );
  inv_x1_sg U8506 ( .A(n10129), .X(n10131) );
  inv_x1_sg U8507 ( .A(n10129), .X(n10132) );
  inv_x1_sg U8508 ( .A(n10218), .X(n10133) );
  inv_x1_sg U8509 ( .A(n10133), .X(n10134) );
  inv_x1_sg U8510 ( .A(n10134), .X(n10135) );
  inv_x1_sg U8511 ( .A(n10134), .X(n10136) );
  inv_x1_sg U8512 ( .A(n10210), .X(n10137) );
  inv_x1_sg U8513 ( .A(n10137), .X(n10138) );
  inv_x1_sg U8514 ( .A(n10137), .X(n10139) );
  inv_x1_sg U8515 ( .A(n10008), .X(n10140) );
  inv_x1_sg U8516 ( .A(n10138), .X(n10141) );
  inv_x1_sg U8517 ( .A(n10252), .X(n10142) );
  inv_x1_sg U8518 ( .A(n10142), .X(n10143) );
  inv_x1_sg U8519 ( .A(n10009), .X(n10144) );
  inv_x1_sg U8520 ( .A(n10143), .X(n10145) );
  inv_x1_sg U8521 ( .A(n10148), .X(n10146) );
  inv_x1_sg U8522 ( .A(n10542), .X(n10147) );
  inv_x1_sg U8523 ( .A(n10493), .X(n10148) );
  inv_x1_sg U8524 ( .A(n10148), .X(n10149) );
  inv_x1_sg U8525 ( .A(n10148), .X(n10150) );
  inv_x1_sg U8526 ( .A(n10150), .X(n10151) );
  inv_x1_sg U8527 ( .A(n10149), .X(n10152) );
  inv_x1_sg U8528 ( .A(n10498), .X(n10153) );
  inv_x1_sg U8529 ( .A(n10153), .X(n10154) );
  inv_x1_sg U8530 ( .A(n10153), .X(n10155) );
  inv_x1_sg U8531 ( .A(n10155), .X(n10156) );
  inv_x1_sg U8532 ( .A(n10154), .X(n10157) );
  inv_x1_sg U8533 ( .A(n10255), .X(n10158) );
  inv_x1_sg U8534 ( .A(n10158), .X(n10159) );
  inv_x1_sg U8535 ( .A(n10158), .X(n10160) );
  inv_x1_sg U8536 ( .A(n10159), .X(n10161) );
  inv_x1_sg U8537 ( .A(n10010), .X(n10162) );
  inv_x1_sg U8538 ( .A(n10588), .X(n10163) );
  inv_x1_sg U8539 ( .A(n10592), .X(n10164) );
  inv_x1_sg U8540 ( .A(n10011), .X(n10165) );
  inv_x1_sg U8541 ( .A(n10011), .X(n10166) );
  inv_x1_sg U8542 ( .A(n10011), .X(n10167) );
  inv_x1_sg U8543 ( .A(n10167), .X(n10168) );
  inv_x1_sg U8544 ( .A(n10167), .X(n10169) );
  inv_x1_sg U8545 ( .A(n10168), .X(n10170) );
  inv_x1_sg U8546 ( .A(n10012), .X(n10171) );
  inv_x1_sg U8547 ( .A(n10221), .X(n10172) );
  inv_x1_sg U8548 ( .A(n10172), .X(n10173) );
  inv_x1_sg U8549 ( .A(n10172), .X(n10174) );
  inv_x1_sg U8550 ( .A(n10139), .X(n10175) );
  inv_x1_sg U8551 ( .A(n10175), .X(n10176) );
  inv_x1_sg U8552 ( .A(n10175), .X(n10177) );
  inv_x1_sg U8553 ( .A(n10176), .X(n10178) );
  inv_x1_sg U8554 ( .A(n10013), .X(n10179) );
  inv_x1_sg U8555 ( .A(n10252), .X(n10180) );
  inv_x1_sg U8556 ( .A(n10180), .X(n10181) );
  inv_x1_sg U8557 ( .A(n10180), .X(n10182) );
  inv_x1_sg U8558 ( .A(n10182), .X(n10183) );
  inv_x1_sg U8559 ( .A(n10014), .X(n10184) );
  inv_x1_sg U8560 ( .A(n10532), .X(n10185) );
  inv_x1_sg U8561 ( .A(n10185), .X(n10186) );
  inv_x1_sg U8562 ( .A(n10185), .X(n10187) );
  inv_x1_sg U8563 ( .A(n10187), .X(n10188) );
  inv_x1_sg U8564 ( .A(n10015), .X(n10189) );
  inv_x1_sg U8565 ( .A(n10213), .X(n10190) );
  inv_x1_sg U8566 ( .A(n10190), .X(n10191) );
  inv_x1_sg U8567 ( .A(n10190), .X(n10192) );
  inv_x1_sg U8568 ( .A(n10542), .X(n10193) );
  inv_x1_sg U8569 ( .A(n10488), .X(n10194) );
  inv_x1_sg U8570 ( .A(n10289), .X(n10195) );
  inv_x1_sg U8571 ( .A(n10195), .X(n10196) );
  inv_x1_sg U8572 ( .A(n10194), .X(n10197) );
  inv_x1_sg U8573 ( .A(n10204), .X(n10198) );
  inv_x1_sg U8574 ( .A(n10198), .X(n10199) );
  inv_x1_sg U8575 ( .A(n10198), .X(n10200) );
  inv_x1_sg U8576 ( .A(n10199), .X(n10201) );
  inv_x1_sg U8577 ( .A(n10200), .X(n10202) );
  inv_x1_sg U8578 ( .A(n10088), .X(n10203) );
  inv_x1_sg U8579 ( .A(n10552), .X(n10204) );
  inv_x1_sg U8580 ( .A(n10203), .X(n10205) );
  inv_x1_sg U8581 ( .A(n10204), .X(n10206) );
  inv_x1_sg U8582 ( .A(n10680), .X(n10207) );
  inv_x1_sg U8583 ( .A(n10678), .X(n10208) );
  inv_x1_sg U8584 ( .A(n10248), .X(n10209) );
  inv_x1_sg U8585 ( .A(n8719), .X(n10210) );
  inv_x1_sg U8586 ( .A(n10569), .X(n10211) );
  inv_x1_sg U8587 ( .A(n10569), .X(n10212) );
  inv_x1_sg U8588 ( .A(n10210), .X(n10213) );
  inv_x1_sg U8589 ( .A(n10573), .X(n10214) );
  inv_x1_sg U8590 ( .A(n10573), .X(n10215) );
  inv_x1_sg U8591 ( .A(n10253), .X(n10216) );
  inv_x1_sg U8592 ( .A(n10577), .X(n10217) );
  inv_x1_sg U8593 ( .A(n10581), .X(n10218) );
  inv_x1_sg U8594 ( .A(n10218), .X(n10219) );
  inv_x1_sg U8595 ( .A(n10583), .X(n10220) );
  inv_x1_sg U8596 ( .A(n10218), .X(n10221) );
  inv_x1_sg U8597 ( .A(n10587), .X(n10222) );
  inv_x1_sg U8598 ( .A(n10071), .X(n10223) );
  inv_x1_sg U8599 ( .A(n10256), .X(n10224) );
  inv_x1_sg U8600 ( .A(n10254), .X(n10225) );
  inv_x1_sg U8601 ( .A(n10063), .X(n10226) );
  inv_x1_sg U8602 ( .A(n10226), .X(n10227) );
  inv_x1_sg U8603 ( .A(n10633), .X(n10228) );
  inv_x1_sg U8604 ( .A(n10110), .X(n10229) );
  inv_x1_sg U8605 ( .A(n10414), .X(n10230) );
  inv_x1_sg U8606 ( .A(n10418), .X(n10231) );
  inv_x1_sg U8607 ( .A(n10418), .X(n10232) );
  inv_x1_sg U8608 ( .A(n10423), .X(n10233) );
  inv_x1_sg U8609 ( .A(n10423), .X(n10234) );
  inv_x1_sg U8610 ( .A(n10427), .X(n10235) );
  inv_x1_sg U8611 ( .A(n10427), .X(n10236) );
  inv_x1_sg U8612 ( .A(n10030), .X(n10237) );
  inv_x1_sg U8613 ( .A(n10030), .X(n10238) );
  inv_x1_sg U8614 ( .A(n10115), .X(n10239) );
  inv_x1_sg U8615 ( .A(n10115), .X(n10240) );
  inv_x1_sg U8616 ( .A(n10438), .X(n10241) );
  inv_x1_sg U8617 ( .A(n10438), .X(n10242) );
  inv_x1_sg U8618 ( .A(n8712), .X(n10243) );
  inv_x1_sg U8619 ( .A(n10243), .X(n10244) );
  inv_x1_sg U8620 ( .A(n10243), .X(n10245) );
  inv_x1_sg U8621 ( .A(n10245), .X(n10246) );
  inv_x1_sg U8622 ( .A(n10016), .X(n10247) );
  inv_x1_sg U8623 ( .A(n10677), .X(n10248) );
  inv_x1_sg U8624 ( .A(n10068), .X(n10249) );
  inv_x1_sg U8625 ( .A(n10564), .X(n10250) );
  inv_x1_sg U8626 ( .A(n10568), .X(n10251) );
  inv_x1_sg U8627 ( .A(n10568), .X(n10252) );
  inv_x1_sg U8628 ( .A(n8719), .X(n10253) );
  inv_x1_sg U8629 ( .A(n10581), .X(n10254) );
  inv_x1_sg U8630 ( .A(n10582), .X(n10255) );
  inv_x1_sg U8631 ( .A(n10582), .X(n10256) );
  inv_x1_sg U8632 ( .A(n10685), .X(n10257) );
  inv_x1_sg U8633 ( .A(n10622), .X(n10258) );
  inv_x1_sg U8634 ( .A(n10072), .X(n10259) );
  inv_x1_sg U8635 ( .A(n10637), .X(n10260) );
  inv_x1_sg U8636 ( .A(n10641), .X(n10261) );
  inv_x1_sg U8637 ( .A(n10260), .X(n10262) );
  inv_x1_sg U8638 ( .A(n10443), .X(n10263) );
  inv_x1_sg U8639 ( .A(n10443), .X(n10264) );
  inv_x1_sg U8640 ( .A(n10210), .X(n10265) );
  inv_x1_sg U8641 ( .A(n10210), .X(n10266) );
  inv_x1_sg U8642 ( .A(n10070), .X(n10267) );
  inv_x1_sg U8643 ( .A(n10573), .X(n10268) );
  inv_x1_sg U8644 ( .A(n10251), .X(n10269) );
  inv_x1_sg U8645 ( .A(n10253), .X(n10270) );
  inv_x1_sg U8646 ( .A(n10218), .X(n10271) );
  inv_x1_sg U8647 ( .A(n10254), .X(n10272) );
  inv_x1_sg U8648 ( .A(n10587), .X(n10273) );
  inv_x1_sg U8649 ( .A(n10587), .X(n10274) );
  inv_x1_sg U8650 ( .A(n10256), .X(n10275) );
  inv_x1_sg U8651 ( .A(n10591), .X(n10276) );
  inv_x1_sg U8652 ( .A(n10120), .X(n10277) );
  inv_x1_sg U8653 ( .A(n10119), .X(n10278) );
  inv_x1_sg U8654 ( .A(n10125), .X(n10279) );
  inv_x1_sg U8655 ( .A(n10124), .X(n10280) );
  inv_x1_sg U8656 ( .A(n10006), .X(n10281) );
  inv_x1_sg U8657 ( .A(n10006), .X(n10282) );
  inv_x1_sg U8658 ( .A(n10007), .X(n10283) );
  inv_x1_sg U8659 ( .A(n10007), .X(n10284) );
  inv_x1_sg U8660 ( .A(n10138), .X(n10285) );
  inv_x1_sg U8661 ( .A(n10008), .X(n10286) );
  inv_x1_sg U8662 ( .A(n10143), .X(n10287) );
  inv_x1_sg U8663 ( .A(n10009), .X(n10288) );
  inv_x1_sg U8664 ( .A(n10542), .X(n10289) );
  inv_x1_sg U8665 ( .A(n10150), .X(n10290) );
  inv_x1_sg U8666 ( .A(n10149), .X(n10291) );
  inv_x1_sg U8667 ( .A(n10154), .X(n10292) );
  inv_x1_sg U8668 ( .A(n10010), .X(n10293) );
  inv_x1_sg U8669 ( .A(n10160), .X(n10294) );
  inv_x1_sg U8670 ( .A(n10164), .X(n10295) );
  inv_x1_sg U8671 ( .A(n10163), .X(n10296) );
  inv_x1_sg U8672 ( .A(n10168), .X(n10297) );
  inv_x1_sg U8673 ( .A(n10169), .X(n10298) );
  inv_x1_sg U8674 ( .A(n10517), .X(n10299) );
  inv_x1_sg U8675 ( .A(n10517), .X(n10300) );
  inv_x1_sg U8676 ( .A(n10177), .X(n10301) );
  inv_x1_sg U8677 ( .A(n10177), .X(n10302) );
  inv_x1_sg U8678 ( .A(n10181), .X(n10303) );
  inv_x1_sg U8679 ( .A(n10181), .X(n10304) );
  inv_x1_sg U8680 ( .A(n10186), .X(n10305) );
  inv_x1_sg U8681 ( .A(n10186), .X(n10306) );
  inv_x1_sg U8682 ( .A(n10537), .X(n10307) );
  inv_x1_sg U8683 ( .A(n10537), .X(n10308) );
  inv_x1_sg U8684 ( .A(n10195), .X(n10309) );
  inv_x1_sg U8685 ( .A(n10194), .X(n10310) );
  inv_x1_sg U8686 ( .A(n10257), .X(n10311) );
  inv_x1_sg U8687 ( .A(n10623), .X(n10312) );
  inv_x1_sg U8688 ( .A(n10651), .X(n10313) );
  inv_x1_sg U8689 ( .A(n10096), .X(n10314) );
  inv_x1_sg U8690 ( .A(n10611), .X(n10315) );
  inv_x1_sg U8691 ( .A(n10082), .X(n10316) );
  inv_x1_sg U8692 ( .A(n10610), .X(n10317) );
  inv_x1_sg U8693 ( .A(n10078), .X(n10318) );
  inv_x1_sg U8694 ( .A(n10617), .X(n10319) );
  inv_x1_sg U8695 ( .A(n10319), .X(n10320) );
  inv_x1_sg U8696 ( .A(n10319), .X(n10321) );
  inv_x1_sg U8697 ( .A(n10319), .X(n10322) );
  inv_x1_sg U8698 ( .A(n10082), .X(n10323) );
  inv_x1_sg U8699 ( .A(n10609), .X(n10324) );
  inv_x1_sg U8700 ( .A(n10620), .X(n10325) );
  inv_x1_sg U8701 ( .A(n10325), .X(n10326) );
  inv_x1_sg U8702 ( .A(n10325), .X(n10327) );
  inv_x1_sg U8703 ( .A(n10325), .X(n10328) );
  inv_x1_sg U8704 ( .A(n10085), .X(n10329) );
  inv_x1_sg U8705 ( .A(n10257), .X(n10330) );
  inv_x1_sg U8706 ( .A(n10626), .X(n10331) );
  inv_x1_sg U8707 ( .A(n10331), .X(n10332) );
  inv_x1_sg U8708 ( .A(n10331), .X(n10333) );
  inv_x1_sg U8709 ( .A(n10331), .X(n10334) );
  inv_x1_sg U8710 ( .A(n10085), .X(n10335) );
  inv_x1_sg U8711 ( .A(n10257), .X(n10336) );
  inv_x1_sg U8712 ( .A(n10629), .X(n10337) );
  inv_x1_sg U8713 ( .A(n10337), .X(n10338) );
  inv_x1_sg U8714 ( .A(n10337), .X(n10339) );
  inv_x1_sg U8715 ( .A(n10337), .X(n10340) );
  inv_x1_sg U8716 ( .A(n10639), .X(n10341) );
  inv_x1_sg U8717 ( .A(n10639), .X(n10342) );
  inv_x1_sg U8718 ( .A(n10103), .X(n10343) );
  inv_x1_sg U8719 ( .A(n10665), .X(n10344) );
  inv_x1_sg U8720 ( .A(n10373), .X(n10345) );
  inv_x1_sg U8721 ( .A(n10345), .X(n10346) );
  inv_x1_sg U8722 ( .A(n10345), .X(n10347) );
  inv_x1_sg U8723 ( .A(n10345), .X(n10348) );
  inv_x1_sg U8724 ( .A(n10099), .X(n10349) );
  inv_x1_sg U8725 ( .A(n10683), .X(n10350) );
  inv_x1_sg U8726 ( .A(n10342), .X(n10351) );
  inv_x1_sg U8727 ( .A(n10351), .X(n10352) );
  inv_x1_sg U8728 ( .A(n10351), .X(n10353) );
  inv_x1_sg U8729 ( .A(n10351), .X(n10354) );
  inv_x1_sg U8730 ( .A(n10103), .X(n10355) );
  inv_x1_sg U8731 ( .A(n10665), .X(n10356) );
  inv_x1_sg U8732 ( .A(n10095), .X(n10357) );
  inv_x1_sg U8733 ( .A(n10357), .X(n10358) );
  inv_x1_sg U8734 ( .A(n10357), .X(n10359) );
  inv_x1_sg U8735 ( .A(n10357), .X(n10360) );
  inv_x1_sg U8736 ( .A(n10683), .X(n10361) );
  inv_x1_sg U8737 ( .A(n10663), .X(n10362) );
  inv_x1_sg U8738 ( .A(n10098), .X(n10363) );
  inv_x1_sg U8739 ( .A(n10363), .X(n10364) );
  inv_x1_sg U8740 ( .A(n10363), .X(n10365) );
  inv_x1_sg U8741 ( .A(n10363), .X(n10366) );
  inv_x1_sg U8742 ( .A(n10653), .X(n10367) );
  inv_x1_sg U8743 ( .A(n10653), .X(n10368) );
  inv_x1_sg U8744 ( .A(n10107), .X(n10369) );
  inv_x1_sg U8745 ( .A(n10369), .X(n10370) );
  inv_x1_sg U8746 ( .A(n10369), .X(n10371) );
  inv_x1_sg U8747 ( .A(n10369), .X(n10372) );
  inv_x1_sg U8748 ( .A(n10640), .X(n10373) );
  inv_x1_sg U8749 ( .A(n10665), .X(n10374) );
  inv_x1_sg U8750 ( .A(n10668), .X(n10375) );
  inv_x1_sg U8751 ( .A(n10375), .X(n10376) );
  inv_x1_sg U8752 ( .A(n10375), .X(n10377) );
  inv_x1_sg U8753 ( .A(n10375), .X(n10378) );
  inv_x1_sg U8754 ( .A(n10103), .X(n10379) );
  inv_x1_sg U8755 ( .A(n10652), .X(n10380) );
  inv_x1_sg U8756 ( .A(n10671), .X(n10381) );
  inv_x1_sg U8757 ( .A(n10381), .X(n10382) );
  inv_x1_sg U8758 ( .A(n10381), .X(n10383) );
  inv_x1_sg U8759 ( .A(n10381), .X(n10384) );
  inv_x1_sg U8760 ( .A(n10612), .X(n10385) );
  inv_x1_sg U8761 ( .A(n10385), .X(n10386) );
  inv_x1_sg U8762 ( .A(n10385), .X(n10387) );
  inv_x1_sg U8763 ( .A(n10385), .X(n10388) );
  inv_x1_sg U8764 ( .A(n10598), .X(n10389) );
  inv_x1_sg U8765 ( .A(n10599), .X(n10390) );
  inv_x1_sg U8766 ( .A(n10606), .X(n10391) );
  inv_x1_sg U8767 ( .A(n10391), .X(n10392) );
  inv_x1_sg U8768 ( .A(n10391), .X(n10393) );
  inv_x1_sg U8769 ( .A(n10391), .X(n10394) );
  inv_x1_sg U8770 ( .A(n10598), .X(n10395) );
  inv_x1_sg U8771 ( .A(n10072), .X(n10396) );
  inv_x1_sg U8772 ( .A(n10603), .X(n10397) );
  inv_x1_sg U8773 ( .A(n10397), .X(n10398) );
  inv_x1_sg U8774 ( .A(n10397), .X(n10399) );
  inv_x1_sg U8775 ( .A(n10397), .X(n10400) );
  inv_x1_sg U8776 ( .A(n10076), .X(n10401) );
  inv_x1_sg U8777 ( .A(n10076), .X(n10402) );
  inv_x1_sg U8778 ( .A(n10642), .X(n10403) );
  inv_x1_sg U8779 ( .A(n10403), .X(n10404) );
  inv_x1_sg U8780 ( .A(n10403), .X(n10405) );
  inv_x1_sg U8781 ( .A(n10403), .X(n10406) );
  inv_x1_sg U8782 ( .A(n10600), .X(n10407) );
  inv_x1_sg U8783 ( .A(n10407), .X(n10408) );
  inv_x1_sg U8784 ( .A(n10407), .X(n10409) );
  inv_x1_sg U8785 ( .A(n10407), .X(n10410) );
  inv_x1_sg U8786 ( .A(n10407), .X(n10411) );
  inv_x1_sg U8787 ( .A(n10680), .X(n10412) );
  inv_x1_sg U8788 ( .A(n10678), .X(n10413) );
  inv_x1_sg U8789 ( .A(n10559), .X(n10414) );
  inv_x1_sg U8790 ( .A(n10110), .X(n10415) );
  inv_x1_sg U8791 ( .A(n10414), .X(n10416) );
  inv_x1_sg U8792 ( .A(n10110), .X(n10417) );
  inv_x1_sg U8793 ( .A(n10416), .X(n10418) );
  inv_x1_sg U8794 ( .A(n10112), .X(n10419) );
  inv_x1_sg U8795 ( .A(n10112), .X(n10420) );
  inv_x1_sg U8796 ( .A(n10112), .X(n10421) );
  inv_x1_sg U8797 ( .A(n10418), .X(n10422) );
  inv_x1_sg U8798 ( .A(n10413), .X(n10423) );
  inv_x1_sg U8799 ( .A(n10114), .X(n10424) );
  inv_x1_sg U8800 ( .A(n10114), .X(n10425) );
  inv_x1_sg U8801 ( .A(n10423), .X(n10426) );
  inv_x1_sg U8802 ( .A(n10560), .X(n10427) );
  inv_x1_sg U8803 ( .A(n10427), .X(n10428) );
  inv_x1_sg U8804 ( .A(n10427), .X(n10429) );
  inv_x1_sg U8805 ( .A(n10118), .X(n10430) );
  inv_x1_sg U8806 ( .A(n10036), .X(n10431) );
  inv_x1_sg U8807 ( .A(n10195), .X(n10432) );
  inv_x1_sg U8808 ( .A(n10123), .X(n10433) );
  inv_x1_sg U8809 ( .A(n10115), .X(n10434) );
  inv_x1_sg U8810 ( .A(n10123), .X(n10435) );
  inv_x1_sg U8811 ( .A(n10199), .X(n10436) );
  inv_x1_sg U8812 ( .A(n10200), .X(n10437) );
  inv_x1_sg U8813 ( .A(n10201), .X(n10438) );
  inv_x1_sg U8814 ( .A(n10116), .X(n10439) );
  inv_x1_sg U8815 ( .A(n10116), .X(n10440) );
  inv_x1_sg U8816 ( .A(n10116), .X(n10441) );
  inv_x1_sg U8817 ( .A(n10438), .X(n10442) );
  inv_x1_sg U8818 ( .A(n10547), .X(n10443) );
  inv_x1_sg U8819 ( .A(n10117), .X(n10444) );
  inv_x1_sg U8820 ( .A(n10117), .X(n10445) );
  inv_x1_sg U8821 ( .A(n10443), .X(n10446) );
  inv_x1_sg U8822 ( .A(n10443), .X(n10447) );
  inv_x1_sg U8823 ( .A(n10226), .X(n10448) );
  inv_x1_sg U8824 ( .A(n10633), .X(n10449) );
  inv_x1_sg U8825 ( .A(n10203), .X(n10450) );
  inv_x1_sg U8826 ( .A(n10204), .X(n10451) );
  inv_x1_sg U8827 ( .A(n10205), .X(n10452) );
  inv_x1_sg U8828 ( .A(n10120), .X(n10453) );
  inv_x1_sg U8829 ( .A(n10119), .X(n10454) );
  inv_x1_sg U8830 ( .A(n10120), .X(n10455) );
  inv_x1_sg U8831 ( .A(n10119), .X(n10456) );
  inv_x1_sg U8832 ( .A(n10125), .X(n10457) );
  inv_x1_sg U8833 ( .A(n10005), .X(n10458) );
  inv_x1_sg U8834 ( .A(n10125), .X(n10459) );
  inv_x1_sg U8835 ( .A(n10005), .X(n10460) );
  inv_x1_sg U8836 ( .A(n10256), .X(n10461) );
  inv_x1_sg U8837 ( .A(n10591), .X(n10462) );
  inv_x1_sg U8838 ( .A(n10129), .X(n10463) );
  inv_x1_sg U8839 ( .A(n10006), .X(n10464) );
  inv_x1_sg U8840 ( .A(n10130), .X(n10465) );
  inv_x1_sg U8841 ( .A(n10129), .X(n10466) );
  inv_x1_sg U8842 ( .A(n10134), .X(n10467) );
  inv_x1_sg U8843 ( .A(n10007), .X(n10468) );
  inv_x1_sg U8844 ( .A(n10130), .X(n10469) );
  inv_x1_sg U8845 ( .A(n10134), .X(n10470) );
  inv_x1_sg U8846 ( .A(n10071), .X(n10471) );
  inv_x1_sg U8847 ( .A(n10071), .X(n10472) );
  inv_x1_sg U8848 ( .A(n10577), .X(n10473) );
  inv_x1_sg U8849 ( .A(n10253), .X(n10474) );
  inv_x1_sg U8850 ( .A(n10138), .X(n10475) );
  inv_x1_sg U8851 ( .A(n10138), .X(n10476) );
  inv_x1_sg U8852 ( .A(n10008), .X(n10477) );
  inv_x1_sg U8853 ( .A(n10139), .X(n10478) );
  inv_x1_sg U8854 ( .A(n10143), .X(n10479) );
  inv_x1_sg U8855 ( .A(n10143), .X(n10480) );
  inv_x1_sg U8856 ( .A(n10009), .X(n10481) );
  inv_x1_sg U8857 ( .A(n10139), .X(n10482) );
  inv_x1_sg U8858 ( .A(n10070), .X(n10483) );
  inv_x1_sg U8859 ( .A(n10070), .X(n10484) );
  inv_x1_sg U8860 ( .A(n10564), .X(n10485) );
  inv_x1_sg U8861 ( .A(n10068), .X(n10486) );
  inv_x1_sg U8862 ( .A(n10068), .X(n10487) );
  inv_x1_sg U8863 ( .A(n10542), .X(n10488) );
  inv_x1_sg U8864 ( .A(n10153), .X(n10489) );
  inv_x1_sg U8865 ( .A(n10148), .X(n10490) );
  inv_x1_sg U8866 ( .A(n10016), .X(n10491) );
  inv_x1_sg U8867 ( .A(n10245), .X(n10492) );
  inv_x1_sg U8868 ( .A(n10492), .X(n10493) );
  inv_x1_sg U8869 ( .A(n10150), .X(n10494) );
  inv_x1_sg U8870 ( .A(n10017), .X(n10495) );
  inv_x1_sg U8871 ( .A(n10150), .X(n10496) );
  inv_x1_sg U8872 ( .A(n10149), .X(n10497) );
  inv_x1_sg U8873 ( .A(n10491), .X(n10498) );
  inv_x1_sg U8874 ( .A(n10155), .X(n10499) );
  inv_x1_sg U8875 ( .A(n10154), .X(n10500) );
  inv_x1_sg U8876 ( .A(n10155), .X(n10501) );
  inv_x1_sg U8877 ( .A(n10154), .X(n10502) );
  inv_x1_sg U8878 ( .A(n10159), .X(n10503) );
  inv_x1_sg U8879 ( .A(n10160), .X(n10504) );
  inv_x1_sg U8880 ( .A(n10160), .X(n10505) );
  inv_x1_sg U8881 ( .A(n10159), .X(n10506) );
  inv_x1_sg U8882 ( .A(n10164), .X(n10507) );
  inv_x1_sg U8883 ( .A(n10163), .X(n10508) );
  inv_x1_sg U8884 ( .A(n10163), .X(n10509) );
  inv_x1_sg U8885 ( .A(n10164), .X(n10510) );
  inv_x1_sg U8886 ( .A(n10583), .X(n10511) );
  inv_x1_sg U8887 ( .A(n10583), .X(n10512) );
  inv_x1_sg U8888 ( .A(n10012), .X(n10513) );
  inv_x1_sg U8889 ( .A(n10168), .X(n10514) );
  inv_x1_sg U8890 ( .A(n10169), .X(n10515) );
  inv_x1_sg U8891 ( .A(n10169), .X(n10516) );
  inv_x1_sg U8892 ( .A(n10584), .X(n10517) );
  inv_x1_sg U8893 ( .A(n10130), .X(n10518) );
  inv_x1_sg U8894 ( .A(n10172), .X(n10519) );
  inv_x1_sg U8895 ( .A(n10172), .X(n10520) );
  inv_x1_sg U8896 ( .A(n10010), .X(n10521) );
  inv_x1_sg U8897 ( .A(n10177), .X(n10522) );
  inv_x1_sg U8898 ( .A(n10176), .X(n10523) );
  inv_x1_sg U8899 ( .A(n10013), .X(n10524) );
  inv_x1_sg U8900 ( .A(n10176), .X(n10525) );
  inv_x1_sg U8901 ( .A(n10181), .X(n10526) );
  inv_x1_sg U8902 ( .A(n10182), .X(n10527) );
  inv_x1_sg U8903 ( .A(n10014), .X(n10528) );
  inv_x1_sg U8904 ( .A(n10182), .X(n10529) );
  inv_x1_sg U8905 ( .A(n10251), .X(n10530) );
  inv_x1_sg U8906 ( .A(n10569), .X(n10531) );
  inv_x1_sg U8907 ( .A(n10571), .X(n10532) );
  inv_x1_sg U8908 ( .A(n10186), .X(n10533) );
  inv_x1_sg U8909 ( .A(n10187), .X(n10534) );
  inv_x1_sg U8910 ( .A(n10015), .X(n10535) );
  inv_x1_sg U8911 ( .A(n10187), .X(n10536) );
  inv_x1_sg U8912 ( .A(n10570), .X(n10537) );
  inv_x1_sg U8913 ( .A(n10190), .X(n10538) );
  inv_x1_sg U8914 ( .A(n10190), .X(n10539) );
  inv_x1_sg U8915 ( .A(n10014), .X(n10540) );
  inv_x1_sg U8916 ( .A(n10181), .X(n10541) );
  inv_x1_sg U8917 ( .A(n10565), .X(n10542) );
  inv_x1_sg U8918 ( .A(n10195), .X(n10543) );
  inv_x1_sg U8919 ( .A(n10194), .X(n10544) );
  inv_x1_sg U8920 ( .A(n10194), .X(n10545) );
  inv_x1_sg U8921 ( .A(n10199), .X(n10546) );
  inv_x1_sg U8922 ( .A(n10200), .X(n10547) );
  inv_x1_sg U8923 ( .A(n10199), .X(n10548) );
  inv_x1_sg U8924 ( .A(n10200), .X(n10549) );
  inv_x1_sg U8925 ( .A(n10035), .X(n10550) );
  inv_x1_sg U8926 ( .A(n10204), .X(n10551) );
  inv_x1_sg U8927 ( .A(n10203), .X(n10552) );
  inv_x1_sg U8928 ( .A(n10244), .X(n10553) );
  inv_x1_sg U8929 ( .A(n10244), .X(n10554) );
  inv_x1_sg U8930 ( .A(n10244), .X(n10555) );
  inv_x1_sg U8931 ( .A(n10016), .X(n10556) );
  inv_x1_sg U8932 ( .A(n10681), .X(n10557) );
  inv_x1_sg U8933 ( .A(n10066), .X(n10558) );
  inv_x1_sg U8934 ( .A(n10066), .X(n10559) );
  inv_x1_sg U8935 ( .A(n10557), .X(n10560) );
  inv_x1_sg U8936 ( .A(n10557), .X(n10561) );
  inv_x1_sg U8937 ( .A(n10678), .X(n10562) );
  inv_x1_sg U8938 ( .A(n10680), .X(n10563) );
  inv_x1_sg U8939 ( .A(n10677), .X(n10564) );
  inv_x1_sg U8940 ( .A(n10564), .X(n10565) );
  inv_x1_sg U8941 ( .A(n10248), .X(n10566) );
  inv_x1_sg U8942 ( .A(n10248), .X(n10567) );
  nor_x1_sg U8943 ( .A(n10682), .B(n10409), .X(n10568) );
  inv_x1_sg U8944 ( .A(n8719), .X(n10569) );
  inv_x1_sg U8945 ( .A(n10251), .X(n10570) );
  inv_x1_sg U8946 ( .A(n10569), .X(n10571) );
  inv_x1_sg U8947 ( .A(n10251), .X(n10572) );
  inv_x1_sg U8948 ( .A(n10568), .X(n10573) );
  inv_x1_sg U8949 ( .A(n10252), .X(n10574) );
  inv_x1_sg U8950 ( .A(n10070), .X(n10575) );
  inv_x1_sg U8951 ( .A(n10573), .X(n10576) );
  inv_x1_sg U8952 ( .A(n8719), .X(n10577) );
  inv_x1_sg U8953 ( .A(n10253), .X(n10578) );
  inv_x1_sg U8954 ( .A(n10577), .X(n10579) );
  inv_x1_sg U8955 ( .A(n10577), .X(n10580) );
  nor_x1_sg U8956 ( .A(n10404), .B(n10684), .X(n10581) );
  nor_x1_sg U8957 ( .A(n10094), .B(n10684), .X(n10582) );
  inv_x1_sg U8958 ( .A(n10581), .X(n10583) );
  inv_x1_sg U8959 ( .A(n10254), .X(n10584) );
  inv_x1_sg U8960 ( .A(n10583), .X(n10585) );
  inv_x1_sg U8961 ( .A(n10254), .X(n10586) );
  inv_x1_sg U8962 ( .A(n10582), .X(n10587) );
  inv_x1_sg U8963 ( .A(n10255), .X(n10588) );
  inv_x1_sg U8964 ( .A(n10071), .X(n10589) );
  inv_x1_sg U8965 ( .A(n10587), .X(n10590) );
  inv_x1_sg U8966 ( .A(n10581), .X(n10591) );
  inv_x1_sg U8967 ( .A(n10256), .X(n10592) );
  inv_x1_sg U8968 ( .A(n10591), .X(n10593) );
  inv_x1_sg U8969 ( .A(n10591), .X(n10594) );
  nor_x1_sg U8970 ( .A(n9359), .B(n8715), .X(n10595) );
  nor_x1_sg U8971 ( .A(n9359), .B(n8715), .X(n10596) );
  inv_x1_sg U8972 ( .A(n10080), .X(n10597) );
  inv_x1_sg U8973 ( .A(n10595), .X(n10598) );
  inv_x1_sg U8974 ( .A(n10595), .X(n10599) );
  inv_x1_sg U8975 ( .A(n10597), .X(n10600) );
  inv_x1_sg U8976 ( .A(n10072), .X(n10601) );
  inv_x1_sg U8977 ( .A(n10597), .X(n10602) );
  inv_x1_sg U8978 ( .A(n10598), .X(n10603) );
  inv_x1_sg U8979 ( .A(n10597), .X(n10604) );
  inv_x1_sg U8980 ( .A(n10599), .X(n10605) );
  inv_x1_sg U8981 ( .A(n10599), .X(n10606) );
  inv_x1_sg U8982 ( .A(n10072), .X(n10607) );
  inv_x1_sg U8983 ( .A(n10076), .X(n10608) );
  inv_x1_sg U8984 ( .A(n10596), .X(n10609) );
  inv_x1_sg U8985 ( .A(n10596), .X(n10610) );
  inv_x1_sg U8986 ( .A(n10021), .X(n10611) );
  inv_x1_sg U8987 ( .A(n10609), .X(n10612) );
  inv_x1_sg U8988 ( .A(n10082), .X(n10613) );
  inv_x1_sg U8989 ( .A(n10078), .X(n10614) );
  inv_x1_sg U8990 ( .A(n10609), .X(n10615) );
  inv_x1_sg U8991 ( .A(n10611), .X(n10616) );
  inv_x1_sg U8992 ( .A(n10610), .X(n10617) );
  inv_x1_sg U8993 ( .A(n10078), .X(n10618) );
  inv_x1_sg U8994 ( .A(n10610), .X(n10619) );
  inv_x1_sg U8995 ( .A(n10611), .X(n10620) );
  inv_x1_sg U8996 ( .A(n10685), .X(n10621) );
  inv_x1_sg U8997 ( .A(n10685), .X(n10622) );
  inv_x1_sg U8998 ( .A(n10685), .X(n10623) );
  inv_x1_sg U8999 ( .A(n10623), .X(n10624) );
  inv_x1_sg U9000 ( .A(n10621), .X(n10625) );
  inv_x1_sg U9001 ( .A(n10337), .X(n10626) );
  inv_x1_sg U9002 ( .A(n10623), .X(n10627) );
  inv_x1_sg U9003 ( .A(n10621), .X(n10628) );
  inv_x1_sg U9004 ( .A(n10622), .X(n10629) );
  inv_x1_sg U9005 ( .A(n10623), .X(n10630) );
  inv_x1_sg U9006 ( .A(n10621), .X(n10631) );
  inv_x1_sg U9007 ( .A(n10085), .X(n10632) );
  inv_x1_sg U9008 ( .A(n10676), .X(n10633) );
  inv_x1_sg U9009 ( .A(n10226), .X(n10634) );
  inv_x1_sg U9010 ( .A(n10226), .X(n10635) );
  inv_x1_sg U9011 ( .A(n10633), .X(n10636) );
  nor_x1_sg U9012 ( .A(n10676), .B(n10682), .X(n10637) );
  nor_x1_sg U9013 ( .A(n10553), .B(n10684), .X(n10638) );
  inv_x1_sg U9014 ( .A(n10637), .X(n10639) );
  inv_x1_sg U9015 ( .A(n10022), .X(n10640) );
  inv_x1_sg U9016 ( .A(n10638), .X(n10641) );
  inv_x1_sg U9017 ( .A(n10639), .X(n10642) );
  inv_x1_sg U9018 ( .A(n10090), .X(n10643) );
  inv_x1_sg U9019 ( .A(n10090), .X(n10644) );
  inv_x1_sg U9020 ( .A(n10651), .X(n10645) );
  inv_x1_sg U9021 ( .A(n10096), .X(n10646) );
  inv_x1_sg U9022 ( .A(n10640), .X(n10647) );
  inv_x1_sg U9023 ( .A(n10641), .X(n10648) );
  inv_x1_sg U9024 ( .A(n10652), .X(n10649) );
  inv_x1_sg U9025 ( .A(n10641), .X(n10650) );
  inv_x1_sg U9026 ( .A(n8716), .X(n10651) );
  inv_x1_sg U9027 ( .A(n10638), .X(n10652) );
  inv_x1_sg U9028 ( .A(n10637), .X(n10653) );
  inv_x1_sg U9029 ( .A(n10651), .X(n10654) );
  inv_x1_sg U9030 ( .A(n10096), .X(n10655) );
  inv_x1_sg U9031 ( .A(n10651), .X(n10656) );
  inv_x1_sg U9032 ( .A(n10652), .X(n10657) );
  inv_x1_sg U9033 ( .A(n10099), .X(n10658) );
  inv_x1_sg U9034 ( .A(n10652), .X(n10659) );
  inv_x1_sg U9035 ( .A(n10101), .X(n10660) );
  inv_x1_sg U9036 ( .A(n10653), .X(n10661) );
  inv_x1_sg U9037 ( .A(n10653), .X(n10662) );
  inv_x1_sg U9038 ( .A(n10638), .X(n10663) );
  inv_x1_sg U9039 ( .A(n10637), .X(n10664) );
  inv_x1_sg U9040 ( .A(n8716), .X(n10665) );
  inv_x1_sg U9041 ( .A(n10663), .X(n10666) );
  inv_x1_sg U9042 ( .A(n10260), .X(n10667) );
  inv_x1_sg U9043 ( .A(n10663), .X(n10668) );
  inv_x1_sg U9044 ( .A(n10664), .X(n10669) );
  inv_x1_sg U9045 ( .A(n10099), .X(n10670) );
  inv_x1_sg U9046 ( .A(n10664), .X(n10671) );
  inv_x1_sg U9047 ( .A(n10664), .X(n10672) );
  inv_x1_sg U9048 ( .A(n10260), .X(n10673) );
  inv_x1_sg U9049 ( .A(n10683), .X(n10674) );
  nor_x1_sg U9050 ( .A(n12286), .B(state[1]), .X(n10675) );
  inv_x1_sg U9051 ( .A(n10675), .X(n10676) );
  inv_x1_sg U9052 ( .A(n10676), .X(n10677) );
  inv_x1_sg U9053 ( .A(n8712), .X(n10678) );
  inv_x1_sg U9054 ( .A(n10678), .X(n10679) );
  inv_x1_sg U9055 ( .A(n10675), .X(n10680) );
  inv_x1_sg U9056 ( .A(n10680), .X(n10681) );
  inv_x1_sg U9057 ( .A(n10638), .X(n10683) );
  inv_x1_sg U9058 ( .A(n8710), .X(n10684) );
  nor_x1_sg U9059 ( .A(n12286), .B(state[1]), .X(n8712) );
  nand_x1_sg U9060 ( .A(n10000), .B(n9999), .X(n3866) );
  nand_x1_sg U9061 ( .A(n9998), .B(n9997), .X(n3867) );
  nand_x1_sg U9062 ( .A(n9996), .B(n9995), .X(n3868) );
  nand_x1_sg U9063 ( .A(n9994), .B(n9993), .X(n3869) );
  nand_x1_sg U9064 ( .A(n9992), .B(n9991), .X(n3870) );
  nand_x1_sg U9065 ( .A(n9990), .B(n9989), .X(n3871) );
  nand_x1_sg U9066 ( .A(n9988), .B(n9987), .X(n3872) );
  nand_x1_sg U9067 ( .A(n9986), .B(n9985), .X(n3873) );
  nand_x1_sg U9068 ( .A(n9984), .B(n9983), .X(n3874) );
  nand_x1_sg U9069 ( .A(n9982), .B(n9981), .X(n3875) );
  nand_x1_sg U9070 ( .A(n9980), .B(n9979), .X(n3876) );
  nand_x1_sg U9071 ( .A(n9978), .B(n9977), .X(n3877) );
  nand_x1_sg U9072 ( .A(n9976), .B(n9975), .X(n3878) );
  nand_x1_sg U9073 ( .A(n9974), .B(n9973), .X(n3879) );
  nand_x1_sg U9074 ( .A(n9972), .B(n9971), .X(n3880) );
  nand_x1_sg U9075 ( .A(n9970), .B(n9969), .X(n3881) );
  nand_x1_sg U9076 ( .A(n9968), .B(n9967), .X(n3882) );
  nand_x1_sg U9077 ( .A(n9966), .B(n9965), .X(n3883) );
  nand_x1_sg U9078 ( .A(n9964), .B(n9963), .X(n3884) );
  nand_x1_sg U9079 ( .A(n9962), .B(n9961), .X(n3885) );
  nand_x1_sg U9080 ( .A(n9960), .B(n9959), .X(n3886) );
  nand_x1_sg U9081 ( .A(n9958), .B(n9957), .X(n3887) );
  nand_x1_sg U9082 ( .A(n9956), .B(n9955), .X(n3888) );
  nand_x1_sg U9083 ( .A(n9954), .B(n9953), .X(n3889) );
  nand_x1_sg U9084 ( .A(n9952), .B(n9951), .X(n3890) );
  nand_x1_sg U9085 ( .A(n9950), .B(n9949), .X(n3891) );
  nand_x1_sg U9086 ( .A(n9948), .B(n9947), .X(n3892) );
  nand_x1_sg U9087 ( .A(n9945), .B(n9946), .X(n3893) );
  nand_x1_sg U9088 ( .A(n9944), .B(n9943), .X(n3894) );
  nand_x1_sg U9089 ( .A(n9942), .B(n9941), .X(n3895) );
  nand_x1_sg U9090 ( .A(n9940), .B(n9939), .X(n3896) );
  nand_x1_sg U9091 ( .A(n9938), .B(n9937), .X(n3897) );
  nand_x1_sg U9092 ( .A(n9936), .B(n9935), .X(n3898) );
  nand_x1_sg U9093 ( .A(n9934), .B(n9933), .X(n3899) );
  nand_x1_sg U9094 ( .A(n9932), .B(n9931), .X(n3900) );
  nand_x1_sg U9095 ( .A(n9930), .B(n9929), .X(n3901) );
  nand_x1_sg U9096 ( .A(n9928), .B(n9927), .X(n3902) );
  nand_x1_sg U9097 ( .A(n9926), .B(n9925), .X(n3903) );
  nand_x1_sg U9098 ( .A(n9924), .B(n9923), .X(n3904) );
  nand_x1_sg U9099 ( .A(n9922), .B(n9921), .X(n3905) );
  nand_x1_sg U9100 ( .A(n9920), .B(n9919), .X(n3906) );
  nand_x1_sg U9101 ( .A(n9918), .B(n9917), .X(n3907) );
  nand_x1_sg U9102 ( .A(n9916), .B(n9915), .X(n3908) );
  nand_x1_sg U9103 ( .A(n9914), .B(n9913), .X(n3909) );
  nand_x1_sg U9104 ( .A(n9912), .B(n9911), .X(n3910) );
  nand_x1_sg U9105 ( .A(n9910), .B(n9909), .X(n3911) );
  nand_x1_sg U9106 ( .A(n9908), .B(n9907), .X(n3912) );
  nand_x1_sg U9107 ( .A(n9906), .B(n9905), .X(n3913) );
  nand_x1_sg U9108 ( .A(n9904), .B(n9903), .X(n3914) );
  nand_x1_sg U9109 ( .A(n9902), .B(n9901), .X(n3915) );
  nand_x1_sg U9110 ( .A(n9900), .B(n9899), .X(n3916) );
  nand_x1_sg U9111 ( .A(n9898), .B(n9897), .X(n3917) );
  nand_x1_sg U9112 ( .A(n9896), .B(n9895), .X(n3918) );
  nand_x1_sg U9113 ( .A(n9894), .B(n9893), .X(n3919) );
  nand_x1_sg U9114 ( .A(n9892), .B(n9891), .X(n3920) );
  nand_x1_sg U9115 ( .A(n9890), .B(n9889), .X(n3921) );
  nand_x1_sg U9116 ( .A(n9888), .B(n9887), .X(n3922) );
  nand_x1_sg U9117 ( .A(n9886), .B(n9885), .X(n3923) );
  nand_x1_sg U9118 ( .A(n9884), .B(n9883), .X(n3924) );
  nand_x1_sg U9119 ( .A(n9882), .B(n9881), .X(n3925) );
  nand_x1_sg U9120 ( .A(n9880), .B(n9879), .X(n3926) );
  nand_x1_sg U9121 ( .A(n9878), .B(n9877), .X(n3927) );
  nand_x1_sg U9122 ( .A(n9876), .B(n9875), .X(n3928) );
  nand_x1_sg U9123 ( .A(n9874), .B(n9873), .X(n3929) );
  nand_x1_sg U9124 ( .A(n9872), .B(n9871), .X(n3930) );
  nand_x1_sg U9125 ( .A(n9870), .B(n9869), .X(n3931) );
  nand_x1_sg U9126 ( .A(n9868), .B(n9867), .X(n3932) );
  nand_x1_sg U9127 ( .A(n9866), .B(n9865), .X(n3933) );
  nand_x1_sg U9128 ( .A(n9864), .B(n9863), .X(n3934) );
  nand_x1_sg U9129 ( .A(n9862), .B(n9861), .X(n3935) );
  nand_x1_sg U9130 ( .A(n9860), .B(n9859), .X(n3936) );
  nand_x1_sg U9131 ( .A(n9858), .B(n9857), .X(n3937) );
  nand_x1_sg U9132 ( .A(n9856), .B(n9855), .X(n3938) );
  nand_x1_sg U9133 ( .A(n9854), .B(n9853), .X(n3939) );
  nand_x1_sg U9134 ( .A(n9852), .B(n9851), .X(n3940) );
  nand_x1_sg U9135 ( .A(n9850), .B(n9849), .X(n3941) );
  nand_x1_sg U9136 ( .A(n9848), .B(n9847), .X(n3942) );
  nand_x1_sg U9137 ( .A(n9846), .B(n9845), .X(n3943) );
  nand_x1_sg U9138 ( .A(n9844), .B(n9843), .X(n3944) );
  nand_x1_sg U9139 ( .A(n9842), .B(n9841), .X(n3945) );
  nand_x1_sg U9140 ( .A(n9840), .B(n9839), .X(n3946) );
  nand_x1_sg U9141 ( .A(n9838), .B(n9837), .X(n3947) );
  nand_x1_sg U9142 ( .A(n9836), .B(n9835), .X(n3948) );
  nand_x1_sg U9143 ( .A(n9834), .B(n9833), .X(n3949) );
  nand_x1_sg U9144 ( .A(n9832), .B(n9831), .X(n3950) );
  nand_x1_sg U9145 ( .A(n9830), .B(n9829), .X(n3951) );
  nand_x1_sg U9146 ( .A(n9828), .B(n9827), .X(n3952) );
  nand_x1_sg U9147 ( .A(n9826), .B(n9825), .X(n3953) );
  nand_x1_sg U9148 ( .A(n9824), .B(n9823), .X(n3954) );
  nand_x1_sg U9149 ( .A(n9822), .B(n9821), .X(n3955) );
  nand_x1_sg U9150 ( .A(n9820), .B(n9819), .X(n3956) );
  nand_x1_sg U9151 ( .A(n9818), .B(n9817), .X(n3957) );
  nand_x1_sg U9152 ( .A(n9816), .B(n9815), .X(n3958) );
  nand_x1_sg U9153 ( .A(n9814), .B(n9813), .X(n3959) );
  nand_x1_sg U9154 ( .A(n9812), .B(n9811), .X(n3960) );
  nand_x1_sg U9155 ( .A(n9810), .B(n9809), .X(n3961) );
  nand_x1_sg U9156 ( .A(n9808), .B(n9807), .X(n3962) );
  nand_x1_sg U9157 ( .A(n9806), .B(n9805), .X(n3963) );
  nand_x1_sg U9158 ( .A(n9804), .B(n9803), .X(n3964) );
  nand_x1_sg U9159 ( .A(n9802), .B(n9801), .X(n3965) );
  nand_x1_sg U9160 ( .A(n9800), .B(n9799), .X(n3966) );
  nand_x1_sg U9161 ( .A(n9798), .B(n9797), .X(n3967) );
  nand_x1_sg U9162 ( .A(n9796), .B(n9795), .X(n3968) );
  nand_x1_sg U9163 ( .A(n9794), .B(n9793), .X(n3969) );
  nand_x1_sg U9164 ( .A(n9792), .B(n9791), .X(n3970) );
  nand_x1_sg U9165 ( .A(n9790), .B(n9789), .X(n3971) );
  nand_x1_sg U9166 ( .A(n9788), .B(n9787), .X(n3972) );
  nand_x1_sg U9167 ( .A(n9786), .B(n9785), .X(n3973) );
  nand_x1_sg U9168 ( .A(n9784), .B(n9783), .X(n3974) );
  nand_x1_sg U9169 ( .A(n9782), .B(n9781), .X(n3975) );
  nand_x1_sg U9170 ( .A(n9780), .B(n9779), .X(n3976) );
  nand_x1_sg U9171 ( .A(n9778), .B(n9777), .X(n3977) );
  nand_x1_sg U9172 ( .A(n9776), .B(n9775), .X(n3978) );
  nand_x1_sg U9173 ( .A(n9774), .B(n9773), .X(n3979) );
  nand_x1_sg U9174 ( .A(n9772), .B(n9771), .X(n3980) );
  nand_x1_sg U9175 ( .A(n9770), .B(n9769), .X(n3981) );
  nand_x1_sg U9176 ( .A(n9768), .B(n9767), .X(n3982) );
  nand_x1_sg U9177 ( .A(n9766), .B(n9765), .X(n3983) );
  nand_x1_sg U9178 ( .A(n9764), .B(n9763), .X(n3984) );
  nand_x1_sg U9179 ( .A(n9762), .B(n9761), .X(n3985) );
  nand_x1_sg U9180 ( .A(n9759), .B(n9760), .X(n3986) );
  nand_x1_sg U9181 ( .A(n9758), .B(n9757), .X(n3987) );
  nand_x1_sg U9182 ( .A(n9756), .B(n9755), .X(n3988) );
  nand_x1_sg U9183 ( .A(n9754), .B(n9753), .X(n3989) );
  nand_x1_sg U9184 ( .A(n9752), .B(n9751), .X(n3990) );
  nand_x1_sg U9185 ( .A(n9750), .B(n9749), .X(n3991) );
  nand_x1_sg U9186 ( .A(n9748), .B(n9747), .X(n3992) );
  nand_x1_sg U9187 ( .A(n9746), .B(n9745), .X(n3993) );
  nand_x1_sg U9188 ( .A(n9744), .B(n9743), .X(n3994) );
  nand_x1_sg U9189 ( .A(n9742), .B(n9741), .X(n3995) );
  nand_x1_sg U9190 ( .A(n9740), .B(n9739), .X(n3996) );
  nand_x1_sg U9191 ( .A(n9738), .B(n9737), .X(n3997) );
  nand_x1_sg U9192 ( .A(n9736), .B(n9735), .X(n3998) );
  nand_x1_sg U9193 ( .A(n9734), .B(n9733), .X(n3999) );
  nand_x1_sg U9194 ( .A(n9732), .B(n9731), .X(n4000) );
  nand_x1_sg U9195 ( .A(n9730), .B(n9729), .X(n4001) );
  nand_x1_sg U9196 ( .A(n9728), .B(n9727), .X(n4002) );
  nand_x1_sg U9197 ( .A(n9726), .B(n9725), .X(n4003) );
  nand_x1_sg U9198 ( .A(n9724), .B(n9723), .X(n4004) );
  nand_x1_sg U9199 ( .A(n9722), .B(n9721), .X(n4005) );
  nand_x1_sg U9200 ( .A(n9720), .B(n9719), .X(n4006) );
  nand_x1_sg U9201 ( .A(n9718), .B(n9717), .X(n4007) );
  nand_x1_sg U9202 ( .A(n9716), .B(n9715), .X(n4008) );
  nand_x1_sg U9203 ( .A(n9714), .B(n9713), .X(n4009) );
  nand_x1_sg U9204 ( .A(n9712), .B(n9711), .X(n4010) );
  nand_x1_sg U9205 ( .A(n9710), .B(n9709), .X(n4011) );
  nand_x1_sg U9206 ( .A(n9708), .B(n9707), .X(n4012) );
  nand_x1_sg U9207 ( .A(n9706), .B(n9705), .X(n4013) );
  nand_x1_sg U9208 ( .A(n9704), .B(n9703), .X(n4014) );
  nand_x1_sg U9209 ( .A(n9702), .B(n9701), .X(n4015) );
  nand_x1_sg U9210 ( .A(n9700), .B(n9699), .X(n4016) );
  nand_x1_sg U9211 ( .A(n9698), .B(n9697), .X(n4017) );
  nand_x1_sg U9212 ( .A(n9696), .B(n9695), .X(n4018) );
  nand_x1_sg U9213 ( .A(n9694), .B(n9693), .X(n4019) );
  nand_x1_sg U9214 ( .A(n9692), .B(n9691), .X(n4020) );
  nand_x1_sg U9215 ( .A(n9690), .B(n9689), .X(n4021) );
  nand_x1_sg U9216 ( .A(n9688), .B(n9687), .X(n4022) );
  nand_x1_sg U9217 ( .A(n9686), .B(n9685), .X(n4023) );
  nand_x1_sg U9218 ( .A(n9684), .B(n9683), .X(n4024) );
  nand_x1_sg U9219 ( .A(n9682), .B(n9681), .X(n4025) );
  nand_x1_sg U9220 ( .A(n9680), .B(n9679), .X(n4026) );
  nand_x1_sg U9221 ( .A(n9678), .B(n9677), .X(n4027) );
  nand_x1_sg U9222 ( .A(n9676), .B(n9675), .X(n4028) );
  nand_x1_sg U9223 ( .A(n9674), .B(n9673), .X(n4029) );
  nand_x1_sg U9224 ( .A(n9672), .B(n9671), .X(n4030) );
  nand_x1_sg U9225 ( .A(n9670), .B(n9669), .X(n4031) );
  nand_x1_sg U9226 ( .A(n9668), .B(n9667), .X(n4032) );
  nand_x1_sg U9227 ( .A(n9666), .B(n9665), .X(n4033) );
  nand_x1_sg U9228 ( .A(n9664), .B(n9663), .X(n4034) );
  nand_x1_sg U9229 ( .A(n9662), .B(n9661), .X(n4035) );
  nand_x1_sg U9230 ( .A(n9660), .B(n9659), .X(n4036) );
  nand_x1_sg U9231 ( .A(n9658), .B(n9657), .X(n4037) );
  nand_x1_sg U9232 ( .A(n9656), .B(n9655), .X(n4038) );
  nand_x1_sg U9233 ( .A(n9654), .B(n9653), .X(n4039) );
  nand_x1_sg U9234 ( .A(n9652), .B(n9651), .X(n4040) );
  nand_x1_sg U9235 ( .A(n9650), .B(n9649), .X(n4041) );
  nand_x1_sg U9236 ( .A(n9648), .B(n9647), .X(n4042) );
  nand_x1_sg U9237 ( .A(n9646), .B(n9645), .X(n4043) );
  nand_x1_sg U9238 ( .A(n9644), .B(n9643), .X(n4044) );
  nand_x1_sg U9239 ( .A(n9642), .B(n9641), .X(n4045) );
  nand_x1_sg U9240 ( .A(n9640), .B(n9639), .X(n4046) );
  nand_x1_sg U9241 ( .A(n9638), .B(n9637), .X(n4047) );
  nand_x1_sg U9242 ( .A(n9636), .B(n9635), .X(n4048) );
  nand_x1_sg U9243 ( .A(n9634), .B(n9633), .X(n4049) );
  nand_x1_sg U9244 ( .A(n9632), .B(n9631), .X(n4050) );
  nand_x1_sg U9245 ( .A(n9630), .B(n9629), .X(n4051) );
  nand_x1_sg U9246 ( .A(n9628), .B(n9627), .X(n4052) );
  nand_x1_sg U9247 ( .A(n9626), .B(n9625), .X(n4053) );
  nand_x1_sg U9248 ( .A(n9624), .B(n9623), .X(n4054) );
  nand_x1_sg U9249 ( .A(n9622), .B(n9621), .X(n4055) );
  nand_x1_sg U9250 ( .A(n9620), .B(n9619), .X(n4056) );
  nand_x1_sg U9251 ( .A(n9618), .B(n9617), .X(n4057) );
  nand_x1_sg U9252 ( .A(n9616), .B(n9615), .X(n4058) );
  nand_x1_sg U9253 ( .A(n9614), .B(n9613), .X(n4059) );
  nand_x1_sg U9254 ( .A(n9612), .B(n9611), .X(n4060) );
  nand_x1_sg U9255 ( .A(n9610), .B(n9609), .X(n4061) );
  nand_x1_sg U9256 ( .A(n9608), .B(n9607), .X(n4062) );
  nand_x1_sg U9257 ( .A(n9606), .B(n9605), .X(n4063) );
  nand_x1_sg U9258 ( .A(n9604), .B(n9603), .X(n4064) );
  nand_x1_sg U9259 ( .A(n9602), .B(n9601), .X(n4065) );
  nand_x1_sg U9260 ( .A(n9600), .B(n9599), .X(n4066) );
  nand_x1_sg U9261 ( .A(n9598), .B(n9597), .X(n4067) );
  nand_x1_sg U9262 ( .A(n9596), .B(n9595), .X(n4068) );
  nand_x1_sg U9263 ( .A(n9594), .B(n9593), .X(n4069) );
  nand_x1_sg U9264 ( .A(n9592), .B(n9591), .X(n4070) );
  nand_x1_sg U9265 ( .A(n9590), .B(n9589), .X(n4071) );
  nand_x1_sg U9266 ( .A(n9588), .B(n9587), .X(n4072) );
  nand_x1_sg U9267 ( .A(n9586), .B(n9585), .X(n4073) );
  nand_x1_sg U9268 ( .A(n9584), .B(n9583), .X(n4074) );
  nand_x1_sg U9269 ( .A(n9582), .B(n9581), .X(n4075) );
  nand_x1_sg U9270 ( .A(n9580), .B(n9579), .X(n4076) );
  nand_x1_sg U9271 ( .A(n9578), .B(n9577), .X(n4077) );
  nand_x1_sg U9272 ( .A(n9576), .B(n9575), .X(n4078) );
  nand_x1_sg U9273 ( .A(n9574), .B(n9573), .X(n4079) );
  nand_x1_sg U9274 ( .A(n9572), .B(n9571), .X(n4080) );
  nand_x1_sg U9275 ( .A(n9570), .B(n9569), .X(n4081) );
  nand_x1_sg U9276 ( .A(n9568), .B(n9567), .X(n4082) );
  nand_x1_sg U9277 ( .A(n9566), .B(n9565), .X(n4083) );
  nand_x1_sg U9278 ( .A(n9564), .B(n9563), .X(n4084) );
  nand_x1_sg U9279 ( .A(n9562), .B(n9561), .X(n4085) );
  nand_x1_sg U9280 ( .A(n9560), .B(n9559), .X(n4086) );
  nand_x1_sg U9281 ( .A(n9558), .B(n9557), .X(n4087) );
  nand_x1_sg U9282 ( .A(n9556), .B(n9555), .X(n4088) );
  nand_x1_sg U9283 ( .A(n9554), .B(n9553), .X(n4089) );
  nand_x1_sg U9284 ( .A(n9552), .B(n9551), .X(n4090) );
  nand_x1_sg U9285 ( .A(n9550), .B(n9549), .X(n4091) );
  nand_x1_sg U9286 ( .A(n9548), .B(n9547), .X(n4092) );
  nand_x1_sg U9287 ( .A(n9546), .B(n9545), .X(n4093) );
  nand_x1_sg U9288 ( .A(n9544), .B(n9543), .X(n4094) );
  nand_x1_sg U9289 ( .A(n9542), .B(n9541), .X(n4095) );
  nand_x1_sg U9290 ( .A(n9540), .B(n9539), .X(n4096) );
  nand_x1_sg U9291 ( .A(n9538), .B(n9537), .X(n4097) );
  nand_x1_sg U9292 ( .A(n9536), .B(n9535), .X(n4098) );
  nand_x1_sg U9293 ( .A(n9534), .B(n9533), .X(n4099) );
  nand_x1_sg U9294 ( .A(n9532), .B(n9531), .X(n4100) );
  nand_x1_sg U9295 ( .A(n9530), .B(n9529), .X(n4101) );
  nand_x1_sg U9296 ( .A(n9528), .B(n9527), .X(n4102) );
  nand_x1_sg U9297 ( .A(n9526), .B(n9525), .X(n4103) );
  nand_x1_sg U9298 ( .A(n9524), .B(n9523), .X(n4104) );
  nand_x1_sg U9299 ( .A(n9522), .B(n9521), .X(n4105) );
  nand_x1_sg U9300 ( .A(n9520), .B(n9519), .X(n4106) );
  nand_x1_sg U9301 ( .A(n9518), .B(n9517), .X(n4107) );
  nand_x1_sg U9302 ( .A(n9516), .B(n9515), .X(n4108) );
  nand_x1_sg U9303 ( .A(n9514), .B(n9513), .X(n4109) );
  nand_x1_sg U9304 ( .A(n9511), .B(n9512), .X(n4110) );
  nand_x1_sg U9305 ( .A(n9510), .B(n9509), .X(n4111) );
  nand_x1_sg U9306 ( .A(n9508), .B(n9507), .X(n4112) );
  nand_x1_sg U9307 ( .A(n9506), .B(n9505), .X(n4113) );
  nand_x1_sg U9308 ( .A(n9504), .B(n9503), .X(n4114) );
  nand_x1_sg U9309 ( .A(n9502), .B(n9501), .X(n4115) );
  nand_x1_sg U9310 ( .A(n9500), .B(n9499), .X(n4116) );
  nand_x1_sg U9311 ( .A(n9498), .B(n9497), .X(n4117) );
  nand_x1_sg U9312 ( .A(n9496), .B(n9495), .X(n4118) );
  nand_x1_sg U9313 ( .A(n9494), .B(n9493), .X(n4119) );
  nand_x1_sg U9314 ( .A(n9492), .B(n9491), .X(n4120) );
  nand_x1_sg U9315 ( .A(n9490), .B(n9489), .X(n4121) );
  nand_x1_sg U9316 ( .A(n9488), .B(n9487), .X(n4122) );
  nand_x1_sg U9317 ( .A(n9486), .B(n9485), .X(n4123) );
  nand_x1_sg U9318 ( .A(n9484), .B(n9483), .X(n4124) );
  nand_x1_sg U9319 ( .A(n9482), .B(n9481), .X(n4125) );
  nand_x1_sg U9320 ( .A(n9480), .B(n9479), .X(n4126) );
  nand_x1_sg U9321 ( .A(n9478), .B(n9477), .X(n4127) );
  nand_x1_sg U9322 ( .A(n9476), .B(n9475), .X(n4128) );
  nand_x1_sg U9323 ( .A(n9474), .B(n9473), .X(n4129) );
  nand_x1_sg U9324 ( .A(n9472), .B(n9471), .X(n4130) );
  nand_x1_sg U9325 ( .A(n9470), .B(n9469), .X(n4131) );
  nand_x1_sg U9326 ( .A(n9468), .B(n9467), .X(n4132) );
  nand_x1_sg U9327 ( .A(n9466), .B(n9465), .X(n4133) );
  nand_x1_sg U9328 ( .A(n9464), .B(n9463), .X(n4134) );
  nand_x1_sg U9329 ( .A(n9462), .B(n9461), .X(n4135) );
  nand_x1_sg U9330 ( .A(n9460), .B(n9459), .X(n4136) );
  nand_x1_sg U9331 ( .A(n9458), .B(n9457), .X(n4137) );
  nand_x1_sg U9332 ( .A(n9456), .B(n9455), .X(n4138) );
  nand_x1_sg U9333 ( .A(n9454), .B(n9453), .X(n4139) );
  nand_x1_sg U9334 ( .A(n9452), .B(n9451), .X(n4140) );
  nand_x1_sg U9335 ( .A(n9450), .B(n9449), .X(n4141) );
  nand_x1_sg U9336 ( .A(n9448), .B(n9447), .X(n4142) );
  nand_x1_sg U9337 ( .A(n9446), .B(n9445), .X(n4143) );
  nand_x1_sg U9338 ( .A(n9444), .B(n9443), .X(n4144) );
  nand_x1_sg U9339 ( .A(n9442), .B(n9441), .X(n4145) );
  nand_x1_sg U9340 ( .A(n9440), .B(n9439), .X(n4146) );
  nand_x1_sg U9341 ( .A(n9438), .B(n9437), .X(n4147) );
  nand_x1_sg U9342 ( .A(n9436), .B(n9435), .X(n4148) );
  nand_x1_sg U9343 ( .A(n9434), .B(n9433), .X(n4149) );
  nand_x1_sg U9344 ( .A(n9432), .B(n9431), .X(n4150) );
  nand_x1_sg U9345 ( .A(n9430), .B(n9429), .X(n4151) );
  nand_x1_sg U9346 ( .A(n9428), .B(n9427), .X(n4152) );
  nand_x1_sg U9347 ( .A(n9426), .B(n9425), .X(n4153) );
  nand_x1_sg U9348 ( .A(n9424), .B(n9423), .X(n4154) );
  nand_x1_sg U9349 ( .A(n9422), .B(n9421), .X(n4155) );
  nand_x1_sg U9350 ( .A(n9420), .B(n9419), .X(n4156) );
  nand_x1_sg U9351 ( .A(n9418), .B(n9417), .X(n4157) );
  nand_x1_sg U9352 ( .A(n9416), .B(n9415), .X(n4158) );
  nand_x1_sg U9353 ( .A(n9414), .B(n9413), .X(n4159) );
  nand_x1_sg U9354 ( .A(n9412), .B(n9411), .X(n4160) );
  nand_x1_sg U9355 ( .A(n9410), .B(n9409), .X(n4161) );
  nand_x1_sg U9356 ( .A(n9408), .B(n9407), .X(n4162) );
  nand_x1_sg U9357 ( .A(n9406), .B(n9405), .X(n4163) );
  nand_x1_sg U9358 ( .A(n9404), .B(n9403), .X(n4164) );
  nand_x1_sg U9359 ( .A(n9402), .B(n9401), .X(n4165) );
  nand_x1_sg U9360 ( .A(n9400), .B(n9399), .X(n4166) );
  nand_x1_sg U9361 ( .A(n9398), .B(n9397), .X(n4167) );
  nand_x1_sg U9362 ( .A(n9396), .B(n9395), .X(n4168) );
  nand_x1_sg U9363 ( .A(n9394), .B(n9393), .X(n4169) );
  nand_x1_sg U9364 ( .A(n9392), .B(n9391), .X(n4170) );
  nand_x1_sg U9365 ( .A(n9390), .B(n9389), .X(n4171) );
  nand_x1_sg U9366 ( .A(n9388), .B(n9387), .X(n4172) );
  nand_x1_sg U9367 ( .A(n9386), .B(n9385), .X(n4173) );
  nand_x1_sg U9368 ( .A(n9384), .B(n9383), .X(n4174) );
  nand_x1_sg U9369 ( .A(n9382), .B(n9381), .X(n4175) );
  nand_x1_sg U9370 ( .A(n9379), .B(n9380), .X(n4176) );
  nand_x1_sg U9371 ( .A(n9378), .B(n9377), .X(n4177) );
  nand_x1_sg U9372 ( .A(n9376), .B(n9375), .X(n4178) );
  nand_x1_sg U9373 ( .A(n9374), .B(n9373), .X(n4179) );
  nand_x1_sg U9374 ( .A(n9372), .B(n9371), .X(n4180) );
  nand_x1_sg U9375 ( .A(n9370), .B(n9369), .X(n4181) );
  nand_x1_sg U9376 ( .A(n9368), .B(n9367), .X(n4182) );
  nand_x1_sg U9377 ( .A(n9366), .B(n9365), .X(n4183) );
  nand_x1_sg U9378 ( .A(n9364), .B(n9363), .X(n4184) );
  nand_x1_sg U9379 ( .A(n9361), .B(n9360), .X(n4185) );
  nand_x1_sg U9380 ( .A(n9357), .B(n9358), .X(n4186) );
  nand_x1_sg U9381 ( .A(n9355), .B(n9356), .X(n4187) );
  nand_x1_sg U9382 ( .A(n9353), .B(n9354), .X(n4188) );
  nand_x1_sg U9383 ( .A(n9351), .B(n9352), .X(n4189) );
  nand_x1_sg U9384 ( .A(n9349), .B(n9350), .X(n4190) );
  nand_x1_sg U9385 ( .A(n9347), .B(n9348), .X(n4191) );
  nand_x1_sg U9386 ( .A(n9345), .B(n9346), .X(n4192) );
  nand_x1_sg U9387 ( .A(n9343), .B(n9344), .X(n4193) );
  nand_x1_sg U9388 ( .A(n9341), .B(n9342), .X(n4194) );
  nand_x1_sg U9389 ( .A(n9339), .B(n9340), .X(n4195) );
  nand_x1_sg U9390 ( .A(n9337), .B(n9338), .X(n4196) );
  nand_x1_sg U9391 ( .A(n9335), .B(n9336), .X(n4197) );
  nand_x1_sg U9392 ( .A(n9333), .B(n9334), .X(n4198) );
  nand_x1_sg U9393 ( .A(n9331), .B(n9332), .X(n4199) );
  nand_x1_sg U9394 ( .A(n9329), .B(n9330), .X(n4200) );
  nand_x1_sg U9395 ( .A(n9327), .B(n9328), .X(n4201) );
  nand_x1_sg U9396 ( .A(n9325), .B(n9326), .X(n4202) );
  nand_x1_sg U9397 ( .A(n9323), .B(n9324), .X(n4203) );
  nand_x1_sg U9398 ( .A(n9321), .B(n9322), .X(n4204) );
  nand_x1_sg U9399 ( .A(n9319), .B(n9320), .X(n4205) );
  nand_x1_sg U9400 ( .A(n9317), .B(n9318), .X(n4206) );
  nand_x1_sg U9401 ( .A(n9315), .B(n9316), .X(n4207) );
  nand_x1_sg U9402 ( .A(n9313), .B(n9314), .X(n4208) );
  nand_x1_sg U9403 ( .A(n9311), .B(n9312), .X(n4209) );
  nand_x1_sg U9404 ( .A(n9309), .B(n9310), .X(n4210) );
  nand_x1_sg U9405 ( .A(n9307), .B(n9308), .X(n4211) );
  nand_x1_sg U9406 ( .A(n9305), .B(n9306), .X(n4212) );
  nand_x1_sg U9407 ( .A(n9303), .B(n9304), .X(n4213) );
  nand_x1_sg U9408 ( .A(n9301), .B(n9302), .X(n4214) );
  nand_x1_sg U9409 ( .A(n9299), .B(n9300), .X(n4215) );
  nand_x1_sg U9410 ( .A(n9297), .B(n9298), .X(n4216) );
  nand_x1_sg U9411 ( .A(n9295), .B(n9296), .X(n4217) );
  nand_x1_sg U9412 ( .A(n9293), .B(n9294), .X(n4218) );
  nand_x1_sg U9413 ( .A(n9291), .B(n9292), .X(n4219) );
  nand_x1_sg U9414 ( .A(n9289), .B(n9290), .X(n4220) );
  nand_x1_sg U9415 ( .A(n9287), .B(n9288), .X(n4221) );
  nand_x1_sg U9416 ( .A(n9285), .B(n9286), .X(n4222) );
  nand_x1_sg U9417 ( .A(n9283), .B(n9284), .X(n4223) );
  nand_x1_sg U9418 ( .A(n9281), .B(n9282), .X(n4224) );
  nand_x1_sg U9419 ( .A(n9279), .B(n9280), .X(n4225) );
  nand_x1_sg U9420 ( .A(n9277), .B(n9278), .X(n4226) );
  nand_x1_sg U9421 ( .A(n9275), .B(n9276), .X(n4227) );
  nand_x1_sg U9422 ( .A(n9273), .B(n9274), .X(n4228) );
  nand_x1_sg U9423 ( .A(n9271), .B(n9272), .X(n4229) );
  nand_x1_sg U9424 ( .A(n9269), .B(n9270), .X(n4230) );
  nand_x1_sg U9425 ( .A(n9267), .B(n9268), .X(n4231) );
  nand_x1_sg U9426 ( .A(n9265), .B(n9266), .X(n4232) );
  nand_x1_sg U9427 ( .A(n9263), .B(n9264), .X(n4233) );
  nand_x1_sg U9428 ( .A(n9261), .B(n9262), .X(n4234) );
  nand_x1_sg U9429 ( .A(n9259), .B(n9260), .X(n4235) );
  nand_x1_sg U9430 ( .A(n9257), .B(n9258), .X(n4236) );
  nand_x1_sg U9431 ( .A(n9255), .B(n9256), .X(n4237) );
  nand_x1_sg U9432 ( .A(n9253), .B(n9254), .X(n4238) );
  nand_x1_sg U9433 ( .A(n9251), .B(n9252), .X(n4239) );
  nand_x1_sg U9434 ( .A(n9249), .B(n9250), .X(n4240) );
  nand_x1_sg U9435 ( .A(n9247), .B(n9248), .X(n4241) );
  nand_x1_sg U9436 ( .A(n9245), .B(n9246), .X(n4242) );
  nand_x1_sg U9437 ( .A(n9243), .B(n9244), .X(n4243) );
  nand_x1_sg U9438 ( .A(n9241), .B(n9242), .X(n4244) );
  nand_x1_sg U9439 ( .A(n9239), .B(n9240), .X(n4245) );
  nand_x1_sg U9440 ( .A(n9237), .B(n9238), .X(n4246) );
  nand_x1_sg U9441 ( .A(n9235), .B(n9236), .X(n4247) );
  nand_x1_sg U9442 ( .A(n9233), .B(n9234), .X(n4248) );
  nand_x1_sg U9443 ( .A(n9231), .B(n9232), .X(n4249) );
  nand_x1_sg U9444 ( .A(n9229), .B(n9230), .X(n4250) );
  nand_x1_sg U9445 ( .A(n9227), .B(n9228), .X(n4251) );
  nand_x1_sg U9446 ( .A(n9225), .B(n9226), .X(n4252) );
  nand_x1_sg U9447 ( .A(n9223), .B(n9224), .X(n4253) );
  nand_x1_sg U9448 ( .A(n9221), .B(n9222), .X(n4254) );
  nand_x1_sg U9449 ( .A(n9219), .B(n9220), .X(n4255) );
  nand_x1_sg U9450 ( .A(n9217), .B(n9218), .X(n4256) );
  nand_x1_sg U9451 ( .A(n9215), .B(n9216), .X(n4257) );
  nand_x1_sg U9452 ( .A(n9213), .B(n9214), .X(n4258) );
  nand_x1_sg U9453 ( .A(n9211), .B(n9212), .X(n4259) );
  nand_x1_sg U9454 ( .A(n9209), .B(n9210), .X(n4260) );
  nand_x1_sg U9455 ( .A(n9207), .B(n9208), .X(n4261) );
  nand_x1_sg U9456 ( .A(n9205), .B(n9206), .X(n4262) );
  nand_x1_sg U9457 ( .A(n9203), .B(n9204), .X(n4263) );
  nand_x1_sg U9458 ( .A(n9201), .B(n9202), .X(n4264) );
  nand_x1_sg U9459 ( .A(n9199), .B(n9200), .X(n4265) );
  nand_x1_sg U9460 ( .A(n9197), .B(n9198), .X(n4266) );
  nand_x1_sg U9461 ( .A(n9195), .B(n9196), .X(n4267) );
  nand_x1_sg U9462 ( .A(n9193), .B(n9194), .X(n4268) );
  nand_x1_sg U9463 ( .A(n9191), .B(n9192), .X(n4269) );
  nand_x1_sg U9464 ( .A(n9189), .B(n9190), .X(n4270) );
  nand_x1_sg U9465 ( .A(n9187), .B(n9188), .X(n4271) );
  nand_x1_sg U9466 ( .A(n9185), .B(n9186), .X(n4272) );
  nand_x1_sg U9467 ( .A(n9183), .B(n9184), .X(n4273) );
  nand_x1_sg U9468 ( .A(n9181), .B(n9182), .X(n4274) );
  nand_x1_sg U9469 ( .A(n9179), .B(n9180), .X(n4275) );
  nand_x1_sg U9470 ( .A(n9177), .B(n9178), .X(n4276) );
  nand_x1_sg U9471 ( .A(n9175), .B(n9176), .X(n4277) );
  nand_x1_sg U9472 ( .A(n9173), .B(n9174), .X(n4278) );
  nand_x1_sg U9473 ( .A(n9171), .B(n9172), .X(n4279) );
  nand_x1_sg U9474 ( .A(n9169), .B(n9170), .X(n4280) );
  nand_x1_sg U9475 ( .A(n9167), .B(n9168), .X(n4281) );
  nand_x1_sg U9476 ( .A(n9165), .B(n9166), .X(n4282) );
  nand_x1_sg U9477 ( .A(n9163), .B(n9164), .X(n4283) );
  nand_x1_sg U9478 ( .A(n9161), .B(n9162), .X(n4284) );
  nand_x1_sg U9479 ( .A(n9159), .B(n9160), .X(n4285) );
  nand_x1_sg U9480 ( .A(n9157), .B(n9158), .X(n4286) );
  nand_x1_sg U9481 ( .A(n9155), .B(n9156), .X(n4287) );
  nand_x1_sg U9482 ( .A(n9153), .B(n9154), .X(n4288) );
  nand_x1_sg U9483 ( .A(n9151), .B(n9152), .X(n4289) );
  nand_x1_sg U9484 ( .A(n9149), .B(n9150), .X(n4290) );
  nand_x1_sg U9485 ( .A(n9147), .B(n9148), .X(n4291) );
  nand_x1_sg U9486 ( .A(n9145), .B(n9146), .X(n4292) );
  nand_x1_sg U9487 ( .A(n9143), .B(n9144), .X(n4293) );
  nand_x1_sg U9488 ( .A(n9141), .B(n9142), .X(n4294) );
  nand_x1_sg U9489 ( .A(n9139), .B(n9140), .X(n4295) );
  nand_x1_sg U9490 ( .A(n9137), .B(n9138), .X(n4296) );
  nand_x1_sg U9491 ( .A(n9135), .B(n9136), .X(n4297) );
  nand_x1_sg U9492 ( .A(n9133), .B(n9134), .X(n4298) );
  nand_x1_sg U9493 ( .A(n9131), .B(n9132), .X(n4299) );
  nand_x1_sg U9494 ( .A(n9129), .B(n9130), .X(n4300) );
  nand_x1_sg U9495 ( .A(n9127), .B(n9128), .X(n4301) );
  nand_x1_sg U9496 ( .A(n9125), .B(n9126), .X(n4302) );
  nand_x1_sg U9497 ( .A(n9123), .B(n9124), .X(n4303) );
  nand_x1_sg U9498 ( .A(n9121), .B(n9122), .X(n4304) );
  nand_x1_sg U9499 ( .A(n9119), .B(n9120), .X(n4305) );
  nand_x1_sg U9500 ( .A(n9117), .B(n9118), .X(n4306) );
  nand_x1_sg U9501 ( .A(n9115), .B(n9116), .X(n4307) );
  nand_x1_sg U9502 ( .A(n9113), .B(n9114), .X(n4308) );
  nand_x1_sg U9503 ( .A(n9111), .B(n9112), .X(n4309) );
  nand_x1_sg U9504 ( .A(n9109), .B(n9110), .X(n4310) );
  nand_x1_sg U9505 ( .A(n9107), .B(n9108), .X(n4311) );
  nand_x1_sg U9506 ( .A(n9105), .B(n9106), .X(n4312) );
  nand_x1_sg U9507 ( .A(n9103), .B(n9104), .X(n4313) );
  nand_x1_sg U9508 ( .A(n9101), .B(n9102), .X(n4314) );
  nand_x1_sg U9509 ( .A(n9099), .B(n9100), .X(n4315) );
  nand_x1_sg U9510 ( .A(n9097), .B(n9098), .X(n4316) );
  nand_x1_sg U9511 ( .A(n9095), .B(n9096), .X(n4317) );
  nand_x1_sg U9512 ( .A(n9093), .B(n9094), .X(n4318) );
  nand_x1_sg U9513 ( .A(n9091), .B(n9092), .X(n4319) );
  nand_x1_sg U9514 ( .A(n9089), .B(n9090), .X(n4320) );
  nand_x1_sg U9515 ( .A(n9087), .B(n9088), .X(n4321) );
  nand_x1_sg U9516 ( .A(n9085), .B(n9086), .X(n4322) );
  nand_x1_sg U9517 ( .A(n9083), .B(n9084), .X(n4323) );
  nand_x1_sg U9518 ( .A(n9081), .B(n9082), .X(n4324) );
  nand_x1_sg U9519 ( .A(n9079), .B(n9080), .X(n4325) );
  nand_x1_sg U9520 ( .A(n9077), .B(n9078), .X(n4326) );
  nand_x1_sg U9521 ( .A(n9075), .B(n9076), .X(n4327) );
  nand_x1_sg U9522 ( .A(n9073), .B(n9074), .X(n4328) );
  nand_x1_sg U9523 ( .A(n9071), .B(n9072), .X(n4329) );
  nand_x1_sg U9524 ( .A(n9069), .B(n9070), .X(n4330) );
  nand_x1_sg U9525 ( .A(n9067), .B(n9068), .X(n4331) );
  nand_x1_sg U9526 ( .A(n9065), .B(n9066), .X(n4332) );
  nand_x1_sg U9527 ( .A(n9063), .B(n9064), .X(n4333) );
  nand_x1_sg U9528 ( .A(n9061), .B(n9062), .X(n4334) );
  nand_x1_sg U9529 ( .A(n9059), .B(n9060), .X(n4335) );
  nand_x1_sg U9530 ( .A(n9057), .B(n9058), .X(n4336) );
  nand_x1_sg U9531 ( .A(n9055), .B(n9056), .X(n4337) );
  nand_x1_sg U9532 ( .A(n9053), .B(n9054), .X(n4338) );
  nand_x1_sg U9533 ( .A(n9051), .B(n9052), .X(n4339) );
  nand_x1_sg U9534 ( .A(n9049), .B(n9050), .X(n4340) );
  nand_x1_sg U9535 ( .A(n9047), .B(n9048), .X(n4341) );
  nand_x1_sg U9536 ( .A(n9045), .B(n9046), .X(n4342) );
  nand_x1_sg U9537 ( .A(n9043), .B(n9044), .X(n4343) );
  nand_x1_sg U9538 ( .A(n9041), .B(n9042), .X(n4344) );
  nand_x1_sg U9539 ( .A(n9039), .B(n9040), .X(n4345) );
  nand_x1_sg U9540 ( .A(n9037), .B(n9038), .X(n4346) );
  nand_x1_sg U9541 ( .A(n9035), .B(n9036), .X(n4347) );
  nand_x1_sg U9542 ( .A(n9033), .B(n9034), .X(n4348) );
  nand_x1_sg U9543 ( .A(n9031), .B(n9032), .X(n4349) );
  nand_x1_sg U9544 ( .A(n9029), .B(n9030), .X(n4350) );
  nand_x1_sg U9545 ( .A(n9027), .B(n9028), .X(n4351) );
  nand_x1_sg U9546 ( .A(n9025), .B(n9026), .X(n4352) );
  nand_x1_sg U9547 ( .A(n9023), .B(n9024), .X(n4353) );
  nand_x1_sg U9548 ( .A(n9021), .B(n9022), .X(n4354) );
  nand_x1_sg U9549 ( .A(n9019), .B(n9020), .X(n4355) );
  nand_x1_sg U9550 ( .A(n9017), .B(n9018), .X(n4356) );
  nand_x1_sg U9551 ( .A(n9015), .B(n9016), .X(n4357) );
  nand_x1_sg U9552 ( .A(n9013), .B(n9014), .X(n4358) );
  nand_x1_sg U9553 ( .A(n9011), .B(n9012), .X(n4359) );
  nand_x1_sg U9554 ( .A(n9009), .B(n9010), .X(n4360) );
  nand_x1_sg U9555 ( .A(n9007), .B(n9008), .X(n4361) );
  nand_x1_sg U9556 ( .A(n9005), .B(n9006), .X(n4362) );
  nand_x1_sg U9557 ( .A(n9003), .B(n9004), .X(n4363) );
  nand_x1_sg U9558 ( .A(n9001), .B(n9002), .X(n4364) );
  nand_x1_sg U9559 ( .A(n8999), .B(n9000), .X(n4365) );
  nand_x1_sg U9560 ( .A(n8997), .B(n8998), .X(n4366) );
  nand_x1_sg U9561 ( .A(n8995), .B(n8996), .X(n4367) );
  nand_x1_sg U9562 ( .A(n8993), .B(n8994), .X(n4368) );
  nand_x1_sg U9563 ( .A(n8991), .B(n8992), .X(n4369) );
  nand_x1_sg U9564 ( .A(n8989), .B(n8990), .X(n4370) );
  nand_x1_sg U9565 ( .A(n8987), .B(n8988), .X(n4371) );
  nand_x1_sg U9566 ( .A(n8985), .B(n8986), .X(n4372) );
  nand_x1_sg U9567 ( .A(n8983), .B(n8984), .X(n4373) );
  nand_x1_sg U9568 ( .A(n8981), .B(n8982), .X(n4374) );
  nand_x1_sg U9569 ( .A(n8979), .B(n8980), .X(n4375) );
  nand_x1_sg U9570 ( .A(n8977), .B(n8978), .X(n4376) );
  nand_x1_sg U9571 ( .A(n8975), .B(n8976), .X(n4377) );
  nand_x1_sg U9572 ( .A(n8973), .B(n8974), .X(n4378) );
  nand_x1_sg U9573 ( .A(n8971), .B(n8972), .X(n4379) );
  nand_x1_sg U9574 ( .A(n8969), .B(n8970), .X(n4380) );
  nand_x1_sg U9575 ( .A(n8967), .B(n8968), .X(n4381) );
  nand_x1_sg U9576 ( .A(n8965), .B(n8966), .X(n4382) );
  nand_x1_sg U9577 ( .A(n8963), .B(n8964), .X(n4383) );
  nand_x1_sg U9578 ( .A(n8961), .B(n8962), .X(n4384) );
  nand_x1_sg U9579 ( .A(n8959), .B(n8960), .X(n4385) );
  nand_x1_sg U9580 ( .A(n8957), .B(n8958), .X(n4386) );
  nand_x1_sg U9581 ( .A(n8955), .B(n8956), .X(n4387) );
  nand_x1_sg U9582 ( .A(n8953), .B(n8954), .X(n4388) );
  nand_x1_sg U9583 ( .A(n8951), .B(n8952), .X(n4389) );
  nand_x1_sg U9584 ( .A(n8949), .B(n8950), .X(n4390) );
  nand_x1_sg U9585 ( .A(n8947), .B(n8948), .X(n4391) );
  nand_x1_sg U9586 ( .A(n8945), .B(n8946), .X(n4392) );
  nand_x1_sg U9587 ( .A(n8943), .B(n8944), .X(n4393) );
  nand_x1_sg U9588 ( .A(n8941), .B(n8942), .X(n4394) );
  nand_x1_sg U9589 ( .A(n8939), .B(n8940), .X(n4395) );
  nand_x1_sg U9590 ( .A(n8937), .B(n8938), .X(n4396) );
  nand_x1_sg U9591 ( .A(n8935), .B(n8936), .X(n4397) );
  nand_x1_sg U9592 ( .A(n8933), .B(n8934), .X(n4398) );
  nand_x1_sg U9593 ( .A(n8931), .B(n8932), .X(n4399) );
  nand_x1_sg U9594 ( .A(n8929), .B(n8930), .X(n4400) );
  nand_x1_sg U9595 ( .A(n8927), .B(n8928), .X(n4401) );
  nand_x1_sg U9596 ( .A(n8925), .B(n8926), .X(n4402) );
  nand_x1_sg U9597 ( .A(n8923), .B(n8924), .X(n4403) );
  nand_x1_sg U9598 ( .A(n8921), .B(n8922), .X(n4404) );
  nand_x1_sg U9599 ( .A(n8919), .B(n8920), .X(n4405) );
  nand_x1_sg U9600 ( .A(n8917), .B(n8918), .X(n4406) );
  nand_x1_sg U9601 ( .A(n8915), .B(n8916), .X(n4407) );
  nand_x1_sg U9602 ( .A(n8913), .B(n8914), .X(n4408) );
  nand_x1_sg U9603 ( .A(n8911), .B(n8912), .X(n4409) );
  nand_x1_sg U9604 ( .A(n8909), .B(n8910), .X(n4410) );
  nand_x1_sg U9605 ( .A(n8907), .B(n8908), .X(n4411) );
  nand_x1_sg U9606 ( .A(n8905), .B(n8906), .X(n4412) );
  nand_x1_sg U9607 ( .A(n8903), .B(n8904), .X(n4413) );
  nand_x1_sg U9608 ( .A(n8901), .B(n8902), .X(n4414) );
  nand_x1_sg U9609 ( .A(n8899), .B(n8900), .X(n4415) );
  nand_x1_sg U9610 ( .A(n8897), .B(n8898), .X(n4416) );
  nand_x1_sg U9611 ( .A(n8895), .B(n8896), .X(n4417) );
  nand_x1_sg U9612 ( .A(n8893), .B(n8894), .X(n4418) );
  nand_x1_sg U9613 ( .A(n8891), .B(n8892), .X(n4419) );
  nand_x1_sg U9614 ( .A(n8889), .B(n8890), .X(n4420) );
  nand_x1_sg U9615 ( .A(n8887), .B(n8888), .X(n4421) );
  nand_x1_sg U9616 ( .A(n8885), .B(n8886), .X(n4422) );
  nand_x1_sg U9617 ( .A(n8883), .B(n8884), .X(n4423) );
  nand_x1_sg U9618 ( .A(n8881), .B(n8882), .X(n4424) );
  nand_x1_sg U9619 ( .A(n8879), .B(n8880), .X(n4425) );
  nand_x1_sg U9620 ( .A(n8877), .B(n8878), .X(n4426) );
  nand_x1_sg U9621 ( .A(n8875), .B(n8876), .X(n4427) );
  nand_x1_sg U9622 ( .A(n8873), .B(n8874), .X(n4428) );
  nand_x1_sg U9623 ( .A(n8871), .B(n8872), .X(n4429) );
  nand_x1_sg U9624 ( .A(n8869), .B(n8870), .X(n4430) );
  nand_x1_sg U9625 ( .A(n8867), .B(n8868), .X(n4431) );
  nand_x1_sg U9626 ( .A(n8865), .B(n8866), .X(n4432) );
  nand_x1_sg U9627 ( .A(n8863), .B(n8864), .X(n4433) );
  nand_x1_sg U9628 ( .A(n8861), .B(n8862), .X(n4434) );
  nand_x1_sg U9629 ( .A(n8859), .B(n8860), .X(n4435) );
  nand_x1_sg U9630 ( .A(n8857), .B(n8858), .X(n4436) );
  nand_x1_sg U9631 ( .A(n8855), .B(n8856), .X(n4437) );
  nand_x1_sg U9632 ( .A(n8853), .B(n8854), .X(n4438) );
  nand_x1_sg U9633 ( .A(n8851), .B(n8852), .X(n4439) );
  nand_x1_sg U9634 ( .A(n8849), .B(n8850), .X(n4440) );
  nand_x1_sg U9635 ( .A(n8847), .B(n8848), .X(n4441) );
  nand_x1_sg U9636 ( .A(n8845), .B(n8846), .X(n4442) );
  nand_x1_sg U9637 ( .A(n8843), .B(n8844), .X(n4443) );
  nand_x1_sg U9638 ( .A(n8841), .B(n8842), .X(n4444) );
  nand_x1_sg U9639 ( .A(n8839), .B(n8840), .X(n4445) );
  nand_x1_sg U9640 ( .A(n8837), .B(n8838), .X(n4446) );
  nand_x1_sg U9641 ( .A(n8835), .B(n8836), .X(n4447) );
  nand_x1_sg U9642 ( .A(n8833), .B(n8834), .X(n4448) );
  nand_x1_sg U9643 ( .A(n8831), .B(n8832), .X(n4449) );
  nand_x1_sg U9644 ( .A(n8829), .B(n8830), .X(n4450) );
  nand_x1_sg U9645 ( .A(n8827), .B(n8828), .X(n4451) );
  nand_x1_sg U9646 ( .A(n8825), .B(n8826), .X(n4452) );
  nand_x1_sg U9647 ( .A(n8823), .B(n8824), .X(n4453) );
  nand_x1_sg U9648 ( .A(n8821), .B(n8822), .X(n4454) );
  nand_x1_sg U9649 ( .A(n8819), .B(n8820), .X(n4455) );
  nand_x1_sg U9650 ( .A(n8817), .B(n8818), .X(n4456) );
  nand_x1_sg U9651 ( .A(n8815), .B(n8816), .X(n4457) );
  nand_x1_sg U9652 ( .A(n8813), .B(n8814), .X(n4458) );
  nand_x1_sg U9653 ( .A(n8811), .B(n8812), .X(n4459) );
  nand_x1_sg U9654 ( .A(n8809), .B(n8810), .X(n4460) );
  nand_x1_sg U9655 ( .A(n8807), .B(n8808), .X(n4461) );
  nand_x1_sg U9656 ( .A(n8805), .B(n8806), .X(n4462) );
  nand_x1_sg U9657 ( .A(n8803), .B(n8804), .X(n4463) );
  nand_x1_sg U9658 ( .A(n8801), .B(n8802), .X(n4464) );
  nand_x1_sg U9659 ( .A(n8799), .B(n8800), .X(n4465) );
  nand_x1_sg U9660 ( .A(n8797), .B(n8798), .X(n4466) );
  nand_x1_sg U9661 ( .A(n8795), .B(n8796), .X(n4467) );
  nand_x1_sg U9662 ( .A(n8793), .B(n8794), .X(n4468) );
  nand_x1_sg U9663 ( .A(n8791), .B(n8792), .X(n4469) );
  nand_x1_sg U9664 ( .A(n8789), .B(n8790), .X(n4470) );
  nand_x1_sg U9665 ( .A(n8787), .B(n8788), .X(n4471) );
  nand_x1_sg U9666 ( .A(n8785), .B(n8786), .X(n4472) );
  nand_x1_sg U9667 ( .A(n8783), .B(n8784), .X(n4473) );
  nand_x1_sg U9668 ( .A(n8781), .B(n8782), .X(n4474) );
  nand_x1_sg U9669 ( .A(n8779), .B(n8780), .X(n4475) );
  nand_x1_sg U9670 ( .A(n8777), .B(n8778), .X(n4476) );
  nand_x1_sg U9671 ( .A(n8775), .B(n8776), .X(n4477) );
  nand_x1_sg U9672 ( .A(n8773), .B(n8774), .X(n4478) );
  nand_x1_sg U9673 ( .A(n8771), .B(n8772), .X(n4479) );
  nand_x1_sg U9674 ( .A(n8769), .B(n8770), .X(n4480) );
  nand_x1_sg U9675 ( .A(n8767), .B(n8768), .X(n4481) );
  nand_x1_sg U9676 ( .A(n8765), .B(n8766), .X(n4482) );
  nand_x1_sg U9677 ( .A(n8763), .B(n8764), .X(n4483) );
  nand_x1_sg U9678 ( .A(n8761), .B(n8762), .X(n4484) );
  nand_x1_sg U9679 ( .A(n8759), .B(n8760), .X(n4485) );
  nand_x1_sg U9680 ( .A(n8757), .B(n8758), .X(n4486) );
  nand_x1_sg U9681 ( .A(n8755), .B(n8756), .X(n4487) );
  nand_x1_sg U9682 ( .A(n8753), .B(n8754), .X(n4488) );
  nand_x1_sg U9683 ( .A(n8751), .B(n8752), .X(n4489) );
  nand_x1_sg U9684 ( .A(n8749), .B(n8750), .X(n4490) );
  nand_x1_sg U9685 ( .A(n8747), .B(n8748), .X(n4491) );
  nand_x1_sg U9686 ( .A(n8745), .B(n8746), .X(n4492) );
  nand_x1_sg U9687 ( .A(n8743), .B(n8744), .X(n4493) );
  nand_x1_sg U9688 ( .A(n8741), .B(n8742), .X(n4494) );
  nand_x1_sg U9689 ( .A(n8739), .B(n8740), .X(n4495) );
  nand_x1_sg U9690 ( .A(n8737), .B(n8738), .X(n4496) );
  nand_x1_sg U9691 ( .A(n8735), .B(n8736), .X(n4497) );
  nand_x1_sg U9692 ( .A(n8733), .B(n8734), .X(n4498) );
  nand_x1_sg U9693 ( .A(n8731), .B(n8732), .X(n4499) );
  nand_x1_sg U9694 ( .A(n8729), .B(n8730), .X(n4500) );
  nand_x1_sg U9695 ( .A(n8727), .B(n8728), .X(n4501) );
  nand_x1_sg U9696 ( .A(n8725), .B(n8726), .X(n4502) );
  nand_x1_sg U9697 ( .A(n8723), .B(n8724), .X(n4503) );
  nand_x1_sg U9698 ( .A(n8721), .B(n8722), .X(n4504) );
  nand_x1_sg U9699 ( .A(n8717), .B(n8718), .X(n4505) );
  nand_x1_sg U9700 ( .A(n10683), .B(n8713), .X(n4506) );
  nand_x1_sg U9701 ( .A(n8707), .B(n8708), .X(n4507) );
  inv_x1_sg U9702 ( .A(n8380), .X(n11967) );
  inv_x1_sg U9703 ( .A(n8379), .X(n11968) );
  inv_x1_sg U9704 ( .A(n8378), .X(n11969) );
  inv_x1_sg U9705 ( .A(n8377), .X(n11970) );
  inv_x1_sg U9706 ( .A(n8376), .X(n11971) );
  inv_x1_sg U9707 ( .A(n8375), .X(n11972) );
  inv_x1_sg U9708 ( .A(n8374), .X(n11973) );
  inv_x1_sg U9709 ( .A(n8368), .X(n11979) );
  inv_x1_sg U9710 ( .A(n8367), .X(n11980) );
  inv_x1_sg U9711 ( .A(n8366), .X(n11981) );
  inv_x1_sg U9712 ( .A(n8365), .X(n11982) );
  inv_x1_sg U9713 ( .A(n8364), .X(n11983) );
  inv_x1_sg U9714 ( .A(n8363), .X(n11984) );
  inv_x1_sg U9715 ( .A(n8362), .X(n11985) );
  inv_x1_sg U9716 ( .A(n8356), .X(n11991) );
  inv_x1_sg U9717 ( .A(n8355), .X(n11992) );
  inv_x1_sg U9718 ( .A(n8354), .X(n11993) );
  inv_x1_sg U9719 ( .A(n8353), .X(n11994) );
  inv_x1_sg U9720 ( .A(n8352), .X(n11995) );
  inv_x1_sg U9721 ( .A(n8351), .X(n11996) );
  inv_x1_sg U9722 ( .A(n8373), .X(n11974) );
  inv_x1_sg U9723 ( .A(n8372), .X(n11975) );
  inv_x1_sg U9724 ( .A(n8371), .X(n11976) );
  inv_x1_sg U9725 ( .A(n8370), .X(n11977) );
  inv_x1_sg U9726 ( .A(n8369), .X(n11978) );
  inv_x1_sg U9727 ( .A(n8361), .X(n11986) );
  inv_x1_sg U9728 ( .A(n8350), .X(n11997) );
  inv_x1_sg U9729 ( .A(n8349), .X(n11998) );
  inv_x1_sg U9730 ( .A(n8348), .X(n11999) );
  inv_x1_sg U9731 ( .A(n8347), .X(n12000) );
  inv_x1_sg U9732 ( .A(n8346), .X(n12001) );
  inv_x1_sg U9733 ( .A(n8345), .X(n12002) );
  inv_x1_sg U9734 ( .A(n8344), .X(n12003) );
  inv_x1_sg U9735 ( .A(n8337), .X(n12010) );
  inv_x1_sg U9736 ( .A(n8334), .X(n12013) );
  inv_x1_sg U9737 ( .A(n8333), .X(n12014) );
  inv_x1_sg U9738 ( .A(n8332), .X(n12015) );
  inv_x1_sg U9739 ( .A(n8328), .X(n12019) );
  inv_x1_sg U9740 ( .A(n8327), .X(n12020) );
  inv_x1_sg U9741 ( .A(n8326), .X(n12021) );
  inv_x1_sg U9742 ( .A(n8325), .X(n12022) );
  inv_x1_sg U9743 ( .A(n8324), .X(n12023) );
  inv_x1_sg U9744 ( .A(n8323), .X(n12024) );
  inv_x1_sg U9745 ( .A(n8322), .X(n12025) );
  inv_x1_sg U9746 ( .A(n8321), .X(n12026) );
  inv_x1_sg U9747 ( .A(n8360), .X(n11987) );
  inv_x1_sg U9748 ( .A(n8359), .X(n11988) );
  inv_x1_sg U9749 ( .A(n8358), .X(n11989) );
  inv_x1_sg U9750 ( .A(n8357), .X(n11990) );
  inv_x1_sg U9751 ( .A(n8343), .X(n12004) );
  inv_x1_sg U9752 ( .A(n8342), .X(n12005) );
  inv_x1_sg U9753 ( .A(n8336), .X(n12011) );
  inv_x1_sg U9754 ( .A(n8331), .X(n12016) );
  inv_x1_sg U9755 ( .A(n8330), .X(n12017) );
  inv_x1_sg U9756 ( .A(n8329), .X(n12018) );
  inv_x1_sg U9757 ( .A(n8320), .X(n12027) );
  inv_x1_sg U9758 ( .A(n8319), .X(n12028) );
  inv_x1_sg U9759 ( .A(n8318), .X(n12029) );
  inv_x1_sg U9760 ( .A(n8317), .X(n12030) );
  inv_x1_sg U9761 ( .A(n8316), .X(n12031) );
  inv_x1_sg U9762 ( .A(n8315), .X(n12032) );
  inv_x1_sg U9763 ( .A(n8314), .X(n12033) );
  inv_x1_sg U9764 ( .A(n8310), .X(n12037) );
  inv_x1_sg U9765 ( .A(n8309), .X(n12038) );
  inv_x1_sg U9766 ( .A(n8308), .X(n12039) );
  inv_x1_sg U9767 ( .A(n8307), .X(n12040) );
  inv_x1_sg U9768 ( .A(n8294), .X(n12053) );
  inv_x1_sg U9769 ( .A(n8293), .X(n12054) );
  inv_x1_sg U9770 ( .A(n8292), .X(n12055) );
  inv_x1_sg U9771 ( .A(n8291), .X(n12056) );
  inv_x1_sg U9772 ( .A(n8341), .X(n12006) );
  inv_x1_sg U9773 ( .A(n8340), .X(n12007) );
  inv_x1_sg U9774 ( .A(n8339), .X(n12008) );
  inv_x1_sg U9775 ( .A(n8338), .X(n12009) );
  inv_x1_sg U9776 ( .A(n8335), .X(n12012) );
  inv_x1_sg U9777 ( .A(n8313), .X(n12034) );
  inv_x1_sg U9778 ( .A(n8312), .X(n12035) );
  inv_x1_sg U9779 ( .A(n8311), .X(n12036) );
  inv_x1_sg U9780 ( .A(n8300), .X(n12047) );
  inv_x1_sg U9781 ( .A(n8299), .X(n12048) );
  inv_x1_sg U9782 ( .A(n8298), .X(n12049) );
  inv_x1_sg U9783 ( .A(n8297), .X(n12050) );
  inv_x1_sg U9784 ( .A(n8296), .X(n12051) );
  inv_x1_sg U9785 ( .A(n8295), .X(n12052) );
  inv_x1_sg U9786 ( .A(n8290), .X(n12057) );
  inv_x1_sg U9787 ( .A(n8289), .X(n12058) );
  inv_x1_sg U9788 ( .A(n8288), .X(n12059) );
  inv_x1_sg U9789 ( .A(n8287), .X(n12060) );
  inv_x1_sg U9790 ( .A(n8285), .X(n12062) );
  inv_x1_sg U9791 ( .A(n8284), .X(n12063) );
  inv_x1_sg U9792 ( .A(n8283), .X(n12064) );
  inv_x1_sg U9793 ( .A(n8282), .X(n12065) );
  inv_x1_sg U9794 ( .A(n8281), .X(n12066) );
  inv_x1_sg U9795 ( .A(n8280), .X(n12067) );
  inv_x1_sg U9796 ( .A(n8279), .X(n12068) );
  inv_x1_sg U9797 ( .A(n8306), .X(n12041) );
  inv_x1_sg U9798 ( .A(n8305), .X(n12042) );
  inv_x1_sg U9799 ( .A(n8304), .X(n12043) );
  inv_x1_sg U9800 ( .A(n8303), .X(n12044) );
  inv_x1_sg U9801 ( .A(n8302), .X(n12045) );
  inv_x1_sg U9802 ( .A(n8301), .X(n12046) );
  inv_x1_sg U9803 ( .A(n8286), .X(n12061) );
  inv_x1_sg U9804 ( .A(n8278), .X(n12069) );
  inv_x1_sg U9805 ( .A(n8277), .X(n12070) );
  inv_x1_sg U9806 ( .A(n8269), .X(n12078) );
  inv_x1_sg U9807 ( .A(n8268), .X(n12079) );
  inv_x1_sg U9808 ( .A(n8267), .X(n12080) );
  inv_x1_sg U9809 ( .A(n8266), .X(n12081) );
  inv_x1_sg U9810 ( .A(n8265), .X(n12082) );
  inv_x1_sg U9811 ( .A(n8264), .X(n12083) );
  inv_x1_sg U9812 ( .A(n8263), .X(n12084) );
  inv_x1_sg U9813 ( .A(n8262), .X(n12085) );
  inv_x1_sg U9814 ( .A(n8260), .X(n12087) );
  inv_x1_sg U9815 ( .A(n8259), .X(n12088) );
  inv_x1_sg U9816 ( .A(n8258), .X(n12089) );
  inv_x1_sg U9817 ( .A(n8257), .X(n12090) );
  inv_x1_sg U9818 ( .A(n8256), .X(n12091) );
  inv_x1_sg U9819 ( .A(n8251), .X(n12096) );
  inv_x1_sg U9820 ( .A(n8250), .X(n12097) );
  inv_x1_sg U9821 ( .A(n8249), .X(n12098) );
  inv_x1_sg U9822 ( .A(n8276), .X(n12071) );
  inv_x1_sg U9823 ( .A(n8275), .X(n12072) );
  inv_x1_sg U9824 ( .A(n8274), .X(n12073) );
  inv_x1_sg U9825 ( .A(n8273), .X(n12074) );
  inv_x1_sg U9826 ( .A(n8272), .X(n12075) );
  inv_x1_sg U9827 ( .A(n8271), .X(n12076) );
  inv_x1_sg U9828 ( .A(n8270), .X(n12077) );
  inv_x1_sg U9829 ( .A(n8261), .X(n12086) );
  inv_x1_sg U9830 ( .A(n8255), .X(n12092) );
  inv_x1_sg U9831 ( .A(n8254), .X(n12093) );
  inv_x1_sg U9832 ( .A(n8253), .X(n12094) );
  inv_x1_sg U9833 ( .A(n8252), .X(n12095) );
  inv_x1_sg U9834 ( .A(n8248), .X(n12099) );
  inv_x1_sg U9835 ( .A(n8247), .X(n12100) );
  inv_x1_sg U9836 ( .A(n8238), .X(n12109) );
  inv_x1_sg U9837 ( .A(n8237), .X(n12110) );
  inv_x1_sg U9838 ( .A(n8235), .X(n12112) );
  inv_x1_sg U9839 ( .A(n8234), .X(n12113) );
  inv_x1_sg U9840 ( .A(n8233), .X(n12114) );
  inv_x1_sg U9841 ( .A(n8231), .X(n12116) );
  inv_x1_sg U9842 ( .A(n8230), .X(n12117) );
  inv_x1_sg U9843 ( .A(n8229), .X(n12118) );
  inv_x1_sg U9844 ( .A(n8228), .X(n12119) );
  inv_x1_sg U9845 ( .A(n8227), .X(n12120) );
  inv_x1_sg U9846 ( .A(n8226), .X(n12121) );
  inv_x1_sg U9847 ( .A(n8246), .X(n12101) );
  inv_x1_sg U9848 ( .A(n8245), .X(n12102) );
  inv_x1_sg U9849 ( .A(n8244), .X(n12103) );
  inv_x1_sg U9850 ( .A(n8243), .X(n12104) );
  inv_x1_sg U9851 ( .A(n8242), .X(n12105) );
  inv_x1_sg U9852 ( .A(n8241), .X(n12106) );
  inv_x1_sg U9853 ( .A(n8240), .X(n12107) );
  inv_x1_sg U9854 ( .A(n8239), .X(n12108) );
  inv_x1_sg U9855 ( .A(n8236), .X(n12111) );
  inv_x1_sg U9856 ( .A(n8232), .X(n12115) );
  inv_x1_sg U9857 ( .A(n8225), .X(n12122) );
  inv_x1_sg U9858 ( .A(n8224), .X(n12123) );
  inv_x1_sg U9859 ( .A(n8223), .X(n12124) );
  inv_x1_sg U9860 ( .A(n8222), .X(n12125) );
  inv_x1_sg U9861 ( .A(n8221), .X(n12126) );
  inv_x1_sg U9862 ( .A(n8220), .X(n12127) );
  inv_x1_sg U9863 ( .A(n8219), .X(n12128) );
  inv_x1_sg U9864 ( .A(n8217), .X(n12130) );
  inv_x1_sg U9865 ( .A(n8211), .X(n12136) );
  inv_x1_sg U9866 ( .A(n8201), .X(n12146) );
  inv_x1_sg U9867 ( .A(n8200), .X(n12147) );
  inv_x1_sg U9868 ( .A(n8199), .X(n12148) );
  inv_x1_sg U9869 ( .A(n8198), .X(n12149) );
  inv_x1_sg U9870 ( .A(n8197), .X(n12150) );
  inv_x1_sg U9871 ( .A(n8196), .X(n12151) );
  inv_x1_sg U9872 ( .A(n8218), .X(n12129) );
  inv_x1_sg U9873 ( .A(n8216), .X(n12131) );
  inv_x1_sg U9874 ( .A(n8215), .X(n12132) );
  inv_x1_sg U9875 ( .A(n8214), .X(n12133) );
  inv_x1_sg U9876 ( .A(n8213), .X(n12134) );
  inv_x1_sg U9877 ( .A(n8212), .X(n12135) );
  inv_x1_sg U9878 ( .A(n8210), .X(n12137) );
  inv_x1_sg U9879 ( .A(n8206), .X(n12141) );
  inv_x1_sg U9880 ( .A(n8205), .X(n12142) );
  inv_x1_sg U9881 ( .A(n8204), .X(n12143) );
  inv_x1_sg U9882 ( .A(n8203), .X(n12144) );
  inv_x1_sg U9883 ( .A(n8202), .X(n12145) );
  inv_x1_sg U9884 ( .A(n8195), .X(n12152) );
  inv_x1_sg U9885 ( .A(n8194), .X(n12153) );
  inv_x1_sg U9886 ( .A(n8193), .X(n12154) );
  inv_x1_sg U9887 ( .A(n8192), .X(n12155) );
  inv_x1_sg U9888 ( .A(n8191), .X(n12156) );
  inv_x1_sg U9889 ( .A(n8190), .X(n12157) );
  inv_x1_sg U9890 ( .A(n8189), .X(n12158) );
  inv_x1_sg U9891 ( .A(n8186), .X(n12161) );
  inv_x1_sg U9892 ( .A(n8170), .X(n12177) );
  inv_x1_sg U9893 ( .A(n8169), .X(n12178) );
  inv_x1_sg U9894 ( .A(n8168), .X(n12179) );
  inv_x1_sg U9895 ( .A(n8167), .X(n12180) );
  inv_x1_sg U9896 ( .A(n8166), .X(n12181) );
  inv_x1_sg U9897 ( .A(n8209), .X(n12138) );
  inv_x1_sg U9898 ( .A(n8208), .X(n12139) );
  inv_x1_sg U9899 ( .A(n8207), .X(n12140) );
  inv_x1_sg U9900 ( .A(n8188), .X(n12159) );
  inv_x1_sg U9901 ( .A(n8187), .X(n12160) );
  inv_x1_sg U9902 ( .A(n8185), .X(n12162) );
  inv_x1_sg U9903 ( .A(n8184), .X(n12163) );
  inv_x1_sg U9904 ( .A(n8183), .X(n12164) );
  inv_x1_sg U9905 ( .A(n8182), .X(n12165) );
  inv_x1_sg U9906 ( .A(n8174), .X(n12173) );
  inv_x1_sg U9907 ( .A(n8173), .X(n12174) );
  inv_x1_sg U9908 ( .A(n8172), .X(n12175) );
  inv_x1_sg U9909 ( .A(n8171), .X(n12176) );
  inv_x1_sg U9910 ( .A(n8165), .X(n12182) );
  inv_x1_sg U9911 ( .A(n8164), .X(n12183) );
  inv_x1_sg U9912 ( .A(n8163), .X(n12184) );
  inv_x1_sg U9913 ( .A(n8162), .X(n12185) );
  inv_x1_sg U9914 ( .A(n8161), .X(n12186) );
  inv_x1_sg U9915 ( .A(n8156), .X(n12191) );
  inv_x1_sg U9916 ( .A(n8155), .X(n12192) );
  inv_x1_sg U9917 ( .A(n8154), .X(n12193) );
  inv_x1_sg U9918 ( .A(n8139), .X(n12208) );
  inv_x1_sg U9919 ( .A(n8138), .X(n12209) );
  inv_x1_sg U9920 ( .A(n8137), .X(n12210) );
  inv_x1_sg U9921 ( .A(n8131), .X(n12216) );
  inv_x1_sg U9922 ( .A(n8181), .X(n12166) );
  inv_x1_sg U9923 ( .A(n8180), .X(n12167) );
  inv_x1_sg U9924 ( .A(n8179), .X(n12168) );
  inv_x1_sg U9925 ( .A(n8178), .X(n12169) );
  inv_x1_sg U9926 ( .A(n8177), .X(n12170) );
  inv_x1_sg U9927 ( .A(n8176), .X(n12171) );
  inv_x1_sg U9928 ( .A(n8175), .X(n12172) );
  inv_x1_sg U9929 ( .A(n8160), .X(n12187) );
  inv_x1_sg U9930 ( .A(n8159), .X(n12188) );
  inv_x1_sg U9931 ( .A(n8158), .X(n12189) );
  inv_x1_sg U9932 ( .A(n8157), .X(n12190) );
  inv_x1_sg U9933 ( .A(n8153), .X(n12194) );
  inv_x1_sg U9934 ( .A(n8152), .X(n12195) );
  inv_x1_sg U9935 ( .A(n8140), .X(n12207) );
  inv_x1_sg U9936 ( .A(n8136), .X(n12211) );
  inv_x1_sg U9937 ( .A(n8133), .X(n12214) );
  inv_x1_sg U9938 ( .A(n8132), .X(n12215) );
  inv_x1_sg U9939 ( .A(n8130), .X(n12217) );
  inv_x1_sg U9940 ( .A(n8129), .X(n12218) );
  inv_x1_sg U9941 ( .A(n8128), .X(n12219) );
  inv_x1_sg U9942 ( .A(n8127), .X(n12220) );
  inv_x1_sg U9943 ( .A(n8126), .X(n12221) );
  inv_x1_sg U9944 ( .A(n8125), .X(n12222) );
  inv_x1_sg U9945 ( .A(n8124), .X(n12223) );
  inv_x1_sg U9946 ( .A(n8110), .X(n12237) );
  inv_x1_sg U9947 ( .A(n8151), .X(n12196) );
  inv_x1_sg U9948 ( .A(n8150), .X(n12197) );
  inv_x1_sg U9949 ( .A(n8149), .X(n12198) );
  inv_x1_sg U9950 ( .A(n8148), .X(n12199) );
  inv_x1_sg U9951 ( .A(n8147), .X(n12200) );
  inv_x1_sg U9952 ( .A(n8146), .X(n12201) );
  inv_x1_sg U9953 ( .A(n8145), .X(n12202) );
  inv_x1_sg U9954 ( .A(n8144), .X(n12203) );
  inv_x1_sg U9955 ( .A(n8143), .X(n12204) );
  inv_x1_sg U9956 ( .A(n8142), .X(n12205) );
  inv_x1_sg U9957 ( .A(n8141), .X(n12206) );
  inv_x1_sg U9958 ( .A(n8135), .X(n12212) );
  inv_x1_sg U9959 ( .A(n8134), .X(n12213) );
  inv_x1_sg U9960 ( .A(n8123), .X(n12224) );
  inv_x1_sg U9961 ( .A(n8122), .X(n12225) );
  inv_x1_sg U9962 ( .A(n8111), .X(n12236) );
  inv_x1_sg U9963 ( .A(n8109), .X(n12238) );
  inv_x1_sg U9964 ( .A(n8108), .X(n12239) );
  inv_x1_sg U9965 ( .A(n8107), .X(n12240) );
  inv_x1_sg U9966 ( .A(n8102), .X(n12245) );
  inv_x1_sg U9967 ( .A(n8101), .X(n12246) );
  inv_x1_sg U9968 ( .A(n8097), .X(n12250) );
  inv_x1_sg U9969 ( .A(n8096), .X(n12251) );
  inv_x1_sg U9970 ( .A(n8095), .X(n12252) );
  inv_x1_sg U9971 ( .A(n8094), .X(n12253) );
  inv_x1_sg U9972 ( .A(n8121), .X(n12226) );
  inv_x1_sg U9973 ( .A(n8120), .X(n12227) );
  inv_x1_sg U9974 ( .A(n8119), .X(n12228) );
  inv_x1_sg U9975 ( .A(n8118), .X(n12229) );
  inv_x1_sg U9976 ( .A(n8117), .X(n12230) );
  inv_x1_sg U9977 ( .A(n8116), .X(n12231) );
  inv_x1_sg U9978 ( .A(n8115), .X(n12232) );
  inv_x1_sg U9979 ( .A(n8114), .X(n12233) );
  inv_x1_sg U9980 ( .A(n8113), .X(n12234) );
  inv_x1_sg U9981 ( .A(n8112), .X(n12235) );
  inv_x1_sg U9982 ( .A(n8106), .X(n12241) );
  inv_x1_sg U9983 ( .A(n8105), .X(n12242) );
  inv_x1_sg U9984 ( .A(n8104), .X(n12243) );
  inv_x1_sg U9985 ( .A(n8103), .X(n12244) );
  inv_x1_sg U9986 ( .A(n8100), .X(n12247) );
  inv_x1_sg U9987 ( .A(n8099), .X(n12248) );
  inv_x1_sg U9988 ( .A(n8098), .X(n12249) );
  inv_x1_sg U9989 ( .A(n8093), .X(n12254) );
  inv_x1_sg U9990 ( .A(n8092), .X(n12255) );
  inv_x1_sg U9991 ( .A(n8086), .X(n12261) );
  inv_x1_sg U9992 ( .A(n8085), .X(n12262) );
  inv_x1_sg U9993 ( .A(n8084), .X(n12263) );
  inv_x1_sg U9994 ( .A(n8083), .X(n12264) );
  inv_x1_sg U9995 ( .A(n8082), .X(n12265) );
  inv_x1_sg U9996 ( .A(n8071), .X(n12276) );
  inv_x1_sg U9997 ( .A(n8091), .X(n12256) );
  inv_x1_sg U9998 ( .A(n8090), .X(n12257) );
  inv_x1_sg U9999 ( .A(n8089), .X(n12258) );
  inv_x1_sg U10000 ( .A(n8088), .X(n12259) );
  inv_x1_sg U10001 ( .A(n8087), .X(n12260) );
  inv_x1_sg U10002 ( .A(n8081), .X(n12266) );
  inv_x1_sg U10003 ( .A(n8080), .X(n12267) );
  inv_x1_sg U10004 ( .A(n8079), .X(n12268) );
  inv_x1_sg U10005 ( .A(n8078), .X(n12269) );
  inv_x1_sg U10006 ( .A(n8077), .X(n12270) );
  inv_x1_sg U10007 ( .A(n8076), .X(n12271) );
  inv_x1_sg U10008 ( .A(n8075), .X(n12272) );
  inv_x1_sg U10009 ( .A(n8074), .X(n12273) );
  inv_x1_sg U10010 ( .A(n8073), .X(n12274) );
  inv_x1_sg U10011 ( .A(n8072), .X(n12275) );
  inv_x1_sg U10012 ( .A(n8070), .X(n12277) );
  inv_x1_sg U10013 ( .A(n8069), .X(n12278) );
  inv_x1_sg U10014 ( .A(n8068), .X(n12279) );
  inv_x1_sg U10015 ( .A(n8067), .X(n12280) );
  inv_x1_sg U10016 ( .A(n8066), .X(n12281) );
  inv_x1_sg U10017 ( .A(n8065), .X(n12282) );
  inv_x1_sg U10018 ( .A(n8064), .X(n12283) );
  inv_x1_sg U10019 ( .A(n8063), .X(n12284) );
  inv_x1_sg U10020 ( .A(n8062), .X(n12285) );
  inv_x1_sg U10021 ( .A(n8381), .X(n11966) );
  nor_x1_sg U10022 ( .A(n9359), .B(n8715), .X(n10685) );
  nor_x1_sg U10023 ( .A(n10550), .B(n10684), .X(n8716) );
  nor_x1_sg U10024 ( .A(n10682), .B(n10410), .X(n8719) );
  nor_x1_sg U10025 ( .A(n10682), .B(n8714), .X(n8711) );
  nand_x1_sg U10026 ( .A(n10546), .B(n8715), .X(n8714) );
  nand_x1_sg U10027 ( .A(n12286), .B(n8710), .X(n9359) );
  nand_x1_sg U10028 ( .A(\out[0][1][7] ), .B(n10053), .X(n9946) );
  nand_x1_sg U10029 ( .A(n10349), .B(n3574), .X(n9943) );
  nand_x1_sg U10030 ( .A(\out[0][1][8] ), .B(n10274), .X(n9944) );
  nand_x1_sg U10031 ( .A(n10355), .B(n3575), .X(n9941) );
  nand_x1_sg U10032 ( .A(\out[0][1][9] ), .B(n10223), .X(n9942) );
  nand_x1_sg U10033 ( .A(n10674), .B(n3603), .X(n9885) );
  nand_x1_sg U10034 ( .A(\out[0][2][17] ), .B(n10222), .X(n9886) );
  nand_x1_sg U10035 ( .A(n10658), .B(n3604), .X(n9883) );
  nand_x1_sg U10036 ( .A(\out[0][2][18] ), .B(n10515), .X(n9884) );
  nand_x1_sg U10037 ( .A(n10658), .B(n3605), .X(n9881) );
  nand_x1_sg U10038 ( .A(\out[0][2][19] ), .B(n10470), .X(n9882) );
  nand_x1_sg U10039 ( .A(n10380), .B(n3633), .X(n9825) );
  nand_x1_sg U10040 ( .A(\out[1][0][7] ), .B(n10470), .X(n9826) );
  nand_x1_sg U10041 ( .A(n10100), .B(n3634), .X(n9823) );
  nand_x1_sg U10042 ( .A(\out[1][0][8] ), .B(n10507), .X(n9824) );
  nand_x1_sg U10043 ( .A(n10368), .B(n3635), .X(n9821) );
  nand_x1_sg U10044 ( .A(\out[1][0][9] ), .B(n10507), .X(n9822) );
  nand_x1_sg U10045 ( .A(n10089), .B(n3643), .X(n9805) );
  nand_x1_sg U10046 ( .A(\out[1][0][17] ), .B(n10463), .X(n9806) );
  nand_x1_sg U10047 ( .A(\out[1][2][0] ), .B(n10052), .X(n9760) );
  nand_x1_sg U10048 ( .A(n10646), .B(n3667), .X(n9757) );
  nand_x1_sg U10049 ( .A(\out[1][2][1] ), .B(n10515), .X(n9758) );
  nand_x1_sg U10050 ( .A(n10644), .B(n3698), .X(n9695) );
  nand_x1_sg U10051 ( .A(\out[1][3][12] ), .B(n10225), .X(n9696) );
  nand_x1_sg U10052 ( .A(n10379), .B(n3699), .X(n9693) );
  nand_x1_sg U10053 ( .A(\out[1][3][13] ), .B(n10276), .X(n9694) );
  nand_x1_sg U10054 ( .A(n10378), .B(n3700), .X(n9691) );
  nand_x1_sg U10055 ( .A(\out[1][3][14] ), .B(n10136), .X(n9692) );
  nand_x1_sg U10056 ( .A(n10313), .B(n3719), .X(n9653) );
  nand_x1_sg U10057 ( .A(\out[2][0][13] ), .B(n10050), .X(n9654) );
  nand_x1_sg U10058 ( .A(n10370), .B(n3720), .X(n9651) );
  nand_x1_sg U10059 ( .A(\out[2][0][14] ), .B(n10593), .X(n9652) );
  nand_x1_sg U10060 ( .A(n10353), .B(n3728), .X(n9635) );
  nand_x1_sg U10061 ( .A(\out[2][1][2] ), .B(n10281), .X(n9636) );
  nand_x1_sg U10062 ( .A(n10657), .B(n3729), .X(n9633) );
  nand_x1_sg U10063 ( .A(\out[2][1][3] ), .B(n10589), .X(n9634) );
  nand_x1_sg U10064 ( .A(n10655), .B(n3730), .X(n9631) );
  nand_x1_sg U10065 ( .A(\out[2][1][4] ), .B(n10464), .X(n9632) );
  nand_x1_sg U10066 ( .A(n10102), .B(n3758), .X(n9575) );
  nand_x1_sg U10067 ( .A(\out[2][2][12] ), .B(n10521), .X(n9576) );
  nand_x1_sg U10068 ( .A(n10102), .B(n3759), .X(n9573) );
  nand_x1_sg U10069 ( .A(\out[2][2][13] ), .B(n10271), .X(n9574) );
  nand_x1_sg U10070 ( .A(n10352), .B(n3760), .X(n9571) );
  nand_x1_sg U10071 ( .A(\out[2][2][14] ), .B(n10039), .X(n9572) );
  nand_x1_sg U10072 ( .A(n10313), .B(n3788), .X(n9515) );
  nand_x1_sg U10073 ( .A(\out[3][0][2] ), .B(n10293), .X(n9516) );
  nand_x1_sg U10074 ( .A(n10646), .B(n3789), .X(n9513) );
  nand_x1_sg U10075 ( .A(\out[3][0][3] ), .B(n10521), .X(n9514) );
  nand_x1_sg U10076 ( .A(\out[3][0][4] ), .B(n10049), .X(n9512) );
  nand_x1_sg U10077 ( .A(n10650), .B(n3853), .X(n9385) );
  nand_x1_sg U10078 ( .A(\out[3][3][7] ), .B(n10469), .X(n9386) );
  nand_x1_sg U10079 ( .A(n10372), .B(n3854), .X(n9383) );
  nand_x1_sg U10080 ( .A(\out[3][3][8] ), .B(n10053), .X(n9384) );
  nand_x1_sg U10081 ( .A(n10352), .B(n3855), .X(n9381) );
  nand_x1_sg U10082 ( .A(\out[3][3][9] ), .B(n10052), .X(n9382) );
  nand_x1_sg U10083 ( .A(n10661), .B(n3546), .X(n9999) );
  nand_x1_sg U10084 ( .A(\out[0][0][0] ), .B(n10510), .X(n10000) );
  nand_x1_sg U10085 ( .A(n10659), .B(n3547), .X(n9997) );
  nand_x1_sg U10086 ( .A(\out[0][0][1] ), .B(n10504), .X(n9998) );
  nand_x1_sg U10087 ( .A(n10377), .B(n3548), .X(n9995) );
  nand_x1_sg U10088 ( .A(\out[0][0][2] ), .B(n10275), .X(n9996) );
  nand_x1_sg U10089 ( .A(n10108), .B(n3549), .X(n9993) );
  nand_x1_sg U10090 ( .A(\out[0][0][3] ), .B(n10135), .X(n9994) );
  nand_x1_sg U10091 ( .A(n10644), .B(n3550), .X(n9991) );
  nand_x1_sg U10092 ( .A(\out[0][0][4] ), .B(n10508), .X(n9992) );
  nand_x1_sg U10093 ( .A(n10647), .B(n3551), .X(n9989) );
  nand_x1_sg U10094 ( .A(\out[0][0][5] ), .B(n10174), .X(n9990) );
  nand_x1_sg U10095 ( .A(n10356), .B(n3552), .X(n9987) );
  nand_x1_sg U10096 ( .A(\out[0][0][6] ), .B(n10166), .X(n9988) );
  nand_x1_sg U10097 ( .A(n10645), .B(n3553), .X(n9985) );
  nand_x1_sg U10098 ( .A(\out[0][0][7] ), .B(n10471), .X(n9986) );
  nand_x1_sg U10099 ( .A(n10091), .B(n3554), .X(n9983) );
  nand_x1_sg U10100 ( .A(\out[0][0][8] ), .B(n10472), .X(n9984) );
  nand_x1_sg U10101 ( .A(n10353), .B(n3557), .X(n9977) );
  nand_x1_sg U10102 ( .A(\out[0][0][11] ), .B(n10273), .X(n9978) );
  nand_x1_sg U10103 ( .A(n10362), .B(n3558), .X(n9975) );
  nand_x1_sg U10104 ( .A(\out[0][0][12] ), .B(n10166), .X(n9976) );
  nand_x1_sg U10105 ( .A(n10672), .B(n3559), .X(n9973) );
  nand_x1_sg U10106 ( .A(\out[0][0][13] ), .B(n10299), .X(n9974) );
  nand_x1_sg U10107 ( .A(n10353), .B(n3560), .X(n9971) );
  nand_x1_sg U10108 ( .A(\out[0][0][14] ), .B(n10284), .X(n9972) );
  nand_x1_sg U10109 ( .A(n10368), .B(n3561), .X(n9969) );
  nand_x1_sg U10110 ( .A(\out[0][0][15] ), .B(n10219), .X(n9970) );
  nand_x1_sg U10111 ( .A(n10661), .B(n3562), .X(n9967) );
  nand_x1_sg U10112 ( .A(\out[0][0][16] ), .B(n10297), .X(n9968) );
  nand_x1_sg U10113 ( .A(n10657), .B(n3563), .X(n9965) );
  nand_x1_sg U10114 ( .A(\out[0][0][17] ), .B(n10038), .X(n9966) );
  nand_x1_sg U10115 ( .A(n10646), .B(n3564), .X(n9963) );
  nand_x1_sg U10116 ( .A(\out[0][0][18] ), .B(n10162), .X(n9964) );
  nand_x1_sg U10117 ( .A(n10105), .B(n3565), .X(n9961) );
  nand_x1_sg U10118 ( .A(\out[0][0][19] ), .B(n10048), .X(n9962) );
  nand_x1_sg U10119 ( .A(n10379), .B(n3566), .X(n9959) );
  nand_x1_sg U10120 ( .A(\out[0][1][0] ), .B(n10465), .X(n9960) );
  nand_x1_sg U10121 ( .A(n10405), .B(n3567), .X(n9957) );
  nand_x1_sg U10122 ( .A(\out[0][1][1] ), .B(n10039), .X(n9958) );
  nand_x1_sg U10123 ( .A(n10355), .B(n3568), .X(n9955) );
  nand_x1_sg U10124 ( .A(\out[0][1][2] ), .B(n10132), .X(n9956) );
  nand_x1_sg U10125 ( .A(n10104), .B(n3570), .X(n9951) );
  nand_x1_sg U10126 ( .A(\out[0][1][4] ), .B(n10505), .X(n9952) );
  nand_x1_sg U10127 ( .A(n10644), .B(n3571), .X(n9949) );
  nand_x1_sg U10128 ( .A(\out[0][1][5] ), .B(n10161), .X(n9950) );
  nand_x1_sg U10129 ( .A(n10371), .B(n3572), .X(n9947) );
  nand_x1_sg U10130 ( .A(\out[0][1][6] ), .B(n10273), .X(n9948) );
  nand_x1_sg U10131 ( .A(n10355), .B(n3576), .X(n9939) );
  nand_x1_sg U10132 ( .A(\out[0][1][10] ), .B(n10298), .X(n9940) );
  nand_x1_sg U10133 ( .A(n10376), .B(n3577), .X(n9937) );
  nand_x1_sg U10134 ( .A(\out[0][1][11] ), .B(n10299), .X(n9938) );
  nand_x1_sg U10135 ( .A(n10107), .B(n3578), .X(n9935) );
  nand_x1_sg U10136 ( .A(\out[0][1][12] ), .B(n10170), .X(n9936) );
  nand_x1_sg U10137 ( .A(n10649), .B(n3579), .X(n9933) );
  nand_x1_sg U10138 ( .A(\out[0][1][13] ), .B(n10584), .X(n9934) );
  nand_x1_sg U10139 ( .A(n10370), .B(n3580), .X(n9931) );
  nand_x1_sg U10140 ( .A(\out[0][1][14] ), .B(n10507), .X(n9932) );
  nand_x1_sg U10141 ( .A(n10346), .B(n3581), .X(n9929) );
  nand_x1_sg U10142 ( .A(\out[0][1][15] ), .B(n10223), .X(n9930) );
  nand_x1_sg U10143 ( .A(n10089), .B(n3587), .X(n9917) );
  nand_x1_sg U10144 ( .A(\out[0][2][1] ), .B(n10171), .X(n9918) );
  nand_x1_sg U10145 ( .A(n10370), .B(n3588), .X(n9915) );
  nand_x1_sg U10146 ( .A(\out[0][2][2] ), .B(n10296), .X(n9916) );
  nand_x1_sg U10147 ( .A(n10671), .B(n3589), .X(n9913) );
  nand_x1_sg U10148 ( .A(\out[0][2][3] ), .B(n10466), .X(n9914) );
  nand_x1_sg U10149 ( .A(n10645), .B(n3590), .X(n9911) );
  nand_x1_sg U10150 ( .A(\out[0][2][4] ), .B(n10590), .X(n9912) );
  nand_x1_sg U10151 ( .A(n10360), .B(n3591), .X(n9909) );
  nand_x1_sg U10152 ( .A(\out[0][2][5] ), .B(n10588), .X(n9910) );
  nand_x1_sg U10153 ( .A(n10361), .B(n3592), .X(n9907) );
  nand_x1_sg U10154 ( .A(\out[0][2][6] ), .B(n10590), .X(n9908) );
  nand_x1_sg U10155 ( .A(n10659), .B(n3593), .X(n9905) );
  nand_x1_sg U10156 ( .A(\out[0][2][7] ), .B(n10515), .X(n9906) );
  nand_x1_sg U10157 ( .A(n10365), .B(n3594), .X(n9903) );
  nand_x1_sg U10158 ( .A(\out[0][2][8] ), .B(n10173), .X(n9904) );
  nand_x1_sg U10159 ( .A(n10384), .B(n3595), .X(n9901) );
  nand_x1_sg U10160 ( .A(\out[0][2][9] ), .B(n10293), .X(n9902) );
  nand_x1_sg U10161 ( .A(n10648), .B(n3596), .X(n9899) );
  nand_x1_sg U10162 ( .A(\out[0][2][10] ), .B(n10585), .X(n9900) );
  nand_x1_sg U10163 ( .A(n10361), .B(n3597), .X(n9897) );
  nand_x1_sg U10164 ( .A(\out[0][2][11] ), .B(n10050), .X(n9898) );
  nand_x1_sg U10165 ( .A(n10102), .B(n3598), .X(n9895) );
  nand_x1_sg U10166 ( .A(\out[0][2][12] ), .B(n10276), .X(n9896) );
  nand_x1_sg U10167 ( .A(n10662), .B(n3599), .X(n9893) );
  nand_x1_sg U10168 ( .A(\out[0][2][13] ), .B(n10515), .X(n9894) );
  nand_x1_sg U10169 ( .A(n10108), .B(n3600), .X(n9891) );
  nand_x1_sg U10170 ( .A(\out[0][2][14] ), .B(n10504), .X(n9892) );
  nand_x1_sg U10171 ( .A(n10365), .B(n3601), .X(n9889) );
  nand_x1_sg U10172 ( .A(\out[0][2][15] ), .B(n10472), .X(n9890) );
  nand_x1_sg U10173 ( .A(n10667), .B(n3602), .X(n9887) );
  nand_x1_sg U10174 ( .A(\out[0][2][16] ), .B(n10594), .X(n9888) );
  nand_x1_sg U10175 ( .A(n10100), .B(n3606), .X(n9879) );
  nand_x1_sg U10176 ( .A(\out[0][3][0] ), .B(n10468), .X(n9880) );
  nand_x1_sg U10177 ( .A(n10314), .B(n3607), .X(n9877) );
  nand_x1_sg U10178 ( .A(\out[0][3][1] ), .B(n10273), .X(n9878) );
  nand_x1_sg U10179 ( .A(n10356), .B(n3608), .X(n9875) );
  nand_x1_sg U10180 ( .A(\out[0][3][2] ), .B(n10047), .X(n9876) );
  nand_x1_sg U10181 ( .A(n10367), .B(n3609), .X(n9873) );
  nand_x1_sg U10182 ( .A(\out[0][3][3] ), .B(n10463), .X(n9874) );
  nand_x1_sg U10183 ( .A(n10383), .B(n3610), .X(n9871) );
  nand_x1_sg U10184 ( .A(\out[0][3][4] ), .B(n10462), .X(n9872) );
  nand_x1_sg U10185 ( .A(n10670), .B(n3611), .X(n9869) );
  nand_x1_sg U10186 ( .A(\out[0][3][5] ), .B(n10275), .X(n9870) );
  nand_x1_sg U10187 ( .A(n10378), .B(n3612), .X(n9867) );
  nand_x1_sg U10188 ( .A(\out[0][3][6] ), .B(n10294), .X(n9868) );
  nand_x1_sg U10189 ( .A(n10673), .B(n3613), .X(n9865) );
  nand_x1_sg U10190 ( .A(\out[0][3][7] ), .B(n10469), .X(n9866) );
  nand_x1_sg U10191 ( .A(n10365), .B(n3614), .X(n9863) );
  nand_x1_sg U10192 ( .A(\out[0][3][8] ), .B(n10282), .X(n9864) );
  nand_x1_sg U10193 ( .A(n10352), .B(n3616), .X(n9859) );
  nand_x1_sg U10194 ( .A(\out[0][3][10] ), .B(n10131), .X(n9860) );
  nand_x1_sg U10195 ( .A(n10371), .B(n3617), .X(n9857) );
  nand_x1_sg U10196 ( .A(\out[0][3][11] ), .B(n10586), .X(n9858) );
  nand_x1_sg U10197 ( .A(n10313), .B(n3618), .X(n9855) );
  nand_x1_sg U10198 ( .A(\out[0][3][12] ), .B(n10520), .X(n9856) );
  nand_x1_sg U10199 ( .A(n10670), .B(n3619), .X(n9853) );
  nand_x1_sg U10200 ( .A(\out[0][3][13] ), .B(n10590), .X(n9854) );
  nand_x1_sg U10201 ( .A(n10662), .B(n3620), .X(n9851) );
  nand_x1_sg U10202 ( .A(\out[0][3][14] ), .B(n10165), .X(n9852) );
  nand_x1_sg U10203 ( .A(n10674), .B(n3626), .X(n9839) );
  nand_x1_sg U10204 ( .A(\out[1][0][0] ), .B(n10047), .X(n9840) );
  nand_x1_sg U10205 ( .A(n10342), .B(n3627), .X(n9837) );
  nand_x1_sg U10206 ( .A(\out[1][0][1] ), .B(n10465), .X(n9838) );
  nand_x1_sg U10207 ( .A(n10348), .B(n3628), .X(n9835) );
  nand_x1_sg U10208 ( .A(\out[1][0][2] ), .B(n10281), .X(n9836) );
  nand_x1_sg U10209 ( .A(n10262), .B(n3629), .X(n9833) );
  nand_x1_sg U10210 ( .A(\out[1][0][3] ), .B(n10471), .X(n9834) );
  nand_x1_sg U10211 ( .A(n10104), .B(n3630), .X(n9831) );
  nand_x1_sg U10212 ( .A(\out[1][0][4] ), .B(n10173), .X(n9832) );
  nand_x1_sg U10213 ( .A(n10374), .B(n3631), .X(n9829) );
  nand_x1_sg U10214 ( .A(\out[1][0][5] ), .B(n10463), .X(n9830) );
  nand_x1_sg U10215 ( .A(n10353), .B(n3632), .X(n9827) );
  nand_x1_sg U10216 ( .A(\out[1][0][6] ), .B(n10298), .X(n9828) );
  nand_x1_sg U10217 ( .A(n10377), .B(n3636), .X(n9819) );
  nand_x1_sg U10218 ( .A(\out[1][0][10] ), .B(n10506), .X(n9820) );
  nand_x1_sg U10219 ( .A(n10376), .B(n3637), .X(n9817) );
  nand_x1_sg U10220 ( .A(\out[1][0][11] ), .B(n10282), .X(n9818) );
  nand_x1_sg U10221 ( .A(n10102), .B(n3638), .X(n9815) );
  nand_x1_sg U10222 ( .A(\out[1][0][12] ), .B(n10513), .X(n9816) );
  nand_x1_sg U10223 ( .A(n10668), .B(n3639), .X(n9813) );
  nand_x1_sg U10224 ( .A(\out[1][0][13] ), .B(n10224), .X(n9814) );
  nand_x1_sg U10225 ( .A(n10649), .B(n3640), .X(n9811) );
  nand_x1_sg U10226 ( .A(\out[1][0][14] ), .B(n10131), .X(n9812) );
  nand_x1_sg U10227 ( .A(n10105), .B(n3641), .X(n9809) );
  nand_x1_sg U10228 ( .A(\out[1][0][15] ), .B(n10506), .X(n9810) );
  nand_x1_sg U10229 ( .A(n10382), .B(n3642), .X(n9807) );
  nand_x1_sg U10230 ( .A(\out[1][0][16] ), .B(n10038), .X(n9808) );
  nand_x1_sg U10231 ( .A(n10406), .B(n3644), .X(n9803) );
  nand_x1_sg U10232 ( .A(\out[1][0][18] ), .B(n10593), .X(n9804) );
  nand_x1_sg U10233 ( .A(n10666), .B(n3645), .X(n9801) );
  nand_x1_sg U10234 ( .A(\out[1][0][19] ), .B(n10466), .X(n9802) );
  nand_x1_sg U10235 ( .A(n10354), .B(n3646), .X(n9799) );
  nand_x1_sg U10236 ( .A(\out[1][1][0] ), .B(n10468), .X(n9800) );
  nand_x1_sg U10237 ( .A(n10350), .B(n3647), .X(n9797) );
  nand_x1_sg U10238 ( .A(\out[1][1][1] ), .B(n10299), .X(n9798) );
  nand_x1_sg U10239 ( .A(n10648), .B(n3648), .X(n9795) );
  nand_x1_sg U10240 ( .A(\out[1][1][2] ), .B(n10276), .X(n9796) );
  nand_x1_sg U10241 ( .A(n10374), .B(n3649), .X(n9793) );
  nand_x1_sg U10242 ( .A(\out[1][1][3] ), .B(n10282), .X(n9794) );
  nand_x1_sg U10243 ( .A(n10378), .B(n3652), .X(n9787) );
  nand_x1_sg U10244 ( .A(\out[1][1][6] ), .B(n10461), .X(n9788) );
  nand_x1_sg U10245 ( .A(n10362), .B(n3653), .X(n9785) );
  nand_x1_sg U10246 ( .A(\out[1][1][7] ), .B(n10300), .X(n9786) );
  nand_x1_sg U10247 ( .A(n10342), .B(n3654), .X(n9783) );
  nand_x1_sg U10248 ( .A(\out[1][1][8] ), .B(n10174), .X(n9784) );
  nand_x1_sg U10249 ( .A(n10344), .B(n3655), .X(n9781) );
  nand_x1_sg U10250 ( .A(\out[1][1][9] ), .B(n10518), .X(n9782) );
  nand_x1_sg U10251 ( .A(n10650), .B(n3656), .X(n9779) );
  nand_x1_sg U10252 ( .A(\out[1][1][10] ), .B(n10221), .X(n9780) );
  nand_x1_sg U10253 ( .A(n10669), .B(n3657), .X(n9777) );
  nand_x1_sg U10254 ( .A(\out[1][1][11] ), .B(n10467), .X(n9778) );
  nand_x1_sg U10255 ( .A(n10660), .B(n3658), .X(n9775) );
  nand_x1_sg U10256 ( .A(\out[1][1][12] ), .B(n10514), .X(n9776) );
  nand_x1_sg U10257 ( .A(n10107), .B(n3659), .X(n9773) );
  nand_x1_sg U10258 ( .A(\out[1][1][13] ), .B(n10516), .X(n9774) );
  nand_x1_sg U10259 ( .A(n10657), .B(n3660), .X(n9771) );
  nand_x1_sg U10260 ( .A(\out[1][1][14] ), .B(n10594), .X(n9772) );
  nand_x1_sg U10261 ( .A(n10661), .B(n3661), .X(n9769) );
  nand_x1_sg U10262 ( .A(\out[1][1][15] ), .B(n10296), .X(n9770) );
  nand_x1_sg U10263 ( .A(n10364), .B(n3668), .X(n9755) );
  nand_x1_sg U10264 ( .A(\out[1][2][2] ), .B(n10053), .X(n9756) );
  nand_x1_sg U10265 ( .A(n10642), .B(n3669), .X(n9753) );
  nand_x1_sg U10266 ( .A(\out[1][2][3] ), .B(n10274), .X(n9754) );
  nand_x1_sg U10267 ( .A(n10642), .B(n3670), .X(n9751) );
  nand_x1_sg U10268 ( .A(\out[1][2][4] ), .B(n10509), .X(n9752) );
  nand_x1_sg U10269 ( .A(n10654), .B(n3671), .X(n9749) );
  nand_x1_sg U10270 ( .A(\out[1][2][5] ), .B(n10048), .X(n9750) );
  nand_x1_sg U10271 ( .A(n10346), .B(n3672), .X(n9747) );
  nand_x1_sg U10272 ( .A(\out[1][2][6] ), .B(n10295), .X(n9748) );
  nand_x1_sg U10273 ( .A(n10647), .B(n3673), .X(n9745) );
  nand_x1_sg U10274 ( .A(\out[1][2][7] ), .B(n10051), .X(n9746) );
  nand_x1_sg U10275 ( .A(n10106), .B(n3674), .X(n9743) );
  nand_x1_sg U10276 ( .A(\out[1][2][8] ), .B(n10220), .X(n9744) );
  nand_x1_sg U10277 ( .A(n10364), .B(n3675), .X(n9741) );
  nand_x1_sg U10278 ( .A(\out[1][2][9] ), .B(n10472), .X(n9742) );
  nand_x1_sg U10279 ( .A(n10341), .B(n3676), .X(n9739) );
  nand_x1_sg U10280 ( .A(\out[1][2][10] ), .B(n10165), .X(n9740) );
  nand_x1_sg U10281 ( .A(n10372), .B(n3677), .X(n9737) );
  nand_x1_sg U10282 ( .A(\out[1][2][11] ), .B(n10471), .X(n9738) );
  nand_x1_sg U10283 ( .A(n10669), .B(n3678), .X(n9735) );
  nand_x1_sg U10284 ( .A(\out[1][2][12] ), .B(n10219), .X(n9736) );
  nand_x1_sg U10285 ( .A(n10261), .B(n3679), .X(n9733) );
  nand_x1_sg U10286 ( .A(\out[1][2][13] ), .B(n10464), .X(n9734) );
  nand_x1_sg U10287 ( .A(n10372), .B(n3682), .X(n9727) );
  nand_x1_sg U10288 ( .A(\out[1][2][16] ), .B(n10132), .X(n9728) );
  nand_x1_sg U10289 ( .A(n10672), .B(n3683), .X(n9725) );
  nand_x1_sg U10290 ( .A(\out[1][2][17] ), .B(n10586), .X(n9726) );
  nand_x1_sg U10291 ( .A(n10650), .B(n3684), .X(n9723) );
  nand_x1_sg U10292 ( .A(\out[1][2][18] ), .B(n10464), .X(n9724) );
  nand_x1_sg U10293 ( .A(n10359), .B(n3685), .X(n9721) );
  nand_x1_sg U10294 ( .A(\out[1][2][19] ), .B(n10512), .X(n9722) );
  nand_x1_sg U10295 ( .A(n10350), .B(n3686), .X(n9719) );
  nand_x1_sg U10296 ( .A(\out[1][3][0] ), .B(n10222), .X(n9720) );
  nand_x1_sg U10297 ( .A(n10370), .B(n3687), .X(n9717) );
  nand_x1_sg U10298 ( .A(\out[1][3][1] ), .B(n10507), .X(n9718) );
  nand_x1_sg U10299 ( .A(n10377), .B(n3688), .X(n9715) );
  nand_x1_sg U10300 ( .A(\out[1][3][2] ), .B(n10273), .X(n9716) );
  nand_x1_sg U10301 ( .A(n10314), .B(n3689), .X(n9713) );
  nand_x1_sg U10302 ( .A(\out[1][3][3] ), .B(n10225), .X(n9714) );
  nand_x1_sg U10303 ( .A(n10368), .B(n3690), .X(n9711) );
  nand_x1_sg U10304 ( .A(\out[1][3][4] ), .B(n10506), .X(n9712) );
  nand_x1_sg U10305 ( .A(n10361), .B(n3691), .X(n9709) );
  nand_x1_sg U10306 ( .A(\out[1][3][5] ), .B(n10462), .X(n9710) );
  nand_x1_sg U10307 ( .A(n10666), .B(n3692), .X(n9707) );
  nand_x1_sg U10308 ( .A(\out[1][3][6] ), .B(n10467), .X(n9708) );
  nand_x1_sg U10309 ( .A(n10361), .B(n3693), .X(n9705) );
  nand_x1_sg U10310 ( .A(\out[1][3][7] ), .B(n10272), .X(n9706) );
  nand_x1_sg U10311 ( .A(n10342), .B(n3694), .X(n9703) );
  nand_x1_sg U10312 ( .A(\out[1][3][8] ), .B(n10297), .X(n9704) );
  nand_x1_sg U10313 ( .A(n10366), .B(n3695), .X(n9701) );
  nand_x1_sg U10314 ( .A(\out[1][3][9] ), .B(n10511), .X(n9702) );
  nand_x1_sg U10315 ( .A(n10105), .B(n3696), .X(n9699) );
  nand_x1_sg U10316 ( .A(\out[1][3][10] ), .B(n10520), .X(n9700) );
  nand_x1_sg U10317 ( .A(n10343), .B(n3697), .X(n9697) );
  nand_x1_sg U10318 ( .A(\out[1][3][11] ), .B(n10297), .X(n9698) );
  nand_x1_sg U10319 ( .A(n10667), .B(n3701), .X(n9689) );
  nand_x1_sg U10320 ( .A(\out[1][3][15] ), .B(n10584), .X(n9690) );
  nand_x1_sg U10321 ( .A(n10374), .B(n3706), .X(n9679) );
  nand_x1_sg U10322 ( .A(\out[2][0][0] ), .B(n10220), .X(n9680) );
  nand_x1_sg U10323 ( .A(n10643), .B(n3707), .X(n9677) );
  nand_x1_sg U10324 ( .A(\out[2][0][1] ), .B(n10171), .X(n9678) );
  nand_x1_sg U10325 ( .A(n10383), .B(n3708), .X(n9675) );
  nand_x1_sg U10326 ( .A(\out[2][0][2] ), .B(n10589), .X(n9676) );
  nand_x1_sg U10327 ( .A(n10655), .B(n3709), .X(n9673) );
  nand_x1_sg U10328 ( .A(\out[2][0][3] ), .B(n10051), .X(n9674) );
  nand_x1_sg U10329 ( .A(n10650), .B(n3712), .X(n9667) );
  nand_x1_sg U10330 ( .A(\out[2][0][6] ), .B(n10586), .X(n9668) );
  nand_x1_sg U10331 ( .A(n10649), .B(n3713), .X(n9665) );
  nand_x1_sg U10332 ( .A(\out[2][0][7] ), .B(n10584), .X(n9666) );
  nand_x1_sg U10333 ( .A(n10654), .B(n3714), .X(n9663) );
  nand_x1_sg U10334 ( .A(\out[2][0][8] ), .B(n10296), .X(n9664) );
  nand_x1_sg U10335 ( .A(n10347), .B(n3715), .X(n9661) );
  nand_x1_sg U10336 ( .A(\out[2][0][9] ), .B(n10508), .X(n9662) );
  nand_x1_sg U10337 ( .A(n10660), .B(n3716), .X(n9659) );
  nand_x1_sg U10338 ( .A(\out[2][0][10] ), .B(n10511), .X(n9660) );
  nand_x1_sg U10339 ( .A(n10405), .B(n3717), .X(n9657) );
  nand_x1_sg U10340 ( .A(\out[2][0][11] ), .B(n10170), .X(n9658) );
  nand_x1_sg U10341 ( .A(n10674), .B(n3718), .X(n9655) );
  nand_x1_sg U10342 ( .A(\out[2][0][12] ), .B(n10282), .X(n9656) );
  nand_x1_sg U10343 ( .A(n10646), .B(n3721), .X(n9649) );
  nand_x1_sg U10344 ( .A(\out[2][0][15] ), .B(n10051), .X(n9650) );
  nand_x1_sg U10345 ( .A(n10376), .B(n3722), .X(n9647) );
  nand_x1_sg U10346 ( .A(\out[2][0][16] ), .B(n10281), .X(n9648) );
  nand_x1_sg U10347 ( .A(n10346), .B(n3723), .X(n9645) );
  nand_x1_sg U10348 ( .A(\out[2][0][17] ), .B(n10503), .X(n9646) );
  nand_x1_sg U10349 ( .A(n10380), .B(n3724), .X(n9643) );
  nand_x1_sg U10350 ( .A(\out[2][0][18] ), .B(n10284), .X(n9644) );
  nand_x1_sg U10351 ( .A(n10377), .B(n3725), .X(n9641) );
  nand_x1_sg U10352 ( .A(\out[2][0][19] ), .B(n10503), .X(n9642) );
  nand_x1_sg U10353 ( .A(n10643), .B(n3726), .X(n9639) );
  nand_x1_sg U10354 ( .A(\out[2][1][0] ), .B(n10592), .X(n9640) );
  nand_x1_sg U10355 ( .A(n10359), .B(n3727), .X(n9637) );
  nand_x1_sg U10356 ( .A(\out[2][1][1] ), .B(n10166), .X(n9638) );
  nand_x1_sg U10357 ( .A(n10360), .B(n3731), .X(n9629) );
  nand_x1_sg U10358 ( .A(\out[2][1][5] ), .B(n10284), .X(n9630) );
  nand_x1_sg U10359 ( .A(n10348), .B(n3732), .X(n9627) );
  nand_x1_sg U10360 ( .A(\out[2][1][6] ), .B(n10468), .X(n9628) );
  nand_x1_sg U10361 ( .A(n10354), .B(n3733), .X(n9625) );
  nand_x1_sg U10362 ( .A(\out[2][1][7] ), .B(n10509), .X(n9626) );
  nand_x1_sg U10363 ( .A(n10097), .B(n3734), .X(n9623) );
  nand_x1_sg U10364 ( .A(\out[2][1][8] ), .B(n10586), .X(n9624) );
  nand_x1_sg U10365 ( .A(n10347), .B(n3735), .X(n9621) );
  nand_x1_sg U10366 ( .A(\out[2][1][9] ), .B(n10135), .X(n9622) );
  nand_x1_sg U10367 ( .A(n10359), .B(n3736), .X(n9619) );
  nand_x1_sg U10368 ( .A(\out[2][1][10] ), .B(n10462), .X(n9620) );
  nand_x1_sg U10369 ( .A(n10364), .B(n3737), .X(n9617) );
  nand_x1_sg U10370 ( .A(\out[2][1][11] ), .B(n10161), .X(n9618) );
  nand_x1_sg U10371 ( .A(n10365), .B(n3738), .X(n9615) );
  nand_x1_sg U10372 ( .A(\out[2][1][12] ), .B(n10504), .X(n9616) );
  nand_x1_sg U10373 ( .A(n10262), .B(n3739), .X(n9613) );
  nand_x1_sg U10374 ( .A(\out[2][1][13] ), .B(n10040), .X(n9614) );
  nand_x1_sg U10375 ( .A(n10022), .B(n3741), .X(n9609) );
  nand_x1_sg U10376 ( .A(\out[2][1][15] ), .B(n10271), .X(n9610) );
  nand_x1_sg U10377 ( .A(n10341), .B(n3747), .X(n9597) );
  nand_x1_sg U10378 ( .A(\out[2][2][1] ), .B(n10594), .X(n9598) );
  nand_x1_sg U10379 ( .A(n10404), .B(n3748), .X(n9595) );
  nand_x1_sg U10380 ( .A(\out[2][2][2] ), .B(n10271), .X(n9596) );
  nand_x1_sg U10381 ( .A(n10358), .B(n3749), .X(n9593) );
  nand_x1_sg U10382 ( .A(\out[2][2][3] ), .B(n10171), .X(n9594) );
  nand_x1_sg U10383 ( .A(n10356), .B(n3750), .X(n9591) );
  nand_x1_sg U10384 ( .A(\out[2][2][4] ), .B(n10165), .X(n9592) );
  nand_x1_sg U10385 ( .A(n10348), .B(n3751), .X(n9589) );
  nand_x1_sg U10386 ( .A(\out[2][2][5] ), .B(n10047), .X(n9590) );
  nand_x1_sg U10387 ( .A(n10092), .B(n3752), .X(n9587) );
  nand_x1_sg U10388 ( .A(\out[2][2][6] ), .B(n10052), .X(n9588) );
  nand_x1_sg U10389 ( .A(n10093), .B(n3753), .X(n9585) );
  nand_x1_sg U10390 ( .A(\out[2][2][7] ), .B(n10592), .X(n9586) );
  nand_x1_sg U10391 ( .A(n10672), .B(n3754), .X(n9583) );
  nand_x1_sg U10392 ( .A(\out[2][2][8] ), .B(n10593), .X(n9584) );
  nand_x1_sg U10393 ( .A(n10659), .B(n3755), .X(n9581) );
  nand_x1_sg U10394 ( .A(\out[2][2][9] ), .B(n10161), .X(n9582) );
  nand_x1_sg U10395 ( .A(n10358), .B(n3756), .X(n9579) );
  nand_x1_sg U10396 ( .A(\out[2][2][10] ), .B(n10516), .X(n9580) );
  nand_x1_sg U10397 ( .A(n10366), .B(n3757), .X(n9577) );
  nand_x1_sg U10398 ( .A(\out[2][2][11] ), .B(n10049), .X(n9578) );
  nand_x1_sg U10399 ( .A(n10658), .B(n3761), .X(n9569) );
  nand_x1_sg U10400 ( .A(\out[2][2][15] ), .B(n10225), .X(n9570) );
  nand_x1_sg U10401 ( .A(n10352), .B(n3762), .X(n9567) );
  nand_x1_sg U10402 ( .A(\out[2][2][16] ), .B(n10300), .X(n9568) );
  nand_x1_sg U10403 ( .A(n10022), .B(n3763), .X(n9565) );
  nand_x1_sg U10404 ( .A(\out[2][2][17] ), .B(n10219), .X(n9566) );
  nand_x1_sg U10405 ( .A(n10656), .B(n3764), .X(n9563) );
  nand_x1_sg U10406 ( .A(\out[2][2][18] ), .B(n10049), .X(n9564) );
  nand_x1_sg U10407 ( .A(n10379), .B(n3765), .X(n9561) );
  nand_x1_sg U10408 ( .A(\out[2][2][19] ), .B(n10225), .X(n9562) );
  nand_x1_sg U10409 ( .A(n10358), .B(n3767), .X(n9557) );
  nand_x1_sg U10410 ( .A(\out[2][3][1] ), .B(n10297), .X(n9558) );
  nand_x1_sg U10411 ( .A(n10373), .B(n3768), .X(n9555) );
  nand_x1_sg U10412 ( .A(\out[2][3][2] ), .B(n10594), .X(n9556) );
  nand_x1_sg U10413 ( .A(n10379), .B(n3769), .X(n9553) );
  nand_x1_sg U10414 ( .A(\out[2][3][3] ), .B(n10220), .X(n9554) );
  nand_x1_sg U10415 ( .A(n10654), .B(n3770), .X(n9551) );
  nand_x1_sg U10416 ( .A(\out[2][3][4] ), .B(n10131), .X(n9552) );
  nand_x1_sg U10417 ( .A(n10313), .B(n3771), .X(n9549) );
  nand_x1_sg U10418 ( .A(\out[2][3][5] ), .B(n10514), .X(n9550) );
  nand_x1_sg U10419 ( .A(n10656), .B(n3772), .X(n9547) );
  nand_x1_sg U10420 ( .A(\out[2][3][6] ), .B(n10224), .X(n9548) );
  nand_x1_sg U10421 ( .A(n10667), .B(n3773), .X(n9545) );
  nand_x1_sg U10422 ( .A(\out[2][3][7] ), .B(n10504), .X(n9546) );
  nand_x1_sg U10423 ( .A(n10655), .B(n3774), .X(n9543) );
  nand_x1_sg U10424 ( .A(\out[2][3][8] ), .B(n10513), .X(n9544) );
  nand_x1_sg U10425 ( .A(n10378), .B(n3777), .X(n9537) );
  nand_x1_sg U10426 ( .A(\out[2][3][11] ), .B(n10283), .X(n9538) );
  nand_x1_sg U10427 ( .A(n10656), .B(n3778), .X(n9535) );
  nand_x1_sg U10428 ( .A(\out[2][3][12] ), .B(n10511), .X(n9536) );
  nand_x1_sg U10429 ( .A(n10362), .B(n3779), .X(n9533) );
  nand_x1_sg U10430 ( .A(\out[2][3][13] ), .B(n10509), .X(n9534) );
  nand_x1_sg U10431 ( .A(n10673), .B(n3780), .X(n9531) );
  nand_x1_sg U10432 ( .A(\out[2][3][14] ), .B(n10516), .X(n9532) );
  nand_x1_sg U10433 ( .A(n10376), .B(n3781), .X(n9529) );
  nand_x1_sg U10434 ( .A(\out[2][3][15] ), .B(n10166), .X(n9530) );
  nand_x1_sg U10435 ( .A(n10349), .B(n3786), .X(n9519) );
  nand_x1_sg U10436 ( .A(\out[3][0][0] ), .B(n10272), .X(n9520) );
  nand_x1_sg U10437 ( .A(n10647), .B(n3787), .X(n9517) );
  nand_x1_sg U10438 ( .A(\out[3][0][1] ), .B(n10468), .X(n9518) );
  nand_x1_sg U10439 ( .A(n10660), .B(n3791), .X(n9509) );
  nand_x1_sg U10440 ( .A(\out[3][0][5] ), .B(n10467), .X(n9510) );
  nand_x1_sg U10441 ( .A(n10107), .B(n3792), .X(n9507) );
  nand_x1_sg U10442 ( .A(\out[3][0][6] ), .B(n10585), .X(n9508) );
  nand_x1_sg U10443 ( .A(n10092), .B(n3793), .X(n9505) );
  nand_x1_sg U10444 ( .A(\out[3][0][7] ), .B(n10503), .X(n9506) );
  nand_x1_sg U10445 ( .A(n10360), .B(n3794), .X(n9503) );
  nand_x1_sg U10446 ( .A(\out[3][0][8] ), .B(n10170), .X(n9504) );
  nand_x1_sg U10447 ( .A(n10100), .B(n3795), .X(n9501) );
  nand_x1_sg U10448 ( .A(\out[3][0][9] ), .B(n10294), .X(n9502) );
  nand_x1_sg U10449 ( .A(n10405), .B(n3796), .X(n9499) );
  nand_x1_sg U10450 ( .A(\out[3][0][10] ), .B(n10588), .X(n9500) );
  nand_x1_sg U10451 ( .A(n10643), .B(n3797), .X(n9497) );
  nand_x1_sg U10452 ( .A(\out[3][0][11] ), .B(n10162), .X(n9498) );
  nand_x1_sg U10453 ( .A(n10662), .B(n3798), .X(n9495) );
  nand_x1_sg U10454 ( .A(\out[3][0][12] ), .B(n10520), .X(n9496) );
  nand_x1_sg U10455 ( .A(n10360), .B(n3799), .X(n9493) );
  nand_x1_sg U10456 ( .A(\out[3][0][13] ), .B(n10050), .X(n9494) );
  nand_x1_sg U10457 ( .A(n10261), .B(n3800), .X(n9491) );
  nand_x1_sg U10458 ( .A(\out[3][0][14] ), .B(n10585), .X(n9492) );
  nand_x1_sg U10459 ( .A(n10354), .B(n3801), .X(n9489) );
  nand_x1_sg U10460 ( .A(\out[3][0][15] ), .B(n10275), .X(n9490) );
  nand_x1_sg U10461 ( .A(n10093), .B(n3802), .X(n9487) );
  nand_x1_sg U10462 ( .A(\out[3][0][16] ), .B(n10518), .X(n9488) );
  nand_x1_sg U10463 ( .A(n10106), .B(n3803), .X(n9485) );
  nand_x1_sg U10464 ( .A(\out[3][0][17] ), .B(n10276), .X(n9486) );
  nand_x1_sg U10465 ( .A(n10669), .B(n3804), .X(n9483) );
  nand_x1_sg U10466 ( .A(\out[3][0][18] ), .B(n10300), .X(n9484) );
  nand_x1_sg U10467 ( .A(n10668), .B(n3807), .X(n9477) );
  nand_x1_sg U10468 ( .A(\out[3][1][1] ), .B(n10461), .X(n9478) );
  nand_x1_sg U10469 ( .A(n10662), .B(n3808), .X(n9475) );
  nand_x1_sg U10470 ( .A(\out[3][1][2] ), .B(n10294), .X(n9476) );
  nand_x1_sg U10471 ( .A(n10643), .B(n3809), .X(n9473) );
  nand_x1_sg U10472 ( .A(\out[3][1][3] ), .B(n10469), .X(n9474) );
  nand_x1_sg U10473 ( .A(n10091), .B(n3810), .X(n9471) );
  nand_x1_sg U10474 ( .A(\out[3][1][4] ), .B(n10585), .X(n9472) );
  nand_x1_sg U10475 ( .A(n10346), .B(n3811), .X(n9469) );
  nand_x1_sg U10476 ( .A(\out[3][1][5] ), .B(n10295), .X(n9470) );
  nand_x1_sg U10477 ( .A(n10344), .B(n3812), .X(n9467) );
  nand_x1_sg U10478 ( .A(\out[3][1][6] ), .B(n10588), .X(n9468) );
  nand_x1_sg U10479 ( .A(n10670), .B(n3813), .X(n9465) );
  nand_x1_sg U10480 ( .A(\out[3][1][7] ), .B(n10521), .X(n9466) );
  nand_x1_sg U10481 ( .A(n10674), .B(n3814), .X(n9463) );
  nand_x1_sg U10482 ( .A(\out[3][1][8] ), .B(n10519), .X(n9464) );
  nand_x1_sg U10483 ( .A(n10644), .B(n3815), .X(n9461) );
  nand_x1_sg U10484 ( .A(\out[3][1][9] ), .B(n10508), .X(n9462) );
  nand_x1_sg U10485 ( .A(n10341), .B(n3816), .X(n9459) );
  nand_x1_sg U10486 ( .A(\out[3][1][10] ), .B(n10284), .X(n9460) );
  nand_x1_sg U10487 ( .A(n10666), .B(n3817), .X(n9457) );
  nand_x1_sg U10488 ( .A(\out[3][1][11] ), .B(n10521), .X(n9458) );
  nand_x1_sg U10489 ( .A(n10384), .B(n3818), .X(n9455) );
  nand_x1_sg U10490 ( .A(\out[3][1][12] ), .B(n10463), .X(n9456) );
  nand_x1_sg U10491 ( .A(n10367), .B(n3819), .X(n9453) );
  nand_x1_sg U10492 ( .A(\out[3][1][13] ), .B(n10040), .X(n9454) );
  nand_x1_sg U10493 ( .A(n10371), .B(n3820), .X(n9451) );
  nand_x1_sg U10494 ( .A(\out[3][1][14] ), .B(n10513), .X(n9452) );
  nand_x1_sg U10495 ( .A(n10368), .B(n3821), .X(n9449) );
  nand_x1_sg U10496 ( .A(\out[3][1][15] ), .B(n10466), .X(n9450) );
  nand_x1_sg U10497 ( .A(n10097), .B(n3826), .X(n9439) );
  nand_x1_sg U10498 ( .A(\out[3][2][0] ), .B(n10299), .X(n9440) );
  nand_x1_sg U10499 ( .A(n10261), .B(n3827), .X(n9437) );
  nand_x1_sg U10500 ( .A(\out[3][2][1] ), .B(n10462), .X(n9438) );
  nand_x1_sg U10501 ( .A(n10350), .B(n3828), .X(n9435) );
  nand_x1_sg U10502 ( .A(\out[3][2][2] ), .B(n10038), .X(n9436) );
  nand_x1_sg U10503 ( .A(n10373), .B(n3829), .X(n9433) );
  nand_x1_sg U10504 ( .A(\out[3][2][3] ), .B(n10514), .X(n9434) );
  nand_x1_sg U10505 ( .A(n10671), .B(n3830), .X(n9431) );
  nand_x1_sg U10506 ( .A(\out[3][2][4] ), .B(n10510), .X(n9432) );
  nand_x1_sg U10507 ( .A(n10669), .B(n3831), .X(n9429) );
  nand_x1_sg U10508 ( .A(\out[3][2][5] ), .B(n10513), .X(n9430) );
  nand_x1_sg U10509 ( .A(n10673), .B(n3832), .X(n9427) );
  nand_x1_sg U10510 ( .A(\out[3][2][6] ), .B(n10272), .X(n9428) );
  nand_x1_sg U10511 ( .A(n10383), .B(n3833), .X(n9425) );
  nand_x1_sg U10512 ( .A(\out[3][2][7] ), .B(n10510), .X(n9426) );
  nand_x1_sg U10513 ( .A(n10347), .B(n3834), .X(n9423) );
  nand_x1_sg U10514 ( .A(\out[3][2][8] ), .B(n10281), .X(n9424) );
  nand_x1_sg U10515 ( .A(n10094), .B(n3837), .X(n9417) );
  nand_x1_sg U10516 ( .A(\out[3][2][11] ), .B(n10512), .X(n9418) );
  nand_x1_sg U10517 ( .A(n10384), .B(n3838), .X(n9415) );
  nand_x1_sg U10518 ( .A(\out[3][2][12] ), .B(n10467), .X(n9416) );
  nand_x1_sg U10519 ( .A(n10371), .B(n3839), .X(n9413) );
  nand_x1_sg U10520 ( .A(\out[3][2][13] ), .B(n10593), .X(n9414) );
  nand_x1_sg U10521 ( .A(n10656), .B(n3840), .X(n9411) );
  nand_x1_sg U10522 ( .A(\out[3][2][14] ), .B(n10519), .X(n9412) );
  nand_x1_sg U10523 ( .A(n10106), .B(n3841), .X(n9409) );
  nand_x1_sg U10524 ( .A(\out[3][2][15] ), .B(n10162), .X(n9410) );
  nand_x1_sg U10525 ( .A(n10642), .B(n3842), .X(n9407) );
  nand_x1_sg U10526 ( .A(\out[3][2][16] ), .B(n10514), .X(n9408) );
  nand_x1_sg U10527 ( .A(n10356), .B(n3843), .X(n9405) );
  nand_x1_sg U10528 ( .A(\out[3][2][17] ), .B(n10589), .X(n9406) );
  nand_x1_sg U10529 ( .A(n10105), .B(n3844), .X(n9403) );
  nand_x1_sg U10530 ( .A(\out[3][2][18] ), .B(n10132), .X(n9404) );
  nand_x1_sg U10531 ( .A(n10261), .B(n3845), .X(n9401) );
  nand_x1_sg U10532 ( .A(\out[3][2][19] ), .B(n10589), .X(n9402) );
  nand_x1_sg U10533 ( .A(n10383), .B(n3846), .X(n9399) );
  nand_x1_sg U10534 ( .A(\out[3][3][0] ), .B(n10293), .X(n9400) );
  nand_x1_sg U10535 ( .A(n10382), .B(n3847), .X(n9397) );
  nand_x1_sg U10536 ( .A(\out[3][3][1] ), .B(n10461), .X(n9398) );
  nand_x1_sg U10537 ( .A(n10314), .B(n3848), .X(n9395) );
  nand_x1_sg U10538 ( .A(\out[3][3][2] ), .B(n10509), .X(n9396) );
  nand_x1_sg U10539 ( .A(n10404), .B(n3849), .X(n9393) );
  nand_x1_sg U10540 ( .A(\out[3][3][3] ), .B(n10136), .X(n9394) );
  nand_x1_sg U10541 ( .A(n10658), .B(n3850), .X(n9391) );
  nand_x1_sg U10542 ( .A(\out[3][3][4] ), .B(n10470), .X(n9392) );
  nand_x1_sg U10543 ( .A(n10367), .B(n3851), .X(n9389) );
  nand_x1_sg U10544 ( .A(\out[3][3][5] ), .B(n10466), .X(n9390) );
  nand_x1_sg U10545 ( .A(n10093), .B(n3852), .X(n9387) );
  nand_x1_sg U10546 ( .A(\out[3][3][6] ), .B(n10136), .X(n9388) );
  nand_x1_sg U10547 ( .A(\out[3][3][10] ), .B(n10221), .X(n9380) );
  nand_x1_sg U10548 ( .A(n10364), .B(n3857), .X(n9377) );
  nand_x1_sg U10549 ( .A(\out[3][3][11] ), .B(n10224), .X(n9378) );
  nand_x1_sg U10550 ( .A(n10104), .B(n3858), .X(n9375) );
  nand_x1_sg U10551 ( .A(\out[3][3][12] ), .B(n10275), .X(n9376) );
  nand_x1_sg U10552 ( .A(n10405), .B(n3859), .X(n9373) );
  nand_x1_sg U10553 ( .A(\out[3][3][13] ), .B(n10518), .X(n9374) );
  nand_x1_sg U10554 ( .A(n10648), .B(n3860), .X(n9371) );
  nand_x1_sg U10555 ( .A(\out[3][3][14] ), .B(n10132), .X(n9372) );
  nand_x1_sg U10556 ( .A(n10406), .B(n3861), .X(n9369) );
  nand_x1_sg U10557 ( .A(\out[3][3][15] ), .B(n10503), .X(n9370) );
  nand_x1_sg U10558 ( .A(n10373), .B(n3555), .X(n9981) );
  nand_x1_sg U10559 ( .A(\out[0][0][9] ), .B(n10219), .X(n9982) );
  nand_x1_sg U10560 ( .A(n10672), .B(n3556), .X(n9979) );
  nand_x1_sg U10561 ( .A(\out[0][0][10] ), .B(n10040), .X(n9980) );
  nand_x1_sg U10562 ( .A(n10262), .B(n3569), .X(n9953) );
  nand_x1_sg U10563 ( .A(\out[0][1][3] ), .B(n10223), .X(n9954) );
  nand_x1_sg U10564 ( .A(n10108), .B(n3586), .X(n9919) );
  nand_x1_sg U10565 ( .A(\out[0][2][0] ), .B(n10222), .X(n9920) );
  nand_x1_sg U10566 ( .A(n10661), .B(n3615), .X(n9861) );
  nand_x1_sg U10567 ( .A(\out[0][3][9] ), .B(n10465), .X(n9862) );
  nand_x1_sg U10568 ( .A(n10660), .B(n3621), .X(n9849) );
  nand_x1_sg U10569 ( .A(\out[0][3][15] ), .B(n10510), .X(n9850) );
  nand_x1_sg U10570 ( .A(n10382), .B(n3650), .X(n9791) );
  nand_x1_sg U10571 ( .A(\out[1][1][4] ), .B(n10295), .X(n9792) );
  nand_x1_sg U10572 ( .A(n10657), .B(n3651), .X(n9789) );
  nand_x1_sg U10573 ( .A(\out[1][1][5] ), .B(n10472), .X(n9790) );
  nand_x1_sg U10574 ( .A(n10404), .B(n3680), .X(n9731) );
  nand_x1_sg U10575 ( .A(\out[1][2][14] ), .B(n10271), .X(n9732) );
  nand_x1_sg U10576 ( .A(n10380), .B(n3681), .X(n9729) );
  nand_x1_sg U10577 ( .A(\out[1][2][15] ), .B(n10224), .X(n9730) );
  nand_x1_sg U10578 ( .A(n10348), .B(n3710), .X(n9671) );
  nand_x1_sg U10579 ( .A(\out[2][0][4] ), .B(n10516), .X(n9672) );
  nand_x1_sg U10580 ( .A(n10671), .B(n3711), .X(n9669) );
  nand_x1_sg U10581 ( .A(\out[2][0][5] ), .B(n10298), .X(n9670) );
  nand_x1_sg U10582 ( .A(n10344), .B(n3740), .X(n9611) );
  nand_x1_sg U10583 ( .A(\out[2][1][14] ), .B(n10520), .X(n9612) );
  nand_x1_sg U10584 ( .A(n10355), .B(n3746), .X(n9599) );
  nand_x1_sg U10585 ( .A(\out[2][2][0] ), .B(n10519), .X(n9600) );
  nand_x1_sg U10586 ( .A(n10648), .B(n3766), .X(n9559) );
  nand_x1_sg U10587 ( .A(\out[2][3][0] ), .B(n10223), .X(n9560) );
  nand_x1_sg U10588 ( .A(n10359), .B(n3775), .X(n9541) );
  nand_x1_sg U10589 ( .A(\out[2][3][9] ), .B(n10283), .X(n9542) );
  nand_x1_sg U10590 ( .A(n10354), .B(n3776), .X(n9539) );
  nand_x1_sg U10591 ( .A(\out[2][3][10] ), .B(n10274), .X(n9540) );
  nand_x1_sg U10592 ( .A(n10406), .B(n3805), .X(n9481) );
  nand_x1_sg U10593 ( .A(\out[3][0][19] ), .B(n10592), .X(n9482) );
  nand_x1_sg U10594 ( .A(n10262), .B(n3806), .X(n9479) );
  nand_x1_sg U10595 ( .A(\out[3][1][0] ), .B(n10518), .X(n9480) );
  nand_x1_sg U10596 ( .A(n10343), .B(n3835), .X(n9421) );
  nand_x1_sg U10597 ( .A(\out[3][2][9] ), .B(n10136), .X(n9422) );
  nand_x1_sg U10598 ( .A(n10374), .B(n3836), .X(n9419) );
  nand_x1_sg U10599 ( .A(\out[3][2][10] ), .B(n10512), .X(n9420) );
  nand_x1_sg U10600 ( .A(n10382), .B(n3663), .X(n9765) );
  nand_x1_sg U10601 ( .A(\out[1][1][17] ), .B(n10173), .X(n9766) );
  nand_x1_sg U10602 ( .A(n10668), .B(n3664), .X(n9763) );
  nand_x1_sg U10603 ( .A(\out[1][1][18] ), .B(n10505), .X(n9764) );
  nand_x1_sg U10604 ( .A(n10406), .B(n3665), .X(n9761) );
  nand_x1_sg U10605 ( .A(\out[1][1][19] ), .B(n10512), .X(n9762) );
  nand_x1_sg U10606 ( .A(n10654), .B(n3744), .X(n9603) );
  nand_x1_sg U10607 ( .A(\out[2][1][18] ), .B(n10506), .X(n9604) );
  nand_x1_sg U10608 ( .A(n10091), .B(n3823), .X(n9445) );
  nand_x1_sg U10609 ( .A(\out[3][1][17] ), .B(n10272), .X(n9446) );
  nand_x1_sg U10610 ( .A(n10341), .B(n3824), .X(n9443) );
  nand_x1_sg U10611 ( .A(\out[3][1][18] ), .B(n10053), .X(n9444) );
  nand_x1_sg U10612 ( .A(n10349), .B(n3825), .X(n9441) );
  nand_x1_sg U10613 ( .A(\out[3][1][19] ), .B(n10464), .X(n9442) );
  nand_x1_sg U10614 ( .A(n10097), .B(n3582), .X(n9927) );
  nand_x1_sg U10615 ( .A(\out[0][1][16] ), .B(n10505), .X(n9928) );
  nand_x1_sg U10616 ( .A(n10649), .B(n3583), .X(n9925) );
  nand_x1_sg U10617 ( .A(\out[0][1][17] ), .B(n10174), .X(n9926) );
  nand_x1_sg U10618 ( .A(n10647), .B(n3584), .X(n9923) );
  nand_x1_sg U10619 ( .A(\out[0][1][18] ), .B(n10508), .X(n9924) );
  nand_x1_sg U10620 ( .A(n10366), .B(n3622), .X(n9847) );
  nand_x1_sg U10621 ( .A(\out[0][3][16] ), .B(n10222), .X(n9848) );
  nand_x1_sg U10622 ( .A(n10362), .B(n3623), .X(n9845) );
  nand_x1_sg U10623 ( .A(\out[0][3][17] ), .B(n10470), .X(n9846) );
  nand_x1_sg U10624 ( .A(n10100), .B(n3624), .X(n9843) );
  nand_x1_sg U10625 ( .A(\out[0][3][18] ), .B(n10221), .X(n9844) );
  nand_x1_sg U10626 ( .A(n10372), .B(n3625), .X(n9841) );
  nand_x1_sg U10627 ( .A(\out[0][3][19] ), .B(n10174), .X(n9842) );
  nand_x1_sg U10628 ( .A(n10091), .B(n3662), .X(n9767) );
  nand_x1_sg U10629 ( .A(\out[1][1][16] ), .B(n10300), .X(n9768) );
  nand_x1_sg U10630 ( .A(n10106), .B(n3702), .X(n9687) );
  nand_x1_sg U10631 ( .A(\out[1][3][16] ), .B(n10171), .X(n9688) );
  nand_x1_sg U10632 ( .A(n10358), .B(n3703), .X(n9685) );
  nand_x1_sg U10633 ( .A(\out[1][3][17] ), .B(n10590), .X(n9686) );
  nand_x1_sg U10634 ( .A(n10343), .B(n3704), .X(n9683) );
  nand_x1_sg U10635 ( .A(\out[1][3][18] ), .B(n10519), .X(n9684) );
  nand_x1_sg U10636 ( .A(n10344), .B(n3705), .X(n9681) );
  nand_x1_sg U10637 ( .A(\out[1][3][19] ), .B(n10283), .X(n9682) );
  nand_x1_sg U10638 ( .A(n10366), .B(n3742), .X(n9607) );
  nand_x1_sg U10639 ( .A(\out[2][1][16] ), .B(n10135), .X(n9608) );
  nand_x1_sg U10640 ( .A(n10380), .B(n3745), .X(n9601) );
  nand_x1_sg U10641 ( .A(\out[2][1][19] ), .B(n10274), .X(n9602) );
  nand_x1_sg U10642 ( .A(n10673), .B(n3782), .X(n9527) );
  nand_x1_sg U10643 ( .A(\out[2][3][16] ), .B(n10293), .X(n9528) );
  nand_x1_sg U10644 ( .A(n10659), .B(n3783), .X(n9525) );
  nand_x1_sg U10645 ( .A(\out[2][3][17] ), .B(n10048), .X(n9526) );
  nand_x1_sg U10646 ( .A(n10347), .B(n3784), .X(n9523) );
  nand_x1_sg U10647 ( .A(\out[2][3][18] ), .B(n10162), .X(n9524) );
  nand_x1_sg U10648 ( .A(n10097), .B(n3785), .X(n9521) );
  nand_x1_sg U10649 ( .A(\out[2][3][19] ), .B(n10173), .X(n9522) );
  nand_x1_sg U10650 ( .A(n10670), .B(n3822), .X(n9447) );
  nand_x1_sg U10651 ( .A(\out[3][1][16] ), .B(n10471), .X(n9448) );
  nand_x1_sg U10652 ( .A(n10367), .B(n3862), .X(n9367) );
  nand_x1_sg U10653 ( .A(\out[3][3][16] ), .B(n10283), .X(n9368) );
  nand_x1_sg U10654 ( .A(n10350), .B(n3863), .X(n9365) );
  nand_x1_sg U10655 ( .A(\out[3][3][17] ), .B(n10461), .X(n9366) );
  nand_x1_sg U10656 ( .A(n10089), .B(n3864), .X(n9363) );
  nand_x1_sg U10657 ( .A(\out[3][3][18] ), .B(n10511), .X(n9364) );
  nand_x1_sg U10658 ( .A(n10343), .B(n3585), .X(n9921) );
  nand_x1_sg U10659 ( .A(\out[0][1][19] ), .B(n10505), .X(n9922) );
  nand_x1_sg U10660 ( .A(n10645), .B(n3743), .X(n9605) );
  nand_x1_sg U10661 ( .A(\out[2][1][17] ), .B(n10165), .X(n9606) );
  nand_x1_sg U10662 ( .A(n10349), .B(n3865), .X(n9360) );
  nand_x1_sg U10663 ( .A(\out[3][3][19] ), .B(n10296), .X(n9361) );
  inv_x1_sg U10664 ( .A(state[0]), .X(n12286) );
  nor_x1_sg U10665 ( .A(n12287), .B(n10002), .X(n10001) );
  nand_x1_sg U10666 ( .A(output_taken), .B(n12286), .X(n10002) );
  inv_x1_sg U10667 ( .A(state[1]), .X(n12287) );
  nand_x1_sg U10668 ( .A(n8711), .B(state[0]), .X(n8707) );
  nor_x1_sg U10669 ( .A(n8711), .B(n10677), .X(n8709) );
  nand_x1_sg U10670 ( .A(n8711), .B(state[1]), .X(n8713) );
  nand_x1_sg U10671 ( .A(\in[0][0][0] ), .B(n10632), .X(n9357) );
  nand_x1_sg U10672 ( .A(\reg_in[0][0][0] ), .B(n10534), .X(n9358) );
  nand_x1_sg U10673 ( .A(\in[0][0][1] ), .B(n10333), .X(n9355) );
  nand_x1_sg U10674 ( .A(\reg_in[0][0][1] ), .B(n10481), .X(n9356) );
  nand_x1_sg U10675 ( .A(\in[0][0][2] ), .B(n10023), .X(n9353) );
  nand_x1_sg U10676 ( .A(\reg_in[0][0][2] ), .B(n10473), .X(n9354) );
  nand_x1_sg U10677 ( .A(\in[0][0][3] ), .B(n10327), .X(n9351) );
  nand_x1_sg U10678 ( .A(\reg_in[0][0][3] ), .B(n10184), .X(n9352) );
  nand_x1_sg U10679 ( .A(\in[0][0][4] ), .B(n10329), .X(n9349) );
  nand_x1_sg U10680 ( .A(\reg_in[0][0][4] ), .B(n10304), .X(n9350) );
  nand_x1_sg U10681 ( .A(\in[0][0][5] ), .B(n10333), .X(n9347) );
  nand_x1_sg U10682 ( .A(\reg_in[0][0][5] ), .B(n10215), .X(n9348) );
  nand_x1_sg U10683 ( .A(\in[0][0][6] ), .B(n10632), .X(n9345) );
  nand_x1_sg U10684 ( .A(\reg_in[0][0][6] ), .B(n10286), .X(n9346) );
  nand_x1_sg U10685 ( .A(\in[0][0][7] ), .B(n10398), .X(n9343) );
  nand_x1_sg U10686 ( .A(\reg_in[0][0][7] ), .B(n10189), .X(n9344) );
  nand_x1_sg U10687 ( .A(\in[0][0][8] ), .B(n10084), .X(n9341) );
  nand_x1_sg U10688 ( .A(\reg_in[0][0][8] ), .B(n10476), .X(n9342) );
  nand_x1_sg U10689 ( .A(\in[0][0][9] ), .B(n10083), .X(n9339) );
  nand_x1_sg U10690 ( .A(\reg_in[0][0][9] ), .B(n10054), .X(n9340) );
  nand_x1_sg U10691 ( .A(\in[0][0][10] ), .B(n10612), .X(n9337) );
  nand_x1_sg U10692 ( .A(\reg_in[0][0][10] ), .B(n10216), .X(n9338) );
  nand_x1_sg U10693 ( .A(\in[0][0][11] ), .B(n10388), .X(n9335) );
  nand_x1_sg U10694 ( .A(\reg_in[0][0][11] ), .B(n10055), .X(n9336) );
  nand_x1_sg U10695 ( .A(\in[0][0][12] ), .B(n10333), .X(n9333) );
  nand_x1_sg U10696 ( .A(\reg_in[0][0][12] ), .B(n10301), .X(n9334) );
  nand_x1_sg U10697 ( .A(\in[0][0][13] ), .B(n10620), .X(n9331) );
  nand_x1_sg U10698 ( .A(\reg_in[0][0][13] ), .B(n10145), .X(n9332) );
  nand_x1_sg U10699 ( .A(\in[0][0][14] ), .B(n10340), .X(n9329) );
  nand_x1_sg U10700 ( .A(\reg_in[0][0][14] ), .B(n10575), .X(n9330) );
  nand_x1_sg U10701 ( .A(\in[0][0][15] ), .B(n10326), .X(n9327) );
  nand_x1_sg U10702 ( .A(\reg_in[0][0][15] ), .B(n10212), .X(n9328) );
  nand_x1_sg U10703 ( .A(\in[0][0][16] ), .B(n10329), .X(n9325) );
  nand_x1_sg U10704 ( .A(\reg_in[0][0][16] ), .B(n10305), .X(n9326) );
  nand_x1_sg U10705 ( .A(\in[0][0][17] ), .B(n10607), .X(n9323) );
  nand_x1_sg U10706 ( .A(\reg_in[0][0][17] ), .B(n10141), .X(n9324) );
  nand_x1_sg U10707 ( .A(\in[0][0][18] ), .B(n10614), .X(n9321) );
  nand_x1_sg U10708 ( .A(\reg_in[0][0][18] ), .B(n10191), .X(n9322) );
  nand_x1_sg U10709 ( .A(\in[0][0][19] ), .B(n10324), .X(n9319) );
  nand_x1_sg U10710 ( .A(\reg_in[0][0][19] ), .B(n10270), .X(n9320) );
  nand_x1_sg U10711 ( .A(\in[0][1][0] ), .B(n10625), .X(n9317) );
  nand_x1_sg U10712 ( .A(\reg_in[0][1][0] ), .B(n10530), .X(n9318) );
  nand_x1_sg U10713 ( .A(\in[0][1][1] ), .B(n10607), .X(n9315) );
  nand_x1_sg U10714 ( .A(\reg_in[0][1][1] ), .B(n10266), .X(n9316) );
  nand_x1_sg U10715 ( .A(\in[0][1][2] ), .B(n10395), .X(n9313) );
  nand_x1_sg U10716 ( .A(\reg_in[0][1][2] ), .B(n10574), .X(n9314) );
  nand_x1_sg U10717 ( .A(\in[0][1][3] ), .B(n10340), .X(n9311) );
  nand_x1_sg U10718 ( .A(\reg_in[0][1][3] ), .B(n10287), .X(n9312) );
  nand_x1_sg U10719 ( .A(\in[0][1][4] ), .B(n10411), .X(n9309) );
  nand_x1_sg U10720 ( .A(\reg_in[0][1][4] ), .B(n10269), .X(n9310) );
  nand_x1_sg U10721 ( .A(\in[0][1][10] ), .B(n10330), .X(n9297) );
  nand_x1_sg U10722 ( .A(\reg_in[0][1][10] ), .B(n10301), .X(n9298) );
  nand_x1_sg U10723 ( .A(\in[0][1][11] ), .B(n10409), .X(n9295) );
  nand_x1_sg U10724 ( .A(\reg_in[0][1][11] ), .B(n10580), .X(n9296) );
  nand_x1_sg U10725 ( .A(\in[0][1][12] ), .B(n10399), .X(n9293) );
  nand_x1_sg U10726 ( .A(\reg_in[0][1][12] ), .B(n10526), .X(n9294) );
  nand_x1_sg U10727 ( .A(\in[0][1][13] ), .B(n10398), .X(n9291) );
  nand_x1_sg U10728 ( .A(\reg_in[0][1][13] ), .B(n10268), .X(n9292) );
  nand_x1_sg U10729 ( .A(\in[0][1][14] ), .B(n10318), .X(n9289) );
  nand_x1_sg U10730 ( .A(\reg_in[0][1][14] ), .B(n10140), .X(n9290) );
  nand_x1_sg U10731 ( .A(\in[0][1][15] ), .B(n10021), .X(n9287) );
  nand_x1_sg U10732 ( .A(\reg_in[0][1][15] ), .B(n10059), .X(n9288) );
  nand_x1_sg U10733 ( .A(\in[0][1][16] ), .B(n10624), .X(n9285) );
  nand_x1_sg U10734 ( .A(\reg_in[0][1][16] ), .B(n10531), .X(n9286) );
  nand_x1_sg U10735 ( .A(\in[0][1][17] ), .B(n10626), .X(n9283) );
  nand_x1_sg U10736 ( .A(\reg_in[0][1][17] ), .B(n10306), .X(n9284) );
  nand_x1_sg U10737 ( .A(\in[0][1][18] ), .B(n10617), .X(n9281) );
  nand_x1_sg U10738 ( .A(\reg_in[0][1][18] ), .B(n10575), .X(n9282) );
  nand_x1_sg U10739 ( .A(\in[0][1][19] ), .B(n10335), .X(n9279) );
  nand_x1_sg U10740 ( .A(\reg_in[0][1][19] ), .B(n10212), .X(n9280) );
  nand_x1_sg U10741 ( .A(\in[0][2][0] ), .B(n10080), .X(n9277) );
  nand_x1_sg U10742 ( .A(\reg_in[0][2][0] ), .B(n10528), .X(n9278) );
  nand_x1_sg U10743 ( .A(\in[0][2][1] ), .B(n10409), .X(n9275) );
  nand_x1_sg U10744 ( .A(\reg_in[0][2][1] ), .B(n10304), .X(n9276) );
  nand_x1_sg U10745 ( .A(\in[0][2][2] ), .B(n10620), .X(n9273) );
  nand_x1_sg U10746 ( .A(\reg_in[0][2][2] ), .B(n10217), .X(n9274) );
  nand_x1_sg U10747 ( .A(\in[0][2][3] ), .B(n10401), .X(n9271) );
  nand_x1_sg U10748 ( .A(\reg_in[0][2][3] ), .B(n10268), .X(n9272) );
  nand_x1_sg U10749 ( .A(\in[0][2][4] ), .B(n10329), .X(n9269) );
  nand_x1_sg U10750 ( .A(\reg_in[0][2][4] ), .B(n10484), .X(n9270) );
  nand_x1_sg U10751 ( .A(\in[0][2][5] ), .B(n10395), .X(n9267) );
  nand_x1_sg U10752 ( .A(\reg_in[0][2][5] ), .B(n10211), .X(n9268) );
  nand_x1_sg U10753 ( .A(\in[0][2][6] ), .B(n10629), .X(n9265) );
  nand_x1_sg U10754 ( .A(\reg_in[0][2][6] ), .B(n10526), .X(n9266) );
  nand_x1_sg U10755 ( .A(\in[0][2][7] ), .B(n10077), .X(n9263) );
  nand_x1_sg U10756 ( .A(\reg_in[0][2][7] ), .B(n10541), .X(n9264) );
  nand_x1_sg U10757 ( .A(\in[0][2][8] ), .B(n10618), .X(n9261) );
  nand_x1_sg U10758 ( .A(\reg_in[0][2][8] ), .B(n10307), .X(n9262) );
  nand_x1_sg U10759 ( .A(\in[0][2][9] ), .B(n10396), .X(n9259) );
  nand_x1_sg U10760 ( .A(\reg_in[0][2][9] ), .B(n10285), .X(n9260) );
  nand_x1_sg U10761 ( .A(\in[0][2][10] ), .B(n10399), .X(n9257) );
  nand_x1_sg U10762 ( .A(\reg_in[0][2][10] ), .B(n10305), .X(n9258) );
  nand_x1_sg U10763 ( .A(\in[0][2][11] ), .B(n10409), .X(n9255) );
  nand_x1_sg U10764 ( .A(\reg_in[0][2][11] ), .B(n10529), .X(n9256) );
  nand_x1_sg U10765 ( .A(\in[0][2][12] ), .B(n10333), .X(n9253) );
  nand_x1_sg U10766 ( .A(\reg_in[0][2][12] ), .B(n10145), .X(n9254) );
  nand_x1_sg U10767 ( .A(\in[0][2][13] ), .B(n10332), .X(n9251) );
  nand_x1_sg U10768 ( .A(\reg_in[0][2][13] ), .B(n10477), .X(n9252) );
  nand_x1_sg U10769 ( .A(\in[0][2][14] ), .B(n10400), .X(n9249) );
  nand_x1_sg U10770 ( .A(\reg_in[0][2][14] ), .B(n10041), .X(n9250) );
  nand_x1_sg U10771 ( .A(\in[0][3][0] ), .B(n10073), .X(n9237) );
  nand_x1_sg U10772 ( .A(\reg_in[0][3][0] ), .B(n10527), .X(n9238) );
  nand_x1_sg U10773 ( .A(\in[0][3][1] ), .B(n10603), .X(n9235) );
  nand_x1_sg U10774 ( .A(\reg_in[0][3][1] ), .B(n10215), .X(n9236) );
  nand_x1_sg U10775 ( .A(\in[0][3][2] ), .B(n10392), .X(n9233) );
  nand_x1_sg U10776 ( .A(\reg_in[0][3][2] ), .B(n10183), .X(n9234) );
  nand_x1_sg U10777 ( .A(\in[0][3][3] ), .B(n10258), .X(n9231) );
  nand_x1_sg U10778 ( .A(\reg_in[0][3][3] ), .B(n10054), .X(n9232) );
  nand_x1_sg U10779 ( .A(\in[0][3][4] ), .B(n10617), .X(n9229) );
  nand_x1_sg U10780 ( .A(\reg_in[0][3][4] ), .B(n10055), .X(n9230) );
  nand_x1_sg U10781 ( .A(\in[0][3][5] ), .B(n10075), .X(n9227) );
  nand_x1_sg U10782 ( .A(\reg_in[0][3][5] ), .B(n10535), .X(n9228) );
  nand_x1_sg U10783 ( .A(\in[0][3][6] ), .B(n10400), .X(n9225) );
  nand_x1_sg U10784 ( .A(\reg_in[0][3][6] ), .B(n10529), .X(n9226) );
  nand_x1_sg U10785 ( .A(\in[0][3][7] ), .B(n10075), .X(n9223) );
  nand_x1_sg U10786 ( .A(\reg_in[0][3][7] ), .B(n10179), .X(n9224) );
  nand_x1_sg U10787 ( .A(\in[0][3][8] ), .B(n10074), .X(n9221) );
  nand_x1_sg U10788 ( .A(\reg_in[0][3][8] ), .B(n10575), .X(n9222) );
  nand_x1_sg U10789 ( .A(\in[0][3][9] ), .B(n10614), .X(n9219) );
  nand_x1_sg U10790 ( .A(\reg_in[0][3][9] ), .B(n10285), .X(n9220) );
  nand_x1_sg U10791 ( .A(\in[0][3][15] ), .B(n10386), .X(n9207) );
  nand_x1_sg U10792 ( .A(\reg_in[0][3][15] ), .B(n10057), .X(n9208) );
  nand_x1_sg U10793 ( .A(\in[0][3][16] ), .B(n10081), .X(n9205) );
  nand_x1_sg U10794 ( .A(\reg_in[0][3][16] ), .B(n10183), .X(n9206) );
  nand_x1_sg U10795 ( .A(\in[0][3][17] ), .B(n10324), .X(n9203) );
  nand_x1_sg U10796 ( .A(\reg_in[0][3][17] ), .B(n10266), .X(n9204) );
  nand_x1_sg U10797 ( .A(\in[0][3][18] ), .B(n10401), .X(n9201) );
  nand_x1_sg U10798 ( .A(\reg_in[0][3][18] ), .B(n10269), .X(n9202) );
  nand_x1_sg U10799 ( .A(\in[0][3][19] ), .B(n10318), .X(n9199) );
  nand_x1_sg U10800 ( .A(\reg_in[0][3][19] ), .B(n10287), .X(n9200) );
  nand_x1_sg U10801 ( .A(\in[1][0][0] ), .B(n10605), .X(n9197) );
  nand_x1_sg U10802 ( .A(\reg_in[1][0][0] ), .B(n10191), .X(n9198) );
  nand_x1_sg U10803 ( .A(\in[1][0][1] ), .B(n10411), .X(n9195) );
  nand_x1_sg U10804 ( .A(\reg_in[1][0][1] ), .B(n10526), .X(n9196) );
  nand_x1_sg U10805 ( .A(\in[1][0][2] ), .B(n10075), .X(n9193) );
  nand_x1_sg U10806 ( .A(\reg_in[1][0][2] ), .B(n10527), .X(n9194) );
  nand_x1_sg U10807 ( .A(\in[1][0][3] ), .B(n10618), .X(n9191) );
  nand_x1_sg U10808 ( .A(\reg_in[1][0][3] ), .B(n10572), .X(n9192) );
  nand_x1_sg U10809 ( .A(\in[1][0][4] ), .B(n10615), .X(n9189) );
  nand_x1_sg U10810 ( .A(\reg_in[1][0][4] ), .B(n10303), .X(n9190) );
  nand_x1_sg U10811 ( .A(\in[1][0][10] ), .B(n10316), .X(n9177) );
  nand_x1_sg U10812 ( .A(\reg_in[1][0][10] ), .B(n10578), .X(n9178) );
  nand_x1_sg U10813 ( .A(\in[1][0][11] ), .B(n10338), .X(n9175) );
  nand_x1_sg U10814 ( .A(\reg_in[1][0][11] ), .B(n10483), .X(n9176) );
  nand_x1_sg U10815 ( .A(\in[1][0][12] ), .B(n10393), .X(n9173) );
  nand_x1_sg U10816 ( .A(\reg_in[1][0][12] ), .B(n10578), .X(n9174) );
  nand_x1_sg U10817 ( .A(\in[1][0][13] ), .B(n10619), .X(n9171) );
  nand_x1_sg U10818 ( .A(\reg_in[1][0][13] ), .B(n10523), .X(n9172) );
  nand_x1_sg U10819 ( .A(\in[1][0][14] ), .B(n10603), .X(n9169) );
  nand_x1_sg U10820 ( .A(\reg_in[1][0][14] ), .B(n10211), .X(n9170) );
  nand_x1_sg U10821 ( .A(\in[1][0][15] ), .B(n10259), .X(n9167) );
  nand_x1_sg U10822 ( .A(\reg_in[1][0][15] ), .B(n10481), .X(n9168) );
  nand_x1_sg U10823 ( .A(\in[1][0][16] ), .B(n10335), .X(n9165) );
  nand_x1_sg U10824 ( .A(\reg_in[1][0][16] ), .B(n10524), .X(n9166) );
  nand_x1_sg U10825 ( .A(\in[1][0][17] ), .B(n10387), .X(n9163) );
  nand_x1_sg U10826 ( .A(\reg_in[1][0][17] ), .B(n10540), .X(n9164) );
  nand_x1_sg U10827 ( .A(\in[1][0][18] ), .B(n10327), .X(n9161) );
  nand_x1_sg U10828 ( .A(\reg_in[1][0][18] ), .B(n10538), .X(n9162) );
  nand_x1_sg U10829 ( .A(\in[1][0][19] ), .B(n10631), .X(n9159) );
  nand_x1_sg U10830 ( .A(\reg_in[1][0][19] ), .B(n10531), .X(n9160) );
  nand_x1_sg U10831 ( .A(\in[1][1][0] ), .B(n10619), .X(n9157) );
  nand_x1_sg U10832 ( .A(\reg_in[1][1][0] ), .B(n10578), .X(n9158) );
  nand_x1_sg U10833 ( .A(\in[1][1][1] ), .B(n10323), .X(n9155) );
  nand_x1_sg U10834 ( .A(\reg_in[1][1][1] ), .B(n10287), .X(n9156) );
  nand_x1_sg U10835 ( .A(\in[1][1][2] ), .B(n10606), .X(n9153) );
  nand_x1_sg U10836 ( .A(\reg_in[1][1][2] ), .B(n10285), .X(n9154) );
  nand_x1_sg U10837 ( .A(\in[1][1][3] ), .B(n10081), .X(n9151) );
  nand_x1_sg U10838 ( .A(\reg_in[1][1][3] ), .B(n10580), .X(n9152) );
  nand_x1_sg U10839 ( .A(\in[1][1][4] ), .B(n10390), .X(n9149) );
  nand_x1_sg U10840 ( .A(\reg_in[1][1][4] ), .B(n10482), .X(n9150) );
  nand_x1_sg U10841 ( .A(\in[1][1][5] ), .B(n10023), .X(n9147) );
  nand_x1_sg U10842 ( .A(\reg_in[1][1][5] ), .B(n10580), .X(n9148) );
  nand_x1_sg U10843 ( .A(\in[1][1][6] ), .B(n10330), .X(n9145) );
  nand_x1_sg U10844 ( .A(\reg_in[1][1][6] ), .B(n10306), .X(n9146) );
  nand_x1_sg U10845 ( .A(\in[1][1][7] ), .B(n10321), .X(n9143) );
  nand_x1_sg U10846 ( .A(\reg_in[1][1][7] ), .B(n10267), .X(n9144) );
  nand_x1_sg U10847 ( .A(\in[1][1][8] ), .B(n10315), .X(n9141) );
  nand_x1_sg U10848 ( .A(\reg_in[1][1][8] ), .B(n10189), .X(n9142) );
  nand_x1_sg U10849 ( .A(\in[1][1][9] ), .B(n10330), .X(n9139) );
  nand_x1_sg U10850 ( .A(\reg_in[1][1][9] ), .B(n10060), .X(n9140) );
  nand_x1_sg U10851 ( .A(\in[1][1][10] ), .B(n10322), .X(n9137) );
  nand_x1_sg U10852 ( .A(\reg_in[1][1][10] ), .B(n10482), .X(n9138) );
  nand_x1_sg U10853 ( .A(\in[1][1][11] ), .B(n10394), .X(n9135) );
  nand_x1_sg U10854 ( .A(\reg_in[1][1][11] ), .B(n10481), .X(n9136) );
  nand_x1_sg U10855 ( .A(\in[1][1][12] ), .B(n10320), .X(n9133) );
  nand_x1_sg U10856 ( .A(\reg_in[1][1][12] ), .B(n10192), .X(n9134) );
  nand_x1_sg U10857 ( .A(\in[1][1][13] ), .B(n10259), .X(n9131) );
  nand_x1_sg U10858 ( .A(\reg_in[1][1][13] ), .B(n10479), .X(n9132) );
  nand_x1_sg U10859 ( .A(\in[1][1][14] ), .B(n10602), .X(n9129) );
  nand_x1_sg U10860 ( .A(\reg_in[1][1][14] ), .B(n10270), .X(n9130) );
  nand_x1_sg U10861 ( .A(\in[1][2][0] ), .B(n10626), .X(n9117) );
  nand_x1_sg U10862 ( .A(\reg_in[1][2][0] ), .B(n10477), .X(n9118) );
  nand_x1_sg U10863 ( .A(\in[1][2][1] ), .B(n10317), .X(n9115) );
  nand_x1_sg U10864 ( .A(\reg_in[1][2][1] ), .B(n10211), .X(n9116) );
  nand_x1_sg U10865 ( .A(\in[1][2][2] ), .B(n10620), .X(n9113) );
  nand_x1_sg U10866 ( .A(\reg_in[1][2][2] ), .B(n10286), .X(n9114) );
  nand_x1_sg U10867 ( .A(\in[1][2][3] ), .B(n10323), .X(n9111) );
  nand_x1_sg U10868 ( .A(\reg_in[1][2][3] ), .B(n10301), .X(n9112) );
  nand_x1_sg U10869 ( .A(\in[1][2][4] ), .B(n10311), .X(n9109) );
  nand_x1_sg U10870 ( .A(\reg_in[1][2][4] ), .B(n10574), .X(n9110) );
  nand_x1_sg U10871 ( .A(\in[1][2][5] ), .B(n10312), .X(n9107) );
  nand_x1_sg U10872 ( .A(\reg_in[1][2][5] ), .B(n10302), .X(n9108) );
  nand_x1_sg U10873 ( .A(\in[1][2][6] ), .B(n10400), .X(n9105) );
  nand_x1_sg U10874 ( .A(\reg_in[1][2][6] ), .B(n10531), .X(n9106) );
  nand_x1_sg U10875 ( .A(\in[1][2][7] ), .B(n10411), .X(n9103) );
  nand_x1_sg U10876 ( .A(\reg_in[1][2][7] ), .B(n10525), .X(n9104) );
  nand_x1_sg U10877 ( .A(\in[1][2][8] ), .B(n10606), .X(n9101) );
  nand_x1_sg U10878 ( .A(\reg_in[1][2][8] ), .B(n10301), .X(n9102) );
  nand_x1_sg U10879 ( .A(\in[1][2][9] ), .B(n10328), .X(n9099) );
  nand_x1_sg U10880 ( .A(\reg_in[1][2][9] ), .B(n10302), .X(n9100) );
  nand_x1_sg U10881 ( .A(\in[1][2][10] ), .B(n10402), .X(n9097) );
  nand_x1_sg U10882 ( .A(\reg_in[1][2][10] ), .B(n10306), .X(n9098) );
  nand_x1_sg U10883 ( .A(\in[1][2][11] ), .B(n10608), .X(n9095) );
  nand_x1_sg U10884 ( .A(\reg_in[1][2][11] ), .B(n10188), .X(n9096) );
  nand_x1_sg U10885 ( .A(\in[1][2][12] ), .B(n10396), .X(n9093) );
  nand_x1_sg U10886 ( .A(\reg_in[1][2][12] ), .B(n10535), .X(n9094) );
  nand_x1_sg U10887 ( .A(\in[1][2][13] ), .B(n10627), .X(n9091) );
  nand_x1_sg U10888 ( .A(\reg_in[1][2][13] ), .B(n10304), .X(n9092) );
  nand_x1_sg U10889 ( .A(\in[1][2][14] ), .B(n10607), .X(n9089) );
  nand_x1_sg U10890 ( .A(\reg_in[1][2][14] ), .B(n10538), .X(n9090) );
  nand_x1_sg U10891 ( .A(\in[1][2][15] ), .B(n10336), .X(n9087) );
  nand_x1_sg U10892 ( .A(\reg_in[1][2][15] ), .B(n10479), .X(n9088) );
  nand_x1_sg U10893 ( .A(\in[1][2][16] ), .B(n10083), .X(n9085) );
  nand_x1_sg U10894 ( .A(\reg_in[1][2][16] ), .B(n10213), .X(n9086) );
  nand_x1_sg U10895 ( .A(\in[1][2][17] ), .B(n10084), .X(n9083) );
  nand_x1_sg U10896 ( .A(\reg_in[1][2][17] ), .B(n10477), .X(n9084) );
  nand_x1_sg U10897 ( .A(\in[1][2][18] ), .B(n10628), .X(n9081) );
  nand_x1_sg U10898 ( .A(\reg_in[1][2][18] ), .B(n10308), .X(n9082) );
  nand_x1_sg U10899 ( .A(\in[1][2][19] ), .B(n10317), .X(n9079) );
  nand_x1_sg U10900 ( .A(\reg_in[1][2][19] ), .B(n10183), .X(n9080) );
  nand_x1_sg U10901 ( .A(\in[1][3][0] ), .B(n10315), .X(n9077) );
  nand_x1_sg U10902 ( .A(\reg_in[1][3][0] ), .B(n10524), .X(n9078) );
  nand_x1_sg U10903 ( .A(\in[1][3][1] ), .B(n10602), .X(n9075) );
  nand_x1_sg U10904 ( .A(\reg_in[1][3][1] ), .B(n10213), .X(n9076) );
  nand_x1_sg U10905 ( .A(\in[1][3][2] ), .B(n10600), .X(n9073) );
  nand_x1_sg U10906 ( .A(\reg_in[1][3][2] ), .B(n10576), .X(n9074) );
  nand_x1_sg U10907 ( .A(\in[1][3][3] ), .B(n10616), .X(n9071) );
  nand_x1_sg U10908 ( .A(\reg_in[1][3][3] ), .B(n10140), .X(n9072) );
  nand_x1_sg U10909 ( .A(\in[1][3][4] ), .B(n10081), .X(n9069) );
  nand_x1_sg U10910 ( .A(\reg_in[1][3][4] ), .B(n10524), .X(n9070) );
  nand_x1_sg U10911 ( .A(\in[1][3][5] ), .B(n10332), .X(n9067) );
  nand_x1_sg U10912 ( .A(\reg_in[1][3][5] ), .B(n10527), .X(n9068) );
  nand_x1_sg U10913 ( .A(\in[1][3][6] ), .B(n10339), .X(n9065) );
  nand_x1_sg U10914 ( .A(\reg_in[1][3][6] ), .B(n10473), .X(n9066) );
  nand_x1_sg U10915 ( .A(\in[1][3][7] ), .B(n10396), .X(n9063) );
  nand_x1_sg U10916 ( .A(\reg_in[1][3][7] ), .B(n10484), .X(n9064) );
  nand_x1_sg U10917 ( .A(\in[1][3][8] ), .B(n10617), .X(n9061) );
  nand_x1_sg U10918 ( .A(\reg_in[1][3][8] ), .B(n10189), .X(n9062) );
  nand_x1_sg U10919 ( .A(\in[1][3][9] ), .B(n10386), .X(n9059) );
  nand_x1_sg U10920 ( .A(\reg_in[1][3][9] ), .B(n10179), .X(n9060) );
  nand_x1_sg U10921 ( .A(\in[1][3][15] ), .B(n10614), .X(n9047) );
  nand_x1_sg U10922 ( .A(\reg_in[1][3][15] ), .B(n10540), .X(n9048) );
  nand_x1_sg U10923 ( .A(\in[1][3][16] ), .B(n10631), .X(n9045) );
  nand_x1_sg U10924 ( .A(\reg_in[1][3][16] ), .B(n10184), .X(n9046) );
  nand_x1_sg U10925 ( .A(\in[1][3][17] ), .B(n10258), .X(n9043) );
  nand_x1_sg U10926 ( .A(\reg_in[1][3][17] ), .B(n10484), .X(n9044) );
  nand_x1_sg U10927 ( .A(\in[1][3][18] ), .B(n10021), .X(n9041) );
  nand_x1_sg U10928 ( .A(\reg_in[1][3][18] ), .B(n10474), .X(n9042) );
  nand_x1_sg U10929 ( .A(\in[1][3][19] ), .B(n10311), .X(n9039) );
  nand_x1_sg U10930 ( .A(\reg_in[1][3][19] ), .B(n10576), .X(n9040) );
  nand_x1_sg U10931 ( .A(\in[2][0][0] ), .B(n10393), .X(n9037) );
  nand_x1_sg U10932 ( .A(\reg_in[2][0][0] ), .B(n10179), .X(n9038) );
  nand_x1_sg U10933 ( .A(\in[2][0][1] ), .B(n10624), .X(n9035) );
  nand_x1_sg U10934 ( .A(\reg_in[2][0][1] ), .B(n10302), .X(n9036) );
  nand_x1_sg U10935 ( .A(\in[2][0][2] ), .B(n10402), .X(n9033) );
  nand_x1_sg U10936 ( .A(\reg_in[2][0][2] ), .B(n10538), .X(n9034) );
  nand_x1_sg U10937 ( .A(\in[2][0][3] ), .B(n10389), .X(n9031) );
  nand_x1_sg U10938 ( .A(\reg_in[2][0][3] ), .B(n10480), .X(n9032) );
  nand_x1_sg U10939 ( .A(\in[2][0][4] ), .B(n10074), .X(n9029) );
  nand_x1_sg U10940 ( .A(\reg_in[2][0][4] ), .B(n10307), .X(n9030) );
  nand_x1_sg U10941 ( .A(\in[2][0][5] ), .B(n10615), .X(n9027) );
  nand_x1_sg U10942 ( .A(\reg_in[2][0][5] ), .B(n10305), .X(n9028) );
  nand_x1_sg U10943 ( .A(\in[2][0][6] ), .B(n10608), .X(n9025) );
  nand_x1_sg U10944 ( .A(\reg_in[2][0][6] ), .B(n10571), .X(n9026) );
  nand_x1_sg U10945 ( .A(\in[2][0][7] ), .B(n10312), .X(n9023) );
  nand_x1_sg U10946 ( .A(\reg_in[2][0][7] ), .B(n10056), .X(n9024) );
  nand_x1_sg U10947 ( .A(\in[2][0][8] ), .B(n10624), .X(n9021) );
  nand_x1_sg U10948 ( .A(\reg_in[2][0][8] ), .B(n10057), .X(n9022) );
  nand_x1_sg U10949 ( .A(\in[2][0][9] ), .B(n10317), .X(n9019) );
  nand_x1_sg U10950 ( .A(\reg_in[2][0][9] ), .B(n10540), .X(n9020) );
  nand_x1_sg U10951 ( .A(\in[2][0][10] ), .B(n10073), .X(n9017) );
  nand_x1_sg U10952 ( .A(\reg_in[2][0][10] ), .B(n10303), .X(n9018) );
  nand_x1_sg U10953 ( .A(\in[2][0][11] ), .B(n10600), .X(n9015) );
  nand_x1_sg U10954 ( .A(\reg_in[2][0][11] ), .B(n10058), .X(n9016) );
  nand_x1_sg U10955 ( .A(\in[2][0][12] ), .B(n10311), .X(n9013) );
  nand_x1_sg U10956 ( .A(\reg_in[2][0][12] ), .B(n10572), .X(n9014) );
  nand_x1_sg U10957 ( .A(\in[2][0][13] ), .B(n10323), .X(n9011) );
  nand_x1_sg U10958 ( .A(\reg_in[2][0][13] ), .B(n10482), .X(n9012) );
  nand_x1_sg U10959 ( .A(\in[2][0][14] ), .B(n10079), .X(n9009) );
  nand_x1_sg U10960 ( .A(\reg_in[2][0][14] ), .B(n10265), .X(n9010) );
  nand_x1_sg U10961 ( .A(\in[2][0][15] ), .B(n10086), .X(n9007) );
  nand_x1_sg U10962 ( .A(\reg_in[2][0][15] ), .B(n10475), .X(n9008) );
  nand_x1_sg U10963 ( .A(\in[2][0][16] ), .B(n10330), .X(n9005) );
  nand_x1_sg U10964 ( .A(\reg_in[2][0][16] ), .B(n10214), .X(n9006) );
  nand_x1_sg U10965 ( .A(\in[2][0][17] ), .B(n10612), .X(n9003) );
  nand_x1_sg U10966 ( .A(\reg_in[2][0][17] ), .B(n10523), .X(n9004) );
  nand_x1_sg U10967 ( .A(\in[2][0][18] ), .B(n10392), .X(n9001) );
  nand_x1_sg U10968 ( .A(\reg_in[2][0][18] ), .B(n10574), .X(n9002) );
  nand_x1_sg U10969 ( .A(\in[2][0][19] ), .B(n10628), .X(n8999) );
  nand_x1_sg U10970 ( .A(\reg_in[2][0][19] ), .B(n10572), .X(n9000) );
  nand_x1_sg U10971 ( .A(\in[2][1][5] ), .B(n10394), .X(n8987) );
  nand_x1_sg U10972 ( .A(\reg_in[2][1][5] ), .B(n10141), .X(n8988) );
  nand_x1_sg U10973 ( .A(\in[2][1][6] ), .B(n10259), .X(n8985) );
  nand_x1_sg U10974 ( .A(\reg_in[2][1][6] ), .B(n10474), .X(n8986) );
  nand_x1_sg U10975 ( .A(\in[2][1][7] ), .B(n10408), .X(n8983) );
  nand_x1_sg U10976 ( .A(\reg_in[2][1][7] ), .B(n10536), .X(n8984) );
  nand_x1_sg U10977 ( .A(\in[2][1][8] ), .B(n10340), .X(n8981) );
  nand_x1_sg U10978 ( .A(\reg_in[2][1][8] ), .B(n10041), .X(n8982) );
  nand_x1_sg U10979 ( .A(\in[2][1][9] ), .B(n10408), .X(n8979) );
  nand_x1_sg U10980 ( .A(\reg_in[2][1][9] ), .B(n10057), .X(n8980) );
  nand_x1_sg U10981 ( .A(\in[2][1][10] ), .B(n10081), .X(n8977) );
  nand_x1_sg U10982 ( .A(\reg_in[2][1][10] ), .B(n10539), .X(n8978) );
  nand_x1_sg U10983 ( .A(\in[2][1][11] ), .B(n10408), .X(n8975) );
  nand_x1_sg U10984 ( .A(\reg_in[2][1][11] ), .B(n10191), .X(n8976) );
  nand_x1_sg U10985 ( .A(\in[2][1][12] ), .B(n10080), .X(n8973) );
  nand_x1_sg U10986 ( .A(\reg_in[2][1][12] ), .B(n10288), .X(n8974) );
  nand_x1_sg U10987 ( .A(\in[2][1][13] ), .B(n10327), .X(n8971) );
  nand_x1_sg U10988 ( .A(\reg_in[2][1][13] ), .B(n10475), .X(n8972) );
  nand_x1_sg U10989 ( .A(\in[2][1][14] ), .B(n10320), .X(n8969) );
  nand_x1_sg U10990 ( .A(\reg_in[2][1][14] ), .B(n10270), .X(n8970) );
  nand_x1_sg U10991 ( .A(\in[2][2][0] ), .B(n10601), .X(n8957) );
  nand_x1_sg U10992 ( .A(\reg_in[2][2][0] ), .B(n10524), .X(n8958) );
  nand_x1_sg U10993 ( .A(\in[2][2][1] ), .B(n10626), .X(n8955) );
  nand_x1_sg U10994 ( .A(\reg_in[2][2][1] ), .B(n10580), .X(n8956) );
  nand_x1_sg U10995 ( .A(\in[2][2][2] ), .B(n10073), .X(n8953) );
  nand_x1_sg U10996 ( .A(\reg_in[2][2][2] ), .B(n10534), .X(n8954) );
  nand_x1_sg U10997 ( .A(\in[2][2][3] ), .B(n10628), .X(n8951) );
  nand_x1_sg U10998 ( .A(\reg_in[2][2][3] ), .B(n10060), .X(n8952) );
  nand_x1_sg U10999 ( .A(\in[2][2][4] ), .B(n10023), .X(n8949) );
  nand_x1_sg U11000 ( .A(\reg_in[2][2][4] ), .B(n10476), .X(n8950) );
  nand_x1_sg U11001 ( .A(\in[2][2][5] ), .B(n10322), .X(n8947) );
  nand_x1_sg U11002 ( .A(\reg_in[2][2][5] ), .B(n10216), .X(n8948) );
  nand_x1_sg U11003 ( .A(\in[2][2][6] ), .B(n10605), .X(n8945) );
  nand_x1_sg U11004 ( .A(\reg_in[2][2][6] ), .B(n10217), .X(n8946) );
  nand_x1_sg U11005 ( .A(\in[2][2][7] ), .B(n10392), .X(n8943) );
  nand_x1_sg U11006 ( .A(\reg_in[2][2][7] ), .B(n10286), .X(n8944) );
  nand_x1_sg U11007 ( .A(\in[2][2][8] ), .B(n10632), .X(n8941) );
  nand_x1_sg U11008 ( .A(\reg_in[2][2][8] ), .B(n10267), .X(n8942) );
  nand_x1_sg U11009 ( .A(\in[2][2][9] ), .B(n10631), .X(n8939) );
  nand_x1_sg U11010 ( .A(\reg_in[2][2][9] ), .B(n10307), .X(n8940) );
  nand_x1_sg U11011 ( .A(\in[2][2][15] ), .B(n10627), .X(n8927) );
  nand_x1_sg U11012 ( .A(\reg_in[2][2][15] ), .B(n10188), .X(n8928) );
  nand_x1_sg U11013 ( .A(\in[2][2][16] ), .B(n10604), .X(n8925) );
  nand_x1_sg U11014 ( .A(\reg_in[2][2][16] ), .B(n10191), .X(n8926) );
  nand_x1_sg U11015 ( .A(\in[2][2][17] ), .B(n10616), .X(n8923) );
  nand_x1_sg U11016 ( .A(\reg_in[2][2][17] ), .B(n10266), .X(n8924) );
  nand_x1_sg U11017 ( .A(\in[2][2][18] ), .B(n10323), .X(n8921) );
  nand_x1_sg U11018 ( .A(\reg_in[2][2][18] ), .B(n10579), .X(n8922) );
  nand_x1_sg U11019 ( .A(\in[2][2][19] ), .B(n10613), .X(n8919) );
  nand_x1_sg U11020 ( .A(\reg_in[2][2][19] ), .B(n10214), .X(n8920) );
  nand_x1_sg U11021 ( .A(\in[2][3][0] ), .B(n10338), .X(n8917) );
  nand_x1_sg U11022 ( .A(\reg_in[2][3][0] ), .B(n10530), .X(n8918) );
  nand_x1_sg U11023 ( .A(\in[2][3][1] ), .B(n10315), .X(n8915) );
  nand_x1_sg U11024 ( .A(\reg_in[2][3][1] ), .B(n10541), .X(n8916) );
  nand_x1_sg U11025 ( .A(\in[2][3][2] ), .B(n10625), .X(n8913) );
  nand_x1_sg U11026 ( .A(\reg_in[2][3][2] ), .B(n10178), .X(n8914) );
  nand_x1_sg U11027 ( .A(\in[2][3][3] ), .B(n10316), .X(n8911) );
  nand_x1_sg U11028 ( .A(\reg_in[2][3][3] ), .B(n10042), .X(n8912) );
  nand_x1_sg U11029 ( .A(\in[2][3][4] ), .B(n10616), .X(n8909) );
  nand_x1_sg U11030 ( .A(\reg_in[2][3][4] ), .B(n10189), .X(n8910) );
  nand_x1_sg U11031 ( .A(\in[2][3][5] ), .B(n10316), .X(n8907) );
  nand_x1_sg U11032 ( .A(\reg_in[2][3][5] ), .B(n10533), .X(n8908) );
  nand_x1_sg U11033 ( .A(\in[2][3][6] ), .B(n10615), .X(n8905) );
  nand_x1_sg U11034 ( .A(\reg_in[2][3][6] ), .B(n10574), .X(n8906) );
  nand_x1_sg U11035 ( .A(\in[2][3][7] ), .B(n10320), .X(n8903) );
  nand_x1_sg U11036 ( .A(\reg_in[2][3][7] ), .B(n10059), .X(n8904) );
  nand_x1_sg U11037 ( .A(\in[2][3][8] ), .B(n10630), .X(n8901) );
  nand_x1_sg U11038 ( .A(\reg_in[2][3][8] ), .B(n10141), .X(n8902) );
  nand_x1_sg U11039 ( .A(\in[2][3][9] ), .B(n10074), .X(n8899) );
  nand_x1_sg U11040 ( .A(\reg_in[2][3][9] ), .B(n10287), .X(n8900) );
  nand_x1_sg U11041 ( .A(\in[2][3][10] ), .B(n10258), .X(n8897) );
  nand_x1_sg U11042 ( .A(\reg_in[2][3][10] ), .B(n10575), .X(n8898) );
  nand_x1_sg U11043 ( .A(\in[2][3][11] ), .B(n10394), .X(n8895) );
  nand_x1_sg U11044 ( .A(\reg_in[2][3][11] ), .B(n10144), .X(n8896) );
  nand_x1_sg U11045 ( .A(\in[2][3][12] ), .B(n10321), .X(n8893) );
  nand_x1_sg U11046 ( .A(\reg_in[2][3][12] ), .B(n10525), .X(n8894) );
  nand_x1_sg U11047 ( .A(\in[2][3][13] ), .B(n10326), .X(n8891) );
  nand_x1_sg U11048 ( .A(\reg_in[2][3][13] ), .B(n10268), .X(n8892) );
  nand_x1_sg U11049 ( .A(\in[2][3][14] ), .B(n10390), .X(n8889) );
  nand_x1_sg U11050 ( .A(\reg_in[2][3][14] ), .B(n10579), .X(n8890) );
  nand_x1_sg U11051 ( .A(\in[2][3][15] ), .B(n10326), .X(n8887) );
  nand_x1_sg U11052 ( .A(\reg_in[2][3][15] ), .B(n10213), .X(n8888) );
  nand_x1_sg U11053 ( .A(\in[2][3][16] ), .B(n10615), .X(n8885) );
  nand_x1_sg U11054 ( .A(\reg_in[2][3][16] ), .B(n10305), .X(n8886) );
  nand_x1_sg U11055 ( .A(\in[2][3][17] ), .B(n10312), .X(n8883) );
  nand_x1_sg U11056 ( .A(\reg_in[2][3][17] ), .B(n10476), .X(n8884) );
  nand_x1_sg U11057 ( .A(\in[2][3][18] ), .B(n10339), .X(n8881) );
  nand_x1_sg U11058 ( .A(\reg_in[2][3][18] ), .B(n10525), .X(n8882) );
  nand_x1_sg U11059 ( .A(\in[2][3][19] ), .B(n10083), .X(n8879) );
  nand_x1_sg U11060 ( .A(\reg_in[2][3][19] ), .B(n10286), .X(n8880) );
  nand_x1_sg U11061 ( .A(\in[3][0][5] ), .B(n10613), .X(n8867) );
  nand_x1_sg U11062 ( .A(\reg_in[3][0][5] ), .B(n10541), .X(n8868) );
  nand_x1_sg U11063 ( .A(\in[3][0][6] ), .B(n10334), .X(n8865) );
  nand_x1_sg U11064 ( .A(\reg_in[3][0][6] ), .B(n10480), .X(n8866) );
  nand_x1_sg U11065 ( .A(\in[3][0][7] ), .B(n10324), .X(n8863) );
  nand_x1_sg U11066 ( .A(\reg_in[3][0][7] ), .B(n10540), .X(n8864) );
  nand_x1_sg U11067 ( .A(\in[3][0][8] ), .B(n10602), .X(n8861) );
  nand_x1_sg U11068 ( .A(\reg_in[3][0][8] ), .B(n10056), .X(n8862) );
  nand_x1_sg U11069 ( .A(\in[3][0][9] ), .B(n10618), .X(n8859) );
  nand_x1_sg U11070 ( .A(\reg_in[3][0][9] ), .B(n10536), .X(n8860) );
  nand_x1_sg U11071 ( .A(\in[3][0][10] ), .B(n10614), .X(n8857) );
  nand_x1_sg U11072 ( .A(\reg_in[3][0][10] ), .B(n10533), .X(n8858) );
  nand_x1_sg U11073 ( .A(\in[3][0][11] ), .B(n10613), .X(n8855) );
  nand_x1_sg U11074 ( .A(\reg_in[3][0][11] ), .B(n10570), .X(n8856) );
  nand_x1_sg U11075 ( .A(\in[3][0][12] ), .B(n10399), .X(n8853) );
  nand_x1_sg U11076 ( .A(\reg_in[3][0][12] ), .B(n10579), .X(n8854) );
  nand_x1_sg U11077 ( .A(\in[3][0][13] ), .B(n10074), .X(n8851) );
  nand_x1_sg U11078 ( .A(\reg_in[3][0][13] ), .B(n10217), .X(n8852) );
  nand_x1_sg U11079 ( .A(\in[3][0][14] ), .B(n10259), .X(n8849) );
  nand_x1_sg U11080 ( .A(\reg_in[3][0][14] ), .B(n10571), .X(n8850) );
  nand_x1_sg U11081 ( .A(\in[3][0][15] ), .B(n10079), .X(n8847) );
  nand_x1_sg U11082 ( .A(\reg_in[3][0][15] ), .B(n10578), .X(n8848) );
  nand_x1_sg U11083 ( .A(\in[3][0][16] ), .B(n10315), .X(n8845) );
  nand_x1_sg U11084 ( .A(\reg_in[3][0][16] ), .B(n10267), .X(n8846) );
  nand_x1_sg U11085 ( .A(\in[3][0][17] ), .B(n10393), .X(n8843) );
  nand_x1_sg U11086 ( .A(\reg_in[3][0][17] ), .B(n10043), .X(n8844) );
  nand_x1_sg U11087 ( .A(\in[3][0][18] ), .B(n10607), .X(n8841) );
  nand_x1_sg U11088 ( .A(\reg_in[3][0][18] ), .B(n10215), .X(n8842) );
  nand_x1_sg U11089 ( .A(\in[3][0][19] ), .B(n10387), .X(n8839) );
  nand_x1_sg U11090 ( .A(\reg_in[3][0][19] ), .B(n10179), .X(n8840) );
  nand_x1_sg U11091 ( .A(\in[3][1][0] ), .B(n10334), .X(n8837) );
  nand_x1_sg U11092 ( .A(\reg_in[3][1][0] ), .B(n10058), .X(n8838) );
  nand_x1_sg U11093 ( .A(\in[3][1][1] ), .B(n10625), .X(n8835) );
  nand_x1_sg U11094 ( .A(\reg_in[3][1][1] ), .B(n10474), .X(n8836) );
  nand_x1_sg U11095 ( .A(\in[3][1][2] ), .B(n10079), .X(n8833) );
  nand_x1_sg U11096 ( .A(\reg_in[3][1][2] ), .B(n10268), .X(n8834) );
  nand_x1_sg U11097 ( .A(\in[3][1][3] ), .B(n10328), .X(n8831) );
  nand_x1_sg U11098 ( .A(\reg_in[3][1][3] ), .B(n10479), .X(n8832) );
  nand_x1_sg U11099 ( .A(\in[3][1][4] ), .B(n10396), .X(n8829) );
  nand_x1_sg U11100 ( .A(\reg_in[3][1][4] ), .B(n10212), .X(n8830) );
  nand_x1_sg U11101 ( .A(\in[3][1][5] ), .B(n10328), .X(n8827) );
  nand_x1_sg U11102 ( .A(\reg_in[3][1][5] ), .B(n10215), .X(n8828) );
  nand_x1_sg U11103 ( .A(\in[3][1][6] ), .B(n10387), .X(n8825) );
  nand_x1_sg U11104 ( .A(\reg_in[3][1][6] ), .B(n10530), .X(n8826) );
  nand_x1_sg U11105 ( .A(\in[3][1][7] ), .B(n10388), .X(n8823) );
  nand_x1_sg U11106 ( .A(\reg_in[3][1][7] ), .B(n10522), .X(n8824) );
  nand_x1_sg U11107 ( .A(\in[3][1][8] ), .B(n10390), .X(n8821) );
  nand_x1_sg U11108 ( .A(\reg_in[3][1][8] ), .B(n10178), .X(n8822) );
  nand_x1_sg U11109 ( .A(\in[3][1][9] ), .B(n10389), .X(n8819) );
  nand_x1_sg U11110 ( .A(\reg_in[3][1][9] ), .B(n10307), .X(n8820) );
  nand_x1_sg U11111 ( .A(\in[3][1][10] ), .B(n10604), .X(n8817) );
  nand_x1_sg U11112 ( .A(\reg_in[3][1][10] ), .B(n10473), .X(n8818) );
  nand_x1_sg U11113 ( .A(\in[3][1][11] ), .B(n10336), .X(n8815) );
  nand_x1_sg U11114 ( .A(\reg_in[3][1][11] ), .B(n10481), .X(n8816) );
  nand_x1_sg U11115 ( .A(\in[3][1][12] ), .B(n10086), .X(n8813) );
  nand_x1_sg U11116 ( .A(\reg_in[3][1][12] ), .B(n10572), .X(n8814) );
  nand_x1_sg U11117 ( .A(\in[3][1][13] ), .B(n10388), .X(n8811) );
  nand_x1_sg U11118 ( .A(\reg_in[3][1][13] ), .B(n10576), .X(n8812) );
  nand_x1_sg U11119 ( .A(\in[3][1][14] ), .B(n10608), .X(n8809) );
  nand_x1_sg U11120 ( .A(\reg_in[3][1][14] ), .B(n10042), .X(n8810) );
  nand_x1_sg U11121 ( .A(\in[3][2][0] ), .B(n10386), .X(n8797) );
  nand_x1_sg U11122 ( .A(\reg_in[3][2][0] ), .B(n10528), .X(n8798) );
  nand_x1_sg U11123 ( .A(\in[3][2][1] ), .B(n10606), .X(n8795) );
  nand_x1_sg U11124 ( .A(\reg_in[3][2][1] ), .B(n10579), .X(n8796) );
  nand_x1_sg U11125 ( .A(\in[3][2][2] ), .B(n10631), .X(n8793) );
  nand_x1_sg U11126 ( .A(\reg_in[3][2][2] ), .B(n10178), .X(n8794) );
  nand_x1_sg U11127 ( .A(\in[3][2][3] ), .B(n10322), .X(n8791) );
  nand_x1_sg U11128 ( .A(\reg_in[3][2][3] ), .B(n10530), .X(n8792) );
  nand_x1_sg U11129 ( .A(\in[3][2][4] ), .B(n10395), .X(n8789) );
  nand_x1_sg U11130 ( .A(\reg_in[3][2][4] ), .B(n10054), .X(n8790) );
  nand_x1_sg U11131 ( .A(\in[3][2][5] ), .B(n10388), .X(n8787) );
  nand_x1_sg U11132 ( .A(\reg_in[3][2][5] ), .B(n10285), .X(n8788) );
  nand_x1_sg U11133 ( .A(\in[3][2][6] ), .B(n10321), .X(n8785) );
  nand_x1_sg U11134 ( .A(\reg_in[3][2][6] ), .B(n10188), .X(n8786) );
  nand_x1_sg U11135 ( .A(\in[3][2][7] ), .B(n10625), .X(n8783) );
  nand_x1_sg U11136 ( .A(\reg_in[3][2][7] ), .B(n10145), .X(n8784) );
  nand_x1_sg U11137 ( .A(\in[3][2][8] ), .B(n10629), .X(n8781) );
  nand_x1_sg U11138 ( .A(\reg_in[3][2][8] ), .B(n10140), .X(n8782) );
  nand_x1_sg U11139 ( .A(\in[3][2][9] ), .B(n10389), .X(n8779) );
  nand_x1_sg U11140 ( .A(\reg_in[3][2][9] ), .B(n10478), .X(n8780) );
  nand_x1_sg U11141 ( .A(\in[3][2][10] ), .B(n10335), .X(n8777) );
  nand_x1_sg U11142 ( .A(\reg_in[3][2][10] ), .B(n10269), .X(n8778) );
  nand_x1_sg U11143 ( .A(\in[3][2][11] ), .B(n10318), .X(n8775) );
  nand_x1_sg U11144 ( .A(\reg_in[3][2][11] ), .B(n10184), .X(n8776) );
  nand_x1_sg U11145 ( .A(\in[3][2][12] ), .B(n10312), .X(n8773) );
  nand_x1_sg U11146 ( .A(\reg_in[3][2][12] ), .B(n10473), .X(n8774) );
  nand_x1_sg U11147 ( .A(\in[3][2][13] ), .B(n10336), .X(n8771) );
  nand_x1_sg U11148 ( .A(\reg_in[3][2][13] ), .B(n10304), .X(n8772) );
  nand_x1_sg U11149 ( .A(\in[3][2][14] ), .B(n10386), .X(n8769) );
  nand_x1_sg U11150 ( .A(\reg_in[3][2][14] ), .B(n10576), .X(n8770) );
  nand_x1_sg U11151 ( .A(\in[3][2][15] ), .B(n10077), .X(n8767) );
  nand_x1_sg U11152 ( .A(\reg_in[3][2][15] ), .B(n10483), .X(n8768) );
  nand_x1_sg U11153 ( .A(\in[3][2][16] ), .B(n10605), .X(n8765) );
  nand_x1_sg U11154 ( .A(\reg_in[3][2][16] ), .B(n10288), .X(n8766) );
  nand_x1_sg U11155 ( .A(\in[3][2][17] ), .B(n10602), .X(n8763) );
  nand_x1_sg U11156 ( .A(\reg_in[3][2][17] ), .B(n10265), .X(n8764) );
  nand_x1_sg U11157 ( .A(\in[3][2][18] ), .B(n10387), .X(n8761) );
  nand_x1_sg U11158 ( .A(\reg_in[3][2][18] ), .B(n10188), .X(n8762) );
  nand_x1_sg U11159 ( .A(\in[3][2][19] ), .B(n10077), .X(n8759) );
  nand_x1_sg U11160 ( .A(\reg_in[3][2][19] ), .B(n10288), .X(n8760) );
  nand_x1_sg U11161 ( .A(\in[3][3][0] ), .B(n10628), .X(n8757) );
  nand_x1_sg U11162 ( .A(\reg_in[3][3][0] ), .B(n10536), .X(n8758) );
  nand_x1_sg U11163 ( .A(\in[3][3][1] ), .B(n10398), .X(n8755) );
  nand_x1_sg U11164 ( .A(\reg_in[3][3][1] ), .B(n10475), .X(n8756) );
  nand_x1_sg U11165 ( .A(\in[3][3][2] ), .B(n10630), .X(n8753) );
  nand_x1_sg U11166 ( .A(\reg_in[3][3][2] ), .B(n10267), .X(n8754) );
  nand_x1_sg U11167 ( .A(\in[3][3][3] ), .B(n10329), .X(n8751) );
  nand_x1_sg U11168 ( .A(\reg_in[3][3][3] ), .B(n10480), .X(n8752) );
  nand_x1_sg U11169 ( .A(\in[3][3][4] ), .B(n10321), .X(n8749) );
  nand_x1_sg U11170 ( .A(\reg_in[3][3][4] ), .B(n10270), .X(n8750) );
  nand_x1_sg U11171 ( .A(\in[3][3][10] ), .B(n10411), .X(n8737) );
  nand_x1_sg U11172 ( .A(\reg_in[3][3][10] ), .B(n10484), .X(n8738) );
  nand_x1_sg U11173 ( .A(\in[3][3][11] ), .B(n10318), .X(n8735) );
  nand_x1_sg U11174 ( .A(\reg_in[3][3][11] ), .B(n10060), .X(n8736) );
  nand_x1_sg U11175 ( .A(\in[3][3][12] ), .B(n10322), .X(n8733) );
  nand_x1_sg U11176 ( .A(\reg_in[3][3][12] ), .B(n10308), .X(n8734) );
  nand_x1_sg U11177 ( .A(\in[3][3][13] ), .B(n10073), .X(n8731) );
  nand_x1_sg U11178 ( .A(\reg_in[3][3][13] ), .B(n10536), .X(n8732) );
  nand_x1_sg U11179 ( .A(\in[3][3][14] ), .B(n10320), .X(n8729) );
  nand_x1_sg U11180 ( .A(\reg_in[3][3][14] ), .B(n10479), .X(n8730) );
  nand_x1_sg U11181 ( .A(\in[3][3][15] ), .B(n10402), .X(n8727) );
  nand_x1_sg U11182 ( .A(\reg_in[3][3][15] ), .B(n10303), .X(n8728) );
  nand_x1_sg U11183 ( .A(\in[3][3][16] ), .B(n10311), .X(n8725) );
  nand_x1_sg U11184 ( .A(\reg_in[3][3][16] ), .B(n10478), .X(n8726) );
  nand_x1_sg U11185 ( .A(\in[3][3][17] ), .B(n10393), .X(n8723) );
  nand_x1_sg U11186 ( .A(\reg_in[3][3][17] ), .B(n10216), .X(n8724) );
  nand_x1_sg U11187 ( .A(\in[3][3][18] ), .B(n10600), .X(n8721) );
  nand_x1_sg U11188 ( .A(\reg_in[3][3][18] ), .B(n10192), .X(n8722) );
  nand_x1_sg U11189 ( .A(\in[3][3][19] ), .B(n10618), .X(n8717) );
  nand_x1_sg U11190 ( .A(\reg_in[3][3][19] ), .B(n10183), .X(n8718) );
  nand_x1_sg U11191 ( .A(\in[0][1][5] ), .B(n10327), .X(n9307) );
  nand_x1_sg U11192 ( .A(\reg_in[0][1][5] ), .B(n10306), .X(n9308) );
  nand_x1_sg U11193 ( .A(\in[0][1][6] ), .B(n10629), .X(n9305) );
  nand_x1_sg U11194 ( .A(\reg_in[0][1][6] ), .B(n10144), .X(n9306) );
  nand_x1_sg U11195 ( .A(\in[0][1][7] ), .B(n10630), .X(n9303) );
  nand_x1_sg U11196 ( .A(\reg_in[0][1][7] ), .B(n10535), .X(n9304) );
  nand_x1_sg U11197 ( .A(\in[0][1][8] ), .B(n10624), .X(n9301) );
  nand_x1_sg U11198 ( .A(\reg_in[0][1][8] ), .B(n10144), .X(n9302) );
  nand_x1_sg U11199 ( .A(\in[0][1][9] ), .B(n10326), .X(n9299) );
  nand_x1_sg U11200 ( .A(\reg_in[0][1][9] ), .B(n10525), .X(n9300) );
  nand_x1_sg U11201 ( .A(\in[0][2][15] ), .B(n10601), .X(n9247) );
  nand_x1_sg U11202 ( .A(\reg_in[0][2][15] ), .B(n10302), .X(n9248) );
  nand_x1_sg U11203 ( .A(\in[0][2][16] ), .B(n10399), .X(n9245) );
  nand_x1_sg U11204 ( .A(\reg_in[0][2][16] ), .B(n10058), .X(n9246) );
  nand_x1_sg U11205 ( .A(\in[0][2][17] ), .B(n10077), .X(n9243) );
  nand_x1_sg U11206 ( .A(\reg_in[0][2][17] ), .B(n10041), .X(n9244) );
  nand_x1_sg U11207 ( .A(\in[0][2][18] ), .B(n10604), .X(n9241) );
  nand_x1_sg U11208 ( .A(\reg_in[0][2][18] ), .B(n10539), .X(n9242) );
  nand_x1_sg U11209 ( .A(\in[0][2][19] ), .B(n10392), .X(n9239) );
  nand_x1_sg U11210 ( .A(\reg_in[0][2][19] ), .B(n10474), .X(n9240) );
  nand_x1_sg U11211 ( .A(\in[0][3][10] ), .B(n10389), .X(n9217) );
  nand_x1_sg U11212 ( .A(\reg_in[0][3][10] ), .B(n10523), .X(n9218) );
  nand_x1_sg U11213 ( .A(\in[0][3][11] ), .B(n10605), .X(n9215) );
  nand_x1_sg U11214 ( .A(\reg_in[0][3][11] ), .B(n10055), .X(n9216) );
  nand_x1_sg U11215 ( .A(\in[0][3][12] ), .B(n10079), .X(n9213) );
  nand_x1_sg U11216 ( .A(\reg_in[0][3][12] ), .B(n10211), .X(n9214) );
  nand_x1_sg U11217 ( .A(\in[0][3][13] ), .B(n10613), .X(n9211) );
  nand_x1_sg U11218 ( .A(\reg_in[0][3][13] ), .B(n10483), .X(n9212) );
  nand_x1_sg U11219 ( .A(\in[0][3][14] ), .B(n10084), .X(n9209) );
  nand_x1_sg U11220 ( .A(\reg_in[0][3][14] ), .B(n10214), .X(n9210) );
  nand_x1_sg U11221 ( .A(\in[1][0][5] ), .B(n10601), .X(n9187) );
  nand_x1_sg U11222 ( .A(\reg_in[1][0][5] ), .B(n10531), .X(n9188) );
  nand_x1_sg U11223 ( .A(\in[1][0][6] ), .B(n10083), .X(n9185) );
  nand_x1_sg U11224 ( .A(\reg_in[1][0][6] ), .B(n10522), .X(n9186) );
  nand_x1_sg U11225 ( .A(\in[1][0][7] ), .B(n10084), .X(n9183) );
  nand_x1_sg U11226 ( .A(\reg_in[1][0][7] ), .B(n10266), .X(n9184) );
  nand_x1_sg U11227 ( .A(\in[1][0][8] ), .B(n10335), .X(n9181) );
  nand_x1_sg U11228 ( .A(\reg_in[1][0][8] ), .B(n10059), .X(n9182) );
  nand_x1_sg U11229 ( .A(\in[1][0][9] ), .B(n10401), .X(n9179) );
  nand_x1_sg U11230 ( .A(\reg_in[1][0][9] ), .B(n10269), .X(n9180) );
  nand_x1_sg U11231 ( .A(\in[1][1][15] ), .B(n10080), .X(n9127) );
  nand_x1_sg U11232 ( .A(\reg_in[1][1][15] ), .B(n10529), .X(n9128) );
  nand_x1_sg U11233 ( .A(\in[1][1][16] ), .B(n10402), .X(n9125) );
  nand_x1_sg U11234 ( .A(\reg_in[1][1][16] ), .B(n10538), .X(n9126) );
  nand_x1_sg U11235 ( .A(\in[1][1][17] ), .B(n10086), .X(n9123) );
  nand_x1_sg U11236 ( .A(\reg_in[1][1][17] ), .B(n10212), .X(n9124) );
  nand_x1_sg U11237 ( .A(\in[1][1][18] ), .B(n10400), .X(n9121) );
  nand_x1_sg U11238 ( .A(\reg_in[1][1][18] ), .B(n10192), .X(n9122) );
  nand_x1_sg U11239 ( .A(\in[1][1][19] ), .B(n10316), .X(n9119) );
  nand_x1_sg U11240 ( .A(\reg_in[1][1][19] ), .B(n10529), .X(n9120) );
  nand_x1_sg U11241 ( .A(\in[1][3][10] ), .B(n10317), .X(n9057) );
  nand_x1_sg U11242 ( .A(\reg_in[1][3][10] ), .B(n10192), .X(n9058) );
  nand_x1_sg U11243 ( .A(\in[1][3][11] ), .B(n10401), .X(n9055) );
  nand_x1_sg U11244 ( .A(\reg_in[1][3][11] ), .B(n10141), .X(n9056) );
  nand_x1_sg U11245 ( .A(\in[1][3][12] ), .B(n10398), .X(n9053) );
  nand_x1_sg U11246 ( .A(\reg_in[1][3][12] ), .B(n10308), .X(n9054) );
  nand_x1_sg U11247 ( .A(\in[1][3][13] ), .B(n10336), .X(n9051) );
  nand_x1_sg U11248 ( .A(\reg_in[1][3][13] ), .B(n10570), .X(n9052) );
  nand_x1_sg U11249 ( .A(\in[1][3][14] ), .B(n10601), .X(n9049) );
  nand_x1_sg U11250 ( .A(\reg_in[1][3][14] ), .B(n10216), .X(n9050) );
  nand_x1_sg U11251 ( .A(\in[2][1][0] ), .B(n10394), .X(n8997) );
  nand_x1_sg U11252 ( .A(\reg_in[2][1][0] ), .B(n10042), .X(n8998) );
  nand_x1_sg U11253 ( .A(\in[2][1][1] ), .B(n10021), .X(n8995) );
  nand_x1_sg U11254 ( .A(\reg_in[2][1][1] ), .B(n10534), .X(n8996) );
  nand_x1_sg U11255 ( .A(\in[2][1][2] ), .B(n10616), .X(n8993) );
  nand_x1_sg U11256 ( .A(\reg_in[2][1][2] ), .B(n10265), .X(n8994) );
  nand_x1_sg U11257 ( .A(\in[2][1][3] ), .B(n10627), .X(n8991) );
  nand_x1_sg U11258 ( .A(\reg_in[2][1][3] ), .B(n10217), .X(n8992) );
  nand_x1_sg U11259 ( .A(\in[2][1][4] ), .B(n10619), .X(n8989) );
  nand_x1_sg U11260 ( .A(\reg_in[2][1][4] ), .B(n10477), .X(n8990) );
  nand_x1_sg U11261 ( .A(\in[2][1][15] ), .B(n10340), .X(n8967) );
  nand_x1_sg U11262 ( .A(\reg_in[2][1][15] ), .B(n10533), .X(n8968) );
  nand_x1_sg U11263 ( .A(\in[2][1][16] ), .B(n10339), .X(n8965) );
  nand_x1_sg U11264 ( .A(\reg_in[2][1][16] ), .B(n10145), .X(n8966) );
  nand_x1_sg U11265 ( .A(\in[2][1][17] ), .B(n10334), .X(n8963) );
  nand_x1_sg U11266 ( .A(\reg_in[2][1][17] ), .B(n10178), .X(n8964) );
  nand_x1_sg U11267 ( .A(\in[2][1][18] ), .B(n10338), .X(n8961) );
  nand_x1_sg U11268 ( .A(\reg_in[2][1][18] ), .B(n10570), .X(n8962) );
  nand_x1_sg U11269 ( .A(\in[2][1][19] ), .B(n10324), .X(n8959) );
  nand_x1_sg U11270 ( .A(\reg_in[2][1][19] ), .B(n10140), .X(n8960) );
  nand_x1_sg U11271 ( .A(\in[2][2][10] ), .B(n10603), .X(n8937) );
  nand_x1_sg U11272 ( .A(\reg_in[2][2][10] ), .B(n10528), .X(n8938) );
  nand_x1_sg U11273 ( .A(\in[2][2][11] ), .B(n10332), .X(n8935) );
  nand_x1_sg U11274 ( .A(\reg_in[2][2][11] ), .B(n10522), .X(n8936) );
  nand_x1_sg U11275 ( .A(\in[2][2][12] ), .B(n10612), .X(n8933) );
  nand_x1_sg U11276 ( .A(\reg_in[2][2][12] ), .B(n10288), .X(n8934) );
  nand_x1_sg U11277 ( .A(\in[2][2][13] ), .B(n10086), .X(n8931) );
  nand_x1_sg U11278 ( .A(\reg_in[2][2][13] ), .B(n10475), .X(n8932) );
  nand_x1_sg U11279 ( .A(\in[2][2][14] ), .B(n10338), .X(n8929) );
  nand_x1_sg U11280 ( .A(\reg_in[2][2][14] ), .B(n10060), .X(n8930) );
  nand_x1_sg U11281 ( .A(\in[3][0][0] ), .B(n10604), .X(n8877) );
  nand_x1_sg U11282 ( .A(\reg_in[3][0][0] ), .B(n10478), .X(n8878) );
  nand_x1_sg U11283 ( .A(\in[3][0][1] ), .B(n10328), .X(n8875) );
  nand_x1_sg U11284 ( .A(\reg_in[3][0][1] ), .B(n10308), .X(n8876) );
  nand_x1_sg U11285 ( .A(\in[3][0][2] ), .B(n10023), .X(n8873) );
  nand_x1_sg U11286 ( .A(\reg_in[3][0][2] ), .B(n10539), .X(n8874) );
  nand_x1_sg U11287 ( .A(\in[3][0][3] ), .B(n10632), .X(n8871) );
  nand_x1_sg U11288 ( .A(\reg_in[3][0][3] ), .B(n10303), .X(n8872) );
  nand_x1_sg U11289 ( .A(\in[3][0][4] ), .B(n10332), .X(n8869) );
  nand_x1_sg U11290 ( .A(\reg_in[3][0][4] ), .B(n10144), .X(n8870) );
  nand_x1_sg U11291 ( .A(\in[3][1][15] ), .B(n10339), .X(n8807) );
  nand_x1_sg U11292 ( .A(\reg_in[3][1][15] ), .B(n10528), .X(n8808) );
  nand_x1_sg U11293 ( .A(\in[3][1][16] ), .B(n10627), .X(n8805) );
  nand_x1_sg U11294 ( .A(\reg_in[3][1][16] ), .B(n10539), .X(n8806) );
  nand_x1_sg U11295 ( .A(\in[3][1][17] ), .B(n10390), .X(n8803) );
  nand_x1_sg U11296 ( .A(\reg_in[3][1][17] ), .B(n10056), .X(n8804) );
  nand_x1_sg U11297 ( .A(\in[3][1][18] ), .B(n10630), .X(n8801) );
  nand_x1_sg U11298 ( .A(\reg_in[3][1][18] ), .B(n10535), .X(n8802) );
  nand_x1_sg U11299 ( .A(\in[3][1][19] ), .B(n10619), .X(n8799) );
  nand_x1_sg U11300 ( .A(\reg_in[3][1][19] ), .B(n10541), .X(n8800) );
  nand_x1_sg U11301 ( .A(\in[3][3][5] ), .B(n10608), .X(n8747) );
  nand_x1_sg U11302 ( .A(\reg_in[3][3][5] ), .B(n10571), .X(n8748) );
  nand_x1_sg U11303 ( .A(\in[3][3][6] ), .B(n10334), .X(n8745) );
  nand_x1_sg U11304 ( .A(\reg_in[3][3][6] ), .B(n10184), .X(n8746) );
  nand_x1_sg U11305 ( .A(\in[3][3][7] ), .B(n10258), .X(n8743) );
  nand_x1_sg U11306 ( .A(\reg_in[3][3][7] ), .B(n10483), .X(n8744) );
  nand_x1_sg U11307 ( .A(\in[3][3][8] ), .B(n10395), .X(n8741) );
  nand_x1_sg U11308 ( .A(\reg_in[3][3][8] ), .B(n10214), .X(n8742) );
  nand_x1_sg U11309 ( .A(\in[3][3][9] ), .B(n10408), .X(n8739) );
  nand_x1_sg U11310 ( .A(\reg_in[3][3][9] ), .B(n10265), .X(n8740) );
  nor_x1_sg U11311 ( .A(\reg_in[0][0][9] ), .B(n10445), .X(n3511) );
  nor_x1_sg U11312 ( .A(\reg_in[0][0][12] ), .B(n10121), .X(n3499) );
  nor_x1_sg U11313 ( .A(\reg_in[0][0][15] ), .B(n10634), .X(n3487) );
  nor_x1_sg U11314 ( .A(\reg_in[0][0][18] ), .B(n10454), .X(n3475) );
  nor_x1_sg U11315 ( .A(\reg_in[1][0][1] ), .B(n10126), .X(n3463) );
  nor_x1_sg U11316 ( .A(\reg_in[1][0][4] ), .B(n10279), .X(n3451) );
  nor_x1_sg U11317 ( .A(\reg_in[1][0][9] ), .B(n10127), .X(n3431) );
  nor_x1_sg U11318 ( .A(\reg_in[1][0][12] ), .B(n10036), .X(n3419) );
  nor_x1_sg U11319 ( .A(\reg_in[1][0][15] ), .B(n10063), .X(n3407) );
  nor_x1_sg U11320 ( .A(\reg_in[1][0][18] ), .B(n10494), .X(n3395) );
  nor_x1_sg U11321 ( .A(\reg_in[2][0][1] ), .B(n10555), .X(n3383) );
  nor_x1_sg U11322 ( .A(\reg_in[2][0][4] ), .B(n10446), .X(n3371) );
  nor_x1_sg U11323 ( .A(\reg_in[2][0][7] ), .B(n10447), .X(n3359) );
  nor_x1_sg U11324 ( .A(\reg_in[2][0][10] ), .B(n10446), .X(n3347) );
  nor_x1_sg U11325 ( .A(\reg_in[2][0][13] ), .B(n10500), .X(n3335) );
  nor_x1_sg U11326 ( .A(\reg_in[2][0][16] ), .B(n10547), .X(n3323) );
  nor_x1_sg U11327 ( .A(\reg_in[2][0][19] ), .B(n10436), .X(n3311) );
  nor_x1_sg U11328 ( .A(\reg_in[3][0][2] ), .B(n10063), .X(n3299) );
  nor_x1_sg U11329 ( .A(\reg_in[3][0][5] ), .B(n10457), .X(n3287) );
  nor_x1_sg U11330 ( .A(\reg_in[3][0][8] ), .B(n10292), .X(n3275) );
  nor_x1_sg U11331 ( .A(\reg_in[3][0][11] ), .B(n10151), .X(n3263) );
  nor_x1_sg U11332 ( .A(\reg_in[3][0][14] ), .B(n10033), .X(n3251) );
  nor_x1_sg U11333 ( .A(\reg_in[3][0][17] ), .B(n10495), .X(n3239) );
  nor_x1_sg U11334 ( .A(\reg_in[0][1][0] ), .B(n10242), .X(n3227) );
  nor_x1_sg U11335 ( .A(\reg_in[0][1][3] ), .B(n10501), .X(n3215) );
  nor_x1_sg U11336 ( .A(\reg_in[0][1][6] ), .B(n10459), .X(n3203) );
  nor_x1_sg U11337 ( .A(\reg_in[0][1][9] ), .B(n10456), .X(n3191) );
  nor_x1_sg U11338 ( .A(\reg_in[0][1][12] ), .B(n10157), .X(n3179) );
  nor_x1_sg U11339 ( .A(\reg_in[0][1][15] ), .B(n10550), .X(n3167) );
  nor_x1_sg U11340 ( .A(\reg_in[0][1][18] ), .B(n10495), .X(n3155) );
  nor_x1_sg U11341 ( .A(\reg_in[1][1][1] ), .B(n10453), .X(n3143) );
  nor_x1_sg U11342 ( .A(\reg_in[1][1][4] ), .B(n10497), .X(n3131) );
  nor_x1_sg U11343 ( .A(\reg_in[1][1][7] ), .B(n10121), .X(n3119) );
  nor_x1_sg U11344 ( .A(\reg_in[1][1][10] ), .B(n10246), .X(n3107) );
  nor_x1_sg U11345 ( .A(\reg_in[1][1][13] ), .B(n10247), .X(n3095) );
  nor_x1_sg U11346 ( .A(\reg_in[1][1][16] ), .B(n10456), .X(n3083) );
  nor_x1_sg U11347 ( .A(\reg_in[1][1][19] ), .B(n10018), .X(n3071) );
  nor_x1_sg U11348 ( .A(\reg_in[2][1][2] ), .B(n10291), .X(n3059) );
  nor_x1_sg U11349 ( .A(\reg_in[2][1][5] ), .B(n10491), .X(n3047) );
  nor_x1_sg U11350 ( .A(\reg_in[2][1][8] ), .B(n10045), .X(n3035) );
  nor_x1_sg U11351 ( .A(\reg_in[2][1][11] ), .B(n10553), .X(n3023) );
  nor_x1_sg U11352 ( .A(\reg_in[2][1][14] ), .B(n10278), .X(n3011) );
  nor_x1_sg U11353 ( .A(\reg_in[2][1][17] ), .B(n10455), .X(n2999) );
  nor_x1_sg U11354 ( .A(\reg_in[3][1][0] ), .B(n10127), .X(n2987) );
  nor_x1_sg U11355 ( .A(\reg_in[3][1][3] ), .B(n10548), .X(n2975) );
  nor_x1_sg U11356 ( .A(\reg_in[3][1][6] ), .B(n10228), .X(n2963) );
  nor_x1_sg U11357 ( .A(\reg_in[3][1][9] ), .B(n10634), .X(n2951) );
  nor_x1_sg U11358 ( .A(\reg_in[3][1][12] ), .B(n10447), .X(n2939) );
  nor_x1_sg U11359 ( .A(\reg_in[3][1][15] ), .B(n10114), .X(n2927) );
  nor_x1_sg U11360 ( .A(\reg_in[3][1][16] ), .B(n10495), .X(n2923) );
  nor_x1_sg U11361 ( .A(\reg_in[3][1][19] ), .B(n10279), .X(n2911) );
  nor_x1_sg U11362 ( .A(\reg_in[0][2][2] ), .B(n10445), .X(n2899) );
  nor_x1_sg U11363 ( .A(\reg_in[0][2][5] ), .B(n10440), .X(n2887) );
  nor_x1_sg U11364 ( .A(\reg_in[0][2][8] ), .B(n10152), .X(n2875) );
  nor_x1_sg U11365 ( .A(\reg_in[0][2][11] ), .B(n10439), .X(n2863) );
  nor_x1_sg U11366 ( .A(\reg_in[0][2][14] ), .B(n10555), .X(n2851) );
  nor_x1_sg U11367 ( .A(\reg_in[0][2][17] ), .B(n10033), .X(n2839) );
  nor_x1_sg U11368 ( .A(\reg_in[1][2][0] ), .B(n10501), .X(n2827) );
  nor_x1_sg U11369 ( .A(\reg_in[1][2][3] ), .B(n10122), .X(n2815) );
  nor_x1_sg U11370 ( .A(\reg_in[1][2][6] ), .B(n10036), .X(n2803) );
  nor_x1_sg U11371 ( .A(\reg_in[1][2][9] ), .B(n10502), .X(n2791) );
  nor_x1_sg U11372 ( .A(\reg_in[1][2][12] ), .B(n10442), .X(n2779) );
  nor_x1_sg U11373 ( .A(\reg_in[1][2][15] ), .B(n10291), .X(n2767) );
  nor_x1_sg U11374 ( .A(\reg_in[1][2][18] ), .B(n10062), .X(n2755) );
  nor_x1_sg U11375 ( .A(\reg_in[2][2][1] ), .B(n10449), .X(n2743) );
  nor_x1_sg U11376 ( .A(\reg_in[2][2][4] ), .B(n10066), .X(n2731) );
  nor_x1_sg U11377 ( .A(\reg_in[2][2][7] ), .B(n10205), .X(n2719) );
  nor_x1_sg U11378 ( .A(\reg_in[2][2][10] ), .B(n10451), .X(n2707) );
  nor_x1_sg U11379 ( .A(\reg_in[2][2][13] ), .B(n10264), .X(n2695) );
  nor_x1_sg U11380 ( .A(\reg_in[2][2][16] ), .B(n10046), .X(n2683) );
  nor_x1_sg U11381 ( .A(\reg_in[2][2][19] ), .B(n10553), .X(n2671) );
  nor_x1_sg U11382 ( .A(\reg_in[3][2][2] ), .B(n10442), .X(n2659) );
  nor_x1_sg U11383 ( .A(\reg_in[3][2][5] ), .B(n10292), .X(n2647) );
  nor_x1_sg U11384 ( .A(\reg_in[3][2][8] ), .B(n10457), .X(n2635) );
  nor_x1_sg U11385 ( .A(\reg_in[3][2][11] ), .B(n10459), .X(n2623) );
  nor_x1_sg U11386 ( .A(\reg_in[3][2][14] ), .B(n10456), .X(n2611) );
  nor_x1_sg U11387 ( .A(\reg_in[3][2][17] ), .B(n10241), .X(n2599) );
  nor_x1_sg U11388 ( .A(\reg_in[0][3][0] ), .B(n10027), .X(n2587) );
  nor_x1_sg U11389 ( .A(\reg_in[0][3][3] ), .B(n10437), .X(n2575) );
  nor_x1_sg U11390 ( .A(\reg_in[0][3][6] ), .B(n10121), .X(n2563) );
  nor_x1_sg U11391 ( .A(\reg_in[0][3][9] ), .B(n10151), .X(n2551) );
  nor_x1_sg U11392 ( .A(\reg_in[0][3][12] ), .B(n10126), .X(n2539) );
  nor_x1_sg U11393 ( .A(\reg_in[0][3][15] ), .B(n10497), .X(n2527) );
  nor_x1_sg U11394 ( .A(\reg_in[0][3][18] ), .B(n10458), .X(n2515) );
  nor_x1_sg U11395 ( .A(\reg_in[1][3][1] ), .B(n10122), .X(n2503) );
  nor_x1_sg U11396 ( .A(\reg_in[1][3][4] ), .B(n10437), .X(n2491) );
  nor_x1_sg U11397 ( .A(\reg_in[1][3][7] ), .B(n10547), .X(n2479) );
  nor_x1_sg U11398 ( .A(\reg_in[1][3][10] ), .B(n10634), .X(n2467) );
  nor_x1_sg U11399 ( .A(\reg_in[1][3][13] ), .B(n10636), .X(n2455) );
  nor_x1_sg U11400 ( .A(\reg_in[1][3][16] ), .B(n10157), .X(n2443) );
  nor_x1_sg U11401 ( .A(\reg_in[1][3][19] ), .B(n10004), .X(n2431) );
  nor_x1_sg U11402 ( .A(\reg_in[2][3][2] ), .B(n10278), .X(n2419) );
  nor_x1_sg U11403 ( .A(\reg_in[2][3][5] ), .B(n10088), .X(n2407) );
  nor_x1_sg U11404 ( .A(\reg_in[2][3][8] ), .B(n10550), .X(n2395) );
  nor_x1_sg U11405 ( .A(\reg_in[2][3][11] ), .B(n10501), .X(n2383) );
  nor_x1_sg U11406 ( .A(\reg_in[2][3][14] ), .B(n10449), .X(n2371) );
  nor_x1_sg U11407 ( .A(\reg_in[2][3][17] ), .B(n10448), .X(n2359) );
  nor_x1_sg U11408 ( .A(\reg_in[3][3][0] ), .B(n10499), .X(n2347) );
  nor_x1_sg U11409 ( .A(\reg_in[3][3][3] ), .B(n10263), .X(n2335) );
  nor_x1_sg U11410 ( .A(\reg_in[3][3][6] ), .B(n10494), .X(n2323) );
  nor_x1_sg U11411 ( .A(\reg_in[3][3][9] ), .B(n10460), .X(n2311) );
  nor_x1_sg U11412 ( .A(\reg_in[3][3][12] ), .B(n10280), .X(n2299) );
  nor_x1_sg U11413 ( .A(\reg_in[3][3][15] ), .B(n10201), .X(n2287) );
  nor_x1_sg U11414 ( .A(\reg_in[3][3][18] ), .B(n10264), .X(n2275) );
  nor_x1_sg U11415 ( .A(\reg_in[0][0][0] ), .B(n10449), .X(n2267) );
  nor_x1_sg U11416 ( .A(\reg_in[0][0][1] ), .B(n10156), .X(n3543) );
  nor_x1_sg U11417 ( .A(\reg_in[0][0][2] ), .B(n10636), .X(n3539) );
  nor_x1_sg U11418 ( .A(\reg_in[0][0][3] ), .B(n10018), .X(n3535) );
  nor_x1_sg U11419 ( .A(\reg_in[0][0][4] ), .B(n10277), .X(n3531) );
  nor_x1_sg U11420 ( .A(\reg_in[0][0][5] ), .B(n10556), .X(n3527) );
  nor_x1_sg U11421 ( .A(\reg_in[0][0][6] ), .B(n10263), .X(n3523) );
  nor_x1_sg U11422 ( .A(\reg_in[0][0][7] ), .B(n10492), .X(n3519) );
  nor_x1_sg U11423 ( .A(\reg_in[0][0][8] ), .B(n10280), .X(n3515) );
  nor_x1_sg U11424 ( .A(\reg_in[0][0][10] ), .B(n10290), .X(n3507) );
  nor_x1_sg U11425 ( .A(\reg_in[0][0][11] ), .B(n10453), .X(n3503) );
  nor_x1_sg U11426 ( .A(\reg_in[0][0][13] ), .B(n10004), .X(n3495) );
  nor_x1_sg U11427 ( .A(\reg_in[0][0][14] ), .B(n10458), .X(n3491) );
  nor_x1_sg U11428 ( .A(\reg_in[0][0][16] ), .B(n10045), .X(n3483) );
  nor_x1_sg U11429 ( .A(\reg_in[0][0][17] ), .B(n10114), .X(n3479) );
  nor_x1_sg U11430 ( .A(\reg_in[0][0][19] ), .B(n10548), .X(n3471) );
  nor_x1_sg U11431 ( .A(\reg_in[1][0][0] ), .B(n10445), .X(n3467) );
  nor_x1_sg U11432 ( .A(\reg_in[1][0][2] ), .B(n10202), .X(n3459) );
  nor_x1_sg U11433 ( .A(\reg_in[1][0][3] ), .B(n10444), .X(n3455) );
  nor_x1_sg U11434 ( .A(\reg_in[1][0][5] ), .B(n10444), .X(n3447) );
  nor_x1_sg U11435 ( .A(\reg_in[1][0][6] ), .B(n10554), .X(n3443) );
  nor_x1_sg U11436 ( .A(\reg_in[1][0][7] ), .B(n10241), .X(n3439) );
  nor_x1_sg U11437 ( .A(\reg_in[1][0][8] ), .B(n10546), .X(n3435) );
  nor_x1_sg U11438 ( .A(\reg_in[1][0][10] ), .B(n10152), .X(n3427) );
  nor_x1_sg U11439 ( .A(\reg_in[1][0][11] ), .B(n10110), .X(n3423) );
  nor_x1_sg U11440 ( .A(\reg_in[1][0][13] ), .B(n10151), .X(n3415) );
  nor_x1_sg U11441 ( .A(\reg_in[1][0][14] ), .B(n10201), .X(n3411) );
  nor_x1_sg U11442 ( .A(\reg_in[1][0][16] ), .B(n10019), .X(n3403) );
  nor_x1_sg U11443 ( .A(\reg_in[1][0][17] ), .B(n10118), .X(n3399) );
  nor_x1_sg U11444 ( .A(\reg_in[1][0][19] ), .B(n10206), .X(n3391) );
  nor_x1_sg U11445 ( .A(\reg_in[2][0][0] ), .B(n10458), .X(n3387) );
  nor_x1_sg U11446 ( .A(\reg_in[2][0][2] ), .B(n10045), .X(n3379) );
  nor_x1_sg U11447 ( .A(\reg_in[2][0][3] ), .B(n10460), .X(n3375) );
  nor_x1_sg U11448 ( .A(\reg_in[2][0][5] ), .B(n10263), .X(n3367) );
  nor_x1_sg U11449 ( .A(\reg_in[2][0][6] ), .B(n10459), .X(n3363) );
  nor_x1_sg U11450 ( .A(\reg_in[2][0][8] ), .B(n10121), .X(n3355) );
  nor_x1_sg U11451 ( .A(\reg_in[2][0][9] ), .B(n10126), .X(n3351) );
  nor_x1_sg U11452 ( .A(\reg_in[2][0][11] ), .B(n10455), .X(n3343) );
  nor_x1_sg U11453 ( .A(\reg_in[2][0][12] ), .B(n10546), .X(n3339) );
  nor_x1_sg U11454 ( .A(\reg_in[2][0][14] ), .B(n10555), .X(n3331) );
  nor_x1_sg U11455 ( .A(\reg_in[2][0][15] ), .B(n10152), .X(n3327) );
  nor_x1_sg U11456 ( .A(\reg_in[2][0][17] ), .B(n10227), .X(n3319) );
  nor_x1_sg U11457 ( .A(\reg_in[2][0][18] ), .B(n10290), .X(n3315) );
  nor_x1_sg U11458 ( .A(\reg_in[3][0][0] ), .B(n10441), .X(n3307) );
  nor_x1_sg U11459 ( .A(\reg_in[3][0][1] ), .B(n10037), .X(n3303) );
  nor_x1_sg U11460 ( .A(\reg_in[3][0][3] ), .B(n10446), .X(n3295) );
  nor_x1_sg U11461 ( .A(\reg_in[3][0][4] ), .B(n10439), .X(n3291) );
  nor_x1_sg U11462 ( .A(\reg_in[3][0][6] ), .B(n10450), .X(n3283) );
  nor_x1_sg U11463 ( .A(\reg_in[3][0][7] ), .B(n10279), .X(n3279) );
  nor_x1_sg U11464 ( .A(\reg_in[3][0][9] ), .B(n10206), .X(n3271) );
  nor_x1_sg U11465 ( .A(\reg_in[3][0][10] ), .B(n10446), .X(n3267) );
  nor_x1_sg U11466 ( .A(\reg_in[3][0][12] ), .B(n10448), .X(n3259) );
  nor_x1_sg U11467 ( .A(\reg_in[3][0][13] ), .B(n10046), .X(n3255) );
  nor_x1_sg U11468 ( .A(\reg_in[3][0][15] ), .B(n10242), .X(n3247) );
  nor_x1_sg U11469 ( .A(\reg_in[3][0][16] ), .B(n10491), .X(n3243) );
  nor_x1_sg U11470 ( .A(\reg_in[3][0][18] ), .B(n10440), .X(n3235) );
  nor_x1_sg U11471 ( .A(\reg_in[3][0][19] ), .B(n10494), .X(n3231) );
  nor_x1_sg U11472 ( .A(\reg_in[0][1][1] ), .B(n10292), .X(n3223) );
  nor_x1_sg U11473 ( .A(\reg_in[0][1][2] ), .B(n10436), .X(n3219) );
  nor_x1_sg U11474 ( .A(\reg_in[0][1][4] ), .B(n10441), .X(n3211) );
  nor_x1_sg U11475 ( .A(\reg_in[0][1][5] ), .B(n10246), .X(n3207) );
  nor_x1_sg U11476 ( .A(\reg_in[0][1][7] ), .B(n10636), .X(n3199) );
  nor_x1_sg U11477 ( .A(\reg_in[0][1][8] ), .B(n10247), .X(n3195) );
  nor_x1_sg U11478 ( .A(\reg_in[0][1][10] ), .B(n10496), .X(n3187) );
  nor_x1_sg U11479 ( .A(\reg_in[0][1][11] ), .B(n10034), .X(n3183) );
  nor_x1_sg U11480 ( .A(\reg_in[0][1][13] ), .B(n10436), .X(n3175) );
  nor_x1_sg U11481 ( .A(\reg_in[0][1][14] ), .B(n10122), .X(n3171) );
  nor_x1_sg U11482 ( .A(\reg_in[0][1][16] ), .B(n10440), .X(n3163) );
  nor_x1_sg U11483 ( .A(\reg_in[0][1][17] ), .B(n10439), .X(n3159) );
  nor_x1_sg U11484 ( .A(\reg_in[0][1][19] ), .B(n10447), .X(n3151) );
  nor_x1_sg U11485 ( .A(\reg_in[1][1][0] ), .B(n10552), .X(n3147) );
  nor_x1_sg U11486 ( .A(\reg_in[1][1][2] ), .B(n10460), .X(n3139) );
  nor_x1_sg U11487 ( .A(\reg_in[1][1][3] ), .B(n10448), .X(n3135) );
  nor_x1_sg U11488 ( .A(\reg_in[1][1][5] ), .B(n10549), .X(n3127) );
  nor_x1_sg U11489 ( .A(\reg_in[1][1][6] ), .B(n10496), .X(n3123) );
  nor_x1_sg U11490 ( .A(\reg_in[1][1][8] ), .B(n10227), .X(n3115) );
  nor_x1_sg U11491 ( .A(\reg_in[1][1][9] ), .B(n10554), .X(n3111) );
  nor_x1_sg U11492 ( .A(\reg_in[1][1][11] ), .B(n10228), .X(n3103) );
  nor_x1_sg U11493 ( .A(\reg_in[1][1][12] ), .B(n10264), .X(n3099) );
  nor_x1_sg U11494 ( .A(\reg_in[1][1][14] ), .B(n10112), .X(n3091) );
  nor_x1_sg U11495 ( .A(\reg_in[1][1][15] ), .B(n10556), .X(n3087) );
  nor_x1_sg U11496 ( .A(\reg_in[1][1][17] ), .B(n10547), .X(n3079) );
  nor_x1_sg U11497 ( .A(\reg_in[1][1][18] ), .B(n10263), .X(n3075) );
  nor_x1_sg U11498 ( .A(\reg_in[2][1][0] ), .B(n10549), .X(n3067) );
  nor_x1_sg U11499 ( .A(\reg_in[2][1][1] ), .B(n10499), .X(n3063) );
  nor_x1_sg U11500 ( .A(\reg_in[2][1][3] ), .B(n10062), .X(n3055) );
  nor_x1_sg U11501 ( .A(\reg_in[2][1][4] ), .B(n10127), .X(n3051) );
  nor_x1_sg U11502 ( .A(\reg_in[2][1][6] ), .B(n10552), .X(n3043) );
  nor_x1_sg U11503 ( .A(\reg_in[2][1][7] ), .B(n10153), .X(n3039) );
  nor_x1_sg U11504 ( .A(\reg_in[2][1][9] ), .B(n10494), .X(n3031) );
  nor_x1_sg U11505 ( .A(\reg_in[2][1][10] ), .B(n10156), .X(n3027) );
  nor_x1_sg U11506 ( .A(\reg_in[2][1][12] ), .B(n10156), .X(n3019) );
  nor_x1_sg U11507 ( .A(\reg_in[2][1][13] ), .B(n10548), .X(n3015) );
  nor_x1_sg U11508 ( .A(\reg_in[2][1][15] ), .B(n10450), .X(n3007) );
  nor_x1_sg U11509 ( .A(\reg_in[2][1][16] ), .B(n10291), .X(n3003) );
  nor_x1_sg U11510 ( .A(\reg_in[2][1][18] ), .B(n10241), .X(n2995) );
  nor_x1_sg U11511 ( .A(\reg_in[2][1][19] ), .B(n10157), .X(n2991) );
  nor_x1_sg U11512 ( .A(\reg_in[3][1][1] ), .B(n10046), .X(n2983) );
  nor_x1_sg U11513 ( .A(\reg_in[3][1][2] ), .B(n10457), .X(n2979) );
  nor_x1_sg U11514 ( .A(\reg_in[3][1][4] ), .B(n10457), .X(n2971) );
  nor_x1_sg U11515 ( .A(\reg_in[3][1][5] ), .B(n10500), .X(n2967) );
  nor_x1_sg U11516 ( .A(\reg_in[3][1][7] ), .B(n10151), .X(n2959) );
  nor_x1_sg U11517 ( .A(\reg_in[3][1][8] ), .B(n10278), .X(n2955) );
  nor_x1_sg U11518 ( .A(\reg_in[3][1][10] ), .B(n10453), .X(n2947) );
  nor_x1_sg U11519 ( .A(\reg_in[3][1][11] ), .B(n10205), .X(n2943) );
  nor_x1_sg U11520 ( .A(\reg_in[3][1][13] ), .B(n10278), .X(n2935) );
  nor_x1_sg U11521 ( .A(\reg_in[3][1][14] ), .B(n10242), .X(n2931) );
  nor_x1_sg U11522 ( .A(\reg_in[3][1][17] ), .B(n10206), .X(n2919) );
  nor_x1_sg U11523 ( .A(\reg_in[3][1][18] ), .B(n10227), .X(n2915) );
  nor_x1_sg U11524 ( .A(\reg_in[0][2][0] ), .B(n10064), .X(n2907) );
  nor_x1_sg U11525 ( .A(\reg_in[0][2][1] ), .B(n10497), .X(n2903) );
  nor_x1_sg U11526 ( .A(\reg_in[0][2][3] ), .B(n10441), .X(n2895) );
  nor_x1_sg U11527 ( .A(\reg_in[0][2][4] ), .B(n10264), .X(n2891) );
  nor_x1_sg U11528 ( .A(\reg_in[0][2][6] ), .B(n10064), .X(n2883) );
  nor_x1_sg U11529 ( .A(\reg_in[0][2][7] ), .B(n10450), .X(n2879) );
  nor_x1_sg U11530 ( .A(\reg_in[0][2][9] ), .B(n10451), .X(n2871) );
  nor_x1_sg U11531 ( .A(\reg_in[0][2][10] ), .B(n10460), .X(n2867) );
  nor_x1_sg U11532 ( .A(\reg_in[0][2][12] ), .B(n10492), .X(n2859) );
  nor_x1_sg U11533 ( .A(\reg_in[0][2][13] ), .B(n10551), .X(n2855) );
  nor_x1_sg U11534 ( .A(\reg_in[0][2][15] ), .B(n10556), .X(n2847) );
  nor_x1_sg U11535 ( .A(\reg_in[0][2][16] ), .B(n10441), .X(n2843) );
  nor_x1_sg U11536 ( .A(\reg_in[0][2][18] ), .B(n10437), .X(n2835) );
  nor_x1_sg U11537 ( .A(\reg_in[0][2][19] ), .B(n10499), .X(n2831) );
  nor_x1_sg U11538 ( .A(\reg_in[1][2][1] ), .B(n10202), .X(n2823) );
  nor_x1_sg U11539 ( .A(\reg_in[1][2][2] ), .B(n10037), .X(n2819) );
  nor_x1_sg U11540 ( .A(\reg_in[1][2][4] ), .B(n10551), .X(n2811) );
  nor_x1_sg U11541 ( .A(\reg_in[1][2][5] ), .B(n10290), .X(n2807) );
  nor_x1_sg U11542 ( .A(\reg_in[1][2][7] ), .B(n10549), .X(n2799) );
  nor_x1_sg U11543 ( .A(\reg_in[1][2][8] ), .B(n10549), .X(n2795) );
  nor_x1_sg U11544 ( .A(\reg_in[1][2][10] ), .B(n10459), .X(n2787) );
  nor_x1_sg U11545 ( .A(\reg_in[1][2][11] ), .B(n10491), .X(n2783) );
  nor_x1_sg U11546 ( .A(\reg_in[1][2][13] ), .B(n10450), .X(n2775) );
  nor_x1_sg U11547 ( .A(\reg_in[1][2][14] ), .B(n10228), .X(n2771) );
  nor_x1_sg U11548 ( .A(\reg_in[1][2][16] ), .B(n10552), .X(n2763) );
  nor_x1_sg U11549 ( .A(\reg_in[1][2][17] ), .B(n10440), .X(n2759) );
  nor_x1_sg U11550 ( .A(\reg_in[1][2][19] ), .B(n10206), .X(n2751) );
  nor_x1_sg U11551 ( .A(\reg_in[2][2][0] ), .B(n10126), .X(n2747) );
  nor_x1_sg U11552 ( .A(\reg_in[2][2][2] ), .B(n10437), .X(n2739) );
  nor_x1_sg U11553 ( .A(\reg_in[2][2][3] ), .B(n10496), .X(n2735) );
  nor_x1_sg U11554 ( .A(\reg_in[2][2][5] ), .B(n10501), .X(n2727) );
  nor_x1_sg U11555 ( .A(\reg_in[2][2][6] ), .B(n10018), .X(n2723) );
  nor_x1_sg U11556 ( .A(\reg_in[2][2][8] ), .B(n10497), .X(n2715) );
  nor_x1_sg U11557 ( .A(\reg_in[2][2][9] ), .B(n10088), .X(n2711) );
  nor_x1_sg U11558 ( .A(\reg_in[2][2][11] ), .B(n10554), .X(n2703) );
  nor_x1_sg U11559 ( .A(\reg_in[2][2][12] ), .B(n10066), .X(n2699) );
  nor_x1_sg U11560 ( .A(\reg_in[2][2][14] ), .B(n10292), .X(n2691) );
  nor_x1_sg U11561 ( .A(\reg_in[2][2][15] ), .B(n10449), .X(n2687) );
  nor_x1_sg U11562 ( .A(\reg_in[2][2][17] ), .B(n10492), .X(n2679) );
  nor_x1_sg U11563 ( .A(\reg_in[2][2][18] ), .B(n10037), .X(n2675) );
  nor_x1_sg U11564 ( .A(\reg_in[3][2][0] ), .B(n10555), .X(n2667) );
  nor_x1_sg U11565 ( .A(\reg_in[3][2][1] ), .B(n10280), .X(n2663) );
  nor_x1_sg U11566 ( .A(\reg_in[3][2][3] ), .B(n10063), .X(n2655) );
  nor_x1_sg U11567 ( .A(\reg_in[3][2][4] ), .B(n10228), .X(n2651) );
  nor_x1_sg U11568 ( .A(\reg_in[3][2][6] ), .B(n10451), .X(n2643) );
  nor_x1_sg U11569 ( .A(\reg_in[3][2][7] ), .B(n10454), .X(n2639) );
  nor_x1_sg U11570 ( .A(\reg_in[3][2][9] ), .B(n10551), .X(n2631) );
  nor_x1_sg U11571 ( .A(\reg_in[3][2][10] ), .B(n10156), .X(n2627) );
  nor_x1_sg U11572 ( .A(\reg_in[3][2][12] ), .B(n10033), .X(n2619) );
  nor_x1_sg U11573 ( .A(\reg_in[3][2][13] ), .B(n10019), .X(n2615) );
  nor_x1_sg U11574 ( .A(\reg_in[3][2][15] ), .B(n10202), .X(n2607) );
  nor_x1_sg U11575 ( .A(\reg_in[3][2][16] ), .B(n10277), .X(n2603) );
  nor_x1_sg U11576 ( .A(\reg_in[3][2][18] ), .B(n10246), .X(n2595) );
  nor_x1_sg U11577 ( .A(\reg_in[3][2][19] ), .B(n10241), .X(n2591) );
  nor_x1_sg U11578 ( .A(\reg_in[0][3][1] ), .B(n10550), .X(n2583) );
  nor_x1_sg U11579 ( .A(\reg_in[0][3][2] ), .B(n10201), .X(n2579) );
  nor_x1_sg U11580 ( .A(\reg_in[0][3][4] ), .B(n10068), .X(n2571) );
  nor_x1_sg U11581 ( .A(\reg_in[0][3][5] ), .B(n10062), .X(n2567) );
  nor_x1_sg U11582 ( .A(\reg_in[0][3][7] ), .B(n10502), .X(n2559) );
  nor_x1_sg U11583 ( .A(\reg_in[0][3][8] ), .B(n10455), .X(n2555) );
  nor_x1_sg U11584 ( .A(\reg_in[0][3][10] ), .B(n10499), .X(n2547) );
  nor_x1_sg U11585 ( .A(\reg_in[0][3][11] ), .B(n10436), .X(n2543) );
  nor_x1_sg U11586 ( .A(\reg_in[0][3][13] ), .B(n10551), .X(n2535) );
  nor_x1_sg U11587 ( .A(\reg_in[0][3][14] ), .B(n10447), .X(n2531) );
  nor_x1_sg U11588 ( .A(\reg_in[0][3][16] ), .B(n10442), .X(n2523) );
  nor_x1_sg U11589 ( .A(\reg_in[0][3][17] ), .B(n10152), .X(n2519) );
  nor_x1_sg U11590 ( .A(\reg_in[0][3][19] ), .B(n10564), .X(n2511) );
  nor_x1_sg U11591 ( .A(\reg_in[1][3][0] ), .B(n10205), .X(n2507) );
  nor_x1_sg U11592 ( .A(\reg_in[1][3][2] ), .B(n10242), .X(n2499) );
  nor_x1_sg U11593 ( .A(\reg_in[1][3][3] ), .B(n10455), .X(n2495) );
  nor_x1_sg U11594 ( .A(\reg_in[1][3][5] ), .B(n10502), .X(n2487) );
  nor_x1_sg U11595 ( .A(\reg_in[1][3][6] ), .B(n10277), .X(n2483) );
  nor_x1_sg U11596 ( .A(\reg_in[1][3][8] ), .B(n10157), .X(n2475) );
  nor_x1_sg U11597 ( .A(\reg_in[1][3][9] ), .B(n10556), .X(n2471) );
  nor_x1_sg U11598 ( .A(\reg_in[1][3][11] ), .B(n10448), .X(n2463) );
  nor_x1_sg U11599 ( .A(\reg_in[1][3][12] ), .B(n10439), .X(n2459) );
  nor_x1_sg U11600 ( .A(\reg_in[1][3][14] ), .B(n10454), .X(n2451) );
  nor_x1_sg U11601 ( .A(\reg_in[1][3][15] ), .B(n10064), .X(n2447) );
  nor_x1_sg U11602 ( .A(\reg_in[1][3][17] ), .B(n10445), .X(n2439) );
  nor_x1_sg U11603 ( .A(\reg_in[1][3][18] ), .B(n10088), .X(n2435) );
  nor_x1_sg U11604 ( .A(\reg_in[2][3][0] ), .B(n10442), .X(n2427) );
  nor_x1_sg U11605 ( .A(\reg_in[2][3][1] ), .B(n10635), .X(n2423) );
  nor_x1_sg U11606 ( .A(\reg_in[2][3][3] ), .B(n10414), .X(n2415) );
  nor_x1_sg U11607 ( .A(\reg_in[2][3][4] ), .B(n10502), .X(n2411) );
  nor_x1_sg U11608 ( .A(\reg_in[2][3][6] ), .B(n10635), .X(n2403) );
  nor_x1_sg U11609 ( .A(\reg_in[2][3][7] ), .B(n10451), .X(n2399) );
  nor_x1_sg U11610 ( .A(\reg_in[2][3][9] ), .B(n10247), .X(n2391) );
  nor_x1_sg U11611 ( .A(\reg_in[2][3][10] ), .B(n10453), .X(n2387) );
  nor_x1_sg U11612 ( .A(\reg_in[2][3][12] ), .B(n10247), .X(n2379) );
  nor_x1_sg U11613 ( .A(\reg_in[2][3][13] ), .B(n10454), .X(n2375) );
  nor_x1_sg U11614 ( .A(\reg_in[2][3][15] ), .B(n10553), .X(n2367) );
  nor_x1_sg U11615 ( .A(\reg_in[2][3][16] ), .B(n10554), .X(n2363) );
  nor_x1_sg U11616 ( .A(\reg_in[2][3][18] ), .B(n10034), .X(n2355) );
  nor_x1_sg U11617 ( .A(\reg_in[2][3][19] ), .B(n10122), .X(n2351) );
  nor_x1_sg U11618 ( .A(\reg_in[3][3][1] ), .B(n10279), .X(n2343) );
  nor_x1_sg U11619 ( .A(\reg_in[3][3][2] ), .B(n10291), .X(n2339) );
  nor_x1_sg U11620 ( .A(\reg_in[3][3][4] ), .B(n10277), .X(n2331) );
  nor_x1_sg U11621 ( .A(\reg_in[3][3][5] ), .B(n10127), .X(n2327) );
  nor_x1_sg U11622 ( .A(\reg_in[3][3][7] ), .B(n10227), .X(n2319) );
  nor_x1_sg U11623 ( .A(\reg_in[3][3][8] ), .B(n10500), .X(n2315) );
  nor_x1_sg U11624 ( .A(\reg_in[3][3][10] ), .B(n10444), .X(n2307) );
  nor_x1_sg U11625 ( .A(\reg_in[3][3][11] ), .B(n10280), .X(n2303) );
  nor_x1_sg U11626 ( .A(\reg_in[3][3][13] ), .B(n10034), .X(n2295) );
  nor_x1_sg U11627 ( .A(\reg_in[3][3][14] ), .B(n10548), .X(n2291) );
  nor_x1_sg U11628 ( .A(\reg_in[3][3][16] ), .B(n10546), .X(n2283) );
  nor_x1_sg U11629 ( .A(\reg_in[3][3][17] ), .B(n10246), .X(n2279) );
  nor_x1_sg U11630 ( .A(\reg_in[3][3][19] ), .B(n10496), .X(n2271) );
  nand_x1_sg U11631 ( .A(n10061), .B(\reg_in[0][0][0] ), .X(n8381) );
  nand_x1_sg U11632 ( .A(n10561), .B(\reg_in[0][0][1] ), .X(n8062) );
  nand_x1_sg U11633 ( .A(n10560), .B(\reg_in[0][0][2] ), .X(n8063) );
  nand_x1_sg U11634 ( .A(n10565), .B(\reg_in[0][0][3] ), .X(n8064) );
  nand_x1_sg U11635 ( .A(n10419), .B(\reg_in[0][0][4] ), .X(n8065) );
  nand_x1_sg U11636 ( .A(n10429), .B(\reg_in[0][0][5] ), .X(n8066) );
  nand_x1_sg U11637 ( .A(n10237), .B(\reg_in[0][0][6] ), .X(n8067) );
  nand_x1_sg U11638 ( .A(n10560), .B(\reg_in[0][0][7] ), .X(n8068) );
  nand_x1_sg U11639 ( .A(n10310), .B(\reg_in[0][0][8] ), .X(n8069) );
  nand_x1_sg U11640 ( .A(n10486), .B(\reg_in[0][0][9] ), .X(n8070) );
  nand_x1_sg U11641 ( .A(n10485), .B(\reg_in[0][0][10] ), .X(n8071) );
  nand_x1_sg U11642 ( .A(n10415), .B(\reg_in[0][0][11] ), .X(n8072) );
  nand_x1_sg U11643 ( .A(n10487), .B(\reg_in[0][0][12] ), .X(n8073) );
  nand_x1_sg U11644 ( .A(n10065), .B(\reg_in[0][0][13] ), .X(n8074) );
  nand_x1_sg U11645 ( .A(n10232), .B(\reg_in[0][0][14] ), .X(n8075) );
  nand_x1_sg U11646 ( .A(n10231), .B(\reg_in[0][0][15] ), .X(n8076) );
  nand_x1_sg U11647 ( .A(n10207), .B(\reg_in[0][0][16] ), .X(n8077) );
  nand_x1_sg U11648 ( .A(n10413), .B(\reg_in[0][0][17] ), .X(n8078) );
  nand_x1_sg U11649 ( .A(n10020), .B(\reg_in[0][0][18] ), .X(n8079) );
  nand_x1_sg U11650 ( .A(n10563), .B(\reg_in[0][0][19] ), .X(n8080) );
  nand_x1_sg U11651 ( .A(n10489), .B(\reg_in[1][0][0] ), .X(n8081) );
  nand_x1_sg U11652 ( .A(n10415), .B(\reg_in[1][0][1] ), .X(n8082) );
  nand_x1_sg U11653 ( .A(n10031), .B(\reg_in[1][0][2] ), .X(n8083) );
  nand_x1_sg U11654 ( .A(n10431), .B(\reg_in[1][0][3] ), .X(n8084) );
  nand_x1_sg U11655 ( .A(n10250), .B(\reg_in[1][0][4] ), .X(n8085) );
  nand_x1_sg U11656 ( .A(n10426), .B(\reg_in[1][0][5] ), .X(n8086) );
  nand_x1_sg U11657 ( .A(n10416), .B(\reg_in[1][0][6] ), .X(n8087) );
  nand_x1_sg U11658 ( .A(n10061), .B(\reg_in[1][0][7] ), .X(n8088) );
  nand_x1_sg U11659 ( .A(n10032), .B(\reg_in[1][0][8] ), .X(n8089) );
  nand_x1_sg U11660 ( .A(n10431), .B(\reg_in[1][0][9] ), .X(n8090) );
  nand_x1_sg U11661 ( .A(n10567), .B(\reg_in[1][0][10] ), .X(n8091) );
  nand_x1_sg U11662 ( .A(n10196), .B(\reg_in[1][0][11] ), .X(n8092) );
  nand_x1_sg U11663 ( .A(n10250), .B(\reg_in[1][0][12] ), .X(n8093) );
  nand_x1_sg U11664 ( .A(n10113), .B(\reg_in[1][0][13] ), .X(n8094) );
  nand_x1_sg U11665 ( .A(n10420), .B(\reg_in[1][0][14] ), .X(n8095) );
  nand_x1_sg U11666 ( .A(n10562), .B(\reg_in[1][0][15] ), .X(n8096) );
  nand_x1_sg U11667 ( .A(n10561), .B(\reg_in[1][0][16] ), .X(n8097) );
  nand_x1_sg U11668 ( .A(n10545), .B(\reg_in[1][0][17] ), .X(n8098) );
  nand_x1_sg U11669 ( .A(n10234), .B(\reg_in[1][0][18] ), .X(n8099) );
  nand_x1_sg U11670 ( .A(n10566), .B(\reg_in[1][0][19] ), .X(n8100) );
  nand_x1_sg U11671 ( .A(n10563), .B(\reg_in[2][0][0] ), .X(n8101) );
  nand_x1_sg U11672 ( .A(n10193), .B(\reg_in[2][0][1] ), .X(n8102) );
  nand_x1_sg U11673 ( .A(n10238), .B(\reg_in[2][0][2] ), .X(n8103) );
  nand_x1_sg U11674 ( .A(n10488), .B(\reg_in[2][0][3] ), .X(n8104) );
  nand_x1_sg U11675 ( .A(n10490), .B(\reg_in[2][0][4] ), .X(n8105) );
  nand_x1_sg U11676 ( .A(n10428), .B(\reg_in[2][0][5] ), .X(n8106) );
  nand_x1_sg U11677 ( .A(n10029), .B(\reg_in[2][0][6] ), .X(n8107) );
  nand_x1_sg U11678 ( .A(n10487), .B(\reg_in[2][0][7] ), .X(n8108) );
  nand_x1_sg U11679 ( .A(n10425), .B(\reg_in[2][0][8] ), .X(n8109) );
  nand_x1_sg U11680 ( .A(n10430), .B(\reg_in[2][0][9] ), .X(n8110) );
  nand_x1_sg U11681 ( .A(n10679), .B(\reg_in[2][0][10] ), .X(n8111) );
  nand_x1_sg U11682 ( .A(n10146), .B(\reg_in[2][0][11] ), .X(n8112) );
  nand_x1_sg U11683 ( .A(n10452), .B(\reg_in[2][0][12] ), .X(n8113) );
  nand_x1_sg U11684 ( .A(n10543), .B(\reg_in[2][0][13] ), .X(n8114) );
  nand_x1_sg U11685 ( .A(n10207), .B(\reg_in[2][0][14] ), .X(n8115) );
  nand_x1_sg U11686 ( .A(n10426), .B(\reg_in[2][0][15] ), .X(n8116) );
  nand_x1_sg U11687 ( .A(n10020), .B(\reg_in[2][0][16] ), .X(n8117) );
  nand_x1_sg U11688 ( .A(n10109), .B(\reg_in[2][0][17] ), .X(n8118) );
  nand_x1_sg U11689 ( .A(n10250), .B(\reg_in[2][0][18] ), .X(n8119) );
  nand_x1_sg U11690 ( .A(n10309), .B(\reg_in[2][0][19] ), .X(n8120) );
  nand_x1_sg U11691 ( .A(n10419), .B(\reg_in[3][0][0] ), .X(n8121) );
  nand_x1_sg U11692 ( .A(n10565), .B(\reg_in[3][0][1] ), .X(n8122) );
  nand_x1_sg U11693 ( .A(n10310), .B(\reg_in[3][0][2] ), .X(n8123) );
  nand_x1_sg U11694 ( .A(n10486), .B(\reg_in[3][0][3] ), .X(n8124) );
  nand_x1_sg U11695 ( .A(n10289), .B(\reg_in[3][0][4] ), .X(n8125) );
  nand_x1_sg U11696 ( .A(n10433), .B(\reg_in[3][0][5] ), .X(n8126) );
  nand_x1_sg U11697 ( .A(n10240), .B(\reg_in[3][0][6] ), .X(n8127) );
  nand_x1_sg U11698 ( .A(n10233), .B(\reg_in[3][0][7] ), .X(n8128) );
  nand_x1_sg U11699 ( .A(n10229), .B(\reg_in[3][0][8] ), .X(n8129) );
  nand_x1_sg U11700 ( .A(n10230), .B(\reg_in[3][0][9] ), .X(n8130) );
  nand_x1_sg U11701 ( .A(n10544), .B(\reg_in[3][0][10] ), .X(n8131) );
  nand_x1_sg U11702 ( .A(n10413), .B(\reg_in[3][0][11] ), .X(n8132) );
  nand_x1_sg U11703 ( .A(n10679), .B(\reg_in[3][0][12] ), .X(n8133) );
  nand_x1_sg U11704 ( .A(n10417), .B(\reg_in[3][0][13] ), .X(n8134) );
  nand_x1_sg U11705 ( .A(n10232), .B(\reg_in[3][0][14] ), .X(n8135) );
  nand_x1_sg U11706 ( .A(n10207), .B(\reg_in[3][0][15] ), .X(n8136) );
  nand_x1_sg U11707 ( .A(n10087), .B(\reg_in[3][0][16] ), .X(n8137) );
  nand_x1_sg U11708 ( .A(n10250), .B(\reg_in[3][0][17] ), .X(n8138) );
  nand_x1_sg U11709 ( .A(n10207), .B(\reg_in[3][0][18] ), .X(n8139) );
  nand_x1_sg U11710 ( .A(n10249), .B(\reg_in[3][0][19] ), .X(n8140) );
  nand_x1_sg U11711 ( .A(n10434), .B(\reg_in[0][1][0] ), .X(n8141) );
  nand_x1_sg U11712 ( .A(n10412), .B(\reg_in[0][1][1] ), .X(n8142) );
  nand_x1_sg U11713 ( .A(n10061), .B(\reg_in[0][1][2] ), .X(n8143) );
  nand_x1_sg U11714 ( .A(n10025), .B(\reg_in[0][1][3] ), .X(n8144) );
  nand_x1_sg U11715 ( .A(n10490), .B(\reg_in[0][1][4] ), .X(n8145) );
  nand_x1_sg U11716 ( .A(n10428), .B(\reg_in[0][1][5] ), .X(n8146) );
  nand_x1_sg U11717 ( .A(n10562), .B(\reg_in[0][1][6] ), .X(n8147) );
  nand_x1_sg U11718 ( .A(n10209), .B(\reg_in[0][1][7] ), .X(n8148) );
  nand_x1_sg U11719 ( .A(n10069), .B(\reg_in[0][1][8] ), .X(n8149) );
  nand_x1_sg U11720 ( .A(n10489), .B(\reg_in[0][1][9] ), .X(n8150) );
  nand_x1_sg U11721 ( .A(n10239), .B(\reg_in[0][1][10] ), .X(n8151) );
  nand_x1_sg U11722 ( .A(n10545), .B(\reg_in[0][1][11] ), .X(n8152) );
  nand_x1_sg U11723 ( .A(n10240), .B(\reg_in[0][1][12] ), .X(n8153) );
  nand_x1_sg U11724 ( .A(n10289), .B(\reg_in[0][1][13] ), .X(n8154) );
  nand_x1_sg U11725 ( .A(n10231), .B(\reg_in[0][1][14] ), .X(n8155) );
  nand_x1_sg U11726 ( .A(n10485), .B(\reg_in[0][1][15] ), .X(n8156) );
  nand_x1_sg U11727 ( .A(n10236), .B(\reg_in[0][1][16] ), .X(n8157) );
  nand_x1_sg U11728 ( .A(n10109), .B(\reg_in[0][1][17] ), .X(n8158) );
  nand_x1_sg U11729 ( .A(n10237), .B(\reg_in[0][1][18] ), .X(n8159) );
  nand_x1_sg U11730 ( .A(n10235), .B(\reg_in[0][1][19] ), .X(n8160) );
  nand_x1_sg U11731 ( .A(n10543), .B(\reg_in[1][1][0] ), .X(n8161) );
  nand_x1_sg U11732 ( .A(n10237), .B(\reg_in[1][1][1] ), .X(n8162) );
  nand_x1_sg U11733 ( .A(n10147), .B(\reg_in[1][1][2] ), .X(n8163) );
  nand_x1_sg U11734 ( .A(n10109), .B(\reg_in[1][1][3] ), .X(n8164) );
  nand_x1_sg U11735 ( .A(n10029), .B(\reg_in[1][1][4] ), .X(n8165) );
  nand_x1_sg U11736 ( .A(n10238), .B(\reg_in[1][1][5] ), .X(n8166) );
  nand_x1_sg U11737 ( .A(n10681), .B(\reg_in[1][1][6] ), .X(n8167) );
  nand_x1_sg U11738 ( .A(n10069), .B(\reg_in[1][1][7] ), .X(n8168) );
  nand_x1_sg U11739 ( .A(n10545), .B(\reg_in[1][1][8] ), .X(n8169) );
  nand_x1_sg U11740 ( .A(n10422), .B(\reg_in[1][1][9] ), .X(n8170) );
  nand_x1_sg U11741 ( .A(n10111), .B(\reg_in[1][1][10] ), .X(n8171) );
  nand_x1_sg U11742 ( .A(n10237), .B(\reg_in[1][1][11] ), .X(n8172) );
  nand_x1_sg U11743 ( .A(n10567), .B(\reg_in[1][1][12] ), .X(n8173) );
  nand_x1_sg U11744 ( .A(n10035), .B(\reg_in[1][1][13] ), .X(n8174) );
  nand_x1_sg U11745 ( .A(n10208), .B(\reg_in[1][1][14] ), .X(n8175) );
  nand_x1_sg U11746 ( .A(n10452), .B(\reg_in[1][1][15] ), .X(n8176) );
  nand_x1_sg U11747 ( .A(n10544), .B(\reg_in[1][1][16] ), .X(n8177) );
  nand_x1_sg U11748 ( .A(n10067), .B(\reg_in[1][1][17] ), .X(n8178) );
  nand_x1_sg U11749 ( .A(n10208), .B(\reg_in[1][1][18] ), .X(n8179) );
  nand_x1_sg U11750 ( .A(n10431), .B(\reg_in[1][1][19] ), .X(n8180) );
  nand_x1_sg U11751 ( .A(n10566), .B(\reg_in[2][1][0] ), .X(n8181) );
  nand_x1_sg U11752 ( .A(n10197), .B(\reg_in[2][1][1] ), .X(n8182) );
  nand_x1_sg U11753 ( .A(n10111), .B(\reg_in[2][1][2] ), .X(n8183) );
  nand_x1_sg U11754 ( .A(n10028), .B(\reg_in[2][1][3] ), .X(n8184) );
  nand_x1_sg U11755 ( .A(n10069), .B(\reg_in[2][1][4] ), .X(n8185) );
  nand_x1_sg U11756 ( .A(n10433), .B(\reg_in[2][1][5] ), .X(n8186) );
  nand_x1_sg U11757 ( .A(n10425), .B(\reg_in[2][1][6] ), .X(n8187) );
  nand_x1_sg U11758 ( .A(n10024), .B(\reg_in[2][1][7] ), .X(n8188) );
  nand_x1_sg U11759 ( .A(n10235), .B(\reg_in[2][1][8] ), .X(n8189) );
  nand_x1_sg U11760 ( .A(n10146), .B(\reg_in[2][1][9] ), .X(n8190) );
  nand_x1_sg U11761 ( .A(n10239), .B(\reg_in[2][1][10] ), .X(n8191) );
  nand_x1_sg U11762 ( .A(n10421), .B(\reg_in[2][1][11] ), .X(n8192) );
  nand_x1_sg U11763 ( .A(n10429), .B(\reg_in[2][1][12] ), .X(n8193) );
  nand_x1_sg U11764 ( .A(n10487), .B(\reg_in[2][1][13] ), .X(n8194) );
  nand_x1_sg U11765 ( .A(n10111), .B(\reg_in[2][1][14] ), .X(n8195) );
  nand_x1_sg U11766 ( .A(n10234), .B(\reg_in[2][1][15] ), .X(n8196) );
  nand_x1_sg U11767 ( .A(n10025), .B(\reg_in[2][1][16] ), .X(n8197) );
  nand_x1_sg U11768 ( .A(n10028), .B(\reg_in[2][1][17] ), .X(n8198) );
  nand_x1_sg U11769 ( .A(n10231), .B(\reg_in[2][1][18] ), .X(n8199) );
  nand_x1_sg U11770 ( .A(n10543), .B(\reg_in[2][1][19] ), .X(n8200) );
  nand_x1_sg U11771 ( .A(n10562), .B(\reg_in[3][1][0] ), .X(n8201) );
  nand_x1_sg U11772 ( .A(n10428), .B(\reg_in[3][1][1] ), .X(n8202) );
  nand_x1_sg U11773 ( .A(n10026), .B(\reg_in[3][1][2] ), .X(n8203) );
  nand_x1_sg U11774 ( .A(n10028), .B(\reg_in[3][1][3] ), .X(n8204) );
  nand_x1_sg U11775 ( .A(n8712), .B(\reg_in[3][1][4] ), .X(n8205) );
  nand_x1_sg U11776 ( .A(n10559), .B(\reg_in[3][1][5] ), .X(n8206) );
  nand_x1_sg U11777 ( .A(n10426), .B(\reg_in[3][1][6] ), .X(n8207) );
  nand_x1_sg U11778 ( .A(n10675), .B(\reg_in[3][1][7] ), .X(n8208) );
  nand_x1_sg U11779 ( .A(n10433), .B(\reg_in[3][1][8] ), .X(n8209) );
  nand_x1_sg U11780 ( .A(n10420), .B(\reg_in[3][1][9] ), .X(n8210) );
  nand_x1_sg U11781 ( .A(n10416), .B(\reg_in[3][1][10] ), .X(n8211) );
  nand_x1_sg U11782 ( .A(n10430), .B(\reg_in[3][1][11] ), .X(n8212) );
  nand_x1_sg U11783 ( .A(n10310), .B(\reg_in[3][1][12] ), .X(n8213) );
  nand_x1_sg U11784 ( .A(n10032), .B(\reg_in[3][1][13] ), .X(n8214) );
  nand_x1_sg U11785 ( .A(n10026), .B(\reg_in[3][1][14] ), .X(n8215) );
  nand_x1_sg U11786 ( .A(n10545), .B(\reg_in[3][1][15] ), .X(n8216) );
  nand_x1_sg U11787 ( .A(n10430), .B(\reg_in[3][1][16] ), .X(n8217) );
  nand_x1_sg U11788 ( .A(n10026), .B(\reg_in[3][1][17] ), .X(n8218) );
  nand_x1_sg U11789 ( .A(n10230), .B(\reg_in[3][1][18] ), .X(n8219) );
  nand_x1_sg U11790 ( .A(n10558), .B(\reg_in[3][1][19] ), .X(n8220) );
  nand_x1_sg U11791 ( .A(n10565), .B(\reg_in[0][2][0] ), .X(n8221) );
  nand_x1_sg U11792 ( .A(n10233), .B(\reg_in[0][2][1] ), .X(n8222) );
  nand_x1_sg U11793 ( .A(n10031), .B(\reg_in[0][2][2] ), .X(n8223) );
  nand_x1_sg U11794 ( .A(n10109), .B(\reg_in[0][2][3] ), .X(n8224) );
  nand_x1_sg U11795 ( .A(n10559), .B(\reg_in[0][2][4] ), .X(n8225) );
  nand_x1_sg U11796 ( .A(n10412), .B(\reg_in[0][2][5] ), .X(n8226) );
  nand_x1_sg U11797 ( .A(n10025), .B(\reg_in[0][2][6] ), .X(n8227) );
  nand_x1_sg U11798 ( .A(n10234), .B(\reg_in[0][2][7] ), .X(n8228) );
  nand_x1_sg U11799 ( .A(n10412), .B(\reg_in[0][2][8] ), .X(n8229) );
  nand_x1_sg U11800 ( .A(n10113), .B(\reg_in[0][2][9] ), .X(n8230) );
  nand_x1_sg U11801 ( .A(n10429), .B(\reg_in[0][2][10] ), .X(n8231) );
  nand_x1_sg U11802 ( .A(n10032), .B(\reg_in[0][2][11] ), .X(n8232) );
  nand_x1_sg U11803 ( .A(n10067), .B(\reg_in[0][2][12] ), .X(n8233) );
  nand_x1_sg U11804 ( .A(n10249), .B(\reg_in[0][2][13] ), .X(n8234) );
  nand_x1_sg U11805 ( .A(n10230), .B(\reg_in[0][2][14] ), .X(n8235) );
  nand_x1_sg U11806 ( .A(n10233), .B(\reg_in[0][2][15] ), .X(n8236) );
  nand_x1_sg U11807 ( .A(n10417), .B(\reg_in[0][2][16] ), .X(n8237) );
  nand_x1_sg U11808 ( .A(n10420), .B(\reg_in[0][2][17] ), .X(n8238) );
  nand_x1_sg U11809 ( .A(n10490), .B(\reg_in[0][2][18] ), .X(n8239) );
  nand_x1_sg U11810 ( .A(n10309), .B(\reg_in[0][2][19] ), .X(n8240) );
  nand_x1_sg U11811 ( .A(n10419), .B(\reg_in[1][2][0] ), .X(n8241) );
  nand_x1_sg U11812 ( .A(n10435), .B(\reg_in[1][2][1] ), .X(n8242) );
  nand_x1_sg U11813 ( .A(n10026), .B(\reg_in[1][2][2] ), .X(n8243) );
  nand_x1_sg U11814 ( .A(n10229), .B(\reg_in[1][2][3] ), .X(n8244) );
  nand_x1_sg U11815 ( .A(n10567), .B(\reg_in[1][2][4] ), .X(n8245) );
  nand_x1_sg U11816 ( .A(n10485), .B(\reg_in[1][2][5] ), .X(n8246) );
  nand_x1_sg U11817 ( .A(n10681), .B(\reg_in[1][2][6] ), .X(n8247) );
  nand_x1_sg U11818 ( .A(n10069), .B(\reg_in[1][2][7] ), .X(n8248) );
  nand_x1_sg U11819 ( .A(n10235), .B(\reg_in[1][2][8] ), .X(n8249) );
  nand_x1_sg U11820 ( .A(n10543), .B(\reg_in[1][2][9] ), .X(n8250) );
  nand_x1_sg U11821 ( .A(n10067), .B(\reg_in[1][2][10] ), .X(n8251) );
  nand_x1_sg U11822 ( .A(n10425), .B(\reg_in[1][2][11] ), .X(n8252) );
  nand_x1_sg U11823 ( .A(n10229), .B(\reg_in[1][2][12] ), .X(n8253) );
  nand_x1_sg U11824 ( .A(n10209), .B(\reg_in[1][2][13] ), .X(n8254) );
  nand_x1_sg U11825 ( .A(n10558), .B(\reg_in[1][2][14] ), .X(n8255) );
  nand_x1_sg U11826 ( .A(n10563), .B(\reg_in[1][2][15] ), .X(n8256) );
  nand_x1_sg U11827 ( .A(n10067), .B(\reg_in[1][2][16] ), .X(n8257) );
  nand_x1_sg U11828 ( .A(n10310), .B(\reg_in[1][2][17] ), .X(n8258) );
  nand_x1_sg U11829 ( .A(n10486), .B(\reg_in[1][2][18] ), .X(n8259) );
  nand_x1_sg U11830 ( .A(n10498), .B(\reg_in[1][2][19] ), .X(n8260) );
  nand_x1_sg U11831 ( .A(n10567), .B(\reg_in[2][2][0] ), .X(n8261) );
  nand_x1_sg U11832 ( .A(n10249), .B(\reg_in[2][2][1] ), .X(n8262) );
  nand_x1_sg U11833 ( .A(n10675), .B(\reg_in[2][2][2] ), .X(n8263) );
  nand_x1_sg U11834 ( .A(n10231), .B(\reg_in[2][2][3] ), .X(n8264) );
  nand_x1_sg U11835 ( .A(n10424), .B(\reg_in[2][2][4] ), .X(n8265) );
  nand_x1_sg U11836 ( .A(n10485), .B(\reg_in[2][2][5] ), .X(n8266) );
  nand_x1_sg U11837 ( .A(n8712), .B(\reg_in[2][2][6] ), .X(n8267) );
  nand_x1_sg U11838 ( .A(n10020), .B(\reg_in[2][2][7] ), .X(n8268) );
  nand_x1_sg U11839 ( .A(n10433), .B(\reg_in[2][2][8] ), .X(n8269) );
  nand_x1_sg U11840 ( .A(n10412), .B(\reg_in[2][2][9] ), .X(n8270) );
  nand_x1_sg U11841 ( .A(n10562), .B(\reg_in[2][2][10] ), .X(n8271) );
  nand_x1_sg U11842 ( .A(n10428), .B(\reg_in[2][2][11] ), .X(n8272) );
  nand_x1_sg U11843 ( .A(n10020), .B(\reg_in[2][2][12] ), .X(n8273) );
  nand_x1_sg U11844 ( .A(n10489), .B(\reg_in[2][2][13] ), .X(n8274) );
  nand_x1_sg U11845 ( .A(n10236), .B(\reg_in[2][2][14] ), .X(n8275) );
  nand_x1_sg U11846 ( .A(n10239), .B(\reg_in[2][2][15] ), .X(n8276) );
  nand_x1_sg U11847 ( .A(n10239), .B(\reg_in[2][2][16] ), .X(n8277) );
  nand_x1_sg U11848 ( .A(n10249), .B(\reg_in[2][2][17] ), .X(n8278) );
  nand_x1_sg U11849 ( .A(n10431), .B(\reg_in[2][2][18] ), .X(n8279) );
  nand_x1_sg U11850 ( .A(n10035), .B(\reg_in[2][2][19] ), .X(n8280) );
  nand_x1_sg U11851 ( .A(n10234), .B(\reg_in[3][2][0] ), .X(n8281) );
  nand_x1_sg U11852 ( .A(n10415), .B(\reg_in[3][2][1] ), .X(n8282) );
  nand_x1_sg U11853 ( .A(n10209), .B(\reg_in[3][2][2] ), .X(n8283) );
  nand_x1_sg U11854 ( .A(n10193), .B(\reg_in[3][2][3] ), .X(n8284) );
  nand_x1_sg U11855 ( .A(n10233), .B(\reg_in[3][2][4] ), .X(n8285) );
  nand_x1_sg U11856 ( .A(n10031), .B(\reg_in[3][2][5] ), .X(n8286) );
  nand_x1_sg U11857 ( .A(n10430), .B(\reg_in[3][2][6] ), .X(n8287) );
  nand_x1_sg U11858 ( .A(n10028), .B(\reg_in[3][2][7] ), .X(n8288) );
  nand_x1_sg U11859 ( .A(n10193), .B(\reg_in[3][2][8] ), .X(n8289) );
  nand_x1_sg U11860 ( .A(n10420), .B(\reg_in[3][2][9] ), .X(n8290) );
  nand_x1_sg U11861 ( .A(n10558), .B(\reg_in[3][2][10] ), .X(n8291) );
  nand_x1_sg U11862 ( .A(n10493), .B(\reg_in[3][2][11] ), .X(n8292) );
  nand_x1_sg U11863 ( .A(n10209), .B(\reg_in[3][2][12] ), .X(n8293) );
  nand_x1_sg U11864 ( .A(n10044), .B(\reg_in[3][2][13] ), .X(n8294) );
  nand_x1_sg U11865 ( .A(n10025), .B(\reg_in[3][2][14] ), .X(n8295) );
  nand_x1_sg U11866 ( .A(n10232), .B(\reg_in[3][2][15] ), .X(n8296) );
  nand_x1_sg U11867 ( .A(n10421), .B(\reg_in[3][2][16] ), .X(n8297) );
  nand_x1_sg U11868 ( .A(n10488), .B(\reg_in[3][2][17] ), .X(n8298) );
  nand_x1_sg U11869 ( .A(n10065), .B(\reg_in[3][2][18] ), .X(n8299) );
  nand_x1_sg U11870 ( .A(n10197), .B(\reg_in[3][2][19] ), .X(n8300) );
  nand_x1_sg U11871 ( .A(n10196), .B(\reg_in[0][3][0] ), .X(n8301) );
  nand_x1_sg U11872 ( .A(n10415), .B(\reg_in[0][3][1] ), .X(n8302) );
  nand_x1_sg U11873 ( .A(n10017), .B(\reg_in[0][3][2] ), .X(n8303) );
  nand_x1_sg U11874 ( .A(n10488), .B(\reg_in[0][3][3] ), .X(n8304) );
  nand_x1_sg U11875 ( .A(n10424), .B(\reg_in[0][3][4] ), .X(n8305) );
  nand_x1_sg U11876 ( .A(n10544), .B(\reg_in[0][3][5] ), .X(n8306) );
  nand_x1_sg U11877 ( .A(n10024), .B(\reg_in[0][3][6] ), .X(n8307) );
  nand_x1_sg U11878 ( .A(n10681), .B(\reg_in[0][3][7] ), .X(n8308) );
  nand_x1_sg U11879 ( .A(n10490), .B(\reg_in[0][3][8] ), .X(n8309) );
  nand_x1_sg U11880 ( .A(n10432), .B(\reg_in[0][3][9] ), .X(n8310) );
  nand_x1_sg U11881 ( .A(n10236), .B(\reg_in[0][3][10] ), .X(n8311) );
  nand_x1_sg U11882 ( .A(n10236), .B(\reg_in[0][3][11] ), .X(n8312) );
  nand_x1_sg U11883 ( .A(n10432), .B(\reg_in[0][3][12] ), .X(n8313) );
  nand_x1_sg U11884 ( .A(n10421), .B(\reg_in[0][3][13] ), .X(n8314) );
  nand_x1_sg U11885 ( .A(n10424), .B(\reg_in[0][3][14] ), .X(n8315) );
  nand_x1_sg U11886 ( .A(n10679), .B(\reg_in[0][3][15] ), .X(n8316) );
  nand_x1_sg U11887 ( .A(n10238), .B(\reg_in[0][3][16] ), .X(n8317) );
  nand_x1_sg U11888 ( .A(n10196), .B(\reg_in[0][3][17] ), .X(n8318) );
  nand_x1_sg U11889 ( .A(n10240), .B(\reg_in[0][3][18] ), .X(n8319) );
  nand_x1_sg U11890 ( .A(n10559), .B(\reg_in[0][3][19] ), .X(n8320) );
  nand_x1_sg U11891 ( .A(n10417), .B(\reg_in[1][3][0] ), .X(n8321) );
  nand_x1_sg U11892 ( .A(n10486), .B(\reg_in[1][3][1] ), .X(n8322) );
  nand_x1_sg U11893 ( .A(n10435), .B(\reg_in[1][3][2] ), .X(n8323) );
  nand_x1_sg U11894 ( .A(n10413), .B(\reg_in[1][3][3] ), .X(n8324) );
  nand_x1_sg U11895 ( .A(n10435), .B(\reg_in[1][3][4] ), .X(n8325) );
  nand_x1_sg U11896 ( .A(n10029), .B(\reg_in[1][3][5] ), .X(n8326) );
  nand_x1_sg U11897 ( .A(n10196), .B(\reg_in[1][3][6] ), .X(n8327) );
  nand_x1_sg U11898 ( .A(n10229), .B(\reg_in[1][3][7] ), .X(n8328) );
  nand_x1_sg U11899 ( .A(n10289), .B(\reg_in[1][3][8] ), .X(n8329) );
  nand_x1_sg U11900 ( .A(n10432), .B(\reg_in[1][3][9] ), .X(n8330) );
  nand_x1_sg U11901 ( .A(n10424), .B(\reg_in[1][3][10] ), .X(n8331) );
  nand_x1_sg U11902 ( .A(n10422), .B(\reg_in[1][3][11] ), .X(n8332) );
  nand_x1_sg U11903 ( .A(n10558), .B(\reg_in[1][3][12] ), .X(n8333) );
  nand_x1_sg U11904 ( .A(n10417), .B(\reg_in[1][3][13] ), .X(n8334) );
  nand_x1_sg U11905 ( .A(n10232), .B(\reg_in[1][3][14] ), .X(n8335) );
  nand_x1_sg U11906 ( .A(n10208), .B(\reg_in[1][3][15] ), .X(n8336) );
  nand_x1_sg U11907 ( .A(n10421), .B(\reg_in[1][3][16] ), .X(n8337) );
  nand_x1_sg U11908 ( .A(n10032), .B(\reg_in[1][3][17] ), .X(n8338) );
  nand_x1_sg U11909 ( .A(n10238), .B(\reg_in[1][3][18] ), .X(n8339) );
  nand_x1_sg U11910 ( .A(n10208), .B(\reg_in[1][3][19] ), .X(n8340) );
  nand_x1_sg U11911 ( .A(n10146), .B(\reg_in[2][3][0] ), .X(n8341) );
  nand_x1_sg U11912 ( .A(n10240), .B(\reg_in[2][3][1] ), .X(n8342) );
  nand_x1_sg U11913 ( .A(n10419), .B(\reg_in[2][3][2] ), .X(n8343) );
  nand_x1_sg U11914 ( .A(n10493), .B(\reg_in[2][3][3] ), .X(n8344) );
  nand_x1_sg U11915 ( .A(n10031), .B(\reg_in[2][3][4] ), .X(n8345) );
  nand_x1_sg U11916 ( .A(n10434), .B(\reg_in[2][3][5] ), .X(n8346) );
  nand_x1_sg U11917 ( .A(n10432), .B(\reg_in[2][3][6] ), .X(n8347) );
  nand_x1_sg U11918 ( .A(n10147), .B(\reg_in[2][3][7] ), .X(n8348) );
  nand_x1_sg U11919 ( .A(n10422), .B(\reg_in[2][3][8] ), .X(n8349) );
  nand_x1_sg U11920 ( .A(n10435), .B(\reg_in[2][3][9] ), .X(n8350) );
  nand_x1_sg U11921 ( .A(n10111), .B(\reg_in[2][3][10] ), .X(n8351) );
  nand_x1_sg U11922 ( .A(n10113), .B(\reg_in[2][3][11] ), .X(n8352) );
  nand_x1_sg U11923 ( .A(n10489), .B(\reg_in[2][3][12] ), .X(n8353) );
  nand_x1_sg U11924 ( .A(n10487), .B(\reg_in[2][3][13] ), .X(n8354) );
  nand_x1_sg U11925 ( .A(n10061), .B(\reg_in[2][3][14] ), .X(n8355) );
  nand_x1_sg U11926 ( .A(n10024), .B(\reg_in[2][3][15] ), .X(n8356) );
  nand_x1_sg U11927 ( .A(n10563), .B(\reg_in[2][3][16] ), .X(n8357) );
  nand_x1_sg U11928 ( .A(n10560), .B(\reg_in[2][3][17] ), .X(n8358) );
  nand_x1_sg U11929 ( .A(n10087), .B(\reg_in[2][3][18] ), .X(n8359) );
  nand_x1_sg U11930 ( .A(n10029), .B(\reg_in[2][3][19] ), .X(n8360) );
  nand_x1_sg U11931 ( .A(n10416), .B(\reg_in[3][3][0] ), .X(n8361) );
  nand_x1_sg U11932 ( .A(n10425), .B(\reg_in[3][3][1] ), .X(n8362) );
  nand_x1_sg U11933 ( .A(n10498), .B(\reg_in[3][3][2] ), .X(n8363) );
  nand_x1_sg U11934 ( .A(n10147), .B(\reg_in[3][3][3] ), .X(n8364) );
  nand_x1_sg U11935 ( .A(n10544), .B(\reg_in[3][3][4] ), .X(n8365) );
  nand_x1_sg U11936 ( .A(n10561), .B(\reg_in[3][3][5] ), .X(n8366) );
  nand_x1_sg U11937 ( .A(n10044), .B(\reg_in[3][3][6] ), .X(n8367) );
  nand_x1_sg U11938 ( .A(n10309), .B(\reg_in[3][3][7] ), .X(n8368) );
  nand_x1_sg U11939 ( .A(n10566), .B(\reg_in[3][3][8] ), .X(n8369) );
  nand_x1_sg U11940 ( .A(n10113), .B(\reg_in[3][3][9] ), .X(n8370) );
  nand_x1_sg U11941 ( .A(n10230), .B(\reg_in[3][3][10] ), .X(n8371) );
  nand_x1_sg U11942 ( .A(n10679), .B(\reg_in[3][3][11] ), .X(n8372) );
  nand_x1_sg U11943 ( .A(n10197), .B(\reg_in[3][3][12] ), .X(n8373) );
  nand_x1_sg U11944 ( .A(n10434), .B(\reg_in[3][3][13] ), .X(n8374) );
  nand_x1_sg U11945 ( .A(n10147), .B(\reg_in[3][3][14] ), .X(n8375) );
  nand_x1_sg U11946 ( .A(n10197), .B(\reg_in[3][3][15] ), .X(n8376) );
  nand_x1_sg U11947 ( .A(n10566), .B(\reg_in[3][3][16] ), .X(n8377) );
  nand_x1_sg U11948 ( .A(n10024), .B(\reg_in[3][3][17] ), .X(n8378) );
  nand_x1_sg U11949 ( .A(n10235), .B(\reg_in[3][3][18] ), .X(n8379) );
  nand_x1_sg U11950 ( .A(n10146), .B(\reg_in[3][3][19] ), .X(n8380) );
endmodule

