
module post_sparsity ( clk, reset, .i_im({\i_im[15][19] , \i_im[15][18] , 
        \i_im[15][17] , \i_im[15][16] , \i_im[15][15] , \i_im[15][14] , 
        \i_im[15][13] , \i_im[15][12] , \i_im[15][11] , \i_im[15][10] , 
        \i_im[15][9] , \i_im[15][8] , \i_im[15][7] , \i_im[15][6] , 
        \i_im[15][5] , \i_im[15][4] , \i_im[15][3] , \i_im[15][2] , 
        \i_im[15][1] , \i_im[15][0] , \i_im[14][19] , \i_im[14][18] , 
        \i_im[14][17] , \i_im[14][16] , \i_im[14][15] , \i_im[14][14] , 
        \i_im[14][13] , \i_im[14][12] , \i_im[14][11] , \i_im[14][10] , 
        \i_im[14][9] , \i_im[14][8] , \i_im[14][7] , \i_im[14][6] , 
        \i_im[14][5] , \i_im[14][4] , \i_im[14][3] , \i_im[14][2] , 
        \i_im[14][1] , \i_im[14][0] , \i_im[13][19] , \i_im[13][18] , 
        \i_im[13][17] , \i_im[13][16] , \i_im[13][15] , \i_im[13][14] , 
        \i_im[13][13] , \i_im[13][12] , \i_im[13][11] , \i_im[13][10] , 
        \i_im[13][9] , \i_im[13][8] , \i_im[13][7] , \i_im[13][6] , 
        \i_im[13][5] , \i_im[13][4] , \i_im[13][3] , \i_im[13][2] , 
        \i_im[13][1] , \i_im[13][0] , \i_im[12][19] , \i_im[12][18] , 
        \i_im[12][17] , \i_im[12][16] , \i_im[12][15] , \i_im[12][14] , 
        \i_im[12][13] , \i_im[12][12] , \i_im[12][11] , \i_im[12][10] , 
        \i_im[12][9] , \i_im[12][8] , \i_im[12][7] , \i_im[12][6] , 
        \i_im[12][5] , \i_im[12][4] , \i_im[12][3] , \i_im[12][2] , 
        \i_im[12][1] , \i_im[12][0] , \i_im[11][19] , \i_im[11][18] , 
        \i_im[11][17] , \i_im[11][16] , \i_im[11][15] , \i_im[11][14] , 
        \i_im[11][13] , \i_im[11][12] , \i_im[11][11] , \i_im[11][10] , 
        \i_im[11][9] , \i_im[11][8] , \i_im[11][7] , \i_im[11][6] , 
        \i_im[11][5] , \i_im[11][4] , \i_im[11][3] , \i_im[11][2] , 
        \i_im[11][1] , \i_im[11][0] , \i_im[10][19] , \i_im[10][18] , 
        \i_im[10][17] , \i_im[10][16] , \i_im[10][15] , \i_im[10][14] , 
        \i_im[10][13] , \i_im[10][12] , \i_im[10][11] , \i_im[10][10] , 
        \i_im[10][9] , \i_im[10][8] , \i_im[10][7] , \i_im[10][6] , 
        \i_im[10][5] , \i_im[10][4] , \i_im[10][3] , \i_im[10][2] , 
        \i_im[10][1] , \i_im[10][0] , \i_im[9][19] , \i_im[9][18] , 
        \i_im[9][17] , \i_im[9][16] , \i_im[9][15] , \i_im[9][14] , 
        \i_im[9][13] , \i_im[9][12] , \i_im[9][11] , \i_im[9][10] , 
        \i_im[9][9] , \i_im[9][8] , \i_im[9][7] , \i_im[9][6] , \i_im[9][5] , 
        \i_im[9][4] , \i_im[9][3] , \i_im[9][2] , \i_im[9][1] , \i_im[9][0] , 
        \i_im[8][19] , \i_im[8][18] , \i_im[8][17] , \i_im[8][16] , 
        \i_im[8][15] , \i_im[8][14] , \i_im[8][13] , \i_im[8][12] , 
        \i_im[8][11] , \i_im[8][10] , \i_im[8][9] , \i_im[8][8] , \i_im[8][7] , 
        \i_im[8][6] , \i_im[8][5] , \i_im[8][4] , \i_im[8][3] , \i_im[8][2] , 
        \i_im[8][1] , \i_im[8][0] , \i_im[7][19] , \i_im[7][18] , 
        \i_im[7][17] , \i_im[7][16] , \i_im[7][15] , \i_im[7][14] , 
        \i_im[7][13] , \i_im[7][12] , \i_im[7][11] , \i_im[7][10] , 
        \i_im[7][9] , \i_im[7][8] , \i_im[7][7] , \i_im[7][6] , \i_im[7][5] , 
        \i_im[7][4] , \i_im[7][3] , \i_im[7][2] , \i_im[7][1] , \i_im[7][0] , 
        \i_im[6][19] , \i_im[6][18] , \i_im[6][17] , \i_im[6][16] , 
        \i_im[6][15] , \i_im[6][14] , \i_im[6][13] , \i_im[6][12] , 
        \i_im[6][11] , \i_im[6][10] , \i_im[6][9] , \i_im[6][8] , \i_im[6][7] , 
        \i_im[6][6] , \i_im[6][5] , \i_im[6][4] , \i_im[6][3] , \i_im[6][2] , 
        \i_im[6][1] , \i_im[6][0] , \i_im[5][19] , \i_im[5][18] , 
        \i_im[5][17] , \i_im[5][16] , \i_im[5][15] , \i_im[5][14] , 
        \i_im[5][13] , \i_im[5][12] , \i_im[5][11] , \i_im[5][10] , 
        \i_im[5][9] , \i_im[5][8] , \i_im[5][7] , \i_im[5][6] , \i_im[5][5] , 
        \i_im[5][4] , \i_im[5][3] , \i_im[5][2] , \i_im[5][1] , \i_im[5][0] , 
        \i_im[4][19] , \i_im[4][18] , \i_im[4][17] , \i_im[4][16] , 
        \i_im[4][15] , \i_im[4][14] , \i_im[4][13] , \i_im[4][12] , 
        \i_im[4][11] , \i_im[4][10] , \i_im[4][9] , \i_im[4][8] , \i_im[4][7] , 
        \i_im[4][6] , \i_im[4][5] , \i_im[4][4] , \i_im[4][3] , \i_im[4][2] , 
        \i_im[4][1] , \i_im[4][0] , \i_im[3][19] , \i_im[3][18] , 
        \i_im[3][17] , \i_im[3][16] , \i_im[3][15] , \i_im[3][14] , 
        \i_im[3][13] , \i_im[3][12] , \i_im[3][11] , \i_im[3][10] , 
        \i_im[3][9] , \i_im[3][8] , \i_im[3][7] , \i_im[3][6] , \i_im[3][5] , 
        \i_im[3][4] , \i_im[3][3] , \i_im[3][2] , \i_im[3][1] , \i_im[3][0] , 
        \i_im[2][19] , \i_im[2][18] , \i_im[2][17] , \i_im[2][16] , 
        \i_im[2][15] , \i_im[2][14] , \i_im[2][13] , \i_im[2][12] , 
        \i_im[2][11] , \i_im[2][10] , \i_im[2][9] , \i_im[2][8] , \i_im[2][7] , 
        \i_im[2][6] , \i_im[2][5] , \i_im[2][4] , \i_im[2][3] , \i_im[2][2] , 
        \i_im[2][1] , \i_im[2][0] , \i_im[1][19] , \i_im[1][18] , 
        \i_im[1][17] , \i_im[1][16] , \i_im[1][15] , \i_im[1][14] , 
        \i_im[1][13] , \i_im[1][12] , \i_im[1][11] , \i_im[1][10] , 
        \i_im[1][9] , \i_im[1][8] , \i_im[1][7] , \i_im[1][6] , \i_im[1][5] , 
        \i_im[1][4] , \i_im[1][3] , \i_im[1][2] , \i_im[1][1] , \i_im[1][0] , 
        \i_im[0][19] , \i_im[0][18] , \i_im[0][17] , \i_im[0][16] , 
        \i_im[0][15] , \i_im[0][14] , \i_im[0][13] , \i_im[0][12] , 
        \i_im[0][11] , \i_im[0][10] , \i_im[0][9] , \i_im[0][8] , \i_im[0][7] , 
        \i_im[0][6] , \i_im[0][5] , \i_im[0][4] , \i_im[0][3] , \i_im[0][2] , 
        \i_im[0][1] , \i_im[0][0] }), i_mask, input_ready, output_taken, 
    .o_im({\o_im[15][19] , \o_im[15][18] , \o_im[15][17] , \o_im[15][16] , 
        \o_im[15][15] , \o_im[15][14] , \o_im[15][13] , \o_im[15][12] , 
        \o_im[15][11] , \o_im[15][10] , \o_im[15][9] , \o_im[15][8] , 
        \o_im[15][7] , \o_im[15][6] , \o_im[15][5] , \o_im[15][4] , 
        \o_im[15][3] , \o_im[15][2] , \o_im[15][1] , \o_im[15][0] , 
        \o_im[14][19] , \o_im[14][18] , \o_im[14][17] , \o_im[14][16] , 
        \o_im[14][15] , \o_im[14][14] , \o_im[14][13] , \o_im[14][12] , 
        \o_im[14][11] , \o_im[14][10] , \o_im[14][9] , \o_im[14][8] , 
        \o_im[14][7] , \o_im[14][6] , \o_im[14][5] , \o_im[14][4] , 
        \o_im[14][3] , \o_im[14][2] , \o_im[14][1] , \o_im[14][0] , 
        \o_im[13][19] , \o_im[13][18] , \o_im[13][17] , \o_im[13][16] , 
        \o_im[13][15] , \o_im[13][14] , \o_im[13][13] , \o_im[13][12] , 
        \o_im[13][11] , \o_im[13][10] , \o_im[13][9] , \o_im[13][8] , 
        \o_im[13][7] , \o_im[13][6] , \o_im[13][5] , \o_im[13][4] , 
        \o_im[13][3] , \o_im[13][2] , \o_im[13][1] , \o_im[13][0] , 
        \o_im[12][19] , \o_im[12][18] , \o_im[12][17] , \o_im[12][16] , 
        \o_im[12][15] , \o_im[12][14] , \o_im[12][13] , \o_im[12][12] , 
        \o_im[12][11] , \o_im[12][10] , \o_im[12][9] , \o_im[12][8] , 
        \o_im[12][7] , \o_im[12][6] , \o_im[12][5] , \o_im[12][4] , 
        \o_im[12][3] , \o_im[12][2] , \o_im[12][1] , \o_im[12][0] , 
        \o_im[11][19] , \o_im[11][18] , \o_im[11][17] , \o_im[11][16] , 
        \o_im[11][15] , \o_im[11][14] , \o_im[11][13] , \o_im[11][12] , 
        \o_im[11][11] , \o_im[11][10] , \o_im[11][9] , \o_im[11][8] , 
        \o_im[11][7] , \o_im[11][6] , \o_im[11][5] , \o_im[11][4] , 
        \o_im[11][3] , \o_im[11][2] , \o_im[11][1] , \o_im[11][0] , 
        \o_im[10][19] , \o_im[10][18] , \o_im[10][17] , \o_im[10][16] , 
        \o_im[10][15] , \o_im[10][14] , \o_im[10][13] , \o_im[10][12] , 
        \o_im[10][11] , \o_im[10][10] , \o_im[10][9] , \o_im[10][8] , 
        \o_im[10][7] , \o_im[10][6] , \o_im[10][5] , \o_im[10][4] , 
        \o_im[10][3] , \o_im[10][2] , \o_im[10][1] , \o_im[10][0] , 
        \o_im[9][19] , \o_im[9][18] , \o_im[9][17] , \o_im[9][16] , 
        \o_im[9][15] , \o_im[9][14] , \o_im[9][13] , \o_im[9][12] , 
        \o_im[9][11] , \o_im[9][10] , \o_im[9][9] , \o_im[9][8] , \o_im[9][7] , 
        \o_im[9][6] , \o_im[9][5] , \o_im[9][4] , \o_im[9][3] , \o_im[9][2] , 
        \o_im[9][1] , \o_im[9][0] , \o_im[8][19] , \o_im[8][18] , 
        \o_im[8][17] , \o_im[8][16] , \o_im[8][15] , \o_im[8][14] , 
        \o_im[8][13] , \o_im[8][12] , \o_im[8][11] , \o_im[8][10] , 
        \o_im[8][9] , \o_im[8][8] , \o_im[8][7] , \o_im[8][6] , \o_im[8][5] , 
        \o_im[8][4] , \o_im[8][3] , \o_im[8][2] , \o_im[8][1] , \o_im[8][0] , 
        \o_im[7][19] , \o_im[7][18] , \o_im[7][17] , \o_im[7][16] , 
        \o_im[7][15] , \o_im[7][14] , \o_im[7][13] , \o_im[7][12] , 
        \o_im[7][11] , \o_im[7][10] , \o_im[7][9] , \o_im[7][8] , \o_im[7][7] , 
        \o_im[7][6] , \o_im[7][5] , \o_im[7][4] , \o_im[7][3] , \o_im[7][2] , 
        \o_im[7][1] , \o_im[7][0] , \o_im[6][19] , \o_im[6][18] , 
        \o_im[6][17] , \o_im[6][16] , \o_im[6][15] , \o_im[6][14] , 
        \o_im[6][13] , \o_im[6][12] , \o_im[6][11] , \o_im[6][10] , 
        \o_im[6][9] , \o_im[6][8] , \o_im[6][7] , \o_im[6][6] , \o_im[6][5] , 
        \o_im[6][4] , \o_im[6][3] , \o_im[6][2] , \o_im[6][1] , \o_im[6][0] , 
        \o_im[5][19] , \o_im[5][18] , \o_im[5][17] , \o_im[5][16] , 
        \o_im[5][15] , \o_im[5][14] , \o_im[5][13] , \o_im[5][12] , 
        \o_im[5][11] , \o_im[5][10] , \o_im[5][9] , \o_im[5][8] , \o_im[5][7] , 
        \o_im[5][6] , \o_im[5][5] , \o_im[5][4] , \o_im[5][3] , \o_im[5][2] , 
        \o_im[5][1] , \o_im[5][0] , \o_im[4][19] , \o_im[4][18] , 
        \o_im[4][17] , \o_im[4][16] , \o_im[4][15] , \o_im[4][14] , 
        \o_im[4][13] , \o_im[4][12] , \o_im[4][11] , \o_im[4][10] , 
        \o_im[4][9] , \o_im[4][8] , \o_im[4][7] , \o_im[4][6] , \o_im[4][5] , 
        \o_im[4][4] , \o_im[4][3] , \o_im[4][2] , \o_im[4][1] , \o_im[4][0] , 
        \o_im[3][19] , \o_im[3][18] , \o_im[3][17] , \o_im[3][16] , 
        \o_im[3][15] , \o_im[3][14] , \o_im[3][13] , \o_im[3][12] , 
        \o_im[3][11] , \o_im[3][10] , \o_im[3][9] , \o_im[3][8] , \o_im[3][7] , 
        \o_im[3][6] , \o_im[3][5] , \o_im[3][4] , \o_im[3][3] , \o_im[3][2] , 
        \o_im[3][1] , \o_im[3][0] , \o_im[2][19] , \o_im[2][18] , 
        \o_im[2][17] , \o_im[2][16] , \o_im[2][15] , \o_im[2][14] , 
        \o_im[2][13] , \o_im[2][12] , \o_im[2][11] , \o_im[2][10] , 
        \o_im[2][9] , \o_im[2][8] , \o_im[2][7] , \o_im[2][6] , \o_im[2][5] , 
        \o_im[2][4] , \o_im[2][3] , \o_im[2][2] , \o_im[2][1] , \o_im[2][0] , 
        \o_im[1][19] , \o_im[1][18] , \o_im[1][17] , \o_im[1][16] , 
        \o_im[1][15] , \o_im[1][14] , \o_im[1][13] , \o_im[1][12] , 
        \o_im[1][11] , \o_im[1][10] , \o_im[1][9] , \o_im[1][8] , \o_im[1][7] , 
        \o_im[1][6] , \o_im[1][5] , \o_im[1][4] , \o_im[1][3] , \o_im[1][2] , 
        \o_im[1][1] , \o_im[1][0] , \o_im[0][19] , \o_im[0][18] , 
        \o_im[0][17] , \o_im[0][16] , \o_im[0][15] , \o_im[0][14] , 
        \o_im[0][13] , \o_im[0][12] , \o_im[0][11] , \o_im[0][10] , 
        \o_im[0][9] , \o_im[0][8] , \o_im[0][7] , \o_im[0][6] , \o_im[0][5] , 
        \o_im[0][4] , \o_im[0][3] , \o_im[0][2] , \o_im[0][1] , \o_im[0][0] }), 
        o_mask, state );
  input [31:0] i_mask;
  output [31:0] o_mask;
  output [1:0] state;
  input clk, reset, \i_im[15][19] , \i_im[15][18] , \i_im[15][17] ,
         \i_im[15][16] , \i_im[15][15] , \i_im[15][14] , \i_im[15][13] ,
         \i_im[15][12] , \i_im[15][11] , \i_im[15][10] , \i_im[15][9] ,
         \i_im[15][8] , \i_im[15][7] , \i_im[15][6] , \i_im[15][5] ,
         \i_im[15][4] , \i_im[15][3] , \i_im[15][2] , \i_im[15][1] ,
         \i_im[15][0] , \i_im[14][19] , \i_im[14][18] , \i_im[14][17] ,
         \i_im[14][16] , \i_im[14][15] , \i_im[14][14] , \i_im[14][13] ,
         \i_im[14][12] , \i_im[14][11] , \i_im[14][10] , \i_im[14][9] ,
         \i_im[14][8] , \i_im[14][7] , \i_im[14][6] , \i_im[14][5] ,
         \i_im[14][4] , \i_im[14][3] , \i_im[14][2] , \i_im[14][1] ,
         \i_im[14][0] , \i_im[13][19] , \i_im[13][18] , \i_im[13][17] ,
         \i_im[13][16] , \i_im[13][15] , \i_im[13][14] , \i_im[13][13] ,
         \i_im[13][12] , \i_im[13][11] , \i_im[13][10] , \i_im[13][9] ,
         \i_im[13][8] , \i_im[13][7] , \i_im[13][6] , \i_im[13][5] ,
         \i_im[13][4] , \i_im[13][3] , \i_im[13][2] , \i_im[13][1] ,
         \i_im[13][0] , \i_im[12][19] , \i_im[12][18] , \i_im[12][17] ,
         \i_im[12][16] , \i_im[12][15] , \i_im[12][14] , \i_im[12][13] ,
         \i_im[12][12] , \i_im[12][11] , \i_im[12][10] , \i_im[12][9] ,
         \i_im[12][8] , \i_im[12][7] , \i_im[12][6] , \i_im[12][5] ,
         \i_im[12][4] , \i_im[12][3] , \i_im[12][2] , \i_im[12][1] ,
         \i_im[12][0] , \i_im[11][19] , \i_im[11][18] , \i_im[11][17] ,
         \i_im[11][16] , \i_im[11][15] , \i_im[11][14] , \i_im[11][13] ,
         \i_im[11][12] , \i_im[11][11] , \i_im[11][10] , \i_im[11][9] ,
         \i_im[11][8] , \i_im[11][7] , \i_im[11][6] , \i_im[11][5] ,
         \i_im[11][4] , \i_im[11][3] , \i_im[11][2] , \i_im[11][1] ,
         \i_im[11][0] , \i_im[10][19] , \i_im[10][18] , \i_im[10][17] ,
         \i_im[10][16] , \i_im[10][15] , \i_im[10][14] , \i_im[10][13] ,
         \i_im[10][12] , \i_im[10][11] , \i_im[10][10] , \i_im[10][9] ,
         \i_im[10][8] , \i_im[10][7] , \i_im[10][6] , \i_im[10][5] ,
         \i_im[10][4] , \i_im[10][3] , \i_im[10][2] , \i_im[10][1] ,
         \i_im[10][0] , \i_im[9][19] , \i_im[9][18] , \i_im[9][17] ,
         \i_im[9][16] , \i_im[9][15] , \i_im[9][14] , \i_im[9][13] ,
         \i_im[9][12] , \i_im[9][11] , \i_im[9][10] , \i_im[9][9] ,
         \i_im[9][8] , \i_im[9][7] , \i_im[9][6] , \i_im[9][5] , \i_im[9][4] ,
         \i_im[9][3] , \i_im[9][2] , \i_im[9][1] , \i_im[9][0] , \i_im[8][19] ,
         \i_im[8][18] , \i_im[8][17] , \i_im[8][16] , \i_im[8][15] ,
         \i_im[8][14] , \i_im[8][13] , \i_im[8][12] , \i_im[8][11] ,
         \i_im[8][10] , \i_im[8][9] , \i_im[8][8] , \i_im[8][7] , \i_im[8][6] ,
         \i_im[8][5] , \i_im[8][4] , \i_im[8][3] , \i_im[8][2] , \i_im[8][1] ,
         \i_im[8][0] , \i_im[7][19] , \i_im[7][18] , \i_im[7][17] ,
         \i_im[7][16] , \i_im[7][15] , \i_im[7][14] , \i_im[7][13] ,
         \i_im[7][12] , \i_im[7][11] , \i_im[7][10] , \i_im[7][9] ,
         \i_im[7][8] , \i_im[7][7] , \i_im[7][6] , \i_im[7][5] , \i_im[7][4] ,
         \i_im[7][3] , \i_im[7][2] , \i_im[7][1] , \i_im[7][0] , \i_im[6][19] ,
         \i_im[6][18] , \i_im[6][17] , \i_im[6][16] , \i_im[6][15] ,
         \i_im[6][14] , \i_im[6][13] , \i_im[6][12] , \i_im[6][11] ,
         \i_im[6][10] , \i_im[6][9] , \i_im[6][8] , \i_im[6][7] , \i_im[6][6] ,
         \i_im[6][5] , \i_im[6][4] , \i_im[6][3] , \i_im[6][2] , \i_im[6][1] ,
         \i_im[6][0] , \i_im[5][19] , \i_im[5][18] , \i_im[5][17] ,
         \i_im[5][16] , \i_im[5][15] , \i_im[5][14] , \i_im[5][13] ,
         \i_im[5][12] , \i_im[5][11] , \i_im[5][10] , \i_im[5][9] ,
         \i_im[5][8] , \i_im[5][7] , \i_im[5][6] , \i_im[5][5] , \i_im[5][4] ,
         \i_im[5][3] , \i_im[5][2] , \i_im[5][1] , \i_im[5][0] , \i_im[4][19] ,
         \i_im[4][18] , \i_im[4][17] , \i_im[4][16] , \i_im[4][15] ,
         \i_im[4][14] , \i_im[4][13] , \i_im[4][12] , \i_im[4][11] ,
         \i_im[4][10] , \i_im[4][9] , \i_im[4][8] , \i_im[4][7] , \i_im[4][6] ,
         \i_im[4][5] , \i_im[4][4] , \i_im[4][3] , \i_im[4][2] , \i_im[4][1] ,
         \i_im[4][0] , \i_im[3][19] , \i_im[3][18] , \i_im[3][17] ,
         \i_im[3][16] , \i_im[3][15] , \i_im[3][14] , \i_im[3][13] ,
         \i_im[3][12] , \i_im[3][11] , \i_im[3][10] , \i_im[3][9] ,
         \i_im[3][8] , \i_im[3][7] , \i_im[3][6] , \i_im[3][5] , \i_im[3][4] ,
         \i_im[3][3] , \i_im[3][2] , \i_im[3][1] , \i_im[3][0] , \i_im[2][19] ,
         \i_im[2][18] , \i_im[2][17] , \i_im[2][16] , \i_im[2][15] ,
         \i_im[2][14] , \i_im[2][13] , \i_im[2][12] , \i_im[2][11] ,
         \i_im[2][10] , \i_im[2][9] , \i_im[2][8] , \i_im[2][7] , \i_im[2][6] ,
         \i_im[2][5] , \i_im[2][4] , \i_im[2][3] , \i_im[2][2] , \i_im[2][1] ,
         \i_im[2][0] , \i_im[1][19] , \i_im[1][18] , \i_im[1][17] ,
         \i_im[1][16] , \i_im[1][15] , \i_im[1][14] , \i_im[1][13] ,
         \i_im[1][12] , \i_im[1][11] , \i_im[1][10] , \i_im[1][9] ,
         \i_im[1][8] , \i_im[1][7] , \i_im[1][6] , \i_im[1][5] , \i_im[1][4] ,
         \i_im[1][3] , \i_im[1][2] , \i_im[1][1] , \i_im[1][0] , \i_im[0][19] ,
         \i_im[0][18] , \i_im[0][17] , \i_im[0][16] , \i_im[0][15] ,
         \i_im[0][14] , \i_im[0][13] , \i_im[0][12] , \i_im[0][11] ,
         \i_im[0][10] , \i_im[0][9] , \i_im[0][8] , \i_im[0][7] , \i_im[0][6] ,
         \i_im[0][5] , \i_im[0][4] , \i_im[0][3] , \i_im[0][2] , \i_im[0][1] ,
         \i_im[0][0] , input_ready, output_taken;
  output \o_im[15][19] , \o_im[15][18] , \o_im[15][17] , \o_im[15][16] ,
         \o_im[15][15] , \o_im[15][14] , \o_im[15][13] , \o_im[15][12] ,
         \o_im[15][11] , \o_im[15][10] , \o_im[15][9] , \o_im[15][8] ,
         \o_im[15][7] , \o_im[15][6] , \o_im[15][5] , \o_im[15][4] ,
         \o_im[15][3] , \o_im[15][2] , \o_im[15][1] , \o_im[15][0] ,
         \o_im[14][19] , \o_im[14][18] , \o_im[14][17] , \o_im[14][16] ,
         \o_im[14][15] , \o_im[14][14] , \o_im[14][13] , \o_im[14][12] ,
         \o_im[14][11] , \o_im[14][10] , \o_im[14][9] , \o_im[14][8] ,
         \o_im[14][7] , \o_im[14][6] , \o_im[14][5] , \o_im[14][4] ,
         \o_im[14][3] , \o_im[14][2] , \o_im[14][1] , \o_im[14][0] ,
         \o_im[13][19] , \o_im[13][18] , \o_im[13][17] , \o_im[13][16] ,
         \o_im[13][15] , \o_im[13][14] , \o_im[13][13] , \o_im[13][12] ,
         \o_im[13][11] , \o_im[13][10] , \o_im[13][9] , \o_im[13][8] ,
         \o_im[13][7] , \o_im[13][6] , \o_im[13][5] , \o_im[13][4] ,
         \o_im[13][3] , \o_im[13][2] , \o_im[13][1] , \o_im[13][0] ,
         \o_im[12][19] , \o_im[12][18] , \o_im[12][17] , \o_im[12][16] ,
         \o_im[12][15] , \o_im[12][14] , \o_im[12][13] , \o_im[12][12] ,
         \o_im[12][11] , \o_im[12][10] , \o_im[12][9] , \o_im[12][8] ,
         \o_im[12][7] , \o_im[12][6] , \o_im[12][5] , \o_im[12][4] ,
         \o_im[12][3] , \o_im[12][2] , \o_im[12][1] , \o_im[12][0] ,
         \o_im[11][19] , \o_im[11][18] , \o_im[11][17] , \o_im[11][16] ,
         \o_im[11][15] , \o_im[11][14] , \o_im[11][13] , \o_im[11][12] ,
         \o_im[11][11] , \o_im[11][10] , \o_im[11][9] , \o_im[11][8] ,
         \o_im[11][7] , \o_im[11][6] , \o_im[11][5] , \o_im[11][4] ,
         \o_im[11][3] , \o_im[11][2] , \o_im[11][1] , \o_im[11][0] ,
         \o_im[10][19] , \o_im[10][18] , \o_im[10][17] , \o_im[10][16] ,
         \o_im[10][15] , \o_im[10][14] , \o_im[10][13] , \o_im[10][12] ,
         \o_im[10][11] , \o_im[10][10] , \o_im[10][9] , \o_im[10][8] ,
         \o_im[10][7] , \o_im[10][6] , \o_im[10][5] , \o_im[10][4] ,
         \o_im[10][3] , \o_im[10][2] , \o_im[10][1] , \o_im[10][0] ,
         \o_im[9][19] , \o_im[9][18] , \o_im[9][17] , \o_im[9][16] ,
         \o_im[9][15] , \o_im[9][14] , \o_im[9][13] , \o_im[9][12] ,
         \o_im[9][11] , \o_im[9][10] , \o_im[9][9] , \o_im[9][8] ,
         \o_im[9][7] , \o_im[9][6] , \o_im[9][5] , \o_im[9][4] , \o_im[9][3] ,
         \o_im[9][2] , \o_im[9][1] , \o_im[9][0] , \o_im[8][19] ,
         \o_im[8][18] , \o_im[8][17] , \o_im[8][16] , \o_im[8][15] ,
         \o_im[8][14] , \o_im[8][13] , \o_im[8][12] , \o_im[8][11] ,
         \o_im[8][10] , \o_im[8][9] , \o_im[8][8] , \o_im[8][7] , \o_im[8][6] ,
         \o_im[8][5] , \o_im[8][4] , \o_im[8][3] , \o_im[8][2] , \o_im[8][1] ,
         \o_im[8][0] , \o_im[7][19] , \o_im[7][18] , \o_im[7][17] ,
         \o_im[7][16] , \o_im[7][15] , \o_im[7][14] , \o_im[7][13] ,
         \o_im[7][12] , \o_im[7][11] , \o_im[7][10] , \o_im[7][9] ,
         \o_im[7][8] , \o_im[7][7] , \o_im[7][6] , \o_im[7][5] , \o_im[7][4] ,
         \o_im[7][3] , \o_im[7][2] , \o_im[7][1] , \o_im[7][0] , \o_im[6][19] ,
         \o_im[6][18] , \o_im[6][17] , \o_im[6][16] , \o_im[6][15] ,
         \o_im[6][14] , \o_im[6][13] , \o_im[6][12] , \o_im[6][11] ,
         \o_im[6][10] , \o_im[6][9] , \o_im[6][8] , \o_im[6][7] , \o_im[6][6] ,
         \o_im[6][5] , \o_im[6][4] , \o_im[6][3] , \o_im[6][2] , \o_im[6][1] ,
         \o_im[6][0] , \o_im[5][19] , \o_im[5][18] , \o_im[5][17] ,
         \o_im[5][16] , \o_im[5][15] , \o_im[5][14] , \o_im[5][13] ,
         \o_im[5][12] , \o_im[5][11] , \o_im[5][10] , \o_im[5][9] ,
         \o_im[5][8] , \o_im[5][7] , \o_im[5][6] , \o_im[5][5] , \o_im[5][4] ,
         \o_im[5][3] , \o_im[5][2] , \o_im[5][1] , \o_im[5][0] , \o_im[4][19] ,
         \o_im[4][18] , \o_im[4][17] , \o_im[4][16] , \o_im[4][15] ,
         \o_im[4][14] , \o_im[4][13] , \o_im[4][12] , \o_im[4][11] ,
         \o_im[4][10] , \o_im[4][9] , \o_im[4][8] , \o_im[4][7] , \o_im[4][6] ,
         \o_im[4][5] , \o_im[4][4] , \o_im[4][3] , \o_im[4][2] , \o_im[4][1] ,
         \o_im[4][0] , \o_im[3][19] , \o_im[3][18] , \o_im[3][17] ,
         \o_im[3][16] , \o_im[3][15] , \o_im[3][14] , \o_im[3][13] ,
         \o_im[3][12] , \o_im[3][11] , \o_im[3][10] , \o_im[3][9] ,
         \o_im[3][8] , \o_im[3][7] , \o_im[3][6] , \o_im[3][5] , \o_im[3][4] ,
         \o_im[3][3] , \o_im[3][2] , \o_im[3][1] , \o_im[3][0] , \o_im[2][19] ,
         \o_im[2][18] , \o_im[2][17] , \o_im[2][16] , \o_im[2][15] ,
         \o_im[2][14] , \o_im[2][13] , \o_im[2][12] , \o_im[2][11] ,
         \o_im[2][10] , \o_im[2][9] , \o_im[2][8] , \o_im[2][7] , \o_im[2][6] ,
         \o_im[2][5] , \o_im[2][4] , \o_im[2][3] , \o_im[2][2] , \o_im[2][1] ,
         \o_im[2][0] , \o_im[1][19] , \o_im[1][18] , \o_im[1][17] ,
         \o_im[1][16] , \o_im[1][15] , \o_im[1][14] , \o_im[1][13] ,
         \o_im[1][12] , \o_im[1][11] , \o_im[1][10] , \o_im[1][9] ,
         \o_im[1][8] , \o_im[1][7] , \o_im[1][6] , \o_im[1][5] , \o_im[1][4] ,
         \o_im[1][3] , \o_im[1][2] , \o_im[1][1] , \o_im[1][0] , \o_im[0][19] ,
         \o_im[0][18] , \o_im[0][17] , \o_im[0][16] , \o_im[0][15] ,
         \o_im[0][14] , \o_im[0][13] , \o_im[0][12] , \o_im[0][11] ,
         \o_im[0][10] , \o_im[0][9] , \o_im[0][8] , \o_im[0][7] , \o_im[0][6] ,
         \o_im[0][5] , \o_im[0][4] , \o_im[0][3] , \o_im[0][2] , \o_im[0][1] ,
         \o_im[0][0] ;
  wire   \mask_state[0] , \output_state[0] , n19, n20, \update_mask_0/n1835 ,
         \update_mask_0/n1442 , \update_mask_0/n1441 , \update_mask_0/n1440 ,
         \update_mask_0/n1439 , \update_mask_0/n1438 , \update_mask_0/n1437 ,
         \update_mask_0/n1436 , \update_mask_0/n1435 , \update_mask_0/n1434 ,
         \update_mask_0/n1433 , \update_mask_0/n1432 , \update_mask_0/n1431 ,
         \update_mask_0/n1430 , \update_mask_0/n1429 , \update_mask_0/n1428 ,
         \update_mask_0/n1427 , \update_mask_0/n1426 , \update_mask_0/n1425 ,
         \update_mask_0/n1424 , \update_mask_0/n1423 , \update_mask_0/n1422 ,
         \update_mask_0/n1421 , \update_mask_0/n1420 , \update_mask_0/n1419 ,
         \update_mask_0/n1418 , \update_mask_0/n1417 , \update_mask_0/n1416 ,
         \update_mask_0/n1415 , \update_mask_0/n1414 , \update_mask_0/n1413 ,
         \update_mask_0/n1412 , \update_mask_0/n1411 , \update_mask_0/n1410 ,
         \update_mask_0/n1409 , \update_mask_0/n1408 , \update_mask_0/n1407 ,
         \update_mask_0/n1406 , \update_mask_0/n1405 , \update_mask_0/n1404 ,
         \update_mask_0/n1403 , \update_mask_0/n1402 , \update_mask_0/n1401 ,
         \update_mask_0/n1400 , \update_mask_0/n1399 , \update_mask_0/n1398 ,
         \update_mask_0/n1397 , \update_mask_0/n1396 , \update_mask_0/n1395 ,
         \update_mask_0/n1394 , \update_mask_0/n1393 , \update_mask_0/n1392 ,
         \update_mask_0/n1391 , \update_mask_0/n1390 , \update_mask_0/n1389 ,
         \update_mask_0/n1388 , \update_mask_0/n1387 , \update_mask_0/n1386 ,
         \update_mask_0/n1385 , \update_mask_0/n1384 , \update_mask_0/n1383 ,
         \update_mask_0/n1382 , \update_mask_0/n1381 , \update_mask_0/n1380 ,
         \update_mask_0/n1379 , \update_mask_0/n1378 , \update_mask_0/n1377 ,
         \update_mask_0/n1376 , \update_mask_0/n1375 , \update_mask_0/n1374 ,
         \update_mask_0/n1373 , \update_mask_0/n1372 , \update_mask_0/n1371 ,
         \update_mask_0/n1370 , \update_mask_0/n1369 , \update_mask_0/n1368 ,
         \update_mask_0/n1367 , \update_mask_0/n1366 , \update_mask_0/n1365 ,
         \update_mask_0/n1364 , \update_mask_0/n1363 , \update_mask_0/n1362 ,
         \update_mask_0/n1361 , \update_mask_0/n1360 , \update_mask_0/n1359 ,
         \update_mask_0/n1358 , \update_mask_0/n1357 , \update_mask_0/n1356 ,
         \update_mask_0/n1355 , \update_mask_0/n1354 , \update_mask_0/n1353 ,
         \update_mask_0/n1352 , \update_mask_0/n1351 , \update_mask_0/n1350 ,
         \update_mask_0/n1349 , \update_mask_0/n1348 , \update_mask_0/n1347 ,
         \update_mask_0/n1346 , \update_mask_0/n1345 , \update_mask_0/n1344 ,
         \update_mask_0/n1343 , \update_mask_0/n1342 , \update_mask_0/n1341 ,
         \update_mask_0/n1340 , \update_mask_0/n1339 , \update_mask_0/n1338 ,
         \update_mask_0/n1337 , \update_mask_0/n1336 , \update_mask_0/n1335 ,
         \update_mask_0/n1334 , \update_mask_0/n1333 , \update_mask_0/n1332 ,
         \update_mask_0/n1331 , \update_mask_0/n1330 , \update_mask_0/n1329 ,
         \update_mask_0/n1328 , \update_mask_0/n1327 , \update_mask_0/n1326 ,
         \update_mask_0/n1325 , \update_mask_0/n1324 , \update_mask_0/n1323 ,
         \update_mask_0/n1322 , \update_mask_0/n1321 , \update_mask_0/n1320 ,
         \update_mask_0/n1319 , \update_mask_0/n1318 , \update_mask_0/n1317 ,
         \update_mask_0/n1316 , \update_mask_0/n1315 , \update_mask_0/n1314 ,
         \update_mask_0/n1313 , \update_mask_0/n1312 , \update_mask_0/n1311 ,
         \update_mask_0/n1310 , \update_mask_0/n1309 , \update_mask_0/n1308 ,
         \update_mask_0/n1307 , \update_mask_0/n1306 , \update_mask_0/n1305 ,
         \update_mask_0/n1304 , \update_mask_0/n1303 , \update_mask_0/n1302 ,
         \update_mask_0/n1301 , \update_mask_0/n1300 , \update_mask_0/n1299 ,
         \update_mask_0/n1298 , \update_mask_0/n1297 , \update_mask_0/n1296 ,
         \update_mask_0/n1295 , \update_mask_0/n1294 , \update_mask_0/n1293 ,
         \update_mask_0/n1292 , \update_mask_0/n1291 , \update_mask_0/n1290 ,
         \update_mask_0/n1289 , \update_mask_0/n1288 , \update_mask_0/n1287 ,
         \update_mask_0/n1286 , \update_mask_0/n1285 , \update_mask_0/n1284 ,
         \update_mask_0/n1283 , \update_mask_0/n1282 , \update_mask_0/n1281 ,
         \update_mask_0/n1280 , \update_mask_0/n1279 , \update_mask_0/n1278 ,
         \update_mask_0/n1277 , \update_mask_0/n1276 , \update_mask_0/n1275 ,
         \update_mask_0/n1274 , \update_mask_0/n1273 , \update_mask_0/n1272 ,
         \update_mask_0/n1271 , \update_mask_0/n1270 , \update_mask_0/n1269 ,
         \update_mask_0/n1268 , \update_mask_0/n1267 , \update_mask_0/n1266 ,
         \update_mask_0/n1265 , \update_mask_0/n1264 , \update_mask_0/n1263 ,
         \update_mask_0/n1262 , \update_mask_0/n1261 , \update_mask_0/n1260 ,
         \update_mask_0/n1259 , \update_mask_0/n1258 , \update_mask_0/n1257 ,
         \update_mask_0/n1256 , \update_mask_0/n1255 , \update_mask_0/n1254 ,
         \update_mask_0/n1253 , \update_mask_0/n1252 , \update_mask_0/n1251 ,
         \update_mask_0/n1250 , \update_mask_0/n1249 , \update_mask_0/n1248 ,
         \update_mask_0/n1247 , \update_mask_0/n1246 , \update_mask_0/n1245 ,
         \update_mask_0/n1244 , \update_mask_0/n1243 , \update_mask_0/n1242 ,
         \update_mask_0/n1241 , \update_mask_0/n1240 , \update_mask_0/n1239 ,
         \update_mask_0/n1238 , \update_mask_0/n1237 , \update_mask_0/n1236 ,
         \update_mask_0/n1235 , \update_mask_0/n1234 , \update_mask_0/n1233 ,
         \update_mask_0/n1232 , \update_mask_0/n1231 , \update_mask_0/n1230 ,
         \update_mask_0/n1229 , \update_mask_0/n1228 , \update_mask_0/n1227 ,
         \update_mask_0/n1226 , \update_mask_0/n1225 , \update_mask_0/n1224 ,
         \update_mask_0/n1223 , \update_mask_0/n1222 , \update_mask_0/n1221 ,
         \update_mask_0/n1220 , \update_mask_0/n1219 , \update_mask_0/n1218 ,
         \update_mask_0/n1217 , \update_mask_0/n1216 , \update_mask_0/n1215 ,
         \update_mask_0/n1214 , \update_mask_0/n1213 , \update_mask_0/n1212 ,
         \update_mask_0/n1211 , \update_mask_0/n1210 , \update_mask_0/n1209 ,
         \update_mask_0/n1208 , \update_mask_0/n1207 , \update_mask_0/n1206 ,
         \update_mask_0/n1205 , \update_mask_0/n1204 , \update_mask_0/n1203 ,
         \update_mask_0/n1202 , \update_mask_0/n1201 , \update_mask_0/n1200 ,
         \update_mask_0/n1199 , \update_mask_0/n1198 , \update_mask_0/n1197 ,
         \update_mask_0/n1196 , \update_mask_0/n1195 , \update_mask_0/n1194 ,
         \update_mask_0/n1193 , \update_mask_0/n1192 , \update_mask_0/n1191 ,
         \update_mask_0/n1190 , \update_mask_0/n1189 , \update_mask_0/n1188 ,
         \update_mask_0/n1187 , \update_mask_0/n1186 , \update_mask_0/n1185 ,
         \update_mask_0/n1184 , \update_mask_0/n1183 , \update_mask_0/n1182 ,
         \update_mask_0/n1181 , \update_mask_0/n1180 , \update_mask_0/n1179 ,
         \update_mask_0/n1178 , \update_mask_0/n1177 , \update_mask_0/n1176 ,
         \update_mask_0/n1175 , \update_mask_0/n1174 , \update_mask_0/n1173 ,
         \update_mask_0/n1172 , \update_mask_0/n1171 , \update_mask_0/n1170 ,
         \update_mask_0/n1169 , \update_mask_0/n1168 , \update_mask_0/n1167 ,
         \update_mask_0/n1166 , \update_mask_0/n1165 , \update_mask_0/n1164 ,
         \update_mask_0/n1163 , \update_mask_0/n1162 , \update_mask_0/n1161 ,
         \update_mask_0/n1160 , \update_mask_0/n1159 , \update_mask_0/n1158 ,
         \update_mask_0/n1157 , \update_mask_0/n1156 , \update_mask_0/n1155 ,
         \update_mask_0/n1154 , \update_mask_0/n1153 , \update_mask_0/n1152 ,
         \update_mask_0/n1151 , \update_mask_0/n1150 , \update_mask_0/n1149 ,
         \update_mask_0/n1148 , \update_mask_0/n1147 , \update_mask_0/n1146 ,
         \update_mask_0/n1145 , \update_mask_0/n1144 , \update_mask_0/n1143 ,
         \update_mask_0/n1142 , \update_mask_0/n1141 , \update_mask_0/n1140 ,
         \update_mask_0/n1139 , \update_mask_0/n1138 , \update_mask_0/n1137 ,
         \update_mask_0/n1136 , \update_mask_0/n1135 , \update_mask_0/n1134 ,
         \update_mask_0/n1133 , \update_mask_0/n1132 , \update_mask_0/n1131 ,
         \update_mask_0/n1130 , \update_mask_0/n1129 , \update_mask_0/n1128 ,
         \update_mask_0/n1127 , \update_mask_0/n1126 , \update_mask_0/n1125 ,
         \update_mask_0/n1124 , \update_mask_0/n1123 , \update_mask_0/n1122 ,
         \update_mask_0/n1121 , \update_mask_0/n1120 , \update_mask_0/n1119 ,
         \update_mask_0/n1118 , \update_mask_0/n1117 , \update_mask_0/n1116 ,
         \update_mask_0/n1115 , \update_mask_0/n1114 , \update_mask_0/n1113 ,
         \update_mask_0/n1112 , \update_mask_0/n1111 , \update_mask_0/n1110 ,
         \update_mask_0/n1109 , \update_mask_0/n1108 , \update_mask_0/n1107 ,
         \update_mask_0/n1106 , \update_mask_0/n1105 , \update_mask_0/n1104 ,
         \update_mask_0/n1103 , \update_mask_0/n1102 , \update_mask_0/n1101 ,
         \update_mask_0/n1100 , \update_mask_0/n1099 , \update_mask_0/n1098 ,
         \update_mask_0/n1097 , \update_mask_0/n1096 , \update_mask_0/n1095 ,
         \update_mask_0/n1094 , \update_mask_0/n1093 , \update_mask_0/n1092 ,
         \update_mask_0/n1091 , \update_mask_0/n1090 , \update_mask_0/n1089 ,
         \update_mask_0/n1088 , \update_mask_0/n1087 , \update_mask_0/n1086 ,
         \update_mask_0/n1085 , \update_mask_0/n1084 , \update_mask_0/n1083 ,
         \update_mask_0/n1082 , \update_mask_0/n1081 ,
         \update_mask_0/reg_out[0][0] , \update_mask_0/reg_out[0][1] ,
         \update_mask_0/reg_out[0][2] , \update_mask_0/reg_out[0][3] ,
         \update_mask_0/reg_out[0][4] , \update_mask_0/reg_out[0][5] ,
         \update_mask_0/reg_out[0][6] , \update_mask_0/reg_out[0][7] ,
         \update_mask_0/reg_out[0][8] , \update_mask_0/reg_out[0][9] ,
         \update_mask_0/reg_out[0][10] , \update_mask_0/reg_out[0][11] ,
         \update_mask_0/reg_out[0][12] , \update_mask_0/reg_out[0][13] ,
         \update_mask_0/reg_out[0][14] , \update_mask_0/reg_out[0][15] ,
         \update_mask_0/reg_out[0][16] , \update_mask_0/reg_out[0][17] ,
         \update_mask_0/reg_out[0][18] , \update_mask_0/reg_out[0][19] ,
         \update_mask_0/reg_out[1][0] , \update_mask_0/reg_out[1][1] ,
         \update_mask_0/reg_out[1][2] , \update_mask_0/reg_out[1][3] ,
         \update_mask_0/reg_out[1][4] , \update_mask_0/reg_out[1][5] ,
         \update_mask_0/reg_out[1][6] , \update_mask_0/reg_out[1][7] ,
         \update_mask_0/reg_out[1][8] , \update_mask_0/reg_out[1][9] ,
         \update_mask_0/reg_out[1][10] , \update_mask_0/reg_out[1][11] ,
         \update_mask_0/reg_out[1][12] , \update_mask_0/reg_out[1][13] ,
         \update_mask_0/reg_out[1][14] , \update_mask_0/reg_out[1][15] ,
         \update_mask_0/reg_out[1][16] , \update_mask_0/reg_out[1][17] ,
         \update_mask_0/reg_out[1][18] , \update_mask_0/reg_out[1][19] ,
         \update_mask_0/reg_out[2][0] , \update_mask_0/reg_out[2][1] ,
         \update_mask_0/reg_out[2][2] , \update_mask_0/reg_out[2][3] ,
         \update_mask_0/reg_out[2][4] , \update_mask_0/reg_out[2][5] ,
         \update_mask_0/reg_out[2][6] , \update_mask_0/reg_out[2][7] ,
         \update_mask_0/reg_out[2][8] , \update_mask_0/reg_out[2][9] ,
         \update_mask_0/reg_out[2][10] , \update_mask_0/reg_out[2][11] ,
         \update_mask_0/reg_out[2][12] , \update_mask_0/reg_out[2][13] ,
         \update_mask_0/reg_out[2][14] , \update_mask_0/reg_out[2][15] ,
         \update_mask_0/reg_out[2][16] , \update_mask_0/reg_out[2][17] ,
         \update_mask_0/reg_out[2][18] , \update_mask_0/reg_out[2][19] ,
         \update_mask_0/reg_out[3][0] , \update_mask_0/reg_out[3][1] ,
         \update_mask_0/reg_out[3][2] , \update_mask_0/reg_out[3][3] ,
         \update_mask_0/reg_out[3][4] , \update_mask_0/reg_out[3][5] ,
         \update_mask_0/reg_out[3][6] , \update_mask_0/reg_out[3][7] ,
         \update_mask_0/reg_out[3][8] , \update_mask_0/reg_out[3][9] ,
         \update_mask_0/reg_out[3][10] , \update_mask_0/reg_out[3][11] ,
         \update_mask_0/reg_out[3][12] , \update_mask_0/reg_out[3][13] ,
         \update_mask_0/reg_out[3][14] , \update_mask_0/reg_out[3][15] ,
         \update_mask_0/reg_out[3][16] , \update_mask_0/reg_out[3][17] ,
         \update_mask_0/reg_out[3][18] , \update_mask_0/reg_out[3][19] ,
         \update_mask_0/reg_out[4][0] , \update_mask_0/reg_out[4][1] ,
         \update_mask_0/reg_out[4][2] , \update_mask_0/reg_out[4][3] ,
         \update_mask_0/reg_out[4][4] , \update_mask_0/reg_out[4][5] ,
         \update_mask_0/reg_out[4][6] , \update_mask_0/reg_out[4][7] ,
         \update_mask_0/reg_out[4][8] , \update_mask_0/reg_out[4][9] ,
         \update_mask_0/reg_out[4][10] , \update_mask_0/reg_out[4][11] ,
         \update_mask_0/reg_out[4][12] , \update_mask_0/reg_out[4][13] ,
         \update_mask_0/reg_out[4][14] , \update_mask_0/reg_out[4][15] ,
         \update_mask_0/reg_out[4][16] , \update_mask_0/reg_out[4][17] ,
         \update_mask_0/reg_out[4][18] , \update_mask_0/reg_out[4][19] ,
         \update_mask_0/reg_out[5][0] , \update_mask_0/reg_out[5][1] ,
         \update_mask_0/reg_out[5][2] , \update_mask_0/reg_out[5][3] ,
         \update_mask_0/reg_out[5][4] , \update_mask_0/reg_out[5][5] ,
         \update_mask_0/reg_out[5][6] , \update_mask_0/reg_out[5][7] ,
         \update_mask_0/reg_out[5][8] , \update_mask_0/reg_out[5][9] ,
         \update_mask_0/reg_out[5][10] , \update_mask_0/reg_out[5][11] ,
         \update_mask_0/reg_out[5][12] , \update_mask_0/reg_out[5][13] ,
         \update_mask_0/reg_out[5][14] , \update_mask_0/reg_out[5][15] ,
         \update_mask_0/reg_out[5][16] , \update_mask_0/reg_out[5][17] ,
         \update_mask_0/reg_out[5][18] , \update_mask_0/reg_out[5][19] ,
         \update_mask_0/reg_out[6][0] , \update_mask_0/reg_out[6][1] ,
         \update_mask_0/reg_out[6][2] , \update_mask_0/reg_out[6][3] ,
         \update_mask_0/reg_out[6][4] , \update_mask_0/reg_out[6][5] ,
         \update_mask_0/reg_out[6][6] , \update_mask_0/reg_out[6][7] ,
         \update_mask_0/reg_out[6][8] , \update_mask_0/reg_out[6][9] ,
         \update_mask_0/reg_out[6][10] , \update_mask_0/reg_out[6][11] ,
         \update_mask_0/reg_out[6][12] , \update_mask_0/reg_out[6][13] ,
         \update_mask_0/reg_out[6][14] , \update_mask_0/reg_out[6][15] ,
         \update_mask_0/reg_out[6][16] , \update_mask_0/reg_out[6][17] ,
         \update_mask_0/reg_out[6][18] , \update_mask_0/reg_out[6][19] ,
         \update_mask_0/reg_out[7][0] , \update_mask_0/reg_out[7][1] ,
         \update_mask_0/reg_out[7][2] , \update_mask_0/reg_out[7][3] ,
         \update_mask_0/reg_out[7][4] , \update_mask_0/reg_out[7][5] ,
         \update_mask_0/reg_out[7][6] , \update_mask_0/reg_out[7][7] ,
         \update_mask_0/reg_out[7][8] , \update_mask_0/reg_out[7][9] ,
         \update_mask_0/reg_out[7][10] , \update_mask_0/reg_out[7][11] ,
         \update_mask_0/reg_out[7][12] , \update_mask_0/reg_out[7][13] ,
         \update_mask_0/reg_out[7][14] , \update_mask_0/reg_out[7][15] ,
         \update_mask_0/reg_out[7][16] , \update_mask_0/reg_out[7][17] ,
         \update_mask_0/reg_out[7][18] , \update_mask_0/reg_out[7][19] ,
         \update_mask_0/reg_out[8][0] , \update_mask_0/reg_out[8][1] ,
         \update_mask_0/reg_out[8][2] , \update_mask_0/reg_out[8][3] ,
         \update_mask_0/reg_out[8][4] , \update_mask_0/reg_out[8][5] ,
         \update_mask_0/reg_out[8][6] , \update_mask_0/reg_out[8][7] ,
         \update_mask_0/reg_out[8][8] , \update_mask_0/reg_out[8][9] ,
         \update_mask_0/reg_out[8][10] , \update_mask_0/reg_out[8][11] ,
         \update_mask_0/reg_out[8][12] , \update_mask_0/reg_out[8][13] ,
         \update_mask_0/reg_out[8][14] , \update_mask_0/reg_out[8][15] ,
         \update_mask_0/reg_out[8][16] , \update_mask_0/reg_out[8][17] ,
         \update_mask_0/reg_out[8][18] , \update_mask_0/reg_out[8][19] ,
         \update_mask_0/reg_out[9][0] , \update_mask_0/reg_out[9][1] ,
         \update_mask_0/reg_out[9][2] , \update_mask_0/reg_out[9][3] ,
         \update_mask_0/reg_out[9][4] , \update_mask_0/reg_out[9][5] ,
         \update_mask_0/reg_out[9][6] , \update_mask_0/reg_out[9][7] ,
         \update_mask_0/reg_out[9][8] , \update_mask_0/reg_out[9][9] ,
         \update_mask_0/reg_out[9][10] , \update_mask_0/reg_out[9][11] ,
         \update_mask_0/reg_out[9][12] , \update_mask_0/reg_out[9][13] ,
         \update_mask_0/reg_out[9][14] , \update_mask_0/reg_out[9][15] ,
         \update_mask_0/reg_out[9][16] , \update_mask_0/reg_out[9][17] ,
         \update_mask_0/reg_out[9][18] , \update_mask_0/reg_out[9][19] ,
         \update_mask_0/reg_out[10][0] , \update_mask_0/reg_out[10][1] ,
         \update_mask_0/reg_out[10][2] , \update_mask_0/reg_out[10][3] ,
         \update_mask_0/reg_out[10][4] , \update_mask_0/reg_out[10][5] ,
         \update_mask_0/reg_out[10][6] , \update_mask_0/reg_out[10][7] ,
         \update_mask_0/reg_out[10][8] , \update_mask_0/reg_out[10][9] ,
         \update_mask_0/reg_out[10][10] , \update_mask_0/reg_out[10][11] ,
         \update_mask_0/reg_out[10][12] , \update_mask_0/reg_out[10][13] ,
         \update_mask_0/reg_out[10][14] , \update_mask_0/reg_out[10][15] ,
         \update_mask_0/reg_out[10][16] , \update_mask_0/reg_out[10][17] ,
         \update_mask_0/reg_out[10][18] , \update_mask_0/reg_out[10][19] ,
         \update_mask_0/reg_out[11][0] , \update_mask_0/reg_out[11][1] ,
         \update_mask_0/reg_out[11][2] , \update_mask_0/reg_out[11][3] ,
         \update_mask_0/reg_out[11][4] , \update_mask_0/reg_out[11][5] ,
         \update_mask_0/reg_out[11][6] , \update_mask_0/reg_out[11][7] ,
         \update_mask_0/reg_out[11][8] , \update_mask_0/reg_out[11][9] ,
         \update_mask_0/reg_out[11][10] , \update_mask_0/reg_out[11][11] ,
         \update_mask_0/reg_out[11][12] , \update_mask_0/reg_out[11][13] ,
         \update_mask_0/reg_out[11][14] , \update_mask_0/reg_out[11][15] ,
         \update_mask_0/reg_out[11][16] , \update_mask_0/reg_out[11][17] ,
         \update_mask_0/reg_out[11][18] , \update_mask_0/reg_out[11][19] ,
         \update_mask_0/reg_out[12][0] , \update_mask_0/reg_out[12][1] ,
         \update_mask_0/reg_out[12][2] , \update_mask_0/reg_out[12][3] ,
         \update_mask_0/reg_out[12][4] , \update_mask_0/reg_out[12][5] ,
         \update_mask_0/reg_out[12][6] , \update_mask_0/reg_out[12][7] ,
         \update_mask_0/reg_out[12][8] , \update_mask_0/reg_out[12][9] ,
         \update_mask_0/reg_out[12][10] , \update_mask_0/reg_out[12][11] ,
         \update_mask_0/reg_out[12][12] , \update_mask_0/reg_out[12][13] ,
         \update_mask_0/reg_out[12][14] , \update_mask_0/reg_out[12][15] ,
         \update_mask_0/reg_out[12][16] , \update_mask_0/reg_out[12][17] ,
         \update_mask_0/reg_out[12][18] , \update_mask_0/reg_out[12][19] ,
         \update_mask_0/reg_out[13][0] , \update_mask_0/reg_out[13][1] ,
         \update_mask_0/reg_out[13][2] , \update_mask_0/reg_out[13][3] ,
         \update_mask_0/reg_out[13][4] , \update_mask_0/reg_out[13][5] ,
         \update_mask_0/reg_out[13][6] , \update_mask_0/reg_out[13][7] ,
         \update_mask_0/reg_out[13][8] , \update_mask_0/reg_out[13][9] ,
         \update_mask_0/reg_out[13][10] , \update_mask_0/reg_out[13][11] ,
         \update_mask_0/reg_out[13][12] , \update_mask_0/reg_out[13][13] ,
         \update_mask_0/reg_out[13][14] , \update_mask_0/reg_out[13][15] ,
         \update_mask_0/reg_out[13][16] , \update_mask_0/reg_out[13][17] ,
         \update_mask_0/reg_out[13][18] , \update_mask_0/reg_out[13][19] ,
         \update_mask_0/reg_out[14][0] , \update_mask_0/reg_out[14][1] ,
         \update_mask_0/reg_out[14][2] , \update_mask_0/reg_out[14][3] ,
         \update_mask_0/reg_out[14][4] , \update_mask_0/reg_out[14][5] ,
         \update_mask_0/reg_out[14][6] , \update_mask_0/reg_out[14][7] ,
         \update_mask_0/reg_out[14][8] , \update_mask_0/reg_out[14][9] ,
         \update_mask_0/reg_out[14][10] , \update_mask_0/reg_out[14][11] ,
         \update_mask_0/reg_out[14][12] , \update_mask_0/reg_out[14][13] ,
         \update_mask_0/reg_out[14][14] , \update_mask_0/reg_out[14][15] ,
         \update_mask_0/reg_out[14][16] , \update_mask_0/reg_out[14][17] ,
         \update_mask_0/reg_out[14][18] , \update_mask_0/reg_out[14][19] ,
         \update_mask_0/reg_out[15][0] , \update_mask_0/reg_out[15][1] ,
         \update_mask_0/reg_out[15][2] , \update_mask_0/reg_out[15][3] ,
         \update_mask_0/reg_out[15][4] , \update_mask_0/reg_out[15][5] ,
         \update_mask_0/reg_out[15][6] , \update_mask_0/reg_out[15][7] ,
         \update_mask_0/reg_out[15][8] , \update_mask_0/reg_out[15][9] ,
         \update_mask_0/reg_out[15][10] , \update_mask_0/reg_out[15][11] ,
         \update_mask_0/reg_out[15][12] , \update_mask_0/reg_out[15][13] ,
         \update_mask_0/reg_out[15][14] , \update_mask_0/reg_out[15][15] ,
         \update_mask_0/reg_out[15][16] , \update_mask_0/reg_out[15][17] ,
         \update_mask_0/reg_out[15][18] , \update_mask_0/reg_out[15][19] ,
         \update_mask_0/reg_i_mask[0] , \update_mask_0/reg_i_mask[1] ,
         \update_mask_0/reg_i_mask[2] , \update_mask_0/reg_i_mask[3] ,
         \update_mask_0/reg_i_mask[4] , \update_mask_0/reg_i_mask[5] ,
         \update_mask_0/reg_i_mask[6] , \update_mask_0/reg_i_mask[7] ,
         \update_mask_0/reg_i_mask[8] , \update_mask_0/reg_i_mask[9] ,
         \update_mask_0/reg_i_mask[10] , \update_mask_0/reg_i_mask[11] ,
         \update_mask_0/reg_i_mask[12] , \update_mask_0/reg_i_mask[13] ,
         \update_mask_0/reg_i_mask[14] , \update_mask_0/reg_i_mask[15] ,
         \update_mask_0/reg_i_mask[16] , \update_mask_0/reg_i_mask[17] ,
         \update_mask_0/reg_i_mask[18] , \update_mask_0/reg_i_mask[19] ,
         \update_mask_0/reg_i_mask[20] , \update_mask_0/reg_i_mask[21] ,
         \update_mask_0/reg_i_mask[22] , \update_mask_0/reg_i_mask[23] ,
         \update_mask_0/reg_i_mask[24] , \update_mask_0/reg_i_mask[25] ,
         \update_mask_0/reg_i_mask[26] , \update_mask_0/reg_i_mask[27] ,
         \update_mask_0/reg_i_mask[28] , \update_mask_0/reg_i_mask[29] ,
         \update_mask_0/reg_i_mask[30] , \update_mask_0/reg_i_mask[31] ,
         \update_mask_0/n2986 , \update_mask_0/N31 , \update_mask_0/N30 ,
         \update_mask_0/N29 , \update_mask_0/N28 , \update_mask_0/N27 ,
         \update_mask_0/N26 , \update_mask_0/N25 , \update_mask_0/N24 ,
         \update_mask_0/N23 , \update_output_0/n3151 , \update_output_0/n3150 ,
         \update_output_0/n3149 , \update_output_0/n3148 ,
         \update_output_0/n3147 , \update_output_0/n3146 ,
         \update_output_0/n3145 , \update_output_0/n3144 ,
         \update_output_0/n3143 , \update_output_0/n3142 ,
         \update_output_0/n3141 , \update_output_0/n3140 ,
         \update_output_0/n3139 , \update_output_0/n3138 ,
         \update_output_0/n3137 , \update_output_0/n3136 ,
         \update_output_0/n3135 , \update_output_0/n3134 ,
         \update_output_0/n3133 , \update_output_0/n3132 ,
         \update_output_0/n3131 , \update_output_0/n3130 ,
         \update_output_0/n3129 , \update_output_0/n3128 ,
         \update_output_0/n3127 , \update_output_0/n3126 ,
         \update_output_0/n3125 , \update_output_0/n3124 ,
         \update_output_0/n3123 , \update_output_0/n3122 ,
         \update_output_0/n3121 , \update_output_0/n3120 ,
         \update_output_0/n3119 , \update_output_0/n3118 ,
         \update_output_0/n3117 , \update_output_0/n3116 ,
         \update_output_0/n3115 , \update_output_0/n3114 ,
         \update_output_0/n3113 , \update_output_0/n3112 ,
         \update_output_0/n3111 , \update_output_0/n3110 ,
         \update_output_0/n3109 , \update_output_0/n3108 ,
         \update_output_0/n3107 , \update_output_0/n3106 ,
         \update_output_0/n3105 , \update_output_0/n3104 ,
         \update_output_0/n3103 , \update_output_0/n3102 ,
         \update_output_0/n3101 , \update_output_0/n3100 ,
         \update_output_0/n3099 , \update_output_0/n3098 ,
         \update_output_0/n3097 , \update_output_0/n3096 ,
         \update_output_0/n3095 , \update_output_0/n3094 ,
         \update_output_0/n3093 , \update_output_0/n3092 ,
         \update_output_0/n3091 , \update_output_0/n3090 ,
         \update_output_0/n3089 , \update_output_0/n3088 ,
         \update_output_0/n3087 , \update_output_0/n3086 ,
         \update_output_0/n3085 , \update_output_0/n3084 ,
         \update_output_0/n3083 , \update_output_0/n3082 ,
         \update_output_0/n3081 , \update_output_0/n3080 ,
         \update_output_0/n3079 , \update_output_0/n3078 ,
         \update_output_0/n3077 , \update_output_0/n3076 ,
         \update_output_0/n3075 , \update_output_0/n3074 ,
         \update_output_0/n3073 , \update_output_0/n3072 ,
         \update_output_0/n3071 , \update_output_0/n3070 ,
         \update_output_0/n3069 , \update_output_0/n3068 ,
         \update_output_0/n3067 , \update_output_0/n3066 ,
         \update_output_0/n3065 , \update_output_0/n3064 ,
         \update_output_0/n3063 , \update_output_0/n3062 ,
         \update_output_0/n3061 , \update_output_0/n3060 ,
         \update_output_0/n3059 , \update_output_0/n3058 ,
         \update_output_0/n3057 , \update_output_0/n3056 ,
         \update_output_0/n3055 , \update_output_0/n3054 ,
         \update_output_0/n3053 , \update_output_0/n3052 ,
         \update_output_0/n3051 , \update_output_0/n3050 ,
         \update_output_0/n3049 , \update_output_0/n3048 ,
         \update_output_0/n3047 , \update_output_0/n3046 ,
         \update_output_0/n3045 , \update_output_0/n3044 ,
         \update_output_0/n3043 , \update_output_0/n3042 ,
         \update_output_0/n3041 , \update_output_0/n3040 ,
         \update_output_0/n3039 , \update_output_0/n3038 ,
         \update_output_0/n3037 , \update_output_0/n3036 ,
         \update_output_0/n3035 , \update_output_0/n3034 ,
         \update_output_0/n3033 , \update_output_0/n3032 ,
         \update_output_0/n3031 , \update_output_0/n3030 ,
         \update_output_0/n3029 , \update_output_0/n3028 ,
         \update_output_0/n3027 , \update_output_0/n3026 ,
         \update_output_0/n3025 , \update_output_0/n3024 ,
         \update_output_0/n3023 , \update_output_0/n3022 ,
         \update_output_0/n3021 , \update_output_0/n3020 ,
         \update_output_0/n3019 , \update_output_0/n3018 ,
         \update_output_0/n3017 , \update_output_0/n3016 ,
         \update_output_0/n3015 , \update_output_0/n3014 ,
         \update_output_0/n3013 , \update_output_0/n3012 ,
         \update_output_0/n3011 , \update_output_0/n3010 ,
         \update_output_0/n3009 , \update_output_0/n3008 ,
         \update_output_0/n3007 , \update_output_0/n3006 ,
         \update_output_0/n3005 , \update_output_0/n3004 ,
         \update_output_0/n3003 , \update_output_0/n3002 ,
         \update_output_0/n3001 , \update_output_0/n3000 ,
         \update_output_0/n2999 , \update_output_0/n2998 ,
         \update_output_0/n2997 , \update_output_0/n2996 ,
         \update_output_0/n2995 , \update_output_0/n2994 ,
         \update_output_0/n2993 , \update_output_0/n2992 ,
         \update_output_0/n2991 , \update_output_0/n2990 ,
         \update_output_0/n2989 , \update_output_0/n2988 ,
         \update_output_0/n2987 , \update_output_0/n2986 ,
         \update_output_0/n2985 , \update_output_0/n2984 ,
         \update_output_0/n2983 , \update_output_0/n2982 ,
         \update_output_0/n2981 , \update_output_0/n2980 ,
         \update_output_0/n2979 , \update_output_0/n2978 ,
         \update_output_0/n2977 , \update_output_0/n2976 ,
         \update_output_0/n2975 , \update_output_0/n2974 ,
         \update_output_0/n2973 , \update_output_0/n2972 ,
         \update_output_0/n2971 , \update_output_0/n2970 ,
         \update_output_0/n2969 , \update_output_0/n2968 ,
         \update_output_0/n2967 , \update_output_0/n2966 ,
         \update_output_0/n2965 , \update_output_0/n2964 ,
         \update_output_0/n2963 , \update_output_0/n2962 ,
         \update_output_0/n2961 , \update_output_0/n2960 ,
         \update_output_0/n2959 , \update_output_0/n2958 ,
         \update_output_0/n2957 , \update_output_0/n2956 ,
         \update_output_0/n2955 , \update_output_0/n2954 ,
         \update_output_0/n2953 , \update_output_0/n2952 ,
         \update_output_0/n2951 , \update_output_0/n2950 ,
         \update_output_0/n2949 , \update_output_0/n2948 ,
         \update_output_0/n2947 , \update_output_0/n2946 ,
         \update_output_0/n2945 , \update_output_0/n2944 ,
         \update_output_0/n2943 , \update_output_0/n2942 ,
         \update_output_0/n2941 , \update_output_0/n2940 ,
         \update_output_0/n2939 , \update_output_0/n2938 ,
         \update_output_0/n2937 , \update_output_0/n2936 ,
         \update_output_0/n2935 , \update_output_0/n2934 ,
         \update_output_0/n2933 , \update_output_0/n2932 ,
         \update_output_0/n2931 , \update_output_0/n2930 ,
         \update_output_0/n2929 , \update_output_0/n2928 ,
         \update_output_0/n2927 , \update_output_0/n2926 ,
         \update_output_0/n2925 , \update_output_0/n2924 ,
         \update_output_0/n2923 , \update_output_0/n2922 ,
         \update_output_0/n2921 , \update_output_0/n2920 ,
         \update_output_0/n2919 , \update_output_0/n2918 ,
         \update_output_0/n2917 , \update_output_0/n2916 ,
         \update_output_0/n2915 , \update_output_0/n2914 ,
         \update_output_0/n2913 , \update_output_0/n2912 ,
         \update_output_0/n2911 , \update_output_0/n2910 ,
         \update_output_0/n2909 , \update_output_0/n2908 ,
         \update_output_0/n2907 , \update_output_0/n2906 ,
         \update_output_0/n2905 , \update_output_0/n2904 ,
         \update_output_0/n2903 , \update_output_0/n2902 ,
         \update_output_0/n2901 , \update_output_0/n2900 ,
         \update_output_0/n2899 , \update_output_0/n2898 ,
         \update_output_0/n2897 , \update_output_0/n2896 ,
         \update_output_0/n2895 , \update_output_0/n2894 ,
         \update_output_0/n2893 , \update_output_0/n2892 ,
         \update_output_0/n2891 , \update_output_0/n2890 ,
         \update_output_0/n2889 , \update_output_0/n2888 ,
         \update_output_0/n2887 , \update_output_0/n2886 ,
         \update_output_0/n2885 , \update_output_0/n2884 ,
         \update_output_0/n2883 , \update_output_0/n2882 ,
         \update_output_0/n2881 , \update_output_0/n2880 ,
         \update_output_0/n2879 , \update_output_0/n2878 ,
         \update_output_0/n2877 , \update_output_0/n2876 ,
         \update_output_0/n2875 , \update_output_0/n2874 ,
         \update_output_0/n2873 , \update_output_0/n2872 ,
         \update_output_0/n2871 , \update_output_0/n2870 ,
         \update_output_0/n2869 , \update_output_0/n2868 ,
         \update_output_0/n2867 , \update_output_0/n2866 ,
         \update_output_0/n2865 , \update_output_0/n2864 ,
         \update_output_0/n2863 , \update_output_0/n2862 ,
         \update_output_0/n2861 , \update_output_0/n2860 ,
         \update_output_0/n2859 , \update_output_0/n2858 ,
         \update_output_0/n2857 , \update_output_0/n2856 ,
         \update_output_0/n2855 , \update_output_0/n2854 ,
         \update_output_0/n2853 , \update_output_0/n2852 ,
         \update_output_0/n2851 , \update_output_0/n2850 ,
         \update_output_0/n2849 , \update_output_0/n2848 ,
         \update_output_0/n2847 , \update_output_0/n2846 ,
         \update_output_0/n2845 , \update_output_0/n2844 ,
         \update_output_0/n2843 , \update_output_0/n2842 ,
         \update_output_0/n2841 , \update_output_0/n2840 ,
         \update_output_0/n2839 , \update_output_0/n2838 ,
         \update_output_0/n2837 , \update_output_0/n2836 ,
         \update_output_0/n2835 , \update_output_0/n2834 ,
         \update_output_0/n2833 , \update_output_0/n2832 ,
         \update_output_0/n2831 , \update_output_0/n2830 ,
         \update_output_0/n2829 , \update_output_0/n2828 ,
         \update_output_0/n2827 , \update_output_0/n2826 ,
         \update_output_0/n2825 , \update_output_0/n2824 ,
         \update_output_0/n2823 , \update_output_0/n2822 ,
         \update_output_0/n2821 , \update_output_0/pre_o_im[13][19] ,
         \update_output_0/pre_o_im[13][18] ,
         \update_output_0/pre_o_im[13][17] ,
         \update_output_0/pre_o_im[13][16] ,
         \update_output_0/pre_o_im[13][15] ,
         \update_output_0/pre_o_im[13][14] ,
         \update_output_0/pre_o_im[13][13] ,
         \update_output_0/pre_o_im[13][12] ,
         \update_output_0/pre_o_im[13][11] ,
         \update_output_0/pre_o_im[13][10] , \update_output_0/pre_o_im[13][9] ,
         \update_output_0/pre_o_im[13][8] , \update_output_0/pre_o_im[13][7] ,
         \update_output_0/pre_o_im[13][6] , \update_output_0/pre_o_im[13][5] ,
         \update_output_0/pre_o_im[13][4] , \update_output_0/pre_o_im[13][3] ,
         \update_output_0/pre_o_im[13][2] , \update_output_0/pre_o_im[13][1] ,
         \update_output_0/pre_o_im[13][0] , \update_output_0/pre_o_im[12][19] ,
         \update_output_0/pre_o_im[12][18] ,
         \update_output_0/pre_o_im[12][17] ,
         \update_output_0/pre_o_im[12][16] ,
         \update_output_0/pre_o_im[12][15] ,
         \update_output_0/pre_o_im[12][14] ,
         \update_output_0/pre_o_im[12][13] ,
         \update_output_0/pre_o_im[12][12] ,
         \update_output_0/pre_o_im[12][11] ,
         \update_output_0/pre_o_im[12][10] , \update_output_0/pre_o_im[12][9] ,
         \update_output_0/pre_o_im[12][8] , \update_output_0/pre_o_im[12][7] ,
         \update_output_0/pre_o_im[12][6] , \update_output_0/pre_o_im[12][5] ,
         \update_output_0/pre_o_im[12][4] , \update_output_0/pre_o_im[12][3] ,
         \update_output_0/pre_o_im[12][2] , \update_output_0/pre_o_im[12][1] ,
         \update_output_0/pre_o_im[12][0] , \update_output_0/pre_o_im[4][19] ,
         \update_output_0/pre_o_im[4][18] , \update_output_0/pre_o_im[4][17] ,
         \update_output_0/pre_o_im[4][16] , \update_output_0/pre_o_im[4][15] ,
         \update_output_0/pre_o_im[4][14] , \update_output_0/pre_o_im[4][13] ,
         \update_output_0/pre_o_im[4][12] , \update_output_0/pre_o_im[4][11] ,
         \update_output_0/pre_o_im[4][10] , \update_output_0/pre_o_im[4][9] ,
         \update_output_0/pre_o_im[4][8] , \update_output_0/pre_o_im[4][7] ,
         \update_output_0/pre_o_im[4][6] , \update_output_0/pre_o_im[4][5] ,
         \update_output_0/pre_o_im[4][4] , \update_output_0/pre_o_im[4][3] ,
         \update_output_0/pre_o_im[4][2] , \update_output_0/pre_o_im[4][1] ,
         \update_output_0/pre_o_im[4][0] , \update_output_0/n6096 ,
         \update_output_0/N34 , \update_output_0/N33 , \update_output_0/N32 ,
         \update_output_0/N31 , \update_output_0/N30 , \update_output_0/N29 ,
         \update_output_0/N28 , \update_output_0/N27 , n3432, n3433, n3434,
         n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445,
         n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455,
         n3456, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467,
         n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477,
         n3478, n3479, n3480, n3481, n3482, n3484, n3485, n3486, n3487, n3488,
         n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498,
         n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508,
         n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518,
         n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3528, n3529,
         n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539,
         n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549,
         n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559,
         n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569,
         n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580,
         n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590,
         n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600,
         n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610,
         n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620,
         n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630,
         n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640,
         n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650,
         n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660,
         n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670,
         n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680,
         n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690,
         n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3700, n3701,
         n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711,
         n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721,
         n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731,
         n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741,
         n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751,
         n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761,
         n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771,
         n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781,
         n3782, n3783, n3784, n3785, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3830, n3831, n3832, n3833,
         n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843,
         n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853,
         n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863,
         n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3873, n3874,
         n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884,
         n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894,
         n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904,
         n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3915,
         n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925,
         n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935,
         n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945,
         n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955,
         n3956, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966,
         n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976,
         n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986,
         n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996,
         n3997, n3998, n3999, n4001, n4002, n4003, n4004, n4005, n4006, n4007,
         n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017,
         n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027,
         n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037,
         n4038, n4039, n4040, n4041, n4042, n4044, n4045, n4046, n4047, n4048,
         n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058,
         n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068,
         n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078,
         n4079, n4080, n4081, n4082, n4083, n4084, n4086, n4087, n4088, n4089,
         n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099,
         n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109,
         n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119,
         n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4130,
         n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140,
         n4141, n4142, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151,
         n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161,
         n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171,
         n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181,
         n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191,
         n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201,
         n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211,
         n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221,
         n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231,
         n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241,
         n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251,
         n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261,
         n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271,
         n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281,
         n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291,
         n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301,
         n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311,
         n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321,
         n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331,
         n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341,
         n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4533,
         n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543,
         n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553,
         n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563,
         n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573,
         n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583,
         n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593,
         n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603,
         n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
         n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
         n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
         n4635, n4636, n4637, n4638, n4639, n4641, n4642, n4643, n4644, n4645,
         n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655,
         n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665,
         n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675,
         n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685,
         n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695,
         n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705,
         n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715,
         n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725,
         n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735,
         n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745,
         n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755,
         n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765,
         n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775,
         n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785,
         n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795,
         n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805,
         n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815,
         n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825,
         n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835,
         n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845,
         n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855,
         n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4865, n4866,
         n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876,
         n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886,
         n4887, n4888, n4889, n4890, n4892, n4893, n4894, n4895, n4896, n4897,
         n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907,
         n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917,
         n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927,
         n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937,
         n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947,
         n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957,
         n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967,
         n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977,
         n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987,
         n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997,
         n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007,
         n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017,
         n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027,
         n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037,
         n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047,
         n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057,
         n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067,
         n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077,
         n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087,
         n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097,
         n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107,
         n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117,
         n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127,
         n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137,
         n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147,
         n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157,
         n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167,
         n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177,
         n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187,
         n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197,
         n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207,
         n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217,
         n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227,
         n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237,
         n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247,
         n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257,
         n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267,
         n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277,
         n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287,
         n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297,
         n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307,
         n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317,
         n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327,
         n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337,
         n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347,
         n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357,
         n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367,
         n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377,
         n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387,
         n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397,
         n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407,
         n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417,
         n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427,
         n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437,
         n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447,
         n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457,
         n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467,
         n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477,
         n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487,
         n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497,
         n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507,
         n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517,
         n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527,
         n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537,
         n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547,
         n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557,
         n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567,
         n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577,
         n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587,
         n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597,
         n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607,
         n5608, n5609, n5610, n5611, n5612, n5614, n5615, n5616, n5617, n5618,
         n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628,
         n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638,
         n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648,
         n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658,
         n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668,
         n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678,
         n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688,
         n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698,
         n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708,
         n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718,
         n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728,
         n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738,
         n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748,
         n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758,
         n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768,
         n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778,
         n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788,
         n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798,
         n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808,
         n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818,
         n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828,
         n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838,
         n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848,
         n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858,
         n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868,
         n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878,
         n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888,
         n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898,
         n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908,
         n5909, n5910, n5911, \update_output_0/n2819 , \update_output_0/n2818 ,
         \update_output_0/n2815 , \update_output_0/n2814 ,
         \update_output_0/n2811 , \update_output_0/n2810 ,
         \update_output_0/n2807 , \update_output_0/n2806 ,
         \update_output_0/n2803 , \update_output_0/n2802 ,
         \update_output_0/n2799 , \update_output_0/n2798 ,
         \update_output_0/n2795 , \update_output_0/n2794 ,
         \update_output_0/n2791 , \update_output_0/n2790 ,
         \update_output_0/n2787 , \update_output_0/n2786 ,
         \update_output_0/n2783 , \update_output_0/n2782 ,
         \update_output_0/n2779 , \update_output_0/n2778 ,
         \update_output_0/n2775 , \update_output_0/n2774 ,
         \update_output_0/n2771 , \update_output_0/n2770 ,
         \update_output_0/n2767 , \update_output_0/n2766 ,
         \update_output_0/n2763 , \update_output_0/n2762 ,
         \update_output_0/n2759 , \update_output_0/n2758 ,
         \update_output_0/n2755 , \update_output_0/n2754 ,
         \update_output_0/n2751 , \update_output_0/n2750 ,
         \update_output_0/n2747 , \update_output_0/n2746 ,
         \update_output_0/n2743 , \update_output_0/n2742 ,
         \update_output_0/n2739 , \update_output_0/n2738 ,
         \update_output_0/n2735 , \update_output_0/n2734 ,
         \update_output_0/n2731 , \update_output_0/n2730 ,
         \update_output_0/n2727 , \update_output_0/n2726 ,
         \update_output_0/n2723 , \update_output_0/n2722 ,
         \update_output_0/n2719 , \update_output_0/n2718 ,
         \update_output_0/n2715 , \update_output_0/n2714 ,
         \update_output_0/n2711 , \update_output_0/n2710 ,
         \update_output_0/n2707 , \update_output_0/n2706 ,
         \update_output_0/n2703 , \update_output_0/n2702 ,
         \update_output_0/n2699 , \update_output_0/n2698 ,
         \update_output_0/n2695 , \update_output_0/n2694 ,
         \update_output_0/n2691 , \update_output_0/n2690 ,
         \update_output_0/n2687 , \update_output_0/n2686 ,
         \update_output_0/n2683 , \update_output_0/n2682 ,
         \update_output_0/n2679 , \update_output_0/n2678 ,
         \update_output_0/n2675 , \update_output_0/n2674 ,
         \update_output_0/n2671 , \update_output_0/n2670 ,
         \update_output_0/n2667 , \update_output_0/n2666 ,
         \update_output_0/n2663 , \update_output_0/n2662 ,
         \update_output_0/n2659 , \update_output_0/n2658 ,
         \update_output_0/n2655 , \update_output_0/n2654 ,
         \update_output_0/n2651 , \update_output_0/n2650 ,
         \update_output_0/n2647 , \update_output_0/n2646 ,
         \update_output_0/n2643 , \update_output_0/n2642 ,
         \update_output_0/n2639 , \update_output_0/n2638 ,
         \update_output_0/n2635 , \update_output_0/n2634 ,
         \update_output_0/n2631 , \update_output_0/n2630 ,
         \update_output_0/n2627 , \update_output_0/n2626 ,
         \update_output_0/n2623 , \update_output_0/n2622 ,
         \update_output_0/n2619 , \update_output_0/n2618 ,
         \update_output_0/n2615 , \update_output_0/n2614 ,
         \update_output_0/n2611 , \update_output_0/n2610 ,
         \update_output_0/n2607 , \update_output_0/n2606 ,
         \update_output_0/n2603 , \update_output_0/n2602 ,
         \update_output_0/n2599 , \update_output_0/n2598 ,
         \update_output_0/n2595 , \update_output_0/n2594 ,
         \update_output_0/n2591 , \update_output_0/n2590 ,
         \update_output_0/n2587 , \update_output_0/n2586 ,
         \update_output_0/n2583 , \update_output_0/n2582 ,
         \update_output_0/n2579 , \update_output_0/n2578 ,
         \update_output_0/n2575 , \update_output_0/n2574 ,
         \update_output_0/n2571 , \update_output_0/n2570 ,
         \update_output_0/n2567 , \update_output_0/n2566 ,
         \update_output_0/n2563 , \update_output_0/n2562 ,
         \update_output_0/n2559 , \update_output_0/n2558 ,
         \update_output_0/n2555 , \update_output_0/n2554 ,
         \update_output_0/n2551 , \update_output_0/n2550 ,
         \update_output_0/n2547 , \update_output_0/n2546 ,
         \update_output_0/n2543 , \update_output_0/n2542 ,
         \update_output_0/n2539 , \update_output_0/n2538 ,
         \update_output_0/n2535 , \update_output_0/n2534 ,
         \update_output_0/n2531 , \update_output_0/n2530 ,
         \update_output_0/n2527 , \update_output_0/n2526 ,
         \update_output_0/n2523 , \update_output_0/n2522 ,
         \update_output_0/n2519 , \update_output_0/n2518 ,
         \update_output_0/n2515 , \update_output_0/n2514 ,
         \update_output_0/n2511 , \update_output_0/n2510 ,
         \update_output_0/n2507 , \update_output_0/n2506 ,
         \update_output_0/n2503 , \update_output_0/n2502 ,
         \update_output_0/n2499 , \update_output_0/n2498 ,
         \update_output_0/n2495 , \update_output_0/n2494 ,
         \update_output_0/n2491 , \update_output_0/n2490 ,
         \update_output_0/n2487 , \update_output_0/n2486 ,
         \update_output_0/n2483 , \update_output_0/n2482 ,
         \update_output_0/n2479 , \update_output_0/n2478 ,
         \update_output_0/n2475 , \update_output_0/n2474 ,
         \update_output_0/n2471 , \update_output_0/n2470 ,
         \update_output_0/n2467 , \update_output_0/n2466 ,
         \update_output_0/n2463 , \update_output_0/n2462 ,
         \update_output_0/n2459 , \update_output_0/n2458 ,
         \update_output_0/n2455 , \update_output_0/n2454 ,
         \update_output_0/n2451 , \update_output_0/n2450 ,
         \update_output_0/n2447 , \update_output_0/n2446 ,
         \update_output_0/n2443 , \update_output_0/n2442 ,
         \update_output_0/n2439 , \update_output_0/n2438 ,
         \update_output_0/n2435 , \update_output_0/n2434 ,
         \update_output_0/n2431 , \update_output_0/n2430 ,
         \update_output_0/n2427 , \update_output_0/n2426 ,
         \update_output_0/n2423 , \update_output_0/n2422 ,
         \update_output_0/n2419 , \update_output_0/n2418 ,
         \update_output_0/n2415 , \update_output_0/n2414 ,
         \update_output_0/n2411 , \update_output_0/n2410 ,
         \update_output_0/n2407 , \update_output_0/n2406 ,
         \update_output_0/n2403 , \update_output_0/n2402 ,
         \update_output_0/n2399 , \update_output_0/n2398 ,
         \update_output_0/n2395 , \update_output_0/n2394 ,
         \update_output_0/n2391 , \update_output_0/n2390 ,
         \update_output_0/n2387 , \update_output_0/n2386 ,
         \update_output_0/n2383 , \update_output_0/n2382 ,
         \update_output_0/n2379 , \update_output_0/n2378 ,
         \update_output_0/n2375 , \update_output_0/n2374 ,
         \update_output_0/n2371 , \update_output_0/n2370 ,
         \update_output_0/n2367 , \update_output_0/n2366 ,
         \update_output_0/n2363 , \update_output_0/n2362 ,
         \update_output_0/n2359 , \update_output_0/n2358 ,
         \update_output_0/n2355 , \update_output_0/n2354 ,
         \update_output_0/n2351 , \update_output_0/n2350 ,
         \update_output_0/n2347 , \update_output_0/n2346 ,
         \update_output_0/n2343 , \update_output_0/n2342 ,
         \update_output_0/n2339 , \update_output_0/n2338 ,
         \update_output_0/n2335 , \update_output_0/n2334 ,
         \update_output_0/n2331 , \update_output_0/n2330 ,
         \update_output_0/n2327 , \update_output_0/n2326 ,
         \update_output_0/n2323 , \update_output_0/n2322 ,
         \update_output_0/n2319 , \update_output_0/n2318 ,
         \update_output_0/n2315 , \update_output_0/n2314 ,
         \update_output_0/n2311 , \update_output_0/n2310 ,
         \update_output_0/n2307 , \update_output_0/n2306 ,
         \update_output_0/n2303 , \update_output_0/n2302 ,
         \update_output_0/n2299 , \update_output_0/n2298 ,
         \update_output_0/n2295 , \update_output_0/n2294 ,
         \update_output_0/n2291 , \update_output_0/n2290 ,
         \update_output_0/n2287 , \update_output_0/n2286 ,
         \update_output_0/n2283 , \update_output_0/n2282 ,
         \update_output_0/n2279 , \update_output_0/n2278 ,
         \update_output_0/n2275 , \update_output_0/n2274 ,
         \update_output_0/n2271 , \update_output_0/n2270 ,
         \update_output_0/n2267 , \update_output_0/n2266 ,
         \update_output_0/n2263 , \update_output_0/n2262 ,
         \update_output_0/n2259 , \update_output_0/n2258 ,
         \update_output_0/n2255 , \update_output_0/n2254 ,
         \update_output_0/n2251 , \update_output_0/n2250 ,
         \update_output_0/n2247 , \update_output_0/n2246 ,
         \update_output_0/n2243 , \update_output_0/n2242 ,
         \update_output_0/n2239 , \update_output_0/n2238 ,
         \update_output_0/n2235 , \update_output_0/n2234 ,
         \update_output_0/n2231 , \update_output_0/n2230 ,
         \update_output_0/n2227 , \update_output_0/n2226 ,
         \update_output_0/n2223 , \update_output_0/n2222 ,
         \update_output_0/n2219 , \update_output_0/n2218 ,
         \update_output_0/n2215 , \update_output_0/n2214 ,
         \update_output_0/n2211 , \update_output_0/n2210 ,
         \update_output_0/n2207 , \update_output_0/n2206 ,
         \update_output_0/n2203 , \update_output_0/n2202 ,
         \update_output_0/n2199 , \update_output_0/n2198 ,
         \update_output_0/n2195 , \update_output_0/n2194 ,
         \update_output_0/n2191 , \update_output_0/n2190 ,
         \update_output_0/n2187 , \update_output_0/n2186 ,
         \update_output_0/n2183 , \update_output_0/n2182 ,
         \update_output_0/n2179 , \update_output_0/n2178 ,
         \update_output_0/n2175 , \update_output_0/n2174 ,
         \update_output_0/n2171 , \update_output_0/n2170 ,
         \update_output_0/n2167 , \update_output_0/n2166 ,
         \update_output_0/n2163 , \update_output_0/n2162 ,
         \update_output_0/n2159 , \update_output_0/n2158 ,
         \update_output_0/n2155 , \update_output_0/n2154 ,
         \update_output_0/n2151 , \update_output_0/n2150 ,
         \update_output_0/n2147 , \update_output_0/n2146 ,
         \update_output_0/n2143 , \update_output_0/n2142 ,
         \update_output_0/n2139 , \update_output_0/n2138 ,
         \update_output_0/n2135 , \update_output_0/n2134 ,
         \update_output_0/n2131 , \update_output_0/n2130 ,
         \update_output_0/n2127 , \update_output_0/n2126 ,
         \update_output_0/n2123 , \update_output_0/n2122 ,
         \update_output_0/n2119 , \update_output_0/n2118 ,
         \update_output_0/n2115 , \update_output_0/n2114 ,
         \update_output_0/n2111 , \update_output_0/n2110 ,
         \update_output_0/n2107 , \update_output_0/n2106 ,
         \update_output_0/n2103 , \update_output_0/n2102 ,
         \update_output_0/n2099 , \update_output_0/n2098 ,
         \update_output_0/n2095 , \update_output_0/n2094 ,
         \update_output_0/n2091 , \update_output_0/n2090 ,
         \update_output_0/n2087 , \update_output_0/n2086 ,
         \update_output_0/n2083 , \update_output_0/n2082 ,
         \update_output_0/n2079 , \update_output_0/n2078 ,
         \update_output_0/n2075 , \update_output_0/n2074 ,
         \update_output_0/n2071 , \update_output_0/n2070 ,
         \update_output_0/n2067 , \update_output_0/n2066 ,
         \update_output_0/n2063 , \update_output_0/n2062 ,
         \update_output_0/n2059 , \update_output_0/n2058 ,
         \update_output_0/n2055 , \update_output_0/n2054 ,
         \update_output_0/n2051 , \update_output_0/n2050 ,
         \update_output_0/n2047 , \update_output_0/n2046 ,
         \update_output_0/n2043 , \update_output_0/n2042 ,
         \update_output_0/n2039 , \update_output_0/n2038 ,
         \update_output_0/n2035 , \update_output_0/n2034 ,
         \update_output_0/n2031 , \update_output_0/n2030 ,
         \update_output_0/n2027 , \update_output_0/n2026 ,
         \update_output_0/n2023 , \update_output_0/n2022 ,
         \update_output_0/n2019 , \update_output_0/n2018 ,
         \update_output_0/n2015 , \update_output_0/n2014 ,
         \update_output_0/n2011 , \update_output_0/n2010 ,
         \update_output_0/n2007 , \update_output_0/n2006 ,
         \update_output_0/n2003 , \update_output_0/n2002 ,
         \update_output_0/n1999 , \update_output_0/n1998 ,
         \update_output_0/n1995 , \update_output_0/n1994 ,
         \update_output_0/n1991 , \update_output_0/n1990 ,
         \update_output_0/n1987 , \update_output_0/n1986 ,
         \update_output_0/n1983 , \update_output_0/n1982 ,
         \update_output_0/n1979 , \update_output_0/n1978 ,
         \update_output_0/n1975 , \update_output_0/n1974 ,
         \update_output_0/n1971 , \update_output_0/n1970 ,
         \update_output_0/n1967 , \update_output_0/n1966 ,
         \update_output_0/n1963 , \update_output_0/n1962 ,
         \update_output_0/n1959 , \update_output_0/n1958 ,
         \update_output_0/n1955 , \update_output_0/n1954 ,
         \update_output_0/n1951 , \update_output_0/n1950 ,
         \update_output_0/n1947 , \update_output_0/n1946 ,
         \update_output_0/n1943 , \update_output_0/n1942 ,
         \update_output_0/n1939 , \update_output_0/n1938 ,
         \update_output_0/n1935 , \update_output_0/n1934 ,
         \update_output_0/n1931 , \update_output_0/n1930 ,
         \update_output_0/n1927 , \update_output_0/n1926 ,
         \update_output_0/n1923 , \update_output_0/n1922 ,
         \update_output_0/n1919 , \update_output_0/n1918 ,
         \update_output_0/n1915 , \update_output_0/n1914 ,
         \update_output_0/n1911 , \update_output_0/n1910 ,
         \update_output_0/n1907 , \update_output_0/n1906 ,
         \update_output_0/n1903 , \update_output_0/n1902 ,
         \update_output_0/n1899 , \update_output_0/n1898 ,
         \update_output_0/n1895 , \update_output_0/n1894 ,
         \update_output_0/n1891 , \update_output_0/n1890 ,
         \update_output_0/n1887 , \update_output_0/n1886 ,
         \update_output_0/n1883 , \update_output_0/n1882 ,
         \update_output_0/n1879 , \update_output_0/n1878 ,
         \update_output_0/n1875 , \update_output_0/n1874 ,
         \update_output_0/n1871 , \update_output_0/n1870 ,
         \update_output_0/n1867 , \update_output_0/n1866 ,
         \update_output_0/n1863 , \update_output_0/n1862 ,
         \update_output_0/n1859 , \update_output_0/n1858 ,
         \update_output_0/n1855 , \update_output_0/n1854 ,
         \update_output_0/n1851 , \update_output_0/n1850 ,
         \update_output_0/n1847 , \update_output_0/n1846 ,
         \update_output_0/n1843 , \update_output_0/n1842 ,
         \update_output_0/n1839 , \update_output_0/n1838 ,
         \update_output_0/n1835 , \update_output_0/n1834 ,
         \update_output_0/n1831 , \update_output_0/n1830 ,
         \update_output_0/n1827 , \update_output_0/n1826 ,
         \update_output_0/n1823 , \update_output_0/n1822 ,
         \update_output_0/n1819 , \update_output_0/n1818 ,
         \update_output_0/n1815 , \update_output_0/n1814 ,
         \update_output_0/n1811 , \update_output_0/n1810 ,
         \update_output_0/n1807 , \update_output_0/n1806 ,
         \update_output_0/n1803 , \update_output_0/n1802 ,
         \update_output_0/n1799 , \update_output_0/n1798 ,
         \update_output_0/n1795 , \update_output_0/n1794 ,
         \update_output_0/n1791 , \update_output_0/n1790 ,
         \update_output_0/n1787 , \update_output_0/n1786 ,
         \update_output_0/n1783 , \update_output_0/n1782 ,
         \update_output_0/n1779 , \update_output_0/n1778 ,
         \update_output_0/n1775 , \update_output_0/n1774 ,
         \update_output_0/n1771 , \update_output_0/n1770 ,
         \update_output_0/n1767 , \update_output_0/n1766 ,
         \update_output_0/n1763 , \update_output_0/n1762 ,
         \update_output_0/n1759 , \update_output_0/n1758 ,
         \update_output_0/n1755 , \update_output_0/n1754 ,
         \update_output_0/n1751 , \update_output_0/n1750 ,
         \update_output_0/n1747 , \update_output_0/n1746 ,
         \update_output_0/n1743 , \update_output_0/n1742 ,
         \update_output_0/n1739 , \update_output_0/n1738 ,
         \update_output_0/n1735 , \update_output_0/n1734 ,
         \update_output_0/n1731 , \update_output_0/n1730 ,
         \update_output_0/n1727 , \update_output_0/n1726 ,
         \update_output_0/n1723 , \update_output_0/n1722 ,
         \update_output_0/n1719 , \update_output_0/n1718 ,
         \update_output_0/n1715 , \update_output_0/n1714 ,
         \update_output_0/n1711 , \update_output_0/n1710 ,
         \update_output_0/n1707 , \update_output_0/n1706 ,
         \update_output_0/n1703 , \update_output_0/n1702 ,
         \update_output_0/n1699 , \update_output_0/n1698 ,
         \update_output_0/n1695 , \update_output_0/n1694 ,
         \update_output_0/n1691 , \update_output_0/n1690 ,
         \update_output_0/n1687 , \update_output_0/n1686 ,
         \update_output_0/n1683 , \update_output_0/n1682 ,
         \update_output_0/n1679 , \update_output_0/n1678 ,
         \update_output_0/n1675 , \update_output_0/n1674 ,
         \update_output_0/n1671 , \update_output_0/n1670 ,
         \update_output_0/n1667 , \update_output_0/n1666 ,
         \update_output_0/n1663 , \update_output_0/n1662 ,
         \update_output_0/n1659 , \update_output_0/n1658 ,
         \update_output_0/n1655 , \update_output_0/n1654 ,
         \update_output_0/n1651 , \update_output_0/n1650 ,
         \update_output_0/n1647 , \update_output_0/n1646 ,
         \update_output_0/n1643 , \update_output_0/n1642 ,
         \update_output_0/n1639 , \update_output_0/n1638 ,
         \update_output_0/n1635 , \update_output_0/n1634 ,
         \update_output_0/n1631 , \update_output_0/n1630 ,
         \update_output_0/n1627 , \update_output_0/n1626 ,
         \update_output_0/n1623 , \update_output_0/n1622 ,
         \update_output_0/n1619 , \update_output_0/n1618 ,
         \update_output_0/n1615 , \update_output_0/n1614 ,
         \update_output_0/n1611 , \update_output_0/n1610 ,
         \update_output_0/n1607 , \update_output_0/n1606 ,
         \update_output_0/n1603 , \update_output_0/n1602 ,
         \update_output_0/n1599 , \update_output_0/n1598 ,
         \update_output_0/n1595 , \update_output_0/n1594 ,
         \update_output_0/n1591 , \update_output_0/n1590 ,
         \update_output_0/n1587 , \update_output_0/n1586 ,
         \update_output_0/n1583 , \update_output_0/n1582 ,
         \update_output_0/n1579 , \update_output_0/n1578 ,
         \update_output_0/n1575 , \update_output_0/n1574 ,
         \update_output_0/n1571 , \update_output_0/n1570 ,
         \update_output_0/n1567 , \update_output_0/n1566 ,
         \update_output_0/n1563 , \update_output_0/n1562 ,
         \update_output_0/n1559 , \update_output_0/n1558 ,
         \update_output_0/n1555 , \update_output_0/n1554 ,
         \update_output_0/n1551 , \update_output_0/n1550 ,
         \update_output_0/n1547 , \update_output_0/n1546 ,
         \update_output_0/n1543 , \update_output_0/n1542 ,
         \update_output_0/n1539 , \update_output_0/n1538 ,
         \update_mask_0/n997 , \update_mask_0/n996 , \update_mask_0/n993 ,
         \update_mask_0/n992 , \update_mask_0/n989 , \update_mask_0/n988 ,
         \update_mask_0/n985 , \update_mask_0/n984 , \update_mask_0/n981 ,
         \update_mask_0/n980 , \update_mask_0/n977 , \update_mask_0/n976 ,
         \update_mask_0/n973 , \update_mask_0/n972 , \update_mask_0/n969 ,
         \update_mask_0/n968 , \update_mask_0/n965 , \update_mask_0/n964 ,
         \update_mask_0/n961 , \update_mask_0/n960 , \update_mask_0/n957 ,
         \update_mask_0/n956 , \update_mask_0/n952 , \update_mask_0/n949 ,
         \update_mask_0/n948 , \update_mask_0/n1077 , \update_mask_0/n1076 ,
         \update_mask_0/n1073 , \update_mask_0/n1072 , \update_mask_0/n1069 ,
         \update_mask_0/n1068 , \update_mask_0/n1065 , \update_mask_0/n1064 ,
         \update_mask_0/n1061 , \update_mask_0/n1060 , \update_mask_0/n1057 ,
         \update_mask_0/n1056 , \update_mask_0/n1053 , \update_mask_0/n1052 ,
         \update_mask_0/n1049 , \update_mask_0/n1048 , \update_mask_0/n1045 ,
         \update_mask_0/n1044 , \update_mask_0/n1041 , \update_mask_0/n1040 ,
         \update_mask_0/n1037 , \update_mask_0/n1036 , \update_mask_0/n1033 ,
         \update_mask_0/n1032 , \update_mask_0/n1029 , \update_mask_0/n1028 ,
         \update_mask_0/n1025 , \update_mask_0/n1024 , \update_mask_0/n1021 ,
         \update_mask_0/n1020 , \update_mask_0/n1017 , \update_mask_0/n1016 ,
         \update_mask_0/n1013 , \update_mask_0/n1012 , \update_mask_0/n1009 ,
         \update_mask_0/n1008 , \update_mask_0/n1005 , \update_mask_0/n1004 ,
         \update_mask_0/n1001 , \update_mask_0/n1000 , n999, n998, n997, n996,
         n995, n994, n993, n992, n991, n990, n989, n988, n987, n986, n985,
         n984, n983, n982, n981, n980, n979, n978, n977, n976, n975, n974,
         n973, n972, n971, n970, n969, n968, n967, n966, n965, n964, n963,
         n962, n961, n960, n959, n958, n957, n956, n955, n954, n953, n952,
         n951, n950, n949, n948, n947, n946, n945, n944, n943, n942, n941,
         n940, n939, n938, n937, n936, n935, n934, n933, n932, n931, n930,
         n929, n928, n927, n926, n925, n924, n923, n922, n921, n920, n919,
         n918, n917, n916, n915, n914, n913, n912, n911, n910, n909, n908,
         n907, n906, n905, n904, n903, n902, n901, n900, n899, n898, n897,
         n896, n895, n894, n893, n892, n891, n890, n889, n888, n887, n886,
         n885, n884, n883, n882, n881, n880, n879, n878, n877, n876, n875,
         n874, n873, n872, n871, n870, n869, n868, n867, n866, n865, n864,
         n863, n862, n861, n860, n859, n858, n857, n856, n855, n854, n853,
         n852, n851, n850, n849, n848, n847, n846, n845, n844, n843, n842,
         n841, n840, n839, n838, n837, n836, n835, n834, n833, n832, n831,
         n830, n829, n828, n827, n826, n825, n824, n823, n822, n821, n820,
         n819, n818, n817, n816, n815, n814, n813, n812, n811, n810, n809,
         n808, n807, n806, n805, n803, n802, n801, n800, n798, n796, n795,
         n793, n792, n791, n790, n789, n788, n787, n786, n785, n784, n783,
         n782, n781, n780, n779, n778, n777, n776, n775, n774, n773, n772,
         n771, n770, n769, n768, n767, n766, n765, n764, n763, n762, n761,
         n760, n759, n758, n757, n756, n755, n754, n753, n752, n751, n750,
         n749, n748, n747, n746, n745, n744, n743, n742, n741, n740, n739,
         n738, n737, n736, n735, n734, n733, n2265, n2264, n2263, n2262, n2261,
         n2260, n2259, n2258, n2257, n2256, n2255, n2254, n2253, n2252, n2251,
         n2250, n2249, n2248, n2247, n2246, n2245, n2244, n2243, n2242, n2241,
         n2240, n2239, n2238, n2237, n2236, n2235, n2234, n2233, n2232, n2231,
         n2230, n2229, n2228, n2227, n2226, n2225, n2224, n2223, n2222, n2221,
         n2220, n2219, n2218, n2217, n2216, n2215, n2214, n2213, n2212, n2211,
         n2210, n2209, n2208, n2207, n2206, n2205, n2204, n2203, n2202, n2201,
         n2200, n2199, n2198, n2197, n2196, n2195, n2194, n2193, n2192, n2191,
         n2190, n2189, n2188, n2187, n2186, n2185, n2184, n2183, n2182, n2181,
         n2180, n2179, n2178, n2177, n2176, n2175, n2174, n2173, n2172, n2171,
         n2170, n2169, n2168, n2167, n2166, n2165, n2164, n2163, n2162, n2161,
         n2160, n2159, n2158, n2157, n2156, n2155, n2154, n2153, n2152, n2151,
         n2150, n2149, n2148, n2147, n2146, n2145, n2144, n2143, n2142, n2141,
         n2140, n2139, n2138, n2137, n2136, n2135, n2134, n2133, n2132, n2131,
         n2130, n2129, n2128, n2127, n2126, n2125, n2124, n2123, n2122, n2121,
         n2120, n2119, n2118, n2117, n2116, n2115, n2114, n2113, n2112, n2111,
         n2110, n2109, n2108, n2107, n2106, n2105, n2104, n2103, n2102, n2101,
         n2100, n2099, n2098, n2097, n2096, n2095, n2094, n2093, n2092, n2091,
         n2090, n2089, n2088, n2087, n2086, n2085, n2084, n2083, n2082, n2081,
         n2080, n2079, n2078, n2077, n2076, n2075, n2074, n2073, n2072, n2071,
         n2070, n2069, n2068, n2067, n2066, n2065, n2064, n2063, n2062, n2061,
         n2060, n2059, n2058, n2057, n2056, n2055, n2054, n2053, n2052, n2051,
         n2050, n2049, n2048, n2047, n2046, n2045, n2044, n2043, n2042, n2041,
         n2040, n2039, n2038, n2037, n2036, n2035, n2034, n2033, n2032, n2031,
         n2030, n2029, n2028, n2027, n2026, n2025, n2024, n2023, n2022, n2021,
         n2020, n2019, n2018, n2017, n2016, n2015, n2014, n2013, n2012, n2011,
         n2010, n2009, n2008, n2007, n2006, n2005, n2004, n2003, n2002, n2001,
         n2000, n1999, n1998, n1997, n1996, n1995, n1994, n1993, n1992, n1991,
         n1990, n1989, n1988, n1987, n1986, n1985, n1984, n1983, n1982, n1981,
         n1980, n1979, n1978, n1977, n1976, n1975, n1974, n1973, n1972, n1971,
         n1970, n1969, n1968, n1967, n1966, n1965, n1964, n1963, n1962, n1961,
         n1960, n1959, n1958, n1957, n1956, n1955, n1954, n1953, n1952, n1951,
         n1950, n1949, n1948, n1947, n1946, n1945, n1944, n1943, n1942, n1941,
         n1940, n1939, n1938, n1937, n1936, n1935, n1934, n1933, n1932, n1931,
         n1930, n1929, n1928, n1927, n1926, n1925, n1924, n1923, n1922, n1921,
         n1920, n1919, n1918, n1917, n1916, n1915, n1914, n1913, n1912, n1911,
         n1910, n1909, n1908, n1907, n1906, n1905, n1904, n1903, n1902, n1901,
         n1900, n1899, n1898, n1897, n1896, n1895, n1894, n1893, n1892, n1891,
         n1890, n1889, n1888, n1887, n1886, n1885, n1884, n1883, n1882, n1881,
         n1880, n1879, n1878, n1877, n1876, n1875, n1874, n1873, n1872, n1871,
         n1870, n1869, n1868, n1867, n1866, n1865, n1864, n1863, n1862, n1861,
         n1860, n1859, n1858, n1857, n1856, n1855, n1854, n1853, n1852, n1851,
         n1850, n1849, n1848, n1847, n1846, n1845, n1844, n1843, n1842, n1841,
         n1840, n1839, n1838, n1837, n1836, n1835, n1834, n1833, n1832, n1831,
         n1830, n1829, n1828, n1827, n1826, n1825, n1824, n1823, n1822, n1821,
         n1820, n1819, n1818, n1817, n1816, n1815, n1814, n1813, n1812, n1811,
         n1810, n1809, n1808, n1807, n1806, n1805, n1804, n1803, n1802, n1801,
         n1800, n1799, n1798, n1797, n1796, n1795, n1794, n1793, n1792, n1791,
         n1790, n1789, n1788, n1787, n1786, n1785, n1784, n1783, n1782, n1781,
         n1780, n1779, n1778, n1777, n1776, n1775, n1774, n1773, n1772, n1771,
         n1770, n1769, n1768, n1767, n1766, n1765, n1764, n1763, n1762, n1761,
         n1760, n1759, n1758, n1757, n1756, n1755, n1754, n1753, n1752, n1751,
         n1750, n1749, n1748, n1747, n1746, n1745, n1744, n1743, n1742, n1741,
         n1740, n1739, n1738, n1737, n1736, n1735, n1734, n1733, n1732, n1731,
         n1730, n1729, n1728, n1727, n1726, n1725, n1724, n1723, n1722, n1721,
         n1720, n1719, n1718, n1717, n1716, n1715, n1714, n1713, n1712, n1711,
         n1710, n1709, n1708, n1707, n1706, n1705, n1704, n1703, n1702, n1701,
         n1700, n1699, n1698, n1697, n1696, n1695, n1694, n1693, n1692, n1691,
         n1690, n1689, n1688, n1687, n1686, n1685, n1684, n1683, n1682, n1681,
         n1680, n1679, n1678, n1677, n1676, n1675, n1674, n1673, n1672, n1671,
         n1670, n1669, n1668, n1667, n1666, n1665, n1664, n1663, n1662, n1661,
         n1660, n1659, n1658, n1657, n1656, n1655, n1654, n1653, n1652, n1651,
         n1650, n1649, n1648, n1647, n1646, n1645, n1644, n1643, n1642, n1641,
         n1640, n1639, n1638, n1637, n1636, n1635, n1634, n1633, n1632, n1631,
         n1630, n1629, n1628, n1627, n1626, n1625, n1624, n1623, n1622, n1621,
         n1620, n1619, n1618, n1617, n1616, n1615, n1614, n1613, n1612, n1611,
         n1610, n1609, n1608, n1607, n1606, n1605, n1604, n1603, n1602, n1601,
         n1600, n1599, n1598, n1597, n1596, n1595, n1594, n1593, n1592, n1591,
         n1590, n1589, n1588, n1587, n1586, n1585, n1584, n1583, n1582, n1581,
         n1580, n1579, n1578, n1577, n1576, n1575, n1574, n1573, n1572, n1571,
         n1570, n1569, n1568, n1567, n1566, n1565, n1564, n1563, n1562, n1561,
         n1560, n1559, n1558, n1557, n1556, n1555, n1554, n1553, n1552, n1551,
         n1550, n1549, n1548, n1547, n1546, n1545, n1544, n1543, n1542, n1541,
         n1540, n1539, n1538, n1537, n1536, n1534, n1533, n1532, n1531, n1530,
         n1529, n1528, n1527, n1526, n1525, n1524, n1523, n1522, n1521, n1520,
         n1519, n1518, n1517, n1516, n1515, n1514, n1513, n1512, n1511, n1510,
         n1509, n1508, n1507, n1506, n1505, n1504, n1503, n1502, n1501, n1500,
         n1499, n1498, n1497, n1496, n1495, n1494, n1493, n1492, n1491, n1490,
         n1489, n1488, n1487, n1486, n1485, n1484, n1482, n1481, n1480, n1479,
         n1478, n1477, n1476, n1475, n1474, n1473, n1471, n1470, n1469, n1468,
         n1467, n1466, n1465, n1464, n1463, n1462, n1460, n1459, n1458, n1456,
         n1455, n1454, n1452, n1451, n1450, n1449, n1448, n1446, n1445, n1444,
         n1443, n1442, n1441, n1440, n1439, n1438, n1437, n1436, n1435, n1434,
         n1433, n1432, n1431, n1430, n1429, n1428, n1427, n1426, n1425, n1424,
         n1423, n1422, n1421, n1420, n1419, n1418, n1417, n1416, n1415, n1414,
         n1413, n1412, n1411, n1410, n1409, n1408, n1407, n1406, n1405, n1404,
         n1403, n1402, n1401, n1400, n1399, n1398, n1397, n1396, n1395, n1394,
         n1393, n1392, n1391, n1390, n1389, n1388, n1387, n1386, n1385, n1384,
         n1383, n1382, n1381, n1380, n1379, n1378, n1377, n1376, n1375, n1374,
         n1373, n1372, n1371, n1370, n1369, n1368, n1367, n1366, n1365, n1364,
         n1363, n1362, n1361, n1360, n1359, n1358, n1357, n1356, n1355, n1354,
         n1353, n1352, n1351, n1350, n1349, n1348, n1347, n1346, n1345, n1344,
         n1343, n1342, n1341, n1340, n1339, n1338, n1337, n1336, n1335, n1334,
         n1333, n1332, n1331, n1330, n1329, n1328, n1327, n1326, n1325, n1324,
         n1323, n1322, n1321, n1320, n1319, n1318, n1317, n1316, n1315, n1314,
         n1313, n1312, n1311, n1310, n1309, n1308, n1307, n1306, n1305, n1304,
         n1303, n1302, n1301, n1300, n1299, n1298, n1297, n1296, n1295, n1294,
         n1293, n1292, n1291, n1290, n1289, n1288, n1287, n1286, n1285, n1284,
         n1283, n1282, n1281, n1280, n1279, n1278, n1277, n1276, n1275, n1274,
         n1273, n1272, n1271, n1270, n1269, n1268, n1267, n1266, n1265, n1264,
         n1263, n1262, n1261, n1260, n1259, n1258, n1257, n1256, n1255, n1254,
         n1253, n1252, n1251, n1250, n1249, n1248, n1247, n1246, n1245, n1244,
         n1243, n1242, n1241, n1240, n1239, n1238, n1237, n1236, n1235, n1234,
         n1233, n1232, n1231, n1230, n1229, n1228, n1227, n1226, n1225, n1224,
         n1223, n1222, n1221, n1220, n1219, n1218, n1217, n1216, n1215, n1214,
         n1213, n1212, n1211, n1210, n1209, n1208, n1207, n1206, n1205, n1204,
         n1203, n1202, n1201, n1200, n1199, n1198, n1197, n1196, n1195, n1194,
         n1193, n1192, n1191, n1190, n1189, n1188, n1187, n1186, n1185, n1184,
         n1183, n1182, n1181, n1180, n1179, n1178, n1177, n1176, n1175, n1174,
         n1173, n1172, n1171, n1170, n1169, n1168, n1167, n1166, n1165, n1164,
         n1163, n1162, n1161, n1160, n1159, n1158, n1157, n1156, n1155, n1154,
         n1153, n1152, n1151, n1150, n1149, n1148, n1147, n1146, n1145, n1144,
         n1143, n1142, n1141, n1140, n1139, n1138, n1137, n1136, n1135, n1134,
         n1133, n1132, n1131, n1130, n1129, n1128, n1127, n1126, n1125, n1124,
         n1123, n1122, n1121, n1120, n1119, n1118, n1117, n1116, n1115, n1114,
         n1113, n1112, n1111, n1110, n1109, n1108, n1107, n1106, n1105, n1104,
         n1103, n1102, n1101, n1100, n1099, n1098, n1097, n1096, n1095, n1094,
         n1093, n1092, n1091, n1090, n1089, n1088, n1087, n1086, n1085, n1084,
         n1083, n1082, n1081, n1080, n1079, n1078, n1077, n1076, n1075, n1074,
         n1073, n1072, n1071, n1070, n1069, n1068, n1067, n1066, n1065, n1064,
         n1063, n1062, n1061, n1060, n1059, n1058, n1057, n1056, n1055, n1054,
         n1053, n1052, n1051, n1050, n1049, n1048, n1047, n1046, n1045, n1044,
         n1043, n1042, n1041, n1040, n1039, n1038, n1037, n1036, n1035, n1034,
         n1033, n1032, n1031, n1030, n1029, n1028, n1027, n1026, n1025, n1024,
         n1023, n1022, n1021, n1020, n1019, n1018, n1017, n1016, n1015, n1014,
         n1013, n1012, n1011, n1010, n1009, n1008, n1007, n1006, n1005, n1004,
         n1003, n1002, n1001, n1000, n5912, n5913, n5914, n5915, n5916, n5917,
         n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927,
         n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937,
         n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947,
         n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957,
         n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967,
         n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977,
         n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987,
         n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997,
         n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007,
         n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017,
         n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027,
         n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037,
         n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047,
         n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057,
         n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067,
         n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077,
         n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087,
         n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097,
         n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107,
         n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117,
         n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127,
         n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137,
         n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147,
         n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157,
         n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167,
         n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177,
         n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187,
         n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197,
         n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207,
         n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217,
         n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227,
         n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237,
         n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247,
         n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257,
         n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267,
         n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277,
         n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287,
         n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297,
         n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307,
         n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317,
         n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327,
         n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337,
         n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347,
         n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357,
         n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367,
         n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377,
         n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387,
         n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397,
         n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407,
         n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417,
         n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427,
         n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437,
         n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447,
         n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457,
         n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467,
         n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477,
         n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487,
         n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497,
         n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507,
         n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517,
         n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527,
         n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537,
         n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547,
         n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557,
         n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567,
         n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577,
         n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587,
         n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597,
         n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607,
         n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617,
         n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627,
         n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637,
         n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647,
         n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657,
         n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667,
         n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677,
         n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687,
         n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697,
         n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707,
         n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717,
         n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727,
         n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737,
         n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747,
         n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757,
         n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767,
         n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777,
         n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787,
         n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797,
         n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807,
         n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817,
         n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827,
         n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837,
         n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847,
         n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857,
         n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867,
         n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877,
         n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887,
         n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897,
         n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907,
         n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917,
         n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927,
         n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937,
         n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947,
         n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957,
         n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967,
         n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977,
         n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987,
         n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997,
         n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007,
         n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017,
         n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027,
         n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037,
         n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047,
         n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057,
         n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067,
         n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077,
         n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087,
         n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097,
         n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107,
         n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117,
         n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127,
         n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137,
         n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147,
         n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157,
         n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167,
         n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177,
         n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187,
         n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197,
         n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207,
         n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217,
         n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227,
         n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237,
         n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247,
         n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257,
         n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267,
         n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277,
         n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287,
         n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297,
         n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307,
         n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317,
         n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327,
         n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337,
         n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347,
         n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357,
         n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367,
         n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377,
         n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387,
         n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397,
         n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407,
         n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417,
         n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427,
         n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437,
         n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447,
         n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457,
         n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467,
         n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477,
         n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903,
         n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913,
         n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923,
         n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933,
         n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943,
         n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953,
         n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963,
         n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973,
         n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983,
         n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993,
         n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003,
         n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013,
         n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023,
         n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033,
         n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043,
         n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053,
         n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063,
         n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073,
         n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083,
         n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093,
         n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103,
         n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113,
         n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123,
         n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133,
         n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143,
         n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153,
         n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163,
         n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173,
         n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183,
         n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193,
         n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203,
         n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213,
         n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223,
         n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233,
         n9234, n9235, n9236, n9237, n9238, n9239;

  dff_sg \state_reg[0]  ( .D(n20), .CP(clk), .Q(state[0]) );
  dff_sg \state_reg[1]  ( .D(n19), .CP(clk), .Q(state[1]) );
  dff_sg \update_mask_0/o_pointer_reg[3]  ( .D(\update_mask_0/n1083 ), .CP(clk), .Q(\update_mask_0/N31 ) );
  dff_sg \update_mask_0/o_pointer_reg[2]  ( .D(\update_mask_0/n1081 ), .CP(clk), .Q(\update_mask_0/N30 ) );
  dff_sg \update_mask_0/o_pointer_reg[1]  ( .D(n5911), .CP(clk), .Q(
        \update_mask_0/N29 ) );
  dff_sg \update_mask_0/o_pointer_reg[0]  ( .D(\update_mask_0/n1082 ), .CP(clk), .Q(\update_mask_0/N28 ) );
  dff_sg \update_mask_0/m_pointer_reg[3]  ( .D(\update_mask_0/n1084 ), .CP(clk), .Q(\update_mask_0/N26 ) );
  dff_sg \update_mask_0/m_pointer_reg[2]  ( .D(\update_mask_0/n1085 ), .CP(clk), .Q(\update_mask_0/N25 ) );
  dff_sg \update_mask_0/m_pointer_reg[1]  ( .D(\update_mask_0/n1086 ), .CP(clk), .Q(\update_mask_0/N24 ) );
  dff_sg \update_mask_0/m_pointer_reg[4]  ( .D(\update_mask_0/n1441 ), .CP(clk), .Q(\update_mask_0/N27 ) );
  dff_sg \update_mask_0/reg_i_mask_reg[0]  ( .D(\update_mask_0/n1438 ), .CP(
        clk), .Q(\update_mask_0/reg_i_mask[0] ) );
  dff_sg \update_mask_0/reg_i_mask_reg[1]  ( .D(\update_mask_0/n1437 ), .CP(
        clk), .Q(\update_mask_0/reg_i_mask[1] ) );
  dff_sg \update_mask_0/reg_i_mask_reg[2]  ( .D(\update_mask_0/n1436 ), .CP(
        clk), .Q(\update_mask_0/reg_i_mask[2] ) );
  dff_sg \update_mask_0/reg_i_mask_reg[3]  ( .D(\update_mask_0/n1435 ), .CP(
        clk), .Q(\update_mask_0/reg_i_mask[3] ) );
  dff_sg \update_mask_0/reg_i_mask_reg[4]  ( .D(\update_mask_0/n1434 ), .CP(
        clk), .Q(\update_mask_0/reg_i_mask[4] ) );
  dff_sg \update_mask_0/reg_i_mask_reg[5]  ( .D(\update_mask_0/n1433 ), .CP(
        clk), .Q(\update_mask_0/reg_i_mask[5] ) );
  dff_sg \update_mask_0/reg_i_mask_reg[6]  ( .D(\update_mask_0/n1432 ), .CP(
        clk), .Q(\update_mask_0/reg_i_mask[6] ) );
  dff_sg \update_mask_0/reg_i_mask_reg[7]  ( .D(\update_mask_0/n1431 ), .CP(
        clk), .Q(\update_mask_0/reg_i_mask[7] ) );
  dff_sg \update_mask_0/reg_i_mask_reg[8]  ( .D(\update_mask_0/n1430 ), .CP(
        clk), .Q(\update_mask_0/reg_i_mask[8] ) );
  dff_sg \update_mask_0/reg_i_mask_reg[9]  ( .D(\update_mask_0/n1429 ), .CP(
        clk), .Q(\update_mask_0/reg_i_mask[9] ) );
  dff_sg \update_mask_0/reg_i_mask_reg[10]  ( .D(\update_mask_0/n1428 ), .CP(
        clk), .Q(\update_mask_0/reg_i_mask[10] ) );
  dff_sg \update_mask_0/reg_i_mask_reg[11]  ( .D(\update_mask_0/n1427 ), .CP(
        clk), .Q(\update_mask_0/reg_i_mask[11] ) );
  dff_sg \update_mask_0/reg_i_mask_reg[12]  ( .D(\update_mask_0/n1426 ), .CP(
        clk), .Q(\update_mask_0/reg_i_mask[12] ) );
  dff_sg \update_mask_0/reg_i_mask_reg[13]  ( .D(\update_mask_0/n1425 ), .CP(
        clk), .Q(\update_mask_0/reg_i_mask[13] ) );
  dff_sg \update_mask_0/reg_i_mask_reg[14]  ( .D(\update_mask_0/n1424 ), .CP(
        clk), .Q(\update_mask_0/reg_i_mask[14] ) );
  dff_sg \update_mask_0/reg_i_mask_reg[15]  ( .D(\update_mask_0/n1423 ), .CP(
        clk), .Q(\update_mask_0/reg_i_mask[15] ) );
  dff_sg \update_mask_0/reg_i_mask_reg[16]  ( .D(\update_mask_0/n1422 ), .CP(
        clk), .Q(\update_mask_0/reg_i_mask[16] ) );
  dff_sg \update_mask_0/reg_i_mask_reg[17]  ( .D(\update_mask_0/n1421 ), .CP(
        clk), .Q(\update_mask_0/reg_i_mask[17] ) );
  dff_sg \update_mask_0/reg_i_mask_reg[18]  ( .D(\update_mask_0/n1420 ), .CP(
        clk), .Q(\update_mask_0/reg_i_mask[18] ) );
  dff_sg \update_mask_0/reg_i_mask_reg[19]  ( .D(\update_mask_0/n1419 ), .CP(
        clk), .Q(\update_mask_0/reg_i_mask[19] ) );
  dff_sg \update_mask_0/reg_i_mask_reg[20]  ( .D(\update_mask_0/n1418 ), .CP(
        clk), .Q(\update_mask_0/reg_i_mask[20] ) );
  dff_sg \update_mask_0/reg_i_mask_reg[21]  ( .D(\update_mask_0/n1417 ), .CP(
        clk), .Q(\update_mask_0/reg_i_mask[21] ) );
  dff_sg \update_mask_0/reg_i_mask_reg[22]  ( .D(\update_mask_0/n1416 ), .CP(
        clk), .Q(\update_mask_0/reg_i_mask[22] ) );
  dff_sg \update_mask_0/reg_i_mask_reg[23]  ( .D(\update_mask_0/n1415 ), .CP(
        clk), .Q(\update_mask_0/reg_i_mask[23] ) );
  dff_sg \update_mask_0/reg_i_mask_reg[24]  ( .D(\update_mask_0/n1414 ), .CP(
        clk), .Q(\update_mask_0/reg_i_mask[24] ) );
  dff_sg \update_mask_0/reg_i_mask_reg[25]  ( .D(\update_mask_0/n1413 ), .CP(
        clk), .Q(\update_mask_0/reg_i_mask[25] ) );
  dff_sg \update_mask_0/reg_i_mask_reg[26]  ( .D(\update_mask_0/n1412 ), .CP(
        clk), .Q(\update_mask_0/reg_i_mask[26] ) );
  dff_sg \update_mask_0/reg_i_mask_reg[27]  ( .D(\update_mask_0/n1411 ), .CP(
        clk), .Q(\update_mask_0/reg_i_mask[27] ) );
  dff_sg \update_mask_0/reg_i_mask_reg[28]  ( .D(\update_mask_0/n1410 ), .CP(
        clk), .Q(\update_mask_0/reg_i_mask[28] ) );
  dff_sg \update_mask_0/reg_i_mask_reg[29]  ( .D(\update_mask_0/n1409 ), .CP(
        clk), .Q(\update_mask_0/reg_i_mask[29] ) );
  dff_sg \update_mask_0/reg_i_mask_reg[30]  ( .D(\update_mask_0/n1408 ), .CP(
        clk), .Q(\update_mask_0/reg_i_mask[30] ) );
  dff_sg \update_mask_0/reg_i_mask_reg[31]  ( .D(\update_mask_0/n1407 ), .CP(
        clk), .Q(\update_mask_0/reg_i_mask[31] ) );
  dff_sg \update_mask_0/reg_out_reg[0][0]  ( .D(\update_mask_0/n1406 ), .CP(
        clk), .Q(\update_mask_0/reg_out[0][0] ) );
  dff_sg \update_mask_0/reg_out_reg[0][1]  ( .D(\update_mask_0/n1405 ), .CP(
        clk), .Q(\update_mask_0/reg_out[0][1] ) );
  dff_sg \update_mask_0/reg_out_reg[0][2]  ( .D(\update_mask_0/n1404 ), .CP(
        clk), .Q(\update_mask_0/reg_out[0][2] ) );
  dff_sg \update_mask_0/reg_out_reg[0][3]  ( .D(\update_mask_0/n1403 ), .CP(
        clk), .Q(\update_mask_0/reg_out[0][3] ) );
  dff_sg \update_mask_0/reg_out_reg[0][4]  ( .D(\update_mask_0/n1402 ), .CP(
        clk), .Q(\update_mask_0/reg_out[0][4] ) );
  dff_sg \update_mask_0/reg_out_reg[0][5]  ( .D(\update_mask_0/n1401 ), .CP(
        clk), .Q(\update_mask_0/reg_out[0][5] ) );
  dff_sg \update_mask_0/reg_out_reg[0][6]  ( .D(\update_mask_0/n1400 ), .CP(
        clk), .Q(\update_mask_0/reg_out[0][6] ) );
  dff_sg \update_mask_0/reg_out_reg[0][7]  ( .D(\update_mask_0/n1399 ), .CP(
        clk), .Q(\update_mask_0/reg_out[0][7] ) );
  dff_sg \update_mask_0/reg_out_reg[0][8]  ( .D(\update_mask_0/n1398 ), .CP(
        clk), .Q(\update_mask_0/reg_out[0][8] ) );
  dff_sg \update_mask_0/reg_out_reg[0][9]  ( .D(\update_mask_0/n1397 ), .CP(
        clk), .Q(\update_mask_0/reg_out[0][9] ) );
  dff_sg \update_mask_0/reg_out_reg[0][10]  ( .D(\update_mask_0/n1396 ), .CP(
        clk), .Q(\update_mask_0/reg_out[0][10] ) );
  dff_sg \update_mask_0/reg_out_reg[0][11]  ( .D(\update_mask_0/n1395 ), .CP(
        clk), .Q(\update_mask_0/reg_out[0][11] ) );
  dff_sg \update_mask_0/reg_out_reg[0][12]  ( .D(\update_mask_0/n1394 ), .CP(
        clk), .Q(\update_mask_0/reg_out[0][12] ) );
  dff_sg \update_mask_0/reg_out_reg[0][13]  ( .D(\update_mask_0/n1393 ), .CP(
        clk), .Q(\update_mask_0/reg_out[0][13] ) );
  dff_sg \update_mask_0/reg_out_reg[0][14]  ( .D(\update_mask_0/n1392 ), .CP(
        clk), .Q(\update_mask_0/reg_out[0][14] ) );
  dff_sg \update_mask_0/reg_out_reg[0][15]  ( .D(\update_mask_0/n1391 ), .CP(
        clk), .Q(\update_mask_0/reg_out[0][15] ) );
  dff_sg \update_mask_0/reg_out_reg[0][16]  ( .D(\update_mask_0/n1390 ), .CP(
        clk), .Q(\update_mask_0/reg_out[0][16] ) );
  dff_sg \update_mask_0/reg_out_reg[0][17]  ( .D(\update_mask_0/n1389 ), .CP(
        clk), .Q(\update_mask_0/reg_out[0][17] ) );
  dff_sg \update_mask_0/reg_out_reg[0][18]  ( .D(\update_mask_0/n1388 ), .CP(
        clk), .Q(\update_mask_0/reg_out[0][18] ) );
  dff_sg \update_mask_0/reg_out_reg[0][19]  ( .D(\update_mask_0/n1387 ), .CP(
        clk), .Q(\update_mask_0/reg_out[0][19] ) );
  dff_sg \update_mask_0/reg_out_reg[1][0]  ( .D(\update_mask_0/n1386 ), .CP(
        clk), .Q(\update_mask_0/reg_out[1][0] ) );
  dff_sg \update_mask_0/reg_out_reg[1][1]  ( .D(\update_mask_0/n1385 ), .CP(
        clk), .Q(\update_mask_0/reg_out[1][1] ) );
  dff_sg \update_mask_0/reg_out_reg[1][2]  ( .D(\update_mask_0/n1384 ), .CP(
        clk), .Q(\update_mask_0/reg_out[1][2] ) );
  dff_sg \update_mask_0/reg_out_reg[1][3]  ( .D(\update_mask_0/n1383 ), .CP(
        clk), .Q(\update_mask_0/reg_out[1][3] ) );
  dff_sg \update_mask_0/reg_out_reg[1][4]  ( .D(\update_mask_0/n1382 ), .CP(
        clk), .Q(\update_mask_0/reg_out[1][4] ) );
  dff_sg \update_mask_0/reg_out_reg[1][5]  ( .D(\update_mask_0/n1381 ), .CP(
        clk), .Q(\update_mask_0/reg_out[1][5] ) );
  dff_sg \update_mask_0/reg_out_reg[1][6]  ( .D(\update_mask_0/n1380 ), .CP(
        clk), .Q(\update_mask_0/reg_out[1][6] ) );
  dff_sg \update_mask_0/reg_out_reg[1][7]  ( .D(\update_mask_0/n1379 ), .CP(
        clk), .Q(\update_mask_0/reg_out[1][7] ) );
  dff_sg \update_mask_0/reg_out_reg[1][8]  ( .D(\update_mask_0/n1378 ), .CP(
        clk), .Q(\update_mask_0/reg_out[1][8] ) );
  dff_sg \update_mask_0/reg_out_reg[1][9]  ( .D(\update_mask_0/n1377 ), .CP(
        clk), .Q(\update_mask_0/reg_out[1][9] ) );
  dff_sg \update_mask_0/reg_out_reg[1][10]  ( .D(\update_mask_0/n1376 ), .CP(
        clk), .Q(\update_mask_0/reg_out[1][10] ) );
  dff_sg \update_mask_0/reg_out_reg[1][11]  ( .D(\update_mask_0/n1375 ), .CP(
        clk), .Q(\update_mask_0/reg_out[1][11] ) );
  dff_sg \update_mask_0/reg_out_reg[1][12]  ( .D(\update_mask_0/n1374 ), .CP(
        clk), .Q(\update_mask_0/reg_out[1][12] ) );
  dff_sg \update_mask_0/reg_out_reg[1][13]  ( .D(\update_mask_0/n1373 ), .CP(
        clk), .Q(\update_mask_0/reg_out[1][13] ) );
  dff_sg \update_mask_0/reg_out_reg[1][14]  ( .D(\update_mask_0/n1372 ), .CP(
        clk), .Q(\update_mask_0/reg_out[1][14] ) );
  dff_sg \update_mask_0/reg_out_reg[1][15]  ( .D(\update_mask_0/n1371 ), .CP(
        clk), .Q(\update_mask_0/reg_out[1][15] ) );
  dff_sg \update_mask_0/reg_out_reg[1][16]  ( .D(\update_mask_0/n1370 ), .CP(
        clk), .Q(\update_mask_0/reg_out[1][16] ) );
  dff_sg \update_mask_0/reg_out_reg[1][17]  ( .D(\update_mask_0/n1369 ), .CP(
        clk), .Q(\update_mask_0/reg_out[1][17] ) );
  dff_sg \update_mask_0/reg_out_reg[1][18]  ( .D(\update_mask_0/n1368 ), .CP(
        clk), .Q(\update_mask_0/reg_out[1][18] ) );
  dff_sg \update_mask_0/reg_out_reg[1][19]  ( .D(\update_mask_0/n1367 ), .CP(
        clk), .Q(\update_mask_0/reg_out[1][19] ) );
  dff_sg \update_mask_0/reg_out_reg[2][0]  ( .D(\update_mask_0/n1366 ), .CP(
        clk), .Q(\update_mask_0/reg_out[2][0] ) );
  dff_sg \update_mask_0/reg_out_reg[2][1]  ( .D(\update_mask_0/n1365 ), .CP(
        clk), .Q(\update_mask_0/reg_out[2][1] ) );
  dff_sg \update_mask_0/reg_out_reg[2][2]  ( .D(\update_mask_0/n1364 ), .CP(
        clk), .Q(\update_mask_0/reg_out[2][2] ) );
  dff_sg \update_mask_0/reg_out_reg[2][3]  ( .D(\update_mask_0/n1363 ), .CP(
        clk), .Q(\update_mask_0/reg_out[2][3] ) );
  dff_sg \update_mask_0/reg_out_reg[2][4]  ( .D(\update_mask_0/n1362 ), .CP(
        clk), .Q(\update_mask_0/reg_out[2][4] ) );
  dff_sg \update_mask_0/reg_out_reg[2][5]  ( .D(\update_mask_0/n1361 ), .CP(
        clk), .Q(\update_mask_0/reg_out[2][5] ) );
  dff_sg \update_mask_0/reg_out_reg[2][6]  ( .D(\update_mask_0/n1360 ), .CP(
        clk), .Q(\update_mask_0/reg_out[2][6] ) );
  dff_sg \update_mask_0/reg_out_reg[2][7]  ( .D(\update_mask_0/n1359 ), .CP(
        clk), .Q(\update_mask_0/reg_out[2][7] ) );
  dff_sg \update_mask_0/reg_out_reg[2][8]  ( .D(\update_mask_0/n1358 ), .CP(
        clk), .Q(\update_mask_0/reg_out[2][8] ) );
  dff_sg \update_mask_0/reg_out_reg[2][9]  ( .D(\update_mask_0/n1357 ), .CP(
        clk), .Q(\update_mask_0/reg_out[2][9] ) );
  dff_sg \update_mask_0/reg_out_reg[2][10]  ( .D(\update_mask_0/n1356 ), .CP(
        clk), .Q(\update_mask_0/reg_out[2][10] ) );
  dff_sg \update_mask_0/reg_out_reg[2][11]  ( .D(\update_mask_0/n1355 ), .CP(
        clk), .Q(\update_mask_0/reg_out[2][11] ) );
  dff_sg \update_mask_0/reg_out_reg[2][12]  ( .D(\update_mask_0/n1354 ), .CP(
        clk), .Q(\update_mask_0/reg_out[2][12] ) );
  dff_sg \update_mask_0/reg_out_reg[2][13]  ( .D(\update_mask_0/n1353 ), .CP(
        clk), .Q(\update_mask_0/reg_out[2][13] ) );
  dff_sg \update_mask_0/reg_out_reg[2][14]  ( .D(\update_mask_0/n1352 ), .CP(
        clk), .Q(\update_mask_0/reg_out[2][14] ) );
  dff_sg \update_mask_0/reg_out_reg[2][15]  ( .D(\update_mask_0/n1351 ), .CP(
        clk), .Q(\update_mask_0/reg_out[2][15] ) );
  dff_sg \update_mask_0/reg_out_reg[2][16]  ( .D(\update_mask_0/n1350 ), .CP(
        clk), .Q(\update_mask_0/reg_out[2][16] ) );
  dff_sg \update_mask_0/reg_out_reg[2][17]  ( .D(\update_mask_0/n1349 ), .CP(
        clk), .Q(\update_mask_0/reg_out[2][17] ) );
  dff_sg \update_mask_0/reg_out_reg[2][18]  ( .D(\update_mask_0/n1348 ), .CP(
        clk), .Q(\update_mask_0/reg_out[2][18] ) );
  dff_sg \update_mask_0/reg_out_reg[2][19]  ( .D(\update_mask_0/n1347 ), .CP(
        clk), .Q(\update_mask_0/reg_out[2][19] ) );
  dff_sg \update_mask_0/reg_out_reg[3][0]  ( .D(\update_mask_0/n1346 ), .CP(
        clk), .Q(\update_mask_0/reg_out[3][0] ) );
  dff_sg \update_mask_0/reg_out_reg[3][1]  ( .D(\update_mask_0/n1345 ), .CP(
        clk), .Q(\update_mask_0/reg_out[3][1] ) );
  dff_sg \update_mask_0/reg_out_reg[3][2]  ( .D(\update_mask_0/n1344 ), .CP(
        clk), .Q(\update_mask_0/reg_out[3][2] ) );
  dff_sg \update_mask_0/reg_out_reg[3][3]  ( .D(\update_mask_0/n1343 ), .CP(
        clk), .Q(\update_mask_0/reg_out[3][3] ) );
  dff_sg \update_mask_0/reg_out_reg[3][4]  ( .D(\update_mask_0/n1342 ), .CP(
        clk), .Q(\update_mask_0/reg_out[3][4] ) );
  dff_sg \update_mask_0/reg_out_reg[3][5]  ( .D(\update_mask_0/n1341 ), .CP(
        clk), .Q(\update_mask_0/reg_out[3][5] ) );
  dff_sg \update_mask_0/reg_out_reg[3][6]  ( .D(\update_mask_0/n1340 ), .CP(
        clk), .Q(\update_mask_0/reg_out[3][6] ) );
  dff_sg \update_mask_0/reg_out_reg[3][7]  ( .D(\update_mask_0/n1339 ), .CP(
        clk), .Q(\update_mask_0/reg_out[3][7] ) );
  dff_sg \update_mask_0/reg_out_reg[3][8]  ( .D(\update_mask_0/n1338 ), .CP(
        clk), .Q(\update_mask_0/reg_out[3][8] ) );
  dff_sg \update_mask_0/reg_out_reg[3][9]  ( .D(\update_mask_0/n1337 ), .CP(
        clk), .Q(\update_mask_0/reg_out[3][9] ) );
  dff_sg \update_mask_0/reg_out_reg[3][10]  ( .D(\update_mask_0/n1336 ), .CP(
        clk), .Q(\update_mask_0/reg_out[3][10] ) );
  dff_sg \update_mask_0/reg_out_reg[3][11]  ( .D(\update_mask_0/n1335 ), .CP(
        clk), .Q(\update_mask_0/reg_out[3][11] ) );
  dff_sg \update_mask_0/reg_out_reg[3][12]  ( .D(\update_mask_0/n1334 ), .CP(
        clk), .Q(\update_mask_0/reg_out[3][12] ) );
  dff_sg \update_mask_0/reg_out_reg[3][13]  ( .D(\update_mask_0/n1333 ), .CP(
        clk), .Q(\update_mask_0/reg_out[3][13] ) );
  dff_sg \update_mask_0/reg_out_reg[3][14]  ( .D(\update_mask_0/n1332 ), .CP(
        clk), .Q(\update_mask_0/reg_out[3][14] ) );
  dff_sg \update_mask_0/reg_out_reg[3][15]  ( .D(\update_mask_0/n1331 ), .CP(
        clk), .Q(\update_mask_0/reg_out[3][15] ) );
  dff_sg \update_mask_0/reg_out_reg[3][16]  ( .D(\update_mask_0/n1330 ), .CP(
        clk), .Q(\update_mask_0/reg_out[3][16] ) );
  dff_sg \update_mask_0/reg_out_reg[3][17]  ( .D(\update_mask_0/n1329 ), .CP(
        clk), .Q(\update_mask_0/reg_out[3][17] ) );
  dff_sg \update_mask_0/reg_out_reg[3][18]  ( .D(\update_mask_0/n1328 ), .CP(
        clk), .Q(\update_mask_0/reg_out[3][18] ) );
  dff_sg \update_mask_0/reg_out_reg[3][19]  ( .D(\update_mask_0/n1327 ), .CP(
        clk), .Q(\update_mask_0/reg_out[3][19] ) );
  dff_sg \update_mask_0/reg_out_reg[4][0]  ( .D(\update_mask_0/n1326 ), .CP(
        clk), .Q(\update_mask_0/reg_out[4][0] ) );
  dff_sg \update_mask_0/reg_out_reg[4][1]  ( .D(\update_mask_0/n1325 ), .CP(
        clk), .Q(\update_mask_0/reg_out[4][1] ) );
  dff_sg \update_mask_0/reg_out_reg[4][2]  ( .D(\update_mask_0/n1324 ), .CP(
        clk), .Q(\update_mask_0/reg_out[4][2] ) );
  dff_sg \update_mask_0/reg_out_reg[4][3]  ( .D(\update_mask_0/n1323 ), .CP(
        clk), .Q(\update_mask_0/reg_out[4][3] ) );
  dff_sg \update_mask_0/reg_out_reg[4][4]  ( .D(\update_mask_0/n1322 ), .CP(
        clk), .Q(\update_mask_0/reg_out[4][4] ) );
  dff_sg \update_mask_0/reg_out_reg[4][5]  ( .D(\update_mask_0/n1321 ), .CP(
        clk), .Q(\update_mask_0/reg_out[4][5] ) );
  dff_sg \update_mask_0/reg_out_reg[4][6]  ( .D(\update_mask_0/n1320 ), .CP(
        clk), .Q(\update_mask_0/reg_out[4][6] ) );
  dff_sg \update_mask_0/reg_out_reg[4][7]  ( .D(\update_mask_0/n1319 ), .CP(
        clk), .Q(\update_mask_0/reg_out[4][7] ) );
  dff_sg \update_mask_0/reg_out_reg[4][8]  ( .D(\update_mask_0/n1318 ), .CP(
        clk), .Q(\update_mask_0/reg_out[4][8] ) );
  dff_sg \update_mask_0/reg_out_reg[4][9]  ( .D(\update_mask_0/n1317 ), .CP(
        clk), .Q(\update_mask_0/reg_out[4][9] ) );
  dff_sg \update_mask_0/reg_out_reg[4][10]  ( .D(\update_mask_0/n1316 ), .CP(
        clk), .Q(\update_mask_0/reg_out[4][10] ) );
  dff_sg \update_mask_0/reg_out_reg[4][11]  ( .D(\update_mask_0/n1315 ), .CP(
        clk), .Q(\update_mask_0/reg_out[4][11] ) );
  dff_sg \update_mask_0/reg_out_reg[4][12]  ( .D(\update_mask_0/n1314 ), .CP(
        clk), .Q(\update_mask_0/reg_out[4][12] ) );
  dff_sg \update_mask_0/reg_out_reg[4][13]  ( .D(\update_mask_0/n1313 ), .CP(
        clk), .Q(\update_mask_0/reg_out[4][13] ) );
  dff_sg \update_mask_0/reg_out_reg[4][14]  ( .D(\update_mask_0/n1312 ), .CP(
        clk), .Q(\update_mask_0/reg_out[4][14] ) );
  dff_sg \update_mask_0/reg_out_reg[4][15]  ( .D(\update_mask_0/n1311 ), .CP(
        clk), .Q(\update_mask_0/reg_out[4][15] ) );
  dff_sg \update_mask_0/reg_out_reg[4][16]  ( .D(\update_mask_0/n1310 ), .CP(
        clk), .Q(\update_mask_0/reg_out[4][16] ) );
  dff_sg \update_mask_0/reg_out_reg[4][17]  ( .D(\update_mask_0/n1309 ), .CP(
        clk), .Q(\update_mask_0/reg_out[4][17] ) );
  dff_sg \update_mask_0/reg_out_reg[4][18]  ( .D(\update_mask_0/n1308 ), .CP(
        clk), .Q(\update_mask_0/reg_out[4][18] ) );
  dff_sg \update_mask_0/reg_out_reg[4][19]  ( .D(\update_mask_0/n1307 ), .CP(
        clk), .Q(\update_mask_0/reg_out[4][19] ) );
  dff_sg \update_mask_0/reg_out_reg[5][0]  ( .D(\update_mask_0/n1306 ), .CP(
        clk), .Q(\update_mask_0/reg_out[5][0] ) );
  dff_sg \update_mask_0/reg_out_reg[5][1]  ( .D(\update_mask_0/n1305 ), .CP(
        clk), .Q(\update_mask_0/reg_out[5][1] ) );
  dff_sg \update_mask_0/reg_out_reg[5][2]  ( .D(\update_mask_0/n1304 ), .CP(
        clk), .Q(\update_mask_0/reg_out[5][2] ) );
  dff_sg \update_mask_0/reg_out_reg[5][3]  ( .D(\update_mask_0/n1303 ), .CP(
        clk), .Q(\update_mask_0/reg_out[5][3] ) );
  dff_sg \update_mask_0/reg_out_reg[5][4]  ( .D(\update_mask_0/n1302 ), .CP(
        clk), .Q(\update_mask_0/reg_out[5][4] ) );
  dff_sg \update_mask_0/reg_out_reg[5][5]  ( .D(\update_mask_0/n1301 ), .CP(
        clk), .Q(\update_mask_0/reg_out[5][5] ) );
  dff_sg \update_mask_0/reg_out_reg[5][6]  ( .D(\update_mask_0/n1300 ), .CP(
        clk), .Q(\update_mask_0/reg_out[5][6] ) );
  dff_sg \update_mask_0/reg_out_reg[5][7]  ( .D(\update_mask_0/n1299 ), .CP(
        clk), .Q(\update_mask_0/reg_out[5][7] ) );
  dff_sg \update_mask_0/reg_out_reg[5][8]  ( .D(\update_mask_0/n1298 ), .CP(
        clk), .Q(\update_mask_0/reg_out[5][8] ) );
  dff_sg \update_mask_0/reg_out_reg[5][9]  ( .D(\update_mask_0/n1297 ), .CP(
        clk), .Q(\update_mask_0/reg_out[5][9] ) );
  dff_sg \update_mask_0/reg_out_reg[5][10]  ( .D(\update_mask_0/n1296 ), .CP(
        clk), .Q(\update_mask_0/reg_out[5][10] ) );
  dff_sg \update_mask_0/reg_out_reg[5][11]  ( .D(\update_mask_0/n1295 ), .CP(
        clk), .Q(\update_mask_0/reg_out[5][11] ) );
  dff_sg \update_mask_0/reg_out_reg[5][12]  ( .D(\update_mask_0/n1294 ), .CP(
        clk), .Q(\update_mask_0/reg_out[5][12] ) );
  dff_sg \update_mask_0/reg_out_reg[5][13]  ( .D(\update_mask_0/n1293 ), .CP(
        clk), .Q(\update_mask_0/reg_out[5][13] ) );
  dff_sg \update_mask_0/reg_out_reg[5][14]  ( .D(\update_mask_0/n1292 ), .CP(
        clk), .Q(\update_mask_0/reg_out[5][14] ) );
  dff_sg \update_mask_0/reg_out_reg[5][15]  ( .D(\update_mask_0/n1291 ), .CP(
        clk), .Q(\update_mask_0/reg_out[5][15] ) );
  dff_sg \update_mask_0/reg_out_reg[5][16]  ( .D(\update_mask_0/n1290 ), .CP(
        clk), .Q(\update_mask_0/reg_out[5][16] ) );
  dff_sg \update_mask_0/reg_out_reg[5][17]  ( .D(\update_mask_0/n1289 ), .CP(
        clk), .Q(\update_mask_0/reg_out[5][17] ) );
  dff_sg \update_mask_0/reg_out_reg[5][18]  ( .D(\update_mask_0/n1288 ), .CP(
        clk), .Q(\update_mask_0/reg_out[5][18] ) );
  dff_sg \update_mask_0/reg_out_reg[5][19]  ( .D(\update_mask_0/n1287 ), .CP(
        clk), .Q(\update_mask_0/reg_out[5][19] ) );
  dff_sg \update_mask_0/reg_out_reg[6][0]  ( .D(\update_mask_0/n1286 ), .CP(
        clk), .Q(\update_mask_0/reg_out[6][0] ) );
  dff_sg \update_mask_0/reg_out_reg[6][1]  ( .D(\update_mask_0/n1285 ), .CP(
        clk), .Q(\update_mask_0/reg_out[6][1] ) );
  dff_sg \update_mask_0/reg_out_reg[6][2]  ( .D(\update_mask_0/n1284 ), .CP(
        clk), .Q(\update_mask_0/reg_out[6][2] ) );
  dff_sg \update_mask_0/reg_out_reg[6][3]  ( .D(\update_mask_0/n1283 ), .CP(
        clk), .Q(\update_mask_0/reg_out[6][3] ) );
  dff_sg \update_mask_0/reg_out_reg[6][4]  ( .D(\update_mask_0/n1282 ), .CP(
        clk), .Q(\update_mask_0/reg_out[6][4] ) );
  dff_sg \update_mask_0/reg_out_reg[6][5]  ( .D(\update_mask_0/n1281 ), .CP(
        clk), .Q(\update_mask_0/reg_out[6][5] ) );
  dff_sg \update_mask_0/reg_out_reg[6][6]  ( .D(\update_mask_0/n1280 ), .CP(
        clk), .Q(\update_mask_0/reg_out[6][6] ) );
  dff_sg \update_mask_0/reg_out_reg[6][7]  ( .D(\update_mask_0/n1279 ), .CP(
        clk), .Q(\update_mask_0/reg_out[6][7] ) );
  dff_sg \update_mask_0/reg_out_reg[6][8]  ( .D(\update_mask_0/n1278 ), .CP(
        clk), .Q(\update_mask_0/reg_out[6][8] ) );
  dff_sg \update_mask_0/reg_out_reg[6][9]  ( .D(\update_mask_0/n1277 ), .CP(
        clk), .Q(\update_mask_0/reg_out[6][9] ) );
  dff_sg \update_mask_0/reg_out_reg[6][10]  ( .D(\update_mask_0/n1276 ), .CP(
        clk), .Q(\update_mask_0/reg_out[6][10] ) );
  dff_sg \update_mask_0/reg_out_reg[6][11]  ( .D(\update_mask_0/n1275 ), .CP(
        clk), .Q(\update_mask_0/reg_out[6][11] ) );
  dff_sg \update_mask_0/reg_out_reg[6][12]  ( .D(\update_mask_0/n1274 ), .CP(
        clk), .Q(\update_mask_0/reg_out[6][12] ) );
  dff_sg \update_mask_0/reg_out_reg[6][13]  ( .D(\update_mask_0/n1273 ), .CP(
        clk), .Q(\update_mask_0/reg_out[6][13] ) );
  dff_sg \update_mask_0/reg_out_reg[6][14]  ( .D(\update_mask_0/n1272 ), .CP(
        clk), .Q(\update_mask_0/reg_out[6][14] ) );
  dff_sg \update_mask_0/reg_out_reg[6][15]  ( .D(\update_mask_0/n1271 ), .CP(
        clk), .Q(\update_mask_0/reg_out[6][15] ) );
  dff_sg \update_mask_0/reg_out_reg[6][16]  ( .D(\update_mask_0/n1270 ), .CP(
        clk), .Q(\update_mask_0/reg_out[6][16] ) );
  dff_sg \update_mask_0/reg_out_reg[6][17]  ( .D(\update_mask_0/n1269 ), .CP(
        clk), .Q(\update_mask_0/reg_out[6][17] ) );
  dff_sg \update_mask_0/reg_out_reg[6][18]  ( .D(\update_mask_0/n1268 ), .CP(
        clk), .Q(\update_mask_0/reg_out[6][18] ) );
  dff_sg \update_mask_0/reg_out_reg[6][19]  ( .D(\update_mask_0/n1267 ), .CP(
        clk), .Q(\update_mask_0/reg_out[6][19] ) );
  dff_sg \update_mask_0/reg_out_reg[7][0]  ( .D(\update_mask_0/n1266 ), .CP(
        clk), .Q(\update_mask_0/reg_out[7][0] ) );
  dff_sg \update_mask_0/reg_out_reg[7][1]  ( .D(\update_mask_0/n1265 ), .CP(
        clk), .Q(\update_mask_0/reg_out[7][1] ) );
  dff_sg \update_mask_0/reg_out_reg[7][2]  ( .D(\update_mask_0/n1264 ), .CP(
        clk), .Q(\update_mask_0/reg_out[7][2] ) );
  dff_sg \update_mask_0/reg_out_reg[7][3]  ( .D(\update_mask_0/n1263 ), .CP(
        clk), .Q(\update_mask_0/reg_out[7][3] ) );
  dff_sg \update_mask_0/reg_out_reg[7][4]  ( .D(\update_mask_0/n1262 ), .CP(
        clk), .Q(\update_mask_0/reg_out[7][4] ) );
  dff_sg \update_mask_0/reg_out_reg[7][5]  ( .D(\update_mask_0/n1261 ), .CP(
        clk), .Q(\update_mask_0/reg_out[7][5] ) );
  dff_sg \update_mask_0/reg_out_reg[7][6]  ( .D(\update_mask_0/n1260 ), .CP(
        clk), .Q(\update_mask_0/reg_out[7][6] ) );
  dff_sg \update_mask_0/reg_out_reg[7][7]  ( .D(\update_mask_0/n1259 ), .CP(
        clk), .Q(\update_mask_0/reg_out[7][7] ) );
  dff_sg \update_mask_0/reg_out_reg[7][8]  ( .D(\update_mask_0/n1258 ), .CP(
        clk), .Q(\update_mask_0/reg_out[7][8] ) );
  dff_sg \update_mask_0/reg_out_reg[7][9]  ( .D(\update_mask_0/n1257 ), .CP(
        clk), .Q(\update_mask_0/reg_out[7][9] ) );
  dff_sg \update_mask_0/reg_out_reg[7][10]  ( .D(\update_mask_0/n1256 ), .CP(
        clk), .Q(\update_mask_0/reg_out[7][10] ) );
  dff_sg \update_mask_0/reg_out_reg[7][11]  ( .D(\update_mask_0/n1255 ), .CP(
        clk), .Q(\update_mask_0/reg_out[7][11] ) );
  dff_sg \update_mask_0/reg_out_reg[7][12]  ( .D(\update_mask_0/n1254 ), .CP(
        clk), .Q(\update_mask_0/reg_out[7][12] ) );
  dff_sg \update_mask_0/reg_out_reg[7][13]  ( .D(\update_mask_0/n1253 ), .CP(
        clk), .Q(\update_mask_0/reg_out[7][13] ) );
  dff_sg \update_mask_0/reg_out_reg[7][14]  ( .D(\update_mask_0/n1252 ), .CP(
        clk), .Q(\update_mask_0/reg_out[7][14] ) );
  dff_sg \update_mask_0/reg_out_reg[7][15]  ( .D(\update_mask_0/n1251 ), .CP(
        clk), .Q(\update_mask_0/reg_out[7][15] ) );
  dff_sg \update_mask_0/reg_out_reg[7][16]  ( .D(\update_mask_0/n1250 ), .CP(
        clk), .Q(\update_mask_0/reg_out[7][16] ) );
  dff_sg \update_mask_0/reg_out_reg[7][17]  ( .D(\update_mask_0/n1249 ), .CP(
        clk), .Q(\update_mask_0/reg_out[7][17] ) );
  dff_sg \update_mask_0/reg_out_reg[7][18]  ( .D(\update_mask_0/n1248 ), .CP(
        clk), .Q(\update_mask_0/reg_out[7][18] ) );
  dff_sg \update_mask_0/reg_out_reg[7][19]  ( .D(\update_mask_0/n1247 ), .CP(
        clk), .Q(\update_mask_0/reg_out[7][19] ) );
  dff_sg \update_mask_0/reg_out_reg[8][0]  ( .D(\update_mask_0/n1246 ), .CP(
        clk), .Q(\update_mask_0/reg_out[8][0] ) );
  dff_sg \update_mask_0/reg_out_reg[8][1]  ( .D(\update_mask_0/n1245 ), .CP(
        clk), .Q(\update_mask_0/reg_out[8][1] ) );
  dff_sg \update_mask_0/reg_out_reg[8][2]  ( .D(\update_mask_0/n1244 ), .CP(
        clk), .Q(\update_mask_0/reg_out[8][2] ) );
  dff_sg \update_mask_0/reg_out_reg[8][3]  ( .D(\update_mask_0/n1243 ), .CP(
        clk), .Q(\update_mask_0/reg_out[8][3] ) );
  dff_sg \update_mask_0/reg_out_reg[8][4]  ( .D(\update_mask_0/n1242 ), .CP(
        clk), .Q(\update_mask_0/reg_out[8][4] ) );
  dff_sg \update_mask_0/reg_out_reg[8][5]  ( .D(\update_mask_0/n1241 ), .CP(
        clk), .Q(\update_mask_0/reg_out[8][5] ) );
  dff_sg \update_mask_0/reg_out_reg[8][6]  ( .D(\update_mask_0/n1240 ), .CP(
        clk), .Q(\update_mask_0/reg_out[8][6] ) );
  dff_sg \update_mask_0/reg_out_reg[8][7]  ( .D(\update_mask_0/n1239 ), .CP(
        clk), .Q(\update_mask_0/reg_out[8][7] ) );
  dff_sg \update_mask_0/reg_out_reg[8][8]  ( .D(\update_mask_0/n1238 ), .CP(
        clk), .Q(\update_mask_0/reg_out[8][8] ) );
  dff_sg \update_mask_0/reg_out_reg[8][9]  ( .D(\update_mask_0/n1237 ), .CP(
        clk), .Q(\update_mask_0/reg_out[8][9] ) );
  dff_sg \update_mask_0/reg_out_reg[8][10]  ( .D(\update_mask_0/n1236 ), .CP(
        clk), .Q(\update_mask_0/reg_out[8][10] ) );
  dff_sg \update_mask_0/reg_out_reg[8][11]  ( .D(\update_mask_0/n1235 ), .CP(
        clk), .Q(\update_mask_0/reg_out[8][11] ) );
  dff_sg \update_mask_0/reg_out_reg[8][12]  ( .D(\update_mask_0/n1234 ), .CP(
        clk), .Q(\update_mask_0/reg_out[8][12] ) );
  dff_sg \update_mask_0/reg_out_reg[8][13]  ( .D(\update_mask_0/n1233 ), .CP(
        clk), .Q(\update_mask_0/reg_out[8][13] ) );
  dff_sg \update_mask_0/reg_out_reg[8][14]  ( .D(\update_mask_0/n1232 ), .CP(
        clk), .Q(\update_mask_0/reg_out[8][14] ) );
  dff_sg \update_mask_0/reg_out_reg[8][15]  ( .D(\update_mask_0/n1231 ), .CP(
        clk), .Q(\update_mask_0/reg_out[8][15] ) );
  dff_sg \update_mask_0/reg_out_reg[8][16]  ( .D(\update_mask_0/n1230 ), .CP(
        clk), .Q(\update_mask_0/reg_out[8][16] ) );
  dff_sg \update_mask_0/reg_out_reg[8][17]  ( .D(\update_mask_0/n1229 ), .CP(
        clk), .Q(\update_mask_0/reg_out[8][17] ) );
  dff_sg \update_mask_0/reg_out_reg[8][18]  ( .D(\update_mask_0/n1228 ), .CP(
        clk), .Q(\update_mask_0/reg_out[8][18] ) );
  dff_sg \update_mask_0/reg_out_reg[8][19]  ( .D(\update_mask_0/n1227 ), .CP(
        clk), .Q(\update_mask_0/reg_out[8][19] ) );
  dff_sg \update_mask_0/reg_out_reg[9][0]  ( .D(\update_mask_0/n1226 ), .CP(
        clk), .Q(\update_mask_0/reg_out[9][0] ) );
  dff_sg \update_mask_0/reg_out_reg[9][1]  ( .D(\update_mask_0/n1225 ), .CP(
        clk), .Q(\update_mask_0/reg_out[9][1] ) );
  dff_sg \update_mask_0/reg_out_reg[9][2]  ( .D(\update_mask_0/n1224 ), .CP(
        clk), .Q(\update_mask_0/reg_out[9][2] ) );
  dff_sg \update_mask_0/reg_out_reg[9][3]  ( .D(\update_mask_0/n1223 ), .CP(
        clk), .Q(\update_mask_0/reg_out[9][3] ) );
  dff_sg \update_mask_0/reg_out_reg[9][4]  ( .D(\update_mask_0/n1222 ), .CP(
        clk), .Q(\update_mask_0/reg_out[9][4] ) );
  dff_sg \update_mask_0/reg_out_reg[9][5]  ( .D(\update_mask_0/n1221 ), .CP(
        clk), .Q(\update_mask_0/reg_out[9][5] ) );
  dff_sg \update_mask_0/reg_out_reg[9][6]  ( .D(\update_mask_0/n1220 ), .CP(
        clk), .Q(\update_mask_0/reg_out[9][6] ) );
  dff_sg \update_mask_0/reg_out_reg[9][7]  ( .D(\update_mask_0/n1219 ), .CP(
        clk), .Q(\update_mask_0/reg_out[9][7] ) );
  dff_sg \update_mask_0/reg_out_reg[9][8]  ( .D(\update_mask_0/n1218 ), .CP(
        clk), .Q(\update_mask_0/reg_out[9][8] ) );
  dff_sg \update_mask_0/reg_out_reg[9][9]  ( .D(\update_mask_0/n1217 ), .CP(
        clk), .Q(\update_mask_0/reg_out[9][9] ) );
  dff_sg \update_mask_0/reg_out_reg[9][10]  ( .D(\update_mask_0/n1216 ), .CP(
        clk), .Q(\update_mask_0/reg_out[9][10] ) );
  dff_sg \update_mask_0/reg_out_reg[9][11]  ( .D(\update_mask_0/n1215 ), .CP(
        clk), .Q(\update_mask_0/reg_out[9][11] ) );
  dff_sg \update_mask_0/reg_out_reg[9][12]  ( .D(\update_mask_0/n1214 ), .CP(
        clk), .Q(\update_mask_0/reg_out[9][12] ) );
  dff_sg \update_mask_0/reg_out_reg[9][13]  ( .D(\update_mask_0/n1213 ), .CP(
        clk), .Q(\update_mask_0/reg_out[9][13] ) );
  dff_sg \update_mask_0/reg_out_reg[9][14]  ( .D(\update_mask_0/n1212 ), .CP(
        clk), .Q(\update_mask_0/reg_out[9][14] ) );
  dff_sg \update_mask_0/reg_out_reg[9][15]  ( .D(\update_mask_0/n1211 ), .CP(
        clk), .Q(\update_mask_0/reg_out[9][15] ) );
  dff_sg \update_mask_0/reg_out_reg[9][16]  ( .D(\update_mask_0/n1210 ), .CP(
        clk), .Q(\update_mask_0/reg_out[9][16] ) );
  dff_sg \update_mask_0/reg_out_reg[9][17]  ( .D(\update_mask_0/n1209 ), .CP(
        clk), .Q(\update_mask_0/reg_out[9][17] ) );
  dff_sg \update_mask_0/reg_out_reg[9][18]  ( .D(\update_mask_0/n1208 ), .CP(
        clk), .Q(\update_mask_0/reg_out[9][18] ) );
  dff_sg \update_mask_0/reg_out_reg[9][19]  ( .D(\update_mask_0/n1207 ), .CP(
        clk), .Q(\update_mask_0/reg_out[9][19] ) );
  dff_sg \update_mask_0/reg_out_reg[10][0]  ( .D(\update_mask_0/n1206 ), .CP(
        clk), .Q(\update_mask_0/reg_out[10][0] ) );
  dff_sg \update_mask_0/reg_out_reg[10][1]  ( .D(\update_mask_0/n1205 ), .CP(
        clk), .Q(\update_mask_0/reg_out[10][1] ) );
  dff_sg \update_mask_0/reg_out_reg[10][2]  ( .D(\update_mask_0/n1204 ), .CP(
        clk), .Q(\update_mask_0/reg_out[10][2] ) );
  dff_sg \update_mask_0/reg_out_reg[10][3]  ( .D(\update_mask_0/n1203 ), .CP(
        clk), .Q(\update_mask_0/reg_out[10][3] ) );
  dff_sg \update_mask_0/reg_out_reg[10][4]  ( .D(\update_mask_0/n1202 ), .CP(
        clk), .Q(\update_mask_0/reg_out[10][4] ) );
  dff_sg \update_mask_0/reg_out_reg[10][5]  ( .D(\update_mask_0/n1201 ), .CP(
        clk), .Q(\update_mask_0/reg_out[10][5] ) );
  dff_sg \update_mask_0/reg_out_reg[10][6]  ( .D(\update_mask_0/n1200 ), .CP(
        clk), .Q(\update_mask_0/reg_out[10][6] ) );
  dff_sg \update_mask_0/reg_out_reg[10][7]  ( .D(\update_mask_0/n1199 ), .CP(
        clk), .Q(\update_mask_0/reg_out[10][7] ) );
  dff_sg \update_mask_0/reg_out_reg[10][8]  ( .D(\update_mask_0/n1198 ), .CP(
        clk), .Q(\update_mask_0/reg_out[10][8] ) );
  dff_sg \update_mask_0/reg_out_reg[10][9]  ( .D(\update_mask_0/n1197 ), .CP(
        clk), .Q(\update_mask_0/reg_out[10][9] ) );
  dff_sg \update_mask_0/reg_out_reg[10][10]  ( .D(\update_mask_0/n1196 ), .CP(
        clk), .Q(\update_mask_0/reg_out[10][10] ) );
  dff_sg \update_mask_0/reg_out_reg[10][11]  ( .D(\update_mask_0/n1195 ), .CP(
        clk), .Q(\update_mask_0/reg_out[10][11] ) );
  dff_sg \update_mask_0/reg_out_reg[10][12]  ( .D(\update_mask_0/n1194 ), .CP(
        clk), .Q(\update_mask_0/reg_out[10][12] ) );
  dff_sg \update_mask_0/reg_out_reg[10][13]  ( .D(\update_mask_0/n1193 ), .CP(
        clk), .Q(\update_mask_0/reg_out[10][13] ) );
  dff_sg \update_mask_0/reg_out_reg[10][14]  ( .D(\update_mask_0/n1192 ), .CP(
        clk), .Q(\update_mask_0/reg_out[10][14] ) );
  dff_sg \update_mask_0/reg_out_reg[10][15]  ( .D(\update_mask_0/n1191 ), .CP(
        clk), .Q(\update_mask_0/reg_out[10][15] ) );
  dff_sg \update_mask_0/reg_out_reg[10][16]  ( .D(\update_mask_0/n1190 ), .CP(
        clk), .Q(\update_mask_0/reg_out[10][16] ) );
  dff_sg \update_mask_0/reg_out_reg[10][17]  ( .D(\update_mask_0/n1189 ), .CP(
        clk), .Q(\update_mask_0/reg_out[10][17] ) );
  dff_sg \update_mask_0/reg_out_reg[10][18]  ( .D(\update_mask_0/n1188 ), .CP(
        clk), .Q(\update_mask_0/reg_out[10][18] ) );
  dff_sg \update_mask_0/reg_out_reg[10][19]  ( .D(\update_mask_0/n1187 ), .CP(
        clk), .Q(\update_mask_0/reg_out[10][19] ) );
  dff_sg \update_mask_0/reg_out_reg[11][0]  ( .D(\update_mask_0/n1186 ), .CP(
        clk), .Q(\update_mask_0/reg_out[11][0] ) );
  dff_sg \update_mask_0/reg_out_reg[11][1]  ( .D(\update_mask_0/n1185 ), .CP(
        clk), .Q(\update_mask_0/reg_out[11][1] ) );
  dff_sg \update_mask_0/reg_out_reg[11][2]  ( .D(\update_mask_0/n1184 ), .CP(
        clk), .Q(\update_mask_0/reg_out[11][2] ) );
  dff_sg \update_mask_0/reg_out_reg[11][3]  ( .D(\update_mask_0/n1183 ), .CP(
        clk), .Q(\update_mask_0/reg_out[11][3] ) );
  dff_sg \update_mask_0/reg_out_reg[11][4]  ( .D(\update_mask_0/n1182 ), .CP(
        clk), .Q(\update_mask_0/reg_out[11][4] ) );
  dff_sg \update_mask_0/reg_out_reg[11][5]  ( .D(\update_mask_0/n1181 ), .CP(
        clk), .Q(\update_mask_0/reg_out[11][5] ) );
  dff_sg \update_mask_0/reg_out_reg[11][6]  ( .D(\update_mask_0/n1180 ), .CP(
        clk), .Q(\update_mask_0/reg_out[11][6] ) );
  dff_sg \update_mask_0/reg_out_reg[11][7]  ( .D(\update_mask_0/n1179 ), .CP(
        clk), .Q(\update_mask_0/reg_out[11][7] ) );
  dff_sg \update_mask_0/reg_out_reg[11][8]  ( .D(\update_mask_0/n1178 ), .CP(
        clk), .Q(\update_mask_0/reg_out[11][8] ) );
  dff_sg \update_mask_0/reg_out_reg[11][9]  ( .D(\update_mask_0/n1177 ), .CP(
        clk), .Q(\update_mask_0/reg_out[11][9] ) );
  dff_sg \update_mask_0/reg_out_reg[11][10]  ( .D(\update_mask_0/n1176 ), .CP(
        clk), .Q(\update_mask_0/reg_out[11][10] ) );
  dff_sg \update_mask_0/reg_out_reg[11][11]  ( .D(\update_mask_0/n1175 ), .CP(
        clk), .Q(\update_mask_0/reg_out[11][11] ) );
  dff_sg \update_mask_0/reg_out_reg[11][12]  ( .D(\update_mask_0/n1174 ), .CP(
        clk), .Q(\update_mask_0/reg_out[11][12] ) );
  dff_sg \update_mask_0/reg_out_reg[11][13]  ( .D(\update_mask_0/n1173 ), .CP(
        clk), .Q(\update_mask_0/reg_out[11][13] ) );
  dff_sg \update_mask_0/reg_out_reg[11][14]  ( .D(\update_mask_0/n1172 ), .CP(
        clk), .Q(\update_mask_0/reg_out[11][14] ) );
  dff_sg \update_mask_0/reg_out_reg[11][15]  ( .D(\update_mask_0/n1171 ), .CP(
        clk), .Q(\update_mask_0/reg_out[11][15] ) );
  dff_sg \update_mask_0/reg_out_reg[11][16]  ( .D(\update_mask_0/n1170 ), .CP(
        clk), .Q(\update_mask_0/reg_out[11][16] ) );
  dff_sg \update_mask_0/reg_out_reg[11][17]  ( .D(\update_mask_0/n1169 ), .CP(
        clk), .Q(\update_mask_0/reg_out[11][17] ) );
  dff_sg \update_mask_0/reg_out_reg[11][18]  ( .D(\update_mask_0/n1168 ), .CP(
        clk), .Q(\update_mask_0/reg_out[11][18] ) );
  dff_sg \update_mask_0/reg_out_reg[11][19]  ( .D(\update_mask_0/n1167 ), .CP(
        clk), .Q(\update_mask_0/reg_out[11][19] ) );
  dff_sg \update_mask_0/reg_out_reg[12][0]  ( .D(\update_mask_0/n1166 ), .CP(
        clk), .Q(\update_mask_0/reg_out[12][0] ) );
  dff_sg \update_mask_0/reg_out_reg[12][1]  ( .D(\update_mask_0/n1165 ), .CP(
        clk), .Q(\update_mask_0/reg_out[12][1] ) );
  dff_sg \update_mask_0/reg_out_reg[12][2]  ( .D(\update_mask_0/n1164 ), .CP(
        clk), .Q(\update_mask_0/reg_out[12][2] ) );
  dff_sg \update_mask_0/reg_out_reg[12][3]  ( .D(\update_mask_0/n1163 ), .CP(
        clk), .Q(\update_mask_0/reg_out[12][3] ) );
  dff_sg \update_mask_0/reg_out_reg[12][4]  ( .D(\update_mask_0/n1162 ), .CP(
        clk), .Q(\update_mask_0/reg_out[12][4] ) );
  dff_sg \update_mask_0/reg_out_reg[12][5]  ( .D(\update_mask_0/n1161 ), .CP(
        clk), .Q(\update_mask_0/reg_out[12][5] ) );
  dff_sg \update_mask_0/reg_out_reg[12][6]  ( .D(\update_mask_0/n1160 ), .CP(
        clk), .Q(\update_mask_0/reg_out[12][6] ) );
  dff_sg \update_mask_0/reg_out_reg[12][7]  ( .D(\update_mask_0/n1159 ), .CP(
        clk), .Q(\update_mask_0/reg_out[12][7] ) );
  dff_sg \update_mask_0/reg_out_reg[12][8]  ( .D(\update_mask_0/n1158 ), .CP(
        clk), .Q(\update_mask_0/reg_out[12][8] ) );
  dff_sg \update_mask_0/reg_out_reg[12][9]  ( .D(\update_mask_0/n1157 ), .CP(
        clk), .Q(\update_mask_0/reg_out[12][9] ) );
  dff_sg \update_mask_0/reg_out_reg[12][10]  ( .D(\update_mask_0/n1156 ), .CP(
        clk), .Q(\update_mask_0/reg_out[12][10] ) );
  dff_sg \update_mask_0/reg_out_reg[12][11]  ( .D(\update_mask_0/n1155 ), .CP(
        clk), .Q(\update_mask_0/reg_out[12][11] ) );
  dff_sg \update_mask_0/reg_out_reg[12][12]  ( .D(\update_mask_0/n1154 ), .CP(
        clk), .Q(\update_mask_0/reg_out[12][12] ) );
  dff_sg \update_mask_0/reg_out_reg[12][13]  ( .D(\update_mask_0/n1153 ), .CP(
        clk), .Q(\update_mask_0/reg_out[12][13] ) );
  dff_sg \update_mask_0/reg_out_reg[12][14]  ( .D(\update_mask_0/n1152 ), .CP(
        clk), .Q(\update_mask_0/reg_out[12][14] ) );
  dff_sg \update_mask_0/reg_out_reg[12][15]  ( .D(\update_mask_0/n1151 ), .CP(
        clk), .Q(\update_mask_0/reg_out[12][15] ) );
  dff_sg \update_mask_0/reg_out_reg[12][16]  ( .D(\update_mask_0/n1150 ), .CP(
        clk), .Q(\update_mask_0/reg_out[12][16] ) );
  dff_sg \update_mask_0/reg_out_reg[12][17]  ( .D(\update_mask_0/n1149 ), .CP(
        clk), .Q(\update_mask_0/reg_out[12][17] ) );
  dff_sg \update_mask_0/reg_out_reg[12][18]  ( .D(\update_mask_0/n1148 ), .CP(
        clk), .Q(\update_mask_0/reg_out[12][18] ) );
  dff_sg \update_mask_0/reg_out_reg[12][19]  ( .D(\update_mask_0/n1147 ), .CP(
        clk), .Q(\update_mask_0/reg_out[12][19] ) );
  dff_sg \update_mask_0/reg_out_reg[13][0]  ( .D(\update_mask_0/n1146 ), .CP(
        clk), .Q(\update_mask_0/reg_out[13][0] ) );
  dff_sg \update_mask_0/reg_out_reg[13][1]  ( .D(\update_mask_0/n1145 ), .CP(
        clk), .Q(\update_mask_0/reg_out[13][1] ) );
  dff_sg \update_mask_0/reg_out_reg[13][2]  ( .D(\update_mask_0/n1144 ), .CP(
        clk), .Q(\update_mask_0/reg_out[13][2] ) );
  dff_sg \update_mask_0/reg_out_reg[13][3]  ( .D(\update_mask_0/n1143 ), .CP(
        clk), .Q(\update_mask_0/reg_out[13][3] ) );
  dff_sg \update_mask_0/reg_out_reg[13][4]  ( .D(\update_mask_0/n1142 ), .CP(
        clk), .Q(\update_mask_0/reg_out[13][4] ) );
  dff_sg \update_mask_0/reg_out_reg[13][5]  ( .D(\update_mask_0/n1141 ), .CP(
        clk), .Q(\update_mask_0/reg_out[13][5] ) );
  dff_sg \update_mask_0/reg_out_reg[13][6]  ( .D(\update_mask_0/n1140 ), .CP(
        clk), .Q(\update_mask_0/reg_out[13][6] ) );
  dff_sg \update_mask_0/reg_out_reg[13][7]  ( .D(\update_mask_0/n1139 ), .CP(
        clk), .Q(\update_mask_0/reg_out[13][7] ) );
  dff_sg \update_mask_0/reg_out_reg[13][8]  ( .D(\update_mask_0/n1138 ), .CP(
        clk), .Q(\update_mask_0/reg_out[13][8] ) );
  dff_sg \update_mask_0/reg_out_reg[13][9]  ( .D(\update_mask_0/n1137 ), .CP(
        clk), .Q(\update_mask_0/reg_out[13][9] ) );
  dff_sg \update_mask_0/reg_out_reg[13][10]  ( .D(\update_mask_0/n1136 ), .CP(
        clk), .Q(\update_mask_0/reg_out[13][10] ) );
  dff_sg \update_mask_0/reg_out_reg[13][11]  ( .D(\update_mask_0/n1135 ), .CP(
        clk), .Q(\update_mask_0/reg_out[13][11] ) );
  dff_sg \update_mask_0/reg_out_reg[13][12]  ( .D(\update_mask_0/n1134 ), .CP(
        clk), .Q(\update_mask_0/reg_out[13][12] ) );
  dff_sg \update_mask_0/reg_out_reg[13][13]  ( .D(\update_mask_0/n1133 ), .CP(
        clk), .Q(\update_mask_0/reg_out[13][13] ) );
  dff_sg \update_mask_0/reg_out_reg[13][14]  ( .D(\update_mask_0/n1132 ), .CP(
        clk), .Q(\update_mask_0/reg_out[13][14] ) );
  dff_sg \update_mask_0/reg_out_reg[13][15]  ( .D(\update_mask_0/n1131 ), .CP(
        clk), .Q(\update_mask_0/reg_out[13][15] ) );
  dff_sg \update_mask_0/reg_out_reg[13][16]  ( .D(\update_mask_0/n1130 ), .CP(
        clk), .Q(\update_mask_0/reg_out[13][16] ) );
  dff_sg \update_mask_0/reg_out_reg[13][17]  ( .D(\update_mask_0/n1129 ), .CP(
        clk), .Q(\update_mask_0/reg_out[13][17] ) );
  dff_sg \update_mask_0/reg_out_reg[13][18]  ( .D(\update_mask_0/n1128 ), .CP(
        clk), .Q(\update_mask_0/reg_out[13][18] ) );
  dff_sg \update_mask_0/reg_out_reg[13][19]  ( .D(\update_mask_0/n1127 ), .CP(
        clk), .Q(\update_mask_0/reg_out[13][19] ) );
  dff_sg \update_mask_0/reg_out_reg[14][0]  ( .D(\update_mask_0/n1126 ), .CP(
        clk), .Q(\update_mask_0/reg_out[14][0] ) );
  dff_sg \update_mask_0/reg_out_reg[14][1]  ( .D(\update_mask_0/n1125 ), .CP(
        clk), .Q(\update_mask_0/reg_out[14][1] ) );
  dff_sg \update_mask_0/reg_out_reg[14][2]  ( .D(\update_mask_0/n1124 ), .CP(
        clk), .Q(\update_mask_0/reg_out[14][2] ) );
  dff_sg \update_mask_0/reg_out_reg[14][3]  ( .D(\update_mask_0/n1123 ), .CP(
        clk), .Q(\update_mask_0/reg_out[14][3] ) );
  dff_sg \update_mask_0/reg_out_reg[14][4]  ( .D(\update_mask_0/n1122 ), .CP(
        clk), .Q(\update_mask_0/reg_out[14][4] ) );
  dff_sg \update_mask_0/reg_out_reg[14][5]  ( .D(\update_mask_0/n1121 ), .CP(
        clk), .Q(\update_mask_0/reg_out[14][5] ) );
  dff_sg \update_mask_0/reg_out_reg[14][6]  ( .D(\update_mask_0/n1120 ), .CP(
        clk), .Q(\update_mask_0/reg_out[14][6] ) );
  dff_sg \update_mask_0/reg_out_reg[14][7]  ( .D(\update_mask_0/n1119 ), .CP(
        clk), .Q(\update_mask_0/reg_out[14][7] ) );
  dff_sg \update_mask_0/reg_out_reg[14][8]  ( .D(\update_mask_0/n1118 ), .CP(
        clk), .Q(\update_mask_0/reg_out[14][8] ) );
  dff_sg \update_mask_0/reg_out_reg[14][9]  ( .D(\update_mask_0/n1117 ), .CP(
        clk), .Q(\update_mask_0/reg_out[14][9] ) );
  dff_sg \update_mask_0/reg_out_reg[14][10]  ( .D(\update_mask_0/n1116 ), .CP(
        clk), .Q(\update_mask_0/reg_out[14][10] ) );
  dff_sg \update_mask_0/reg_out_reg[14][11]  ( .D(\update_mask_0/n1115 ), .CP(
        clk), .Q(\update_mask_0/reg_out[14][11] ) );
  dff_sg \update_mask_0/reg_out_reg[14][12]  ( .D(\update_mask_0/n1114 ), .CP(
        clk), .Q(\update_mask_0/reg_out[14][12] ) );
  dff_sg \update_mask_0/reg_out_reg[14][13]  ( .D(\update_mask_0/n1113 ), .CP(
        clk), .Q(\update_mask_0/reg_out[14][13] ) );
  dff_sg \update_mask_0/reg_out_reg[14][14]  ( .D(\update_mask_0/n1112 ), .CP(
        clk), .Q(\update_mask_0/reg_out[14][14] ) );
  dff_sg \update_mask_0/reg_out_reg[14][15]  ( .D(\update_mask_0/n1111 ), .CP(
        clk), .Q(\update_mask_0/reg_out[14][15] ) );
  dff_sg \update_mask_0/reg_out_reg[14][16]  ( .D(\update_mask_0/n1110 ), .CP(
        clk), .Q(\update_mask_0/reg_out[14][16] ) );
  dff_sg \update_mask_0/reg_out_reg[14][17]  ( .D(\update_mask_0/n1109 ), .CP(
        clk), .Q(\update_mask_0/reg_out[14][17] ) );
  dff_sg \update_mask_0/reg_out_reg[14][18]  ( .D(\update_mask_0/n1108 ), .CP(
        clk), .Q(\update_mask_0/reg_out[14][18] ) );
  dff_sg \update_mask_0/reg_out_reg[14][19]  ( .D(\update_mask_0/n1107 ), .CP(
        clk), .Q(\update_mask_0/reg_out[14][19] ) );
  dff_sg \update_mask_0/reg_out_reg[15][0]  ( .D(\update_mask_0/n1106 ), .CP(
        clk), .Q(\update_mask_0/reg_out[15][0] ) );
  dff_sg \update_mask_0/reg_out_reg[15][1]  ( .D(\update_mask_0/n1105 ), .CP(
        clk), .Q(\update_mask_0/reg_out[15][1] ) );
  dff_sg \update_mask_0/reg_out_reg[15][2]  ( .D(\update_mask_0/n1104 ), .CP(
        clk), .Q(\update_mask_0/reg_out[15][2] ) );
  dff_sg \update_mask_0/reg_out_reg[15][3]  ( .D(\update_mask_0/n1103 ), .CP(
        clk), .Q(\update_mask_0/reg_out[15][3] ) );
  dff_sg \update_mask_0/reg_out_reg[15][4]  ( .D(\update_mask_0/n1102 ), .CP(
        clk), .Q(\update_mask_0/reg_out[15][4] ) );
  dff_sg \update_mask_0/reg_out_reg[15][5]  ( .D(\update_mask_0/n1101 ), .CP(
        clk), .Q(\update_mask_0/reg_out[15][5] ) );
  dff_sg \update_mask_0/reg_out_reg[15][6]  ( .D(\update_mask_0/n1100 ), .CP(
        clk), .Q(\update_mask_0/reg_out[15][6] ) );
  dff_sg \update_mask_0/reg_out_reg[15][7]  ( .D(\update_mask_0/n1099 ), .CP(
        clk), .Q(\update_mask_0/reg_out[15][7] ) );
  dff_sg \update_mask_0/reg_out_reg[15][8]  ( .D(\update_mask_0/n1098 ), .CP(
        clk), .Q(\update_mask_0/reg_out[15][8] ) );
  dff_sg \update_mask_0/reg_out_reg[15][9]  ( .D(\update_mask_0/n1097 ), .CP(
        clk), .Q(\update_mask_0/reg_out[15][9] ) );
  dff_sg \update_mask_0/reg_out_reg[15][10]  ( .D(\update_mask_0/n1096 ), .CP(
        clk), .Q(\update_mask_0/reg_out[15][10] ) );
  dff_sg \update_mask_0/reg_out_reg[15][11]  ( .D(\update_mask_0/n1095 ), .CP(
        clk), .Q(\update_mask_0/reg_out[15][11] ) );
  dff_sg \update_mask_0/reg_out_reg[15][12]  ( .D(\update_mask_0/n1094 ), .CP(
        clk), .Q(\update_mask_0/reg_out[15][12] ) );
  dff_sg \update_mask_0/reg_out_reg[15][13]  ( .D(\update_mask_0/n1093 ), .CP(
        clk), .Q(\update_mask_0/reg_out[15][13] ) );
  dff_sg \update_mask_0/reg_out_reg[15][14]  ( .D(\update_mask_0/n1092 ), .CP(
        clk), .Q(\update_mask_0/reg_out[15][14] ) );
  dff_sg \update_mask_0/reg_out_reg[15][15]  ( .D(\update_mask_0/n1091 ), .CP(
        clk), .Q(\update_mask_0/reg_out[15][15] ) );
  dff_sg \update_mask_0/reg_out_reg[15][16]  ( .D(\update_mask_0/n1090 ), .CP(
        clk), .Q(\update_mask_0/reg_out[15][16] ) );
  dff_sg \update_mask_0/reg_out_reg[15][17]  ( .D(\update_mask_0/n1089 ), .CP(
        clk), .Q(\update_mask_0/reg_out[15][17] ) );
  dff_sg \update_mask_0/reg_out_reg[15][18]  ( .D(\update_mask_0/n1088 ), .CP(
        clk), .Q(\update_mask_0/reg_out[15][18] ) );
  dff_sg \update_mask_0/reg_out_reg[15][19]  ( .D(\update_mask_0/n1087 ), .CP(
        clk), .Q(\update_mask_0/reg_out[15][19] ) );
  dff_sg \update_mask_0/state_reg[0]  ( .D(\update_mask_0/n1439 ), .CP(clk), 
        .Q(\mask_state[0] ) );
  dff_sg \update_mask_0/state_reg[1]  ( .D(\update_mask_0/n1440 ), .CP(clk), 
        .Q(\update_mask_0/n2986 ) );
  dff_sg \update_mask_0/m_pointer_reg[0]  ( .D(\update_mask_0/n1442 ), .CP(clk), .Q(\update_mask_0/N23 ) );
  dff_sg \update_output_0/o_im_reg[11][0]  ( .D(\update_output_0/n2922 ), .CP(
        clk), .Q(\o_im[11][0] ) );
  dff_sg \update_output_0/o_im_reg[11][1]  ( .D(\update_output_0/n2921 ), .CP(
        clk), .Q(\o_im[11][1] ) );
  dff_sg \update_output_0/o_im_reg[11][2]  ( .D(\update_output_0/n2920 ), .CP(
        clk), .Q(\o_im[11][2] ) );
  dff_sg \update_output_0/o_im_reg[11][3]  ( .D(\update_output_0/n2919 ), .CP(
        clk), .Q(\o_im[11][3] ) );
  dff_sg \update_output_0/o_im_reg[11][4]  ( .D(\update_output_0/n2918 ), .CP(
        clk), .Q(\o_im[11][4] ) );
  dff_sg \update_output_0/o_im_reg[11][5]  ( .D(\update_output_0/n2917 ), .CP(
        clk), .Q(\o_im[11][5] ) );
  dff_sg \update_output_0/o_im_reg[11][6]  ( .D(\update_output_0/n2916 ), .CP(
        clk), .Q(\o_im[11][6] ) );
  dff_sg \update_output_0/o_im_reg[11][7]  ( .D(\update_output_0/n2915 ), .CP(
        clk), .Q(\o_im[11][7] ) );
  dff_sg \update_output_0/o_im_reg[11][8]  ( .D(\update_output_0/n2914 ), .CP(
        clk), .Q(\o_im[11][8] ) );
  dff_sg \update_output_0/o_im_reg[11][9]  ( .D(\update_output_0/n2913 ), .CP(
        clk), .Q(\o_im[11][9] ) );
  dff_sg \update_output_0/o_im_reg[11][10]  ( .D(\update_output_0/n2912 ), 
        .CP(clk), .Q(\o_im[11][10] ) );
  dff_sg \update_output_0/o_im_reg[11][11]  ( .D(\update_output_0/n2911 ), 
        .CP(clk), .Q(\o_im[11][11] ) );
  dff_sg \update_output_0/o_im_reg[11][12]  ( .D(\update_output_0/n2910 ), 
        .CP(clk), .Q(\o_im[11][12] ) );
  dff_sg \update_output_0/o_im_reg[11][13]  ( .D(\update_output_0/n2909 ), 
        .CP(clk), .Q(\o_im[11][13] ) );
  dff_sg \update_output_0/o_im_reg[11][14]  ( .D(\update_output_0/n2908 ), 
        .CP(clk), .Q(\o_im[11][14] ) );
  dff_sg \update_output_0/o_im_reg[11][15]  ( .D(\update_output_0/n2907 ), 
        .CP(clk), .Q(\o_im[11][15] ) );
  dff_sg \update_output_0/o_im_reg[11][16]  ( .D(\update_output_0/n2906 ), 
        .CP(clk), .Q(\o_im[11][16] ) );
  dff_sg \update_output_0/o_im_reg[11][17]  ( .D(\update_output_0/n2905 ), 
        .CP(clk), .Q(\o_im[11][17] ) );
  dff_sg \update_output_0/o_im_reg[11][18]  ( .D(\update_output_0/n2904 ), 
        .CP(clk), .Q(\o_im[11][18] ) );
  dff_sg \update_output_0/o_im_reg[11][19]  ( .D(\update_output_0/n2903 ), 
        .CP(clk), .Q(\o_im[11][19] ) );
  dff_sg \update_output_0/o_im_reg[15][0]  ( .D(\update_output_0/n2842 ), .CP(
        clk), .Q(\o_im[15][0] ) );
  dff_sg \update_output_0/o_im_reg[15][1]  ( .D(\update_output_0/n2841 ), .CP(
        clk), .Q(\o_im[15][1] ) );
  dff_sg \update_output_0/o_im_reg[15][2]  ( .D(\update_output_0/n2840 ), .CP(
        clk), .Q(\o_im[15][2] ) );
  dff_sg \update_output_0/o_im_reg[15][3]  ( .D(\update_output_0/n2839 ), .CP(
        clk), .Q(\o_im[15][3] ) );
  dff_sg \update_output_0/o_im_reg[15][4]  ( .D(\update_output_0/n2838 ), .CP(
        clk), .Q(\o_im[15][4] ) );
  dff_sg \update_output_0/o_im_reg[15][5]  ( .D(\update_output_0/n2837 ), .CP(
        clk), .Q(\o_im[15][5] ) );
  dff_sg \update_output_0/o_im_reg[15][6]  ( .D(\update_output_0/n2836 ), .CP(
        clk), .Q(\o_im[15][6] ) );
  dff_sg \update_output_0/o_im_reg[15][7]  ( .D(\update_output_0/n2835 ), .CP(
        clk), .Q(\o_im[15][7] ) );
  dff_sg \update_output_0/o_im_reg[15][8]  ( .D(\update_output_0/n2834 ), .CP(
        clk), .Q(\o_im[15][8] ) );
  dff_sg \update_output_0/o_im_reg[15][9]  ( .D(\update_output_0/n2833 ), .CP(
        clk), .Q(\o_im[15][9] ) );
  dff_sg \update_output_0/o_im_reg[15][10]  ( .D(\update_output_0/n2832 ), 
        .CP(clk), .Q(\o_im[15][10] ) );
  dff_sg \update_output_0/o_im_reg[15][11]  ( .D(\update_output_0/n2831 ), 
        .CP(clk), .Q(\o_im[15][11] ) );
  dff_sg \update_output_0/o_im_reg[15][12]  ( .D(\update_output_0/n2830 ), 
        .CP(clk), .Q(\o_im[15][12] ) );
  dff_sg \update_output_0/o_im_reg[15][13]  ( .D(\update_output_0/n2829 ), 
        .CP(clk), .Q(\o_im[15][13] ) );
  dff_sg \update_output_0/o_im_reg[15][14]  ( .D(\update_output_0/n2828 ), 
        .CP(clk), .Q(\o_im[15][14] ) );
  dff_sg \update_output_0/o_im_reg[15][15]  ( .D(\update_output_0/n2827 ), 
        .CP(clk), .Q(\o_im[15][15] ) );
  dff_sg \update_output_0/o_im_reg[15][16]  ( .D(\update_output_0/n2826 ), 
        .CP(clk), .Q(\o_im[15][16] ) );
  dff_sg \update_output_0/o_im_reg[15][17]  ( .D(\update_output_0/n2825 ), 
        .CP(clk), .Q(\o_im[15][17] ) );
  dff_sg \update_output_0/o_im_reg[15][18]  ( .D(\update_output_0/n2824 ), 
        .CP(clk), .Q(\o_im[15][18] ) );
  dff_sg \update_output_0/o_im_reg[15][19]  ( .D(\update_output_0/n2823 ), 
        .CP(clk), .Q(\o_im[15][19] ) );
  dff_sg \update_output_0/o_im_reg[10][0]  ( .D(\update_output_0/n2942 ), .CP(
        clk), .Q(\o_im[10][0] ) );
  dff_sg \update_output_0/o_im_reg[10][1]  ( .D(\update_output_0/n2941 ), .CP(
        clk), .Q(\o_im[10][1] ) );
  dff_sg \update_output_0/o_im_reg[10][2]  ( .D(\update_output_0/n2940 ), .CP(
        clk), .Q(\o_im[10][2] ) );
  dff_sg \update_output_0/o_im_reg[10][3]  ( .D(\update_output_0/n2939 ), .CP(
        clk), .Q(\o_im[10][3] ) );
  dff_sg \update_output_0/o_im_reg[10][4]  ( .D(\update_output_0/n2938 ), .CP(
        clk), .Q(\o_im[10][4] ) );
  dff_sg \update_output_0/o_im_reg[10][5]  ( .D(\update_output_0/n2937 ), .CP(
        clk), .Q(\o_im[10][5] ) );
  dff_sg \update_output_0/o_im_reg[10][6]  ( .D(\update_output_0/n2936 ), .CP(
        clk), .Q(\o_im[10][6] ) );
  dff_sg \update_output_0/o_im_reg[10][7]  ( .D(\update_output_0/n2935 ), .CP(
        clk), .Q(\o_im[10][7] ) );
  dff_sg \update_output_0/o_im_reg[10][8]  ( .D(\update_output_0/n2934 ), .CP(
        clk), .Q(\o_im[10][8] ) );
  dff_sg \update_output_0/o_im_reg[10][9]  ( .D(\update_output_0/n2933 ), .CP(
        clk), .Q(\o_im[10][9] ) );
  dff_sg \update_output_0/o_im_reg[10][10]  ( .D(\update_output_0/n2932 ), 
        .CP(clk), .Q(\o_im[10][10] ) );
  dff_sg \update_output_0/o_im_reg[10][11]  ( .D(\update_output_0/n2931 ), 
        .CP(clk), .Q(\o_im[10][11] ) );
  dff_sg \update_output_0/o_im_reg[10][12]  ( .D(\update_output_0/n2930 ), 
        .CP(clk), .Q(\o_im[10][12] ) );
  dff_sg \update_output_0/o_im_reg[10][13]  ( .D(\update_output_0/n2929 ), 
        .CP(clk), .Q(\o_im[10][13] ) );
  dff_sg \update_output_0/o_im_reg[10][14]  ( .D(\update_output_0/n2928 ), 
        .CP(clk), .Q(\o_im[10][14] ) );
  dff_sg \update_output_0/o_im_reg[10][15]  ( .D(\update_output_0/n2927 ), 
        .CP(clk), .Q(\o_im[10][15] ) );
  dff_sg \update_output_0/o_im_reg[10][16]  ( .D(\update_output_0/n2926 ), 
        .CP(clk), .Q(\o_im[10][16] ) );
  dff_sg \update_output_0/o_im_reg[10][17]  ( .D(\update_output_0/n2925 ), 
        .CP(clk), .Q(\o_im[10][17] ) );
  dff_sg \update_output_0/o_im_reg[10][18]  ( .D(\update_output_0/n2924 ), 
        .CP(clk), .Q(\o_im[10][18] ) );
  dff_sg \update_output_0/o_im_reg[10][19]  ( .D(\update_output_0/n2923 ), 
        .CP(clk), .Q(\o_im[10][19] ) );
  dff_sg \update_output_0/o_im_reg[14][0]  ( .D(\update_output_0/n2862 ), .CP(
        clk), .Q(\o_im[14][0] ) );
  dff_sg \update_output_0/o_im_reg[14][1]  ( .D(\update_output_0/n2861 ), .CP(
        clk), .Q(\o_im[14][1] ) );
  dff_sg \update_output_0/o_im_reg[14][2]  ( .D(\update_output_0/n2860 ), .CP(
        clk), .Q(\o_im[14][2] ) );
  dff_sg \update_output_0/o_im_reg[14][3]  ( .D(\update_output_0/n2859 ), .CP(
        clk), .Q(\o_im[14][3] ) );
  dff_sg \update_output_0/o_im_reg[14][4]  ( .D(\update_output_0/n2858 ), .CP(
        clk), .Q(\o_im[14][4] ) );
  dff_sg \update_output_0/o_im_reg[14][5]  ( .D(\update_output_0/n2857 ), .CP(
        clk), .Q(\o_im[14][5] ) );
  dff_sg \update_output_0/o_im_reg[14][6]  ( .D(\update_output_0/n2856 ), .CP(
        clk), .Q(\o_im[14][6] ) );
  dff_sg \update_output_0/o_im_reg[14][7]  ( .D(\update_output_0/n2855 ), .CP(
        clk), .Q(\o_im[14][7] ) );
  dff_sg \update_output_0/o_im_reg[14][8]  ( .D(\update_output_0/n2854 ), .CP(
        clk), .Q(\o_im[14][8] ) );
  dff_sg \update_output_0/o_im_reg[14][9]  ( .D(\update_output_0/n2853 ), .CP(
        clk), .Q(\o_im[14][9] ) );
  dff_sg \update_output_0/o_im_reg[14][10]  ( .D(\update_output_0/n2852 ), 
        .CP(clk), .Q(\o_im[14][10] ) );
  dff_sg \update_output_0/o_im_reg[14][11]  ( .D(\update_output_0/n2851 ), 
        .CP(clk), .Q(\o_im[14][11] ) );
  dff_sg \update_output_0/o_im_reg[14][12]  ( .D(\update_output_0/n2850 ), 
        .CP(clk), .Q(\o_im[14][12] ) );
  dff_sg \update_output_0/o_im_reg[14][13]  ( .D(\update_output_0/n2849 ), 
        .CP(clk), .Q(\o_im[14][13] ) );
  dff_sg \update_output_0/o_im_reg[14][14]  ( .D(\update_output_0/n2848 ), 
        .CP(clk), .Q(\o_im[14][14] ) );
  dff_sg \update_output_0/o_im_reg[14][15]  ( .D(\update_output_0/n2847 ), 
        .CP(clk), .Q(\o_im[14][15] ) );
  dff_sg \update_output_0/o_im_reg[14][16]  ( .D(\update_output_0/n2846 ), 
        .CP(clk), .Q(\o_im[14][16] ) );
  dff_sg \update_output_0/o_im_reg[14][17]  ( .D(\update_output_0/n2845 ), 
        .CP(clk), .Q(\o_im[14][17] ) );
  dff_sg \update_output_0/o_im_reg[14][18]  ( .D(\update_output_0/n2844 ), 
        .CP(clk), .Q(\o_im[14][18] ) );
  dff_sg \update_output_0/o_im_reg[14][19]  ( .D(\update_output_0/n2843 ), 
        .CP(clk), .Q(\o_im[14][19] ) );
  dff_sg \update_output_0/o_im_reg[8][0]  ( .D(\update_output_0/n2982 ), .CP(
        clk), .Q(\o_im[8][0] ) );
  dff_sg \update_output_0/o_im_reg[8][1]  ( .D(\update_output_0/n2981 ), .CP(
        clk), .Q(\o_im[8][1] ) );
  dff_sg \update_output_0/o_im_reg[8][2]  ( .D(\update_output_0/n2980 ), .CP(
        clk), .Q(\o_im[8][2] ) );
  dff_sg \update_output_0/o_im_reg[8][3]  ( .D(\update_output_0/n2979 ), .CP(
        clk), .Q(\o_im[8][3] ) );
  dff_sg \update_output_0/o_im_reg[8][4]  ( .D(\update_output_0/n2978 ), .CP(
        clk), .Q(\o_im[8][4] ) );
  dff_sg \update_output_0/o_im_reg[8][5]  ( .D(\update_output_0/n2977 ), .CP(
        clk), .Q(\o_im[8][5] ) );
  dff_sg \update_output_0/o_im_reg[8][6]  ( .D(\update_output_0/n2976 ), .CP(
        clk), .Q(\o_im[8][6] ) );
  dff_sg \update_output_0/o_im_reg[8][7]  ( .D(\update_output_0/n2975 ), .CP(
        clk), .Q(\o_im[8][7] ) );
  dff_sg \update_output_0/o_im_reg[8][8]  ( .D(\update_output_0/n2974 ), .CP(
        clk), .Q(\o_im[8][8] ) );
  dff_sg \update_output_0/o_im_reg[8][9]  ( .D(\update_output_0/n2973 ), .CP(
        clk), .Q(\o_im[8][9] ) );
  dff_sg \update_output_0/o_im_reg[8][10]  ( .D(\update_output_0/n2972 ), .CP(
        clk), .Q(\o_im[8][10] ) );
  dff_sg \update_output_0/o_im_reg[8][11]  ( .D(\update_output_0/n2971 ), .CP(
        clk), .Q(\o_im[8][11] ) );
  dff_sg \update_output_0/o_im_reg[8][12]  ( .D(\update_output_0/n2970 ), .CP(
        clk), .Q(\o_im[8][12] ) );
  dff_sg \update_output_0/o_im_reg[8][13]  ( .D(\update_output_0/n2969 ), .CP(
        clk), .Q(\o_im[8][13] ) );
  dff_sg \update_output_0/o_im_reg[8][14]  ( .D(\update_output_0/n2968 ), .CP(
        clk), .Q(\o_im[8][14] ) );
  dff_sg \update_output_0/o_im_reg[8][15]  ( .D(\update_output_0/n2967 ), .CP(
        clk), .Q(\o_im[8][15] ) );
  dff_sg \update_output_0/o_im_reg[8][16]  ( .D(\update_output_0/n2966 ), .CP(
        clk), .Q(\o_im[8][16] ) );
  dff_sg \update_output_0/o_im_reg[8][17]  ( .D(\update_output_0/n2965 ), .CP(
        clk), .Q(\o_im[8][17] ) );
  dff_sg \update_output_0/o_im_reg[8][18]  ( .D(\update_output_0/n2964 ), .CP(
        clk), .Q(\o_im[8][18] ) );
  dff_sg \update_output_0/o_im_reg[8][19]  ( .D(\update_output_0/n2963 ), .CP(
        clk), .Q(\o_im[8][19] ) );
  dff_sg \update_output_0/o_im_reg[12][0]  ( .D(\update_output_0/n2902 ), .CP(
        clk), .Q(\o_im[12][0] ) );
  dff_sg \update_output_0/o_im_reg[12][1]  ( .D(\update_output_0/n2901 ), .CP(
        clk), .Q(\o_im[12][1] ) );
  dff_sg \update_output_0/o_im_reg[12][2]  ( .D(\update_output_0/n2900 ), .CP(
        clk), .Q(\o_im[12][2] ) );
  dff_sg \update_output_0/o_im_reg[12][3]  ( .D(\update_output_0/n2899 ), .CP(
        clk), .Q(\o_im[12][3] ) );
  dff_sg \update_output_0/o_im_reg[12][4]  ( .D(\update_output_0/n2898 ), .CP(
        clk), .Q(\o_im[12][4] ) );
  dff_sg \update_output_0/o_im_reg[12][5]  ( .D(\update_output_0/n2897 ), .CP(
        clk), .Q(\o_im[12][5] ) );
  dff_sg \update_output_0/o_im_reg[12][6]  ( .D(\update_output_0/n2896 ), .CP(
        clk), .Q(\o_im[12][6] ) );
  dff_sg \update_output_0/o_im_reg[12][7]  ( .D(\update_output_0/n2895 ), .CP(
        clk), .Q(\o_im[12][7] ) );
  dff_sg \update_output_0/o_im_reg[12][8]  ( .D(\update_output_0/n2894 ), .CP(
        clk), .Q(\o_im[12][8] ) );
  dff_sg \update_output_0/o_im_reg[12][9]  ( .D(\update_output_0/n2893 ), .CP(
        clk), .Q(\o_im[12][9] ) );
  dff_sg \update_output_0/o_im_reg[12][10]  ( .D(\update_output_0/n2892 ), 
        .CP(clk), .Q(\o_im[12][10] ) );
  dff_sg \update_output_0/o_im_reg[12][11]  ( .D(\update_output_0/n2891 ), 
        .CP(clk), .Q(\o_im[12][11] ) );
  dff_sg \update_output_0/o_im_reg[12][12]  ( .D(\update_output_0/n2890 ), 
        .CP(clk), .Q(\o_im[12][12] ) );
  dff_sg \update_output_0/o_im_reg[12][13]  ( .D(\update_output_0/n2889 ), 
        .CP(clk), .Q(\o_im[12][13] ) );
  dff_sg \update_output_0/o_im_reg[12][14]  ( .D(\update_output_0/n2888 ), 
        .CP(clk), .Q(\o_im[12][14] ) );
  dff_sg \update_output_0/o_im_reg[12][15]  ( .D(\update_output_0/n2887 ), 
        .CP(clk), .Q(\o_im[12][15] ) );
  dff_sg \update_output_0/o_im_reg[12][16]  ( .D(\update_output_0/n2886 ), 
        .CP(clk), .Q(\o_im[12][16] ) );
  dff_sg \update_output_0/o_im_reg[12][17]  ( .D(\update_output_0/n2885 ), 
        .CP(clk), .Q(\o_im[12][17] ) );
  dff_sg \update_output_0/o_im_reg[12][18]  ( .D(\update_output_0/n2884 ), 
        .CP(clk), .Q(\o_im[12][18] ) );
  dff_sg \update_output_0/o_im_reg[12][19]  ( .D(\update_output_0/n2883 ), 
        .CP(clk), .Q(\o_im[12][19] ) );
  dff_sg \update_output_0/o_im_reg[9][0]  ( .D(\update_output_0/n2962 ), .CP(
        clk), .Q(\o_im[9][0] ) );
  dff_sg \update_output_0/o_im_reg[9][1]  ( .D(\update_output_0/n2961 ), .CP(
        clk), .Q(\o_im[9][1] ) );
  dff_sg \update_output_0/o_im_reg[9][2]  ( .D(\update_output_0/n2960 ), .CP(
        clk), .Q(\o_im[9][2] ) );
  dff_sg \update_output_0/o_im_reg[9][3]  ( .D(\update_output_0/n2959 ), .CP(
        clk), .Q(\o_im[9][3] ) );
  dff_sg \update_output_0/o_im_reg[9][4]  ( .D(\update_output_0/n2958 ), .CP(
        clk), .Q(\o_im[9][4] ) );
  dff_sg \update_output_0/o_im_reg[9][5]  ( .D(\update_output_0/n2957 ), .CP(
        clk), .Q(\o_im[9][5] ) );
  dff_sg \update_output_0/o_im_reg[9][6]  ( .D(\update_output_0/n2956 ), .CP(
        clk), .Q(\o_im[9][6] ) );
  dff_sg \update_output_0/o_im_reg[9][7]  ( .D(\update_output_0/n2955 ), .CP(
        clk), .Q(\o_im[9][7] ) );
  dff_sg \update_output_0/o_im_reg[9][8]  ( .D(\update_output_0/n2954 ), .CP(
        clk), .Q(\o_im[9][8] ) );
  dff_sg \update_output_0/o_im_reg[9][9]  ( .D(\update_output_0/n2953 ), .CP(
        clk), .Q(\o_im[9][9] ) );
  dff_sg \update_output_0/o_im_reg[9][10]  ( .D(\update_output_0/n2952 ), .CP(
        clk), .Q(\o_im[9][10] ) );
  dff_sg \update_output_0/o_im_reg[9][11]  ( .D(\update_output_0/n2951 ), .CP(
        clk), .Q(\o_im[9][11] ) );
  dff_sg \update_output_0/o_im_reg[9][12]  ( .D(\update_output_0/n2950 ), .CP(
        clk), .Q(\o_im[9][12] ) );
  dff_sg \update_output_0/o_im_reg[9][13]  ( .D(\update_output_0/n2949 ), .CP(
        clk), .Q(\o_im[9][13] ) );
  dff_sg \update_output_0/o_im_reg[9][14]  ( .D(\update_output_0/n2948 ), .CP(
        clk), .Q(\o_im[9][14] ) );
  dff_sg \update_output_0/o_im_reg[9][15]  ( .D(\update_output_0/n2947 ), .CP(
        clk), .Q(\o_im[9][15] ) );
  dff_sg \update_output_0/o_im_reg[9][16]  ( .D(\update_output_0/n2946 ), .CP(
        clk), .Q(\o_im[9][16] ) );
  dff_sg \update_output_0/o_im_reg[9][17]  ( .D(\update_output_0/n2945 ), .CP(
        clk), .Q(\o_im[9][17] ) );
  dff_sg \update_output_0/o_im_reg[9][18]  ( .D(\update_output_0/n2944 ), .CP(
        clk), .Q(\o_im[9][18] ) );
  dff_sg \update_output_0/o_im_reg[9][19]  ( .D(\update_output_0/n2943 ), .CP(
        clk), .Q(\o_im[9][19] ) );
  dff_sg \update_output_0/o_im_reg[13][0]  ( .D(\update_output_0/n2882 ), .CP(
        clk), .Q(\o_im[13][0] ) );
  dff_sg \update_output_0/o_im_reg[13][1]  ( .D(\update_output_0/n2881 ), .CP(
        clk), .Q(\o_im[13][1] ) );
  dff_sg \update_output_0/o_im_reg[13][2]  ( .D(\update_output_0/n2880 ), .CP(
        clk), .Q(\o_im[13][2] ) );
  dff_sg \update_output_0/o_im_reg[13][3]  ( .D(\update_output_0/n2879 ), .CP(
        clk), .Q(\o_im[13][3] ) );
  dff_sg \update_output_0/o_im_reg[13][4]  ( .D(\update_output_0/n2878 ), .CP(
        clk), .Q(\o_im[13][4] ) );
  dff_sg \update_output_0/o_im_reg[13][5]  ( .D(\update_output_0/n2877 ), .CP(
        clk), .Q(\o_im[13][5] ) );
  dff_sg \update_output_0/o_im_reg[13][6]  ( .D(\update_output_0/n2876 ), .CP(
        clk), .Q(\o_im[13][6] ) );
  dff_sg \update_output_0/o_im_reg[13][7]  ( .D(\update_output_0/n2875 ), .CP(
        clk), .Q(\o_im[13][7] ) );
  dff_sg \update_output_0/o_im_reg[13][8]  ( .D(\update_output_0/n2874 ), .CP(
        clk), .Q(\o_im[13][8] ) );
  dff_sg \update_output_0/o_im_reg[13][9]  ( .D(\update_output_0/n2873 ), .CP(
        clk), .Q(\o_im[13][9] ) );
  dff_sg \update_output_0/o_im_reg[13][10]  ( .D(\update_output_0/n2872 ), 
        .CP(clk), .Q(\o_im[13][10] ) );
  dff_sg \update_output_0/o_im_reg[13][11]  ( .D(\update_output_0/n2871 ), 
        .CP(clk), .Q(\o_im[13][11] ) );
  dff_sg \update_output_0/o_im_reg[13][12]  ( .D(\update_output_0/n2870 ), 
        .CP(clk), .Q(\o_im[13][12] ) );
  dff_sg \update_output_0/o_im_reg[13][13]  ( .D(\update_output_0/n2869 ), 
        .CP(clk), .Q(\o_im[13][13] ) );
  dff_sg \update_output_0/o_im_reg[13][14]  ( .D(\update_output_0/n2868 ), 
        .CP(clk), .Q(\o_im[13][14] ) );
  dff_sg \update_output_0/o_im_reg[13][15]  ( .D(\update_output_0/n2867 ), 
        .CP(clk), .Q(\o_im[13][15] ) );
  dff_sg \update_output_0/o_im_reg[13][16]  ( .D(\update_output_0/n2866 ), 
        .CP(clk), .Q(\o_im[13][16] ) );
  dff_sg \update_output_0/o_im_reg[13][17]  ( .D(\update_output_0/n2865 ), 
        .CP(clk), .Q(\o_im[13][17] ) );
  dff_sg \update_output_0/o_im_reg[13][18]  ( .D(\update_output_0/n2864 ), 
        .CP(clk), .Q(\o_im[13][18] ) );
  dff_sg \update_output_0/o_im_reg[13][19]  ( .D(\update_output_0/n2863 ), 
        .CP(clk), .Q(\o_im[13][19] ) );
  dff_sg \update_output_0/o_im_reg[1][0]  ( .D(\update_output_0/n3122 ), .CP(
        clk), .Q(\o_im[1][0] ) );
  dff_sg \update_output_0/o_im_reg[1][1]  ( .D(\update_output_0/n3121 ), .CP(
        clk), .Q(\o_im[1][1] ) );
  dff_sg \update_output_0/o_im_reg[1][2]  ( .D(\update_output_0/n3120 ), .CP(
        clk), .Q(\o_im[1][2] ) );
  dff_sg \update_output_0/o_im_reg[1][3]  ( .D(\update_output_0/n3119 ), .CP(
        clk), .Q(\o_im[1][3] ) );
  dff_sg \update_output_0/o_im_reg[1][4]  ( .D(\update_output_0/n3118 ), .CP(
        clk), .Q(\o_im[1][4] ) );
  dff_sg \update_output_0/o_im_reg[1][5]  ( .D(\update_output_0/n3117 ), .CP(
        clk), .Q(\o_im[1][5] ) );
  dff_sg \update_output_0/o_im_reg[1][6]  ( .D(\update_output_0/n3116 ), .CP(
        clk), .Q(\o_im[1][6] ) );
  dff_sg \update_output_0/o_im_reg[1][7]  ( .D(\update_output_0/n3115 ), .CP(
        clk), .Q(\o_im[1][7] ) );
  dff_sg \update_output_0/o_im_reg[1][8]  ( .D(\update_output_0/n3114 ), .CP(
        clk), .Q(\o_im[1][8] ) );
  dff_sg \update_output_0/o_im_reg[1][9]  ( .D(\update_output_0/n3113 ), .CP(
        clk), .Q(\o_im[1][9] ) );
  dff_sg \update_output_0/o_im_reg[1][10]  ( .D(\update_output_0/n3112 ), .CP(
        clk), .Q(\o_im[1][10] ) );
  dff_sg \update_output_0/o_im_reg[1][11]  ( .D(\update_output_0/n3111 ), .CP(
        clk), .Q(\o_im[1][11] ) );
  dff_sg \update_output_0/o_im_reg[1][12]  ( .D(\update_output_0/n3110 ), .CP(
        clk), .Q(\o_im[1][12] ) );
  dff_sg \update_output_0/o_im_reg[1][13]  ( .D(\update_output_0/n3109 ), .CP(
        clk), .Q(\o_im[1][13] ) );
  dff_sg \update_output_0/o_im_reg[1][14]  ( .D(\update_output_0/n3108 ), .CP(
        clk), .Q(\o_im[1][14] ) );
  dff_sg \update_output_0/o_im_reg[1][15]  ( .D(\update_output_0/n3107 ), .CP(
        clk), .Q(\o_im[1][15] ) );
  dff_sg \update_output_0/o_im_reg[1][16]  ( .D(\update_output_0/n3106 ), .CP(
        clk), .Q(\o_im[1][16] ) );
  dff_sg \update_output_0/o_im_reg[1][17]  ( .D(\update_output_0/n3105 ), .CP(
        clk), .Q(\o_im[1][17] ) );
  dff_sg \update_output_0/o_im_reg[1][18]  ( .D(\update_output_0/n3104 ), .CP(
        clk), .Q(\o_im[1][18] ) );
  dff_sg \update_output_0/o_im_reg[1][19]  ( .D(\update_output_0/n3103 ), .CP(
        clk), .Q(\o_im[1][19] ) );
  dff_sg \update_output_0/o_im_reg[3][0]  ( .D(\update_output_0/n3082 ), .CP(
        clk), .Q(\o_im[3][0] ) );
  dff_sg \update_output_0/o_im_reg[3][1]  ( .D(\update_output_0/n3081 ), .CP(
        clk), .Q(\o_im[3][1] ) );
  dff_sg \update_output_0/o_im_reg[3][2]  ( .D(\update_output_0/n3080 ), .CP(
        clk), .Q(\o_im[3][2] ) );
  dff_sg \update_output_0/o_im_reg[3][3]  ( .D(\update_output_0/n3079 ), .CP(
        clk), .Q(\o_im[3][3] ) );
  dff_sg \update_output_0/o_im_reg[3][4]  ( .D(\update_output_0/n3078 ), .CP(
        clk), .Q(\o_im[3][4] ) );
  dff_sg \update_output_0/o_im_reg[3][5]  ( .D(\update_output_0/n3077 ), .CP(
        clk), .Q(\o_im[3][5] ) );
  dff_sg \update_output_0/o_im_reg[3][6]  ( .D(\update_output_0/n3076 ), .CP(
        clk), .Q(\o_im[3][6] ) );
  dff_sg \update_output_0/o_im_reg[3][7]  ( .D(\update_output_0/n3075 ), .CP(
        clk), .Q(\o_im[3][7] ) );
  dff_sg \update_output_0/o_im_reg[3][8]  ( .D(\update_output_0/n3074 ), .CP(
        clk), .Q(\o_im[3][8] ) );
  dff_sg \update_output_0/o_im_reg[3][9]  ( .D(\update_output_0/n3073 ), .CP(
        clk), .Q(\o_im[3][9] ) );
  dff_sg \update_output_0/o_im_reg[3][10]  ( .D(\update_output_0/n3072 ), .CP(
        clk), .Q(\o_im[3][10] ) );
  dff_sg \update_output_0/o_im_reg[3][11]  ( .D(\update_output_0/n3071 ), .CP(
        clk), .Q(\o_im[3][11] ) );
  dff_sg \update_output_0/o_im_reg[3][12]  ( .D(\update_output_0/n3070 ), .CP(
        clk), .Q(\o_im[3][12] ) );
  dff_sg \update_output_0/o_im_reg[3][13]  ( .D(\update_output_0/n3069 ), .CP(
        clk), .Q(\o_im[3][13] ) );
  dff_sg \update_output_0/o_im_reg[3][14]  ( .D(\update_output_0/n3068 ), .CP(
        clk), .Q(\o_im[3][14] ) );
  dff_sg \update_output_0/o_im_reg[3][15]  ( .D(\update_output_0/n3067 ), .CP(
        clk), .Q(\o_im[3][15] ) );
  dff_sg \update_output_0/o_im_reg[3][16]  ( .D(\update_output_0/n3066 ), .CP(
        clk), .Q(\o_im[3][16] ) );
  dff_sg \update_output_0/o_im_reg[3][17]  ( .D(\update_output_0/n3065 ), .CP(
        clk), .Q(\o_im[3][17] ) );
  dff_sg \update_output_0/o_im_reg[3][18]  ( .D(\update_output_0/n3064 ), .CP(
        clk), .Q(\o_im[3][18] ) );
  dff_sg \update_output_0/o_im_reg[3][19]  ( .D(\update_output_0/n3063 ), .CP(
        clk), .Q(\o_im[3][19] ) );
  dff_sg \update_output_0/o_im_reg[5][0]  ( .D(\update_output_0/n3042 ), .CP(
        clk), .Q(\o_im[5][0] ) );
  dff_sg \update_output_0/o_im_reg[5][1]  ( .D(\update_output_0/n3041 ), .CP(
        clk), .Q(\o_im[5][1] ) );
  dff_sg \update_output_0/o_im_reg[5][2]  ( .D(\update_output_0/n3040 ), .CP(
        clk), .Q(\o_im[5][2] ) );
  dff_sg \update_output_0/o_im_reg[5][3]  ( .D(\update_output_0/n3039 ), .CP(
        clk), .Q(\o_im[5][3] ) );
  dff_sg \update_output_0/o_im_reg[5][4]  ( .D(\update_output_0/n3038 ), .CP(
        clk), .Q(\o_im[5][4] ) );
  dff_sg \update_output_0/o_im_reg[5][5]  ( .D(\update_output_0/n3037 ), .CP(
        clk), .Q(\o_im[5][5] ) );
  dff_sg \update_output_0/o_im_reg[5][6]  ( .D(\update_output_0/n3036 ), .CP(
        clk), .Q(\o_im[5][6] ) );
  dff_sg \update_output_0/o_im_reg[5][7]  ( .D(\update_output_0/n3035 ), .CP(
        clk), .Q(\o_im[5][7] ) );
  dff_sg \update_output_0/o_im_reg[5][8]  ( .D(\update_output_0/n3034 ), .CP(
        clk), .Q(\o_im[5][8] ) );
  dff_sg \update_output_0/o_im_reg[5][9]  ( .D(\update_output_0/n3033 ), .CP(
        clk), .Q(\o_im[5][9] ) );
  dff_sg \update_output_0/o_im_reg[5][10]  ( .D(\update_output_0/n3032 ), .CP(
        clk), .Q(\o_im[5][10] ) );
  dff_sg \update_output_0/o_im_reg[5][11]  ( .D(\update_output_0/n3031 ), .CP(
        clk), .Q(\o_im[5][11] ) );
  dff_sg \update_output_0/o_im_reg[5][12]  ( .D(\update_output_0/n3030 ), .CP(
        clk), .Q(\o_im[5][12] ) );
  dff_sg \update_output_0/o_im_reg[5][13]  ( .D(\update_output_0/n3029 ), .CP(
        clk), .Q(\o_im[5][13] ) );
  dff_sg \update_output_0/o_im_reg[5][14]  ( .D(\update_output_0/n3028 ), .CP(
        clk), .Q(\o_im[5][14] ) );
  dff_sg \update_output_0/o_im_reg[5][15]  ( .D(\update_output_0/n3027 ), .CP(
        clk), .Q(\o_im[5][15] ) );
  dff_sg \update_output_0/o_im_reg[5][16]  ( .D(\update_output_0/n3026 ), .CP(
        clk), .Q(\o_im[5][16] ) );
  dff_sg \update_output_0/o_im_reg[5][17]  ( .D(\update_output_0/n3025 ), .CP(
        clk), .Q(\o_im[5][17] ) );
  dff_sg \update_output_0/o_im_reg[5][18]  ( .D(\update_output_0/n3024 ), .CP(
        clk), .Q(\o_im[5][18] ) );
  dff_sg \update_output_0/o_im_reg[5][19]  ( .D(\update_output_0/n3023 ), .CP(
        clk), .Q(\o_im[5][19] ) );
  dff_sg \update_output_0/o_im_reg[7][0]  ( .D(\update_output_0/n3002 ), .CP(
        clk), .Q(\o_im[7][0] ) );
  dff_sg \update_output_0/o_im_reg[7][1]  ( .D(\update_output_0/n3001 ), .CP(
        clk), .Q(\o_im[7][1] ) );
  dff_sg \update_output_0/o_im_reg[7][2]  ( .D(\update_output_0/n3000 ), .CP(
        clk), .Q(\o_im[7][2] ) );
  dff_sg \update_output_0/o_im_reg[7][3]  ( .D(\update_output_0/n2999 ), .CP(
        clk), .Q(\o_im[7][3] ) );
  dff_sg \update_output_0/o_im_reg[7][4]  ( .D(\update_output_0/n2998 ), .CP(
        clk), .Q(\o_im[7][4] ) );
  dff_sg \update_output_0/o_im_reg[7][5]  ( .D(\update_output_0/n2997 ), .CP(
        clk), .Q(\o_im[7][5] ) );
  dff_sg \update_output_0/o_im_reg[7][6]  ( .D(\update_output_0/n2996 ), .CP(
        clk), .Q(\o_im[7][6] ) );
  dff_sg \update_output_0/o_im_reg[7][7]  ( .D(\update_output_0/n2995 ), .CP(
        clk), .Q(\o_im[7][7] ) );
  dff_sg \update_output_0/o_im_reg[7][8]  ( .D(\update_output_0/n2994 ), .CP(
        clk), .Q(\o_im[7][8] ) );
  dff_sg \update_output_0/o_im_reg[7][9]  ( .D(\update_output_0/n2993 ), .CP(
        clk), .Q(\o_im[7][9] ) );
  dff_sg \update_output_0/o_im_reg[7][10]  ( .D(\update_output_0/n2992 ), .CP(
        clk), .Q(\o_im[7][10] ) );
  dff_sg \update_output_0/o_im_reg[7][11]  ( .D(\update_output_0/n2991 ), .CP(
        clk), .Q(\o_im[7][11] ) );
  dff_sg \update_output_0/o_im_reg[7][12]  ( .D(\update_output_0/n2990 ), .CP(
        clk), .Q(\o_im[7][12] ) );
  dff_sg \update_output_0/o_im_reg[7][13]  ( .D(\update_output_0/n2989 ), .CP(
        clk), .Q(\o_im[7][13] ) );
  dff_sg \update_output_0/o_im_reg[7][14]  ( .D(\update_output_0/n2988 ), .CP(
        clk), .Q(\o_im[7][14] ) );
  dff_sg \update_output_0/o_im_reg[7][15]  ( .D(\update_output_0/n2987 ), .CP(
        clk), .Q(\o_im[7][15] ) );
  dff_sg \update_output_0/o_im_reg[7][16]  ( .D(\update_output_0/n2986 ), .CP(
        clk), .Q(\o_im[7][16] ) );
  dff_sg \update_output_0/o_im_reg[7][17]  ( .D(\update_output_0/n2985 ), .CP(
        clk), .Q(\o_im[7][17] ) );
  dff_sg \update_output_0/o_im_reg[7][18]  ( .D(\update_output_0/n2984 ), .CP(
        clk), .Q(\o_im[7][18] ) );
  dff_sg \update_output_0/o_im_reg[7][19]  ( .D(\update_output_0/n2983 ), .CP(
        clk), .Q(\o_im[7][19] ) );
  dff_sg \update_output_0/o_im_reg[4][0]  ( .D(\update_output_0/n3062 ), .CP(
        clk), .Q(\o_im[4][0] ) );
  dff_sg \update_output_0/o_im_reg[4][1]  ( .D(\update_output_0/n3061 ), .CP(
        clk), .Q(\o_im[4][1] ) );
  dff_sg \update_output_0/o_im_reg[4][2]  ( .D(\update_output_0/n3060 ), .CP(
        clk), .Q(\o_im[4][2] ) );
  dff_sg \update_output_0/o_im_reg[4][3]  ( .D(\update_output_0/n3059 ), .CP(
        clk), .Q(\o_im[4][3] ) );
  dff_sg \update_output_0/o_im_reg[4][4]  ( .D(\update_output_0/n3058 ), .CP(
        clk), .Q(\o_im[4][4] ) );
  dff_sg \update_output_0/o_im_reg[4][5]  ( .D(\update_output_0/n3057 ), .CP(
        clk), .Q(\o_im[4][5] ) );
  dff_sg \update_output_0/o_im_reg[4][6]  ( .D(\update_output_0/n3056 ), .CP(
        clk), .Q(\o_im[4][6] ) );
  dff_sg \update_output_0/o_im_reg[4][7]  ( .D(\update_output_0/n3055 ), .CP(
        clk), .Q(\o_im[4][7] ) );
  dff_sg \update_output_0/o_im_reg[4][8]  ( .D(\update_output_0/n3054 ), .CP(
        clk), .Q(\o_im[4][8] ) );
  dff_sg \update_output_0/o_im_reg[4][9]  ( .D(\update_output_0/n3053 ), .CP(
        clk), .Q(\o_im[4][9] ) );
  dff_sg \update_output_0/o_im_reg[4][10]  ( .D(\update_output_0/n3052 ), .CP(
        clk), .Q(\o_im[4][10] ) );
  dff_sg \update_output_0/o_im_reg[4][11]  ( .D(\update_output_0/n3051 ), .CP(
        clk), .Q(\o_im[4][11] ) );
  dff_sg \update_output_0/o_im_reg[4][12]  ( .D(\update_output_0/n3050 ), .CP(
        clk), .Q(\o_im[4][12] ) );
  dff_sg \update_output_0/o_im_reg[4][13]  ( .D(\update_output_0/n3049 ), .CP(
        clk), .Q(\o_im[4][13] ) );
  dff_sg \update_output_0/o_im_reg[4][14]  ( .D(\update_output_0/n3048 ), .CP(
        clk), .Q(\o_im[4][14] ) );
  dff_sg \update_output_0/o_im_reg[4][15]  ( .D(\update_output_0/n3047 ), .CP(
        clk), .Q(\o_im[4][15] ) );
  dff_sg \update_output_0/o_im_reg[4][16]  ( .D(\update_output_0/n3046 ), .CP(
        clk), .Q(\o_im[4][16] ) );
  dff_sg \update_output_0/o_im_reg[4][17]  ( .D(\update_output_0/n3045 ), .CP(
        clk), .Q(\o_im[4][17] ) );
  dff_sg \update_output_0/o_im_reg[4][18]  ( .D(\update_output_0/n3044 ), .CP(
        clk), .Q(\o_im[4][18] ) );
  dff_sg \update_output_0/o_im_reg[4][19]  ( .D(\update_output_0/n3043 ), .CP(
        clk), .Q(\o_im[4][19] ) );
  dff_sg \update_output_0/o_im_reg[0][0]  ( .D(\update_output_0/n3142 ), .CP(
        clk), .Q(\o_im[0][0] ) );
  dff_sg \update_output_0/o_im_reg[0][1]  ( .D(\update_output_0/n3141 ), .CP(
        clk), .Q(\o_im[0][1] ) );
  dff_sg \update_output_0/o_im_reg[0][2]  ( .D(\update_output_0/n3140 ), .CP(
        clk), .Q(\o_im[0][2] ) );
  dff_sg \update_output_0/o_im_reg[0][3]  ( .D(\update_output_0/n3139 ), .CP(
        clk), .Q(\o_im[0][3] ) );
  dff_sg \update_output_0/o_im_reg[0][4]  ( .D(\update_output_0/n3138 ), .CP(
        clk), .Q(\o_im[0][4] ) );
  dff_sg \update_output_0/o_im_reg[0][5]  ( .D(\update_output_0/n3137 ), .CP(
        clk), .Q(\o_im[0][5] ) );
  dff_sg \update_output_0/o_im_reg[0][6]  ( .D(\update_output_0/n3136 ), .CP(
        clk), .Q(\o_im[0][6] ) );
  dff_sg \update_output_0/o_im_reg[0][7]  ( .D(\update_output_0/n3135 ), .CP(
        clk), .Q(\o_im[0][7] ) );
  dff_sg \update_output_0/o_im_reg[0][8]  ( .D(\update_output_0/n3134 ), .CP(
        clk), .Q(\o_im[0][8] ) );
  dff_sg \update_output_0/o_im_reg[0][9]  ( .D(\update_output_0/n3133 ), .CP(
        clk), .Q(\o_im[0][9] ) );
  dff_sg \update_output_0/o_im_reg[0][10]  ( .D(\update_output_0/n3132 ), .CP(
        clk), .Q(\o_im[0][10] ) );
  dff_sg \update_output_0/o_im_reg[0][11]  ( .D(\update_output_0/n3131 ), .CP(
        clk), .Q(\o_im[0][11] ) );
  dff_sg \update_output_0/o_im_reg[0][12]  ( .D(\update_output_0/n3130 ), .CP(
        clk), .Q(\o_im[0][12] ) );
  dff_sg \update_output_0/o_im_reg[0][13]  ( .D(\update_output_0/n3129 ), .CP(
        clk), .Q(\o_im[0][13] ) );
  dff_sg \update_output_0/o_im_reg[0][14]  ( .D(\update_output_0/n3128 ), .CP(
        clk), .Q(\o_im[0][14] ) );
  dff_sg \update_output_0/o_im_reg[0][15]  ( .D(\update_output_0/n3127 ), .CP(
        clk), .Q(\o_im[0][15] ) );
  dff_sg \update_output_0/o_im_reg[0][16]  ( .D(\update_output_0/n3126 ), .CP(
        clk), .Q(\o_im[0][16] ) );
  dff_sg \update_output_0/o_im_reg[0][17]  ( .D(\update_output_0/n3125 ), .CP(
        clk), .Q(\o_im[0][17] ) );
  dff_sg \update_output_0/o_im_reg[0][18]  ( .D(\update_output_0/n3124 ), .CP(
        clk), .Q(\o_im[0][18] ) );
  dff_sg \update_output_0/o_im_reg[0][19]  ( .D(\update_output_0/n3123 ), .CP(
        clk), .Q(\o_im[0][19] ) );
  dff_sg \update_output_0/o_im_reg[2][0]  ( .D(\update_output_0/n3102 ), .CP(
        clk), .Q(\o_im[2][0] ) );
  dff_sg \update_output_0/o_im_reg[2][1]  ( .D(\update_output_0/n3101 ), .CP(
        clk), .Q(\o_im[2][1] ) );
  dff_sg \update_output_0/o_im_reg[2][2]  ( .D(\update_output_0/n3100 ), .CP(
        clk), .Q(\o_im[2][2] ) );
  dff_sg \update_output_0/o_im_reg[2][3]  ( .D(\update_output_0/n3099 ), .CP(
        clk), .Q(\o_im[2][3] ) );
  dff_sg \update_output_0/o_im_reg[2][4]  ( .D(\update_output_0/n3098 ), .CP(
        clk), .Q(\o_im[2][4] ) );
  dff_sg \update_output_0/o_im_reg[2][5]  ( .D(\update_output_0/n3097 ), .CP(
        clk), .Q(\o_im[2][5] ) );
  dff_sg \update_output_0/o_im_reg[2][6]  ( .D(\update_output_0/n3096 ), .CP(
        clk), .Q(\o_im[2][6] ) );
  dff_sg \update_output_0/o_im_reg[2][7]  ( .D(\update_output_0/n3095 ), .CP(
        clk), .Q(\o_im[2][7] ) );
  dff_sg \update_output_0/o_im_reg[2][8]  ( .D(\update_output_0/n3094 ), .CP(
        clk), .Q(\o_im[2][8] ) );
  dff_sg \update_output_0/o_im_reg[2][9]  ( .D(\update_output_0/n3093 ), .CP(
        clk), .Q(\o_im[2][9] ) );
  dff_sg \update_output_0/o_im_reg[2][10]  ( .D(\update_output_0/n3092 ), .CP(
        clk), .Q(\o_im[2][10] ) );
  dff_sg \update_output_0/o_im_reg[2][11]  ( .D(\update_output_0/n3091 ), .CP(
        clk), .Q(\o_im[2][11] ) );
  dff_sg \update_output_0/o_im_reg[2][12]  ( .D(\update_output_0/n3090 ), .CP(
        clk), .Q(\o_im[2][12] ) );
  dff_sg \update_output_0/o_im_reg[2][13]  ( .D(\update_output_0/n3089 ), .CP(
        clk), .Q(\o_im[2][13] ) );
  dff_sg \update_output_0/o_im_reg[2][14]  ( .D(\update_output_0/n3088 ), .CP(
        clk), .Q(\o_im[2][14] ) );
  dff_sg \update_output_0/o_im_reg[2][15]  ( .D(\update_output_0/n3087 ), .CP(
        clk), .Q(\o_im[2][15] ) );
  dff_sg \update_output_0/o_im_reg[2][16]  ( .D(\update_output_0/n3086 ), .CP(
        clk), .Q(\o_im[2][16] ) );
  dff_sg \update_output_0/o_im_reg[2][17]  ( .D(\update_output_0/n3085 ), .CP(
        clk), .Q(\o_im[2][17] ) );
  dff_sg \update_output_0/o_im_reg[2][18]  ( .D(\update_output_0/n3084 ), .CP(
        clk), .Q(\o_im[2][18] ) );
  dff_sg \update_output_0/o_im_reg[2][19]  ( .D(\update_output_0/n3083 ), .CP(
        clk), .Q(\o_im[2][19] ) );
  dff_sg \update_output_0/o_im_reg[6][0]  ( .D(\update_output_0/n3022 ), .CP(
        clk), .Q(\o_im[6][0] ) );
  dff_sg \update_output_0/o_im_reg[6][1]  ( .D(\update_output_0/n3021 ), .CP(
        clk), .Q(\o_im[6][1] ) );
  dff_sg \update_output_0/o_im_reg[6][2]  ( .D(\update_output_0/n3020 ), .CP(
        clk), .Q(\o_im[6][2] ) );
  dff_sg \update_output_0/o_im_reg[6][3]  ( .D(\update_output_0/n3019 ), .CP(
        clk), .Q(\o_im[6][3] ) );
  dff_sg \update_output_0/o_im_reg[6][4]  ( .D(\update_output_0/n3018 ), .CP(
        clk), .Q(\o_im[6][4] ) );
  dff_sg \update_output_0/o_im_reg[6][5]  ( .D(\update_output_0/n3017 ), .CP(
        clk), .Q(\o_im[6][5] ) );
  dff_sg \update_output_0/o_im_reg[6][6]  ( .D(\update_output_0/n3016 ), .CP(
        clk), .Q(\o_im[6][6] ) );
  dff_sg \update_output_0/o_im_reg[6][7]  ( .D(\update_output_0/n3015 ), .CP(
        clk), .Q(\o_im[6][7] ) );
  dff_sg \update_output_0/o_im_reg[6][8]  ( .D(\update_output_0/n3014 ), .CP(
        clk), .Q(\o_im[6][8] ) );
  dff_sg \update_output_0/o_im_reg[6][9]  ( .D(\update_output_0/n3013 ), .CP(
        clk), .Q(\o_im[6][9] ) );
  dff_sg \update_output_0/o_im_reg[6][10]  ( .D(\update_output_0/n3012 ), .CP(
        clk), .Q(\o_im[6][10] ) );
  dff_sg \update_output_0/o_im_reg[6][11]  ( .D(\update_output_0/n3011 ), .CP(
        clk), .Q(\o_im[6][11] ) );
  dff_sg \update_output_0/o_im_reg[6][12]  ( .D(\update_output_0/n3010 ), .CP(
        clk), .Q(\o_im[6][12] ) );
  dff_sg \update_output_0/o_im_reg[6][13]  ( .D(\update_output_0/n3009 ), .CP(
        clk), .Q(\o_im[6][13] ) );
  dff_sg \update_output_0/o_im_reg[6][14]  ( .D(\update_output_0/n3008 ), .CP(
        clk), .Q(\o_im[6][14] ) );
  dff_sg \update_output_0/o_im_reg[6][15]  ( .D(\update_output_0/n3007 ), .CP(
        clk), .Q(\o_im[6][15] ) );
  dff_sg \update_output_0/o_im_reg[6][16]  ( .D(\update_output_0/n3006 ), .CP(
        clk), .Q(\o_im[6][16] ) );
  dff_sg \update_output_0/o_im_reg[6][17]  ( .D(\update_output_0/n3005 ), .CP(
        clk), .Q(\o_im[6][17] ) );
  dff_sg \update_output_0/o_im_reg[6][18]  ( .D(\update_output_0/n3004 ), .CP(
        clk), .Q(\o_im[6][18] ) );
  dff_sg \update_output_0/o_im_reg[6][19]  ( .D(\update_output_0/n3003 ), .CP(
        clk), .Q(\o_im[6][19] ) );
  dff_sg \update_output_0/o_pointer_reg[3]  ( .D(\update_output_0/n3146 ), 
        .CP(clk), .Q(\update_output_0/N34 ) );
  dff_sg \update_output_0/o_pointer_reg[2]  ( .D(\update_output_0/n3143 ), 
        .CP(clk), .Q(\update_output_0/N33 ) );
  dff_sg \update_output_0/o_pointer_reg[1]  ( .D(\update_output_0/n3144 ), 
        .CP(clk), .Q(\update_output_0/N32 ) );
  dff_sg \update_output_0/o_pointer_reg[0]  ( .D(\update_output_0/n3145 ), 
        .CP(clk), .Q(\update_output_0/N31 ) );
  dff_sg \update_output_0/i_pointer_reg[2]  ( .D(\update_output_0/n3147 ), 
        .CP(clk), .Q(\update_output_0/N29 ) );
  dff_sg \update_output_0/i_pointer_reg[1]  ( .D(\update_output_0/n2822 ), 
        .CP(clk), .Q(\update_output_0/N28 ) );
  dff_sg \update_output_0/state_reg[0]  ( .D(\update_output_0/n3148 ), .CP(clk), .Q(\output_state[0] ) );
  dff_sg \update_output_0/state_reg[1]  ( .D(\update_output_0/n3149 ), .CP(clk), .Q(\update_output_0/n6096 ) );
  dff_sg \update_output_0/i_pointer_reg[3]  ( .D(\update_output_0/n3150 ), 
        .CP(clk), .Q(\update_output_0/N30 ) );
  dff_sg \update_output_0/i_pointer_reg[0]  ( .D(\update_output_0/n3151 ), 
        .CP(clk), .Q(\update_output_0/N27 ) );
  \**FFGEN**  \update_mask_0/increment_reg  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\update_mask_0/n952 ), .force_10(
        n733), .force_11(1'b0), .QN(\update_mask_0/n1835 ) );
  \**FFGEN**  \update_mask_0/o_mask_reg[31]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\update_mask_0/n956 ), .force_10(
        \update_mask_0/n957 ), .force_11(1'b0), .Q(o_mask[31]) );
  \**FFGEN**  \update_mask_0/o_mask_reg[30]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\update_mask_0/n960 ), .force_10(
        \update_mask_0/n961 ), .force_11(1'b0), .Q(o_mask[30]) );
  \**FFGEN**  \update_mask_0/o_mask_reg[29]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\update_mask_0/n964 ), .force_10(
        \update_mask_0/n965 ), .force_11(1'b0), .Q(o_mask[29]) );
  \**FFGEN**  \update_mask_0/o_mask_reg[28]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\update_mask_0/n968 ), .force_10(
        \update_mask_0/n969 ), .force_11(1'b0), .Q(o_mask[28]) );
  \**FFGEN**  \update_mask_0/o_mask_reg[27]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\update_mask_0/n972 ), .force_10(
        \update_mask_0/n973 ), .force_11(1'b0), .Q(o_mask[27]) );
  \**FFGEN**  \update_mask_0/o_mask_reg[26]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\update_mask_0/n976 ), .force_10(
        \update_mask_0/n977 ), .force_11(1'b0), .Q(o_mask[26]) );
  \**FFGEN**  \update_mask_0/o_mask_reg[25]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\update_mask_0/n980 ), .force_10(
        \update_mask_0/n981 ), .force_11(1'b0), .Q(o_mask[25]) );
  \**FFGEN**  \update_mask_0/o_mask_reg[24]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\update_mask_0/n984 ), .force_10(
        \update_mask_0/n985 ), .force_11(1'b0), .Q(o_mask[24]) );
  \**FFGEN**  \update_mask_0/o_mask_reg[23]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\update_mask_0/n988 ), .force_10(
        \update_mask_0/n989 ), .force_11(1'b0), .Q(o_mask[23]) );
  \**FFGEN**  \update_mask_0/o_mask_reg[22]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\update_mask_0/n992 ), .force_10(
        \update_mask_0/n993 ), .force_11(1'b0), .Q(o_mask[22]) );
  \**FFGEN**  \update_mask_0/o_mask_reg[21]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\update_mask_0/n996 ), .force_10(
        \update_mask_0/n997 ), .force_11(1'b0), .Q(o_mask[21]) );
  \**FFGEN**  \update_mask_0/o_mask_reg[20]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\update_mask_0/n1000 ), .force_10(
        \update_mask_0/n1001 ), .force_11(1'b0), .Q(o_mask[20]) );
  \**FFGEN**  \update_mask_0/o_mask_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\update_mask_0/n1004 ), .force_10(
        \update_mask_0/n1005 ), .force_11(1'b0), .Q(o_mask[19]) );
  \**FFGEN**  \update_mask_0/o_mask_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\update_mask_0/n1008 ), .force_10(
        \update_mask_0/n1009 ), .force_11(1'b0), .Q(o_mask[18]) );
  \**FFGEN**  \update_mask_0/o_mask_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\update_mask_0/n1012 ), .force_10(
        \update_mask_0/n1013 ), .force_11(1'b0), .Q(o_mask[17]) );
  \**FFGEN**  \update_mask_0/o_mask_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\update_mask_0/n1016 ), .force_10(
        \update_mask_0/n1017 ), .force_11(1'b0), .Q(o_mask[16]) );
  \**FFGEN**  \update_mask_0/o_mask_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\update_mask_0/n1020 ), .force_10(
        \update_mask_0/n1021 ), .force_11(1'b0), .Q(o_mask[15]) );
  \**FFGEN**  \update_mask_0/o_mask_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\update_mask_0/n1024 ), .force_10(
        \update_mask_0/n1025 ), .force_11(1'b0), .Q(o_mask[14]) );
  \**FFGEN**  \update_mask_0/o_mask_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\update_mask_0/n1028 ), .force_10(
        \update_mask_0/n1029 ), .force_11(1'b0), .Q(o_mask[13]) );
  \**FFGEN**  \update_mask_0/o_mask_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\update_mask_0/n1032 ), .force_10(
        \update_mask_0/n1033 ), .force_11(1'b0), .Q(o_mask[12]) );
  \**FFGEN**  \update_mask_0/o_mask_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\update_mask_0/n1036 ), .force_10(
        \update_mask_0/n1037 ), .force_11(1'b0), .Q(o_mask[11]) );
  \**FFGEN**  \update_mask_0/o_mask_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\update_mask_0/n1040 ), .force_10(
        \update_mask_0/n1041 ), .force_11(1'b0), .Q(o_mask[10]) );
  \**FFGEN**  \update_mask_0/o_mask_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\update_mask_0/n1044 ), .force_10(
        \update_mask_0/n1045 ), .force_11(1'b0), .Q(o_mask[9]) );
  \**FFGEN**  \update_mask_0/o_mask_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\update_mask_0/n1048 ), .force_10(
        \update_mask_0/n1049 ), .force_11(1'b0), .Q(o_mask[8]) );
  \**FFGEN**  \update_mask_0/o_mask_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\update_mask_0/n1052 ), .force_10(
        \update_mask_0/n1053 ), .force_11(1'b0), .Q(o_mask[7]) );
  \**FFGEN**  \update_mask_0/o_mask_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\update_mask_0/n1056 ), .force_10(
        \update_mask_0/n1057 ), .force_11(1'b0), .Q(o_mask[6]) );
  \**FFGEN**  \update_mask_0/o_mask_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\update_mask_0/n1060 ), .force_10(
        \update_mask_0/n1061 ), .force_11(1'b0), .Q(o_mask[5]) );
  \**FFGEN**  \update_mask_0/o_mask_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\update_mask_0/n1064 ), .force_10(
        \update_mask_0/n1065 ), .force_11(1'b0), .Q(o_mask[4]) );
  \**FFGEN**  \update_mask_0/o_mask_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\update_mask_0/n1068 ), .force_10(
        \update_mask_0/n1069 ), .force_11(1'b0), .Q(o_mask[3]) );
  \**FFGEN**  \update_mask_0/o_mask_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\update_mask_0/n1072 ), .force_10(
        \update_mask_0/n1073 ), .force_11(1'b0), .Q(o_mask[2]) );
  \**FFGEN**  \update_mask_0/o_mask_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\update_mask_0/n1076 ), .force_10(
        \update_mask_0/n1077 ), .force_11(1'b0), .Q(o_mask[1]) );
  \**FFGEN**  \update_mask_0/o_mask_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\update_mask_0/n948 ), .force_10(
        \update_mask_0/n949 ), .force_11(1'b0), .Q(o_mask[0]) );
  \**FFGEN**  \update_output_0/increment_reg  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1542 ), 
        .force_10(\update_output_0/n1543 ), .force_11(1'b0), .Q(
        \update_output_0/n2821 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[15][19]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1546 ), 
        .force_10(\update_output_0/n1547 ), .force_11(1'b0), .QN(n5816) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[15][18]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1550 ), 
        .force_10(\update_output_0/n1551 ), .force_11(1'b0), .QN(n5687) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[15][17]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1554 ), 
        .force_10(\update_output_0/n1555 ), .force_11(1'b0), .QN(n5783) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[15][16]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1558 ), 
        .force_10(\update_output_0/n1559 ), .force_11(1'b0), .QN(n5826) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[15][15]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1562 ), 
        .force_10(\update_output_0/n1563 ), .force_11(1'b0), .QN(n5689) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[15][14]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1566 ), 
        .force_10(\update_output_0/n1567 ), .force_11(1'b0), .QN(n5798) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[15][13]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1570 ), 
        .force_10(\update_output_0/n1571 ), .force_11(1'b0), .QN(n5832) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[15][12]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1574 ), 
        .force_10(\update_output_0/n1575 ), .force_11(1'b0), .QN(n5691) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[15][11]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1578 ), 
        .force_10(\update_output_0/n1579 ), .force_11(1'b0), .QN(n5803) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[15][10]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1582 ), 
        .force_10(\update_output_0/n1583 ), .force_11(1'b0), .QN(n5804) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[15][9]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1586 ), 
        .force_10(\update_output_0/n1587 ), .force_11(1'b0), .QN(n5693) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[15][8]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1590 ), 
        .force_10(\update_output_0/n1591 ), .force_11(1'b0), .QN(n5833) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[15][7]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1594 ), 
        .force_10(\update_output_0/n1595 ), .force_11(1'b0), .QN(n5884) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[15][6]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1598 ), 
        .force_10(\update_output_0/n1599 ), .force_11(1'b0), .QN(n5695) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[15][5]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1602 ), 
        .force_10(\update_output_0/n1603 ), .force_11(1'b0), .QN(n5827) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[15][4]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1606 ), 
        .force_10(\update_output_0/n1607 ), .force_11(1'b0), .QN(n5785) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[15][3]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1610 ), 
        .force_10(\update_output_0/n1611 ), .force_11(1'b0), .QN(n5697) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[15][2]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1614 ), 
        .force_10(\update_output_0/n1615 ), .force_11(1'b0), .QN(n5799) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[15][1]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1618 ), 
        .force_10(\update_output_0/n1619 ), .force_11(1'b0), .QN(n5797) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[15][0]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1622 ), 
        .force_10(\update_output_0/n1623 ), .force_11(1'b0), .QN(n5652) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[14][19]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1626 ), 
        .force_10(\update_output_0/n1627 ), .force_11(1'b0), .QN(n5886) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[14][18]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1630 ), 
        .force_10(\update_output_0/n1631 ), .force_11(1'b0), .QN(n5716) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[14][17]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1634 ), 
        .force_10(\update_output_0/n1635 ), .force_11(1'b0), .QN(n5862) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[14][16]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1638 ), 
        .force_10(\update_output_0/n1639 ), .force_11(1'b0), .QN(n5879) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[14][15]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1642 ), 
        .force_10(\update_output_0/n1643 ), .force_11(1'b0), .QN(n5722) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[14][14]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1646 ), 
        .force_10(\update_output_0/n1647 ), .force_11(1'b0), .QN(n5841) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[14][13]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1650 ), 
        .force_10(\update_output_0/n1651 ), .force_11(1'b0), .QN(n5885) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[14][12]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1654 ), 
        .force_10(\update_output_0/n1655 ), .force_11(1'b0), .QN(n5728) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[14][11]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1658 ), 
        .force_10(\update_output_0/n1659 ), .force_11(1'b0), .QN(n5868) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[14][10]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1662 ), 
        .force_10(\update_output_0/n1663 ), .force_11(1'b0), .QN(n5844) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[14][9]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1666 ), 
        .force_10(\update_output_0/n1667 ), .force_11(1'b0), .QN(n5732) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[14][8]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1670 ), 
        .force_10(\update_output_0/n1671 ), .force_11(1'b0), .QN(n5904) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[14][7]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1674 ), 
        .force_10(\update_output_0/n1675 ), .force_11(1'b0), .QN(n5847) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[14][6]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1678 ), 
        .force_10(\update_output_0/n1679 ), .force_11(1'b0), .QN(n5736) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[14][5]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1682 ), 
        .force_10(\update_output_0/n1683 ), .force_11(1'b0), .QN(n5902) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[14][4]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1686 ), 
        .force_10(\update_output_0/n1687 ), .force_11(1'b0), .QN(n5883) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[14][3]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1690 ), 
        .force_10(\update_output_0/n1691 ), .force_11(1'b0), .QN(n5740) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[14][2]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1694 ), 
        .force_10(\update_output_0/n1695 ), .force_11(1'b0), .QN(n5842) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[14][1]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1698 ), 
        .force_10(\update_output_0/n1699 ), .force_11(1'b0), .QN(n5882) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[14][0]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1702 ), 
        .force_10(\update_output_0/n1703 ), .force_11(1'b0), .QN(n5712) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[13][19]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1706 ), 
        .force_10(\update_output_0/n1707 ), .force_11(1'b0), .Q(
        \update_output_0/pre_o_im[13][19] ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[13][18]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1710 ), 
        .force_10(\update_output_0/n1711 ), .force_11(1'b0), .Q(
        \update_output_0/pre_o_im[13][18] ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[13][17]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1714 ), 
        .force_10(\update_output_0/n1715 ), .force_11(1'b0), .Q(
        \update_output_0/pre_o_im[13][17] ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[13][16]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1718 ), 
        .force_10(\update_output_0/n1719 ), .force_11(1'b0), .Q(
        \update_output_0/pre_o_im[13][16] ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[13][15]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1722 ), 
        .force_10(\update_output_0/n1723 ), .force_11(1'b0), .Q(
        \update_output_0/pre_o_im[13][15] ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[13][14]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1726 ), 
        .force_10(\update_output_0/n1727 ), .force_11(1'b0), .Q(
        \update_output_0/pre_o_im[13][14] ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[13][13]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1730 ), 
        .force_10(\update_output_0/n1731 ), .force_11(1'b0), .Q(
        \update_output_0/pre_o_im[13][13] ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[13][12]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1734 ), 
        .force_10(\update_output_0/n1735 ), .force_11(1'b0), .Q(
        \update_output_0/pre_o_im[13][12] ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[13][11]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1738 ), 
        .force_10(\update_output_0/n1739 ), .force_11(1'b0), .Q(
        \update_output_0/pre_o_im[13][11] ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[13][10]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1742 ), 
        .force_10(\update_output_0/n1743 ), .force_11(1'b0), .Q(
        \update_output_0/pre_o_im[13][10] ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[13][9]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1746 ), 
        .force_10(\update_output_0/n1747 ), .force_11(1'b0), .Q(
        \update_output_0/pre_o_im[13][9] ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[13][8]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1750 ), 
        .force_10(\update_output_0/n1751 ), .force_11(1'b0), .Q(
        \update_output_0/pre_o_im[13][8] ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[13][7]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1754 ), 
        .force_10(\update_output_0/n1755 ), .force_11(1'b0), .Q(
        \update_output_0/pre_o_im[13][7] ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[13][6]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1758 ), 
        .force_10(\update_output_0/n1759 ), .force_11(1'b0), .Q(
        \update_output_0/pre_o_im[13][6] ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[13][5]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1762 ), 
        .force_10(\update_output_0/n1763 ), .force_11(1'b0), .Q(
        \update_output_0/pre_o_im[13][5] ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[13][4]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1766 ), 
        .force_10(\update_output_0/n1767 ), .force_11(1'b0), .Q(
        \update_output_0/pre_o_im[13][4] ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[13][3]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1770 ), 
        .force_10(\update_output_0/n1771 ), .force_11(1'b0), .Q(
        \update_output_0/pre_o_im[13][3] ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[13][2]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1774 ), 
        .force_10(\update_output_0/n1775 ), .force_11(1'b0), .Q(
        \update_output_0/pre_o_im[13][2] ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[13][1]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1778 ), 
        .force_10(\update_output_0/n1779 ), .force_11(1'b0), .Q(
        \update_output_0/pre_o_im[13][1] ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[13][0]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1782 ), 
        .force_10(\update_output_0/n1783 ), .force_11(1'b0), .Q(
        \update_output_0/pre_o_im[13][0] ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[12][19]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1786 ), 
        .force_10(\update_output_0/n1787 ), .force_11(1'b0), .Q(
        \update_output_0/pre_o_im[12][19] ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[12][18]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1790 ), 
        .force_10(\update_output_0/n1791 ), .force_11(1'b0), .Q(
        \update_output_0/pre_o_im[12][18] ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[12][17]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1794 ), 
        .force_10(\update_output_0/n1795 ), .force_11(1'b0), .Q(
        \update_output_0/pre_o_im[12][17] ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[12][16]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1798 ), 
        .force_10(\update_output_0/n1799 ), .force_11(1'b0), .Q(
        \update_output_0/pre_o_im[12][16] ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[12][15]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1802 ), 
        .force_10(\update_output_0/n1803 ), .force_11(1'b0), .Q(
        \update_output_0/pre_o_im[12][15] ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[12][14]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1806 ), 
        .force_10(\update_output_0/n1807 ), .force_11(1'b0), .Q(
        \update_output_0/pre_o_im[12][14] ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[12][13]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1810 ), 
        .force_10(\update_output_0/n1811 ), .force_11(1'b0), .Q(
        \update_output_0/pre_o_im[12][13] ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[12][12]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1814 ), 
        .force_10(\update_output_0/n1815 ), .force_11(1'b0), .Q(
        \update_output_0/pre_o_im[12][12] ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[12][11]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1818 ), 
        .force_10(\update_output_0/n1819 ), .force_11(1'b0), .Q(
        \update_output_0/pre_o_im[12][11] ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[12][10]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1822 ), 
        .force_10(\update_output_0/n1823 ), .force_11(1'b0), .Q(
        \update_output_0/pre_o_im[12][10] ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[12][9]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1826 ), 
        .force_10(\update_output_0/n1827 ), .force_11(1'b0), .Q(
        \update_output_0/pre_o_im[12][9] ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[12][8]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1830 ), 
        .force_10(\update_output_0/n1831 ), .force_11(1'b0), .Q(
        \update_output_0/pre_o_im[12][8] ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[12][7]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1834 ), 
        .force_10(\update_output_0/n1835 ), .force_11(1'b0), .Q(
        \update_output_0/pre_o_im[12][7] ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[12][6]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1838 ), 
        .force_10(\update_output_0/n1839 ), .force_11(1'b0), .Q(
        \update_output_0/pre_o_im[12][6] ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[12][5]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1842 ), 
        .force_10(\update_output_0/n1843 ), .force_11(1'b0), .Q(
        \update_output_0/pre_o_im[12][5] ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[12][4]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1846 ), 
        .force_10(\update_output_0/n1847 ), .force_11(1'b0), .Q(
        \update_output_0/pre_o_im[12][4] ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[12][3]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1850 ), 
        .force_10(\update_output_0/n1851 ), .force_11(1'b0), .Q(
        \update_output_0/pre_o_im[12][3] ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[12][2]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1854 ), 
        .force_10(\update_output_0/n1855 ), .force_11(1'b0), .Q(
        \update_output_0/pre_o_im[12][2] ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[12][1]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1858 ), 
        .force_10(\update_output_0/n1859 ), .force_11(1'b0), .Q(
        \update_output_0/pre_o_im[12][1] ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[12][0]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1862 ), 
        .force_10(\update_output_0/n1863 ), .force_11(1'b0), .Q(
        \update_output_0/pre_o_im[12][0] ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[11][19]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1866 ), 
        .force_10(\update_output_0/n1867 ), .force_11(1'b0), .QN(n5686) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[11][18]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1870 ), 
        .force_10(\update_output_0/n1871 ), .force_11(1'b0), .QN(n5794) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[11][17]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1874 ), 
        .force_10(\update_output_0/n1875 ), .force_11(1'b0), .QN(n5769) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[11][16]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1878 ), 
        .force_10(\update_output_0/n1879 ), .force_11(1'b0), .QN(n5688) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[11][15]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1882 ), 
        .force_10(\update_output_0/n1883 ), .force_11(1'b0), .QN(n5786) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[11][14]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1886 ), 
        .force_10(\update_output_0/n1887 ), .force_11(1'b0), .QN(n5808) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[11][13]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1890 ), 
        .force_10(\update_output_0/n1891 ), .force_11(1'b0), .QN(n5690) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[11][12]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1894 ), 
        .force_10(\update_output_0/n1895 ), .force_11(1'b0), .QN(n5795) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[11][11]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1898 ), 
        .force_10(\update_output_0/n1899 ), .force_11(1'b0), .QN(n5812) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[11][10]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1902 ), 
        .force_10(\update_output_0/n1903 ), .force_11(1'b0), .QN(n5692) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[11][9]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1906 ), 
        .force_10(\update_output_0/n1907 ), .force_11(1'b0), .QN(n5876) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[11][8]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1910 ), 
        .force_10(\update_output_0/n1911 ), .force_11(1'b0), .QN(n5771) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[11][7]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1914 ), 
        .force_10(\update_output_0/n1915 ), .force_11(1'b0), .QN(n5694) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[11][6]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1918 ), 
        .force_10(\update_output_0/n1919 ), .force_11(1'b0), .QN(n5903) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[11][5]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1922 ), 
        .force_10(\update_output_0/n1923 ), .force_11(1'b0), .QN(n5777) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[11][4]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1926 ), 
        .force_10(\update_output_0/n1927 ), .force_11(1'b0), .QN(n5696) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[11][3]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1930 ), 
        .force_10(\update_output_0/n1931 ), .force_11(1'b0), .QN(n5873) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[11][2]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1934 ), 
        .force_10(\update_output_0/n1935 ), .force_11(1'b0), .QN(n5815) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[11][1]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1938 ), 
        .force_10(\update_output_0/n1939 ), .force_11(1'b0), .QN(n5698) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[11][0]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1942 ), 
        .force_10(\update_output_0/n1943 ), .force_11(1'b0), .QN(n5766) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[10][19]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1946 ), 
        .force_10(\update_output_0/n1947 ), .force_11(1'b0), .QN(n5714) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[10][18]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1950 ), 
        .force_10(\update_output_0/n1951 ), .force_11(1'b0), .QN(n5905) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[10][17]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1954 ), 
        .force_10(\update_output_0/n1955 ), .force_11(1'b0), .QN(n5821) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[10][16]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1958 ), 
        .force_10(\update_output_0/n1959 ), .force_11(1'b0), .QN(n5720) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[10][15]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1962 ), 
        .force_10(\update_output_0/n1963 ), .force_11(1'b0), .QN(n5875) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[10][14]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1966 ), 
        .force_10(\update_output_0/n1967 ), .force_11(1'b0), .QN(n5859) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[10][13]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1970 ), 
        .force_10(\update_output_0/n1971 ), .force_11(1'b0), .QN(n5726) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[10][12]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1974 ), 
        .force_10(\update_output_0/n1975 ), .force_11(1'b0), .QN(n5869) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[10][11]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1978 ), 
        .force_10(\update_output_0/n1979 ), .force_11(1'b0), .QN(n5867) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[10][10]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1982 ), 
        .force_10(\update_output_0/n1983 ), .force_11(1'b0), .QN(n5730) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[10][9]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1986 ), 
        .force_10(\update_output_0/n1987 ), .force_11(1'b0), .QN(n5857) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[10][8]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1990 ), 
        .force_10(\update_output_0/n1991 ), .force_11(1'b0), .QN(n5890) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[10][7]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1994 ), 
        .force_10(\update_output_0/n1995 ), .force_11(1'b0), .QN(n5734) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[10][6]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1998 ), 
        .force_10(\update_output_0/n1999 ), .force_11(1'b0), .QN(n5852) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[10][5]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2002 ), 
        .force_10(\update_output_0/n2003 ), .force_11(1'b0), .QN(n5865) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[10][4]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2006 ), 
        .force_10(\update_output_0/n2007 ), .force_11(1'b0), .QN(n5738) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[10][3]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2010 ), 
        .force_10(\update_output_0/n2011 ), .force_11(1'b0), .QN(n5901) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[10][2]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2014 ), 
        .force_10(\update_output_0/n2015 ), .force_11(1'b0), .QN(n5881) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[10][1]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2018 ), 
        .force_10(\update_output_0/n2019 ), .force_11(1'b0), .QN(n5742) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[10][0]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2022 ), 
        .force_10(\update_output_0/n2023 ), .force_11(1'b0), .QN(n5851) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[9][19]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2026 ), 
        .force_10(\update_output_0/n2027 ), .force_11(1'b0), .QN(n5791) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[9][18]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2030 ), 
        .force_10(\update_output_0/n2031 ), .force_11(1'b0), .QN(n5781) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[9][17]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2034 ), 
        .force_10(\update_output_0/n2035 ), .force_11(1'b0), .QN(n5657) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[9][16]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2038 ), 
        .force_10(\update_output_0/n2039 ), .force_11(1'b0), .QN(n5802) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[9][15]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2042 ), 
        .force_10(\update_output_0/n2043 ), .force_11(1'b0), .QN(n5871) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[9][14]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2046 ), 
        .force_10(\update_output_0/n2047 ), .force_11(1'b0), .QN(n5662) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[9][13]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2050 ), 
        .force_10(\update_output_0/n2051 ), .force_11(1'b0), .QN(n5824) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[9][12]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2054 ), 
        .force_10(\update_output_0/n2055 ), .force_11(1'b0), .QN(n5776) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[9][11]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2058 ), 
        .force_10(\update_output_0/n2059 ), .force_11(1'b0), .QN(n5667) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[9][10]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2062 ), 
        .force_10(\update_output_0/n2063 ), .force_11(1'b0), .QN(n5834) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[9][9]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2066 ), 
        .force_10(\update_output_0/n2067 ), .force_11(1'b0), .QN(n5805) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[9][8]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2070 ), 
        .force_10(\update_output_0/n2071 ), .force_11(1'b0), .QN(n5672) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[9][7]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2074 ), 
        .force_10(\update_output_0/n2075 ), .force_11(1'b0), .QN(n5779) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[9][6]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2078 ), 
        .force_10(\update_output_0/n2079 ), .force_11(1'b0), .QN(n5792) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[9][5]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2082 ), 
        .force_10(\update_output_0/n2083 ), .force_11(1'b0), .QN(n5677) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[9][4]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2086 ), 
        .force_10(\update_output_0/n2087 ), .force_11(1'b0), .QN(n5835) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[9][3]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2090 ), 
        .force_10(\update_output_0/n2091 ), .force_11(1'b0), .QN(n5817) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[9][2]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2094 ), 
        .force_10(\update_output_0/n2095 ), .force_11(1'b0), .QN(n5682) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[9][1]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2098 ), 
        .force_10(\update_output_0/n2099 ), .force_11(1'b0), .QN(n5811) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[9][0]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2102 ), 
        .force_10(\update_output_0/n2103 ), .force_11(1'b0), .QN(n5910) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[8][19]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2106 ), 
        .force_10(\update_output_0/n2107 ), .force_11(1'b0), .QN(n5897) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[8][18]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2110 ), 
        .force_10(\update_output_0/n2111 ), .force_11(1'b0), .QN(n5863) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[8][17]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2114 ), 
        .force_10(\update_output_0/n2115 ), .force_11(1'b0), .QN(n5717) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[8][16]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2118 ), 
        .force_10(\update_output_0/n2119 ), .force_11(1'b0), .QN(n5894) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[8][15]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2122 ), 
        .force_10(\update_output_0/n2123 ), .force_11(1'b0), .QN(n5908) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[8][14]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2126 ), 
        .force_10(\update_output_0/n2127 ), .force_11(1'b0), .QN(n5723) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[8][13]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2130 ), 
        .force_10(\update_output_0/n2131 ), .force_11(1'b0), .QN(n5866) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[8][12]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2134 ), 
        .force_10(\update_output_0/n2135 ), .force_11(1'b0), .QN(n5907) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[8][11]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2138 ), 
        .force_10(\update_output_0/n2139 ), .force_11(1'b0), .QN(n5729) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[8][10]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2142 ), 
        .force_10(\update_output_0/n2143 ), .force_11(1'b0), .QN(n5843) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[8][9]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2146 ), 
        .force_10(\update_output_0/n2147 ), .force_11(1'b0), .QN(n5906) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[8][8]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2150 ), 
        .force_10(\update_output_0/n2151 ), .force_11(1'b0), .QN(n5733) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[8][7]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2154 ), 
        .force_10(\update_output_0/n2155 ), .force_11(1'b0), .QN(n5818) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[8][6]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2158 ), 
        .force_10(\update_output_0/n2159 ), .force_11(1'b0), .QN(n5846) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[8][5]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2162 ), 
        .force_10(\update_output_0/n2163 ), .force_11(1'b0), .QN(n5737) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[8][4]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2166 ), 
        .force_10(\update_output_0/n2167 ), .force_11(1'b0), .QN(n5820) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[8][3]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2170 ), 
        .force_10(\update_output_0/n2171 ), .force_11(1'b0), .QN(n5861) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[8][2]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2174 ), 
        .force_10(\update_output_0/n2175 ), .force_11(1'b0), .QN(n5741) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[8][1]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2178 ), 
        .force_10(\update_output_0/n2179 ), .force_11(1'b0), .QN(n5836) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[8][0]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2182 ), 
        .force_10(\update_output_0/n2183 ), .force_11(1'b0), .QN(n5711) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[7][19]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2186 ), 
        .force_10(\update_output_0/n2187 ), .force_11(1'b0), .QN(n5654) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[7][18]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2190 ), 
        .force_10(\update_output_0/n2191 ), .force_11(1'b0), .QN(n5774) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[7][17]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2194 ), 
        .force_10(\update_output_0/n2195 ), .force_11(1'b0), .QN(n5700) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[7][16]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2198 ), 
        .force_10(\update_output_0/n2199 ), .force_11(1'b0), .QN(n5659) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[7][15]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2202 ), 
        .force_10(\update_output_0/n2203 ), .force_11(1'b0), .QN(n5829) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[7][14]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2206 ), 
        .force_10(\update_output_0/n2207 ), .force_11(1'b0), .QN(n5702) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[7][13]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2210 ), 
        .force_10(\update_output_0/n2211 ), .force_11(1'b0), .QN(n5664) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[7][12]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2214 ), 
        .force_10(\update_output_0/n2215 ), .force_11(1'b0), .QN(n5767) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[7][11]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2218 ), 
        .force_10(\update_output_0/n2219 ), .force_11(1'b0), .QN(n5704) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[7][10]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2222 ), 
        .force_10(\update_output_0/n2223 ), .force_11(1'b0), .QN(n5669) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[7][9]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2226 ), 
        .force_10(\update_output_0/n2227 ), .force_11(1'b0), .QN(n5788) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[7][8]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2230 ), 
        .force_10(\update_output_0/n2231 ), .force_11(1'b0), .QN(n5706) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[7][7]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2234 ), 
        .force_10(\update_output_0/n2235 ), .force_11(1'b0), .QN(n5674) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[7][6]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2238 ), 
        .force_10(\update_output_0/n2239 ), .force_11(1'b0), .QN(n5828) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[7][5]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2242 ), 
        .force_10(\update_output_0/n2243 ), .force_11(1'b0), .QN(n5708) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[7][4]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2246 ), 
        .force_10(\update_output_0/n2247 ), .force_11(1'b0), .QN(n5679) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[7][3]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2250 ), 
        .force_10(\update_output_0/n2251 ), .force_11(1'b0), .QN(n5801) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[7][2]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2254 ), 
        .force_10(\update_output_0/n2255 ), .force_11(1'b0), .QN(n5710) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[7][1]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2258 ), 
        .force_10(\update_output_0/n2259 ), .force_11(1'b0), .QN(n5684) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[7][0]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2262 ), 
        .force_10(\update_output_0/n2263 ), .force_11(1'b0), .QN(n5772) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[6][19]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2266 ), 
        .force_10(\update_output_0/n2267 ), .force_11(1'b0), .QN(n5715) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[6][18]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2270 ), 
        .force_10(\update_output_0/n2271 ), .force_11(1'b0), .QN(n5896) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[6][17]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2274 ), 
        .force_10(\update_output_0/n2275 ), .force_11(1'b0), .QN(n5719) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[6][16]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2278 ), 
        .force_10(\update_output_0/n2279 ), .force_11(1'b0), .QN(n5721) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[6][15]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2282 ), 
        .force_10(\update_output_0/n2283 ), .force_11(1'b0), .QN(n5860) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[6][14]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2286 ), 
        .force_10(\update_output_0/n2287 ), .force_11(1'b0), .QN(n5725) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[6][13]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2290 ), 
        .force_10(\update_output_0/n2291 ), .force_11(1'b0), .QN(n5727) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[6][12]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2294 ), 
        .force_10(\update_output_0/n2295 ), .force_11(1'b0), .QN(n5839) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[6][11]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2298 ), 
        .force_10(\update_output_0/n2299 ), .force_11(1'b0), .QN(n5751) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[6][10]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2302 ), 
        .force_10(\update_output_0/n2303 ), .force_11(1'b0), .QN(n5731) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[6][9]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2306 ), 
        .force_10(\update_output_0/n2307 ), .force_11(1'b0), .QN(n5840) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[6][8]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2310 ), 
        .force_10(\update_output_0/n2311 ), .force_11(1'b0), .QN(n5755) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[6][7]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2314 ), 
        .force_10(\update_output_0/n2315 ), .force_11(1'b0), .QN(n5735) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[6][6]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2318 ), 
        .force_10(\update_output_0/n2319 ), .force_11(1'b0), .QN(n5845) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[6][5]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2322 ), 
        .force_10(\update_output_0/n2323 ), .force_11(1'b0), .QN(n5759) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[6][4]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2326 ), 
        .force_10(\update_output_0/n2327 ), .force_11(1'b0), .QN(n5739) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[6][3]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2330 ), 
        .force_10(\update_output_0/n2331 ), .force_11(1'b0), .QN(n5887) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[6][2]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2334 ), 
        .force_10(\update_output_0/n2335 ), .force_11(1'b0), .QN(n5763) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[6][1]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2338 ), 
        .force_10(\update_output_0/n2339 ), .force_11(1'b0), .QN(n5743) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[6][0]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2342 ), 
        .force_10(\update_output_0/n2343 ), .force_11(1'b0), .QN(n5909) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[5][19]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2346 ), 
        .force_10(\update_output_0/n2347 ), .force_11(1'b0), .QN(n5814) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[5][18]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2350 ), 
        .force_10(\update_output_0/n2351 ), .force_11(1'b0), .QN(n5656) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[5][17]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2354 ), 
        .force_10(\update_output_0/n2355 ), .force_11(1'b0), .QN(n5895) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[5][16]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2358 ), 
        .force_10(\update_output_0/n2359 ), .force_11(1'b0), .QN(n5809) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[5][15]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2362 ), 
        .force_10(\update_output_0/n2363 ), .force_11(1'b0), .QN(n5661) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[5][14]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2366 ), 
        .force_10(\update_output_0/n2367 ), .force_11(1'b0), .QN(n5806) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[5][13]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2370 ), 
        .force_10(\update_output_0/n2371 ), .force_11(1'b0), .QN(n5898) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[5][12]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2374 ), 
        .force_10(\update_output_0/n2375 ), .force_11(1'b0), .QN(n5666) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[5][11]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2378 ), 
        .force_10(\update_output_0/n2379 ), .force_11(1'b0), .QN(n5892) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[5][10]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2382 ), 
        .force_10(\update_output_0/n2383 ), .force_11(1'b0), .QN(n5800) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[5][9]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2386 ), 
        .force_10(\update_output_0/n2387 ), .force_11(1'b0), .QN(n5671) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[5][8]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2390 ), 
        .force_10(\update_output_0/n2391 ), .force_11(1'b0), .QN(n5793) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[5][7]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2394 ), 
        .force_10(\update_output_0/n2395 ), .force_11(1'b0), .QN(n5787) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[5][6]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2398 ), 
        .force_10(\update_output_0/n2399 ), .force_11(1'b0), .QN(n5676) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[5][5]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2402 ), 
        .force_10(\update_output_0/n2403 ), .force_11(1'b0), .QN(n5790) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[5][4]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2406 ), 
        .force_10(\update_output_0/n2407 ), .force_11(1'b0), .QN(n5782) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[5][3]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2410 ), 
        .force_10(\update_output_0/n2411 ), .force_11(1'b0), .QN(n5681) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[5][2]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2414 ), 
        .force_10(\update_output_0/n2415 ), .force_11(1'b0), .QN(n5780) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[5][1]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2418 ), 
        .force_10(\update_output_0/n2419 ), .force_11(1'b0), .QN(n5789) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[5][0]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2422 ), 
        .force_10(\update_output_0/n2423 ), .force_11(1'b0), .QN(n5651) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[4][19]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2426 ), 
        .force_10(\update_output_0/n2427 ), .force_11(1'b0), .Q(
        \update_output_0/pre_o_im[4][19] ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[4][18]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2430 ), 
        .force_10(\update_output_0/n2431 ), .force_11(1'b0), .Q(
        \update_output_0/pre_o_im[4][18] ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[4][17]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2434 ), 
        .force_10(\update_output_0/n2435 ), .force_11(1'b0), .Q(
        \update_output_0/pre_o_im[4][17] ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[4][16]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2438 ), 
        .force_10(\update_output_0/n2439 ), .force_11(1'b0), .Q(
        \update_output_0/pre_o_im[4][16] ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[4][15]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2442 ), 
        .force_10(\update_output_0/n2443 ), .force_11(1'b0), .Q(
        \update_output_0/pre_o_im[4][15] ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[4][14]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2446 ), 
        .force_10(\update_output_0/n2447 ), .force_11(1'b0), .Q(
        \update_output_0/pre_o_im[4][14] ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[4][13]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2450 ), 
        .force_10(\update_output_0/n2451 ), .force_11(1'b0), .Q(
        \update_output_0/pre_o_im[4][13] ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[4][12]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2454 ), 
        .force_10(\update_output_0/n2455 ), .force_11(1'b0), .Q(
        \update_output_0/pre_o_im[4][12] ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[4][11]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2458 ), 
        .force_10(\update_output_0/n2459 ), .force_11(1'b0), .Q(
        \update_output_0/pre_o_im[4][11] ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[4][10]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2462 ), 
        .force_10(\update_output_0/n2463 ), .force_11(1'b0), .Q(
        \update_output_0/pre_o_im[4][10] ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[4][9]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2466 ), 
        .force_10(\update_output_0/n2467 ), .force_11(1'b0), .Q(
        \update_output_0/pre_o_im[4][9] ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[4][8]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2470 ), 
        .force_10(\update_output_0/n2471 ), .force_11(1'b0), .Q(
        \update_output_0/pre_o_im[4][8] ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[4][7]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2474 ), 
        .force_10(\update_output_0/n2475 ), .force_11(1'b0), .Q(
        \update_output_0/pre_o_im[4][7] ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[4][6]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2478 ), 
        .force_10(\update_output_0/n2479 ), .force_11(1'b0), .Q(
        \update_output_0/pre_o_im[4][6] ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[4][5]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2482 ), 
        .force_10(\update_output_0/n2483 ), .force_11(1'b0), .Q(
        \update_output_0/pre_o_im[4][5] ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[4][4]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2486 ), 
        .force_10(\update_output_0/n2487 ), .force_11(1'b0), .Q(
        \update_output_0/pre_o_im[4][4] ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[4][3]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2490 ), 
        .force_10(\update_output_0/n2491 ), .force_11(1'b0), .Q(
        \update_output_0/pre_o_im[4][3] ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[4][2]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2494 ), 
        .force_10(\update_output_0/n2495 ), .force_11(1'b0), .Q(
        \update_output_0/pre_o_im[4][2] ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[4][1]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2498 ), 
        .force_10(\update_output_0/n2499 ), .force_11(1'b0), .Q(
        \update_output_0/pre_o_im[4][1] ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[4][0]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2502 ), 
        .force_10(\update_output_0/n2503 ), .force_11(1'b0), .Q(
        \update_output_0/pre_o_im[4][0] ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[3][19]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2506 ), 
        .force_10(\update_output_0/n2507 ), .force_11(1'b0), .QN(n5773) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[3][18]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2510 ), 
        .force_10(\update_output_0/n2511 ), .force_11(1'b0), .QN(n5699) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[3][17]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2514 ), 
        .force_10(\update_output_0/n2515 ), .force_11(1'b0), .QN(n5658) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[3][16]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2518 ), 
        .force_10(\update_output_0/n2519 ), .force_11(1'b0), .QN(n5870) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[3][15]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2522 ), 
        .force_10(\update_output_0/n2523 ), .force_11(1'b0), .QN(n5701) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[3][14]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2526 ), 
        .force_10(\update_output_0/n2527 ), .force_11(1'b0), .QN(n5663) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[3][13]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2530 ), 
        .force_10(\update_output_0/n2531 ), .force_11(1'b0), .QN(n5784) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[3][12]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2534 ), 
        .force_10(\update_output_0/n2535 ), .force_11(1'b0), .QN(n5703) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[3][11]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2538 ), 
        .force_10(\update_output_0/n2539 ), .force_11(1'b0), .QN(n5668) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[3][10]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2542 ), 
        .force_10(\update_output_0/n2543 ), .force_11(1'b0), .QN(n5775) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[3][9]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2546 ), 
        .force_10(\update_output_0/n2547 ), .force_11(1'b0), .QN(n5705) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[3][8]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2550 ), 
        .force_10(\update_output_0/n2551 ), .force_11(1'b0), .QN(n5673) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[3][7]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2554 ), 
        .force_10(\update_output_0/n2555 ), .force_11(1'b0), .QN(n5810) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[3][6]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2558 ), 
        .force_10(\update_output_0/n2559 ), .force_11(1'b0), .QN(n5707) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[3][5]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2562 ), 
        .force_10(\update_output_0/n2563 ), .force_11(1'b0), .QN(n5678) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[3][4]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2566 ), 
        .force_10(\update_output_0/n2567 ), .force_11(1'b0), .QN(n5888) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[3][3]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2570 ), 
        .force_10(\update_output_0/n2571 ), .force_11(1'b0), .QN(n5709) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[3][2]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2574 ), 
        .force_10(\update_output_0/n2575 ), .force_11(1'b0), .QN(n5683) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[3][1]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2578 ), 
        .force_10(\update_output_0/n2579 ), .force_11(1'b0), .QN(n5823) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[3][0]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2582 ), 
        .force_10(\update_output_0/n2583 ), .force_11(1'b0), .QN(n5653) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[2][19]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2586 ), 
        .force_10(\update_output_0/n2587 ), .force_11(1'b0), .QN(n5849) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[2][18]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2590 ), 
        .force_10(\update_output_0/n2591 ), .force_11(1'b0), .QN(n5745) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[2][17]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2594 ), 
        .force_10(\update_output_0/n2595 ), .force_11(1'b0), .QN(n5718) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[2][16]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2598 ), 
        .force_10(\update_output_0/n2599 ), .force_11(1'b0), .QN(n5878) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[2][15]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2602 ), 
        .force_10(\update_output_0/n2603 ), .force_11(1'b0), .QN(n5747) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[2][14]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2606 ), 
        .force_10(\update_output_0/n2607 ), .force_11(1'b0), .QN(n5724) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[2][13]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2610 ), 
        .force_10(\update_output_0/n2611 ), .force_11(1'b0), .QN(n5837) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[2][12]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2614 ), 
        .force_10(\update_output_0/n2615 ), .force_11(1'b0), .QN(n5749) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[2][11]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2618 ), 
        .force_10(\update_output_0/n2619 ), .force_11(1'b0), .QN(n5750) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[2][10]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2622 ), 
        .force_10(\update_output_0/n2623 ), .force_11(1'b0), .QN(n5891) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[2][9]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2626 ), 
        .force_10(\update_output_0/n2627 ), .force_11(1'b0), .QN(n5753) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[2][8]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2630 ), 
        .force_10(\update_output_0/n2631 ), .force_11(1'b0), .QN(n5754) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[2][7]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2634 ), 
        .force_10(\update_output_0/n2635 ), .force_11(1'b0), .QN(n5858) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[2][6]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2638 ), 
        .force_10(\update_output_0/n2639 ), .force_11(1'b0), .QN(n5757) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[2][5]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2642 ), 
        .force_10(\update_output_0/n2643 ), .force_11(1'b0), .QN(n5758) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[2][4]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2646 ), 
        .force_10(\update_output_0/n2647 ), .force_11(1'b0), .QN(n5854) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[2][3]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2650 ), 
        .force_10(\update_output_0/n2651 ), .force_11(1'b0), .QN(n5761) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[2][2]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2654 ), 
        .force_10(\update_output_0/n2655 ), .force_11(1'b0), .QN(n5762) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[2][1]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2658 ), 
        .force_10(\update_output_0/n2659 ), .force_11(1'b0), .QN(n5880) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[2][0]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2662 ), 
        .force_10(\update_output_0/n2663 ), .force_11(1'b0), .QN(n5713) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[1][19]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2666 ), 
        .force_10(\update_output_0/n2667 ), .force_11(1'b0), .QN(n5655) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[1][18]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2670 ), 
        .force_10(\update_output_0/n2671 ), .force_11(1'b0), .QN(n5872) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[1][17]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2674 ), 
        .force_10(\update_output_0/n2675 ), .force_11(1'b0), .QN(n5899) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[1][16]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2678 ), 
        .force_10(\update_output_0/n2679 ), .force_11(1'b0), .QN(n5660) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[1][15]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2682 ), 
        .force_10(\update_output_0/n2683 ), .force_11(1'b0), .QN(n5770) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[1][14]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2686 ), 
        .force_10(\update_output_0/n2687 ), .force_11(1'b0), .QN(n5765) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[1][13]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2690 ), 
        .force_10(\update_output_0/n2691 ), .force_11(1'b0), .QN(n5665) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[1][12]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2694 ), 
        .force_10(\update_output_0/n2695 ), .force_11(1'b0), .QN(n5825) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[1][11]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2698 ), 
        .force_10(\update_output_0/n2699 ), .force_11(1'b0), .QN(n5778) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[1][10]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2702 ), 
        .force_10(\update_output_0/n2703 ), .force_11(1'b0), .QN(n5670) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[1][9]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2706 ), 
        .force_10(\update_output_0/n2707 ), .force_11(1'b0), .QN(n5807) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[1][8]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2710 ), 
        .force_10(\update_output_0/n2711 ), .force_11(1'b0), .QN(n5796) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[1][7]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2714 ), 
        .force_10(\update_output_0/n2715 ), .force_11(1'b0), .QN(n5675) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[1][6]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2718 ), 
        .force_10(\update_output_0/n2719 ), .force_11(1'b0), .QN(n5889) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[1][5]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2722 ), 
        .force_10(\update_output_0/n2723 ), .force_11(1'b0), .QN(n5830) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[1][4]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2726 ), 
        .force_10(\update_output_0/n2727 ), .force_11(1'b0), .QN(n5680) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[1][3]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2730 ), 
        .force_10(\update_output_0/n2731 ), .force_11(1'b0), .QN(n5768) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[1][2]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2734 ), 
        .force_10(\update_output_0/n2735 ), .force_11(1'b0), .QN(n5813) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[1][1]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2738 ), 
        .force_10(\update_output_0/n2739 ), .force_11(1'b0), .QN(n5685) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[1][0]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2742 ), 
        .force_10(\update_output_0/n2743 ), .force_11(1'b0), .QN(n5831) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[0][19]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2746 ), 
        .force_10(\update_output_0/n2747 ), .force_11(1'b0), .QN(n5744) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[0][18]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2750 ), 
        .force_10(\update_output_0/n2751 ), .force_11(1'b0), .QN(n5819) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[0][17]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2754 ), 
        .force_10(\update_output_0/n2755 ), .force_11(1'b0), .QN(n5900) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[0][16]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2758 ), 
        .force_10(\update_output_0/n2759 ), .force_11(1'b0), .QN(n5746) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[0][15]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2762 ), 
        .force_10(\update_output_0/n2763 ), .force_11(1'b0), .QN(n5893) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[0][14]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2766 ), 
        .force_10(\update_output_0/n2767 ), .force_11(1'b0), .QN(n5850) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[0][13]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2770 ), 
        .force_10(\update_output_0/n2771 ), .force_11(1'b0), .QN(n5748) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[0][12]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2774 ), 
        .force_10(\update_output_0/n2775 ), .force_11(1'b0), .QN(n5848) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[0][11]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2778 ), 
        .force_10(\update_output_0/n2779 ), .force_11(1'b0), .QN(n5855) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[0][10]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2782 ), 
        .force_10(\update_output_0/n2783 ), .force_11(1'b0), .QN(n5752) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[0][9]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2786 ), 
        .force_10(\update_output_0/n2787 ), .force_11(1'b0), .QN(n5856) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[0][8]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2790 ), 
        .force_10(\update_output_0/n2791 ), .force_11(1'b0), .QN(n5838) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[0][7]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2794 ), 
        .force_10(\update_output_0/n2795 ), .force_11(1'b0), .QN(n5756) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[0][6]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2798 ), 
        .force_10(\update_output_0/n2799 ), .force_11(1'b0), .QN(n5877) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[0][5]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2802 ), 
        .force_10(\update_output_0/n2803 ), .force_11(1'b0), .QN(n5864) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[0][4]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2806 ), 
        .force_10(\update_output_0/n2807 ), .force_11(1'b0), .QN(n5760) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[0][3]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2810 ), 
        .force_10(\update_output_0/n2811 ), .force_11(1'b0), .QN(n5874) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[0][2]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2814 ), 
        .force_10(\update_output_0/n2815 ), .force_11(1'b0), .QN(n5853) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[0][1]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2818 ), 
        .force_10(\update_output_0/n2819 ), .force_11(1'b0), .QN(n5764) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[0][0]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n1538 ), 
        .force_10(\update_output_0/n1539 ), .force_11(1'b0), .QN(n5822) );
  nor_x2_sg U3975 ( .A(n1503), .B(n1504), .X(n1502) );
  nand_x4_sg U7051 ( .A(n1505), .B(n1506), .X(n1504) );
  nand_x4_sg U7052 ( .A(n1849), .B(n1850), .X(n1503) );
  nand_x1_sg U7053 ( .A(n1513), .B(n1514), .X(n1512) );
  nand_x1_sg U7054 ( .A(n1857), .B(n1858), .X(n1856) );
  nand_x1_sg U7055 ( .A(n7268), .B(n9193), .X(n1048) );
  inv_x2_sg U7056 ( .A(\i_im[14][11] ), .X(n9193) );
  nand_x1_sg U7057 ( .A(n1687), .B(n1688), .X(n1686) );
  nand_x1_sg U7058 ( .A(n1602), .B(n1603), .X(n1601) );
  nand_x1_sg U7059 ( .A(n1770), .B(n1771), .X(n1769) );
  nand_x1_sg U7060 ( .A(n2025), .B(n2026), .X(n2024) );
  nand_x1_sg U7061 ( .A(n1940), .B(n1941), .X(n1939) );
  nand_x1_sg U7062 ( .A(n2108), .B(n2109), .X(n2107) );
  nand_x1_sg U7063 ( .A(n7264), .B(n9194), .X(n984) );
  inv_x2_sg U7064 ( .A(\i_im[14][12] ), .X(n9194) );
  nand_x1_sg U7065 ( .A(n7270), .B(n9192), .X(n1016) );
  inv_x2_sg U7066 ( .A(\i_im[14][10] ), .X(n9192) );
  nand_x1_sg U7067 ( .A(n1048), .B(n9133), .X(n1045) );
  nand_x1_sg U7068 ( .A(n949), .B(n9141), .X(n946) );
  nand_x1_sg U7069 ( .A(n7269), .B(n9201), .X(n949) );
  inv_x2_sg U7070 ( .A(\i_im[14][19] ), .X(n9201) );
  nor_x1_sg U7071 ( .A(n1681), .B(n1682), .X(n1505) );
  nor_x1_sg U7072 ( .A(n1507), .B(n1508), .X(n1506) );
  nor_x1_sg U7073 ( .A(n2019), .B(n2020), .X(n1849) );
  nor_x1_sg U7074 ( .A(n1851), .B(n1852), .X(n1850) );
  nand_x1_sg U7075 ( .A(n984), .B(n9134), .X(n981) );
  nand_x1_sg U7076 ( .A(n1410), .B(n1411), .X(n755) );
  nand_x1_sg U7077 ( .A(n1412), .B(n1413), .X(n1411) );
  nand_x1_sg U7078 ( .A(n1215), .B(n1216), .X(n737) );
  nand_x1_sg U7079 ( .A(n1183), .B(n1184), .X(n738) );
  nand_x1_sg U7080 ( .A(n1200), .B(n1201), .X(n1183) );
  nand_x1_sg U7081 ( .A(n1314), .B(n1315), .X(n741) );
  nand_x1_sg U7082 ( .A(n1346), .B(n1347), .X(n742) );
  nand_x1_sg U7083 ( .A(n1363), .B(n1364), .X(n1346) );
  nand_x1_sg U7084 ( .A(n1016), .B(n9132), .X(n1013) );
  nand_x1_sg U7085 ( .A(n1018), .B(n1019), .X(n745) );
  nand_x1_sg U7086 ( .A(n1050), .B(n1051), .X(n747) );
  nand_x1_sg U7087 ( .A(n1052), .B(n1053), .X(n1051) );
  nand_x1_sg U7088 ( .A(n1082), .B(n1083), .X(n748) );
  nand_x1_sg U7089 ( .A(n1099), .B(n1100), .X(n1082) );
  nand_x1_sg U7090 ( .A(n855), .B(n856), .X(n751) );
  nand_x1_sg U7091 ( .A(n857), .B(n858), .X(n856) );
  nand_x1_sg U7092 ( .A(n887), .B(n888), .X(n752) );
  nand_x1_sg U7093 ( .A(n889), .B(n890), .X(n888) );
  nand_x1_sg U7094 ( .A(n919), .B(n920), .X(n753) );
  nand_x1_sg U7095 ( .A(n936), .B(n937), .X(n919) );
  nand_x1_sg U7096 ( .A(n1378), .B(n1379), .X(n743) );
  nand_x1_sg U7097 ( .A(n1250), .B(n1251), .X(n739) );
  nand_x1_sg U7098 ( .A(n1282), .B(n1283), .X(n740) );
  nand_x1_sg U7099 ( .A(n6830), .B(n3695), .X(n3656) );
  nand_x1_sg U7100 ( .A(n8959), .B(n1772), .X(n1771) );
  nand_x1_sg U7101 ( .A(n7438), .B(n1536), .X(n1513) );
  nand_x1_sg U7102 ( .A(n7437), .B(n1515), .X(n1514) );
  nand_x1_sg U7103 ( .A(n1674), .B(n1675), .X(n1666) );
  nand_x1_sg U7104 ( .A(n7436), .B(n1619), .X(n1602) );
  nand_x1_sg U7105 ( .A(n7435), .B(n1604), .X(n1603) );
  nand_x1_sg U7106 ( .A(n7434), .B(n1704), .X(n1687) );
  nand_x1_sg U7107 ( .A(n7433), .B(n1689), .X(n1688) );
  nand_x1_sg U7108 ( .A(n8960), .B(n2110), .X(n2109) );
  nand_x1_sg U7109 ( .A(n7429), .B(n1874), .X(n1857) );
  nand_x1_sg U7110 ( .A(n7432), .B(n1859), .X(n1858) );
  nand_x1_sg U7111 ( .A(n2012), .B(n2013), .X(n2004) );
  nand_x1_sg U7112 ( .A(n7427), .B(n1957), .X(n1940) );
  nand_x1_sg U7113 ( .A(n7430), .B(n1942), .X(n1941) );
  nand_x1_sg U7114 ( .A(n7425), .B(n2042), .X(n2025) );
  nand_x1_sg U7115 ( .A(n7428), .B(n2027), .X(n2026) );
  nand_x1_sg U7116 ( .A(n7431), .B(n1787), .X(n1770) );
  nor_x1_sg U7117 ( .A(n1834), .B(n1835), .X(n1817) );
  nor_x1_sg U7118 ( .A(n1819), .B(n1820), .X(n1818) );
  nand_x1_sg U7119 ( .A(n1842), .B(n1843), .X(n1834) );
  nand_x2_sg U7120 ( .A(n1509), .B(n1510), .X(n1508) );
  nor_x1_sg U7121 ( .A(n1583), .B(n1584), .X(n1566) );
  nand_x2_sg U7122 ( .A(n1598), .B(n1599), .X(n1507) );
  nor_x1_sg U7123 ( .A(n1666), .B(n1667), .X(n1649) );
  nand_x2_sg U7124 ( .A(n1683), .B(n1684), .X(n1682) );
  nor_x1_sg U7125 ( .A(n1751), .B(n1752), .X(n1734) );
  nand_x1_sg U7126 ( .A(n7426), .B(n2125), .X(n2108) );
  nor_x1_sg U7127 ( .A(n2172), .B(n2173), .X(n2155) );
  nor_x1_sg U7128 ( .A(n2157), .B(n2158), .X(n2156) );
  nand_x1_sg U7129 ( .A(n2181), .B(n2182), .X(n2172) );
  nand_x2_sg U7130 ( .A(n1853), .B(n1854), .X(n1852) );
  nor_x1_sg U7131 ( .A(n1921), .B(n1922), .X(n1904) );
  nand_x2_sg U7132 ( .A(n1936), .B(n1937), .X(n1851) );
  nor_x1_sg U7133 ( .A(n2004), .B(n2005), .X(n1987) );
  nand_x2_sg U7134 ( .A(n2021), .B(n2022), .X(n2020) );
  nor_x1_sg U7135 ( .A(n2089), .B(n2090), .X(n2072) );
  nand_x1_sg U7136 ( .A(n9021), .B(n934), .X(n930) );
  nand_x2_sg U7137 ( .A(n1766), .B(n1767), .X(n1681) );
  nand_x2_sg U7138 ( .A(n2104), .B(n2105), .X(n2019) );
  nand_x2_sg U7139 ( .A(n5980), .B(n5814), .X(n4848) );
  nand_x2_sg U7140 ( .A(n6894), .B(n5895), .X(n4774) );
  nand_x2_sg U7141 ( .A(n6895), .B(n5809), .X(n4738) );
  nand_x2_sg U7142 ( .A(n6893), .B(n5806), .X(n4666) );
  nand_x2_sg U7143 ( .A(n6894), .B(n5898), .X(n4630) );
  nand_x2_sg U7144 ( .A(n6896), .B(n5666), .X(n4594) );
  nand_x2_sg U7145 ( .A(n6895), .B(n5892), .X(n4558) );
  nand_x2_sg U7146 ( .A(n6895), .B(n5800), .X(n4522) );
  nand_x2_sg U7147 ( .A(n6894), .B(n5793), .X(n4450) );
  nand_x2_sg U7148 ( .A(n7136), .B(n5737), .X(n4327) );
  nand_x2_sg U7149 ( .A(n5980), .B(n5780), .X(n4234) );
  nand_x2_sg U7150 ( .A(n6893), .B(n5789), .X(n4198) );
  nand_x2_sg U7151 ( .A(n6896), .B(n5651), .X(n4162) );
  nand_x1_sg U7152 ( .A(n9014), .B(n969), .X(n965) );
  nand_x1_sg U7153 ( .A(n1427), .B(n1428), .X(n1410) );
  nand_x1_sg U7154 ( .A(n1217), .B(n1218), .X(n1216) );
  nand_x1_sg U7155 ( .A(n1232), .B(n1233), .X(n1215) );
  nand_x1_sg U7156 ( .A(n1185), .B(n1186), .X(n1184) );
  nand_x1_sg U7157 ( .A(n1316), .B(n1317), .X(n1315) );
  nand_x1_sg U7158 ( .A(n1331), .B(n1332), .X(n1314) );
  nand_x1_sg U7159 ( .A(n1348), .B(n1349), .X(n1347) );
  nand_x1_sg U7160 ( .A(n9012), .B(n1001), .X(n997) );
  nand_x1_sg U7161 ( .A(n1035), .B(n1036), .X(n1018) );
  nand_x1_sg U7162 ( .A(n1020), .B(n1021), .X(n1019) );
  nand_x1_sg U7163 ( .A(n1067), .B(n1068), .X(n1050) );
  nand_x1_sg U7164 ( .A(n1084), .B(n1085), .X(n1083) );
  nand_x1_sg U7165 ( .A(n872), .B(n873), .X(n855) );
  nand_x1_sg U7166 ( .A(n904), .B(n905), .X(n887) );
  nand_x1_sg U7167 ( .A(n921), .B(n922), .X(n920) );
  nand_x1_sg U7168 ( .A(n1395), .B(n1396), .X(n1378) );
  nand_x1_sg U7169 ( .A(n1380), .B(n1381), .X(n1379) );
  nand_x2_sg U7170 ( .A(n5980), .B(n5656), .X(n4810) );
  nand_x2_sg U7171 ( .A(n5980), .B(n5661), .X(n4702) );
  nand_x2_sg U7172 ( .A(n6896), .B(n5671), .X(n4486) );
  nand_x2_sg U7173 ( .A(n7137), .B(n5846), .X(n4363) );
  nand_x2_sg U7174 ( .A(n7141), .B(n5820), .X(n4291) );
  nand_x2_sg U7175 ( .A(n6893), .B(n5681), .X(n4270) );
  nand_x1_sg U7176 ( .A(n1252), .B(n1253), .X(n1251) );
  nand_x1_sg U7177 ( .A(n1267), .B(n1268), .X(n1250) );
  nand_x1_sg U7178 ( .A(n1299), .B(n1300), .X(n1282) );
  nand_x1_sg U7179 ( .A(n1284), .B(n1285), .X(n1283) );
  nand_x2_sg U7180 ( .A(n2205), .B(n2206), .X(n2204) );
  nor_x1_sg U7181 ( .A(n2230), .B(n2231), .X(n2229) );
  nand_x1_sg U7182 ( .A(n2238), .B(n2239), .X(n2230) );
  nand_x1_sg U7183 ( .A(n3696), .B(n9226), .X(n3695) );
  nand_x2_sg U7184 ( .A(n778), .B(n779), .X(n777) );
  nand_x1_sg U7185 ( .A(n2192), .B(n2193), .X(n1471) );
  nand_x4_sg U7186 ( .A(n4863), .B(input_ready), .X(n4862) );
  nand_x1_sg U7187 ( .A(\i_im[1][17] ), .B(n7369), .X(n5029) );
  nand_x4_sg U7188 ( .A(n840), .B(n841), .X(n823) );
  nand_x4_sg U7189 ( .A(n808), .B(n809), .X(n785) );
  nand_x4_sg U7190 ( .A(n971), .B(n972), .X(n954) );
  nand_x4_sg U7191 ( .A(n988), .B(n989), .X(n987) );
  nand_x4_sg U7192 ( .A(n1136), .B(n1137), .X(n1119) );
  inv_x1_sg U7193 ( .A(n740), .X(n5912) );
  inv_x1_sg U7194 ( .A(n740), .X(n5913) );
  nand_x4_sg U7195 ( .A(n986), .B(n987), .X(n744) );
  inv_x1_sg U7196 ( .A(n739), .X(n5914) );
  inv_x1_sg U7197 ( .A(n739), .X(n5915) );
  nand_x4_sg U7198 ( .A(n954), .B(n955), .X(n746) );
  nand_x4_sg U7199 ( .A(n785), .B(n786), .X(n749) );
  nand_x4_sg U7200 ( .A(n823), .B(n824), .X(n750) );
  nand_x4_sg U7201 ( .A(n1119), .B(n1120), .X(n735) );
  nor_x1_sg U7202 ( .A(n4885), .B(reset), .X(n5916) );
  nand_x8_sg U7203 ( .A(n5633), .B(input_ready), .X(n4885) );
  nor_x1_sg U7204 ( .A(n6160), .B(reset), .X(n5917) );
  nand_x16_sg U7205 ( .A(n5633), .B(input_ready), .X(n6160) );
  inv_x1_sg U7206 ( .A(n7373), .X(n5918) );
  inv_x1_sg U7207 ( .A(n1466), .X(n5919) );
  inv_x1_sg U7208 ( .A(n5919), .X(n5920) );
  inv_x1_sg U7209 ( .A(n7374), .X(n5921) );
  inv_x1_sg U7210 ( .A(n6155), .X(n5922) );
  inv_x1_sg U7211 ( .A(n6273), .X(n5923) );
  inv_x1_sg U7212 ( .A(n6278), .X(n5924) );
  inv_x1_sg U7213 ( .A(n6283), .X(n5925) );
  inv_x1_sg U7214 ( .A(n6288), .X(n5926) );
  inv_x1_sg U7215 ( .A(n6238), .X(n5927) );
  inv_x1_sg U7216 ( .A(n6729), .X(n5928) );
  inv_x1_sg U7217 ( .A(n5928), .X(n5929) );
  inv_x1_sg U7218 ( .A(n6734), .X(n5930) );
  inv_x1_sg U7219 ( .A(n5930), .X(n5931) );
  inv_x1_sg U7220 ( .A(n6739), .X(n5932) );
  inv_x1_sg U7221 ( .A(n5932), .X(n5933) );
  inv_x1_sg U7222 ( .A(n6744), .X(n5934) );
  inv_x1_sg U7223 ( .A(n5934), .X(n5935) );
  inv_x1_sg U7224 ( .A(n5915), .X(n5936) );
  inv_x1_sg U7225 ( .A(n6754), .X(n5937) );
  inv_x1_sg U7226 ( .A(n5937), .X(n5938) );
  inv_x1_sg U7227 ( .A(n6759), .X(n5939) );
  inv_x1_sg U7228 ( .A(n5939), .X(n5940) );
  inv_x1_sg U7229 ( .A(n5913), .X(n5941) );
  inv_x2_sg U7230 ( .A(n748), .X(n5942) );
  inv_x1_sg U7231 ( .A(n5942), .X(n5943) );
  inv_x2_sg U7232 ( .A(n745), .X(n5944) );
  inv_x1_sg U7233 ( .A(n5944), .X(n5945) );
  inv_x2_sg U7234 ( .A(n742), .X(n5946) );
  inv_x1_sg U7235 ( .A(n5946), .X(n5947) );
  inv_x2_sg U7236 ( .A(n753), .X(n5948) );
  inv_x1_sg U7237 ( .A(n5948), .X(n5949) );
  inv_x2_sg U7238 ( .A(n755), .X(n5950) );
  inv_x1_sg U7239 ( .A(n5950), .X(n5951) );
  inv_x2_sg U7240 ( .A(n747), .X(n5952) );
  inv_x1_sg U7241 ( .A(n5952), .X(n5953) );
  inv_x2_sg U7242 ( .A(n752), .X(n5954) );
  inv_x1_sg U7243 ( .A(n5954), .X(n5955) );
  inv_x2_sg U7244 ( .A(n751), .X(n5956) );
  inv_x1_sg U7245 ( .A(n5956), .X(n5957) );
  inv_x2_sg U7246 ( .A(n738), .X(n5958) );
  inv_x1_sg U7247 ( .A(n5958), .X(n5959) );
  inv_x2_sg U7248 ( .A(n741), .X(n5960) );
  inv_x1_sg U7249 ( .A(n5960), .X(n5961) );
  inv_x1_sg U7250 ( .A(n6819), .X(n5962) );
  inv_x1_sg U7251 ( .A(n5962), .X(n5963) );
  inv_x2_sg U7252 ( .A(n737), .X(n5964) );
  inv_x1_sg U7253 ( .A(n5964), .X(n5965) );
  inv_x1_sg U7254 ( .A(n5967), .X(n5966) );
  inv_x1_sg U7255 ( .A(n6828), .X(n5967) );
  inv_x1_sg U7256 ( .A(n3656), .X(n5968) );
  inv_x1_sg U7257 ( .A(n7464), .X(n5969) );
  inv_x1_sg U7258 ( .A(n7476), .X(n5970) );
  inv_x1_sg U7259 ( .A(n7466), .X(n5971) );
  inv_x1_sg U7260 ( .A(n7470), .X(n5972) );
  inv_x1_sg U7261 ( .A(n7467), .X(n5973) );
  inv_x1_sg U7262 ( .A(n7468), .X(n5974) );
  inv_x1_sg U7263 ( .A(n7472), .X(n5975) );
  inv_x1_sg U7264 ( .A(n7474), .X(n5976) );
  inv_x1_sg U7265 ( .A(n7465), .X(n5977) );
  inv_x1_sg U7266 ( .A(n7475), .X(n5978) );
  inv_x1_sg U7267 ( .A(n7477), .X(n5979) );
  inv_x1_sg U7268 ( .A(n4146), .X(n5980) );
  inv_x1_sg U7269 ( .A(n3613), .X(n5981) );
  inv_x1_sg U7270 ( .A(n7471), .X(n5982) );
  inv_x1_sg U7271 ( .A(n7469), .X(n5983) );
  inv_x1_sg U7272 ( .A(n4884), .X(n5984) );
  inv_x1_sg U7273 ( .A(n4884), .X(n5985) );
  inv_x1_sg U7274 ( .A(n6289), .X(n5986) );
  inv_x1_sg U7275 ( .A(n6290), .X(n5987) );
  inv_x1_sg U7276 ( .A(n6285), .X(n5988) );
  inv_x1_sg U7277 ( .A(n6284), .X(n5989) );
  inv_x1_sg U7278 ( .A(n6280), .X(n5990) );
  inv_x1_sg U7279 ( .A(n6279), .X(n5991) );
  inv_x1_sg U7280 ( .A(n6274), .X(n5992) );
  inv_x1_sg U7281 ( .A(n6275), .X(n5993) );
  inv_x1_sg U7282 ( .A(n6269), .X(n5994) );
  inv_x1_sg U7283 ( .A(n6270), .X(n5995) );
  inv_x1_sg U7284 ( .A(n6266), .X(n5996) );
  inv_x1_sg U7285 ( .A(n6142), .X(n5997) );
  inv_x1_sg U7286 ( .A(n1521), .X(n5998) );
  inv_x1_sg U7287 ( .A(n5998), .X(n5999) );
  inv_x1_sg U7288 ( .A(n7053), .X(n6000) );
  inv_x1_sg U7289 ( .A(n1520), .X(n6001) );
  inv_x1_sg U7290 ( .A(n6001), .X(n6002) );
  inv_x1_sg U7291 ( .A(n7058), .X(n6003) );
  inv_x1_sg U7292 ( .A(n7063), .X(n6004) );
  inv_x1_sg U7293 ( .A(n6123), .X(n6005) );
  inv_x1_sg U7294 ( .A(n792), .X(n6006) );
  inv_x1_sg U7295 ( .A(n6169), .X(n6007) );
  inv_x1_sg U7296 ( .A(n6169), .X(n6008) );
  inv_x1_sg U7297 ( .A(n1534), .X(n6009) );
  inv_x1_sg U7298 ( .A(n6009), .X(n6010) );
  inv_x1_sg U7299 ( .A(n7087), .X(n6011) );
  inv_x1_sg U7300 ( .A(n1524), .X(n6012) );
  inv_x1_sg U7301 ( .A(n6012), .X(n6013) );
  inv_x1_sg U7302 ( .A(n7092), .X(n6014) );
  inv_x1_sg U7303 ( .A(n1526), .X(n6015) );
  inv_x1_sg U7304 ( .A(n6015), .X(n6016) );
  inv_x1_sg U7305 ( .A(n7097), .X(n6017) );
  inv_x1_sg U7306 ( .A(n734), .X(n6018) );
  inv_x1_sg U7307 ( .A(n6018), .X(n6019) );
  inv_x1_sg U7308 ( .A(n7102), .X(n6020) );
  inv_x1_sg U7309 ( .A(n772), .X(n6021) );
  inv_x1_sg U7310 ( .A(n6021), .X(n6022) );
  inv_x1_sg U7311 ( .A(n7107), .X(n6023) );
  inv_x1_sg U7312 ( .A(n766), .X(n6024) );
  inv_x1_sg U7313 ( .A(n6024), .X(n6025) );
  inv_x1_sg U7314 ( .A(n7112), .X(n6026) );
  inv_x1_sg U7315 ( .A(n759), .X(n6027) );
  inv_x1_sg U7316 ( .A(n6027), .X(n6028) );
  inv_x1_sg U7317 ( .A(n7117), .X(n6029) );
  inv_x1_sg U7318 ( .A(n4151), .X(n6030) );
  inv_x1_sg U7319 ( .A(n6193), .X(n6031) );
  inv_x1_sg U7320 ( .A(n6030), .X(n6032) );
  inv_x1_sg U7321 ( .A(n806), .X(n6033) );
  inv_x1_sg U7322 ( .A(n7143), .X(n6034) );
  inv_x1_sg U7323 ( .A(n6033), .X(n6035) );
  inv_x1_sg U7324 ( .A(n770), .X(n6036) );
  inv_x1_sg U7325 ( .A(n6036), .X(n6037) );
  inv_x1_sg U7326 ( .A(n7163), .X(n6038) );
  inv_x1_sg U7327 ( .A(n768), .X(n6039) );
  inv_x1_sg U7328 ( .A(n6039), .X(n6040) );
  inv_x1_sg U7329 ( .A(n7168), .X(n6041) );
  inv_x1_sg U7330 ( .A(n758), .X(n6042) );
  inv_x1_sg U7331 ( .A(n6042), .X(n6043) );
  inv_x1_sg U7332 ( .A(n7173), .X(n6044) );
  inv_x1_sg U7333 ( .A(n754), .X(n6045) );
  inv_x1_sg U7334 ( .A(n6045), .X(n6046) );
  inv_x1_sg U7335 ( .A(n7178), .X(n6047) );
  inv_x1_sg U7336 ( .A(n776), .X(n6048) );
  inv_x1_sg U7337 ( .A(n6048), .X(n6049) );
  inv_x1_sg U7338 ( .A(n7183), .X(n6050) );
  inv_x1_sg U7339 ( .A(n775), .X(n6051) );
  inv_x1_sg U7340 ( .A(n6051), .X(n6052) );
  inv_x1_sg U7341 ( .A(n7188), .X(n6053) );
  inv_x1_sg U7342 ( .A(n774), .X(n6054) );
  inv_x1_sg U7343 ( .A(n6054), .X(n6055) );
  inv_x1_sg U7344 ( .A(n7193), .X(n6056) );
  inv_x1_sg U7345 ( .A(n764), .X(n6057) );
  inv_x1_sg U7346 ( .A(n6057), .X(n6058) );
  inv_x1_sg U7347 ( .A(n7198), .X(n6059) );
  inv_x1_sg U7348 ( .A(n763), .X(n6060) );
  inv_x1_sg U7349 ( .A(n6060), .X(n6061) );
  inv_x1_sg U7350 ( .A(n7203), .X(n6062) );
  inv_x1_sg U7351 ( .A(n762), .X(n6063) );
  inv_x1_sg U7352 ( .A(n6063), .X(n6064) );
  inv_x1_sg U7353 ( .A(n7208), .X(n6065) );
  inv_x1_sg U7354 ( .A(n769), .X(n6066) );
  inv_x1_sg U7355 ( .A(n6066), .X(n6067) );
  inv_x1_sg U7356 ( .A(n7213), .X(n6068) );
  inv_x1_sg U7357 ( .A(n757), .X(n6069) );
  inv_x1_sg U7358 ( .A(n6069), .X(n6070) );
  inv_x1_sg U7359 ( .A(n7218), .X(n6071) );
  inv_x1_sg U7360 ( .A(n7444), .X(n6072) );
  inv_x1_sg U7361 ( .A(n6072), .X(n6073) );
  inv_x1_sg U7362 ( .A(n7223), .X(n6074) );
  inv_x1_sg U7363 ( .A(n4140), .X(n6075) );
  inv_x1_sg U7364 ( .A(n6075), .X(n6076) );
  inv_x1_sg U7365 ( .A(n6235), .X(n6077) );
  inv_x1_sg U7366 ( .A(n7462), .X(n6078) );
  inv_x1_sg U7367 ( .A(n7313), .X(n6079) );
  inv_x1_sg U7368 ( .A(n6079), .X(n6080) );
  inv_x1_sg U7369 ( .A(n6471), .X(n6081) );
  inv_x1_sg U7370 ( .A(n7317), .X(n6082) );
  inv_x1_sg U7371 ( .A(n6239), .X(n6083) );
  inv_x1_sg U7372 ( .A(n6162), .X(n6084) );
  inv_x1_sg U7373 ( .A(n6089), .X(n6085) );
  inv_x1_sg U7374 ( .A(n5916), .X(n6086) );
  inv_x1_sg U7375 ( .A(n6086), .X(n6087) );
  inv_x1_sg U7376 ( .A(n6533), .X(n6088) );
  inv_x1_sg U7377 ( .A(n5917), .X(n6089) );
  inv_x1_sg U7378 ( .A(n6304), .X(n6090) );
  inv_x1_sg U7379 ( .A(n6161), .X(n6091) );
  inv_x1_sg U7380 ( .A(n6252), .X(n6092) );
  inv_x1_sg U7381 ( .A(n4855), .X(n6093) );
  inv_x1_sg U7382 ( .A(\output_state[0] ), .X(n6094) );
  inv_x1_sg U7383 ( .A(n6094), .X(n6095) );
  inv_x1_sg U7384 ( .A(n7395), .X(n6096) );
  inv_x1_sg U7385 ( .A(\update_mask_0/N23 ), .X(n6097) );
  inv_x1_sg U7386 ( .A(n6097), .X(n6098) );
  inv_x1_sg U7387 ( .A(\update_mask_0/N28 ), .X(n6099) );
  inv_x1_sg U7388 ( .A(n6099), .X(n6100) );
  inv_x1_sg U7389 ( .A(n7396), .X(n6101) );
  inv_x1_sg U7390 ( .A(n6921), .X(n6102) );
  inv_x1_sg U7391 ( .A(n6926), .X(n6103) );
  inv_x1_sg U7392 ( .A(n7380), .X(n6104) );
  inv_x1_sg U7393 ( .A(n6936), .X(n6105) );
  inv_x1_sg U7394 ( .A(n6941), .X(n6106) );
  inv_x1_sg U7395 ( .A(n6946), .X(n6107) );
  inv_x1_sg U7396 ( .A(n6951), .X(n6108) );
  inv_x1_sg U7397 ( .A(n6956), .X(n6109) );
  inv_x1_sg U7398 ( .A(n6961), .X(n6110) );
  inv_x1_sg U7399 ( .A(n6966), .X(n6111) );
  inv_x1_sg U7400 ( .A(n6971), .X(n6112) );
  inv_x1_sg U7401 ( .A(n6976), .X(n6113) );
  inv_x1_sg U7402 ( .A(n6981), .X(n6114) );
  inv_x1_sg U7403 ( .A(n6986), .X(n6115) );
  inv_x1_sg U7404 ( .A(n6991), .X(n6116) );
  inv_x1_sg U7405 ( .A(n7417), .X(n6117) );
  inv_x1_sg U7406 ( .A(n6117), .X(n6118) );
  inv_x1_sg U7407 ( .A(n7010), .X(n6119) );
  inv_x1_sg U7408 ( .A(n5985), .X(n6120) );
  inv_x1_sg U7409 ( .A(n6120), .X(n6121) );
  inv_x1_sg U7410 ( .A(n7015), .X(n6122) );
  inv_x1_sg U7411 ( .A(n4154), .X(n6123) );
  inv_x1_sg U7412 ( .A(n6126), .X(n6124) );
  inv_x1_sg U7413 ( .A(n6124), .X(n6125) );
  inv_x1_sg U7414 ( .A(n7272), .X(n6126) );
  inv_x1_sg U7415 ( .A(n6129), .X(n6127) );
  inv_x1_sg U7416 ( .A(n6127), .X(n6128) );
  inv_x1_sg U7417 ( .A(n7277), .X(n6129) );
  inv_x1_sg U7418 ( .A(n6132), .X(n6130) );
  inv_x1_sg U7419 ( .A(n6130), .X(n6131) );
  inv_x1_sg U7420 ( .A(n7282), .X(n6132) );
  inv_x1_sg U7421 ( .A(n6484), .X(n6133) );
  inv_x1_sg U7422 ( .A(n7302), .X(n6134) );
  inv_x1_sg U7423 ( .A(n7302), .X(n6135) );
  inv_x1_sg U7424 ( .A(n6480), .X(n6136) );
  inv_x1_sg U7425 ( .A(n7307), .X(n6137) );
  inv_x1_sg U7426 ( .A(n7307), .X(n6138) );
  inv_x1_sg U7427 ( .A(\update_output_0/N34 ), .X(n6139) );
  inv_x1_sg U7428 ( .A(n7312), .X(n6140) );
  inv_x1_sg U7429 ( .A(n6139), .X(n6141) );
  inv_x1_sg U7430 ( .A(n6149), .X(n6142) );
  inv_x1_sg U7431 ( .A(n6142), .X(n6143) );
  inv_x1_sg U7432 ( .A(n6142), .X(n6144) );
  inv_x1_sg U7433 ( .A(n6242), .X(n6145) );
  inv_x1_sg U7434 ( .A(n7324), .X(n6146) );
  inv_x1_sg U7435 ( .A(n7323), .X(n6147) );
  inv_x1_sg U7436 ( .A(n6147), .X(n6148) );
  inv_x1_sg U7437 ( .A(n6147), .X(n6149) );
  inv_x1_sg U7438 ( .A(n6243), .X(n6150) );
  inv_x1_sg U7439 ( .A(n7328), .X(n6151) );
  inv_x1_sg U7440 ( .A(n7463), .X(n6152) );
  inv_x1_sg U7441 ( .A(n6152), .X(n6153) );
  inv_x1_sg U7442 ( .A(n6152), .X(n6154) );
  inv_x1_sg U7443 ( .A(n6244), .X(n6155) );
  inv_x1_sg U7444 ( .A(n7332), .X(n6156) );
  inv_x1_sg U7445 ( .A(n3479), .X(n6157) );
  inv_x1_sg U7446 ( .A(n6510), .X(n6158) );
  nand_x8_sg U7447 ( .A(n5633), .B(input_ready), .X(n6159) );
  nor_x1_sg U7448 ( .A(n6160), .B(reset), .X(n6161) );
  nor_x1_sg U7449 ( .A(n6159), .B(reset), .X(n6162) );
  inv_x1_sg U7450 ( .A(n1521), .X(n6163) );
  inv_x1_sg U7451 ( .A(n7053), .X(n6164) );
  inv_x1_sg U7452 ( .A(n6163), .X(n6165) );
  inv_x1_sg U7453 ( .A(n1520), .X(n6166) );
  inv_x1_sg U7454 ( .A(n7058), .X(n6167) );
  inv_x1_sg U7455 ( .A(n6166), .X(n6168) );
  inv_x1_sg U7456 ( .A(n792), .X(n6169) );
  inv_x1_sg U7457 ( .A(n6006), .X(n6170) );
  inv_x1_sg U7458 ( .A(n6169), .X(n6171) );
  inv_x1_sg U7459 ( .A(n1534), .X(n6172) );
  inv_x1_sg U7460 ( .A(n7087), .X(n6173) );
  inv_x1_sg U7461 ( .A(n6172), .X(n6174) );
  inv_x1_sg U7462 ( .A(n1524), .X(n6175) );
  inv_x1_sg U7463 ( .A(n7092), .X(n6176) );
  inv_x1_sg U7464 ( .A(n6175), .X(n6177) );
  inv_x1_sg U7465 ( .A(n1526), .X(n6178) );
  inv_x1_sg U7466 ( .A(n7097), .X(n6179) );
  inv_x1_sg U7467 ( .A(n6178), .X(n6180) );
  inv_x1_sg U7468 ( .A(n734), .X(n6181) );
  inv_x1_sg U7469 ( .A(n7102), .X(n6182) );
  inv_x1_sg U7470 ( .A(n6181), .X(n6183) );
  inv_x1_sg U7471 ( .A(n772), .X(n6184) );
  inv_x1_sg U7472 ( .A(n7107), .X(n6185) );
  inv_x1_sg U7473 ( .A(n6184), .X(n6186) );
  inv_x1_sg U7474 ( .A(n766), .X(n6187) );
  inv_x1_sg U7475 ( .A(n7112), .X(n6188) );
  inv_x1_sg U7476 ( .A(n6187), .X(n6189) );
  inv_x1_sg U7477 ( .A(n759), .X(n6190) );
  inv_x1_sg U7478 ( .A(n7117), .X(n6191) );
  inv_x1_sg U7479 ( .A(n6190), .X(n6192) );
  inv_x1_sg U7480 ( .A(n4151), .X(n6193) );
  inv_x1_sg U7481 ( .A(n6193), .X(n6194) );
  inv_x1_sg U7482 ( .A(n7122), .X(n6195) );
  inv_x1_sg U7483 ( .A(n770), .X(n6196) );
  inv_x1_sg U7484 ( .A(n7163), .X(n6197) );
  inv_x1_sg U7485 ( .A(n6196), .X(n6198) );
  inv_x1_sg U7486 ( .A(n768), .X(n6199) );
  inv_x1_sg U7487 ( .A(n7168), .X(n6200) );
  inv_x1_sg U7488 ( .A(n6199), .X(n6201) );
  inv_x1_sg U7489 ( .A(n758), .X(n6202) );
  inv_x1_sg U7490 ( .A(n7173), .X(n6203) );
  inv_x1_sg U7491 ( .A(n6202), .X(n6204) );
  inv_x1_sg U7492 ( .A(n754), .X(n6205) );
  inv_x1_sg U7493 ( .A(n7178), .X(n6206) );
  inv_x1_sg U7494 ( .A(n6205), .X(n6207) );
  inv_x1_sg U7495 ( .A(n776), .X(n6208) );
  inv_x1_sg U7496 ( .A(n7183), .X(n6209) );
  inv_x1_sg U7497 ( .A(n6208), .X(n6210) );
  inv_x1_sg U7498 ( .A(n775), .X(n6211) );
  inv_x1_sg U7499 ( .A(n7188), .X(n6212) );
  inv_x1_sg U7500 ( .A(n6211), .X(n6213) );
  inv_x1_sg U7501 ( .A(n774), .X(n6214) );
  inv_x1_sg U7502 ( .A(n7193), .X(n6215) );
  inv_x1_sg U7503 ( .A(n6214), .X(n6216) );
  inv_x1_sg U7504 ( .A(n764), .X(n6217) );
  inv_x1_sg U7505 ( .A(n7198), .X(n6218) );
  inv_x1_sg U7506 ( .A(n6217), .X(n6219) );
  inv_x1_sg U7507 ( .A(n763), .X(n6220) );
  inv_x1_sg U7508 ( .A(n7203), .X(n6221) );
  inv_x1_sg U7509 ( .A(n6220), .X(n6222) );
  inv_x1_sg U7510 ( .A(n762), .X(n6223) );
  inv_x1_sg U7511 ( .A(n7208), .X(n6224) );
  inv_x1_sg U7512 ( .A(n6223), .X(n6225) );
  inv_x1_sg U7513 ( .A(n769), .X(n6226) );
  inv_x1_sg U7514 ( .A(n7213), .X(n6227) );
  inv_x1_sg U7515 ( .A(n6226), .X(n6228) );
  inv_x1_sg U7516 ( .A(n757), .X(n6229) );
  inv_x1_sg U7517 ( .A(n7218), .X(n6230) );
  inv_x1_sg U7518 ( .A(n6229), .X(n6231) );
  inv_x1_sg U7519 ( .A(n7444), .X(n6232) );
  inv_x1_sg U7520 ( .A(n7223), .X(n6233) );
  inv_x1_sg U7521 ( .A(n6232), .X(n6234) );
  inv_x1_sg U7522 ( .A(n4140), .X(n6235) );
  inv_x1_sg U7523 ( .A(n6235), .X(n6236) );
  inv_x1_sg U7524 ( .A(n7254), .X(n6237) );
  inv_x1_sg U7525 ( .A(\update_output_0/N30 ), .X(n6238) );
  inv_x1_sg U7526 ( .A(\update_output_0/N30 ), .X(n6239) );
  inv_x1_sg U7527 ( .A(n6238), .X(n6240) );
  inv_x1_sg U7528 ( .A(n6239), .X(n6241) );
  inv_x1_sg U7529 ( .A(n7463), .X(n6242) );
  inv_x1_sg U7530 ( .A(n7323), .X(n6243) );
  inv_x1_sg U7531 ( .A(n7463), .X(n6244) );
  inv_x1_sg U7532 ( .A(n5917), .X(n6245) );
  inv_x1_sg U7533 ( .A(n7336), .X(n6246) );
  inv_x1_sg U7534 ( .A(n7337), .X(n6247) );
  inv_x1_sg U7535 ( .A(n7339), .X(n6248) );
  inv_x1_sg U7536 ( .A(n6246), .X(n6249) );
  inv_x1_sg U7537 ( .A(n7355), .X(n6250) );
  inv_x1_sg U7538 ( .A(n6162), .X(n6251) );
  inv_x1_sg U7539 ( .A(n4892), .X(n6252) );
  inv_x1_sg U7540 ( .A(n6251), .X(n6253) );
  inv_x1_sg U7541 ( .A(n6299), .X(n6254) );
  inv_x1_sg U7542 ( .A(n6245), .X(n6255) );
  inv_x1_sg U7543 ( .A(n6252), .X(n6256) );
  inv_x1_sg U7544 ( .A(n6303), .X(n6257) );
  inv_x1_sg U7545 ( .A(n7355), .X(n6258) );
  inv_x1_sg U7546 ( .A(n6303), .X(n6259) );
  inv_x1_sg U7547 ( .A(n6091), .X(n6260) );
  inv_x1_sg U7548 ( .A(n6084), .X(n6261) );
  inv_x1_sg U7549 ( .A(n6252), .X(n6262) );
  inv_x1_sg U7550 ( .A(n7002), .X(n6263) );
  inv_x1_sg U7551 ( .A(n7048), .X(n6264) );
  inv_x1_sg U7552 ( .A(n6264), .X(n6265) );
  inv_x1_sg U7553 ( .A(n6264), .X(n6266) );
  inv_x1_sg U7554 ( .A(n6265), .X(n6267) );
  inv_x1_sg U7555 ( .A(n6265), .X(n6268) );
  inv_x1_sg U7556 ( .A(n6156), .X(n6269) );
  inv_x1_sg U7557 ( .A(n6154), .X(n6270) );
  inv_x1_sg U7558 ( .A(n6270), .X(n6271) );
  inv_x1_sg U7559 ( .A(n6270), .X(n6272) );
  inv_x1_sg U7560 ( .A(n7037), .X(n6273) );
  inv_x1_sg U7561 ( .A(n6273), .X(n6274) );
  inv_x1_sg U7562 ( .A(n6273), .X(n6275) );
  inv_x1_sg U7563 ( .A(n6275), .X(n6276) );
  inv_x1_sg U7564 ( .A(n6275), .X(n6277) );
  inv_x1_sg U7565 ( .A(n7032), .X(n6278) );
  inv_x1_sg U7566 ( .A(n6278), .X(n6279) );
  inv_x1_sg U7567 ( .A(n6278), .X(n6280) );
  inv_x1_sg U7568 ( .A(n6279), .X(n6281) );
  inv_x1_sg U7569 ( .A(n6279), .X(n6282) );
  inv_x1_sg U7570 ( .A(n5922), .X(n6283) );
  inv_x1_sg U7571 ( .A(n6283), .X(n6284) );
  inv_x1_sg U7572 ( .A(n6283), .X(n6285) );
  inv_x1_sg U7573 ( .A(n6284), .X(n6286) );
  inv_x1_sg U7574 ( .A(n6284), .X(n6287) );
  inv_x1_sg U7575 ( .A(n6269), .X(n6288) );
  inv_x1_sg U7576 ( .A(n6288), .X(n6289) );
  inv_x1_sg U7577 ( .A(n6288), .X(n6290) );
  inv_x1_sg U7578 ( .A(n6290), .X(n6291) );
  inv_x1_sg U7579 ( .A(n6290), .X(n6292) );
  inv_x1_sg U7580 ( .A(n6086), .X(n6293) );
  inv_x1_sg U7581 ( .A(n6251), .X(n6294) );
  inv_x1_sg U7582 ( .A(n6246), .X(n6295) );
  inv_x1_sg U7583 ( .A(n6084), .X(n6296) );
  inv_x1_sg U7584 ( .A(n7357), .X(n6297) );
  inv_x1_sg U7585 ( .A(n6089), .X(n6298) );
  inv_x1_sg U7586 ( .A(n4892), .X(n6299) );
  inv_x1_sg U7587 ( .A(n5916), .X(n6300) );
  inv_x1_sg U7588 ( .A(n6300), .X(n6301) );
  inv_x1_sg U7589 ( .A(n7337), .X(n6302) );
  inv_x1_sg U7590 ( .A(n4892), .X(n6303) );
  inv_x1_sg U7591 ( .A(n6162), .X(n6304) );
  inv_x1_sg U7592 ( .A(n6091), .X(n6305) );
  inv_x1_sg U7593 ( .A(n6304), .X(n6306) );
  inv_x1_sg U7594 ( .A(\update_mask_0/N26 ), .X(n6307) );
  inv_x1_sg U7595 ( .A(n6307), .X(n6308) );
  inv_x1_sg U7596 ( .A(n7403), .X(n6309) );
  inv_x1_sg U7597 ( .A(n7402), .X(n6310) );
  inv_x1_sg U7598 ( .A(\update_output_0/N33 ), .X(n6311) );
  inv_x1_sg U7599 ( .A(n7401), .X(n6312) );
  inv_x1_sg U7600 ( .A(n7399), .X(n6313) );
  inv_x1_sg U7601 ( .A(n3524), .X(n6314) );
  inv_x1_sg U7602 ( .A(n6314), .X(n6315) );
  inv_x1_sg U7603 ( .A(n1482), .X(n6316) );
  inv_x1_sg U7604 ( .A(n1493), .X(n6317) );
  inv_x1_sg U7605 ( .A(n1500), .X(n6318) );
  inv_x1_sg U7606 ( .A(n1468), .X(n6319) );
  inv_x1_sg U7607 ( .A(n4821), .X(n6320) );
  inv_x1_sg U7608 ( .A(n7473), .X(n6321) );
  inv_x1_sg U7609 ( .A(n806), .X(n6322) );
  inv_x1_sg U7610 ( .A(n6322), .X(n6323) );
  inv_x1_sg U7611 ( .A(n7143), .X(n6324) );
  inv_x1_sg U7612 ( .A(n6117), .X(n6325) );
  inv_x1_sg U7613 ( .A(n7010), .X(n6326) );
  inv_x1_sg U7614 ( .A(n7407), .X(n6327) );
  inv_x1_sg U7615 ( .A(\update_mask_0/n2986 ), .X(n6328) );
  inv_x1_sg U7616 ( .A(n6328), .X(n6329) );
  inv_x1_sg U7617 ( .A(n6328), .X(n6330) );
  inv_x1_sg U7618 ( .A(\update_output_0/N31 ), .X(n6331) );
  inv_x1_sg U7619 ( .A(n6331), .X(n6332) );
  inv_x1_sg U7620 ( .A(n6331), .X(n6333) );
  inv_x1_sg U7621 ( .A(n7473), .X(n6334) );
  inv_x1_sg U7622 ( .A(n6334), .X(n6335) );
  inv_x1_sg U7623 ( .A(n6334), .X(n6336) );
  inv_x1_sg U7624 ( .A(n7455), .X(n6337) );
  inv_x1_sg U7625 ( .A(n6337), .X(n6338) );
  inv_x1_sg U7626 ( .A(n6337), .X(n6339) );
  inv_x1_sg U7627 ( .A(n7454), .X(n6340) );
  inv_x1_sg U7628 ( .A(n6340), .X(n6341) );
  inv_x1_sg U7629 ( .A(n6340), .X(n6342) );
  inv_x1_sg U7630 ( .A(n7453), .X(n6343) );
  inv_x1_sg U7631 ( .A(n6343), .X(n6344) );
  inv_x1_sg U7632 ( .A(n6343), .X(n6345) );
  inv_x1_sg U7633 ( .A(n1446), .X(n6346) );
  inv_x1_sg U7634 ( .A(n6346), .X(n6347) );
  inv_x1_sg U7635 ( .A(n6346), .X(n6348) );
  inv_x1_sg U7636 ( .A(n7443), .X(n6349) );
  inv_x1_sg U7637 ( .A(n6349), .X(n6350) );
  inv_x1_sg U7638 ( .A(n6349), .X(n6351) );
  inv_x1_sg U7639 ( .A(n1449), .X(n6352) );
  inv_x1_sg U7640 ( .A(n6352), .X(n6353) );
  inv_x1_sg U7641 ( .A(n6352), .X(n6354) );
  inv_x1_sg U7642 ( .A(n6244), .X(n6355) );
  inv_x1_sg U7643 ( .A(n7332), .X(n6356) );
  inv_x1_sg U7644 ( .A(n6243), .X(n6357) );
  inv_x1_sg U7645 ( .A(n7328), .X(n6358) );
  inv_x1_sg U7646 ( .A(n6242), .X(n6359) );
  inv_x1_sg U7647 ( .A(n7324), .X(n6360) );
  inv_x1_sg U7648 ( .A(n6238), .X(n6361) );
  inv_x1_sg U7649 ( .A(n6238), .X(n6362) );
  inv_x1_sg U7650 ( .A(n6120), .X(n6363) );
  inv_x1_sg U7651 ( .A(n7015), .X(n6364) );
  inv_x1_sg U7652 ( .A(\update_mask_0/N24 ), .X(n6365) );
  inv_x1_sg U7653 ( .A(n6365), .X(n6366) );
  inv_x1_sg U7654 ( .A(n6365), .X(n6367) );
  inv_x1_sg U7655 ( .A(\update_output_0/N27 ), .X(n6368) );
  inv_x1_sg U7656 ( .A(n6368), .X(n6369) );
  inv_x1_sg U7657 ( .A(n1452), .X(n6370) );
  inv_x1_sg U7658 ( .A(n6370), .X(n6371) );
  inv_x1_sg U7659 ( .A(n6370), .X(n6372) );
  inv_x1_sg U7660 ( .A(n1455), .X(n6373) );
  inv_x1_sg U7661 ( .A(n6373), .X(n6374) );
  inv_x1_sg U7662 ( .A(n6373), .X(n6375) );
  inv_x1_sg U7663 ( .A(n1459), .X(n6376) );
  inv_x1_sg U7664 ( .A(n6376), .X(n6377) );
  inv_x1_sg U7665 ( .A(n6376), .X(n6378) );
  inv_x1_sg U7666 ( .A(n7442), .X(n6379) );
  inv_x1_sg U7667 ( .A(n6379), .X(n6380) );
  inv_x1_sg U7668 ( .A(n6379), .X(n6381) );
  inv_x1_sg U7669 ( .A(n7446), .X(n6382) );
  inv_x1_sg U7670 ( .A(n6382), .X(n6383) );
  inv_x1_sg U7671 ( .A(n6382), .X(n6384) );
  inv_x1_sg U7672 ( .A(n6133), .X(n6385) );
  inv_x1_sg U7673 ( .A(n7302), .X(n6386) );
  inv_x1_sg U7674 ( .A(n6130), .X(n6387) );
  inv_x1_sg U7675 ( .A(n7282), .X(n6388) );
  inv_x1_sg U7676 ( .A(n6127), .X(n6389) );
  inv_x1_sg U7677 ( .A(n6127), .X(n6390) );
  inv_x1_sg U7678 ( .A(n6124), .X(n6391) );
  inv_x1_sg U7679 ( .A(n6124), .X(n6392) );
  inv_x1_sg U7680 ( .A(n6235), .X(n6393) );
  inv_x1_sg U7681 ( .A(n7254), .X(n6394) );
  inv_x1_sg U7682 ( .A(n6072), .X(n6395) );
  inv_x1_sg U7683 ( .A(n6072), .X(n6396) );
  inv_x1_sg U7684 ( .A(n6069), .X(n6397) );
  inv_x1_sg U7685 ( .A(n6069), .X(n6398) );
  inv_x1_sg U7686 ( .A(n6066), .X(n6399) );
  inv_x1_sg U7687 ( .A(n6066), .X(n6400) );
  inv_x1_sg U7688 ( .A(n6063), .X(n6401) );
  inv_x1_sg U7689 ( .A(n6063), .X(n6402) );
  inv_x1_sg U7690 ( .A(n6060), .X(n6403) );
  inv_x1_sg U7691 ( .A(n6060), .X(n6404) );
  inv_x1_sg U7692 ( .A(n6057), .X(n6405) );
  inv_x1_sg U7693 ( .A(n6057), .X(n6406) );
  inv_x1_sg U7694 ( .A(n6054), .X(n6407) );
  inv_x1_sg U7695 ( .A(n6054), .X(n6408) );
  inv_x1_sg U7696 ( .A(n6051), .X(n6409) );
  inv_x1_sg U7697 ( .A(n6051), .X(n6410) );
  inv_x1_sg U7698 ( .A(n6048), .X(n6411) );
  inv_x1_sg U7699 ( .A(n6048), .X(n6412) );
  inv_x1_sg U7700 ( .A(n6045), .X(n6413) );
  inv_x1_sg U7701 ( .A(n6045), .X(n6414) );
  inv_x1_sg U7702 ( .A(n6042), .X(n6415) );
  inv_x1_sg U7703 ( .A(n6042), .X(n6416) );
  inv_x1_sg U7704 ( .A(n6039), .X(n6417) );
  inv_x1_sg U7705 ( .A(n6039), .X(n6418) );
  inv_x1_sg U7706 ( .A(n6036), .X(n6419) );
  inv_x1_sg U7707 ( .A(n6036), .X(n6420) );
  inv_x1_sg U7708 ( .A(n7143), .X(n6421) );
  inv_x1_sg U7709 ( .A(n7143), .X(n6422) );
  inv_x1_sg U7710 ( .A(n7122), .X(n6423) );
  inv_x1_sg U7711 ( .A(n6193), .X(n6424) );
  inv_x1_sg U7712 ( .A(n6027), .X(n6425) );
  inv_x1_sg U7713 ( .A(n6027), .X(n6426) );
  inv_x1_sg U7714 ( .A(n6024), .X(n6427) );
  inv_x1_sg U7715 ( .A(n6024), .X(n6428) );
  inv_x1_sg U7716 ( .A(n6021), .X(n6429) );
  inv_x1_sg U7717 ( .A(n6021), .X(n6430) );
  inv_x1_sg U7718 ( .A(n6018), .X(n6431) );
  inv_x1_sg U7719 ( .A(n6018), .X(n6432) );
  inv_x1_sg U7720 ( .A(n6015), .X(n6433) );
  inv_x1_sg U7721 ( .A(n6015), .X(n6434) );
  inv_x1_sg U7722 ( .A(n6012), .X(n6435) );
  inv_x1_sg U7723 ( .A(n6012), .X(n6436) );
  inv_x1_sg U7724 ( .A(n6009), .X(n6437) );
  inv_x1_sg U7725 ( .A(n6009), .X(n6438) );
  inv_x1_sg U7726 ( .A(n6006), .X(n6439) );
  inv_x1_sg U7727 ( .A(n6169), .X(n6440) );
  inv_x1_sg U7728 ( .A(n6001), .X(n6441) );
  inv_x1_sg U7729 ( .A(n6001), .X(n6442) );
  inv_x1_sg U7730 ( .A(n5998), .X(n6443) );
  inv_x1_sg U7731 ( .A(n5998), .X(n6444) );
  inv_x1_sg U7732 ( .A(n6152), .X(n6445) );
  inv_x1_sg U7733 ( .A(n6266), .X(n6446) );
  inv_x1_sg U7734 ( .A(n5922), .X(n6447) );
  inv_x1_sg U7735 ( .A(n6270), .X(n6448) );
  inv_x1_sg U7736 ( .A(n5923), .X(n6449) );
  inv_x1_sg U7737 ( .A(n6275), .X(n6450) );
  inv_x1_sg U7738 ( .A(n5924), .X(n6451) );
  inv_x1_sg U7739 ( .A(n6279), .X(n6452) );
  inv_x1_sg U7740 ( .A(n5925), .X(n6453) );
  inv_x1_sg U7741 ( .A(n6284), .X(n6454) );
  inv_x1_sg U7742 ( .A(n5926), .X(n6455) );
  inv_x1_sg U7743 ( .A(n6290), .X(n6456) );
  inv_x1_sg U7744 ( .A(\update_output_0/N27 ), .X(n6457) );
  inv_x1_sg U7745 ( .A(\update_output_0/N27 ), .X(n6458) );
  inv_x1_sg U7746 ( .A(n7419), .X(n6459) );
  inv_x1_sg U7747 ( .A(n6459), .X(n6460) );
  inv_x1_sg U7748 ( .A(n6459), .X(n6461) );
  inv_x1_sg U7749 ( .A(n6459), .X(n6462) );
  inv_x1_sg U7750 ( .A(n7356), .X(n6463) );
  inv_x1_sg U7751 ( .A(n6303), .X(n6464) );
  inv_x1_sg U7752 ( .A(n6161), .X(n6465) );
  inv_x1_sg U7753 ( .A(n6465), .X(n6466) );
  inv_x1_sg U7754 ( .A(n6465), .X(n6467) );
  inv_x1_sg U7755 ( .A(n6465), .X(n6468) );
  inv_x1_sg U7756 ( .A(n7312), .X(n6469) );
  inv_x1_sg U7757 ( .A(n6139), .X(n6470) );
  inv_x1_sg U7758 ( .A(n7313), .X(n6471) );
  inv_x1_sg U7759 ( .A(n6471), .X(n6472) );
  inv_x1_sg U7760 ( .A(n6471), .X(n6473) );
  inv_x1_sg U7761 ( .A(n6471), .X(n6474) );
  inv_x1_sg U7762 ( .A(n6136), .X(n6475) );
  inv_x1_sg U7763 ( .A(n6136), .X(n6476) );
  inv_x1_sg U7764 ( .A(n7308), .X(n6477) );
  inv_x1_sg U7765 ( .A(n6477), .X(n6478) );
  inv_x1_sg U7766 ( .A(n6477), .X(n6479) );
  inv_x1_sg U7767 ( .A(n6477), .X(n6480) );
  inv_x1_sg U7768 ( .A(n7303), .X(n6481) );
  inv_x1_sg U7769 ( .A(n6481), .X(n6482) );
  inv_x1_sg U7770 ( .A(n6481), .X(n6483) );
  inv_x1_sg U7771 ( .A(n6481), .X(n6484) );
  inv_x1_sg U7772 ( .A(n7283), .X(n6485) );
  inv_x1_sg U7773 ( .A(n6485), .X(n6486) );
  inv_x1_sg U7774 ( .A(n6485), .X(n6487) );
  inv_x1_sg U7775 ( .A(n6485), .X(n6488) );
  inv_x1_sg U7776 ( .A(n7278), .X(n6489) );
  inv_x1_sg U7777 ( .A(n6489), .X(n6490) );
  inv_x1_sg U7778 ( .A(n6489), .X(n6491) );
  inv_x1_sg U7779 ( .A(n6489), .X(n6492) );
  inv_x1_sg U7780 ( .A(n7273), .X(n6493) );
  inv_x1_sg U7781 ( .A(n6493), .X(n6494) );
  inv_x1_sg U7782 ( .A(n6493), .X(n6495) );
  inv_x1_sg U7783 ( .A(n6493), .X(n6496) );
  inv_x1_sg U7784 ( .A(n6123), .X(n6497) );
  inv_x1_sg U7785 ( .A(n6123), .X(n6498) );
  inv_x1_sg U7786 ( .A(n7066), .X(n6499) );
  inv_x1_sg U7787 ( .A(n6499), .X(n6500) );
  inv_x1_sg U7788 ( .A(n6499), .X(n6501) );
  inv_x1_sg U7789 ( .A(n6499), .X(n6502) );
  inv_x1_sg U7790 ( .A(\update_mask_0/N31 ), .X(n6503) );
  inv_x1_sg U7791 ( .A(n6503), .X(n6504) );
  inv_x1_sg U7792 ( .A(n6503), .X(n6505) );
  inv_x1_sg U7793 ( .A(n6503), .X(n6506) );
  inv_x1_sg U7794 ( .A(\update_output_0/N32 ), .X(n6507) );
  inv_x1_sg U7795 ( .A(n6507), .X(n6508) );
  inv_x1_sg U7796 ( .A(n6507), .X(n6509) );
  inv_x1_sg U7797 ( .A(n6507), .X(n6510) );
  inv_x1_sg U7798 ( .A(n3742), .X(n6511) );
  inv_x1_sg U7799 ( .A(n3742), .X(n6512) );
  inv_x1_sg U7800 ( .A(n3742), .X(n6513) );
  inv_x1_sg U7801 ( .A(n6304), .X(n6514) );
  inv_x1_sg U7802 ( .A(n6091), .X(n6515) );
  inv_x1_sg U7803 ( .A(n6161), .X(n6516) );
  inv_x1_sg U7804 ( .A(n6516), .X(n6517) );
  inv_x1_sg U7805 ( .A(n6516), .X(n6518) );
  inv_x1_sg U7806 ( .A(n6516), .X(n6519) );
  inv_x1_sg U7807 ( .A(n6252), .X(n6520) );
  inv_x1_sg U7808 ( .A(n7357), .X(n6521) );
  inv_x1_sg U7809 ( .A(n6091), .X(n6522) );
  inv_x1_sg U7810 ( .A(n6465), .X(n6523) );
  inv_x1_sg U7811 ( .A(n6516), .X(n6524) );
  inv_x1_sg U7812 ( .A(n7355), .X(n6525) );
  inv_x1_sg U7813 ( .A(n7339), .X(n6526) );
  inv_x1_sg U7814 ( .A(n6090), .X(n6527) );
  inv_x1_sg U7815 ( .A(n6527), .X(n6528) );
  inv_x1_sg U7816 ( .A(n6527), .X(n6529) );
  inv_x1_sg U7817 ( .A(n6527), .X(n6530) );
  inv_x1_sg U7818 ( .A(n7357), .X(n6531) );
  inv_x1_sg U7819 ( .A(n6246), .X(n6532) );
  inv_x1_sg U7820 ( .A(n6087), .X(n6533) );
  inv_x1_sg U7821 ( .A(n6533), .X(n6534) );
  inv_x1_sg U7822 ( .A(n6533), .X(n6535) );
  inv_x1_sg U7823 ( .A(n6533), .X(n6536) );
  inv_x1_sg U7824 ( .A(n6300), .X(n6537) );
  inv_x1_sg U7825 ( .A(n7338), .X(n6538) );
  inv_x1_sg U7826 ( .A(n7460), .X(n6539) );
  inv_x1_sg U7827 ( .A(n6539), .X(n6540) );
  inv_x1_sg U7828 ( .A(n6539), .X(n6541) );
  inv_x1_sg U7829 ( .A(n6539), .X(n6542) );
  inv_x1_sg U7830 ( .A(n7340), .X(n6543) );
  inv_x1_sg U7831 ( .A(n6543), .X(n6544) );
  inv_x1_sg U7832 ( .A(n6543), .X(n6545) );
  inv_x1_sg U7833 ( .A(n6543), .X(n6546) );
  inv_x1_sg U7834 ( .A(n6543), .X(n6547) );
  inv_x1_sg U7835 ( .A(n3742), .X(n6548) );
  inv_x1_sg U7836 ( .A(n6548), .X(n6549) );
  inv_x1_sg U7837 ( .A(n6548), .X(n6550) );
  inv_x1_sg U7838 ( .A(n6548), .X(n6551) );
  inv_x1_sg U7839 ( .A(n6548), .X(n6552) );
  inv_x1_sg U7840 ( .A(n6788), .X(n6553) );
  inv_x1_sg U7841 ( .A(n6553), .X(n6554) );
  inv_x1_sg U7842 ( .A(n6553), .X(n6555) );
  inv_x1_sg U7843 ( .A(n6553), .X(n6556) );
  inv_x1_sg U7844 ( .A(n6553), .X(n6557) );
  inv_x1_sg U7845 ( .A(n7445), .X(n6558) );
  inv_x1_sg U7846 ( .A(n7445), .X(n6559) );
  inv_x1_sg U7847 ( .A(n7445), .X(n6560) );
  inv_x1_sg U7848 ( .A(n7445), .X(n6561) );
  inv_x1_sg U7849 ( .A(n7450), .X(n6562) );
  inv_x1_sg U7850 ( .A(n7450), .X(n6563) );
  inv_x1_sg U7851 ( .A(n7450), .X(n6564) );
  inv_x1_sg U7852 ( .A(n7450), .X(n6565) );
  inv_x1_sg U7853 ( .A(n7449), .X(n6566) );
  inv_x1_sg U7854 ( .A(n7449), .X(n6567) );
  inv_x1_sg U7855 ( .A(n7449), .X(n6568) );
  inv_x1_sg U7856 ( .A(n7449), .X(n6569) );
  inv_x1_sg U7857 ( .A(n7448), .X(n6570) );
  inv_x1_sg U7858 ( .A(n7448), .X(n6571) );
  inv_x1_sg U7859 ( .A(n7448), .X(n6572) );
  inv_x1_sg U7860 ( .A(n7448), .X(n6573) );
  inv_x1_sg U7861 ( .A(n4244), .X(n6574) );
  inv_x1_sg U7862 ( .A(n4244), .X(n6575) );
  inv_x1_sg U7863 ( .A(n4244), .X(n6576) );
  inv_x1_sg U7864 ( .A(n4244), .X(n6577) );
  inv_x1_sg U7865 ( .A(n4208), .X(n6578) );
  inv_x1_sg U7866 ( .A(n4208), .X(n6579) );
  inv_x1_sg U7867 ( .A(n4208), .X(n6580) );
  inv_x1_sg U7868 ( .A(n4208), .X(n6581) );
  inv_x1_sg U7869 ( .A(n6778), .X(n6582) );
  inv_x1_sg U7870 ( .A(n6582), .X(n6583) );
  inv_x1_sg U7871 ( .A(n6582), .X(n6584) );
  inv_x1_sg U7872 ( .A(n6582), .X(n6585) );
  inv_x1_sg U7873 ( .A(n6582), .X(n6586) );
  inv_x1_sg U7874 ( .A(n6773), .X(n6587) );
  inv_x1_sg U7875 ( .A(n6587), .X(n6588) );
  inv_x1_sg U7876 ( .A(n6587), .X(n6589) );
  inv_x1_sg U7877 ( .A(n6587), .X(n6590) );
  inv_x1_sg U7878 ( .A(n6587), .X(n6591) );
  inv_x1_sg U7879 ( .A(n6783), .X(n6592) );
  inv_x1_sg U7880 ( .A(n6592), .X(n6593) );
  inv_x1_sg U7881 ( .A(n6592), .X(n6594) );
  inv_x1_sg U7882 ( .A(n6592), .X(n6595) );
  inv_x1_sg U7883 ( .A(n6592), .X(n6596) );
  inv_x1_sg U7884 ( .A(n6813), .X(n6597) );
  inv_x1_sg U7885 ( .A(n6597), .X(n6598) );
  inv_x1_sg U7886 ( .A(n6597), .X(n6599) );
  inv_x1_sg U7887 ( .A(n6597), .X(n6600) );
  inv_x1_sg U7888 ( .A(n6597), .X(n6601) );
  inv_x1_sg U7889 ( .A(n6768), .X(n6602) );
  inv_x1_sg U7890 ( .A(n6602), .X(n6603) );
  inv_x1_sg U7891 ( .A(n6602), .X(n6604) );
  inv_x1_sg U7892 ( .A(n6602), .X(n6605) );
  inv_x1_sg U7893 ( .A(n6602), .X(n6606) );
  inv_x1_sg U7894 ( .A(n4130), .X(n6607) );
  inv_x1_sg U7895 ( .A(n4130), .X(n6608) );
  inv_x1_sg U7896 ( .A(n4130), .X(n6609) );
  inv_x1_sg U7897 ( .A(n4130), .X(n6610) );
  inv_x1_sg U7898 ( .A(n4172), .X(n6611) );
  inv_x1_sg U7899 ( .A(n4172), .X(n6612) );
  inv_x1_sg U7900 ( .A(n4172), .X(n6613) );
  inv_x1_sg U7901 ( .A(n4172), .X(n6614) );
  inv_x1_sg U7902 ( .A(n4280), .X(n6615) );
  inv_x1_sg U7903 ( .A(n4280), .X(n6616) );
  inv_x1_sg U7904 ( .A(n4280), .X(n6617) );
  inv_x1_sg U7905 ( .A(n4280), .X(n6618) );
  inv_x1_sg U7906 ( .A(n4316), .X(n6619) );
  inv_x1_sg U7907 ( .A(n4316), .X(n6620) );
  inv_x1_sg U7908 ( .A(n4316), .X(n6621) );
  inv_x1_sg U7909 ( .A(n4316), .X(n6622) );
  inv_x1_sg U7910 ( .A(n4388), .X(n6623) );
  inv_x1_sg U7911 ( .A(n4388), .X(n6624) );
  inv_x1_sg U7912 ( .A(n4388), .X(n6625) );
  inv_x1_sg U7913 ( .A(n4388), .X(n6626) );
  inv_x1_sg U7914 ( .A(n4424), .X(n6627) );
  inv_x1_sg U7915 ( .A(n4424), .X(n6628) );
  inv_x1_sg U7916 ( .A(n4424), .X(n6629) );
  inv_x1_sg U7917 ( .A(n4424), .X(n6630) );
  inv_x1_sg U7918 ( .A(n4460), .X(n6631) );
  inv_x1_sg U7919 ( .A(n4460), .X(n6632) );
  inv_x1_sg U7920 ( .A(n4460), .X(n6633) );
  inv_x1_sg U7921 ( .A(n4460), .X(n6634) );
  inv_x1_sg U7922 ( .A(n4496), .X(n6635) );
  inv_x1_sg U7923 ( .A(n4496), .X(n6636) );
  inv_x1_sg U7924 ( .A(n4496), .X(n6637) );
  inv_x1_sg U7925 ( .A(n4496), .X(n6638) );
  inv_x1_sg U7926 ( .A(n4568), .X(n6639) );
  inv_x1_sg U7927 ( .A(n4568), .X(n6640) );
  inv_x1_sg U7928 ( .A(n4568), .X(n6641) );
  inv_x1_sg U7929 ( .A(n4568), .X(n6642) );
  inv_x1_sg U7930 ( .A(n4676), .X(n6643) );
  inv_x1_sg U7931 ( .A(n4676), .X(n6644) );
  inv_x1_sg U7932 ( .A(n4676), .X(n6645) );
  inv_x1_sg U7933 ( .A(n4676), .X(n6646) );
  inv_x1_sg U7934 ( .A(n4712), .X(n6647) );
  inv_x1_sg U7935 ( .A(n4712), .X(n6648) );
  inv_x1_sg U7936 ( .A(n4712), .X(n6649) );
  inv_x1_sg U7937 ( .A(n4712), .X(n6650) );
  inv_x1_sg U7938 ( .A(n4748), .X(n6651) );
  inv_x1_sg U7939 ( .A(n4748), .X(n6652) );
  inv_x1_sg U7940 ( .A(n4748), .X(n6653) );
  inv_x1_sg U7941 ( .A(n4748), .X(n6654) );
  inv_x1_sg U7942 ( .A(n4784), .X(n6655) );
  inv_x1_sg U7943 ( .A(n4784), .X(n6656) );
  inv_x1_sg U7944 ( .A(n4784), .X(n6657) );
  inv_x1_sg U7945 ( .A(n4784), .X(n6658) );
  inv_x1_sg U7946 ( .A(n4822), .X(n6659) );
  inv_x1_sg U7947 ( .A(n4822), .X(n6660) );
  inv_x1_sg U7948 ( .A(n4822), .X(n6661) );
  inv_x1_sg U7949 ( .A(n4822), .X(n6662) );
  inv_x1_sg U7950 ( .A(n6793), .X(n6663) );
  inv_x1_sg U7951 ( .A(n6663), .X(n6664) );
  inv_x1_sg U7952 ( .A(n6663), .X(n6665) );
  inv_x1_sg U7953 ( .A(n6663), .X(n6666) );
  inv_x1_sg U7954 ( .A(n6663), .X(n6667) );
  inv_x1_sg U7955 ( .A(n6798), .X(n6668) );
  inv_x1_sg U7956 ( .A(n6668), .X(n6669) );
  inv_x1_sg U7957 ( .A(n6668), .X(n6670) );
  inv_x1_sg U7958 ( .A(n6668), .X(n6671) );
  inv_x1_sg U7959 ( .A(n6668), .X(n6672) );
  inv_x1_sg U7960 ( .A(n6803), .X(n6673) );
  inv_x1_sg U7961 ( .A(n6673), .X(n6674) );
  inv_x1_sg U7962 ( .A(n6673), .X(n6675) );
  inv_x1_sg U7963 ( .A(n6673), .X(n6676) );
  inv_x1_sg U7964 ( .A(n6673), .X(n6677) );
  inv_x1_sg U7965 ( .A(n6808), .X(n6678) );
  inv_x1_sg U7966 ( .A(n6678), .X(n6679) );
  inv_x1_sg U7967 ( .A(n6678), .X(n6680) );
  inv_x1_sg U7968 ( .A(n6678), .X(n6681) );
  inv_x1_sg U7969 ( .A(n6678), .X(n6682) );
  inv_x1_sg U7970 ( .A(n7420), .X(n6683) );
  inv_x1_sg U7971 ( .A(n6683), .X(n6684) );
  inv_x1_sg U7972 ( .A(n6683), .X(n6685) );
  inv_x1_sg U7973 ( .A(n6683), .X(n6686) );
  inv_x1_sg U7974 ( .A(n6823), .X(n6687) );
  inv_x1_sg U7975 ( .A(n6687), .X(n6688) );
  inv_x1_sg U7976 ( .A(n6687), .X(n6689) );
  inv_x1_sg U7977 ( .A(n6687), .X(n6690) );
  inv_x1_sg U7978 ( .A(n6687), .X(n6691) );
  inv_x1_sg U7979 ( .A(n6749), .X(n6692) );
  inv_x1_sg U7980 ( .A(n5936), .X(n6693) );
  inv_x1_sg U7981 ( .A(n6749), .X(n6694) );
  inv_x1_sg U7982 ( .A(n6764), .X(n6695) );
  inv_x1_sg U7983 ( .A(n5941), .X(n6696) );
  inv_x1_sg U7984 ( .A(n5941), .X(n6697) );
  inv_x1_sg U7985 ( .A(n5932), .X(n6698) );
  inv_x1_sg U7986 ( .A(n6698), .X(n6699) );
  inv_x1_sg U7987 ( .A(n6698), .X(n6700) );
  inv_x1_sg U7988 ( .A(n6698), .X(n6701) );
  inv_x1_sg U7989 ( .A(n6698), .X(n6702) );
  inv_x1_sg U7990 ( .A(n5937), .X(n6703) );
  inv_x1_sg U7991 ( .A(n6703), .X(n6704) );
  inv_x1_sg U7992 ( .A(n6703), .X(n6705) );
  inv_x1_sg U7993 ( .A(n6703), .X(n6706) );
  inv_x1_sg U7994 ( .A(n6703), .X(n6707) );
  inv_x1_sg U7995 ( .A(n5930), .X(n6708) );
  inv_x1_sg U7996 ( .A(n6708), .X(n6709) );
  inv_x1_sg U7997 ( .A(n6708), .X(n6710) );
  inv_x1_sg U7998 ( .A(n6708), .X(n6711) );
  inv_x1_sg U7999 ( .A(n6708), .X(n6712) );
  inv_x1_sg U8000 ( .A(n5928), .X(n6713) );
  inv_x1_sg U8001 ( .A(n6713), .X(n6714) );
  inv_x1_sg U8002 ( .A(n6713), .X(n6715) );
  inv_x1_sg U8003 ( .A(n6713), .X(n6716) );
  inv_x1_sg U8004 ( .A(n6713), .X(n6717) );
  inv_x1_sg U8005 ( .A(n5934), .X(n6718) );
  inv_x1_sg U8006 ( .A(n6718), .X(n6719) );
  inv_x1_sg U8007 ( .A(n6718), .X(n6720) );
  inv_x1_sg U8008 ( .A(n6718), .X(n6721) );
  inv_x1_sg U8009 ( .A(n6718), .X(n6722) );
  inv_x1_sg U8010 ( .A(n5939), .X(n6723) );
  inv_x1_sg U8011 ( .A(n6723), .X(n6724) );
  inv_x1_sg U8012 ( .A(n6723), .X(n6725) );
  inv_x1_sg U8013 ( .A(n6723), .X(n6726) );
  inv_x1_sg U8014 ( .A(n6723), .X(n6727) );
  inv_x1_sg U8015 ( .A(n735), .X(n6728) );
  inv_x1_sg U8016 ( .A(n6728), .X(n6729) );
  inv_x1_sg U8017 ( .A(n6728), .X(n6730) );
  inv_x1_sg U8018 ( .A(n6728), .X(n6731) );
  inv_x1_sg U8019 ( .A(n6728), .X(n6732) );
  inv_x1_sg U8020 ( .A(n750), .X(n6733) );
  inv_x1_sg U8021 ( .A(n6733), .X(n6734) );
  inv_x1_sg U8022 ( .A(n6733), .X(n6735) );
  inv_x1_sg U8023 ( .A(n6733), .X(n6736) );
  inv_x1_sg U8024 ( .A(n6733), .X(n6737) );
  inv_x1_sg U8025 ( .A(n749), .X(n6738) );
  inv_x1_sg U8026 ( .A(n6738), .X(n6739) );
  inv_x1_sg U8027 ( .A(n6738), .X(n6740) );
  inv_x1_sg U8028 ( .A(n6738), .X(n6741) );
  inv_x1_sg U8029 ( .A(n6738), .X(n6742) );
  inv_x1_sg U8030 ( .A(n746), .X(n6743) );
  inv_x1_sg U8031 ( .A(n6743), .X(n6744) );
  inv_x1_sg U8032 ( .A(n6743), .X(n6745) );
  inv_x1_sg U8033 ( .A(n6743), .X(n6746) );
  inv_x1_sg U8034 ( .A(n6743), .X(n6747) );
  inv_x1_sg U8035 ( .A(n739), .X(n6748) );
  inv_x1_sg U8036 ( .A(n6748), .X(n6749) );
  inv_x1_sg U8037 ( .A(n6748), .X(n6750) );
  inv_x1_sg U8038 ( .A(n5915), .X(n6751) );
  inv_x1_sg U8039 ( .A(n5914), .X(n6752) );
  inv_x1_sg U8040 ( .A(n744), .X(n6753) );
  inv_x1_sg U8041 ( .A(n6753), .X(n6754) );
  inv_x1_sg U8042 ( .A(n6753), .X(n6755) );
  inv_x1_sg U8043 ( .A(n6753), .X(n6756) );
  inv_x1_sg U8044 ( .A(n6753), .X(n6757) );
  inv_x1_sg U8045 ( .A(n736), .X(n6758) );
  inv_x1_sg U8046 ( .A(n6758), .X(n6759) );
  inv_x1_sg U8047 ( .A(n6758), .X(n6760) );
  inv_x1_sg U8048 ( .A(n6758), .X(n6761) );
  inv_x1_sg U8049 ( .A(n6758), .X(n6762) );
  inv_x1_sg U8050 ( .A(n740), .X(n6763) );
  inv_x1_sg U8051 ( .A(n6763), .X(n6764) );
  inv_x1_sg U8052 ( .A(n6763), .X(n6765) );
  inv_x1_sg U8053 ( .A(n5913), .X(n6766) );
  inv_x1_sg U8054 ( .A(n5912), .X(n6767) );
  inv_x1_sg U8055 ( .A(n748), .X(n6768) );
  inv_x1_sg U8056 ( .A(n6768), .X(n6769) );
  inv_x1_sg U8057 ( .A(n5942), .X(n6770) );
  inv_x1_sg U8058 ( .A(n5942), .X(n6771) );
  inv_x1_sg U8059 ( .A(n5942), .X(n6772) );
  inv_x1_sg U8060 ( .A(n745), .X(n6773) );
  inv_x1_sg U8061 ( .A(n6773), .X(n6774) );
  inv_x1_sg U8062 ( .A(n5944), .X(n6775) );
  inv_x1_sg U8063 ( .A(n5944), .X(n6776) );
  inv_x1_sg U8064 ( .A(n5944), .X(n6777) );
  inv_x1_sg U8065 ( .A(n742), .X(n6778) );
  inv_x1_sg U8066 ( .A(n6778), .X(n6779) );
  inv_x1_sg U8067 ( .A(n5946), .X(n6780) );
  inv_x1_sg U8068 ( .A(n5946), .X(n6781) );
  inv_x1_sg U8069 ( .A(n5946), .X(n6782) );
  inv_x1_sg U8070 ( .A(n753), .X(n6783) );
  inv_x1_sg U8071 ( .A(n6783), .X(n6784) );
  inv_x1_sg U8072 ( .A(n5948), .X(n6785) );
  inv_x1_sg U8073 ( .A(n5948), .X(n6786) );
  inv_x1_sg U8074 ( .A(n5948), .X(n6787) );
  inv_x1_sg U8075 ( .A(n755), .X(n6788) );
  inv_x1_sg U8076 ( .A(n6788), .X(n6789) );
  inv_x1_sg U8077 ( .A(n5950), .X(n6790) );
  inv_x1_sg U8078 ( .A(n5950), .X(n6791) );
  inv_x1_sg U8079 ( .A(n5950), .X(n6792) );
  inv_x1_sg U8080 ( .A(n747), .X(n6793) );
  inv_x1_sg U8081 ( .A(n6793), .X(n6794) );
  inv_x1_sg U8082 ( .A(n5952), .X(n6795) );
  inv_x1_sg U8083 ( .A(n5952), .X(n6796) );
  inv_x1_sg U8084 ( .A(n5952), .X(n6797) );
  inv_x1_sg U8085 ( .A(n752), .X(n6798) );
  inv_x1_sg U8086 ( .A(n6798), .X(n6799) );
  inv_x1_sg U8087 ( .A(n5954), .X(n6800) );
  inv_x1_sg U8088 ( .A(n5954), .X(n6801) );
  inv_x1_sg U8089 ( .A(n5954), .X(n6802) );
  inv_x1_sg U8090 ( .A(n751), .X(n6803) );
  inv_x1_sg U8091 ( .A(n6803), .X(n6804) );
  inv_x1_sg U8092 ( .A(n5956), .X(n6805) );
  inv_x1_sg U8093 ( .A(n5956), .X(n6806) );
  inv_x1_sg U8094 ( .A(n5956), .X(n6807) );
  inv_x1_sg U8095 ( .A(n738), .X(n6808) );
  inv_x1_sg U8096 ( .A(n6808), .X(n6809) );
  inv_x1_sg U8097 ( .A(n5958), .X(n6810) );
  inv_x1_sg U8098 ( .A(n5958), .X(n6811) );
  inv_x1_sg U8099 ( .A(n5958), .X(n6812) );
  inv_x1_sg U8100 ( .A(n741), .X(n6813) );
  inv_x1_sg U8101 ( .A(n6813), .X(n6814) );
  inv_x1_sg U8102 ( .A(n5960), .X(n6815) );
  inv_x1_sg U8103 ( .A(n5960), .X(n6816) );
  inv_x1_sg U8104 ( .A(n5960), .X(n6817) );
  inv_x1_sg U8105 ( .A(n743), .X(n6818) );
  inv_x1_sg U8106 ( .A(n6818), .X(n6819) );
  inv_x1_sg U8107 ( .A(n6818), .X(n6820) );
  inv_x1_sg U8108 ( .A(n6818), .X(n6821) );
  inv_x1_sg U8109 ( .A(n6818), .X(n6822) );
  inv_x1_sg U8110 ( .A(n737), .X(n6823) );
  inv_x1_sg U8111 ( .A(n6823), .X(n6824) );
  inv_x1_sg U8112 ( .A(n5964), .X(n6825) );
  inv_x1_sg U8113 ( .A(n5964), .X(n6826) );
  inv_x1_sg U8114 ( .A(n5964), .X(n6827) );
  inv_x1_sg U8115 ( .A(n7375), .X(n6828) );
  inv_x1_sg U8116 ( .A(n5966), .X(n6829) );
  inv_x1_sg U8117 ( .A(n6828), .X(n6830) );
  inv_x1_sg U8118 ( .A(n6828), .X(n6831) );
  inv_x1_sg U8119 ( .A(n6828), .X(n6832) );
  inv_x1_sg U8120 ( .A(n7422), .X(n6833) );
  inv_x1_sg U8121 ( .A(n6833), .X(n6834) );
  inv_x1_sg U8122 ( .A(n6833), .X(n6835) );
  inv_x1_sg U8123 ( .A(n6833), .X(n6836) );
  inv_x1_sg U8124 ( .A(n6833), .X(n6837) );
  inv_x1_sg U8125 ( .A(n7421), .X(n6838) );
  inv_x1_sg U8126 ( .A(n6838), .X(n6839) );
  inv_x1_sg U8127 ( .A(n6838), .X(n6840) );
  inv_x1_sg U8128 ( .A(n6838), .X(n6841) );
  inv_x1_sg U8129 ( .A(n6838), .X(n6842) );
  inv_x1_sg U8130 ( .A(n7388), .X(n6843) );
  inv_x1_sg U8131 ( .A(n6843), .X(n6844) );
  inv_x1_sg U8132 ( .A(n6843), .X(n6845) );
  inv_x1_sg U8133 ( .A(n6843), .X(n6846) );
  inv_x1_sg U8134 ( .A(n6843), .X(n6847) );
  inv_x1_sg U8135 ( .A(n7387), .X(n6848) );
  inv_x1_sg U8136 ( .A(n6848), .X(n6849) );
  inv_x1_sg U8137 ( .A(n6848), .X(n6850) );
  inv_x1_sg U8138 ( .A(n6848), .X(n6851) );
  inv_x1_sg U8139 ( .A(n6848), .X(n6852) );
  inv_x1_sg U8140 ( .A(n7386), .X(n6853) );
  inv_x1_sg U8141 ( .A(n6853), .X(n6854) );
  inv_x1_sg U8142 ( .A(n6853), .X(n6855) );
  inv_x1_sg U8143 ( .A(n6853), .X(n6856) );
  inv_x1_sg U8144 ( .A(n6853), .X(n6857) );
  inv_x1_sg U8145 ( .A(n7385), .X(n6858) );
  inv_x1_sg U8146 ( .A(n6858), .X(n6859) );
  inv_x1_sg U8147 ( .A(n6858), .X(n6860) );
  inv_x1_sg U8148 ( .A(n6858), .X(n6861) );
  inv_x1_sg U8149 ( .A(n6858), .X(n6862) );
  inv_x1_sg U8150 ( .A(n7384), .X(n6863) );
  inv_x1_sg U8151 ( .A(n6863), .X(n6864) );
  inv_x1_sg U8152 ( .A(n6863), .X(n6865) );
  inv_x1_sg U8153 ( .A(n6863), .X(n6866) );
  inv_x1_sg U8154 ( .A(n6863), .X(n6867) );
  inv_x1_sg U8155 ( .A(n7383), .X(n6868) );
  inv_x1_sg U8156 ( .A(n6868), .X(n6869) );
  inv_x1_sg U8157 ( .A(n6868), .X(n6870) );
  inv_x1_sg U8158 ( .A(n6868), .X(n6871) );
  inv_x1_sg U8159 ( .A(n6868), .X(n6872) );
  inv_x1_sg U8160 ( .A(n7382), .X(n6873) );
  inv_x1_sg U8161 ( .A(n6873), .X(n6874) );
  inv_x1_sg U8162 ( .A(n6873), .X(n6875) );
  inv_x1_sg U8163 ( .A(n6873), .X(n6876) );
  inv_x1_sg U8164 ( .A(n6873), .X(n6877) );
  inv_x1_sg U8165 ( .A(n7381), .X(n6878) );
  inv_x1_sg U8166 ( .A(n6878), .X(n6879) );
  inv_x1_sg U8167 ( .A(n6878), .X(n6880) );
  inv_x1_sg U8168 ( .A(n6878), .X(n6881) );
  inv_x1_sg U8169 ( .A(n6878), .X(n6882) );
  inv_x1_sg U8170 ( .A(n7380), .X(n6883) );
  inv_x1_sg U8171 ( .A(n6883), .X(n6884) );
  inv_x1_sg U8172 ( .A(n6883), .X(n6885) );
  inv_x1_sg U8173 ( .A(n6883), .X(n6886) );
  inv_x1_sg U8174 ( .A(n6883), .X(n6887) );
  inv_x1_sg U8175 ( .A(n7379), .X(n6888) );
  inv_x1_sg U8176 ( .A(n6888), .X(n6889) );
  inv_x1_sg U8177 ( .A(n6888), .X(n6890) );
  inv_x1_sg U8178 ( .A(n6888), .X(n6891) );
  inv_x1_sg U8179 ( .A(n6888), .X(n6892) );
  inv_x1_sg U8180 ( .A(n6912), .X(n6893) );
  inv_x1_sg U8181 ( .A(n6912), .X(n6894) );
  inv_x1_sg U8182 ( .A(n6918), .X(n6895) );
  inv_x1_sg U8183 ( .A(n6912), .X(n6896) );
  inv_x1_sg U8184 ( .A(n7378), .X(n6897) );
  inv_x1_sg U8185 ( .A(n6897), .X(n6898) );
  inv_x1_sg U8186 ( .A(n6897), .X(n6899) );
  inv_x1_sg U8187 ( .A(n6897), .X(n6900) );
  inv_x1_sg U8188 ( .A(n6897), .X(n6901) );
  inv_x1_sg U8189 ( .A(n7377), .X(n6902) );
  inv_x1_sg U8190 ( .A(n6902), .X(n6903) );
  inv_x1_sg U8191 ( .A(n6902), .X(n6904) );
  inv_x1_sg U8192 ( .A(n6902), .X(n6905) );
  inv_x1_sg U8193 ( .A(n6902), .X(n6906) );
  inv_x1_sg U8194 ( .A(n7376), .X(n6907) );
  inv_x1_sg U8195 ( .A(n6907), .X(n6908) );
  inv_x1_sg U8196 ( .A(n6907), .X(n6909) );
  inv_x1_sg U8197 ( .A(n6907), .X(n6910) );
  inv_x1_sg U8198 ( .A(n6907), .X(n6911) );
  nand_x1_sg U8199 ( .A(n4849), .B(n6332), .X(n6912) );
  inv_x1_sg U8200 ( .A(n6912), .X(n6913) );
  inv_x1_sg U8201 ( .A(n6913), .X(n6914) );
  inv_x1_sg U8202 ( .A(n6913), .X(n6915) );
  inv_x1_sg U8203 ( .A(n4146), .X(n6916) );
  inv_x1_sg U8204 ( .A(n6916), .X(n6917) );
  inv_x1_sg U8205 ( .A(n6916), .X(n6918) );
  inv_x1_sg U8206 ( .A(n6916), .X(n6919) );
  inv_x1_sg U8207 ( .A(n6916), .X(n6920) );
  inv_x1_sg U8208 ( .A(n7467), .X(n6921) );
  inv_x1_sg U8209 ( .A(n7385), .X(n6922) );
  inv_x1_sg U8210 ( .A(n6921), .X(n6923) );
  inv_x1_sg U8211 ( .A(n6921), .X(n6924) );
  inv_x1_sg U8212 ( .A(n6921), .X(n6925) );
  inv_x1_sg U8213 ( .A(n7470), .X(n6926) );
  inv_x1_sg U8214 ( .A(n7386), .X(n6927) );
  inv_x1_sg U8215 ( .A(n6926), .X(n6928) );
  inv_x1_sg U8216 ( .A(n6926), .X(n6929) );
  inv_x1_sg U8217 ( .A(n6926), .X(n6930) );
  inv_x1_sg U8218 ( .A(n7475), .X(n6931) );
  inv_x1_sg U8219 ( .A(n6931), .X(n6932) );
  inv_x1_sg U8220 ( .A(n6931), .X(n6933) );
  inv_x1_sg U8221 ( .A(n6931), .X(n6934) );
  inv_x1_sg U8222 ( .A(n6931), .X(n6935) );
  inv_x1_sg U8223 ( .A(n7472), .X(n6936) );
  inv_x1_sg U8224 ( .A(n7383), .X(n6937) );
  inv_x1_sg U8225 ( .A(n6936), .X(n6938) );
  inv_x1_sg U8226 ( .A(n6936), .X(n6939) );
  inv_x1_sg U8227 ( .A(n6936), .X(n6940) );
  inv_x1_sg U8228 ( .A(n7466), .X(n6941) );
  inv_x1_sg U8229 ( .A(n7387), .X(n6942) );
  inv_x1_sg U8230 ( .A(n6941), .X(n6943) );
  inv_x1_sg U8231 ( .A(n6941), .X(n6944) );
  inv_x1_sg U8232 ( .A(n6941), .X(n6945) );
  inv_x1_sg U8233 ( .A(n7469), .X(n6946) );
  inv_x1_sg U8234 ( .A(n7376), .X(n6947) );
  inv_x1_sg U8235 ( .A(n6946), .X(n6948) );
  inv_x1_sg U8236 ( .A(n6946), .X(n6949) );
  inv_x1_sg U8237 ( .A(n6946), .X(n6950) );
  inv_x1_sg U8238 ( .A(n7474), .X(n6951) );
  inv_x1_sg U8239 ( .A(n7382), .X(n6952) );
  inv_x1_sg U8240 ( .A(n6951), .X(n6953) );
  inv_x1_sg U8241 ( .A(n6951), .X(n6954) );
  inv_x1_sg U8242 ( .A(n6951), .X(n6955) );
  inv_x1_sg U8243 ( .A(n7471), .X(n6956) );
  inv_x1_sg U8244 ( .A(n7377), .X(n6957) );
  inv_x1_sg U8245 ( .A(n6956), .X(n6958) );
  inv_x1_sg U8246 ( .A(n6956), .X(n6959) );
  inv_x1_sg U8247 ( .A(n6956), .X(n6960) );
  inv_x1_sg U8248 ( .A(n7465), .X(n6961) );
  inv_x1_sg U8249 ( .A(n7381), .X(n6962) );
  inv_x1_sg U8250 ( .A(n6961), .X(n6963) );
  inv_x1_sg U8251 ( .A(n6961), .X(n6964) );
  inv_x1_sg U8252 ( .A(n6961), .X(n6965) );
  inv_x1_sg U8253 ( .A(n3613), .X(n6966) );
  inv_x1_sg U8254 ( .A(n7378), .X(n6967) );
  inv_x1_sg U8255 ( .A(n6966), .X(n6968) );
  inv_x1_sg U8256 ( .A(n6966), .X(n6969) );
  inv_x1_sg U8257 ( .A(n6966), .X(n6970) );
  inv_x1_sg U8258 ( .A(n7476), .X(n6971) );
  inv_x1_sg U8259 ( .A(n7388), .X(n6972) );
  inv_x1_sg U8260 ( .A(n6971), .X(n6973) );
  inv_x1_sg U8261 ( .A(n6971), .X(n6974) );
  inv_x1_sg U8262 ( .A(n6971), .X(n6975) );
  inv_x1_sg U8263 ( .A(n7468), .X(n6976) );
  inv_x1_sg U8264 ( .A(n7384), .X(n6977) );
  inv_x1_sg U8265 ( .A(n6976), .X(n6978) );
  inv_x1_sg U8266 ( .A(n6976), .X(n6979) );
  inv_x1_sg U8267 ( .A(n6976), .X(n6980) );
  inv_x1_sg U8268 ( .A(n7477), .X(n6981) );
  inv_x1_sg U8269 ( .A(n7379), .X(n6982) );
  inv_x1_sg U8270 ( .A(n6981), .X(n6983) );
  inv_x1_sg U8271 ( .A(n6981), .X(n6984) );
  inv_x1_sg U8272 ( .A(n6981), .X(n6985) );
  inv_x1_sg U8273 ( .A(n7464), .X(n6986) );
  inv_x1_sg U8274 ( .A(n7421), .X(n6987) );
  inv_x1_sg U8275 ( .A(n6986), .X(n6988) );
  inv_x1_sg U8276 ( .A(n6986), .X(n6989) );
  inv_x1_sg U8277 ( .A(n6986), .X(n6990) );
  inv_x1_sg U8278 ( .A(n3656), .X(n6991) );
  inv_x1_sg U8279 ( .A(n7422), .X(n6992) );
  inv_x1_sg U8280 ( .A(n6991), .X(n6993) );
  inv_x1_sg U8281 ( .A(n6991), .X(n6994) );
  inv_x1_sg U8282 ( .A(n6991), .X(n6995) );
  inv_x1_sg U8283 ( .A(n7458), .X(n6996) );
  inv_x1_sg U8284 ( .A(n7458), .X(n6997) );
  inv_x1_sg U8285 ( .A(n7458), .X(n6998) );
  inv_x1_sg U8286 ( .A(n6997), .X(n6999) );
  inv_x1_sg U8287 ( .A(n6263), .X(n7000) );
  inv_x1_sg U8288 ( .A(n6996), .X(n7001) );
  inv_x1_sg U8289 ( .A(n6996), .X(n7002) );
  inv_x1_sg U8290 ( .A(n6996), .X(n7003) );
  inv_x1_sg U8291 ( .A(n6997), .X(n7004) );
  inv_x1_sg U8292 ( .A(n6997), .X(n7005) );
  inv_x1_sg U8293 ( .A(n6997), .X(n7006) );
  inv_x1_sg U8294 ( .A(n6998), .X(n7007) );
  inv_x1_sg U8295 ( .A(n6998), .X(n7008) );
  inv_x1_sg U8296 ( .A(n6998), .X(n7009) );
  inv_x1_sg U8297 ( .A(n7417), .X(n7010) );
  inv_x1_sg U8298 ( .A(n6117), .X(n7011) );
  inv_x1_sg U8299 ( .A(n7010), .X(n7012) );
  inv_x1_sg U8300 ( .A(n6117), .X(n7013) );
  inv_x1_sg U8301 ( .A(n7010), .X(n7014) );
  inv_x1_sg U8302 ( .A(n5985), .X(n7015) );
  inv_x1_sg U8303 ( .A(n6120), .X(n7016) );
  inv_x1_sg U8304 ( .A(n7015), .X(n7017) );
  inv_x1_sg U8305 ( .A(n6120), .X(n7018) );
  inv_x1_sg U8306 ( .A(n7015), .X(n7019) );
  inv_x1_sg U8307 ( .A(n6152), .X(n7020) );
  inv_x1_sg U8308 ( .A(n6244), .X(n7021) );
  inv_x1_sg U8309 ( .A(n5926), .X(n7022) );
  inv_x1_sg U8310 ( .A(n5926), .X(n7023) );
  inv_x1_sg U8311 ( .A(n6289), .X(n7024) );
  inv_x1_sg U8312 ( .A(n6289), .X(n7025) );
  inv_x1_sg U8313 ( .A(n5925), .X(n7026) );
  inv_x1_sg U8314 ( .A(n5925), .X(n7027) );
  inv_x1_sg U8315 ( .A(n6285), .X(n7028) );
  inv_x1_sg U8316 ( .A(n6285), .X(n7029) );
  inv_x1_sg U8317 ( .A(n6147), .X(n7030) );
  inv_x1_sg U8318 ( .A(n6243), .X(n7031) );
  inv_x1_sg U8319 ( .A(n7330), .X(n7032) );
  inv_x1_sg U8320 ( .A(n5924), .X(n7033) );
  inv_x1_sg U8321 ( .A(n5924), .X(n7034) );
  inv_x1_sg U8322 ( .A(n6280), .X(n7035) );
  inv_x1_sg U8323 ( .A(n6280), .X(n7036) );
  inv_x1_sg U8324 ( .A(n7329), .X(n7037) );
  inv_x1_sg U8325 ( .A(n5923), .X(n7038) );
  inv_x1_sg U8326 ( .A(n5923), .X(n7039) );
  inv_x1_sg U8327 ( .A(n6274), .X(n7040) );
  inv_x1_sg U8328 ( .A(n6274), .X(n7041) );
  inv_x1_sg U8329 ( .A(n6142), .X(n7042) );
  inv_x1_sg U8330 ( .A(n6242), .X(n7043) );
  inv_x1_sg U8331 ( .A(n5922), .X(n7044) );
  inv_x1_sg U8332 ( .A(n5922), .X(n7045) );
  inv_x1_sg U8333 ( .A(n6269), .X(n7046) );
  inv_x1_sg U8334 ( .A(n6269), .X(n7047) );
  inv_x1_sg U8335 ( .A(n7325), .X(n7048) );
  inv_x1_sg U8336 ( .A(n6265), .X(n7049) );
  inv_x1_sg U8337 ( .A(n6266), .X(n7050) );
  inv_x1_sg U8338 ( .A(n6266), .X(n7051) );
  inv_x1_sg U8339 ( .A(n6147), .X(n7052) );
  inv_x1_sg U8340 ( .A(n1521), .X(n7053) );
  inv_x1_sg U8341 ( .A(n7053), .X(n7054) );
  inv_x1_sg U8342 ( .A(n6163), .X(n7055) );
  inv_x1_sg U8343 ( .A(n6163), .X(n7056) );
  inv_x1_sg U8344 ( .A(n7053), .X(n7057) );
  inv_x1_sg U8345 ( .A(n1520), .X(n7058) );
  inv_x1_sg U8346 ( .A(n7058), .X(n7059) );
  inv_x1_sg U8347 ( .A(n6166), .X(n7060) );
  inv_x1_sg U8348 ( .A(n6166), .X(n7061) );
  inv_x1_sg U8349 ( .A(n7058), .X(n7062) );
  inv_x1_sg U8350 ( .A(n4154), .X(n7063) );
  inv_x1_sg U8351 ( .A(n7063), .X(n7064) );
  inv_x1_sg U8352 ( .A(n7063), .X(n7065) );
  inv_x1_sg U8353 ( .A(n7063), .X(n7066) );
  inv_x1_sg U8354 ( .A(n6123), .X(n7067) );
  nand_x1_sg U8355 ( .A(n1433), .B(n6369), .X(n7068) );
  inv_x1_sg U8356 ( .A(n7068), .X(n7069) );
  inv_x1_sg U8357 ( .A(n7069), .X(n7070) );
  inv_x1_sg U8358 ( .A(n7069), .X(n7071) );
  inv_x1_sg U8359 ( .A(n7069), .X(n7072) );
  inv_x1_sg U8360 ( .A(n7069), .X(n7073) );
  inv_x1_sg U8361 ( .A(n7071), .X(n7074) );
  inv_x1_sg U8362 ( .A(n7074), .X(n7075) );
  inv_x1_sg U8363 ( .A(n7074), .X(n7076) );
  inv_x1_sg U8364 ( .A(n7074), .X(n7077) );
  inv_x1_sg U8365 ( .A(n7074), .X(n7078) );
  inv_x1_sg U8366 ( .A(n7068), .X(n7079) );
  inv_x1_sg U8367 ( .A(n7079), .X(n7080) );
  inv_x1_sg U8368 ( .A(n7079), .X(n7081) );
  inv_x1_sg U8369 ( .A(n792), .X(n7082) );
  inv_x1_sg U8370 ( .A(n6006), .X(n7083) );
  inv_x1_sg U8371 ( .A(n6006), .X(n7084) );
  inv_x1_sg U8372 ( .A(n7082), .X(n7085) );
  inv_x1_sg U8373 ( .A(n7082), .X(n7086) );
  inv_x1_sg U8374 ( .A(n1534), .X(n7087) );
  inv_x1_sg U8375 ( .A(n7087), .X(n7088) );
  inv_x1_sg U8376 ( .A(n6172), .X(n7089) );
  inv_x1_sg U8377 ( .A(n6172), .X(n7090) );
  inv_x1_sg U8378 ( .A(n7087), .X(n7091) );
  inv_x1_sg U8379 ( .A(n1524), .X(n7092) );
  inv_x1_sg U8380 ( .A(n7092), .X(n7093) );
  inv_x1_sg U8381 ( .A(n6175), .X(n7094) );
  inv_x1_sg U8382 ( .A(n6175), .X(n7095) );
  inv_x1_sg U8383 ( .A(n7092), .X(n7096) );
  inv_x1_sg U8384 ( .A(n1526), .X(n7097) );
  inv_x1_sg U8385 ( .A(n7097), .X(n7098) );
  inv_x1_sg U8386 ( .A(n6178), .X(n7099) );
  inv_x1_sg U8387 ( .A(n6178), .X(n7100) );
  inv_x1_sg U8388 ( .A(n7097), .X(n7101) );
  inv_x1_sg U8389 ( .A(n734), .X(n7102) );
  inv_x1_sg U8390 ( .A(n7102), .X(n7103) );
  inv_x1_sg U8391 ( .A(n6181), .X(n7104) );
  inv_x1_sg U8392 ( .A(n6181), .X(n7105) );
  inv_x1_sg U8393 ( .A(n7102), .X(n7106) );
  inv_x1_sg U8394 ( .A(n772), .X(n7107) );
  inv_x1_sg U8395 ( .A(n7107), .X(n7108) );
  inv_x1_sg U8396 ( .A(n6184), .X(n7109) );
  inv_x1_sg U8397 ( .A(n6184), .X(n7110) );
  inv_x1_sg U8398 ( .A(n7107), .X(n7111) );
  inv_x1_sg U8399 ( .A(n766), .X(n7112) );
  inv_x1_sg U8400 ( .A(n7112), .X(n7113) );
  inv_x1_sg U8401 ( .A(n6187), .X(n7114) );
  inv_x1_sg U8402 ( .A(n6187), .X(n7115) );
  inv_x1_sg U8403 ( .A(n7112), .X(n7116) );
  inv_x1_sg U8404 ( .A(n759), .X(n7117) );
  inv_x1_sg U8405 ( .A(n7117), .X(n7118) );
  inv_x1_sg U8406 ( .A(n6190), .X(n7119) );
  inv_x1_sg U8407 ( .A(n6190), .X(n7120) );
  inv_x1_sg U8408 ( .A(n7117), .X(n7121) );
  inv_x1_sg U8409 ( .A(n4151), .X(n7122) );
  inv_x1_sg U8410 ( .A(n7122), .X(n7123) );
  inv_x1_sg U8411 ( .A(n6030), .X(n7124) );
  inv_x1_sg U8412 ( .A(n7122), .X(n7125) );
  inv_x1_sg U8413 ( .A(n6030), .X(n7126) );
  nor_x1_sg U8414 ( .A(n3954), .B(n6510), .X(n7127) );
  inv_x1_sg U8415 ( .A(n7127), .X(n7128) );
  inv_x1_sg U8416 ( .A(n7128), .X(n7129) );
  inv_x1_sg U8417 ( .A(n7128), .X(n7130) );
  inv_x1_sg U8418 ( .A(n7128), .X(n7131) );
  inv_x1_sg U8419 ( .A(n7128), .X(n7132) );
  inv_x1_sg U8420 ( .A(n7127), .X(n7133) );
  inv_x1_sg U8421 ( .A(n7133), .X(n7134) );
  inv_x1_sg U8422 ( .A(n7133), .X(n7135) );
  inv_x1_sg U8423 ( .A(n7133), .X(n7136) );
  inv_x1_sg U8424 ( .A(n7133), .X(n7137) );
  inv_x1_sg U8425 ( .A(n7127), .X(n7138) );
  inv_x1_sg U8426 ( .A(n7138), .X(n7139) );
  inv_x1_sg U8427 ( .A(n7138), .X(n7140) );
  inv_x1_sg U8428 ( .A(n7138), .X(n7141) );
  inv_x1_sg U8429 ( .A(n7138), .X(n7142) );
  inv_x1_sg U8430 ( .A(n806), .X(n7143) );
  inv_x1_sg U8431 ( .A(n6033), .X(n7144) );
  inv_x1_sg U8432 ( .A(n6033), .X(n7145) );
  inv_x1_sg U8433 ( .A(n6322), .X(n7146) );
  inv_x1_sg U8434 ( .A(n6322), .X(n7147) );
  nand_x1_sg U8435 ( .A(n1433), .B(n6458), .X(n7148) );
  inv_x1_sg U8436 ( .A(n7148), .X(n7149) );
  inv_x1_sg U8437 ( .A(n7149), .X(n7150) );
  inv_x1_sg U8438 ( .A(n7149), .X(n7151) );
  inv_x1_sg U8439 ( .A(n7149), .X(n7152) );
  inv_x1_sg U8440 ( .A(n7149), .X(n7153) );
  inv_x1_sg U8441 ( .A(n7148), .X(n7154) );
  inv_x1_sg U8442 ( .A(n7154), .X(n7155) );
  inv_x1_sg U8443 ( .A(n7154), .X(n7156) );
  inv_x1_sg U8444 ( .A(n7154), .X(n7157) );
  inv_x1_sg U8445 ( .A(n7148), .X(n7158) );
  inv_x1_sg U8446 ( .A(n7158), .X(n7159) );
  inv_x1_sg U8447 ( .A(n7158), .X(n7160) );
  inv_x1_sg U8448 ( .A(n7158), .X(n7161) );
  inv_x1_sg U8449 ( .A(n7158), .X(n7162) );
  inv_x1_sg U8450 ( .A(n770), .X(n7163) );
  inv_x1_sg U8451 ( .A(n7163), .X(n7164) );
  inv_x1_sg U8452 ( .A(n6196), .X(n7165) );
  inv_x1_sg U8453 ( .A(n6196), .X(n7166) );
  inv_x1_sg U8454 ( .A(n7163), .X(n7167) );
  inv_x1_sg U8455 ( .A(n768), .X(n7168) );
  inv_x1_sg U8456 ( .A(n7168), .X(n7169) );
  inv_x1_sg U8457 ( .A(n6199), .X(n7170) );
  inv_x1_sg U8458 ( .A(n6199), .X(n7171) );
  inv_x1_sg U8459 ( .A(n7168), .X(n7172) );
  inv_x1_sg U8460 ( .A(n758), .X(n7173) );
  inv_x1_sg U8461 ( .A(n7173), .X(n7174) );
  inv_x1_sg U8462 ( .A(n6202), .X(n7175) );
  inv_x1_sg U8463 ( .A(n6202), .X(n7176) );
  inv_x1_sg U8464 ( .A(n7173), .X(n7177) );
  inv_x1_sg U8465 ( .A(n754), .X(n7178) );
  inv_x1_sg U8466 ( .A(n7178), .X(n7179) );
  inv_x1_sg U8467 ( .A(n6205), .X(n7180) );
  inv_x1_sg U8468 ( .A(n6205), .X(n7181) );
  inv_x1_sg U8469 ( .A(n7178), .X(n7182) );
  inv_x1_sg U8470 ( .A(n776), .X(n7183) );
  inv_x1_sg U8471 ( .A(n7183), .X(n7184) );
  inv_x1_sg U8472 ( .A(n6208), .X(n7185) );
  inv_x1_sg U8473 ( .A(n6208), .X(n7186) );
  inv_x1_sg U8474 ( .A(n7183), .X(n7187) );
  inv_x1_sg U8475 ( .A(n775), .X(n7188) );
  inv_x1_sg U8476 ( .A(n7188), .X(n7189) );
  inv_x1_sg U8477 ( .A(n6211), .X(n7190) );
  inv_x1_sg U8478 ( .A(n6211), .X(n7191) );
  inv_x1_sg U8479 ( .A(n7188), .X(n7192) );
  inv_x1_sg U8480 ( .A(n774), .X(n7193) );
  inv_x1_sg U8481 ( .A(n7193), .X(n7194) );
  inv_x1_sg U8482 ( .A(n6214), .X(n7195) );
  inv_x1_sg U8483 ( .A(n6214), .X(n7196) );
  inv_x1_sg U8484 ( .A(n7193), .X(n7197) );
  inv_x1_sg U8485 ( .A(n764), .X(n7198) );
  inv_x1_sg U8486 ( .A(n7198), .X(n7199) );
  inv_x1_sg U8487 ( .A(n6217), .X(n7200) );
  inv_x1_sg U8488 ( .A(n6217), .X(n7201) );
  inv_x1_sg U8489 ( .A(n7198), .X(n7202) );
  inv_x1_sg U8490 ( .A(n763), .X(n7203) );
  inv_x1_sg U8491 ( .A(n7203), .X(n7204) );
  inv_x1_sg U8492 ( .A(n6220), .X(n7205) );
  inv_x1_sg U8493 ( .A(n6220), .X(n7206) );
  inv_x1_sg U8494 ( .A(n7203), .X(n7207) );
  inv_x1_sg U8495 ( .A(n762), .X(n7208) );
  inv_x1_sg U8496 ( .A(n7208), .X(n7209) );
  inv_x1_sg U8497 ( .A(n6223), .X(n7210) );
  inv_x1_sg U8498 ( .A(n6223), .X(n7211) );
  inv_x1_sg U8499 ( .A(n7208), .X(n7212) );
  inv_x1_sg U8500 ( .A(n769), .X(n7213) );
  inv_x1_sg U8501 ( .A(n7213), .X(n7214) );
  inv_x1_sg U8502 ( .A(n6226), .X(n7215) );
  inv_x1_sg U8503 ( .A(n6226), .X(n7216) );
  inv_x1_sg U8504 ( .A(n7213), .X(n7217) );
  inv_x1_sg U8505 ( .A(n757), .X(n7218) );
  inv_x1_sg U8506 ( .A(n7218), .X(n7219) );
  inv_x1_sg U8507 ( .A(n6229), .X(n7220) );
  inv_x1_sg U8508 ( .A(n6229), .X(n7221) );
  inv_x1_sg U8509 ( .A(n7218), .X(n7222) );
  inv_x1_sg U8510 ( .A(n7444), .X(n7223) );
  inv_x1_sg U8511 ( .A(n7223), .X(n7224) );
  inv_x1_sg U8512 ( .A(n6232), .X(n7225) );
  inv_x1_sg U8513 ( .A(n6232), .X(n7226) );
  inv_x1_sg U8514 ( .A(n7223), .X(n7227) );
  inv_x1_sg U8515 ( .A(n7461), .X(n7228) );
  inv_x1_sg U8516 ( .A(n7228), .X(n7229) );
  inv_x1_sg U8517 ( .A(n7228), .X(n7230) );
  inv_x1_sg U8518 ( .A(n7228), .X(n7231) );
  inv_x1_sg U8519 ( .A(n7228), .X(n7232) );
  inv_x1_sg U8520 ( .A(n7461), .X(n7233) );
  inv_x1_sg U8521 ( .A(n7233), .X(n7234) );
  inv_x1_sg U8522 ( .A(n7233), .X(n7235) );
  inv_x1_sg U8523 ( .A(n7233), .X(n7236) );
  inv_x1_sg U8524 ( .A(n7461), .X(n7237) );
  inv_x1_sg U8525 ( .A(n7237), .X(n7238) );
  inv_x1_sg U8526 ( .A(n7237), .X(n7239) );
  inv_x1_sg U8527 ( .A(n7237), .X(n7240) );
  inv_x1_sg U8528 ( .A(n4147), .X(n7241) );
  inv_x1_sg U8529 ( .A(n7243), .X(n7242) );
  inv_x1_sg U8530 ( .A(n4147), .X(n7243) );
  inv_x1_sg U8531 ( .A(n7248), .X(n7244) );
  inv_x1_sg U8532 ( .A(n7241), .X(n7245) );
  inv_x1_sg U8533 ( .A(n7241), .X(n7246) );
  inv_x1_sg U8534 ( .A(n7243), .X(n7247) );
  inv_x1_sg U8535 ( .A(n4147), .X(n7248) );
  inv_x1_sg U8536 ( .A(n7248), .X(n7249) );
  inv_x1_sg U8537 ( .A(n7243), .X(n7250) );
  inv_x1_sg U8538 ( .A(n7248), .X(n7251) );
  inv_x1_sg U8539 ( .A(n7241), .X(n7252) );
  inv_x1_sg U8540 ( .A(n7241), .X(n7253) );
  inv_x1_sg U8541 ( .A(n4140), .X(n7254) );
  inv_x1_sg U8542 ( .A(n6075), .X(n7255) );
  inv_x1_sg U8543 ( .A(n6075), .X(n7256) );
  inv_x1_sg U8544 ( .A(n7254), .X(n7257) );
  inv_x1_sg U8545 ( .A(n6235), .X(n7258) );
  inv_x1_sg U8546 ( .A(n7462), .X(n7259) );
  inv_x1_sg U8547 ( .A(n7259), .X(n7260) );
  inv_x1_sg U8548 ( .A(n6078), .X(n7261) );
  inv_x1_sg U8549 ( .A(n7259), .X(n7262) );
  inv_x1_sg U8550 ( .A(n7259), .X(n7263) );
  inv_x1_sg U8551 ( .A(n6078), .X(n7264) );
  inv_x1_sg U8552 ( .A(n7462), .X(n7265) );
  inv_x1_sg U8553 ( .A(n7265), .X(n7266) );
  inv_x1_sg U8554 ( .A(n7265), .X(n7267) );
  inv_x1_sg U8555 ( .A(n7265), .X(n7268) );
  inv_x1_sg U8556 ( .A(n7265), .X(n7269) );
  inv_x1_sg U8557 ( .A(n7259), .X(n7270) );
  inv_x1_sg U8558 ( .A(n6078), .X(n7271) );
  inv_x1_sg U8559 ( .A(n7418), .X(n7272) );
  inv_x1_sg U8560 ( .A(n7272), .X(n7273) );
  inv_x1_sg U8561 ( .A(n7272), .X(n7274) );
  inv_x1_sg U8562 ( .A(n6124), .X(n7275) );
  inv_x1_sg U8563 ( .A(n7272), .X(n7276) );
  inv_x1_sg U8564 ( .A(n7416), .X(n7277) );
  inv_x1_sg U8565 ( .A(n7277), .X(n7278) );
  inv_x1_sg U8566 ( .A(n7277), .X(n7279) );
  inv_x1_sg U8567 ( .A(n7277), .X(n7280) );
  inv_x1_sg U8568 ( .A(n6127), .X(n7281) );
  inv_x1_sg U8569 ( .A(n7415), .X(n7282) );
  inv_x1_sg U8570 ( .A(n7282), .X(n7283) );
  inv_x1_sg U8571 ( .A(n7282), .X(n7284) );
  inv_x1_sg U8572 ( .A(n6130), .X(n7285) );
  inv_x1_sg U8573 ( .A(n6130), .X(n7286) );
  nand_x1_sg U8574 ( .A(n1438), .B(n6369), .X(n7287) );
  inv_x1_sg U8575 ( .A(n7287), .X(n7288) );
  inv_x1_sg U8576 ( .A(n7288), .X(n7289) );
  inv_x1_sg U8577 ( .A(n7288), .X(n7290) );
  inv_x1_sg U8578 ( .A(n7288), .X(n7291) );
  inv_x1_sg U8579 ( .A(n7287), .X(n7292) );
  inv_x1_sg U8580 ( .A(n7292), .X(n7293) );
  inv_x1_sg U8581 ( .A(n7292), .X(n7294) );
  inv_x1_sg U8582 ( .A(n7292), .X(n7295) );
  inv_x1_sg U8583 ( .A(n7292), .X(n7296) );
  inv_x1_sg U8584 ( .A(n7287), .X(n7297) );
  inv_x1_sg U8585 ( .A(n7297), .X(n7298) );
  inv_x1_sg U8586 ( .A(n7297), .X(n7299) );
  inv_x1_sg U8587 ( .A(n7297), .X(n7300) );
  inv_x1_sg U8588 ( .A(n7297), .X(n7301) );
  inv_x1_sg U8589 ( .A(n5625), .X(n7302) );
  inv_x1_sg U8590 ( .A(n7302), .X(n7303) );
  inv_x1_sg U8591 ( .A(n6133), .X(n7304) );
  inv_x1_sg U8592 ( .A(n6133), .X(n7305) );
  inv_x1_sg U8593 ( .A(n6133), .X(n7306) );
  inv_x1_sg U8594 ( .A(n5611), .X(n7307) );
  inv_x1_sg U8595 ( .A(n7307), .X(n7308) );
  inv_x1_sg U8596 ( .A(n7307), .X(n7309) );
  inv_x1_sg U8597 ( .A(n6136), .X(n7310) );
  inv_x1_sg U8598 ( .A(n6136), .X(n7311) );
  inv_x1_sg U8599 ( .A(\update_output_0/N34 ), .X(n7312) );
  inv_x1_sg U8600 ( .A(n7312), .X(n7313) );
  inv_x1_sg U8601 ( .A(n6139), .X(n7314) );
  inv_x1_sg U8602 ( .A(n7312), .X(n7315) );
  inv_x1_sg U8603 ( .A(n6139), .X(n7316) );
  inv_x1_sg U8604 ( .A(\update_output_0/N30 ), .X(n7317) );
  inv_x1_sg U8605 ( .A(n7317), .X(n7318) );
  inv_x1_sg U8606 ( .A(n7317), .X(n7319) );
  inv_x1_sg U8607 ( .A(n7317), .X(n7320) );
  inv_x1_sg U8608 ( .A(n6239), .X(n7321) );
  inv_x1_sg U8609 ( .A(n6239), .X(n7322) );
  nor_x1_sg U8610 ( .A(n6544), .B(reset), .X(n7323) );
  inv_x1_sg U8611 ( .A(n6151), .X(n7324) );
  inv_x1_sg U8612 ( .A(n6242), .X(n7325) );
  inv_x1_sg U8613 ( .A(n7324), .X(n7326) );
  inv_x1_sg U8614 ( .A(n7324), .X(n7327) );
  inv_x1_sg U8615 ( .A(n7323), .X(n7328) );
  inv_x1_sg U8616 ( .A(n6243), .X(n7329) );
  inv_x1_sg U8617 ( .A(n7328), .X(n7330) );
  inv_x1_sg U8618 ( .A(n7328), .X(n7331) );
  inv_x1_sg U8619 ( .A(n7463), .X(n7332) );
  inv_x1_sg U8620 ( .A(n6244), .X(n7333) );
  inv_x1_sg U8621 ( .A(n7332), .X(n7334) );
  inv_x1_sg U8622 ( .A(n7332), .X(n7335) );
  nor_x1_sg U8623 ( .A(n4885), .B(reset), .X(n7336) );
  inv_x1_sg U8624 ( .A(n7336), .X(n7337) );
  inv_x1_sg U8625 ( .A(n7336), .X(n7338) );
  inv_x1_sg U8626 ( .A(n6162), .X(n7339) );
  inv_x1_sg U8627 ( .A(n7337), .X(n7340) );
  inv_x1_sg U8628 ( .A(n6299), .X(n7341) );
  inv_x1_sg U8629 ( .A(n6086), .X(n7342) );
  inv_x1_sg U8630 ( .A(n6246), .X(n7343) );
  inv_x1_sg U8631 ( .A(n7337), .X(n7344) );
  inv_x1_sg U8632 ( .A(n7338), .X(n7345) );
  inv_x1_sg U8633 ( .A(n6245), .X(n7346) );
  inv_x1_sg U8634 ( .A(n6245), .X(n7347) );
  inv_x1_sg U8635 ( .A(n6086), .X(n7348) );
  inv_x1_sg U8636 ( .A(n7338), .X(n7349) );
  inv_x1_sg U8637 ( .A(n7339), .X(n7350) );
  inv_x1_sg U8638 ( .A(n6299), .X(n7351) );
  inv_x1_sg U8639 ( .A(n6300), .X(n7352) );
  inv_x1_sg U8640 ( .A(n7338), .X(n7353) );
  inv_x1_sg U8641 ( .A(n6300), .X(n7354) );
  inv_x1_sg U8642 ( .A(n4892), .X(n7355) );
  inv_x1_sg U8643 ( .A(n5917), .X(n7356) );
  inv_x1_sg U8644 ( .A(n5917), .X(n7357) );
  inv_x1_sg U8645 ( .A(n7356), .X(n7358) );
  inv_x1_sg U8646 ( .A(n7357), .X(n7359) );
  inv_x1_sg U8647 ( .A(n7355), .X(n7360) );
  inv_x1_sg U8648 ( .A(n7339), .X(n7361) );
  inv_x1_sg U8649 ( .A(n7356), .X(n7362) );
  inv_x1_sg U8650 ( .A(n6089), .X(n7363) );
  inv_x1_sg U8651 ( .A(n6251), .X(n7364) );
  inv_x1_sg U8652 ( .A(n6304), .X(n7365) );
  inv_x1_sg U8653 ( .A(n6084), .X(n7366) );
  inv_x1_sg U8654 ( .A(n6089), .X(n7367) );
  inv_x1_sg U8655 ( .A(n6299), .X(n7368) );
  inv_x1_sg U8656 ( .A(n6303), .X(n7369) );
  inv_x1_sg U8657 ( .A(n6251), .X(n7370) );
  inv_x1_sg U8658 ( .A(n6245), .X(n7371) );
  inv_x1_sg U8659 ( .A(n7356), .X(n7372) );
  nor_x1_sg U8660 ( .A(n6160), .B(reset), .X(n4892) );
  nor_x1_sg U8661 ( .A(n1445), .B(n7399), .X(n7462) );
  nor_x1_sg U8662 ( .A(n3954), .B(n7414), .X(n4140) );
  inv_x1_sg U8663 ( .A(n3452), .X(n7373) );
  inv_x1_sg U8664 ( .A(\update_output_0/n6096 ), .X(n7374) );
  inv_x1_sg U8665 ( .A(n3436), .X(n7375) );
  inv_x1_sg U8666 ( .A(n7469), .X(n7376) );
  inv_x1_sg U8667 ( .A(n7471), .X(n7377) );
  inv_x1_sg U8668 ( .A(n3613), .X(n7378) );
  inv_x1_sg U8669 ( .A(n7477), .X(n7379) );
  inv_x1_sg U8670 ( .A(n7475), .X(n7380) );
  inv_x1_sg U8671 ( .A(n7465), .X(n7381) );
  inv_x1_sg U8672 ( .A(n7474), .X(n7382) );
  inv_x1_sg U8673 ( .A(n7472), .X(n7383) );
  inv_x1_sg U8674 ( .A(n7468), .X(n7384) );
  inv_x1_sg U8675 ( .A(n7467), .X(n7385) );
  inv_x1_sg U8676 ( .A(n7470), .X(n7386) );
  inv_x1_sg U8677 ( .A(n7466), .X(n7387) );
  inv_x1_sg U8678 ( .A(n7476), .X(n7388) );
  inv_x1_sg U8679 ( .A(\update_mask_0/N23 ), .X(n7389) );
  inv_x1_sg U8680 ( .A(n6540), .X(n7390) );
  inv_x1_sg U8681 ( .A(n4855), .X(n7391) );
  inv_x1_sg U8682 ( .A(n6348), .X(n7392) );
  inv_x1_sg U8683 ( .A(n6354), .X(n7393) );
  inv_x1_sg U8684 ( .A(\update_mask_0/N28 ), .X(n7394) );
  inv_x1_sg U8685 ( .A(\update_output_0/N28 ), .X(n7395) );
  inv_x1_sg U8686 ( .A(\update_mask_0/N30 ), .X(n7396) );
  inv_x1_sg U8687 ( .A(n3479), .X(n7397) );
  inv_x1_sg U8688 ( .A(n3524), .X(n7398) );
  inv_x1_sg U8689 ( .A(\update_output_0/N29 ), .X(n7399) );
  inv_x1_sg U8690 ( .A(n6333), .X(n7400) );
  inv_x1_sg U8691 ( .A(\update_output_0/N33 ), .X(n7401) );
  inv_x1_sg U8692 ( .A(\mask_state[0] ), .X(n7402) );
  inv_x1_sg U8693 ( .A(\update_mask_0/N25 ), .X(n7403) );
  inv_x1_sg U8694 ( .A(n7007), .X(n7404) );
  inv_x1_sg U8695 ( .A(\update_mask_0/N26 ), .X(n7405) );
  inv_x1_sg U8696 ( .A(n6335), .X(n7406) );
  inv_x1_sg U8697 ( .A(\update_mask_0/N27 ), .X(n7407) );
  inv_x1_sg U8698 ( .A(n4821), .X(n7408) );
  inv_x1_sg U8699 ( .A(n1468), .X(n7409) );
  inv_x1_sg U8700 ( .A(n1500), .X(n7410) );
  inv_x1_sg U8701 ( .A(n1493), .X(n7411) );
  inv_x1_sg U8702 ( .A(n1482), .X(n7412) );
  inv_x1_sg U8703 ( .A(n6377), .X(n7413) );
  inv_x1_sg U8704 ( .A(n6508), .X(n7414) );
  inv_x1_sg U8705 ( .A(n3997), .X(n7415) );
  inv_x1_sg U8706 ( .A(n3453), .X(n7416) );
  inv_x1_sg U8707 ( .A(n6505), .X(n7417) );
  inv_x1_sg U8708 ( .A(n3466), .X(n7418) );
  inv_x1_sg U8709 ( .A(n4872), .X(n7419) );
  inv_x1_sg U8710 ( .A(n6819), .X(n7420) );
  inv_x1_sg U8711 ( .A(n7464), .X(n7421) );
  inv_x1_sg U8712 ( .A(n3656), .X(n7422) );
  nand_x1_sg U8713 ( .A(n3451), .B(n7321), .X(n7423) );
  nand_x4_sg U8714 ( .A(n5632), .B(n6159), .X(n7424) );
  nand_x2_sg U8715 ( .A(n6498), .B(n5680), .X(n4311) );
  nand_x2_sg U8716 ( .A(n6031), .B(n5739), .X(n4310) );
  nand_x2_sg U8717 ( .A(n2190), .B(n9227), .X(n4884) );
  nand_x2_sg U8718 ( .A(n2191), .B(n6330), .X(n2190) );
  nand_x4_sg U8719 ( .A(n1442), .B(n6313), .X(n3453) );
  nor_x1_sg U8720 ( .A(n6546), .B(reset), .X(n7463) );
  nand_x4_sg U8721 ( .A(n2254), .B(n6309), .X(n7446) );
  inv_x1_sg U8722 ( .A(n6372), .X(n7457) );
  inv_x1_sg U8723 ( .A(n6375), .X(n7456) );
  nand_x1_sg U8724 ( .A(n2180), .B(n7396), .X(n5625) );
  nand_x4_sg U8725 ( .A(n2252), .B(n6367), .X(n7442) );
  nand_x1_sg U8726 ( .A(n4849), .B(n7400), .X(n4147) );
  nand_x4_sg U8727 ( .A(n2262), .B(\update_mask_0/N24 ), .X(n7460) );
  nand_x4_sg U8728 ( .A(n1151), .B(n1152), .X(n736) );
  nand_x4_sg U8729 ( .A(n2189), .B(n6310), .X(n1470) );
  nand_x4_sg U8730 ( .A(n5635), .B(\mask_state[0] ), .X(n4872) );
  nand_x1_sg U8731 ( .A(n6831), .B(n4820), .X(n7464) );
  nand_x1_sg U8732 ( .A(n6831), .B(n3781), .X(n3742) );
  nand_x1_sg U8733 ( .A(n1438), .B(n6458), .X(n7461) );
  nand_x4_sg U8734 ( .A(n2261), .B(n6366), .X(n1449) );
  nand_x4_sg U8735 ( .A(n2251), .B(n6367), .X(n1459) );
  inv_x1_sg U8736 ( .A(n2051), .X(n7425) );
  inv_x1_sg U8737 ( .A(n2133), .X(n7426) );
  inv_x1_sg U8738 ( .A(n1965), .X(n7427) );
  inv_x1_sg U8739 ( .A(n2035), .X(n7428) );
  inv_x1_sg U8740 ( .A(n1883), .X(n7429) );
  inv_x1_sg U8741 ( .A(n1951), .X(n7430) );
  inv_x1_sg U8742 ( .A(n1795), .X(n7431) );
  inv_x1_sg U8743 ( .A(n1867), .X(n7432) );
  inv_x1_sg U8744 ( .A(n1697), .X(n7433) );
  inv_x1_sg U8745 ( .A(n1713), .X(n7434) );
  inv_x1_sg U8746 ( .A(n1613), .X(n7435) );
  inv_x1_sg U8747 ( .A(n1627), .X(n7436) );
  inv_x1_sg U8748 ( .A(n1527), .X(n7437) );
  inv_x1_sg U8749 ( .A(n1545), .X(n7438) );
  nor_x1_sg U8750 ( .A(n1114), .B(n1115), .X(n778) );
  nor_x1_sg U8751 ( .A(n1429), .B(n1430), .X(n1428) );
  nor_x1_sg U8752 ( .A(n1350), .B(n1351), .X(n1349) );
  nor_x1_sg U8753 ( .A(n1389), .B(n1390), .X(n1380) );
  nor_x1_sg U8754 ( .A(n1293), .B(n1294), .X(n1284) );
  nor_x1_sg U8755 ( .A(n1325), .B(n1326), .X(n1316) );
  nor_x1_sg U8756 ( .A(n1226), .B(n1227), .X(n1217) );
  nor_x1_sg U8757 ( .A(n1277), .B(n1278), .X(n1267) );
  nor_x1_sg U8758 ( .A(n1138), .B(n1139), .X(n1137) );
  nor_x1_sg U8759 ( .A(n1187), .B(n1188), .X(n1186) );
  nor_x1_sg U8760 ( .A(n1069), .B(n1070), .X(n1068) );
  nor_x1_sg U8761 ( .A(n1086), .B(n1087), .X(n1085) );
  nor_x1_sg U8762 ( .A(n990), .B(n991), .X(n989) );
  nor_x1_sg U8763 ( .A(n1029), .B(n1030), .X(n1020) );
  nor_x1_sg U8764 ( .A(n923), .B(n924), .X(n922) );
  nor_x1_sg U8765 ( .A(n973), .B(n974), .X(n972) );
  nor_x1_sg U8766 ( .A(n874), .B(n875), .X(n873) );
  nor_x1_sg U8767 ( .A(n906), .B(n907), .X(n905) );
  nor_x1_sg U8768 ( .A(n810), .B(n811), .X(n809) );
  nor_x1_sg U8769 ( .A(n842), .B(n843), .X(n841) );
  nor_x1_sg U8770 ( .A(n2106), .B(n2107), .X(n2105) );
  nor_x1_sg U8771 ( .A(n2023), .B(n2024), .X(n2022) );
  nor_x1_sg U8772 ( .A(n1855), .B(n1856), .X(n1854) );
  nor_x1_sg U8773 ( .A(n1938), .B(n1939), .X(n1937) );
  nor_x1_sg U8774 ( .A(n1768), .B(n1769), .X(n1767) );
  nor_x1_sg U8775 ( .A(n1685), .B(n1686), .X(n1684) );
  nor_x1_sg U8776 ( .A(n1511), .B(n1512), .X(n1510) );
  nor_x1_sg U8777 ( .A(n1600), .B(n1601), .X(n1599) );
  nand_x8_sg U8778 ( .A(n9227), .B(n4862), .X(n3436) );
  inv_x16_sg U8779 ( .A(reset), .X(n9227) );
  nor_x1_sg U8780 ( .A(n2140), .B(n2141), .X(n2106) );
  nor_x1_sg U8781 ( .A(n1802), .B(n1803), .X(n1768) );
  inv_x1_sg U8782 ( .A(n3464), .X(n7439) );
  inv_x1_sg U8783 ( .A(\update_mask_0/N29 ), .X(n7440) );
  inv_x1_sg U8784 ( .A(n6381), .X(n7441) );
  nand_x1_sg U8785 ( .A(n1498), .B(n1466), .X(n7443) );
  nand_x1_sg U8786 ( .A(n5626), .B(n6101), .X(n7444) );
  nand_x2_sg U8787 ( .A(n7000), .B(n4569), .X(n4568) );
  nand_x2_sg U8788 ( .A(n7009), .B(n4677), .X(n4676) );
  nand_x2_sg U8789 ( .A(n7003), .B(n4281), .X(n4280) );
  nand_x2_sg U8790 ( .A(n7001), .B(n4389), .X(n4388) );
  nand_x2_sg U8791 ( .A(n7009), .B(n4823), .X(n4822) );
  nand_x2_sg U8792 ( .A(n7008), .B(n4425), .X(n4424) );
  nand_x2_sg U8793 ( .A(n7009), .B(n4173), .X(n4172) );
  nand_x1_sg U8794 ( .A(n5967), .B(n3522), .X(n7477) );
  nand_x1_sg U8795 ( .A(n7003), .B(n4641), .X(n7445) );
  inv_x8_sg U8796 ( .A(output_taken), .X(n7447) );
  inv_x16_sg U8797 ( .A(output_taken), .X(n9234) );
  nand_x2_sg U8798 ( .A(n6999), .B(n4353), .X(n7448) );
  nand_x2_sg U8799 ( .A(n7006), .B(n4533), .X(n7449) );
  nand_x2_sg U8800 ( .A(n7008), .B(n4605), .X(n7450) );
  nand_x1_sg U8801 ( .A(n5967), .B(n3996), .X(n7468) );
  nand_x1_sg U8802 ( .A(n3782), .B(n9226), .X(n7451) );
  nand_x2_sg U8803 ( .A(n7007), .B(n4497), .X(n4496) );
  nand_x2_sg U8804 ( .A(n7008), .B(n4245), .X(n4244) );
  nand_x2_sg U8805 ( .A(n7009), .B(n4317), .X(n4316) );
  nand_x1_sg U8806 ( .A(n6831), .B(n3566), .X(n7476) );
  nand_x1_sg U8807 ( .A(n3826), .B(n7408), .X(n4820) );
  nand_x1_sg U8808 ( .A(n5597), .B(n6309), .X(n1446) );
  nand_x1_sg U8809 ( .A(n6829), .B(n3652), .X(n3613) );
  nand_x1_sg U8810 ( .A(n6830), .B(n4124), .X(n7465) );
  nand_x1_sg U8811 ( .A(n6832), .B(n3868), .X(n7471) );
  nand_x1_sg U8812 ( .A(n6832), .B(n3738), .X(n7474) );
  inv_x1_sg U8813 ( .A(n7424), .X(n7452) );
  nand_x1_sg U8814 ( .A(n1465), .B(n5920), .X(n7453) );
  nand_x1_sg U8815 ( .A(n1491), .B(n1466), .X(n7454) );
  nand_x1_sg U8816 ( .A(n1480), .B(n5920), .X(n7455) );
  nand_x1_sg U8817 ( .A(n6830), .B(n3953), .X(n7469) );
  nand_x1_sg U8818 ( .A(n6832), .B(n4082), .X(n7466) );
  nand_x1_sg U8819 ( .A(n6830), .B(n3825), .X(n7472) );
  nor_x1_sg U8820 ( .A(n5918), .B(n5966), .X(n7458) );
  nand_x1_sg U8821 ( .A(n2265), .B(n6098), .X(n1455) );
  inv_x8_sg U8822 ( .A(input_ready), .X(n9233) );
  nand_x1_sg U8823 ( .A(n2265), .B(n7389), .X(n1452) );
  nand_x1_sg U8824 ( .A(n6829), .B(n3609), .X(n7475) );
  nand_x4_sg U8825 ( .A(n825), .B(n826), .X(n824) );
  nand_x4_sg U8826 ( .A(n787), .B(n788), .X(n786) );
  nand_x4_sg U8827 ( .A(n956), .B(n957), .X(n955) );
  nand_x4_sg U8828 ( .A(n1003), .B(n1004), .X(n986) );
  nand_x4_sg U8829 ( .A(n1168), .B(n1169), .X(n1151) );
  nand_x4_sg U8830 ( .A(n1153), .B(n1154), .X(n1152) );
  nand_x4_sg U8831 ( .A(n1121), .B(n1122), .X(n1120) );
  nand_x1_sg U8832 ( .A(n1777), .B(n8918), .X(n1773) );
  inv_x1_sg U8833 ( .A(n1542), .X(n8915) );
  inv_x1_sg U8834 ( .A(n1523), .X(n8939) );
  inv_x1_sg U8835 ( .A(n1610), .X(n8916) );
  inv_x1_sg U8836 ( .A(n1625), .X(n8941) );
  inv_x1_sg U8837 ( .A(n1710), .X(n8917) );
  inv_x1_sg U8838 ( .A(n1695), .X(n8944) );
  nand_x1_sg U8839 ( .A(n2115), .B(n8922), .X(n2111) );
  inv_x1_sg U8840 ( .A(n1880), .X(n8919) );
  inv_x1_sg U8841 ( .A(n1865), .X(n8949) );
  inv_x1_sg U8842 ( .A(n1948), .X(n8920) );
  inv_x1_sg U8843 ( .A(n1963), .X(n8951) );
  inv_x1_sg U8844 ( .A(n2048), .X(n8921) );
  inv_x1_sg U8845 ( .A(n2033), .X(n8954) );
  nor_x1_sg U8846 ( .A(n1844), .B(n1845), .X(n1843) );
  nand_x2_sg U8847 ( .A(n1821), .B(n1822), .X(n1820) );
  nand_x2_sg U8848 ( .A(n1826), .B(n1827), .X(n1819) );
  nand_x2_sg U8849 ( .A(n1836), .B(n1837), .X(n1835) );
  inv_x1_sg U8850 ( .A(n1793), .X(n8946) );
  nand_x2_sg U8851 ( .A(n1796), .B(n1797), .X(n1795) );
  nand_x2_sg U8852 ( .A(n1804), .B(n1805), .X(n1803) );
  nand_x2_sg U8853 ( .A(n1809), .B(n1810), .X(n1802) );
  inv_x1_sg U8854 ( .A(n1781), .X(n8959) );
  nand_x2_sg U8855 ( .A(n1782), .B(n1783), .X(n1781) );
  nand_x2_sg U8856 ( .A(n1546), .B(n1547), .X(n1545) );
  nand_x2_sg U8857 ( .A(n1528), .B(n1529), .X(n1527) );
  nor_x1_sg U8858 ( .A(n1568), .B(n1569), .X(n1567) );
  nand_x1_sg U8859 ( .A(n1576), .B(n1577), .X(n1568) );
  nor_x1_sg U8860 ( .A(n1578), .B(n1579), .X(n1577) );
  nand_x2_sg U8861 ( .A(n1590), .B(n1591), .X(n1583) );
  nand_x2_sg U8862 ( .A(n1585), .B(n1586), .X(n1584) );
  nor_x1_sg U8863 ( .A(n1551), .B(n1552), .X(n1511) );
  nand_x1_sg U8864 ( .A(n1559), .B(n1560), .X(n1551) );
  nor_x1_sg U8865 ( .A(n1561), .B(n1562), .X(n1560) );
  nand_x2_sg U8866 ( .A(n1614), .B(n1615), .X(n1613) );
  nand_x2_sg U8867 ( .A(n1628), .B(n1629), .X(n1627) );
  nor_x1_sg U8868 ( .A(n1651), .B(n1652), .X(n1650) );
  nand_x1_sg U8869 ( .A(n1658), .B(n1659), .X(n1651) );
  nand_x2_sg U8870 ( .A(n1668), .B(n1669), .X(n1667) );
  nor_x1_sg U8871 ( .A(n1676), .B(n1677), .X(n1675) );
  nor_x1_sg U8872 ( .A(n1634), .B(n1635), .X(n1600) );
  nand_x1_sg U8873 ( .A(n1641), .B(n1642), .X(n1634) );
  nand_x2_sg U8874 ( .A(n1714), .B(n1715), .X(n1713) );
  nand_x2_sg U8875 ( .A(n1698), .B(n1699), .X(n1697) );
  nor_x1_sg U8876 ( .A(n1736), .B(n1737), .X(n1735) );
  nand_x1_sg U8877 ( .A(n1744), .B(n1745), .X(n1736) );
  nor_x1_sg U8878 ( .A(n1746), .B(n1747), .X(n1745) );
  nand_x2_sg U8879 ( .A(n1758), .B(n1759), .X(n1751) );
  nand_x2_sg U8880 ( .A(n1753), .B(n1754), .X(n1752) );
  nor_x1_sg U8881 ( .A(n1719), .B(n1720), .X(n1685) );
  nand_x1_sg U8882 ( .A(n1727), .B(n1728), .X(n1719) );
  nor_x1_sg U8883 ( .A(n1729), .B(n1730), .X(n1728) );
  nor_x1_sg U8884 ( .A(n2183), .B(n2184), .X(n2182) );
  nand_x2_sg U8885 ( .A(n2159), .B(n2160), .X(n2158) );
  nand_x2_sg U8886 ( .A(n2164), .B(n2165), .X(n2157) );
  nand_x2_sg U8887 ( .A(n2174), .B(n2175), .X(n2173) );
  inv_x1_sg U8888 ( .A(n2131), .X(n8956) );
  nand_x2_sg U8889 ( .A(n2134), .B(n2135), .X(n2133) );
  nand_x2_sg U8890 ( .A(n2142), .B(n2143), .X(n2141) );
  nand_x2_sg U8891 ( .A(n2147), .B(n2148), .X(n2140) );
  inv_x1_sg U8892 ( .A(n2119), .X(n8960) );
  nand_x2_sg U8893 ( .A(n2120), .B(n2121), .X(n2119) );
  nand_x2_sg U8894 ( .A(n1884), .B(n1885), .X(n1883) );
  nand_x2_sg U8895 ( .A(n1868), .B(n1869), .X(n1867) );
  nor_x1_sg U8896 ( .A(n1906), .B(n1907), .X(n1905) );
  nand_x1_sg U8897 ( .A(n1914), .B(n1915), .X(n1906) );
  nor_x1_sg U8898 ( .A(n1916), .B(n1917), .X(n1915) );
  nand_x2_sg U8899 ( .A(n1928), .B(n1929), .X(n1921) );
  nand_x2_sg U8900 ( .A(n1923), .B(n1924), .X(n1922) );
  nor_x1_sg U8901 ( .A(n1889), .B(n1890), .X(n1855) );
  nand_x1_sg U8902 ( .A(n1897), .B(n1898), .X(n1889) );
  nor_x1_sg U8903 ( .A(n1899), .B(n1900), .X(n1898) );
  nand_x2_sg U8904 ( .A(n1952), .B(n1953), .X(n1951) );
  nand_x2_sg U8905 ( .A(n1966), .B(n1967), .X(n1965) );
  nor_x1_sg U8906 ( .A(n1989), .B(n1990), .X(n1988) );
  nand_x1_sg U8907 ( .A(n1996), .B(n1997), .X(n1989) );
  nand_x2_sg U8908 ( .A(n2006), .B(n2007), .X(n2005) );
  nor_x1_sg U8909 ( .A(n2014), .B(n2015), .X(n2013) );
  nor_x1_sg U8910 ( .A(n1972), .B(n1973), .X(n1938) );
  nand_x1_sg U8911 ( .A(n1979), .B(n1980), .X(n1972) );
  nand_x2_sg U8912 ( .A(n2052), .B(n2053), .X(n2051) );
  nand_x2_sg U8913 ( .A(n2036), .B(n2037), .X(n2035) );
  nor_x1_sg U8914 ( .A(n2074), .B(n2075), .X(n2073) );
  nand_x1_sg U8915 ( .A(n2082), .B(n2083), .X(n2074) );
  nor_x1_sg U8916 ( .A(n2084), .B(n2085), .X(n2083) );
  nand_x2_sg U8917 ( .A(n2096), .B(n2097), .X(n2089) );
  nand_x2_sg U8918 ( .A(n2091), .B(n2092), .X(n2090) );
  nor_x1_sg U8919 ( .A(n2057), .B(n2058), .X(n2023) );
  nand_x1_sg U8920 ( .A(n2065), .B(n2066), .X(n2057) );
  nor_x1_sg U8921 ( .A(n2067), .B(n2068), .X(n2066) );
  nand_x1_sg U8922 ( .A(n6005), .B(n5805), .X(n4477) );
  nand_x1_sg U8923 ( .A(n7066), .B(n5796), .X(n4455) );
  nand_x1_sg U8924 ( .A(n6393), .B(n5858), .X(n4411) );
  nand_x1_sg U8925 ( .A(n6424), .B(n5735), .X(n4418) );
  nand_x1_sg U8926 ( .A(n7131), .B(n5818), .X(n4399) );
  nand_x1_sg U8927 ( .A(n6394), .B(n5734), .X(n4397) );
  nand_x1_sg U8928 ( .A(n7132), .B(n5877), .X(n4376) );
  nand_x1_sg U8929 ( .A(n6031), .B(n5845), .X(n4382) );
  nand_x1_sg U8930 ( .A(n7256), .B(n5852), .X(n4361) );
  nand_x1_sg U8931 ( .A(n7131), .B(n5864), .X(n4340) );
  nand_x1_sg U8932 ( .A(n7126), .B(n5759), .X(n4346) );
  nand_x1_sg U8933 ( .A(n7255), .B(n5865), .X(n4325) );
  nand_x1_sg U8934 ( .A(n7139), .B(n5760), .X(n4304) );
  inv_x2_sg U8935 ( .A(\i_im[6][0] ), .X(n9062) );
  inv_x1_sg U8936 ( .A(n1426), .X(n9002) );
  inv_x2_sg U8937 ( .A(\i_im[6][1] ), .X(n9063) );
  inv_x1_sg U8938 ( .A(n1135), .X(n9003) );
  inv_x2_sg U8939 ( .A(\i_im[15][1] ), .X(n9203) );
  inv_x2_sg U8940 ( .A(\i_im[6][2] ), .X(n9064) );
  inv_x1_sg U8941 ( .A(n1167), .X(n9004) );
  inv_x1_sg U8942 ( .A(n1237), .X(n9105) );
  inv_x2_sg U8943 ( .A(\i_im[13][3] ), .X(n9165) );
  inv_x2_sg U8944 ( .A(\i_im[7][3] ), .X(n9085) );
  inv_x2_sg U8945 ( .A(\i_im[6][4] ), .X(n9066) );
  inv_x1_sg U8946 ( .A(n1199), .X(n9006) );
  inv_x2_sg U8947 ( .A(\i_im[4][4] ), .X(n9026) );
  inv_x2_sg U8948 ( .A(\i_im[15][4] ), .X(n9206) );
  inv_x2_sg U8949 ( .A(\i_im[6][5] ), .X(n9067) );
  inv_x1_sg U8950 ( .A(n1266), .X(n9007) );
  inv_x1_sg U8951 ( .A(n1304), .X(n9108) );
  inv_x2_sg U8952 ( .A(\i_im[13][6] ), .X(n9168) );
  inv_x2_sg U8953 ( .A(\i_im[7][6] ), .X(n9088) );
  inv_x1_sg U8954 ( .A(n1336), .X(n9109) );
  inv_x2_sg U8955 ( .A(\i_im[13][7] ), .X(n9169) );
  inv_x2_sg U8956 ( .A(\i_im[7][7] ), .X(n9089) );
  inv_x2_sg U8957 ( .A(\i_im[6][8] ), .X(n9070) );
  inv_x1_sg U8958 ( .A(n1362), .X(n9010) );
  inv_x2_sg U8959 ( .A(\i_im[4][8] ), .X(n9030) );
  inv_x2_sg U8960 ( .A(\i_im[7][9] ), .X(n9091) );
  inv_x2_sg U8961 ( .A(\i_im[6][10] ), .X(n9072) );
  inv_x1_sg U8962 ( .A(n1002), .X(n9012) );
  nand_x1_sg U8963 ( .A(n6324), .B(n9052), .X(n1001) );
  inv_x2_sg U8964 ( .A(\i_im[5][10] ), .X(n9052) );
  inv_x2_sg U8965 ( .A(\i_im[4][10] ), .X(n9032) );
  inv_x2_sg U8966 ( .A(\i_im[15][10] ), .X(n9212) );
  inv_x2_sg U8967 ( .A(\i_im[15][11] ), .X(n9213) );
  inv_x1_sg U8968 ( .A(n1040), .X(n9113) );
  nand_x1_sg U8969 ( .A(n6422), .B(n9173), .X(n1039) );
  inv_x2_sg U8970 ( .A(\i_im[13][11] ), .X(n9173) );
  inv_x2_sg U8971 ( .A(\i_im[5][11] ), .X(n9053) );
  inv_x2_sg U8972 ( .A(\i_im[7][11] ), .X(n9093) );
  nand_x1_sg U8973 ( .A(n7264), .B(n9073), .X(n1032) );
  inv_x2_sg U8974 ( .A(\i_im[6][11] ), .X(n9073) );
  inv_x2_sg U8975 ( .A(\i_im[6][12] ), .X(n9074) );
  inv_x1_sg U8976 ( .A(n970), .X(n9014) );
  nand_x1_sg U8977 ( .A(n7146), .B(n9054), .X(n969) );
  inv_x2_sg U8978 ( .A(\i_im[5][12] ), .X(n9054) );
  inv_x2_sg U8979 ( .A(\i_im[15][12] ), .X(n9214) );
  inv_x2_sg U8980 ( .A(\i_im[12][13] ), .X(n9155) );
  inv_x2_sg U8981 ( .A(\i_im[6][13] ), .X(n9075) );
  inv_x1_sg U8982 ( .A(n1066), .X(n9015) );
  inv_x2_sg U8983 ( .A(\i_im[15][13] ), .X(n9215) );
  inv_x2_sg U8984 ( .A(\i_im[6][14] ), .X(n9076) );
  inv_x1_sg U8985 ( .A(n1098), .X(n9016) );
  nand_x1_sg U8986 ( .A(n6440), .B(n9036), .X(n1088) );
  inv_x2_sg U8987 ( .A(\i_im[4][14] ), .X(n9036) );
  inv_x2_sg U8988 ( .A(\i_im[15][14] ), .X(n9216) );
  inv_x2_sg U8989 ( .A(\i_im[12][15] ), .X(n9157) );
  inv_x2_sg U8990 ( .A(\i_im[6][15] ), .X(n9077) );
  inv_x1_sg U8991 ( .A(n807), .X(n9017) );
  inv_x2_sg U8992 ( .A(\i_im[15][15] ), .X(n9217) );
  inv_x2_sg U8993 ( .A(\i_im[6][16] ), .X(n9078) );
  inv_x1_sg U8994 ( .A(n839), .X(n9018) );
  inv_x2_sg U8995 ( .A(\i_im[15][16] ), .X(n9218) );
  inv_x2_sg U8996 ( .A(\i_im[6][17] ), .X(n9079) );
  inv_x1_sg U8997 ( .A(n871), .X(n9019) );
  inv_x2_sg U8998 ( .A(\i_im[15][17] ), .X(n9219) );
  inv_x2_sg U8999 ( .A(\i_im[6][18] ), .X(n9080) );
  inv_x1_sg U9000 ( .A(n903), .X(n9020) );
  inv_x2_sg U9001 ( .A(\i_im[15][18] ), .X(n9220) );
  inv_x2_sg U9002 ( .A(\i_im[15][19] ), .X(n9221) );
  inv_x2_sg U9003 ( .A(\i_im[13][19] ), .X(n9181) );
  inv_x1_sg U9004 ( .A(n941), .X(n9121) );
  inv_x2_sg U9005 ( .A(\i_im[6][19] ), .X(n9081) );
  inv_x1_sg U9006 ( .A(n935), .X(n9021) );
  nand_x1_sg U9007 ( .A(n6034), .B(n9061), .X(n934) );
  inv_x2_sg U9008 ( .A(\i_im[5][19] ), .X(n9061) );
  nand_x1_sg U9009 ( .A(n2247), .B(n2248), .X(n2246) );
  nor_x1_sg U9010 ( .A(n2240), .B(n2241), .X(n2239) );
  nor_x1_sg U9011 ( .A(n4843), .B(n4844), .X(n4842) );
  nand_x1_sg U9012 ( .A(n4845), .B(n4846), .X(n4844) );
  nor_x1_sg U9013 ( .A(n4851), .B(n4852), .X(n4841) );
  nand_x1_sg U9014 ( .A(n4853), .B(n4854), .X(n4852) );
  nor_x1_sg U9015 ( .A(n4828), .B(n4829), .X(n4827) );
  nand_x1_sg U9016 ( .A(n4830), .B(n4831), .X(n4829) );
  nand_x1_sg U9017 ( .A(n4832), .B(n4833), .X(n4828) );
  nor_x1_sg U9018 ( .A(n4836), .B(n4837), .X(n4826) );
  nand_x1_sg U9019 ( .A(n4839), .B(n4840), .X(n4836) );
  nor_x1_sg U9020 ( .A(n4805), .B(n4806), .X(n4804) );
  nand_x1_sg U9021 ( .A(n4807), .B(n4808), .X(n4806) );
  nor_x1_sg U9022 ( .A(n4812), .B(n4813), .X(n4803) );
  nand_x1_sg U9023 ( .A(n4814), .B(n4815), .X(n4813) );
  nor_x1_sg U9024 ( .A(n4790), .B(n4791), .X(n4789) );
  nand_x1_sg U9025 ( .A(n4792), .B(n4793), .X(n4791) );
  nand_x1_sg U9026 ( .A(n4794), .B(n4795), .X(n4790) );
  nor_x1_sg U9027 ( .A(n4798), .B(n4799), .X(n4788) );
  nand_x1_sg U9028 ( .A(n4801), .B(n4802), .X(n4798) );
  nor_x1_sg U9029 ( .A(n4754), .B(n4755), .X(n4753) );
  nand_x1_sg U9030 ( .A(n4756), .B(n4757), .X(n4755) );
  nand_x1_sg U9031 ( .A(n4758), .B(n4759), .X(n4754) );
  nor_x1_sg U9032 ( .A(n4762), .B(n4763), .X(n4752) );
  nand_x1_sg U9033 ( .A(n4765), .B(n4766), .X(n4762) );
  nor_x1_sg U9034 ( .A(n4769), .B(n4770), .X(n4768) );
  nand_x1_sg U9035 ( .A(n4771), .B(n4772), .X(n4770) );
  nor_x1_sg U9036 ( .A(n4776), .B(n4777), .X(n4767) );
  nand_x1_sg U9037 ( .A(n4778), .B(n4779), .X(n4777) );
  nor_x1_sg U9038 ( .A(n4733), .B(n4734), .X(n4732) );
  nand_x1_sg U9039 ( .A(n4735), .B(n4736), .X(n4734) );
  nor_x1_sg U9040 ( .A(n4740), .B(n4741), .X(n4731) );
  nand_x1_sg U9041 ( .A(n4742), .B(n4743), .X(n4741) );
  nor_x1_sg U9042 ( .A(n4718), .B(n4719), .X(n4717) );
  nand_x1_sg U9043 ( .A(n4720), .B(n4721), .X(n4719) );
  nand_x1_sg U9044 ( .A(n4722), .B(n4723), .X(n4718) );
  nor_x1_sg U9045 ( .A(n4726), .B(n4727), .X(n4716) );
  nand_x1_sg U9046 ( .A(n4729), .B(n4730), .X(n4726) );
  nor_x1_sg U9047 ( .A(n4682), .B(n4683), .X(n4681) );
  nand_x1_sg U9048 ( .A(n4684), .B(n4685), .X(n4683) );
  nand_x1_sg U9049 ( .A(n4686), .B(n4687), .X(n4682) );
  nor_x1_sg U9050 ( .A(n4690), .B(n4691), .X(n4680) );
  nand_x1_sg U9051 ( .A(n4693), .B(n4694), .X(n4690) );
  nor_x1_sg U9052 ( .A(n4697), .B(n4698), .X(n4696) );
  nand_x1_sg U9053 ( .A(n4699), .B(n4700), .X(n4698) );
  nor_x1_sg U9054 ( .A(n4704), .B(n4705), .X(n4695) );
  nand_x1_sg U9055 ( .A(n4706), .B(n4707), .X(n4705) );
  nor_x1_sg U9056 ( .A(n4661), .B(n4662), .X(n4660) );
  nand_x1_sg U9057 ( .A(n4663), .B(n4664), .X(n4662) );
  nor_x1_sg U9058 ( .A(n4668), .B(n4669), .X(n4659) );
  nand_x1_sg U9059 ( .A(n4670), .B(n4671), .X(n4669) );
  nor_x1_sg U9060 ( .A(n4646), .B(n4647), .X(n4645) );
  nand_x1_sg U9061 ( .A(n4650), .B(n4651), .X(n4646) );
  nand_x1_sg U9062 ( .A(n4648), .B(n4649), .X(n4647) );
  nor_x1_sg U9063 ( .A(n4654), .B(n4655), .X(n4644) );
  nand_x1_sg U9064 ( .A(n4657), .B(n4658), .X(n4654) );
  nor_x1_sg U9065 ( .A(n4610), .B(n4611), .X(n4609) );
  nand_x1_sg U9066 ( .A(n4612), .B(n4613), .X(n4611) );
  nand_x1_sg U9067 ( .A(n4614), .B(n4615), .X(n4610) );
  nor_x1_sg U9068 ( .A(n4618), .B(n4619), .X(n4608) );
  nand_x1_sg U9069 ( .A(n4621), .B(n4622), .X(n4618) );
  nor_x1_sg U9070 ( .A(n4625), .B(n4626), .X(n4624) );
  nand_x1_sg U9071 ( .A(n4627), .B(n4628), .X(n4626) );
  nor_x1_sg U9072 ( .A(n4632), .B(n4633), .X(n4623) );
  nand_x1_sg U9073 ( .A(n4634), .B(n4635), .X(n4633) );
  nor_x1_sg U9074 ( .A(n4574), .B(n4575), .X(n4573) );
  nand_x1_sg U9075 ( .A(n4578), .B(n4579), .X(n4574) );
  nand_x1_sg U9076 ( .A(n4576), .B(n4577), .X(n4575) );
  nor_x1_sg U9077 ( .A(n4582), .B(n4583), .X(n4572) );
  nand_x1_sg U9078 ( .A(n4585), .B(n4586), .X(n4582) );
  nor_x1_sg U9079 ( .A(n4589), .B(n4590), .X(n4588) );
  nand_x1_sg U9080 ( .A(n4591), .B(n4592), .X(n4590) );
  nor_x1_sg U9081 ( .A(n4596), .B(n4597), .X(n4587) );
  nand_x1_sg U9082 ( .A(n4598), .B(n4599), .X(n4597) );
  nor_x1_sg U9083 ( .A(n4538), .B(n4539), .X(n4537) );
  nand_x1_sg U9084 ( .A(n4540), .B(n4541), .X(n4539) );
  nand_x1_sg U9085 ( .A(n4542), .B(n4543), .X(n4538) );
  nor_x1_sg U9086 ( .A(n4546), .B(n4547), .X(n4536) );
  nand_x1_sg U9087 ( .A(n4549), .B(n4550), .X(n4546) );
  nor_x1_sg U9088 ( .A(n4553), .B(n4554), .X(n4552) );
  nand_x1_sg U9089 ( .A(n4555), .B(n4556), .X(n4554) );
  nor_x1_sg U9090 ( .A(n4560), .B(n4561), .X(n4551) );
  nand_x1_sg U9091 ( .A(n4562), .B(n4563), .X(n4561) );
  nor_x1_sg U9092 ( .A(n4517), .B(n4518), .X(n4516) );
  nand_x1_sg U9093 ( .A(n4519), .B(n4520), .X(n4518) );
  nor_x1_sg U9094 ( .A(n4524), .B(n4525), .X(n4515) );
  nand_x1_sg U9095 ( .A(n4526), .B(n4527), .X(n4525) );
  nor_x1_sg U9096 ( .A(n4502), .B(n4503), .X(n4501) );
  nand_x1_sg U9097 ( .A(n4506), .B(n4507), .X(n4502) );
  nand_x1_sg U9098 ( .A(n4504), .B(n4505), .X(n4503) );
  nor_x1_sg U9099 ( .A(n4510), .B(n4511), .X(n4500) );
  nand_x1_sg U9100 ( .A(n4513), .B(n4514), .X(n4510) );
  nor_x1_sg U9101 ( .A(n4466), .B(n4467), .X(n4465) );
  nand_x1_sg U9102 ( .A(n4468), .B(n4469), .X(n4467) );
  nand_x1_sg U9103 ( .A(n4470), .B(n4471), .X(n4466) );
  nor_x1_sg U9104 ( .A(n4474), .B(n4475), .X(n4464) );
  nand_x1_sg U9105 ( .A(n4477), .B(n4478), .X(n4474) );
  nor_x1_sg U9106 ( .A(n4481), .B(n4482), .X(n4480) );
  nand_x1_sg U9107 ( .A(n4483), .B(n4484), .X(n4482) );
  nor_x1_sg U9108 ( .A(n4488), .B(n4489), .X(n4479) );
  nand_x1_sg U9109 ( .A(n4490), .B(n4491), .X(n4489) );
  nor_x1_sg U9110 ( .A(n4430), .B(n4431), .X(n4429) );
  nand_x1_sg U9111 ( .A(n4434), .B(n4435), .X(n4430) );
  nand_x1_sg U9112 ( .A(n4432), .B(n4433), .X(n4431) );
  nor_x1_sg U9113 ( .A(n4438), .B(n4439), .X(n4428) );
  nand_x1_sg U9114 ( .A(n4441), .B(n4442), .X(n4438) );
  nor_x1_sg U9115 ( .A(n4445), .B(n4446), .X(n4444) );
  nand_x1_sg U9116 ( .A(n4447), .B(n4448), .X(n4446) );
  nor_x1_sg U9117 ( .A(n4452), .B(n4453), .X(n4443) );
  nand_x1_sg U9118 ( .A(n4454), .B(n4455), .X(n4453) );
  nor_x1_sg U9119 ( .A(n4409), .B(n4410), .X(n4408) );
  nand_x1_sg U9120 ( .A(n4411), .B(n4412), .X(n4410) );
  nand_x1_sg U9121 ( .A(n4413), .B(n4414), .X(n4409) );
  nand_x1_sg U9122 ( .A(n7129), .B(n5756), .X(n4412) );
  nor_x1_sg U9123 ( .A(n4416), .B(n4417), .X(n4407) );
  nand_x1_sg U9124 ( .A(n4420), .B(n4421), .X(n4416) );
  nand_x1_sg U9125 ( .A(n4418), .B(n4419), .X(n4417) );
  nor_x1_sg U9126 ( .A(n4394), .B(n4395), .X(n4393) );
  nand_x1_sg U9127 ( .A(n4396), .B(n4397), .X(n4395) );
  nor_x1_sg U9128 ( .A(n4402), .B(n4403), .X(n4392) );
  nand_x1_sg U9129 ( .A(n4405), .B(n4406), .X(n4402) );
  nor_x1_sg U9130 ( .A(n4373), .B(n4374), .X(n4372) );
  nand_x1_sg U9131 ( .A(n4375), .B(n4376), .X(n4374) );
  nand_x1_sg U9132 ( .A(n4377), .B(n4378), .X(n4373) );
  nand_x1_sg U9133 ( .A(n7258), .B(n5757), .X(n4375) );
  nor_x1_sg U9134 ( .A(n4380), .B(n4381), .X(n4371) );
  nand_x1_sg U9135 ( .A(n4384), .B(n4385), .X(n4380) );
  nand_x1_sg U9136 ( .A(n4382), .B(n4383), .X(n4381) );
  nor_x1_sg U9137 ( .A(n4358), .B(n4359), .X(n4357) );
  nand_x1_sg U9138 ( .A(n4360), .B(n4361), .X(n4359) );
  nor_x1_sg U9139 ( .A(n4366), .B(n4367), .X(n4356) );
  nand_x1_sg U9140 ( .A(n4369), .B(n4370), .X(n4366) );
  nor_x1_sg U9141 ( .A(n4337), .B(n4338), .X(n4336) );
  nand_x1_sg U9142 ( .A(n4339), .B(n4340), .X(n4338) );
  nand_x1_sg U9143 ( .A(n4341), .B(n4342), .X(n4337) );
  nand_x1_sg U9144 ( .A(n6394), .B(n5758), .X(n4339) );
  nor_x1_sg U9145 ( .A(n4344), .B(n4345), .X(n4335) );
  nand_x1_sg U9146 ( .A(n4346), .B(n4347), .X(n4345) );
  nand_x1_sg U9147 ( .A(n4348), .B(n4349), .X(n4344) );
  nor_x1_sg U9148 ( .A(n4322), .B(n4323), .X(n4321) );
  nand_x1_sg U9149 ( .A(n4324), .B(n4325), .X(n4323) );
  nor_x1_sg U9150 ( .A(n4330), .B(n4331), .X(n4320) );
  nand_x1_sg U9151 ( .A(n4333), .B(n4334), .X(n4330) );
  nor_x1_sg U9152 ( .A(n4301), .B(n4302), .X(n4300) );
  nand_x1_sg U9153 ( .A(n4303), .B(n4304), .X(n4302) );
  nand_x1_sg U9154 ( .A(n4305), .B(n4306), .X(n4301) );
  nand_x1_sg U9155 ( .A(n6076), .B(n5854), .X(n4303) );
  nor_x1_sg U9156 ( .A(n4308), .B(n4309), .X(n4299) );
  nand_x1_sg U9157 ( .A(n4312), .B(n4313), .X(n4308) );
  nor_x1_sg U9158 ( .A(n4286), .B(n4287), .X(n4285) );
  nand_x1_sg U9159 ( .A(n4288), .B(n4289), .X(n4287) );
  nand_x1_sg U9160 ( .A(n6393), .B(n5738), .X(n4289) );
  nor_x1_sg U9161 ( .A(n4294), .B(n4295), .X(n4284) );
  nand_x1_sg U9162 ( .A(n4297), .B(n4298), .X(n4294) );
  nor_x1_sg U9163 ( .A(n4250), .B(n4251), .X(n4249) );
  nand_x1_sg U9164 ( .A(n4252), .B(n4253), .X(n4251) );
  nand_x1_sg U9165 ( .A(n4254), .B(n4255), .X(n4250) );
  nor_x1_sg U9166 ( .A(n4258), .B(n4259), .X(n4248) );
  nand_x1_sg U9167 ( .A(n4261), .B(n4262), .X(n4258) );
  nor_x1_sg U9168 ( .A(n4265), .B(n4266), .X(n4264) );
  nand_x1_sg U9169 ( .A(n4267), .B(n4268), .X(n4266) );
  nor_x1_sg U9170 ( .A(n4272), .B(n4273), .X(n4263) );
  nand_x1_sg U9171 ( .A(n4274), .B(n4275), .X(n4273) );
  nor_x1_sg U9172 ( .A(n4229), .B(n4230), .X(n4228) );
  nand_x1_sg U9173 ( .A(n4231), .B(n4232), .X(n4230) );
  nor_x1_sg U9174 ( .A(n4236), .B(n4237), .X(n4227) );
  nand_x1_sg U9175 ( .A(n4238), .B(n4239), .X(n4237) );
  nor_x1_sg U9176 ( .A(n4214), .B(n4215), .X(n4213) );
  nand_x1_sg U9177 ( .A(n4216), .B(n4217), .X(n4215) );
  nand_x1_sg U9178 ( .A(n4218), .B(n4219), .X(n4214) );
  nor_x1_sg U9179 ( .A(n4222), .B(n4223), .X(n4212) );
  nand_x1_sg U9180 ( .A(n4225), .B(n4226), .X(n4222) );
  nor_x1_sg U9181 ( .A(n4178), .B(n4179), .X(n4177) );
  nand_x1_sg U9182 ( .A(n4180), .B(n4181), .X(n4179) );
  nand_x1_sg U9183 ( .A(n4182), .B(n4183), .X(n4178) );
  nor_x1_sg U9184 ( .A(n4186), .B(n4187), .X(n4176) );
  nand_x1_sg U9185 ( .A(n4189), .B(n4190), .X(n4186) );
  nor_x1_sg U9186 ( .A(n4193), .B(n4194), .X(n4192) );
  nand_x1_sg U9187 ( .A(n4195), .B(n4196), .X(n4194) );
  nor_x1_sg U9188 ( .A(n4200), .B(n4201), .X(n4191) );
  nand_x1_sg U9189 ( .A(n4202), .B(n4203), .X(n4201) );
  nor_x1_sg U9190 ( .A(n4157), .B(n4158), .X(n4156) );
  nand_x1_sg U9191 ( .A(n4159), .B(n4160), .X(n4158) );
  nor_x1_sg U9192 ( .A(n4164), .B(n4165), .X(n4155) );
  nand_x1_sg U9193 ( .A(n4166), .B(n4167), .X(n4165) );
  nor_x1_sg U9194 ( .A(n4136), .B(n4137), .X(n4135) );
  nand_x1_sg U9195 ( .A(n4138), .B(n4139), .X(n4137) );
  nand_x1_sg U9196 ( .A(n4141), .B(n4142), .X(n4136) );
  nor_x1_sg U9197 ( .A(n4148), .B(n4149), .X(n4134) );
  nand_x1_sg U9198 ( .A(n4152), .B(n4153), .X(n4148) );
  nand_x1_sg U9199 ( .A(n1431), .B(n9102), .X(n1430) );
  nand_x1_sg U9200 ( .A(n1434), .B(n1435), .X(n1429) );
  inv_x2_sg U9201 ( .A(\i_im[12][0] ), .X(n9142) );
  nor_x1_sg U9202 ( .A(n1421), .B(n1422), .X(n1412) );
  nand_x1_sg U9203 ( .A(n1423), .B(n1424), .X(n1422) );
  nor_x1_sg U9204 ( .A(n1414), .B(n1415), .X(n1413) );
  nor_x1_sg U9205 ( .A(n1439), .B(n1440), .X(n1427) );
  nand_x1_sg U9206 ( .A(n1140), .B(n9103), .X(n1139) );
  nand_x1_sg U9207 ( .A(n1142), .B(n1143), .X(n1138) );
  nor_x1_sg U9208 ( .A(n1130), .B(n1131), .X(n1121) );
  nand_x1_sg U9209 ( .A(n1132), .B(n1133), .X(n1131) );
  nor_x1_sg U9210 ( .A(n1123), .B(n1124), .X(n1122) );
  nor_x1_sg U9211 ( .A(n1146), .B(n1147), .X(n1136) );
  nand_x1_sg U9212 ( .A(n1172), .B(n9104), .X(n1171) );
  inv_x1_sg U9213 ( .A(n1173), .X(n9104) );
  inv_x2_sg U9214 ( .A(\i_im[13][2] ), .X(n9164) );
  nor_x1_sg U9215 ( .A(n1162), .B(n1163), .X(n1153) );
  nand_x1_sg U9216 ( .A(n1165), .B(n1164), .X(n1163) );
  nor_x1_sg U9217 ( .A(n1155), .B(n1156), .X(n1154) );
  nand_x1_sg U9218 ( .A(n1181), .B(n9124), .X(n1178) );
  inv_x1_sg U9219 ( .A(n1222), .X(n8965) );
  nand_x1_sg U9220 ( .A(n1223), .B(n8985), .X(n1219) );
  nor_x1_sg U9221 ( .A(n1242), .B(n1243), .X(n1232) );
  nor_x1_sg U9222 ( .A(n1234), .B(n1235), .X(n1233) );
  nand_x1_sg U9223 ( .A(n1236), .B(n9105), .X(n1235) );
  nand_x1_sg U9224 ( .A(n1228), .B(n1229), .X(n1227) );
  nand_x1_sg U9225 ( .A(n9005), .B(n1230), .X(n1226) );
  nand_x1_sg U9226 ( .A(n1204), .B(n9106), .X(n1203) );
  inv_x1_sg U9227 ( .A(n1205), .X(n9106) );
  inv_x2_sg U9228 ( .A(\i_im[13][4] ), .X(n9166) );
  nor_x1_sg U9229 ( .A(n1194), .B(n1195), .X(n1185) );
  nand_x1_sg U9230 ( .A(n1196), .B(n1197), .X(n1195) );
  nand_x1_sg U9231 ( .A(n1191), .B(n8986), .X(n1187) );
  nand_x1_sg U9232 ( .A(n8966), .B(n1189), .X(n1188) );
  nor_x1_sg U9233 ( .A(n1210), .B(n1211), .X(n1200) );
  nand_x1_sg U9234 ( .A(n1271), .B(n9107), .X(n1270) );
  inv_x1_sg U9235 ( .A(n1272), .X(n9107) );
  inv_x2_sg U9236 ( .A(\i_im[13][5] ), .X(n9167) );
  nor_x1_sg U9237 ( .A(n1261), .B(n1262), .X(n1252) );
  nand_x1_sg U9238 ( .A(n1263), .B(n1264), .X(n1262) );
  nor_x1_sg U9239 ( .A(n1254), .B(n1255), .X(n1253) );
  nand_x1_sg U9240 ( .A(n7320), .B(n1279), .X(n1278) );
  nand_x1_sg U9241 ( .A(n1280), .B(n9127), .X(n1277) );
  inv_x1_sg U9242 ( .A(n1289), .X(n8968) );
  nand_x1_sg U9243 ( .A(n1290), .B(n8988), .X(n1286) );
  nor_x1_sg U9244 ( .A(n1309), .B(n1310), .X(n1299) );
  nor_x1_sg U9245 ( .A(n1301), .B(n1302), .X(n1300) );
  nand_x1_sg U9246 ( .A(n1303), .B(n9108), .X(n1302) );
  nand_x1_sg U9247 ( .A(n1295), .B(n1296), .X(n1294) );
  nand_x1_sg U9248 ( .A(n9008), .B(n1297), .X(n1293) );
  inv_x1_sg U9249 ( .A(n1321), .X(n8969) );
  nand_x1_sg U9250 ( .A(n1322), .B(n8989), .X(n1318) );
  nor_x1_sg U9251 ( .A(n1341), .B(n1342), .X(n1331) );
  nor_x1_sg U9252 ( .A(n1333), .B(n1334), .X(n1332) );
  nand_x1_sg U9253 ( .A(n1335), .B(n9109), .X(n1334) );
  nand_x1_sg U9254 ( .A(n1327), .B(n1328), .X(n1326) );
  nand_x1_sg U9255 ( .A(n9009), .B(n1329), .X(n1325) );
  nand_x1_sg U9256 ( .A(n1367), .B(n9110), .X(n1366) );
  inv_x1_sg U9257 ( .A(n1368), .X(n9110) );
  inv_x2_sg U9258 ( .A(\i_im[13][8] ), .X(n9170) );
  nor_x1_sg U9259 ( .A(n1357), .B(n1358), .X(n1348) );
  nand_x1_sg U9260 ( .A(n1359), .B(n1360), .X(n1358) );
  nand_x1_sg U9261 ( .A(n1354), .B(n8990), .X(n1350) );
  nand_x1_sg U9262 ( .A(n8970), .B(n1352), .X(n1351) );
  nor_x1_sg U9263 ( .A(n1373), .B(n1374), .X(n1363) );
  inv_x1_sg U9264 ( .A(n1385), .X(n8971) );
  nand_x1_sg U9265 ( .A(n1386), .B(n8991), .X(n1382) );
  nor_x1_sg U9266 ( .A(n1405), .B(n1406), .X(n1395) );
  nor_x1_sg U9267 ( .A(n1397), .B(n1398), .X(n1396) );
  nand_x1_sg U9268 ( .A(n1391), .B(n1392), .X(n1390) );
  nand_x1_sg U9269 ( .A(n9011), .B(n1393), .X(n1389) );
  nand_x1_sg U9270 ( .A(n1007), .B(n9112), .X(n1006) );
  nand_x1_sg U9271 ( .A(n6421), .B(n9172), .X(n1007) );
  inv_x1_sg U9272 ( .A(n1008), .X(n9112) );
  inv_x2_sg U9273 ( .A(\i_im[13][10] ), .X(n9172) );
  nor_x1_sg U9274 ( .A(n997), .B(n998), .X(n988) );
  nand_x1_sg U9275 ( .A(n999), .B(n1000), .X(n998) );
  nand_x1_sg U9276 ( .A(n7263), .B(n9072), .X(n1000) );
  nand_x1_sg U9277 ( .A(n994), .B(n8992), .X(n990) );
  nand_x1_sg U9278 ( .A(n8972), .B(n992), .X(n991) );
  nor_x1_sg U9279 ( .A(n1013), .B(n1014), .X(n1003) );
  inv_x1_sg U9280 ( .A(n1025), .X(n8973) );
  nand_x1_sg U9281 ( .A(n1026), .B(n8993), .X(n1022) );
  nor_x1_sg U9282 ( .A(n1045), .B(n1046), .X(n1035) );
  nor_x1_sg U9283 ( .A(n1037), .B(n1038), .X(n1036) );
  nand_x1_sg U9284 ( .A(n1039), .B(n9113), .X(n1038) );
  nand_x1_sg U9285 ( .A(n9013), .B(n1033), .X(n1029) );
  nand_x1_sg U9286 ( .A(n1031), .B(n1032), .X(n1030) );
  nand_x1_sg U9287 ( .A(n6034), .B(n9053), .X(n1033) );
  nand_x1_sg U9288 ( .A(n975), .B(n9114), .X(n974) );
  nand_x1_sg U9289 ( .A(n7147), .B(n9174), .X(n975) );
  inv_x2_sg U9290 ( .A(\i_im[13][12] ), .X(n9174) );
  nand_x1_sg U9291 ( .A(n977), .B(n978), .X(n973) );
  inv_x2_sg U9292 ( .A(\i_im[12][12] ), .X(n9154) );
  nor_x1_sg U9293 ( .A(n965), .B(n966), .X(n956) );
  nand_x1_sg U9294 ( .A(n967), .B(n968), .X(n966) );
  nand_x1_sg U9295 ( .A(n7266), .B(n9074), .X(n968) );
  nor_x1_sg U9296 ( .A(n958), .B(n959), .X(n957) );
  nor_x1_sg U9297 ( .A(n981), .B(n982), .X(n971) );
  nand_x1_sg U9298 ( .A(n1071), .B(n9115), .X(n1070) );
  nand_x4_sg U9299 ( .A(n1073), .B(n1074), .X(n1069) );
  nand_x1_sg U9300 ( .A(n6171), .B(n9155), .X(n1074) );
  nor_x1_sg U9301 ( .A(n1061), .B(n1062), .X(n1052) );
  nand_x1_sg U9302 ( .A(n1063), .B(n1064), .X(n1062) );
  nor_x1_sg U9303 ( .A(n1054), .B(n1055), .X(n1053) );
  nor_x1_sg U9304 ( .A(n1077), .B(n1078), .X(n1067) );
  nand_x1_sg U9305 ( .A(n1103), .B(n9116), .X(n1102) );
  inv_x1_sg U9306 ( .A(n1104), .X(n9116) );
  inv_x2_sg U9307 ( .A(\i_im[13][14] ), .X(n9176) );
  nor_x1_sg U9308 ( .A(n1093), .B(n1094), .X(n1084) );
  nand_x1_sg U9309 ( .A(n1095), .B(n1096), .X(n1094) );
  nand_x1_sg U9310 ( .A(n1090), .B(n8996), .X(n1086) );
  nand_x1_sg U9311 ( .A(n8976), .B(n1088), .X(n1087) );
  nor_x1_sg U9312 ( .A(n1109), .B(n1110), .X(n1099) );
  nand_x1_sg U9313 ( .A(n814), .B(n815), .X(n810) );
  nand_x1_sg U9314 ( .A(n812), .B(n9117), .X(n811) );
  nor_x1_sg U9315 ( .A(n800), .B(n801), .X(n787) );
  nand_x1_sg U9316 ( .A(n802), .B(n803), .X(n801) );
  nor_x1_sg U9317 ( .A(n789), .B(n790), .X(n788) );
  nor_x1_sg U9318 ( .A(n818), .B(n819), .X(n808) );
  nand_x1_sg U9319 ( .A(n844), .B(n9118), .X(n843) );
  nand_x1_sg U9320 ( .A(n846), .B(n847), .X(n842) );
  inv_x2_sg U9321 ( .A(\i_im[12][16] ), .X(n9158) );
  nor_x1_sg U9322 ( .A(n834), .B(n835), .X(n825) );
  nand_x1_sg U9323 ( .A(n836), .B(n837), .X(n835) );
  nor_x1_sg U9324 ( .A(n827), .B(n828), .X(n826) );
  nor_x1_sg U9325 ( .A(n850), .B(n851), .X(n840) );
  nand_x1_sg U9326 ( .A(n876), .B(n9119), .X(n875) );
  nand_x1_sg U9327 ( .A(n878), .B(n879), .X(n874) );
  inv_x2_sg U9328 ( .A(\i_im[12][17] ), .X(n9159) );
  nor_x1_sg U9329 ( .A(n866), .B(n867), .X(n857) );
  nand_x1_sg U9330 ( .A(n868), .B(n869), .X(n867) );
  nor_x1_sg U9331 ( .A(n859), .B(n860), .X(n858) );
  nor_x1_sg U9332 ( .A(n882), .B(n883), .X(n872) );
  nand_x1_sg U9333 ( .A(n908), .B(n9120), .X(n907) );
  nand_x1_sg U9334 ( .A(n910), .B(n911), .X(n906) );
  inv_x2_sg U9335 ( .A(\i_im[12][18] ), .X(n9160) );
  nor_x1_sg U9336 ( .A(n898), .B(n899), .X(n889) );
  nand_x1_sg U9337 ( .A(n900), .B(n901), .X(n899) );
  nor_x1_sg U9338 ( .A(n891), .B(n892), .X(n890) );
  nor_x1_sg U9339 ( .A(n914), .B(n915), .X(n904) );
  nand_x1_sg U9340 ( .A(n8981), .B(n925), .X(n924) );
  inv_x2_sg U9341 ( .A(\i_im[4][19] ), .X(n9041) );
  nand_x1_sg U9342 ( .A(n927), .B(n9001), .X(n923) );
  nor_x1_sg U9343 ( .A(n946), .B(n947), .X(n936) );
  nor_x1_sg U9344 ( .A(n938), .B(n939), .X(n937) );
  nand_x1_sg U9345 ( .A(n940), .B(n9121), .X(n939) );
  nand_x1_sg U9346 ( .A(n7147), .B(n9181), .X(n940) );
  nor_x1_sg U9347 ( .A(n930), .B(n931), .X(n921) );
  nand_x1_sg U9348 ( .A(n932), .B(n933), .X(n931) );
  nand_x1_sg U9349 ( .A(n7262), .B(n9081), .X(n933) );
  nand_x2_sg U9350 ( .A(n1247), .B(n1248), .X(n1114) );
  nand_x2_sg U9351 ( .A(n1116), .B(n1117), .X(n1115) );
  inv_x1_sg U9352 ( .A(n2204), .X(n8898) );
  nor_x1_sg U9353 ( .A(n2245), .B(n2246), .X(n2228) );
  nand_x2_sg U9354 ( .A(n2232), .B(n2233), .X(n2231) );
  nor_x1_sg U9355 ( .A(n2212), .B(n2213), .X(n2211) );
  nand_x1_sg U9356 ( .A(n3782), .B(n9226), .X(n3781) );
  nand_x2_sg U9357 ( .A(n4824), .B(n4825), .X(n4823) );
  nand_x2_sg U9358 ( .A(n4826), .B(n4827), .X(n4825) );
  nand_x2_sg U9359 ( .A(n4841), .B(n4842), .X(n4824) );
  nand_x2_sg U9360 ( .A(n4786), .B(n4787), .X(n4785) );
  nand_x2_sg U9361 ( .A(n4788), .B(n4789), .X(n4787) );
  nand_x2_sg U9362 ( .A(n4803), .B(n4804), .X(n4786) );
  nand_x2_sg U9363 ( .A(n4750), .B(n4751), .X(n4749) );
  nand_x2_sg U9364 ( .A(n4767), .B(n4768), .X(n4750) );
  nand_x2_sg U9365 ( .A(n4752), .B(n4753), .X(n4751) );
  nand_x2_sg U9366 ( .A(n4714), .B(n4715), .X(n4713) );
  nand_x2_sg U9367 ( .A(n4716), .B(n4717), .X(n4715) );
  nand_x2_sg U9368 ( .A(n4731), .B(n4732), .X(n4714) );
  nand_x2_sg U9369 ( .A(n4678), .B(n4679), .X(n4677) );
  nand_x2_sg U9370 ( .A(n4695), .B(n4696), .X(n4678) );
  nand_x2_sg U9371 ( .A(n4680), .B(n4681), .X(n4679) );
  nand_x2_sg U9372 ( .A(n4642), .B(n4643), .X(n4641) );
  nand_x2_sg U9373 ( .A(n4644), .B(n4645), .X(n4643) );
  nand_x2_sg U9374 ( .A(n4659), .B(n4660), .X(n4642) );
  nand_x2_sg U9375 ( .A(n4606), .B(n4607), .X(n4605) );
  nand_x2_sg U9376 ( .A(n4623), .B(n4624), .X(n4606) );
  nand_x2_sg U9377 ( .A(n4608), .B(n4609), .X(n4607) );
  nand_x2_sg U9378 ( .A(n4570), .B(n4571), .X(n4569) );
  nand_x2_sg U9379 ( .A(n4587), .B(n4588), .X(n4570) );
  nand_x2_sg U9380 ( .A(n4572), .B(n4573), .X(n4571) );
  nand_x2_sg U9381 ( .A(n4534), .B(n4535), .X(n4533) );
  nand_x2_sg U9382 ( .A(n4551), .B(n4552), .X(n4534) );
  nand_x2_sg U9383 ( .A(n4536), .B(n4537), .X(n4535) );
  nand_x2_sg U9384 ( .A(n4498), .B(n4499), .X(n4497) );
  nand_x2_sg U9385 ( .A(n4500), .B(n4501), .X(n4499) );
  nand_x2_sg U9386 ( .A(n4515), .B(n4516), .X(n4498) );
  nand_x2_sg U9387 ( .A(n4462), .B(n4463), .X(n4461) );
  nand_x2_sg U9388 ( .A(n4479), .B(n4480), .X(n4462) );
  nand_x2_sg U9389 ( .A(n4464), .B(n4465), .X(n4463) );
  nand_x2_sg U9390 ( .A(n4426), .B(n4427), .X(n4425) );
  nand_x2_sg U9391 ( .A(n4443), .B(n4444), .X(n4426) );
  nand_x2_sg U9392 ( .A(n4428), .B(n4429), .X(n4427) );
  nand_x2_sg U9393 ( .A(n4390), .B(n4391), .X(n4389) );
  nand_x2_sg U9394 ( .A(n4392), .B(n4393), .X(n4391) );
  nand_x2_sg U9395 ( .A(n4407), .B(n4408), .X(n4390) );
  nand_x2_sg U9396 ( .A(n4354), .B(n4355), .X(n4353) );
  nand_x2_sg U9397 ( .A(n4356), .B(n4357), .X(n4355) );
  nand_x2_sg U9398 ( .A(n4371), .B(n4372), .X(n4354) );
  nand_x2_sg U9399 ( .A(n4318), .B(n4319), .X(n4317) );
  nand_x2_sg U9400 ( .A(n4320), .B(n4321), .X(n4319) );
  nand_x2_sg U9401 ( .A(n4335), .B(n4336), .X(n4318) );
  nand_x2_sg U9402 ( .A(n4282), .B(n4283), .X(n4281) );
  nand_x2_sg U9403 ( .A(n4284), .B(n4285), .X(n4283) );
  nand_x2_sg U9404 ( .A(n4299), .B(n4300), .X(n4282) );
  nand_x2_sg U9405 ( .A(n4246), .B(n4247), .X(n4245) );
  nand_x2_sg U9406 ( .A(n4263), .B(n4264), .X(n4246) );
  nand_x2_sg U9407 ( .A(n4248), .B(n4249), .X(n4247) );
  nand_x2_sg U9408 ( .A(n4210), .B(n4211), .X(n4209) );
  nand_x2_sg U9409 ( .A(n4212), .B(n4213), .X(n4211) );
  nand_x2_sg U9410 ( .A(n4227), .B(n4228), .X(n4210) );
  nand_x2_sg U9411 ( .A(n4174), .B(n4175), .X(n4173) );
  nand_x2_sg U9412 ( .A(n4191), .B(n4192), .X(n4174) );
  nand_x2_sg U9413 ( .A(n4176), .B(n4177), .X(n4175) );
  nand_x2_sg U9414 ( .A(n4132), .B(n4133), .X(n4131) );
  nand_x2_sg U9415 ( .A(n4134), .B(n4135), .X(n4133) );
  nand_x2_sg U9416 ( .A(n4155), .B(n4156), .X(n4132) );
  nor_x1_sg U9417 ( .A(n1170), .B(n1171), .X(n1169) );
  nor_x1_sg U9418 ( .A(n1219), .B(n1220), .X(n1218) );
  nor_x1_sg U9419 ( .A(n1202), .B(n1203), .X(n1201) );
  nor_x1_sg U9420 ( .A(n1269), .B(n1270), .X(n1268) );
  nor_x1_sg U9421 ( .A(n1286), .B(n1287), .X(n1285) );
  nor_x1_sg U9422 ( .A(n1318), .B(n1319), .X(n1317) );
  nor_x1_sg U9423 ( .A(n1365), .B(n1366), .X(n1364) );
  nor_x1_sg U9424 ( .A(n1382), .B(n1383), .X(n1381) );
  nor_x1_sg U9425 ( .A(n1005), .B(n1006), .X(n1004) );
  nor_x1_sg U9426 ( .A(n1022), .B(n1023), .X(n1021) );
  nor_x1_sg U9427 ( .A(n1101), .B(n1102), .X(n1100) );
  nor_x1_sg U9428 ( .A(n780), .B(n781), .X(n779) );
  nand_x1_sg U9429 ( .A(n951), .B(n952), .X(n780) );
  nand_x1_sg U9430 ( .A(n2194), .B(n2195), .X(n2193) );
  nand_x1_sg U9431 ( .A(n8898), .B(n2196), .X(n2195) );
  inv_x1_sg U9432 ( .A(n3443), .X(n9223) );
  inv_x1_sg U9433 ( .A(n7423), .X(n9239) );
  nand_x1_sg U9434 ( .A(n3451), .B(n6240), .X(n3448) );
  nand_x1_sg U9435 ( .A(n3432), .B(n4861), .X(n3443) );
  nor_x1_sg U9436 ( .A(n4886), .B(n4887), .X(n4879) );
  nor_x1_sg U9437 ( .A(n5640), .B(n5641), .X(n5639) );
  inv_x1_sg U9438 ( .A(n5630), .X(n9230) );
  nand_x2_sg U9439 ( .A(n5607), .B(n6160), .X(n4867) );
  nand_x1_sg U9440 ( .A(\update_output_0/N29 ), .B(n7395), .X(n7459) );
  nand_x1_sg U9441 ( .A(\output_state[0] ), .B(n7374), .X(n3452) );
  nor_x1_sg U9442 ( .A(n9222), .B(n6081), .X(n3524) );
  nand_x1_sg U9443 ( .A(n3469), .B(n9224), .X(\update_output_0/n3144 ) );
  inv_x1_sg U9444 ( .A(n3470), .X(n9224) );
  nand_x1_sg U9445 ( .A(n1399), .B(n9111), .X(n1398) );
  nand_x2_sg U9446 ( .A(n4310), .B(n4311), .X(n4309) );
  nand_x1_sg U9447 ( .A(n3459), .B(n3460), .X(\update_output_0/n3146 ) );
  nand_x1_sg U9448 ( .A(n3437), .B(n3438), .X(\update_output_0/n3150 ) );
  nand_x1_sg U9449 ( .A(n9231), .B(n4874), .X(n4873) );
  inv_x1_sg U9450 ( .A(n4875), .X(n9231) );
  nand_x1_sg U9451 ( .A(n5595), .B(n5596), .X(\update_mask_0/n1086 ) );
  nand_x1_sg U9452 ( .A(n5608), .B(n5609), .X(\update_mask_0/n1083 ) );
  nand_x1_sg U9453 ( .A(n5610), .B(n9228), .X(n5609) );
  inv_x1_sg U9454 ( .A(n2198), .X(n8901) );
  inv_x1_sg U9455 ( .A(n1789), .X(n8930) );
  inv_x1_sg U9456 ( .A(n2127), .X(n8938) );
  inv_x1_sg U9457 ( .A(n1517), .X(n8923) );
  inv_x1_sg U9458 ( .A(n1621), .X(n8926) );
  inv_x1_sg U9459 ( .A(n1691), .X(n8927) );
  inv_x1_sg U9460 ( .A(n1861), .X(n8931) );
  inv_x1_sg U9461 ( .A(n1959), .X(n8934) );
  inv_x1_sg U9462 ( .A(n2029), .X(n8935) );
  inv_x1_sg U9463 ( .A(n1538), .X(n8924) );
  inv_x1_sg U9464 ( .A(n1606), .X(n8925) );
  inv_x1_sg U9465 ( .A(n1706), .X(n8928) );
  inv_x1_sg U9466 ( .A(n1876), .X(n8932) );
  inv_x1_sg U9467 ( .A(n1944), .X(n8933) );
  inv_x1_sg U9468 ( .A(n2044), .X(n8936) );
  inv_x1_sg U9469 ( .A(n1501), .X(n8961) );
  nand_x1_sg U9470 ( .A(n4080), .B(n4081), .X(\update_output_0/n2863 ) );
  nand_x1_sg U9471 ( .A(n4078), .B(n4079), .X(\update_output_0/n2864 ) );
  nand_x1_sg U9472 ( .A(n4074), .B(n4075), .X(\update_output_0/n2866 ) );
  nand_x1_sg U9473 ( .A(n4070), .B(n4071), .X(\update_output_0/n2868 ) );
  nand_x1_sg U9474 ( .A(n4066), .B(n4067), .X(\update_output_0/n2870 ) );
  nand_x1_sg U9475 ( .A(n4062), .B(n4063), .X(\update_output_0/n2872 ) );
  nand_x1_sg U9476 ( .A(n4058), .B(n4059), .X(\update_output_0/n2874 ) );
  nand_x1_sg U9477 ( .A(n4054), .B(n4055), .X(\update_output_0/n2876 ) );
  nand_x1_sg U9478 ( .A(n4050), .B(n4051), .X(\update_output_0/n2878 ) );
  nand_x1_sg U9479 ( .A(n4046), .B(n4047), .X(\update_output_0/n2880 ) );
  nand_x1_sg U9480 ( .A(n4041), .B(n4042), .X(\update_output_0/n2882 ) );
  nand_x1_sg U9481 ( .A(n3951), .B(n3952), .X(\update_output_0/n2923 ) );
  nand_x1_sg U9482 ( .A(n3949), .B(n3950), .X(\update_output_0/n2924 ) );
  nand_x1_sg U9483 ( .A(n3945), .B(n3946), .X(\update_output_0/n2926 ) );
  nand_x1_sg U9484 ( .A(n3941), .B(n3942), .X(\update_output_0/n2928 ) );
  nand_x1_sg U9485 ( .A(n3937), .B(n3938), .X(\update_output_0/n2930 ) );
  nand_x1_sg U9486 ( .A(n3933), .B(n3934), .X(\update_output_0/n2932 ) );
  nand_x1_sg U9487 ( .A(n3929), .B(n3930), .X(\update_output_0/n2934 ) );
  nand_x1_sg U9488 ( .A(n3925), .B(n3926), .X(\update_output_0/n2936 ) );
  nand_x1_sg U9489 ( .A(n3921), .B(n3922), .X(\update_output_0/n2938 ) );
  nand_x1_sg U9490 ( .A(n3917), .B(n3918), .X(\update_output_0/n2940 ) );
  nand_x1_sg U9491 ( .A(n3912), .B(n3913), .X(\update_output_0/n2942 ) );
  nand_x1_sg U9492 ( .A(n3984), .B(n3985), .X(\update_output_0/n2908 ) );
  nand_x1_sg U9493 ( .A(n3982), .B(n3983), .X(\update_output_0/n2909 ) );
  nand_x1_sg U9494 ( .A(n3980), .B(n3981), .X(\update_output_0/n2910 ) );
  nand_x1_sg U9495 ( .A(n3978), .B(n3979), .X(\update_output_0/n2911 ) );
  nand_x1_sg U9496 ( .A(n3976), .B(n3977), .X(\update_output_0/n2912 ) );
  nand_x1_sg U9497 ( .A(n3974), .B(n3975), .X(\update_output_0/n2913 ) );
  nand_x1_sg U9498 ( .A(n3972), .B(n3973), .X(\update_output_0/n2914 ) );
  nand_x1_sg U9499 ( .A(n3970), .B(n3971), .X(\update_output_0/n2915 ) );
  nand_x1_sg U9500 ( .A(n3968), .B(n3969), .X(\update_output_0/n2916 ) );
  nand_x1_sg U9501 ( .A(n3966), .B(n3967), .X(\update_output_0/n2917 ) );
  nand_x1_sg U9502 ( .A(n3964), .B(n3965), .X(\update_output_0/n2918 ) );
  nand_x1_sg U9503 ( .A(n3962), .B(n3963), .X(\update_output_0/n2919 ) );
  nand_x1_sg U9504 ( .A(n3960), .B(n3961), .X(\update_output_0/n2920 ) );
  nand_x1_sg U9505 ( .A(n3958), .B(n3959), .X(\update_output_0/n2921 ) );
  nand_x1_sg U9506 ( .A(n3955), .B(n3956), .X(\update_output_0/n2922 ) );
  nand_x1_sg U9507 ( .A(n3866), .B(n3867), .X(\update_output_0/n2963 ) );
  nand_x1_sg U9508 ( .A(n3864), .B(n3865), .X(\update_output_0/n2964 ) );
  nand_x1_sg U9509 ( .A(n3862), .B(n3863), .X(\update_output_0/n2965 ) );
  nand_x1_sg U9510 ( .A(n3860), .B(n3861), .X(\update_output_0/n2966 ) );
  nand_x1_sg U9511 ( .A(n3858), .B(n3859), .X(\update_output_0/n2967 ) );
  nand_x1_sg U9512 ( .A(n3856), .B(n3857), .X(\update_output_0/n2968 ) );
  nand_x1_sg U9513 ( .A(n3854), .B(n3855), .X(\update_output_0/n2969 ) );
  nand_x1_sg U9514 ( .A(n3852), .B(n3853), .X(\update_output_0/n2970 ) );
  nand_x1_sg U9515 ( .A(n3850), .B(n3851), .X(\update_output_0/n2971 ) );
  nand_x1_sg U9516 ( .A(n3848), .B(n3849), .X(\update_output_0/n2972 ) );
  nand_x1_sg U9517 ( .A(n3846), .B(n3847), .X(\update_output_0/n2973 ) );
  nand_x1_sg U9518 ( .A(n3844), .B(n3845), .X(\update_output_0/n2974 ) );
  nand_x1_sg U9519 ( .A(n3842), .B(n3843), .X(\update_output_0/n2975 ) );
  nand_x1_sg U9520 ( .A(n3840), .B(n3841), .X(\update_output_0/n2976 ) );
  nand_x1_sg U9521 ( .A(n3838), .B(n3839), .X(\update_output_0/n2977 ) );
  nand_x1_sg U9522 ( .A(n3836), .B(n3837), .X(\update_output_0/n2978 ) );
  nand_x1_sg U9523 ( .A(n3834), .B(n3835), .X(\update_output_0/n2979 ) );
  nand_x1_sg U9524 ( .A(n3832), .B(n3833), .X(\update_output_0/n2980 ) );
  nand_x1_sg U9525 ( .A(n3830), .B(n3831), .X(\update_output_0/n2981 ) );
  nand_x1_sg U9526 ( .A(n3827), .B(n3828), .X(\update_output_0/n2982 ) );
  nand_x1_sg U9527 ( .A(n4122), .B(n4123), .X(\update_output_0/n2843 ) );
  nand_x1_sg U9528 ( .A(n4120), .B(n4121), .X(\update_output_0/n2844 ) );
  nand_x1_sg U9529 ( .A(n4118), .B(n4119), .X(\update_output_0/n2845 ) );
  nand_x1_sg U9530 ( .A(n4116), .B(n4117), .X(\update_output_0/n2846 ) );
  nand_x1_sg U9531 ( .A(n4114), .B(n4115), .X(\update_output_0/n2847 ) );
  nand_x1_sg U9532 ( .A(n4112), .B(n4113), .X(\update_output_0/n2848 ) );
  nand_x1_sg U9533 ( .A(n4110), .B(n4111), .X(\update_output_0/n2849 ) );
  nand_x1_sg U9534 ( .A(n4108), .B(n4109), .X(\update_output_0/n2850 ) );
  nand_x1_sg U9535 ( .A(n4106), .B(n4107), .X(\update_output_0/n2851 ) );
  nand_x1_sg U9536 ( .A(n4104), .B(n4105), .X(\update_output_0/n2852 ) );
  nand_x1_sg U9537 ( .A(n4102), .B(n4103), .X(\update_output_0/n2853 ) );
  nand_x1_sg U9538 ( .A(n4100), .B(n4101), .X(\update_output_0/n2854 ) );
  nand_x1_sg U9539 ( .A(n4098), .B(n4099), .X(\update_output_0/n2855 ) );
  nand_x1_sg U9540 ( .A(n4096), .B(n4097), .X(\update_output_0/n2856 ) );
  nand_x1_sg U9541 ( .A(n4094), .B(n4095), .X(\update_output_0/n2857 ) );
  nand_x1_sg U9542 ( .A(n4092), .B(n4093), .X(\update_output_0/n2858 ) );
  nand_x1_sg U9543 ( .A(n4090), .B(n4091), .X(\update_output_0/n2859 ) );
  nand_x1_sg U9544 ( .A(n4088), .B(n4089), .X(\update_output_0/n2860 ) );
  nand_x1_sg U9545 ( .A(n4086), .B(n4087), .X(\update_output_0/n2861 ) );
  nand_x1_sg U9546 ( .A(n4083), .B(n4084), .X(\update_output_0/n2862 ) );
  nand_x1_sg U9547 ( .A(n3994), .B(n3995), .X(\update_output_0/n2903 ) );
  nand_x1_sg U9548 ( .A(n3992), .B(n3993), .X(\update_output_0/n2904 ) );
  nand_x1_sg U9549 ( .A(n3990), .B(n3991), .X(\update_output_0/n2905 ) );
  nand_x1_sg U9550 ( .A(n3988), .B(n3989), .X(\update_output_0/n2906 ) );
  nand_x1_sg U9551 ( .A(n3986), .B(n3987), .X(\update_output_0/n2907 ) );
  nand_x1_sg U9552 ( .A(n4076), .B(n4077), .X(\update_output_0/n2865 ) );
  nand_x1_sg U9553 ( .A(n4072), .B(n4073), .X(\update_output_0/n2867 ) );
  nand_x1_sg U9554 ( .A(n4068), .B(n4069), .X(\update_output_0/n2869 ) );
  nand_x1_sg U9555 ( .A(n4064), .B(n4065), .X(\update_output_0/n2871 ) );
  nand_x1_sg U9556 ( .A(n4060), .B(n4061), .X(\update_output_0/n2873 ) );
  nand_x1_sg U9557 ( .A(n4056), .B(n4057), .X(\update_output_0/n2875 ) );
  nand_x1_sg U9558 ( .A(n4052), .B(n4053), .X(\update_output_0/n2877 ) );
  nand_x1_sg U9559 ( .A(n4048), .B(n4049), .X(\update_output_0/n2879 ) );
  nand_x1_sg U9560 ( .A(n4044), .B(n4045), .X(\update_output_0/n2881 ) );
  nand_x1_sg U9561 ( .A(n3947), .B(n3948), .X(\update_output_0/n2925 ) );
  nand_x1_sg U9562 ( .A(n3943), .B(n3944), .X(\update_output_0/n2927 ) );
  nand_x1_sg U9563 ( .A(n3939), .B(n3940), .X(\update_output_0/n2929 ) );
  nand_x1_sg U9564 ( .A(n3935), .B(n3936), .X(\update_output_0/n2931 ) );
  nand_x1_sg U9565 ( .A(n3931), .B(n3932), .X(\update_output_0/n2933 ) );
  nand_x1_sg U9566 ( .A(n3927), .B(n3928), .X(\update_output_0/n2935 ) );
  nand_x1_sg U9567 ( .A(n3923), .B(n3924), .X(\update_output_0/n2937 ) );
  nand_x1_sg U9568 ( .A(n3919), .B(n3920), .X(\update_output_0/n2939 ) );
  nand_x1_sg U9569 ( .A(n3915), .B(n3916), .X(\update_output_0/n2941 ) );
  nand_x1_sg U9570 ( .A(n3905), .B(n3906), .X(\update_output_0/n2945 ) );
  nand_x1_sg U9571 ( .A(n3901), .B(n3902), .X(\update_output_0/n2947 ) );
  nand_x1_sg U9572 ( .A(n3897), .B(n3898), .X(\update_output_0/n2949 ) );
  nand_x1_sg U9573 ( .A(n3893), .B(n3894), .X(\update_output_0/n2951 ) );
  nand_x1_sg U9574 ( .A(n3889), .B(n3890), .X(\update_output_0/n2953 ) );
  nand_x1_sg U9575 ( .A(n3885), .B(n3886), .X(\update_output_0/n2955 ) );
  nand_x1_sg U9576 ( .A(n3881), .B(n3882), .X(\update_output_0/n2957 ) );
  nand_x1_sg U9577 ( .A(n3877), .B(n3878), .X(\update_output_0/n2959 ) );
  nand_x1_sg U9578 ( .A(n3873), .B(n3874), .X(\update_output_0/n2961 ) );
  nand_x1_sg U9579 ( .A(n4033), .B(n4034), .X(\update_output_0/n2885 ) );
  nand_x1_sg U9580 ( .A(n4029), .B(n4030), .X(\update_output_0/n2887 ) );
  nand_x1_sg U9581 ( .A(n4025), .B(n4026), .X(\update_output_0/n2889 ) );
  nand_x1_sg U9582 ( .A(n4021), .B(n4022), .X(\update_output_0/n2891 ) );
  nand_x1_sg U9583 ( .A(n4017), .B(n4018), .X(\update_output_0/n2893 ) );
  nand_x1_sg U9584 ( .A(n4013), .B(n4014), .X(\update_output_0/n2895 ) );
  nand_x1_sg U9585 ( .A(n4009), .B(n4010), .X(\update_output_0/n2897 ) );
  nand_x1_sg U9586 ( .A(n4005), .B(n4006), .X(\update_output_0/n2899 ) );
  nand_x1_sg U9587 ( .A(n4001), .B(n4002), .X(\update_output_0/n2901 ) );
  nand_x1_sg U9588 ( .A(n3909), .B(n3910), .X(\update_output_0/n2943 ) );
  nand_x1_sg U9589 ( .A(n3907), .B(n3908), .X(\update_output_0/n2944 ) );
  nand_x1_sg U9590 ( .A(n3903), .B(n3904), .X(\update_output_0/n2946 ) );
  nand_x1_sg U9591 ( .A(n3899), .B(n3900), .X(\update_output_0/n2948 ) );
  nand_x1_sg U9592 ( .A(n3895), .B(n3896), .X(\update_output_0/n2950 ) );
  nand_x1_sg U9593 ( .A(n3891), .B(n3892), .X(\update_output_0/n2952 ) );
  nand_x1_sg U9594 ( .A(n3887), .B(n3888), .X(\update_output_0/n2954 ) );
  nand_x1_sg U9595 ( .A(n3883), .B(n3884), .X(\update_output_0/n2956 ) );
  nand_x1_sg U9596 ( .A(n3879), .B(n3880), .X(\update_output_0/n2958 ) );
  nand_x1_sg U9597 ( .A(n3875), .B(n3876), .X(\update_output_0/n2960 ) );
  nand_x1_sg U9598 ( .A(n3870), .B(n3871), .X(\update_output_0/n2962 ) );
  nand_x1_sg U9599 ( .A(n4037), .B(n4038), .X(\update_output_0/n2883 ) );
  nand_x1_sg U9600 ( .A(n4035), .B(n4036), .X(\update_output_0/n2884 ) );
  nand_x1_sg U9601 ( .A(n4031), .B(n4032), .X(\update_output_0/n2886 ) );
  nand_x1_sg U9602 ( .A(n4027), .B(n4028), .X(\update_output_0/n2888 ) );
  nand_x1_sg U9603 ( .A(n4023), .B(n4024), .X(\update_output_0/n2890 ) );
  nand_x1_sg U9604 ( .A(n4019), .B(n4020), .X(\update_output_0/n2892 ) );
  nand_x1_sg U9605 ( .A(n4015), .B(n4016), .X(\update_output_0/n2894 ) );
  nand_x1_sg U9606 ( .A(n4011), .B(n4012), .X(\update_output_0/n2896 ) );
  nand_x1_sg U9607 ( .A(n4007), .B(n4008), .X(\update_output_0/n2898 ) );
  nand_x1_sg U9608 ( .A(n4003), .B(n4004), .X(\update_output_0/n2900 ) );
  nand_x1_sg U9609 ( .A(n3998), .B(n3999), .X(\update_output_0/n2902 ) );
  nand_x1_sg U9610 ( .A(n4818), .B(n4819), .X(\update_output_0/n2823 ) );
  nand_x1_sg U9611 ( .A(n4782), .B(n4783), .X(\update_output_0/n2824 ) );
  nand_x1_sg U9612 ( .A(n4746), .B(n4747), .X(\update_output_0/n2825 ) );
  nand_x1_sg U9613 ( .A(n4710), .B(n4711), .X(\update_output_0/n2826 ) );
  nand_x1_sg U9614 ( .A(n4674), .B(n4675), .X(\update_output_0/n2827 ) );
  nand_x1_sg U9615 ( .A(n4638), .B(n4639), .X(\update_output_0/n2828 ) );
  nand_x1_sg U9616 ( .A(n4603), .B(n4602), .X(\update_output_0/n2829 ) );
  nand_x1_sg U9617 ( .A(n4566), .B(n4567), .X(\update_output_0/n2830 ) );
  nand_x1_sg U9618 ( .A(n4531), .B(n4530), .X(\update_output_0/n2831 ) );
  nand_x1_sg U9619 ( .A(n4494), .B(n4495), .X(\update_output_0/n2832 ) );
  nand_x1_sg U9620 ( .A(n4458), .B(n4459), .X(\update_output_0/n2833 ) );
  nand_x1_sg U9621 ( .A(n4422), .B(n4423), .X(\update_output_0/n2834 ) );
  nand_x1_sg U9622 ( .A(n4386), .B(n4387), .X(\update_output_0/n2835 ) );
  nand_x1_sg U9623 ( .A(n4350), .B(n4351), .X(\update_output_0/n2836 ) );
  nand_x1_sg U9624 ( .A(n4314), .B(n4315), .X(\update_output_0/n2837 ) );
  nand_x1_sg U9625 ( .A(n4278), .B(n4279), .X(\update_output_0/n2838 ) );
  nand_x1_sg U9626 ( .A(n4242), .B(n4243), .X(\update_output_0/n2839 ) );
  nand_x1_sg U9627 ( .A(n4206), .B(n4207), .X(\update_output_0/n2840 ) );
  nand_x1_sg U9628 ( .A(n4170), .B(n4171), .X(\update_output_0/n2841 ) );
  nand_x1_sg U9629 ( .A(n4127), .B(n4128), .X(\update_output_0/n2842 ) );
  nand_x1_sg U9630 ( .A(n3689), .B(n3690), .X(\update_output_0/n3045 ) );
  nand_x1_sg U9631 ( .A(n3685), .B(n3686), .X(\update_output_0/n3047 ) );
  nand_x1_sg U9632 ( .A(n3681), .B(n3682), .X(\update_output_0/n3049 ) );
  nand_x1_sg U9633 ( .A(n3677), .B(n3678), .X(\update_output_0/n3051 ) );
  nand_x1_sg U9634 ( .A(n3673), .B(n3674), .X(\update_output_0/n3053 ) );
  nand_x1_sg U9635 ( .A(n3669), .B(n3670), .X(\update_output_0/n3055 ) );
  nand_x1_sg U9636 ( .A(n3665), .B(n3666), .X(\update_output_0/n3057 ) );
  nand_x1_sg U9637 ( .A(n3661), .B(n3662), .X(\update_output_0/n3059 ) );
  nand_x1_sg U9638 ( .A(n3657), .B(n3658), .X(\update_output_0/n3061 ) );
  nand_x1_sg U9639 ( .A(n3693), .B(n3694), .X(\update_output_0/n3043 ) );
  nand_x1_sg U9640 ( .A(n3691), .B(n3692), .X(\update_output_0/n3044 ) );
  nand_x1_sg U9641 ( .A(n3687), .B(n3688), .X(\update_output_0/n3046 ) );
  nand_x1_sg U9642 ( .A(n3683), .B(n3684), .X(\update_output_0/n3048 ) );
  nand_x1_sg U9643 ( .A(n3679), .B(n3680), .X(\update_output_0/n3050 ) );
  nand_x1_sg U9644 ( .A(n3675), .B(n3676), .X(\update_output_0/n3052 ) );
  nand_x1_sg U9645 ( .A(n3671), .B(n3672), .X(\update_output_0/n3054 ) );
  nand_x1_sg U9646 ( .A(n3667), .B(n3668), .X(\update_output_0/n3056 ) );
  nand_x1_sg U9647 ( .A(n3663), .B(n3664), .X(\update_output_0/n3058 ) );
  nand_x1_sg U9648 ( .A(n3659), .B(n3660), .X(\update_output_0/n3060 ) );
  nand_x1_sg U9649 ( .A(n3654), .B(n3655), .X(\update_output_0/n3062 ) );
  nand_x1_sg U9650 ( .A(n3823), .B(n3824), .X(\update_output_0/n2983 ) );
  nand_x1_sg U9651 ( .A(n3821), .B(n3822), .X(\update_output_0/n2984 ) );
  nand_x1_sg U9652 ( .A(n3817), .B(n3818), .X(\update_output_0/n2986 ) );
  nand_x1_sg U9653 ( .A(n3813), .B(n3814), .X(\update_output_0/n2988 ) );
  nand_x1_sg U9654 ( .A(n3809), .B(n3810), .X(\update_output_0/n2990 ) );
  nand_x1_sg U9655 ( .A(n3805), .B(n3806), .X(\update_output_0/n2992 ) );
  nand_x1_sg U9656 ( .A(n3801), .B(n3802), .X(\update_output_0/n2994 ) );
  nand_x1_sg U9657 ( .A(n3797), .B(n3798), .X(\update_output_0/n2996 ) );
  nand_x1_sg U9658 ( .A(n3793), .B(n3794), .X(\update_output_0/n2998 ) );
  nand_x1_sg U9659 ( .A(n3789), .B(n3790), .X(\update_output_0/n3000 ) );
  nand_x1_sg U9660 ( .A(n3784), .B(n3785), .X(\update_output_0/n3002 ) );
  nand_x1_sg U9661 ( .A(n3564), .B(n3565), .X(\update_output_0/n3103 ) );
  nand_x1_sg U9662 ( .A(n3562), .B(n3563), .X(\update_output_0/n3104 ) );
  nand_x1_sg U9663 ( .A(n3558), .B(n3559), .X(\update_output_0/n3106 ) );
  nand_x1_sg U9664 ( .A(n3554), .B(n3555), .X(\update_output_0/n3108 ) );
  nand_x1_sg U9665 ( .A(n3550), .B(n3551), .X(\update_output_0/n3110 ) );
  nand_x1_sg U9666 ( .A(n3546), .B(n3547), .X(\update_output_0/n3112 ) );
  nand_x1_sg U9667 ( .A(n3542), .B(n3543), .X(\update_output_0/n3114 ) );
  nand_x1_sg U9668 ( .A(n3538), .B(n3539), .X(\update_output_0/n3116 ) );
  nand_x1_sg U9669 ( .A(n3534), .B(n3535), .X(\update_output_0/n3118 ) );
  nand_x1_sg U9670 ( .A(n3530), .B(n3531), .X(\update_output_0/n3120 ) );
  nand_x1_sg U9671 ( .A(n3525), .B(n3526), .X(\update_output_0/n3122 ) );
  nand_x1_sg U9672 ( .A(n3736), .B(n3737), .X(\update_output_0/n3023 ) );
  nand_x1_sg U9673 ( .A(n3734), .B(n3735), .X(\update_output_0/n3024 ) );
  nand_x1_sg U9674 ( .A(n3732), .B(n3733), .X(\update_output_0/n3025 ) );
  nand_x1_sg U9675 ( .A(n3730), .B(n3731), .X(\update_output_0/n3026 ) );
  nand_x1_sg U9676 ( .A(n3728), .B(n3729), .X(\update_output_0/n3027 ) );
  nand_x1_sg U9677 ( .A(n3726), .B(n3727), .X(\update_output_0/n3028 ) );
  nand_x1_sg U9678 ( .A(n3724), .B(n3725), .X(\update_output_0/n3029 ) );
  nand_x1_sg U9679 ( .A(n3722), .B(n3723), .X(\update_output_0/n3030 ) );
  nand_x1_sg U9680 ( .A(n3720), .B(n3721), .X(\update_output_0/n3031 ) );
  nand_x1_sg U9681 ( .A(n3718), .B(n3719), .X(\update_output_0/n3032 ) );
  nand_x1_sg U9682 ( .A(n3716), .B(n3717), .X(\update_output_0/n3033 ) );
  nand_x1_sg U9683 ( .A(n3714), .B(n3715), .X(\update_output_0/n3034 ) );
  nand_x1_sg U9684 ( .A(n3712), .B(n3713), .X(\update_output_0/n3035 ) );
  nand_x1_sg U9685 ( .A(n3710), .B(n3711), .X(\update_output_0/n3036 ) );
  nand_x1_sg U9686 ( .A(n3708), .B(n3709), .X(\update_output_0/n3037 ) );
  nand_x1_sg U9687 ( .A(n3706), .B(n3707), .X(\update_output_0/n3038 ) );
  nand_x1_sg U9688 ( .A(n3704), .B(n3705), .X(\update_output_0/n3039 ) );
  nand_x1_sg U9689 ( .A(n3702), .B(n3703), .X(\update_output_0/n3040 ) );
  nand_x1_sg U9690 ( .A(n3700), .B(n3701), .X(\update_output_0/n3041 ) );
  nand_x1_sg U9691 ( .A(n3697), .B(n3698), .X(\update_output_0/n3042 ) );
  nand_x1_sg U9692 ( .A(n3819), .B(n3820), .X(\update_output_0/n2985 ) );
  nand_x1_sg U9693 ( .A(n3815), .B(n3816), .X(\update_output_0/n2987 ) );
  nand_x1_sg U9694 ( .A(n3811), .B(n3812), .X(\update_output_0/n2989 ) );
  nand_x1_sg U9695 ( .A(n3807), .B(n3808), .X(\update_output_0/n2991 ) );
  nand_x1_sg U9696 ( .A(n3803), .B(n3804), .X(\update_output_0/n2993 ) );
  nand_x1_sg U9697 ( .A(n3799), .B(n3800), .X(\update_output_0/n2995 ) );
  nand_x1_sg U9698 ( .A(n3795), .B(n3796), .X(\update_output_0/n2997 ) );
  nand_x1_sg U9699 ( .A(n3791), .B(n3792), .X(\update_output_0/n2999 ) );
  nand_x1_sg U9700 ( .A(n3787), .B(n3788), .X(\update_output_0/n3001 ) );
  nand_x1_sg U9701 ( .A(n3560), .B(n3561), .X(\update_output_0/n3105 ) );
  nand_x1_sg U9702 ( .A(n3556), .B(n3557), .X(\update_output_0/n3107 ) );
  nand_x1_sg U9703 ( .A(n3552), .B(n3553), .X(\update_output_0/n3109 ) );
  nand_x1_sg U9704 ( .A(n3548), .B(n3549), .X(\update_output_0/n3111 ) );
  nand_x1_sg U9705 ( .A(n3544), .B(n3545), .X(\update_output_0/n3113 ) );
  nand_x1_sg U9706 ( .A(n3540), .B(n3541), .X(\update_output_0/n3115 ) );
  nand_x1_sg U9707 ( .A(n3536), .B(n3537), .X(\update_output_0/n3117 ) );
  nand_x1_sg U9708 ( .A(n3532), .B(n3533), .X(\update_output_0/n3119 ) );
  nand_x1_sg U9709 ( .A(n3528), .B(n3529), .X(\update_output_0/n3121 ) );
  nand_x1_sg U9710 ( .A(n3607), .B(n3608), .X(\update_output_0/n3083 ) );
  nand_x1_sg U9711 ( .A(n3605), .B(n3606), .X(\update_output_0/n3084 ) );
  nand_x1_sg U9712 ( .A(n3603), .B(n3604), .X(\update_output_0/n3085 ) );
  nand_x1_sg U9713 ( .A(n3601), .B(n3602), .X(\update_output_0/n3086 ) );
  nand_x1_sg U9714 ( .A(n3599), .B(n3600), .X(\update_output_0/n3087 ) );
  nand_x1_sg U9715 ( .A(n3597), .B(n3598), .X(\update_output_0/n3088 ) );
  nand_x1_sg U9716 ( .A(n3595), .B(n3596), .X(\update_output_0/n3089 ) );
  nand_x1_sg U9717 ( .A(n3593), .B(n3594), .X(\update_output_0/n3090 ) );
  nand_x1_sg U9718 ( .A(n3591), .B(n3592), .X(\update_output_0/n3091 ) );
  nand_x1_sg U9719 ( .A(n3589), .B(n3590), .X(\update_output_0/n3092 ) );
  nand_x1_sg U9720 ( .A(n3587), .B(n3588), .X(\update_output_0/n3093 ) );
  nand_x1_sg U9721 ( .A(n3585), .B(n3586), .X(\update_output_0/n3094 ) );
  nand_x1_sg U9722 ( .A(n3583), .B(n3584), .X(\update_output_0/n3095 ) );
  nand_x1_sg U9723 ( .A(n3581), .B(n3582), .X(\update_output_0/n3096 ) );
  nand_x1_sg U9724 ( .A(n3579), .B(n3580), .X(\update_output_0/n3097 ) );
  nand_x1_sg U9725 ( .A(n3577), .B(n3578), .X(\update_output_0/n3098 ) );
  nand_x1_sg U9726 ( .A(n3575), .B(n3576), .X(\update_output_0/n3099 ) );
  nand_x1_sg U9727 ( .A(n3573), .B(n3574), .X(\update_output_0/n3100 ) );
  nand_x1_sg U9728 ( .A(n3571), .B(n3572), .X(\update_output_0/n3101 ) );
  nand_x1_sg U9729 ( .A(n3568), .B(n3569), .X(\update_output_0/n3102 ) );
  nand_x1_sg U9730 ( .A(n3779), .B(n3780), .X(\update_output_0/n3003 ) );
  nand_x1_sg U9731 ( .A(n3777), .B(n3778), .X(\update_output_0/n3004 ) );
  nand_x1_sg U9732 ( .A(n3773), .B(n3774), .X(\update_output_0/n3006 ) );
  nand_x1_sg U9733 ( .A(n3769), .B(n3770), .X(\update_output_0/n3008 ) );
  nand_x1_sg U9734 ( .A(n3765), .B(n3766), .X(\update_output_0/n3010 ) );
  nand_x1_sg U9735 ( .A(n3761), .B(n3762), .X(\update_output_0/n3012 ) );
  nand_x1_sg U9736 ( .A(n3757), .B(n3758), .X(\update_output_0/n3014 ) );
  nand_x1_sg U9737 ( .A(n3753), .B(n3754), .X(\update_output_0/n3016 ) );
  nand_x1_sg U9738 ( .A(n3749), .B(n3750), .X(\update_output_0/n3018 ) );
  nand_x1_sg U9739 ( .A(n3745), .B(n3746), .X(\update_output_0/n3020 ) );
  nand_x1_sg U9740 ( .A(n3740), .B(n3741), .X(\update_output_0/n3022 ) );
  nand_x1_sg U9741 ( .A(n3775), .B(n3776), .X(\update_output_0/n3005 ) );
  nand_x1_sg U9742 ( .A(n3771), .B(n3772), .X(\update_output_0/n3007 ) );
  nand_x1_sg U9743 ( .A(n3767), .B(n3768), .X(\update_output_0/n3009 ) );
  nand_x1_sg U9744 ( .A(n3763), .B(n3764), .X(\update_output_0/n3011 ) );
  nand_x1_sg U9745 ( .A(n3759), .B(n3760), .X(\update_output_0/n3013 ) );
  nand_x1_sg U9746 ( .A(n3755), .B(n3756), .X(\update_output_0/n3015 ) );
  nand_x1_sg U9747 ( .A(n3751), .B(n3752), .X(\update_output_0/n3017 ) );
  nand_x1_sg U9748 ( .A(n3747), .B(n3748), .X(\update_output_0/n3019 ) );
  nand_x1_sg U9749 ( .A(n3743), .B(n3744), .X(\update_output_0/n3021 ) );
  nand_x1_sg U9750 ( .A(n3516), .B(n3517), .X(\update_output_0/n3125 ) );
  nand_x1_sg U9751 ( .A(n3512), .B(n3513), .X(\update_output_0/n3127 ) );
  nand_x1_sg U9752 ( .A(n3508), .B(n3509), .X(\update_output_0/n3129 ) );
  nand_x1_sg U9753 ( .A(n3504), .B(n3505), .X(\update_output_0/n3131 ) );
  nand_x1_sg U9754 ( .A(n3500), .B(n3501), .X(\update_output_0/n3133 ) );
  nand_x1_sg U9755 ( .A(n3496), .B(n3497), .X(\update_output_0/n3135 ) );
  nand_x1_sg U9756 ( .A(n3492), .B(n3493), .X(\update_output_0/n3137 ) );
  nand_x1_sg U9757 ( .A(n3488), .B(n3489), .X(\update_output_0/n3139 ) );
  nand_x1_sg U9758 ( .A(n3484), .B(n3485), .X(\update_output_0/n3141 ) );
  nand_x1_sg U9759 ( .A(n3646), .B(n3647), .X(\update_output_0/n3065 ) );
  nand_x1_sg U9760 ( .A(n3642), .B(n3643), .X(\update_output_0/n3067 ) );
  nand_x1_sg U9761 ( .A(n3638), .B(n3639), .X(\update_output_0/n3069 ) );
  nand_x1_sg U9762 ( .A(n3634), .B(n3635), .X(\update_output_0/n3071 ) );
  nand_x1_sg U9763 ( .A(n3630), .B(n3631), .X(\update_output_0/n3073 ) );
  nand_x1_sg U9764 ( .A(n3626), .B(n3627), .X(\update_output_0/n3075 ) );
  nand_x1_sg U9765 ( .A(n3622), .B(n3623), .X(\update_output_0/n3077 ) );
  nand_x1_sg U9766 ( .A(n3618), .B(n3619), .X(\update_output_0/n3079 ) );
  nand_x1_sg U9767 ( .A(n3614), .B(n3615), .X(\update_output_0/n3081 ) );
  nand_x1_sg U9768 ( .A(n3520), .B(n3521), .X(\update_output_0/n3123 ) );
  nand_x1_sg U9769 ( .A(n3518), .B(n3519), .X(\update_output_0/n3124 ) );
  nand_x1_sg U9770 ( .A(n3514), .B(n3515), .X(\update_output_0/n3126 ) );
  nand_x1_sg U9771 ( .A(n3510), .B(n3511), .X(\update_output_0/n3128 ) );
  nand_x1_sg U9772 ( .A(n3506), .B(n3507), .X(\update_output_0/n3130 ) );
  nand_x1_sg U9773 ( .A(n3502), .B(n3503), .X(\update_output_0/n3132 ) );
  nand_x1_sg U9774 ( .A(n3498), .B(n3499), .X(\update_output_0/n3134 ) );
  nand_x1_sg U9775 ( .A(n3494), .B(n3495), .X(\update_output_0/n3136 ) );
  nand_x1_sg U9776 ( .A(n3490), .B(n3491), .X(\update_output_0/n3138 ) );
  nand_x1_sg U9777 ( .A(n3486), .B(n3487), .X(\update_output_0/n3140 ) );
  nand_x1_sg U9778 ( .A(n3481), .B(n3482), .X(\update_output_0/n3142 ) );
  nand_x1_sg U9779 ( .A(n3650), .B(n3651), .X(\update_output_0/n3063 ) );
  nand_x1_sg U9780 ( .A(n3648), .B(n3649), .X(\update_output_0/n3064 ) );
  nand_x1_sg U9781 ( .A(n3644), .B(n3645), .X(\update_output_0/n3066 ) );
  nand_x1_sg U9782 ( .A(n3640), .B(n3641), .X(\update_output_0/n3068 ) );
  nand_x1_sg U9783 ( .A(n3636), .B(n3637), .X(\update_output_0/n3070 ) );
  nand_x1_sg U9784 ( .A(n3632), .B(n3633), .X(\update_output_0/n3072 ) );
  nand_x1_sg U9785 ( .A(n3628), .B(n3629), .X(\update_output_0/n3074 ) );
  nand_x1_sg U9786 ( .A(n3624), .B(n3625), .X(\update_output_0/n3076 ) );
  nand_x1_sg U9787 ( .A(n3620), .B(n3621), .X(\update_output_0/n3078 ) );
  nand_x1_sg U9788 ( .A(n3616), .B(n3617), .X(\update_output_0/n3080 ) );
  nand_x1_sg U9789 ( .A(n3611), .B(n3612), .X(\update_output_0/n3082 ) );
  inv_x1_sg U9790 ( .A(n995), .X(n8992) );
  inv_x1_sg U9791 ( .A(n1313), .X(n9128) );
  inv_x1_sg U9792 ( .A(n1150), .X(n9123) );
  inv_x1_sg U9793 ( .A(n854), .X(n9138) );
  inv_x1_sg U9794 ( .A(n822), .X(n9137) );
  inv_x1_sg U9795 ( .A(n993), .X(n8972) );
  inv_x1_sg U9796 ( .A(n1182), .X(n9124) );
  inv_x1_sg U9797 ( .A(n1017), .X(n9132) );
  inv_x1_sg U9798 ( .A(n1298), .X(n9008) );
  inv_x1_sg U9799 ( .A(n1281), .X(n9127) );
  inv_x1_sg U9800 ( .A(n985), .X(n9134) );
  inv_x1_sg U9801 ( .A(n1141), .X(n9103) );
  inv_x1_sg U9802 ( .A(n1291), .X(n8988) );
  inv_x1_sg U9803 ( .A(n845), .X(n9118) );
  inv_x1_sg U9804 ( .A(n813), .X(n9117) );
  inv_x1_sg U9805 ( .A(n1257), .X(n8967) );
  inv_x1_sg U9806 ( .A(n1158), .X(n8964) );
  inv_x1_sg U9807 ( .A(n961), .X(n8974) );
  inv_x1_sg U9808 ( .A(n1126), .X(n8963) );
  inv_x1_sg U9809 ( .A(n830), .X(n8978) );
  inv_x1_sg U9810 ( .A(n793), .X(n8977) );
  inv_x1_sg U9811 ( .A(n976), .X(n9114) );
  inv_x1_sg U9812 ( .A(n1355), .X(n8990) );
  inv_x1_sg U9813 ( .A(n1192), .X(n8986) );
  inv_x1_sg U9814 ( .A(n928), .X(n9001) );
  inv_x1_sg U9815 ( .A(n1091), .X(n8996) );
  inv_x1_sg U9816 ( .A(n1409), .X(n9131) );
  inv_x1_sg U9817 ( .A(n1113), .X(n9136) );
  inv_x1_sg U9818 ( .A(n1345), .X(n9129) );
  inv_x1_sg U9819 ( .A(n1377), .X(n9130) );
  inv_x1_sg U9820 ( .A(n1246), .X(n9125) );
  inv_x1_sg U9821 ( .A(n1214), .X(n9126) );
  inv_x1_sg U9822 ( .A(n1081), .X(n9135) );
  inv_x1_sg U9823 ( .A(n1444), .X(n9122) );
  inv_x1_sg U9824 ( .A(n886), .X(n9139) );
  inv_x1_sg U9825 ( .A(n918), .X(n9140) );
  inv_x1_sg U9826 ( .A(n1353), .X(n8970) );
  inv_x1_sg U9827 ( .A(n1394), .X(n9011) );
  inv_x1_sg U9828 ( .A(n1190), .X(n8966) );
  inv_x1_sg U9829 ( .A(n1049), .X(n9133) );
  inv_x1_sg U9830 ( .A(n1330), .X(n9009) );
  inv_x1_sg U9831 ( .A(n926), .X(n8981) );
  inv_x1_sg U9832 ( .A(n1034), .X(n9013) );
  inv_x1_sg U9833 ( .A(n1231), .X(n9005) );
  inv_x1_sg U9834 ( .A(n950), .X(n9141) );
  inv_x1_sg U9835 ( .A(n1089), .X(n8976) );
  inv_x1_sg U9836 ( .A(n1072), .X(n9115) );
  inv_x1_sg U9837 ( .A(n1432), .X(n9102) );
  inv_x1_sg U9838 ( .A(n1387), .X(n8991) );
  inv_x1_sg U9839 ( .A(n909), .X(n9120) );
  inv_x1_sg U9840 ( .A(n877), .X(n9119) );
  inv_x1_sg U9841 ( .A(n1323), .X(n8989) );
  inv_x1_sg U9842 ( .A(n1224), .X(n8985) );
  inv_x1_sg U9843 ( .A(n1027), .X(n8993) );
  inv_x1_sg U9844 ( .A(n1057), .X(n8975) );
  inv_x1_sg U9845 ( .A(n1417), .X(n8962) );
  inv_x1_sg U9846 ( .A(n862), .X(n8979) );
  inv_x1_sg U9847 ( .A(n894), .X(n8980) );
  nand_x1_sg U9848 ( .A(n3467), .B(n3468), .X(\update_output_0/n3145 ) );
  nand_x1_sg U9849 ( .A(n3475), .B(n3476), .X(\update_output_0/n3143 ) );
  nand_x1_sg U9850 ( .A(n9223), .B(n3441), .X(n3440) );
  nand_x1_sg U9851 ( .A(n4858), .B(n4859), .X(\update_output_0/n2822 ) );
  nand_x1_sg U9852 ( .A(n3454), .B(n3455), .X(\update_output_0/n3147 ) );
  nand_x1_sg U9853 ( .A(n4880), .B(n4881), .X(\update_mask_0/n1439 ) );
  nand_x1_sg U9854 ( .A(n4876), .B(n4877), .X(\update_mask_0/n1440 ) );
  nand_x1_sg U9855 ( .A(n4933), .B(n4934), .X(\update_mask_0/n1417 ) );
  nand_x1_sg U9856 ( .A(n4903), .B(n4904), .X(\update_mask_0/n1432 ) );
  nand_x1_sg U9857 ( .A(n5567), .B(n5568), .X(\update_mask_0/n1100 ) );
  nand_x1_sg U9858 ( .A(n5565), .B(n5566), .X(\update_mask_0/n1101 ) );
  nand_x1_sg U9859 ( .A(n5563), .B(n5564), .X(\update_mask_0/n1102 ) );
  nand_x1_sg U9860 ( .A(n5443), .B(n5444), .X(\update_mask_0/n1162 ) );
  nand_x1_sg U9861 ( .A(n5441), .B(n5442), .X(\update_mask_0/n1163 ) );
  nand_x1_sg U9862 ( .A(n5439), .B(n5440), .X(\update_mask_0/n1164 ) );
  nand_x1_sg U9863 ( .A(n5375), .B(n5376), .X(\update_mask_0/n1196 ) );
  nand_x1_sg U9864 ( .A(n5373), .B(n5374), .X(\update_mask_0/n1197 ) );
  nand_x1_sg U9865 ( .A(n5371), .B(n5372), .X(\update_mask_0/n1198 ) );
  nand_x1_sg U9866 ( .A(n5247), .B(n5248), .X(\update_mask_0/n1260 ) );
  nand_x1_sg U9867 ( .A(n5245), .B(n5246), .X(\update_mask_0/n1261 ) );
  nand_x1_sg U9868 ( .A(n5243), .B(n5244), .X(\update_mask_0/n1262 ) );
  nand_x1_sg U9869 ( .A(n5087), .B(n5088), .X(\update_mask_0/n1340 ) );
  nand_x1_sg U9870 ( .A(n5085), .B(n5086), .X(\update_mask_0/n1341 ) );
  nand_x1_sg U9871 ( .A(n5083), .B(n5084), .X(\update_mask_0/n1342 ) );
  nand_x1_sg U9872 ( .A(n5071), .B(n5072), .X(\update_mask_0/n1348 ) );
  nand_x1_sg U9873 ( .A(n5069), .B(n5070), .X(\update_mask_0/n1349 ) );
  nand_x1_sg U9874 ( .A(n5067), .B(n5068), .X(\update_mask_0/n1350 ) );
  nand_x1_sg U9875 ( .A(n4927), .B(n4928), .X(\update_mask_0/n1420 ) );
  nand_x1_sg U9876 ( .A(n4925), .B(n4926), .X(\update_mask_0/n1421 ) );
  nand_x1_sg U9877 ( .A(n4923), .B(n4924), .X(\update_mask_0/n1422 ) );
  nand_x1_sg U9878 ( .A(n5593), .B(n5594), .X(\update_mask_0/n1087 ) );
  nand_x1_sg U9879 ( .A(n5591), .B(n5592), .X(\update_mask_0/n1088 ) );
  nand_x1_sg U9880 ( .A(n5589), .B(n5590), .X(\update_mask_0/n1089 ) );
  nand_x1_sg U9881 ( .A(n5587), .B(n5588), .X(\update_mask_0/n1090 ) );
  nand_x1_sg U9882 ( .A(n5585), .B(n5586), .X(\update_mask_0/n1091 ) );
  nand_x1_sg U9883 ( .A(n5583), .B(n5584), .X(\update_mask_0/n1092 ) );
  nand_x1_sg U9884 ( .A(n5581), .B(n5582), .X(\update_mask_0/n1093 ) );
  nand_x1_sg U9885 ( .A(n5579), .B(n5580), .X(\update_mask_0/n1094 ) );
  nand_x1_sg U9886 ( .A(n5561), .B(n5562), .X(\update_mask_0/n1103 ) );
  nand_x1_sg U9887 ( .A(n5559), .B(n5560), .X(\update_mask_0/n1104 ) );
  nand_x1_sg U9888 ( .A(n5557), .B(n5558), .X(\update_mask_0/n1105 ) );
  nand_x1_sg U9889 ( .A(n5555), .B(n5556), .X(\update_mask_0/n1106 ) );
  nand_x1_sg U9890 ( .A(n5553), .B(n5554), .X(\update_mask_0/n1107 ) );
  nand_x1_sg U9891 ( .A(n5551), .B(n5552), .X(\update_mask_0/n1108 ) );
  nand_x1_sg U9892 ( .A(n5549), .B(n5550), .X(\update_mask_0/n1109 ) );
  nand_x1_sg U9893 ( .A(n5547), .B(n5548), .X(\update_mask_0/n1110 ) );
  nand_x1_sg U9894 ( .A(n5545), .B(n5546), .X(\update_mask_0/n1111 ) );
  nand_x1_sg U9895 ( .A(n5543), .B(n5544), .X(\update_mask_0/n1112 ) );
  nand_x1_sg U9896 ( .A(n5541), .B(n5542), .X(\update_mask_0/n1113 ) );
  nand_x1_sg U9897 ( .A(n5539), .B(n5540), .X(\update_mask_0/n1114 ) );
  nand_x1_sg U9898 ( .A(n5537), .B(n5538), .X(\update_mask_0/n1115 ) );
  nand_x1_sg U9899 ( .A(n5535), .B(n5536), .X(\update_mask_0/n1116 ) );
  nand_x1_sg U9900 ( .A(n5533), .B(n5534), .X(\update_mask_0/n1117 ) );
  nand_x1_sg U9901 ( .A(n5531), .B(n5532), .X(\update_mask_0/n1118 ) );
  nand_x1_sg U9902 ( .A(n5529), .B(n5530), .X(\update_mask_0/n1119 ) );
  nand_x1_sg U9903 ( .A(n5527), .B(n5528), .X(\update_mask_0/n1120 ) );
  nand_x1_sg U9904 ( .A(n5525), .B(n5526), .X(\update_mask_0/n1121 ) );
  nand_x1_sg U9905 ( .A(n5513), .B(n5514), .X(\update_mask_0/n1127 ) );
  nand_x1_sg U9906 ( .A(n5511), .B(n5512), .X(\update_mask_0/n1128 ) );
  nand_x1_sg U9907 ( .A(n5509), .B(n5510), .X(\update_mask_0/n1129 ) );
  nand_x1_sg U9908 ( .A(n5507), .B(n5508), .X(\update_mask_0/n1130 ) );
  nand_x1_sg U9909 ( .A(n5505), .B(n5506), .X(\update_mask_0/n1131 ) );
  nand_x1_sg U9910 ( .A(n5503), .B(n5504), .X(\update_mask_0/n1132 ) );
  nand_x1_sg U9911 ( .A(n5501), .B(n5502), .X(\update_mask_0/n1133 ) );
  nand_x1_sg U9912 ( .A(n5499), .B(n5500), .X(\update_mask_0/n1134 ) );
  nand_x1_sg U9913 ( .A(n5497), .B(n5498), .X(\update_mask_0/n1135 ) );
  nand_x1_sg U9914 ( .A(n5495), .B(n5496), .X(\update_mask_0/n1136 ) );
  nand_x1_sg U9915 ( .A(n5493), .B(n5494), .X(\update_mask_0/n1137 ) );
  nand_x1_sg U9916 ( .A(n5491), .B(n5492), .X(\update_mask_0/n1138 ) );
  nand_x1_sg U9917 ( .A(n5489), .B(n5490), .X(\update_mask_0/n1139 ) );
  nand_x1_sg U9918 ( .A(n5487), .B(n5488), .X(\update_mask_0/n1140 ) );
  nand_x1_sg U9919 ( .A(n5485), .B(n5486), .X(\update_mask_0/n1141 ) );
  nand_x1_sg U9920 ( .A(n5483), .B(n5484), .X(\update_mask_0/n1142 ) );
  nand_x1_sg U9921 ( .A(n5481), .B(n5482), .X(\update_mask_0/n1143 ) );
  nand_x1_sg U9922 ( .A(n5479), .B(n5480), .X(\update_mask_0/n1144 ) );
  nand_x1_sg U9923 ( .A(n5477), .B(n5478), .X(\update_mask_0/n1145 ) );
  nand_x1_sg U9924 ( .A(n5475), .B(n5476), .X(\update_mask_0/n1146 ) );
  nand_x1_sg U9925 ( .A(n5473), .B(n5474), .X(\update_mask_0/n1147 ) );
  nand_x1_sg U9926 ( .A(n5471), .B(n5472), .X(\update_mask_0/n1148 ) );
  nand_x1_sg U9927 ( .A(n5469), .B(n5470), .X(\update_mask_0/n1149 ) );
  nand_x1_sg U9928 ( .A(n5467), .B(n5468), .X(\update_mask_0/n1150 ) );
  nand_x1_sg U9929 ( .A(n5465), .B(n5466), .X(\update_mask_0/n1151 ) );
  nand_x1_sg U9930 ( .A(n5463), .B(n5464), .X(\update_mask_0/n1152 ) );
  nand_x1_sg U9931 ( .A(n5461), .B(n5462), .X(\update_mask_0/n1153 ) );
  nand_x1_sg U9932 ( .A(n5459), .B(n5460), .X(\update_mask_0/n1154 ) );
  nand_x1_sg U9933 ( .A(n5457), .B(n5458), .X(\update_mask_0/n1155 ) );
  nand_x1_sg U9934 ( .A(n5455), .B(n5456), .X(\update_mask_0/n1156 ) );
  nand_x1_sg U9935 ( .A(n5453), .B(n5454), .X(\update_mask_0/n1157 ) );
  nand_x1_sg U9936 ( .A(n5451), .B(n5452), .X(\update_mask_0/n1158 ) );
  nand_x1_sg U9937 ( .A(n5449), .B(n5450), .X(\update_mask_0/n1159 ) );
  nand_x1_sg U9938 ( .A(n5447), .B(n5448), .X(\update_mask_0/n1160 ) );
  nand_x1_sg U9939 ( .A(n5445), .B(n5446), .X(\update_mask_0/n1161 ) );
  nand_x1_sg U9940 ( .A(n5437), .B(n5438), .X(\update_mask_0/n1165 ) );
  nand_x1_sg U9941 ( .A(n5435), .B(n5436), .X(\update_mask_0/n1166 ) );
  nand_x1_sg U9942 ( .A(n5433), .B(n5434), .X(\update_mask_0/n1167 ) );
  nand_x1_sg U9943 ( .A(n5431), .B(n5432), .X(\update_mask_0/n1168 ) );
  nand_x1_sg U9944 ( .A(n5429), .B(n5430), .X(\update_mask_0/n1169 ) );
  nand_x1_sg U9945 ( .A(n5427), .B(n5428), .X(\update_mask_0/n1170 ) );
  nand_x1_sg U9946 ( .A(n5425), .B(n5426), .X(\update_mask_0/n1171 ) );
  nand_x1_sg U9947 ( .A(n5423), .B(n5424), .X(\update_mask_0/n1172 ) );
  nand_x1_sg U9948 ( .A(n5421), .B(n5422), .X(\update_mask_0/n1173 ) );
  nand_x1_sg U9949 ( .A(n5419), .B(n5420), .X(\update_mask_0/n1174 ) );
  nand_x1_sg U9950 ( .A(n5397), .B(n5398), .X(\update_mask_0/n1185 ) );
  nand_x1_sg U9951 ( .A(n5395), .B(n5396), .X(\update_mask_0/n1186 ) );
  nand_x1_sg U9952 ( .A(n5393), .B(n5394), .X(\update_mask_0/n1187 ) );
  nand_x1_sg U9953 ( .A(n5391), .B(n5392), .X(\update_mask_0/n1188 ) );
  nand_x1_sg U9954 ( .A(n5389), .B(n5390), .X(\update_mask_0/n1189 ) );
  nand_x1_sg U9955 ( .A(n5387), .B(n5388), .X(\update_mask_0/n1190 ) );
  nand_x1_sg U9956 ( .A(n5369), .B(n5370), .X(\update_mask_0/n1199 ) );
  nand_x1_sg U9957 ( .A(n5367), .B(n5368), .X(\update_mask_0/n1200 ) );
  nand_x1_sg U9958 ( .A(n5365), .B(n5366), .X(\update_mask_0/n1201 ) );
  nand_x1_sg U9959 ( .A(n5363), .B(n5364), .X(\update_mask_0/n1202 ) );
  nand_x1_sg U9960 ( .A(n5361), .B(n5362), .X(\update_mask_0/n1203 ) );
  nand_x1_sg U9961 ( .A(n5359), .B(n5360), .X(\update_mask_0/n1204 ) );
  nand_x1_sg U9962 ( .A(n5357), .B(n5358), .X(\update_mask_0/n1205 ) );
  nand_x1_sg U9963 ( .A(n5355), .B(n5356), .X(\update_mask_0/n1206 ) );
  nand_x1_sg U9964 ( .A(n5353), .B(n5354), .X(\update_mask_0/n1207 ) );
  nand_x1_sg U9965 ( .A(n5351), .B(n5352), .X(\update_mask_0/n1208 ) );
  nand_x1_sg U9966 ( .A(n5349), .B(n5350), .X(\update_mask_0/n1209 ) );
  nand_x1_sg U9967 ( .A(n5347), .B(n5348), .X(\update_mask_0/n1210 ) );
  nand_x1_sg U9968 ( .A(n5345), .B(n5346), .X(\update_mask_0/n1211 ) );
  nand_x1_sg U9969 ( .A(n5343), .B(n5344), .X(\update_mask_0/n1212 ) );
  nand_x1_sg U9970 ( .A(n5341), .B(n5342), .X(\update_mask_0/n1213 ) );
  nand_x1_sg U9971 ( .A(n5339), .B(n5340), .X(\update_mask_0/n1214 ) );
  nand_x1_sg U9972 ( .A(n5337), .B(n5338), .X(\update_mask_0/n1215 ) );
  nand_x1_sg U9973 ( .A(n5335), .B(n5336), .X(\update_mask_0/n1216 ) );
  nand_x1_sg U9974 ( .A(n5333), .B(n5334), .X(\update_mask_0/n1217 ) );
  nand_x1_sg U9975 ( .A(n5331), .B(n5332), .X(\update_mask_0/n1218 ) );
  nand_x1_sg U9976 ( .A(n5329), .B(n5330), .X(\update_mask_0/n1219 ) );
  nand_x1_sg U9977 ( .A(n5327), .B(n5328), .X(\update_mask_0/n1220 ) );
  nand_x1_sg U9978 ( .A(n5325), .B(n5326), .X(\update_mask_0/n1221 ) );
  nand_x1_sg U9979 ( .A(n5323), .B(n5324), .X(\update_mask_0/n1222 ) );
  nand_x1_sg U9980 ( .A(n5321), .B(n5322), .X(\update_mask_0/n1223 ) );
  nand_x1_sg U9981 ( .A(n5319), .B(n5320), .X(\update_mask_0/n1224 ) );
  nand_x1_sg U9982 ( .A(n5317), .B(n5318), .X(\update_mask_0/n1225 ) );
  nand_x1_sg U9983 ( .A(n5315), .B(n5316), .X(\update_mask_0/n1226 ) );
  nand_x1_sg U9984 ( .A(n5313), .B(n5314), .X(\update_mask_0/n1227 ) );
  nand_x1_sg U9985 ( .A(n5311), .B(n5312), .X(\update_mask_0/n1228 ) );
  nand_x1_sg U9986 ( .A(n5309), .B(n5310), .X(\update_mask_0/n1229 ) );
  nand_x1_sg U9987 ( .A(n5307), .B(n5308), .X(\update_mask_0/n1230 ) );
  nand_x1_sg U9988 ( .A(n5305), .B(n5306), .X(\update_mask_0/n1231 ) );
  nand_x1_sg U9989 ( .A(n5303), .B(n5304), .X(\update_mask_0/n1232 ) );
  nand_x1_sg U9990 ( .A(n5301), .B(n5302), .X(\update_mask_0/n1233 ) );
  nand_x1_sg U9991 ( .A(n5299), .B(n5300), .X(\update_mask_0/n1234 ) );
  nand_x1_sg U9992 ( .A(n5297), .B(n5298), .X(\update_mask_0/n1235 ) );
  nand_x1_sg U9993 ( .A(n5295), .B(n5296), .X(\update_mask_0/n1236 ) );
  nand_x1_sg U9994 ( .A(n5293), .B(n5294), .X(\update_mask_0/n1237 ) );
  nand_x1_sg U9995 ( .A(n5291), .B(n5292), .X(\update_mask_0/n1238 ) );
  nand_x1_sg U9996 ( .A(n5289), .B(n5290), .X(\update_mask_0/n1239 ) );
  nand_x1_sg U9997 ( .A(n5287), .B(n5288), .X(\update_mask_0/n1240 ) );
  nand_x1_sg U9998 ( .A(n5285), .B(n5286), .X(\update_mask_0/n1241 ) );
  nand_x1_sg U9999 ( .A(n5283), .B(n5284), .X(\update_mask_0/n1242 ) );
  nand_x1_sg U10000 ( .A(n5281), .B(n5282), .X(\update_mask_0/n1243 ) );
  nand_x1_sg U10001 ( .A(n5279), .B(n5280), .X(\update_mask_0/n1244 ) );
  nand_x1_sg U10002 ( .A(n5277), .B(n5278), .X(\update_mask_0/n1245 ) );
  nand_x1_sg U10003 ( .A(n5275), .B(n5276), .X(\update_mask_0/n1246 ) );
  nand_x1_sg U10004 ( .A(n5273), .B(n5274), .X(\update_mask_0/n1247 ) );
  nand_x1_sg U10005 ( .A(n5271), .B(n5272), .X(\update_mask_0/n1248 ) );
  nand_x1_sg U10006 ( .A(n5269), .B(n5270), .X(\update_mask_0/n1249 ) );
  nand_x1_sg U10007 ( .A(n5267), .B(n5268), .X(\update_mask_0/n1250 ) );
  nand_x1_sg U10008 ( .A(n5265), .B(n5266), .X(\update_mask_0/n1251 ) );
  nand_x1_sg U10009 ( .A(n5263), .B(n5264), .X(\update_mask_0/n1252 ) );
  nand_x1_sg U10010 ( .A(n5261), .B(n5262), .X(\update_mask_0/n1253 ) );
  nand_x1_sg U10011 ( .A(n5259), .B(n5260), .X(\update_mask_0/n1254 ) );
  nand_x1_sg U10012 ( .A(n5241), .B(n5242), .X(\update_mask_0/n1263 ) );
  nand_x1_sg U10013 ( .A(n5239), .B(n5240), .X(\update_mask_0/n1264 ) );
  nand_x1_sg U10014 ( .A(n5237), .B(n5238), .X(\update_mask_0/n1265 ) );
  nand_x1_sg U10015 ( .A(n5235), .B(n5236), .X(\update_mask_0/n1266 ) );
  nand_x1_sg U10016 ( .A(n5233), .B(n5234), .X(\update_mask_0/n1267 ) );
  nand_x1_sg U10017 ( .A(n5231), .B(n5232), .X(\update_mask_0/n1268 ) );
  nand_x1_sg U10018 ( .A(n5229), .B(n5230), .X(\update_mask_0/n1269 ) );
  nand_x1_sg U10019 ( .A(n5227), .B(n5228), .X(\update_mask_0/n1270 ) );
  nand_x1_sg U10020 ( .A(n5225), .B(n5226), .X(\update_mask_0/n1271 ) );
  nand_x1_sg U10021 ( .A(n5223), .B(n5224), .X(\update_mask_0/n1272 ) );
  nand_x1_sg U10022 ( .A(n5221), .B(n5222), .X(\update_mask_0/n1273 ) );
  nand_x1_sg U10023 ( .A(n5219), .B(n5220), .X(\update_mask_0/n1274 ) );
  nand_x1_sg U10024 ( .A(n5201), .B(n5202), .X(\update_mask_0/n1283 ) );
  nand_x1_sg U10025 ( .A(n5199), .B(n5200), .X(\update_mask_0/n1284 ) );
  nand_x1_sg U10026 ( .A(n5197), .B(n5198), .X(\update_mask_0/n1285 ) );
  nand_x1_sg U10027 ( .A(n5195), .B(n5196), .X(\update_mask_0/n1286 ) );
  nand_x1_sg U10028 ( .A(n5193), .B(n5194), .X(\update_mask_0/n1287 ) );
  nand_x1_sg U10029 ( .A(n5191), .B(n5192), .X(\update_mask_0/n1288 ) );
  nand_x1_sg U10030 ( .A(n5189), .B(n5190), .X(\update_mask_0/n1289 ) );
  nand_x1_sg U10031 ( .A(n5187), .B(n5188), .X(\update_mask_0/n1290 ) );
  nand_x1_sg U10032 ( .A(n5185), .B(n5186), .X(\update_mask_0/n1291 ) );
  nand_x1_sg U10033 ( .A(n5183), .B(n5184), .X(\update_mask_0/n1292 ) );
  nand_x1_sg U10034 ( .A(n5181), .B(n5182), .X(\update_mask_0/n1293 ) );
  nand_x1_sg U10035 ( .A(n5179), .B(n5180), .X(\update_mask_0/n1294 ) );
  nand_x1_sg U10036 ( .A(n5177), .B(n5178), .X(\update_mask_0/n1295 ) );
  nand_x1_sg U10037 ( .A(n5175), .B(n5176), .X(\update_mask_0/n1296 ) );
  nand_x1_sg U10038 ( .A(n5173), .B(n5174), .X(\update_mask_0/n1297 ) );
  nand_x1_sg U10039 ( .A(n5171), .B(n5172), .X(\update_mask_0/n1298 ) );
  nand_x1_sg U10040 ( .A(n5169), .B(n5170), .X(\update_mask_0/n1299 ) );
  nand_x1_sg U10041 ( .A(n5167), .B(n5168), .X(\update_mask_0/n1300 ) );
  nand_x1_sg U10042 ( .A(n5165), .B(n5166), .X(\update_mask_0/n1301 ) );
  nand_x1_sg U10043 ( .A(n5163), .B(n5164), .X(\update_mask_0/n1302 ) );
  nand_x1_sg U10044 ( .A(n5161), .B(n5162), .X(\update_mask_0/n1303 ) );
  nand_x1_sg U10045 ( .A(n5159), .B(n5160), .X(\update_mask_0/n1304 ) );
  nand_x1_sg U10046 ( .A(n5157), .B(n5158), .X(\update_mask_0/n1305 ) );
  nand_x1_sg U10047 ( .A(n5155), .B(n5156), .X(\update_mask_0/n1306 ) );
  nand_x1_sg U10048 ( .A(n5153), .B(n5154), .X(\update_mask_0/n1307 ) );
  nand_x1_sg U10049 ( .A(n5151), .B(n5152), .X(\update_mask_0/n1308 ) );
  nand_x1_sg U10050 ( .A(n5149), .B(n5150), .X(\update_mask_0/n1309 ) );
  nand_x1_sg U10051 ( .A(n5147), .B(n5148), .X(\update_mask_0/n1310 ) );
  nand_x1_sg U10052 ( .A(n5145), .B(n5146), .X(\update_mask_0/n1311 ) );
  nand_x1_sg U10053 ( .A(n5143), .B(n5144), .X(\update_mask_0/n1312 ) );
  nand_x1_sg U10054 ( .A(n5141), .B(n5142), .X(\update_mask_0/n1313 ) );
  nand_x1_sg U10055 ( .A(n5139), .B(n5140), .X(\update_mask_0/n1314 ) );
  nand_x1_sg U10056 ( .A(n5129), .B(n5130), .X(\update_mask_0/n1319 ) );
  nand_x1_sg U10057 ( .A(n5127), .B(n5128), .X(\update_mask_0/n1320 ) );
  nand_x1_sg U10058 ( .A(n5125), .B(n5126), .X(\update_mask_0/n1321 ) );
  nand_x1_sg U10059 ( .A(n5123), .B(n5124), .X(\update_mask_0/n1322 ) );
  nand_x1_sg U10060 ( .A(n5121), .B(n5122), .X(\update_mask_0/n1323 ) );
  nand_x1_sg U10061 ( .A(n5119), .B(n5120), .X(\update_mask_0/n1324 ) );
  nand_x1_sg U10062 ( .A(n5117), .B(n5118), .X(\update_mask_0/n1325 ) );
  nand_x1_sg U10063 ( .A(n5115), .B(n5116), .X(\update_mask_0/n1326 ) );
  nand_x1_sg U10064 ( .A(n5113), .B(n5114), .X(\update_mask_0/n1327 ) );
  nand_x1_sg U10065 ( .A(n5111), .B(n5112), .X(\update_mask_0/n1328 ) );
  nand_x1_sg U10066 ( .A(n5109), .B(n5110), .X(\update_mask_0/n1329 ) );
  nand_x1_sg U10067 ( .A(n5107), .B(n5108), .X(\update_mask_0/n1330 ) );
  nand_x1_sg U10068 ( .A(n5105), .B(n5106), .X(\update_mask_0/n1331 ) );
  nand_x1_sg U10069 ( .A(n5103), .B(n5104), .X(\update_mask_0/n1332 ) );
  nand_x1_sg U10070 ( .A(n5101), .B(n5102), .X(\update_mask_0/n1333 ) );
  nand_x1_sg U10071 ( .A(n5099), .B(n5100), .X(\update_mask_0/n1334 ) );
  nand_x1_sg U10072 ( .A(n5081), .B(n5082), .X(\update_mask_0/n1343 ) );
  nand_x1_sg U10073 ( .A(n5079), .B(n5080), .X(\update_mask_0/n1344 ) );
  nand_x1_sg U10074 ( .A(n5077), .B(n5078), .X(\update_mask_0/n1345 ) );
  nand_x1_sg U10075 ( .A(n5075), .B(n5076), .X(\update_mask_0/n1346 ) );
  nand_x1_sg U10076 ( .A(n5065), .B(n5066), .X(\update_mask_0/n1351 ) );
  nand_x1_sg U10077 ( .A(n5063), .B(n5064), .X(\update_mask_0/n1352 ) );
  nand_x1_sg U10078 ( .A(n5061), .B(n5062), .X(\update_mask_0/n1353 ) );
  nand_x1_sg U10079 ( .A(n5059), .B(n5060), .X(\update_mask_0/n1354 ) );
  nand_x1_sg U10080 ( .A(n5057), .B(n5058), .X(\update_mask_0/n1355 ) );
  nand_x1_sg U10081 ( .A(n5055), .B(n5056), .X(\update_mask_0/n1356 ) );
  nand_x1_sg U10082 ( .A(n5053), .B(n5054), .X(\update_mask_0/n1357 ) );
  nand_x1_sg U10083 ( .A(n5051), .B(n5052), .X(\update_mask_0/n1358 ) );
  nand_x1_sg U10084 ( .A(n5049), .B(n5050), .X(\update_mask_0/n1359 ) );
  nand_x1_sg U10085 ( .A(n5047), .B(n5048), .X(\update_mask_0/n1360 ) );
  nand_x1_sg U10086 ( .A(n5045), .B(n5046), .X(\update_mask_0/n1361 ) );
  nand_x1_sg U10087 ( .A(n5043), .B(n5044), .X(\update_mask_0/n1362 ) );
  nand_x1_sg U10088 ( .A(n5041), .B(n5042), .X(\update_mask_0/n1363 ) );
  nand_x1_sg U10089 ( .A(n5039), .B(n5040), .X(\update_mask_0/n1364 ) );
  nand_x1_sg U10090 ( .A(n5037), .B(n5038), .X(\update_mask_0/n1365 ) );
  nand_x1_sg U10091 ( .A(n5035), .B(n5036), .X(\update_mask_0/n1366 ) );
  nand_x1_sg U10092 ( .A(n5033), .B(n5034), .X(\update_mask_0/n1367 ) );
  nand_x1_sg U10093 ( .A(n5031), .B(n5032), .X(\update_mask_0/n1368 ) );
  nand_x1_sg U10094 ( .A(n5029), .B(n5030), .X(\update_mask_0/n1369 ) );
  nand_x1_sg U10095 ( .A(n5027), .B(n5028), .X(\update_mask_0/n1370 ) );
  nand_x1_sg U10096 ( .A(n5025), .B(n5026), .X(\update_mask_0/n1371 ) );
  nand_x1_sg U10097 ( .A(n5023), .B(n5024), .X(\update_mask_0/n1372 ) );
  nand_x1_sg U10098 ( .A(n5005), .B(n5006), .X(\update_mask_0/n1381 ) );
  nand_x1_sg U10099 ( .A(n5003), .B(n5004), .X(\update_mask_0/n1382 ) );
  nand_x1_sg U10100 ( .A(n5001), .B(n5002), .X(\update_mask_0/n1383 ) );
  nand_x1_sg U10101 ( .A(n4999), .B(n5000), .X(\update_mask_0/n1384 ) );
  nand_x1_sg U10102 ( .A(n4997), .B(n4998), .X(\update_mask_0/n1385 ) );
  nand_x1_sg U10103 ( .A(n4995), .B(n4996), .X(\update_mask_0/n1386 ) );
  nand_x1_sg U10104 ( .A(n4993), .B(n4994), .X(\update_mask_0/n1387 ) );
  nand_x1_sg U10105 ( .A(n4991), .B(n4992), .X(\update_mask_0/n1388 ) );
  nand_x1_sg U10106 ( .A(n4989), .B(n4990), .X(\update_mask_0/n1389 ) );
  nand_x1_sg U10107 ( .A(n4987), .B(n4988), .X(\update_mask_0/n1390 ) );
  nand_x1_sg U10108 ( .A(n4985), .B(n4986), .X(\update_mask_0/n1391 ) );
  nand_x1_sg U10109 ( .A(n4983), .B(n4984), .X(\update_mask_0/n1392 ) );
  nand_x1_sg U10110 ( .A(n4981), .B(n4982), .X(\update_mask_0/n1393 ) );
  nand_x1_sg U10111 ( .A(n4979), .B(n4980), .X(\update_mask_0/n1394 ) );
  nand_x1_sg U10112 ( .A(n4977), .B(n4978), .X(\update_mask_0/n1395 ) );
  nand_x1_sg U10113 ( .A(n4975), .B(n4976), .X(\update_mask_0/n1396 ) );
  nand_x1_sg U10114 ( .A(n4973), .B(n4974), .X(\update_mask_0/n1397 ) );
  nand_x1_sg U10115 ( .A(n4971), .B(n4972), .X(\update_mask_0/n1398 ) );
  nand_x1_sg U10116 ( .A(n4969), .B(n4970), .X(\update_mask_0/n1399 ) );
  nand_x1_sg U10117 ( .A(n4967), .B(n4968), .X(\update_mask_0/n1400 ) );
  nand_x1_sg U10118 ( .A(n4965), .B(n4966), .X(\update_mask_0/n1401 ) );
  nand_x1_sg U10119 ( .A(n4963), .B(n4964), .X(\update_mask_0/n1402 ) );
  nand_x1_sg U10120 ( .A(n4961), .B(n4962), .X(\update_mask_0/n1403 ) );
  nand_x1_sg U10121 ( .A(n4959), .B(n4960), .X(\update_mask_0/n1404 ) );
  nand_x1_sg U10122 ( .A(n4957), .B(n4958), .X(\update_mask_0/n1405 ) );
  nand_x1_sg U10123 ( .A(n4955), .B(n4956), .X(\update_mask_0/n1406 ) );
  nand_x1_sg U10124 ( .A(n4953), .B(n4954), .X(\update_mask_0/n1407 ) );
  nand_x1_sg U10125 ( .A(n4951), .B(n4952), .X(\update_mask_0/n1408 ) );
  nand_x1_sg U10126 ( .A(n4949), .B(n4950), .X(\update_mask_0/n1409 ) );
  nand_x1_sg U10127 ( .A(n4947), .B(n4948), .X(\update_mask_0/n1410 ) );
  nand_x1_sg U10128 ( .A(n4945), .B(n4946), .X(\update_mask_0/n1411 ) );
  nand_x1_sg U10129 ( .A(n4943), .B(n4944), .X(\update_mask_0/n1412 ) );
  nand_x1_sg U10130 ( .A(n4941), .B(n4942), .X(\update_mask_0/n1413 ) );
  nand_x1_sg U10131 ( .A(n4939), .B(n4940), .X(\update_mask_0/n1414 ) );
  nand_x1_sg U10132 ( .A(n4921), .B(n4922), .X(\update_mask_0/n1423 ) );
  nand_x1_sg U10133 ( .A(n4919), .B(n4920), .X(\update_mask_0/n1424 ) );
  nand_x1_sg U10134 ( .A(n4917), .B(n4918), .X(\update_mask_0/n1425 ) );
  nand_x1_sg U10135 ( .A(n4915), .B(n4916), .X(\update_mask_0/n1426 ) );
  nand_x1_sg U10136 ( .A(n4913), .B(n4914), .X(\update_mask_0/n1427 ) );
  nand_x1_sg U10137 ( .A(n4911), .B(n4912), .X(\update_mask_0/n1428 ) );
  nand_x1_sg U10138 ( .A(n4909), .B(n4910), .X(\update_mask_0/n1429 ) );
  nand_x1_sg U10139 ( .A(n4907), .B(n4908), .X(\update_mask_0/n1430 ) );
  nand_x1_sg U10140 ( .A(n4905), .B(n4906), .X(\update_mask_0/n1431 ) );
  nand_x1_sg U10141 ( .A(n4901), .B(n4902), .X(\update_mask_0/n1433 ) );
  nand_x1_sg U10142 ( .A(n4899), .B(n4900), .X(\update_mask_0/n1434 ) );
  nand_x1_sg U10143 ( .A(n4897), .B(n4898), .X(\update_mask_0/n1435 ) );
  nand_x1_sg U10144 ( .A(n4895), .B(n4896), .X(\update_mask_0/n1436 ) );
  nand_x1_sg U10145 ( .A(n4893), .B(n4894), .X(\update_mask_0/n1437 ) );
  nand_x1_sg U10146 ( .A(n4889), .B(n4890), .X(\update_mask_0/n1438 ) );
  nand_x1_sg U10147 ( .A(n5577), .B(n5578), .X(\update_mask_0/n1095 ) );
  nand_x1_sg U10148 ( .A(n5575), .B(n5576), .X(\update_mask_0/n1096 ) );
  nand_x1_sg U10149 ( .A(n5573), .B(n5574), .X(\update_mask_0/n1097 ) );
  nand_x1_sg U10150 ( .A(n5571), .B(n5572), .X(\update_mask_0/n1098 ) );
  nand_x1_sg U10151 ( .A(n5569), .B(n5570), .X(\update_mask_0/n1099 ) );
  nand_x1_sg U10152 ( .A(n5523), .B(n5524), .X(\update_mask_0/n1122 ) );
  nand_x1_sg U10153 ( .A(n5521), .B(n5522), .X(\update_mask_0/n1123 ) );
  nand_x1_sg U10154 ( .A(n5519), .B(n5520), .X(\update_mask_0/n1124 ) );
  nand_x1_sg U10155 ( .A(n5517), .B(n5518), .X(\update_mask_0/n1125 ) );
  nand_x1_sg U10156 ( .A(n5515), .B(n5516), .X(\update_mask_0/n1126 ) );
  nand_x1_sg U10157 ( .A(n5417), .B(n5418), .X(\update_mask_0/n1175 ) );
  nand_x1_sg U10158 ( .A(n5415), .B(n5416), .X(\update_mask_0/n1176 ) );
  nand_x1_sg U10159 ( .A(n5385), .B(n5386), .X(\update_mask_0/n1191 ) );
  nand_x1_sg U10160 ( .A(n5383), .B(n5384), .X(\update_mask_0/n1192 ) );
  nand_x1_sg U10161 ( .A(n5381), .B(n5382), .X(\update_mask_0/n1193 ) );
  nand_x1_sg U10162 ( .A(n5379), .B(n5380), .X(\update_mask_0/n1194 ) );
  nand_x1_sg U10163 ( .A(n5377), .B(n5378), .X(\update_mask_0/n1195 ) );
  nand_x1_sg U10164 ( .A(n5257), .B(n5258), .X(\update_mask_0/n1255 ) );
  nand_x1_sg U10165 ( .A(n5255), .B(n5256), .X(\update_mask_0/n1256 ) );
  nand_x1_sg U10166 ( .A(n5253), .B(n5254), .X(\update_mask_0/n1257 ) );
  nand_x1_sg U10167 ( .A(n5251), .B(n5252), .X(\update_mask_0/n1258 ) );
  nand_x1_sg U10168 ( .A(n5249), .B(n5250), .X(\update_mask_0/n1259 ) );
  nand_x1_sg U10169 ( .A(n5137), .B(n5138), .X(\update_mask_0/n1315 ) );
  nand_x1_sg U10170 ( .A(n5135), .B(n5136), .X(\update_mask_0/n1316 ) );
  nand_x1_sg U10171 ( .A(n5133), .B(n5134), .X(\update_mask_0/n1317 ) );
  nand_x1_sg U10172 ( .A(n5131), .B(n5132), .X(\update_mask_0/n1318 ) );
  nand_x1_sg U10173 ( .A(n5097), .B(n5098), .X(\update_mask_0/n1335 ) );
  nand_x1_sg U10174 ( .A(n5095), .B(n5096), .X(\update_mask_0/n1336 ) );
  nand_x1_sg U10175 ( .A(n5093), .B(n5094), .X(\update_mask_0/n1337 ) );
  nand_x1_sg U10176 ( .A(n5091), .B(n5092), .X(\update_mask_0/n1338 ) );
  nand_x1_sg U10177 ( .A(n5089), .B(n5090), .X(\update_mask_0/n1339 ) );
  nand_x1_sg U10178 ( .A(n5073), .B(n5074), .X(\update_mask_0/n1347 ) );
  nand_x1_sg U10179 ( .A(n4937), .B(n4938), .X(\update_mask_0/n1415 ) );
  nand_x1_sg U10180 ( .A(n4935), .B(n4936), .X(\update_mask_0/n1416 ) );
  nand_x1_sg U10181 ( .A(n4931), .B(n4932), .X(\update_mask_0/n1418 ) );
  nand_x1_sg U10182 ( .A(n4929), .B(n4930), .X(\update_mask_0/n1419 ) );
  nand_x1_sg U10183 ( .A(n5407), .B(n5408), .X(\update_mask_0/n1180 ) );
  nand_x1_sg U10184 ( .A(n5405), .B(n5406), .X(\update_mask_0/n1181 ) );
  nand_x1_sg U10185 ( .A(n5403), .B(n5404), .X(\update_mask_0/n1182 ) );
  nand_x1_sg U10186 ( .A(n5401), .B(n5402), .X(\update_mask_0/n1183 ) );
  nand_x1_sg U10187 ( .A(n5399), .B(n5400), .X(\update_mask_0/n1184 ) );
  nand_x1_sg U10188 ( .A(n5217), .B(n5218), .X(\update_mask_0/n1275 ) );
  nand_x1_sg U10189 ( .A(n5215), .B(n5216), .X(\update_mask_0/n1276 ) );
  nand_x1_sg U10190 ( .A(n5213), .B(n5214), .X(\update_mask_0/n1277 ) );
  nand_x1_sg U10191 ( .A(n5211), .B(n5212), .X(\update_mask_0/n1278 ) );
  nand_x1_sg U10192 ( .A(n5209), .B(n5210), .X(\update_mask_0/n1279 ) );
  nand_x1_sg U10193 ( .A(n5207), .B(n5208), .X(\update_mask_0/n1280 ) );
  nand_x1_sg U10194 ( .A(n5205), .B(n5206), .X(\update_mask_0/n1281 ) );
  nand_x1_sg U10195 ( .A(n5203), .B(n5204), .X(\update_mask_0/n1282 ) );
  nand_x1_sg U10196 ( .A(n5021), .B(n5022), .X(\update_mask_0/n1373 ) );
  nand_x1_sg U10197 ( .A(n5019), .B(n5020), .X(\update_mask_0/n1374 ) );
  nand_x1_sg U10198 ( .A(n5017), .B(n5018), .X(\update_mask_0/n1375 ) );
  nand_x1_sg U10199 ( .A(n5015), .B(n5016), .X(\update_mask_0/n1376 ) );
  nand_x1_sg U10200 ( .A(n5013), .B(n5014), .X(\update_mask_0/n1377 ) );
  nand_x1_sg U10201 ( .A(n5011), .B(n5012), .X(\update_mask_0/n1378 ) );
  nand_x1_sg U10202 ( .A(n5009), .B(n5010), .X(\update_mask_0/n1379 ) );
  nand_x1_sg U10203 ( .A(n5007), .B(n5008), .X(\update_mask_0/n1380 ) );
  nand_x1_sg U10204 ( .A(n5413), .B(n5414), .X(\update_mask_0/n1177 ) );
  nand_x1_sg U10205 ( .A(n5411), .B(n5412), .X(\update_mask_0/n1178 ) );
  nand_x1_sg U10206 ( .A(n5409), .B(n5410), .X(\update_mask_0/n1179 ) );
  nand_x1_sg U10207 ( .A(n4868), .B(n4869), .X(\update_mask_0/n1441 ) );
  nand_x2_sg U10208 ( .A(n4870), .B(n4871), .X(n4869) );
  nand_x1_sg U10209 ( .A(n5599), .B(n5600), .X(\update_mask_0/n1085 ) );
  inv_x1_sg U10210 ( .A(n5601), .X(n9229) );
  nand_x1_sg U10211 ( .A(n5603), .B(n5604), .X(\update_mask_0/n1084 ) );
  nand_x1_sg U10212 ( .A(n5618), .B(n5619), .X(\update_mask_0/n1081 ) );
  nand_x1_sg U10213 ( .A(n5627), .B(n5628), .X(n5911) );
  nand_x1_sg U10214 ( .A(n5615), .B(n5616), .X(\update_mask_0/n1082 ) );
  nand_x1_sg U10215 ( .A(n3444), .B(n3445), .X(\update_output_0/n3149 ) );
  inv_x1_sg U10216 ( .A(n1678), .X(n8905) );
  inv_x1_sg U10217 ( .A(n2016), .X(n8911) );
  inv_x1_sg U10218 ( .A(n1644), .X(n8942) );
  inv_x1_sg U10219 ( .A(n1661), .X(n8943) );
  inv_x1_sg U10220 ( .A(n1982), .X(n8952) );
  inv_x1_sg U10221 ( .A(n1999), .X(n8953) );
  inv_x1_sg U10222 ( .A(n1563), .X(n8903) );
  inv_x1_sg U10223 ( .A(n1580), .X(n8904) );
  inv_x1_sg U10224 ( .A(n1731), .X(n8906) );
  inv_x1_sg U10225 ( .A(n1748), .X(n8907) );
  inv_x1_sg U10226 ( .A(n1901), .X(n8909) );
  inv_x1_sg U10227 ( .A(n1918), .X(n8910) );
  inv_x1_sg U10228 ( .A(n2069), .X(n8912) );
  inv_x1_sg U10229 ( .A(n2086), .X(n8913) );
  inv_x1_sg U10230 ( .A(n1846), .X(n8908) );
  inv_x1_sg U10231 ( .A(n2185), .X(n8914) );
  inv_x1_sg U10232 ( .A(n2258), .X(n8900) );
  inv_x1_sg U10233 ( .A(n2222), .X(n8899) );
  inv_x1_sg U10234 ( .A(n1778), .X(n8918) );
  inv_x1_sg U10235 ( .A(n2116), .X(n8922) );
  inv_x1_sg U10236 ( .A(n1774), .X(n8929) );
  inv_x1_sg U10237 ( .A(n2112), .X(n8937) );
  inv_x1_sg U10238 ( .A(n1593), .X(n8940) );
  inv_x1_sg U10239 ( .A(n1761), .X(n8945) );
  inv_x1_sg U10240 ( .A(n1812), .X(n8947) );
  inv_x1_sg U10241 ( .A(n1829), .X(n8948) );
  inv_x1_sg U10242 ( .A(n1931), .X(n8950) );
  inv_x1_sg U10243 ( .A(n2099), .X(n8955) );
  inv_x1_sg U10244 ( .A(n2150), .X(n8957) );
  inv_x1_sg U10245 ( .A(n2167), .X(n8958) );
  nand_x4_sg U10246 ( .A(n4398), .B(n4399), .X(n4394) );
  nand_x4_sg U10247 ( .A(n4362), .B(n4363), .X(n4358) );
  nand_x4_sg U10248 ( .A(n4326), .B(n4327), .X(n4322) );
  nand_x4_sg U10249 ( .A(n4290), .B(n4291), .X(n4286) );
  inv_x1_sg U10250 ( .A(n777), .X(n9222) );
  nand_x4_sg U10251 ( .A(n782), .B(n783), .X(n781) );
  nand_x1_sg U10252 ( .A(n6831), .B(n7451), .X(n7473) );
  nand_x1_sg U10253 ( .A(n3653), .B(n6315), .X(n3652) );
  nand_x1_sg U10254 ( .A(n3610), .B(n3524), .X(n3609) );
  nand_x1_sg U10255 ( .A(n3610), .B(n7408), .X(n3953) );
  nand_x1_sg U10256 ( .A(n3653), .B(n7408), .X(n3996) );
  nand_x1_sg U10257 ( .A(n756), .B(n8894), .X(n757) );
  nand_x1_sg U10258 ( .A(n767), .B(n8894), .X(n769) );
  nor_x1_sg U10259 ( .A(n6716), .B(n7105), .X(\update_output_0/n2819 ) );
  nor_x1_sg U10260 ( .A(n6724), .B(n6182), .X(\update_output_0/n2815 ) );
  nor_x1_sg U10261 ( .A(n6692), .B(n7103), .X(\update_output_0/n2803 ) );
  nor_x1_sg U10262 ( .A(n6695), .B(n6182), .X(\update_output_0/n2799 ) );
  nor_x1_sg U10263 ( .A(n6706), .B(n7106), .X(\update_output_0/n2783 ) );
  nor_x1_sg U10264 ( .A(n6720), .B(n6431), .X(\update_output_0/n2775 ) );
  nor_x1_sg U10265 ( .A(n6700), .B(n6019), .X(\update_output_0/n2763 ) );
  nor_x1_sg U10266 ( .A(n6712), .B(n7104), .X(\update_output_0/n2759 ) );
  nor_x1_sg U10267 ( .A(n6714), .B(n7181), .X(\update_output_0/n2739 ) );
  nor_x1_sg U10268 ( .A(n6725), .B(n6047), .X(\update_output_0/n2735 ) );
  nor_x1_sg U10269 ( .A(n6693), .B(n6047), .X(\update_output_0/n2723 ) );
  nor_x1_sg U10270 ( .A(n6696), .B(n6206), .X(\update_output_0/n2719 ) );
  nor_x1_sg U10271 ( .A(n6704), .B(n7179), .X(\update_output_0/n2703 ) );
  nor_x1_sg U10272 ( .A(n6721), .B(n6207), .X(\update_output_0/n2695 ) );
  nor_x1_sg U10273 ( .A(n6699), .B(n7179), .X(\update_output_0/n2683 ) );
  nor_x1_sg U10274 ( .A(n6709), .B(n7182), .X(\update_output_0/n2679 ) );
  nor_x1_sg U10275 ( .A(n6717), .B(n6398), .X(\update_output_0/n2659 ) );
  nor_x1_sg U10276 ( .A(n6725), .B(n7219), .X(\update_output_0/n2655 ) );
  nor_x1_sg U10277 ( .A(n5915), .B(n7222), .X(\update_output_0/n2643 ) );
  nor_x1_sg U10278 ( .A(n6696), .B(n7221), .X(\update_output_0/n2639 ) );
  nor_x1_sg U10279 ( .A(n6705), .B(n6397), .X(\update_output_0/n2623 ) );
  nor_x1_sg U10280 ( .A(n6720), .B(n6397), .X(\update_output_0/n2615 ) );
  nor_x1_sg U10281 ( .A(n6702), .B(n6070), .X(\update_output_0/n2603 ) );
  nor_x1_sg U10282 ( .A(n6712), .B(n6397), .X(\update_output_0/n2599 ) );
  nor_x1_sg U10283 ( .A(n6714), .B(n6415), .X(\update_output_0/n2579 ) );
  nor_x1_sg U10284 ( .A(n6727), .B(n7176), .X(\update_output_0/n2575 ) );
  nor_x1_sg U10285 ( .A(n6693), .B(n6204), .X(\update_output_0/n2563 ) );
  nor_x1_sg U10286 ( .A(n6697), .B(n6204), .X(\update_output_0/n2559 ) );
  nor_x1_sg U10287 ( .A(n6707), .B(n6415), .X(\update_output_0/n2543 ) );
  nor_x1_sg U10288 ( .A(n6719), .B(n6043), .X(\update_output_0/n2535 ) );
  nor_x1_sg U10289 ( .A(n6702), .B(n6044), .X(\update_output_0/n2523 ) );
  nor_x1_sg U10290 ( .A(n6711), .B(n7177), .X(\update_output_0/n2519 ) );
  nor_x1_sg U10291 ( .A(n6715), .B(n7120), .X(\update_output_0/n2499 ) );
  nor_x1_sg U10292 ( .A(n6726), .B(n6425), .X(\update_output_0/n2495 ) );
  nor_x1_sg U10293 ( .A(n6692), .B(n6028), .X(\update_output_0/n2483 ) );
  nor_x1_sg U10294 ( .A(n6697), .B(n7120), .X(\update_output_0/n2479 ) );
  nor_x1_sg U10295 ( .A(n6706), .B(n6191), .X(\update_output_0/n2463 ) );
  nor_x1_sg U10296 ( .A(n6719), .B(n7118), .X(\update_output_0/n2455 ) );
  nor_x1_sg U10297 ( .A(n6701), .B(n6426), .X(\update_output_0/n2443 ) );
  nor_x1_sg U10298 ( .A(n6712), .B(n6029), .X(\update_output_0/n2439 ) );
  nor_x1_sg U10299 ( .A(n6716), .B(n7211), .X(\update_output_0/n2419 ) );
  nor_x1_sg U10300 ( .A(n6726), .B(n7211), .X(\update_output_0/n2415 ) );
  nor_x1_sg U10301 ( .A(n6694), .B(n6225), .X(\update_output_0/n2403 ) );
  nor_x1_sg U10302 ( .A(n6763), .B(n6224), .X(\update_output_0/n2399 ) );
  nor_x1_sg U10303 ( .A(n6706), .B(n6224), .X(\update_output_0/n2383 ) );
  nor_x1_sg U10304 ( .A(n6722), .B(n6064), .X(\update_output_0/n2375 ) );
  nor_x1_sg U10305 ( .A(n6702), .B(n6401), .X(\update_output_0/n2363 ) );
  nor_x1_sg U10306 ( .A(n6711), .B(n7212), .X(\update_output_0/n2359 ) );
  nor_x1_sg U10307 ( .A(n6715), .B(n6061), .X(\update_output_0/n2339 ) );
  nor_x1_sg U10308 ( .A(n6724), .B(n7204), .X(\update_output_0/n2335 ) );
  nor_x1_sg U10309 ( .A(n6748), .B(n6404), .X(\update_output_0/n2323 ) );
  nor_x1_sg U10310 ( .A(n5913), .B(n6061), .X(\update_output_0/n2319 ) );
  nor_x1_sg U10311 ( .A(n6707), .B(n6062), .X(\update_output_0/n2303 ) );
  nor_x1_sg U10312 ( .A(n6721), .B(n6061), .X(\update_output_0/n2295 ) );
  nor_x1_sg U10313 ( .A(n6701), .B(n6222), .X(\update_output_0/n2283 ) );
  nor_x1_sg U10314 ( .A(n6711), .B(n6062), .X(\update_output_0/n2279 ) );
  nor_x1_sg U10315 ( .A(n6715), .B(n7201), .X(\update_output_0/n2259 ) );
  nor_x1_sg U10316 ( .A(n6725), .B(n6059), .X(\update_output_0/n2255 ) );
  nor_x1_sg U10317 ( .A(n6692), .B(n6059), .X(\update_output_0/n2243 ) );
  nor_x1_sg U10318 ( .A(n6695), .B(n6218), .X(\update_output_0/n2239 ) );
  nor_x1_sg U10319 ( .A(n6707), .B(n7199), .X(\update_output_0/n2223 ) );
  nor_x1_sg U10320 ( .A(n6721), .B(n6219), .X(\update_output_0/n2215 ) );
  nor_x1_sg U10321 ( .A(n6701), .B(n7199), .X(\update_output_0/n2203 ) );
  nor_x1_sg U10322 ( .A(n6710), .B(n7202), .X(\update_output_0/n2199 ) );
  nor_x1_sg U10323 ( .A(n6716), .B(n6188), .X(\update_output_0/n2179 ) );
  nor_x1_sg U10324 ( .A(n6724), .B(n7114), .X(\update_output_0/n2175 ) );
  nor_x1_sg U10325 ( .A(n6693), .B(n6428), .X(\update_output_0/n2163 ) );
  nor_x1_sg U10326 ( .A(n6695), .B(n6427), .X(\update_output_0/n2159 ) );
  nor_x1_sg U10327 ( .A(n6706), .B(n7115), .X(\update_output_0/n2143 ) );
  nor_x1_sg U10328 ( .A(n6722), .B(n7116), .X(\update_output_0/n2135 ) );
  nor_x1_sg U10329 ( .A(n6700), .B(n7113), .X(\update_output_0/n2123 ) );
  nor_x1_sg U10330 ( .A(n6712), .B(n6189), .X(\update_output_0/n2119 ) );
  nor_x1_sg U10331 ( .A(n6714), .B(n6040), .X(\update_output_0/n2099 ) );
  nor_x1_sg U10332 ( .A(n6726), .B(n7169), .X(\update_output_0/n2095 ) );
  nor_x1_sg U10333 ( .A(n6694), .B(n6418), .X(\update_output_0/n2083 ) );
  nor_x1_sg U10334 ( .A(n6697), .B(n6040), .X(\update_output_0/n2079 ) );
  nor_x1_sg U10335 ( .A(n6704), .B(n6041), .X(\update_output_0/n2063 ) );
  nor_x1_sg U10336 ( .A(n6720), .B(n6040), .X(\update_output_0/n2055 ) );
  nor_x1_sg U10337 ( .A(n6699), .B(n6201), .X(\update_output_0/n2043 ) );
  nor_x1_sg U10338 ( .A(n6710), .B(n6041), .X(\update_output_0/n2039 ) );
  nor_x1_sg U10339 ( .A(n6717), .B(n6228), .X(\update_output_0/n2019 ) );
  nor_x1_sg U10340 ( .A(n6724), .B(n6400), .X(\update_output_0/n2015 ) );
  nor_x1_sg U10341 ( .A(n6693), .B(n6399), .X(\update_output_0/n2003 ) );
  nor_x1_sg U10342 ( .A(n6696), .B(n7217), .X(\update_output_0/n1999 ) );
  nor_x1_sg U10343 ( .A(n6704), .B(n7215), .X(\update_output_0/n1983 ) );
  nor_x1_sg U10344 ( .A(n6722), .B(n6399), .X(\update_output_0/n1975 ) );
  nor_x1_sg U10345 ( .A(n6700), .B(n6228), .X(\update_output_0/n1963 ) );
  nor_x1_sg U10346 ( .A(n6709), .B(n6067), .X(\update_output_0/n1959 ) );
  nor_x1_sg U10347 ( .A(n6714), .B(n6198), .X(\update_output_0/n1939 ) );
  nor_x1_sg U10348 ( .A(n6727), .B(n6037), .X(\update_output_0/n1935 ) );
  nor_x1_sg U10349 ( .A(n6748), .B(n6037), .X(\update_output_0/n1923 ) );
  nor_x1_sg U10350 ( .A(n6696), .B(n6419), .X(\update_output_0/n1919 ) );
  nor_x1_sg U10351 ( .A(n6704), .B(n6038), .X(\update_output_0/n1903 ) );
  nor_x1_sg U10352 ( .A(n6719), .B(n6038), .X(\update_output_0/n1895 ) );
  nor_x1_sg U10353 ( .A(n6702), .B(n6197), .X(\update_output_0/n1883 ) );
  nor_x1_sg U10354 ( .A(n6711), .B(n6197), .X(\update_output_0/n1879 ) );
  nor_x1_sg U10355 ( .A(n6717), .B(n6022), .X(\update_output_0/n1859 ) );
  nor_x1_sg U10356 ( .A(n6726), .B(n7108), .X(\update_output_0/n1855 ) );
  nor_x1_sg U10357 ( .A(n6692), .B(n6430), .X(\update_output_0/n1843 ) );
  nor_x1_sg U10358 ( .A(n6695), .B(n6022), .X(\update_output_0/n1839 ) );
  nor_x1_sg U10359 ( .A(n6707), .B(n6023), .X(\update_output_0/n1823 ) );
  nor_x1_sg U10360 ( .A(n6720), .B(n6022), .X(\update_output_0/n1815 ) );
  nor_x1_sg U10361 ( .A(n6699), .B(n6186), .X(\update_output_0/n1803 ) );
  nor_x1_sg U10362 ( .A(n6710), .B(n6023), .X(\update_output_0/n1799 ) );
  nor_x1_sg U10363 ( .A(n6716), .B(n6056), .X(\update_output_0/n1779 ) );
  nor_x1_sg U10364 ( .A(n6727), .B(n7194), .X(\update_output_0/n1775 ) );
  nor_x1_sg U10365 ( .A(n6694), .B(n7196), .X(\update_output_0/n1763 ) );
  nor_x1_sg U10366 ( .A(n6763), .B(n6055), .X(\update_output_0/n1759 ) );
  nor_x1_sg U10367 ( .A(n6705), .B(n6215), .X(\update_output_0/n1743 ) );
  nor_x1_sg U10368 ( .A(n6719), .B(n6056), .X(\update_output_0/n1735 ) );
  nor_x1_sg U10369 ( .A(n6699), .B(n7195), .X(\update_output_0/n1723 ) );
  nor_x1_sg U10370 ( .A(n6709), .B(n7195), .X(\update_output_0/n1719 ) );
  nor_x1_sg U10371 ( .A(n6717), .B(n7190), .X(\update_output_0/n1699 ) );
  nor_x1_sg U10372 ( .A(n6725), .B(n6409), .X(\update_output_0/n1695 ) );
  nor_x1_sg U10373 ( .A(n6694), .B(n6410), .X(\update_output_0/n1683 ) );
  nor_x1_sg U10374 ( .A(n6697), .B(n6213), .X(\update_output_0/n1679 ) );
  nor_x1_sg U10375 ( .A(n6705), .B(n7191), .X(\update_output_0/n1663 ) );
  nor_x1_sg U10376 ( .A(n6722), .B(n6212), .X(\update_output_0/n1655 ) );
  nor_x1_sg U10377 ( .A(n6701), .B(n6052), .X(\update_output_0/n1643 ) );
  nor_x1_sg U10378 ( .A(n6710), .B(n7190), .X(\update_output_0/n1639 ) );
  nor_x1_sg U10379 ( .A(n6715), .B(n7186), .X(\update_output_0/n1619 ) );
  nor_x1_sg U10380 ( .A(n6727), .B(n7184), .X(\update_output_0/n1615 ) );
  nor_x1_sg U10381 ( .A(n5915), .B(n6050), .X(\update_output_0/n1603 ) );
  nor_x1_sg U10382 ( .A(n5913), .B(n7184), .X(\update_output_0/n1599 ) );
  nor_x1_sg U10383 ( .A(n6705), .B(n7186), .X(\update_output_0/n1583 ) );
  nor_x1_sg U10384 ( .A(n6721), .B(n6049), .X(\update_output_0/n1575 ) );
  nor_x1_sg U10385 ( .A(n6700), .B(n6210), .X(\update_output_0/n1563 ) );
  nor_x1_sg U10386 ( .A(n6709), .B(n6049), .X(\update_output_0/n1559 ) );
  nor_x1_sg U10387 ( .A(n6557), .B(n7105), .X(\update_output_0/n1539 ) );
  nor_x1_sg U10388 ( .A(n6689), .B(n6020), .X(\update_output_0/n2811 ) );
  nor_x1_sg U10389 ( .A(n6679), .B(n7105), .X(\update_output_0/n2807 ) );
  nor_x1_sg U10390 ( .A(n6600), .B(n6432), .X(\update_output_0/n2795 ) );
  nor_x1_sg U10391 ( .A(n6585), .B(n6019), .X(\update_output_0/n2791 ) );
  nor_x1_sg U10392 ( .A(n6686), .B(n6020), .X(\update_output_0/n2787 ) );
  nor_x1_sg U10393 ( .A(n6590), .B(n6431), .X(\update_output_0/n2779 ) );
  nor_x1_sg U10394 ( .A(n6667), .B(n7105), .X(\update_output_0/n2771 ) );
  nor_x1_sg U10395 ( .A(n6605), .B(n7104), .X(\update_output_0/n2767 ) );
  nor_x1_sg U10396 ( .A(n6677), .B(n7103), .X(\update_output_0/n2755 ) );
  nor_x1_sg U10397 ( .A(n6672), .B(n7106), .X(\update_output_0/n2751 ) );
  nor_x1_sg U10398 ( .A(n6595), .B(n6432), .X(\update_output_0/n2747 ) );
  nor_x1_sg U10399 ( .A(n6555), .B(n6414), .X(\update_output_0/n2743 ) );
  nor_x1_sg U10400 ( .A(n6688), .B(n6413), .X(\update_output_0/n2731 ) );
  nor_x1_sg U10401 ( .A(n6682), .B(n6414), .X(\update_output_0/n2727 ) );
  nor_x1_sg U10402 ( .A(n6599), .B(n6046), .X(\update_output_0/n2715 ) );
  nor_x1_sg U10403 ( .A(n6586), .B(n6046), .X(\update_output_0/n2711 ) );
  nor_x1_sg U10404 ( .A(n6684), .B(n7181), .X(\update_output_0/n2707 ) );
  nor_x1_sg U10405 ( .A(n6589), .B(n6413), .X(\update_output_0/n2699 ) );
  nor_x1_sg U10406 ( .A(n6665), .B(n6413), .X(\update_output_0/n2691 ) );
  nor_x1_sg U10407 ( .A(n6606), .B(n7182), .X(\update_output_0/n2687 ) );
  nor_x1_sg U10408 ( .A(n6675), .B(n6046), .X(\update_output_0/n2675 ) );
  nor_x1_sg U10409 ( .A(n6670), .B(n6206), .X(\update_output_0/n2671 ) );
  nor_x1_sg U10410 ( .A(n6595), .B(n7180), .X(\update_output_0/n2667 ) );
  nor_x1_sg U10411 ( .A(n6557), .B(n6070), .X(\update_output_0/n2663 ) );
  nor_x1_sg U10412 ( .A(n6689), .B(n6397), .X(\update_output_0/n2651 ) );
  nor_x1_sg U10413 ( .A(n6680), .B(n7220), .X(\update_output_0/n2647 ) );
  nor_x1_sg U10414 ( .A(n6600), .B(n6071), .X(\update_output_0/n2635 ) );
  nor_x1_sg U10415 ( .A(n6583), .B(n7219), .X(\update_output_0/n2631 ) );
  nor_x1_sg U10416 ( .A(n6685), .B(n6231), .X(\update_output_0/n2627 ) );
  nor_x1_sg U10417 ( .A(n6590), .B(n7221), .X(\update_output_0/n2619 ) );
  nor_x1_sg U10418 ( .A(n6666), .B(n6230), .X(\update_output_0/n2611 ) );
  nor_x1_sg U10419 ( .A(n6606), .B(n6230), .X(\update_output_0/n2607 ) );
  nor_x1_sg U10420 ( .A(n6676), .B(n6071), .X(\update_output_0/n2595 ) );
  nor_x1_sg U10421 ( .A(n6671), .B(n7221), .X(\update_output_0/n2591 ) );
  nor_x1_sg U10422 ( .A(n6596), .B(n6071), .X(\update_output_0/n2587 ) );
  nor_x1_sg U10423 ( .A(n6556), .B(n7176), .X(\update_output_0/n2583 ) );
  nor_x1_sg U10424 ( .A(n6689), .B(n7174), .X(\update_output_0/n2571 ) );
  nor_x1_sg U10425 ( .A(n6679), .B(n7174), .X(\update_output_0/n2567 ) );
  nor_x1_sg U10426 ( .A(n6598), .B(n6416), .X(\update_output_0/n2555 ) );
  nor_x1_sg U10427 ( .A(n6586), .B(n6203), .X(\update_output_0/n2551 ) );
  nor_x1_sg U10428 ( .A(n6685), .B(n7174), .X(\update_output_0/n2547 ) );
  nor_x1_sg U10429 ( .A(n6591), .B(n6203), .X(\update_output_0/n2539 ) );
  nor_x1_sg U10430 ( .A(n6664), .B(n6416), .X(\update_output_0/n2531 ) );
  nor_x1_sg U10431 ( .A(n6605), .B(n6043), .X(\update_output_0/n2527 ) );
  nor_x1_sg U10432 ( .A(n6674), .B(n6416), .X(\update_output_0/n2515 ) );
  nor_x1_sg U10433 ( .A(n6669), .B(n6415), .X(\update_output_0/n2511 ) );
  nor_x1_sg U10434 ( .A(n6596), .B(n6043), .X(\update_output_0/n2507 ) );
  nor_x1_sg U10435 ( .A(n6557), .B(n7119), .X(\update_output_0/n2503 ) );
  nor_x1_sg U10436 ( .A(n6688), .B(n6028), .X(\update_output_0/n2491 ) );
  nor_x1_sg U10437 ( .A(n6680), .B(n6426), .X(\update_output_0/n2487 ) );
  nor_x1_sg U10438 ( .A(n6601), .B(n6029), .X(\update_output_0/n2475 ) );
  nor_x1_sg U10439 ( .A(n6584), .B(n6191), .X(\update_output_0/n2471 ) );
  nor_x1_sg U10440 ( .A(n6686), .B(n6191), .X(\update_output_0/n2467 ) );
  nor_x1_sg U10441 ( .A(n6589), .B(n7121), .X(\update_output_0/n2459 ) );
  nor_x1_sg U10442 ( .A(n6666), .B(n6425), .X(\update_output_0/n2451 ) );
  nor_x1_sg U10443 ( .A(n6603), .B(n7121), .X(\update_output_0/n2447 ) );
  nor_x1_sg U10444 ( .A(n6676), .B(n6029), .X(\update_output_0/n2435 ) );
  nor_x1_sg U10445 ( .A(n6671), .B(n6191), .X(\update_output_0/n2431 ) );
  nor_x1_sg U10446 ( .A(n6593), .B(n7121), .X(\update_output_0/n2427 ) );
  nor_x1_sg U10447 ( .A(n6555), .B(n7209), .X(\update_output_0/n2423 ) );
  nor_x1_sg U10448 ( .A(n6690), .B(n6225), .X(\update_output_0/n2411 ) );
  nor_x1_sg U10449 ( .A(n6682), .B(n7209), .X(\update_output_0/n2407 ) );
  nor_x1_sg U10450 ( .A(n6599), .B(n7212), .X(\update_output_0/n2395 ) );
  nor_x1_sg U10451 ( .A(n6585), .B(n7211), .X(\update_output_0/n2391 ) );
  nor_x1_sg U10452 ( .A(n5962), .B(n7212), .X(\update_output_0/n2387 ) );
  nor_x1_sg U10453 ( .A(n6588), .B(n6401), .X(\update_output_0/n2379 ) );
  nor_x1_sg U10454 ( .A(n6664), .B(n6065), .X(\update_output_0/n2371 ) );
  nor_x1_sg U10455 ( .A(n6603), .B(n6224), .X(\update_output_0/n2367 ) );
  nor_x1_sg U10456 ( .A(n6674), .B(n6402), .X(\update_output_0/n2355 ) );
  nor_x1_sg U10457 ( .A(n6669), .B(n7210), .X(\update_output_0/n2351 ) );
  nor_x1_sg U10458 ( .A(n6595), .B(n6225), .X(\update_output_0/n2347 ) );
  nor_x1_sg U10459 ( .A(n6556), .B(n6222), .X(\update_output_0/n2343 ) );
  nor_x1_sg U10460 ( .A(n6688), .B(n6061), .X(\update_output_0/n2331 ) );
  nor_x1_sg U10461 ( .A(n6681), .B(n6221), .X(\update_output_0/n2327 ) );
  nor_x1_sg U10462 ( .A(n6601), .B(n7204), .X(\update_output_0/n2315 ) );
  nor_x1_sg U10463 ( .A(n6585), .B(n7207), .X(\update_output_0/n2311 ) );
  nor_x1_sg U10464 ( .A(n6684), .B(n7206), .X(\update_output_0/n2307 ) );
  nor_x1_sg U10465 ( .A(n6591), .B(n7204), .X(\update_output_0/n2299 ) );
  nor_x1_sg U10466 ( .A(n6665), .B(n7204), .X(\update_output_0/n2291 ) );
  nor_x1_sg U10467 ( .A(n6603), .B(n6062), .X(\update_output_0/n2287 ) );
  nor_x1_sg U10468 ( .A(n6675), .B(n6403), .X(\update_output_0/n2275 ) );
  nor_x1_sg U10469 ( .A(n6670), .B(n7207), .X(\update_output_0/n2271 ) );
  nor_x1_sg U10470 ( .A(n6593), .B(n7205), .X(\update_output_0/n2267 ) );
  nor_x1_sg U10471 ( .A(n6555), .B(n6406), .X(\update_output_0/n2263 ) );
  nor_x1_sg U10472 ( .A(n6691), .B(n6405), .X(\update_output_0/n2251 ) );
  nor_x1_sg U10473 ( .A(n6681), .B(n6406), .X(\update_output_0/n2247 ) );
  nor_x1_sg U10474 ( .A(n6601), .B(n6058), .X(\update_output_0/n2235 ) );
  nor_x1_sg U10475 ( .A(n6584), .B(n6058), .X(\update_output_0/n2231 ) );
  nor_x1_sg U10476 ( .A(n5962), .B(n7201), .X(\update_output_0/n2227 ) );
  nor_x1_sg U10477 ( .A(n6590), .B(n6405), .X(\update_output_0/n2219 ) );
  nor_x1_sg U10478 ( .A(n6664), .B(n6405), .X(\update_output_0/n2211 ) );
  nor_x1_sg U10479 ( .A(n6605), .B(n7202), .X(\update_output_0/n2207 ) );
  nor_x1_sg U10480 ( .A(n6674), .B(n6058), .X(\update_output_0/n2195 ) );
  nor_x1_sg U10481 ( .A(n6669), .B(n6218), .X(\update_output_0/n2191 ) );
  nor_x1_sg U10482 ( .A(n6593), .B(n7200), .X(\update_output_0/n2187 ) );
  nor_x1_sg U10483 ( .A(n6554), .B(n6025), .X(\update_output_0/n2183 ) );
  nor_x1_sg U10484 ( .A(n6691), .B(n7113), .X(\update_output_0/n2171 ) );
  nor_x1_sg U10485 ( .A(n6682), .B(n7116), .X(\update_output_0/n2167 ) );
  nor_x1_sg U10486 ( .A(n6599), .B(n7114), .X(\update_output_0/n2155 ) );
  nor_x1_sg U10487 ( .A(n6584), .B(n6026), .X(\update_output_0/n2151 ) );
  nor_x1_sg U10488 ( .A(n6684), .B(n7116), .X(\update_output_0/n2147 ) );
  nor_x1_sg U10489 ( .A(n6588), .B(n6025), .X(\update_output_0/n2139 ) );
  nor_x1_sg U10490 ( .A(n6667), .B(n6026), .X(\update_output_0/n2131 ) );
  nor_x1_sg U10491 ( .A(n6604), .B(n6427), .X(\update_output_0/n2127 ) );
  nor_x1_sg U10492 ( .A(n6677), .B(n6189), .X(\update_output_0/n2115 ) );
  nor_x1_sg U10493 ( .A(n6672), .B(n6428), .X(\update_output_0/n2111 ) );
  nor_x1_sg U10494 ( .A(n6594), .B(n7116), .X(\update_output_0/n2107 ) );
  nor_x1_sg U10495 ( .A(n6554), .B(n6201), .X(\update_output_0/n2103 ) );
  nor_x1_sg U10496 ( .A(n6690), .B(n6040), .X(\update_output_0/n2091 ) );
  nor_x1_sg U10497 ( .A(n6680), .B(n6200), .X(\update_output_0/n2087 ) );
  nor_x1_sg U10498 ( .A(n6600), .B(n7169), .X(\update_output_0/n2075 ) );
  nor_x1_sg U10499 ( .A(n6583), .B(n7172), .X(\update_output_0/n2071 ) );
  nor_x1_sg U10500 ( .A(n7420), .B(n7171), .X(\update_output_0/n2067 ) );
  nor_x1_sg U10501 ( .A(n6591), .B(n7169), .X(\update_output_0/n2059 ) );
  nor_x1_sg U10502 ( .A(n6665), .B(n7169), .X(\update_output_0/n2051 ) );
  nor_x1_sg U10503 ( .A(n6606), .B(n6041), .X(\update_output_0/n2047 ) );
  nor_x1_sg U10504 ( .A(n6675), .B(n7172), .X(\update_output_0/n2035 ) );
  nor_x1_sg U10505 ( .A(n6670), .B(n6417), .X(\update_output_0/n2031 ) );
  nor_x1_sg U10506 ( .A(n6596), .B(n7170), .X(\update_output_0/n2027 ) );
  nor_x1_sg U10507 ( .A(n6554), .B(n6227), .X(\update_output_0/n2023 ) );
  nor_x1_sg U10508 ( .A(n6690), .B(n7216), .X(\update_output_0/n2011 ) );
  nor_x1_sg U10509 ( .A(n6679), .B(n7215), .X(\update_output_0/n2007 ) );
  nor_x1_sg U10510 ( .A(n6598), .B(n6227), .X(\update_output_0/n1995 ) );
  nor_x1_sg U10511 ( .A(n6586), .B(n7216), .X(\update_output_0/n1991 ) );
  nor_x1_sg U10512 ( .A(n6684), .B(n6400), .X(\update_output_0/n1987 ) );
  nor_x1_sg U10513 ( .A(n6588), .B(n7217), .X(\update_output_0/n1979 ) );
  nor_x1_sg U10514 ( .A(n6665), .B(n7214), .X(\update_output_0/n1971 ) );
  nor_x1_sg U10515 ( .A(n6605), .B(n7216), .X(\update_output_0/n1967 ) );
  nor_x1_sg U10516 ( .A(n6675), .B(n6068), .X(\update_output_0/n1955 ) );
  nor_x1_sg U10517 ( .A(n6670), .B(n6400), .X(\update_output_0/n1951 ) );
  nor_x1_sg U10518 ( .A(n6594), .B(n7217), .X(\update_output_0/n1947 ) );
  nor_x1_sg U10519 ( .A(n6557), .B(n6419), .X(\update_output_0/n1943 ) );
  nor_x1_sg U10520 ( .A(n6688), .B(n7167), .X(\update_output_0/n1931 ) );
  nor_x1_sg U10521 ( .A(n6682), .B(n7165), .X(\update_output_0/n1927 ) );
  nor_x1_sg U10522 ( .A(n6601), .B(n7166), .X(\update_output_0/n1915 ) );
  nor_x1_sg U10523 ( .A(n6583), .B(n7164), .X(\update_output_0/n1911 ) );
  nor_x1_sg U10524 ( .A(n6686), .B(n7166), .X(\update_output_0/n1907 ) );
  nor_x1_sg U10525 ( .A(n6590), .B(n6037), .X(\update_output_0/n1899 ) );
  nor_x1_sg U10526 ( .A(n6664), .B(n6038), .X(\update_output_0/n1891 ) );
  nor_x1_sg U10527 ( .A(n6604), .B(n7165), .X(\update_output_0/n1887 ) );
  nor_x1_sg U10528 ( .A(n6674), .B(n7166), .X(\update_output_0/n1875 ) );
  nor_x1_sg U10529 ( .A(n6669), .B(n6198), .X(\update_output_0/n1871 ) );
  nor_x1_sg U10530 ( .A(n6594), .B(n7164), .X(\update_output_0/n1867 ) );
  nor_x1_sg U10531 ( .A(n6556), .B(n6186), .X(\update_output_0/n1863 ) );
  nor_x1_sg U10532 ( .A(n6689), .B(n6022), .X(\update_output_0/n1851 ) );
  nor_x1_sg U10533 ( .A(n6681), .B(n6185), .X(\update_output_0/n1847 ) );
  nor_x1_sg U10534 ( .A(n6600), .B(n7108), .X(\update_output_0/n1835 ) );
  nor_x1_sg U10535 ( .A(n6585), .B(n7111), .X(\update_output_0/n1831 ) );
  nor_x1_sg U10536 ( .A(n6685), .B(n7110), .X(\update_output_0/n1827 ) );
  nor_x1_sg U10537 ( .A(n6589), .B(n7108), .X(\update_output_0/n1819 ) );
  nor_x1_sg U10538 ( .A(n6667), .B(n7108), .X(\update_output_0/n1811 ) );
  nor_x1_sg U10539 ( .A(n6604), .B(n6023), .X(\update_output_0/n1807 ) );
  nor_x1_sg U10540 ( .A(n6677), .B(n6429), .X(\update_output_0/n1795 ) );
  nor_x1_sg U10541 ( .A(n6672), .B(n7111), .X(\update_output_0/n1791 ) );
  nor_x1_sg U10542 ( .A(n6593), .B(n7109), .X(\update_output_0/n1787 ) );
  nor_x1_sg U10543 ( .A(n6556), .B(n6215), .X(\update_output_0/n1783 ) );
  nor_x1_sg U10544 ( .A(n6690), .B(n7197), .X(\update_output_0/n1771 ) );
  nor_x1_sg U10545 ( .A(n6680), .B(n7194), .X(\update_output_0/n1767 ) );
  nor_x1_sg U10546 ( .A(n6599), .B(n7196), .X(\update_output_0/n1755 ) );
  nor_x1_sg U10547 ( .A(n6586), .B(n7197), .X(\update_output_0/n1751 ) );
  nor_x1_sg U10548 ( .A(n7420), .B(n6408), .X(\update_output_0/n1747 ) );
  nor_x1_sg U10549 ( .A(n6591), .B(n7194), .X(\update_output_0/n1739 ) );
  nor_x1_sg U10550 ( .A(n6666), .B(n6408), .X(\update_output_0/n1731 ) );
  nor_x1_sg U10551 ( .A(n6604), .B(n6056), .X(\update_output_0/n1727 ) );
  nor_x1_sg U10552 ( .A(n6676), .B(n6055), .X(\update_output_0/n1715 ) );
  nor_x1_sg U10553 ( .A(n6671), .B(n6407), .X(\update_output_0/n1711 ) );
  nor_x1_sg U10554 ( .A(n6596), .B(n6055), .X(\update_output_0/n1707 ) );
  nor_x1_sg U10555 ( .A(n6555), .B(n7191), .X(\update_output_0/n1703 ) );
  nor_x1_sg U10556 ( .A(n6691), .B(n7190), .X(\update_output_0/n1691 ) );
  nor_x1_sg U10557 ( .A(n6679), .B(n6212), .X(\update_output_0/n1687 ) );
  nor_x1_sg U10558 ( .A(n6598), .B(n6053), .X(\update_output_0/n1675 ) );
  nor_x1_sg U10559 ( .A(n6584), .B(n6409), .X(\update_output_0/n1671 ) );
  nor_x1_sg U10560 ( .A(n6685), .B(n6213), .X(\update_output_0/n1667 ) );
  nor_x1_sg U10561 ( .A(n6588), .B(n7189), .X(\update_output_0/n1659 ) );
  nor_x1_sg U10562 ( .A(n6667), .B(n6052), .X(\update_output_0/n1651 ) );
  nor_x1_sg U10563 ( .A(n6603), .B(n7192), .X(\update_output_0/n1647 ) );
  nor_x1_sg U10564 ( .A(n6677), .B(n7189), .X(\update_output_0/n1635 ) );
  nor_x1_sg U10565 ( .A(n6672), .B(n6213), .X(\update_output_0/n1631 ) );
  nor_x1_sg U10566 ( .A(n6595), .B(n6213), .X(\update_output_0/n1627 ) );
  nor_x1_sg U10567 ( .A(n6554), .B(n7184), .X(\update_output_0/n1623 ) );
  nor_x1_sg U10568 ( .A(n6691), .B(n6411), .X(\update_output_0/n1611 ) );
  nor_x1_sg U10569 ( .A(n6681), .B(n6411), .X(\update_output_0/n1607 ) );
  nor_x1_sg U10570 ( .A(n6598), .B(n6210), .X(\update_output_0/n1595 ) );
  nor_x1_sg U10571 ( .A(n6583), .B(n6209), .X(\update_output_0/n1591 ) );
  nor_x1_sg U10572 ( .A(n6686), .B(n7187), .X(\update_output_0/n1587 ) );
  nor_x1_sg U10573 ( .A(n6589), .B(n6050), .X(\update_output_0/n1579 ) );
  nor_x1_sg U10574 ( .A(n6666), .B(n6049), .X(\update_output_0/n1571 ) );
  nor_x1_sg U10575 ( .A(n6606), .B(n6209), .X(\update_output_0/n1567 ) );
  nor_x1_sg U10576 ( .A(n6676), .B(n7185), .X(\update_output_0/n1555 ) );
  nor_x1_sg U10577 ( .A(n6671), .B(n7187), .X(\update_output_0/n1551 ) );
  nor_x1_sg U10578 ( .A(n6594), .B(n6412), .X(\update_output_0/n1547 ) );
  nor_x1_sg U10579 ( .A(n6158), .B(n7398), .X(n3782) );
  nor_x1_sg U10580 ( .A(n743), .B(n6779), .X(n1247) );
  nor_x1_sg U10581 ( .A(n6814), .B(n1249), .X(n1248) );
  nand_x1_sg U10582 ( .A(n5912), .B(n5914), .X(n1249) );
  nor_x1_sg U10583 ( .A(n6769), .B(n6794), .X(n951) );
  nor_x1_sg U10584 ( .A(n6774), .B(n953), .X(n952) );
  nand_x1_sg U10585 ( .A(n5937), .B(n5934), .X(n953) );
  nor_x1_sg U10586 ( .A(n6804), .B(n784), .X(n783) );
  nand_x1_sg U10587 ( .A(n5930), .B(n5932), .X(n784) );
  nor_x1_sg U10588 ( .A(n6824), .B(n6789), .X(n1116) );
  nor_x1_sg U10589 ( .A(n6809), .B(n1118), .X(n1117) );
  nand_x1_sg U10590 ( .A(n5939), .B(n5928), .X(n1118) );
  nand_x1_sg U10591 ( .A(n3523), .B(n6315), .X(n3522) );
  nand_x1_sg U10592 ( .A(n3826), .B(n3524), .X(n3825) );
  nand_x1_sg U10593 ( .A(n3739), .B(n6315), .X(n3738) );
  nor_x1_sg U10594 ( .A(n6784), .B(n6799), .X(n782) );
  nand_x1_sg U10595 ( .A(n3739), .B(n6320), .X(n4082) );
  nand_x1_sg U10596 ( .A(n3523), .B(n6320), .X(n3868) );
  nand_x1_sg U10597 ( .A(n6829), .B(n3911), .X(n7470) );
  nand_x1_sg U10598 ( .A(n5967), .B(n4039), .X(n7467) );
  nor_x1_sg U10599 ( .A(n7404), .B(n3997), .X(n3653) );
  nand_x1_sg U10600 ( .A(n6093), .B(n7001), .X(n3471) );
  nor_x1_sg U10601 ( .A(n6263), .B(n7439), .X(n3462) );
  nor_x1_sg U10602 ( .A(n6080), .B(n9225), .X(n3461) );
  inv_x1_sg U10603 ( .A(n3462), .X(n9225) );
  nor_x1_sg U10604 ( .A(n7414), .B(n3869), .X(n3610) );
  nand_x1_sg U10605 ( .A(n9238), .B(n7003), .X(n3869) );
  inv_x1_sg U10606 ( .A(n3954), .X(n9238) );
  nor_x1_sg U10607 ( .A(n3471), .B(n7439), .X(n3470) );
  nor_x1_sg U10608 ( .A(n3472), .B(n3473), .X(n3469) );
  nor_x1_sg U10609 ( .A(n6263), .B(n3474), .X(n3472) );
  nand_x1_sg U10610 ( .A(n6832), .B(n7404), .X(n4861) );
  inv_x1_sg U10611 ( .A(n5617), .X(n9228) );
  nand_x1_sg U10612 ( .A(n6460), .B(n6478), .X(n5614) );
  nor_x1_sg U10613 ( .A(n771), .B(n7398), .X(n756) );
  nor_x1_sg U10614 ( .A(n771), .B(n4821), .X(n767) );
  nand_x1_sg U10615 ( .A(n1465), .B(n1469), .X(n1468) );
  inv_x1_sg U10616 ( .A(n3474), .X(n8894) );
  nand_x1_sg U10617 ( .A(n760), .B(n7391), .X(n762) );
  nand_x1_sg U10618 ( .A(n760), .B(n8894), .X(n763) );
  nand_x1_sg U10619 ( .A(n760), .B(n7397), .X(n764) );
  nand_x1_sg U10620 ( .A(n773), .B(n7391), .X(n774) );
  nand_x1_sg U10621 ( .A(n773), .B(n8894), .X(n775) );
  nand_x1_sg U10622 ( .A(n773), .B(n7397), .X(n776) );
  nand_x1_sg U10623 ( .A(n756), .B(n7391), .X(n754) );
  nand_x1_sg U10624 ( .A(n756), .B(n6157), .X(n758) );
  nand_x1_sg U10625 ( .A(n767), .B(n7391), .X(n768) );
  nand_x1_sg U10626 ( .A(n767), .B(n6157), .X(n770) );
  nor_x1_sg U10627 ( .A(n6790), .B(n7103), .X(\update_output_0/n1538 ) );
  nor_x1_sg U10628 ( .A(n6827), .B(n6432), .X(\update_output_0/n2810 ) );
  nor_x1_sg U10629 ( .A(n6811), .B(n6431), .X(\update_output_0/n2806 ) );
  nor_x1_sg U10630 ( .A(n6815), .B(n6183), .X(\update_output_0/n2794 ) );
  nor_x1_sg U10631 ( .A(n6782), .B(n6020), .X(\update_output_0/n2790 ) );
  nor_x1_sg U10632 ( .A(n6820), .B(n7103), .X(\update_output_0/n2786 ) );
  nor_x1_sg U10633 ( .A(n6777), .B(n7106), .X(\update_output_0/n2778 ) );
  nor_x1_sg U10634 ( .A(n6797), .B(n6183), .X(\update_output_0/n2770 ) );
  nor_x1_sg U10635 ( .A(n6771), .B(n6019), .X(\update_output_0/n2766 ) );
  nor_x1_sg U10636 ( .A(n6807), .B(n6182), .X(\update_output_0/n2754 ) );
  nor_x1_sg U10637 ( .A(n6802), .B(n6431), .X(\update_output_0/n2750 ) );
  nor_x1_sg U10638 ( .A(n5949), .B(n7106), .X(\update_output_0/n2746 ) );
  nor_x1_sg U10639 ( .A(n6792), .B(n7182), .X(\update_output_0/n2742 ) );
  nor_x1_sg U10640 ( .A(n6826), .B(n6207), .X(\update_output_0/n2730 ) );
  nor_x1_sg U10641 ( .A(n6812), .B(n6414), .X(\update_output_0/n2726 ) );
  nor_x1_sg U10642 ( .A(n6815), .B(n7179), .X(\update_output_0/n2714 ) );
  nor_x1_sg U10643 ( .A(n6782), .B(n6206), .X(\update_output_0/n2710 ) );
  nor_x1_sg U10644 ( .A(n6822), .B(n6047), .X(\update_output_0/n2706 ) );
  nor_x1_sg U10645 ( .A(n6774), .B(n6413), .X(\update_output_0/n2698 ) );
  nor_x1_sg U10646 ( .A(n6796), .B(n6207), .X(\update_output_0/n2690 ) );
  nor_x1_sg U10647 ( .A(n6769), .B(n7181), .X(\update_output_0/n2686 ) );
  nor_x1_sg U10648 ( .A(n6806), .B(n6047), .X(\update_output_0/n2674 ) );
  nor_x1_sg U10649 ( .A(n6801), .B(n7181), .X(\update_output_0/n2670 ) );
  nor_x1_sg U10650 ( .A(n6785), .B(n6207), .X(\update_output_0/n2666 ) );
  nor_x1_sg U10651 ( .A(n6792), .B(n7221), .X(\update_output_0/n2662 ) );
  nor_x1_sg U10652 ( .A(n5965), .B(n6398), .X(\update_output_0/n2650 ) );
  nor_x1_sg U10653 ( .A(n6810), .B(n6231), .X(\update_output_0/n2646 ) );
  nor_x1_sg U10654 ( .A(n6815), .B(n6230), .X(\update_output_0/n2634 ) );
  nor_x1_sg U10655 ( .A(n5947), .B(n6231), .X(\update_output_0/n2630 ) );
  nor_x1_sg U10656 ( .A(n6822), .B(n7220), .X(\update_output_0/n2626 ) );
  nor_x1_sg U10657 ( .A(n6776), .B(n6398), .X(\update_output_0/n2618 ) );
  nor_x1_sg U10658 ( .A(n5953), .B(n7220), .X(\update_output_0/n2610 ) );
  nor_x1_sg U10659 ( .A(n6772), .B(n7222), .X(\update_output_0/n2606 ) );
  nor_x1_sg U10660 ( .A(n5957), .B(n7222), .X(\update_output_0/n2594 ) );
  nor_x1_sg U10661 ( .A(n5955), .B(n7219), .X(\update_output_0/n2590 ) );
  nor_x1_sg U10662 ( .A(n6787), .B(n7222), .X(\update_output_0/n2586 ) );
  nor_x1_sg U10663 ( .A(n6789), .B(n6044), .X(\update_output_0/n2582 ) );
  nor_x1_sg U10664 ( .A(n6825), .B(n7176), .X(\update_output_0/n2570 ) );
  nor_x1_sg U10665 ( .A(n6811), .B(n7175), .X(\update_output_0/n2566 ) );
  nor_x1_sg U10666 ( .A(n6815), .B(n6415), .X(\update_output_0/n2554 ) );
  nor_x1_sg U10667 ( .A(n6780), .B(n6203), .X(\update_output_0/n2550 ) );
  nor_x1_sg U10668 ( .A(n6819), .B(n7176), .X(\update_output_0/n2546 ) );
  nor_x1_sg U10669 ( .A(n6777), .B(n7175), .X(\update_output_0/n2538 ) );
  nor_x1_sg U10670 ( .A(n6795), .B(n6044), .X(\update_output_0/n2530 ) );
  nor_x1_sg U10671 ( .A(n6770), .B(n6416), .X(\update_output_0/n2526 ) );
  nor_x1_sg U10672 ( .A(n6805), .B(n7177), .X(\update_output_0/n2514 ) );
  nor_x1_sg U10673 ( .A(n6800), .B(n6203), .X(\update_output_0/n2510 ) );
  nor_x1_sg U10674 ( .A(n5949), .B(n7174), .X(\update_output_0/n2506 ) );
  nor_x1_sg U10675 ( .A(n5951), .B(n7120), .X(\update_output_0/n2502 ) );
  nor_x1_sg U10676 ( .A(n6826), .B(n6425), .X(\update_output_0/n2490 ) );
  nor_x1_sg U10677 ( .A(n6810), .B(n6426), .X(\update_output_0/n2486 ) );
  nor_x1_sg U10678 ( .A(n5961), .B(n6192), .X(\update_output_0/n2474 ) );
  nor_x1_sg U10679 ( .A(n6780), .B(n6028), .X(\update_output_0/n2470 ) );
  nor_x1_sg U10680 ( .A(n6821), .B(n6029), .X(\update_output_0/n2466 ) );
  nor_x1_sg U10681 ( .A(n5945), .B(n6028), .X(\update_output_0/n2458 ) );
  nor_x1_sg U10682 ( .A(n5953), .B(n7120), .X(\update_output_0/n2450 ) );
  nor_x1_sg U10683 ( .A(n6769), .B(n7119), .X(\update_output_0/n2446 ) );
  nor_x1_sg U10684 ( .A(n5957), .B(n6426), .X(\update_output_0/n2434 ) );
  nor_x1_sg U10685 ( .A(n5955), .B(n7118), .X(\update_output_0/n2430 ) );
  nor_x1_sg U10686 ( .A(n6785), .B(n7119), .X(\update_output_0/n2426 ) );
  nor_x1_sg U10687 ( .A(n6791), .B(n6401), .X(\update_output_0/n2422 ) );
  nor_x1_sg U10688 ( .A(n6824), .B(n7210), .X(\update_output_0/n2410 ) );
  nor_x1_sg U10689 ( .A(n6812), .B(n6065), .X(\update_output_0/n2406 ) );
  nor_x1_sg U10690 ( .A(n5961), .B(n6065), .X(\update_output_0/n2394 ) );
  nor_x1_sg U10691 ( .A(n6781), .B(n6224), .X(\update_output_0/n2390 ) );
  nor_x1_sg U10692 ( .A(n6821), .B(n7211), .X(\update_output_0/n2386 ) );
  nor_x1_sg U10693 ( .A(n6776), .B(n6064), .X(\update_output_0/n2378 ) );
  nor_x1_sg U10694 ( .A(n6794), .B(n7212), .X(\update_output_0/n2370 ) );
  nor_x1_sg U10695 ( .A(n6771), .B(n6225), .X(\update_output_0/n2366 ) );
  nor_x1_sg U10696 ( .A(n6804), .B(n7210), .X(\update_output_0/n2354 ) );
  nor_x1_sg U10697 ( .A(n6799), .B(n6402), .X(\update_output_0/n2350 ) );
  nor_x1_sg U10698 ( .A(n6786), .B(n7210), .X(\update_output_0/n2346 ) );
  nor_x1_sg U10699 ( .A(n6790), .B(n6062), .X(\update_output_0/n2342 ) );
  nor_x1_sg U10700 ( .A(n6825), .B(n7205), .X(\update_output_0/n2330 ) );
  nor_x1_sg U10701 ( .A(n5959), .B(n6221), .X(\update_output_0/n2326 ) );
  nor_x1_sg U10702 ( .A(n6814), .B(n6222), .X(\update_output_0/n2314 ) );
  nor_x1_sg U10703 ( .A(n6782), .B(n6403), .X(\update_output_0/n2310 ) );
  nor_x1_sg U10704 ( .A(n6820), .B(n7207), .X(\update_output_0/n2306 ) );
  nor_x1_sg U10705 ( .A(n6775), .B(n6221), .X(\update_output_0/n2298 ) );
  nor_x1_sg U10706 ( .A(n6796), .B(n6404), .X(\update_output_0/n2290 ) );
  nor_x1_sg U10707 ( .A(n6769), .B(n6403), .X(\update_output_0/n2286 ) );
  nor_x1_sg U10708 ( .A(n6806), .B(n7207), .X(\update_output_0/n2274 ) );
  nor_x1_sg U10709 ( .A(n6801), .B(n7205), .X(\update_output_0/n2270 ) );
  nor_x1_sg U10710 ( .A(n6787), .B(n6404), .X(\update_output_0/n2266 ) );
  nor_x1_sg U10711 ( .A(n6790), .B(n7202), .X(\update_output_0/n2262 ) );
  nor_x1_sg U10712 ( .A(n5965), .B(n6219), .X(\update_output_0/n2250 ) );
  nor_x1_sg U10713 ( .A(n6809), .B(n6406), .X(\update_output_0/n2246 ) );
  nor_x1_sg U10714 ( .A(n6817), .B(n7199), .X(\update_output_0/n2234 ) );
  nor_x1_sg U10715 ( .A(n6780), .B(n6218), .X(\update_output_0/n2230 ) );
  nor_x1_sg U10716 ( .A(n5963), .B(n6059), .X(\update_output_0/n2226 ) );
  nor_x1_sg U10717 ( .A(n6777), .B(n6405), .X(\update_output_0/n2218 ) );
  nor_x1_sg U10718 ( .A(n6794), .B(n6219), .X(\update_output_0/n2210 ) );
  nor_x1_sg U10719 ( .A(n5943), .B(n7201), .X(\update_output_0/n2206 ) );
  nor_x1_sg U10720 ( .A(n6804), .B(n6059), .X(\update_output_0/n2194 ) );
  nor_x1_sg U10721 ( .A(n6799), .B(n7201), .X(\update_output_0/n2190 ) );
  nor_x1_sg U10722 ( .A(n6785), .B(n6219), .X(\update_output_0/n2186 ) );
  nor_x1_sg U10723 ( .A(n6790), .B(n6189), .X(\update_output_0/n2182 ) );
  nor_x1_sg U10724 ( .A(n6824), .B(n6026), .X(\update_output_0/n2170 ) );
  nor_x1_sg U10725 ( .A(n6809), .B(n7115), .X(\update_output_0/n2166 ) );
  nor_x1_sg U10726 ( .A(n6817), .B(n7113), .X(\update_output_0/n2154 ) );
  nor_x1_sg U10727 ( .A(n6779), .B(n6427), .X(\update_output_0/n2150 ) );
  nor_x1_sg U10728 ( .A(n6821), .B(n6025), .X(\update_output_0/n2146 ) );
  nor_x1_sg U10729 ( .A(n6774), .B(n7114), .X(\update_output_0/n2138 ) );
  nor_x1_sg U10730 ( .A(n6794), .B(n7115), .X(\update_output_0/n2130 ) );
  nor_x1_sg U10731 ( .A(n6771), .B(n6427), .X(\update_output_0/n2126 ) );
  nor_x1_sg U10732 ( .A(n6804), .B(n6026), .X(\update_output_0/n2114 ) );
  nor_x1_sg U10733 ( .A(n6799), .B(n7113), .X(\update_output_0/n2110 ) );
  nor_x1_sg U10734 ( .A(n6784), .B(n6189), .X(\update_output_0/n2106 ) );
  nor_x1_sg U10735 ( .A(n6792), .B(n6041), .X(\update_output_0/n2102 ) );
  nor_x1_sg U10736 ( .A(n6825), .B(n7170), .X(\update_output_0/n2090 ) );
  nor_x1_sg U10737 ( .A(n5959), .B(n6200), .X(\update_output_0/n2086 ) );
  nor_x1_sg U10738 ( .A(n6814), .B(n6201), .X(\update_output_0/n2074 ) );
  nor_x1_sg U10739 ( .A(n5947), .B(n6417), .X(\update_output_0/n2070 ) );
  nor_x1_sg U10740 ( .A(n6820), .B(n7172), .X(\update_output_0/n2066 ) );
  nor_x1_sg U10741 ( .A(n6775), .B(n6200), .X(\update_output_0/n2058 ) );
  nor_x1_sg U10742 ( .A(n6796), .B(n6418), .X(\update_output_0/n2050 ) );
  nor_x1_sg U10743 ( .A(n6770), .B(n6417), .X(\update_output_0/n2046 ) );
  nor_x1_sg U10744 ( .A(n6806), .B(n7170), .X(\update_output_0/n2034 ) );
  nor_x1_sg U10745 ( .A(n6801), .B(n6200), .X(\update_output_0/n2030 ) );
  nor_x1_sg U10746 ( .A(n6784), .B(n6418), .X(\update_output_0/n2026 ) );
  nor_x1_sg U10747 ( .A(n6791), .B(n6067), .X(\update_output_0/n2022 ) );
  nor_x1_sg U10748 ( .A(n6827), .B(n6228), .X(\update_output_0/n2010 ) );
  nor_x1_sg U10749 ( .A(n6809), .B(n7216), .X(\update_output_0/n2006 ) );
  nor_x1_sg U10750 ( .A(n6817), .B(n6227), .X(\update_output_0/n1994 ) );
  nor_x1_sg U10751 ( .A(n6779), .B(n6068), .X(\update_output_0/n1990 ) );
  nor_x1_sg U10752 ( .A(n6822), .B(n6399), .X(\update_output_0/n1986 ) );
  nor_x1_sg U10753 ( .A(n6776), .B(n7215), .X(\update_output_0/n1978 ) );
  nor_x1_sg U10754 ( .A(n6797), .B(n7214), .X(\update_output_0/n1970 ) );
  nor_x1_sg U10755 ( .A(n5943), .B(n7214), .X(\update_output_0/n1966 ) );
  nor_x1_sg U10756 ( .A(n6807), .B(n6067), .X(\update_output_0/n1954 ) );
  nor_x1_sg U10757 ( .A(n6802), .B(n7215), .X(\update_output_0/n1950 ) );
  nor_x1_sg U10758 ( .A(n5949), .B(n7217), .X(\update_output_0/n1946 ) );
  nor_x1_sg U10759 ( .A(n6791), .B(n6198), .X(\update_output_0/n1942 ) );
  nor_x1_sg U10760 ( .A(n6824), .B(n7165), .X(\update_output_0/n1930 ) );
  nor_x1_sg U10761 ( .A(n6812), .B(n7167), .X(\update_output_0/n1926 ) );
  nor_x1_sg U10762 ( .A(n6814), .B(n6198), .X(\update_output_0/n1914 ) );
  nor_x1_sg U10763 ( .A(n6781), .B(n7164), .X(\update_output_0/n1910 ) );
  nor_x1_sg U10764 ( .A(n6820), .B(n6420), .X(\update_output_0/n1906 ) );
  nor_x1_sg U10765 ( .A(n6775), .B(n6419), .X(\update_output_0/n1898 ) );
  nor_x1_sg U10766 ( .A(n6795), .B(n6419), .X(\update_output_0/n1890 ) );
  nor_x1_sg U10767 ( .A(n6770), .B(n7165), .X(\update_output_0/n1886 ) );
  nor_x1_sg U10768 ( .A(n6805), .B(n6197), .X(\update_output_0/n1874 ) );
  nor_x1_sg U10769 ( .A(n6800), .B(n6038), .X(\update_output_0/n1870 ) );
  nor_x1_sg U10770 ( .A(n6787), .B(n7167), .X(\update_output_0/n1866 ) );
  nor_x1_sg U10771 ( .A(n6789), .B(n6023), .X(\update_output_0/n1862 ) );
  nor_x1_sg U10772 ( .A(n6826), .B(n7109), .X(\update_output_0/n1850 ) );
  nor_x1_sg U10773 ( .A(n6810), .B(n6185), .X(\update_output_0/n1846 ) );
  nor_x1_sg U10774 ( .A(n6816), .B(n6186), .X(\update_output_0/n1834 ) );
  nor_x1_sg U10775 ( .A(n6780), .B(n6429), .X(\update_output_0/n1830 ) );
  nor_x1_sg U10776 ( .A(n6819), .B(n7111), .X(\update_output_0/n1826 ) );
  nor_x1_sg U10777 ( .A(n6774), .B(n6185), .X(\update_output_0/n1818 ) );
  nor_x1_sg U10778 ( .A(n6795), .B(n6430), .X(\update_output_0/n1810 ) );
  nor_x1_sg U10779 ( .A(n6772), .B(n6429), .X(\update_output_0/n1806 ) );
  nor_x1_sg U10780 ( .A(n6805), .B(n7111), .X(\update_output_0/n1794 ) );
  nor_x1_sg U10781 ( .A(n6800), .B(n7109), .X(\update_output_0/n1790 ) );
  nor_x1_sg U10782 ( .A(n6786), .B(n6430), .X(\update_output_0/n1786 ) );
  nor_x1_sg U10783 ( .A(n5951), .B(n6215), .X(\update_output_0/n1782 ) );
  nor_x1_sg U10784 ( .A(n5965), .B(n7195), .X(\update_output_0/n1770 ) );
  nor_x1_sg U10785 ( .A(n5959), .B(n7195), .X(\update_output_0/n1766 ) );
  nor_x1_sg U10786 ( .A(n5961), .B(n7194), .X(\update_output_0/n1754 ) );
  nor_x1_sg U10787 ( .A(n5947), .B(n6055), .X(\update_output_0/n1750 ) );
  nor_x1_sg U10788 ( .A(n6822), .B(n6216), .X(\update_output_0/n1746 ) );
  nor_x1_sg U10789 ( .A(n5945), .B(n7196), .X(\update_output_0/n1738 ) );
  nor_x1_sg U10790 ( .A(n5953), .B(n6407), .X(\update_output_0/n1730 ) );
  nor_x1_sg U10791 ( .A(n5943), .B(n6216), .X(\update_output_0/n1726 ) );
  nor_x1_sg U10792 ( .A(n5957), .B(n6407), .X(\update_output_0/n1714 ) );
  nor_x1_sg U10793 ( .A(n5955), .B(n7197), .X(\update_output_0/n1710 ) );
  nor_x1_sg U10794 ( .A(n6785), .B(n6408), .X(\update_output_0/n1706 ) );
  nor_x1_sg U10795 ( .A(n6789), .B(n6053), .X(\update_output_0/n1702 ) );
  nor_x1_sg U10796 ( .A(n6827), .B(n6053), .X(\update_output_0/n1690 ) );
  nor_x1_sg U10797 ( .A(n6810), .B(n6410), .X(\update_output_0/n1686 ) );
  nor_x1_sg U10798 ( .A(n6816), .B(n6212), .X(\update_output_0/n1674 ) );
  nor_x1_sg U10799 ( .A(n6781), .B(n6410), .X(\update_output_0/n1670 ) );
  nor_x1_sg U10800 ( .A(n6821), .B(n7191), .X(\update_output_0/n1666 ) );
  nor_x1_sg U10801 ( .A(n5945), .B(n7192), .X(\update_output_0/n1658 ) );
  nor_x1_sg U10802 ( .A(n6797), .B(n7189), .X(\update_output_0/n1650 ) );
  nor_x1_sg U10803 ( .A(n6772), .B(n6052), .X(\update_output_0/n1646 ) );
  nor_x1_sg U10804 ( .A(n6807), .B(n7192), .X(\update_output_0/n1634 ) );
  nor_x1_sg U10805 ( .A(n6802), .B(n6409), .X(\update_output_0/n1630 ) );
  nor_x1_sg U10806 ( .A(n6786), .B(n7192), .X(\update_output_0/n1626 ) );
  nor_x1_sg U10807 ( .A(n5951), .B(n7184), .X(\update_output_0/n1622 ) );
  nor_x1_sg U10808 ( .A(n6825), .B(n6412), .X(\update_output_0/n1610 ) );
  nor_x1_sg U10809 ( .A(n6811), .B(n6210), .X(\update_output_0/n1606 ) );
  nor_x1_sg U10810 ( .A(n6816), .B(n7187), .X(\update_output_0/n1594 ) );
  nor_x1_sg U10811 ( .A(n6779), .B(n6209), .X(\update_output_0/n1590 ) );
  nor_x1_sg U10812 ( .A(n5963), .B(n7185), .X(\update_output_0/n1586 ) );
  nor_x1_sg U10813 ( .A(n6775), .B(n7186), .X(\update_output_0/n1578 ) );
  nor_x1_sg U10814 ( .A(n6795), .B(n6050), .X(\update_output_0/n1570 ) );
  nor_x1_sg U10815 ( .A(n6770), .B(n6412), .X(\update_output_0/n1566 ) );
  nor_x1_sg U10816 ( .A(n6805), .B(n6411), .X(\update_output_0/n1554 ) );
  nor_x1_sg U10817 ( .A(n6800), .B(n6049), .X(\update_output_0/n1550 ) );
  nor_x1_sg U10818 ( .A(n6784), .B(n7185), .X(\update_output_0/n1546 ) );
  nor_x1_sg U10819 ( .A(n6732), .B(n6182), .X(\update_output_0/n2818 ) );
  nor_x1_sg U10820 ( .A(n5940), .B(n6183), .X(\update_output_0/n2814 ) );
  nor_x1_sg U10821 ( .A(n6750), .B(n7104), .X(\update_output_0/n2802 ) );
  nor_x1_sg U10822 ( .A(n6764), .B(n6183), .X(\update_output_0/n2798 ) );
  nor_x1_sg U10823 ( .A(n6755), .B(n6020), .X(\update_output_0/n2782 ) );
  nor_x1_sg U10824 ( .A(n6745), .B(n7104), .X(\update_output_0/n2774 ) );
  nor_x1_sg U10825 ( .A(n6741), .B(n6432), .X(\update_output_0/n2762 ) );
  nor_x1_sg U10826 ( .A(n6737), .B(n6019), .X(\update_output_0/n2758 ) );
  nor_x1_sg U10827 ( .A(n6730), .B(n6206), .X(\update_output_0/n2738 ) );
  nor_x1_sg U10828 ( .A(n6762), .B(n6046), .X(\update_output_0/n2734 ) );
  nor_x1_sg U10829 ( .A(n6751), .B(n7182), .X(\update_output_0/n2722 ) );
  nor_x1_sg U10830 ( .A(n5941), .B(n7180), .X(\update_output_0/n2718 ) );
  nor_x1_sg U10831 ( .A(n6757), .B(n6414), .X(\update_output_0/n2702 ) );
  nor_x1_sg U10832 ( .A(n6744), .B(n7180), .X(\update_output_0/n2694 ) );
  nor_x1_sg U10833 ( .A(n6740), .B(n7179), .X(\update_output_0/n2682 ) );
  nor_x1_sg U10834 ( .A(n6735), .B(n7180), .X(\update_output_0/n2678 ) );
  nor_x1_sg U10835 ( .A(n6731), .B(n7220), .X(\update_output_0/n2658 ) );
  nor_x1_sg U10836 ( .A(n6760), .B(n6398), .X(\update_output_0/n2654 ) );
  nor_x1_sg U10837 ( .A(n6751), .B(n6070), .X(\update_output_0/n2642 ) );
  nor_x1_sg U10838 ( .A(n5941), .B(n7219), .X(\update_output_0/n2638 ) );
  nor_x1_sg U10839 ( .A(n6757), .B(n6071), .X(\update_output_0/n2622 ) );
  nor_x1_sg U10840 ( .A(n6747), .B(n6070), .X(\update_output_0/n2614 ) );
  nor_x1_sg U10841 ( .A(n6739), .B(n6231), .X(\update_output_0/n2602 ) );
  nor_x1_sg U10842 ( .A(n6736), .B(n6230), .X(\update_output_0/n2598 ) );
  nor_x1_sg U10843 ( .A(n5929), .B(n7177), .X(\update_output_0/n2578 ) );
  nor_x1_sg U10844 ( .A(n6761), .B(n7175), .X(\update_output_0/n2574 ) );
  nor_x1_sg U10845 ( .A(n6749), .B(n7177), .X(\update_output_0/n2562 ) );
  nor_x1_sg U10846 ( .A(n6765), .B(n6204), .X(\update_output_0/n2558 ) );
  nor_x1_sg U10847 ( .A(n6755), .B(n6043), .X(\update_output_0/n2542 ) );
  nor_x1_sg U10848 ( .A(n5935), .B(n6204), .X(\update_output_0/n2534 ) );
  nor_x1_sg U10849 ( .A(n6742), .B(n7175), .X(\update_output_0/n2522 ) );
  nor_x1_sg U10850 ( .A(n5931), .B(n6044), .X(\update_output_0/n2518 ) );
  nor_x1_sg U10851 ( .A(n6731), .B(n7118), .X(\update_output_0/n2498 ) );
  nor_x1_sg U10852 ( .A(n6760), .B(n7121), .X(\update_output_0/n2494 ) );
  nor_x1_sg U10853 ( .A(n6751), .B(n6192), .X(\update_output_0/n2482 ) );
  nor_x1_sg U10854 ( .A(n6766), .B(n6425), .X(\update_output_0/n2478 ) );
  nor_x1_sg U10855 ( .A(n6754), .B(n6192), .X(\update_output_0/n2462 ) );
  nor_x1_sg U10856 ( .A(n6745), .B(n6192), .X(\update_output_0/n2454 ) );
  nor_x1_sg U10857 ( .A(n6740), .B(n7119), .X(\update_output_0/n2442 ) );
  nor_x1_sg U10858 ( .A(n6737), .B(n7118), .X(\update_output_0/n2438 ) );
  nor_x1_sg U10859 ( .A(n6730), .B(n6401), .X(\update_output_0/n2418 ) );
  nor_x1_sg U10860 ( .A(n6761), .B(n7209), .X(\update_output_0/n2414 ) );
  nor_x1_sg U10861 ( .A(n6750), .B(n6065), .X(\update_output_0/n2402 ) );
  nor_x1_sg U10862 ( .A(n6764), .B(n6064), .X(\update_output_0/n2398 ) );
  nor_x1_sg U10863 ( .A(n5938), .B(n6402), .X(\update_output_0/n2382 ) );
  nor_x1_sg U10864 ( .A(n6745), .B(n6064), .X(\update_output_0/n2374 ) );
  nor_x1_sg U10865 ( .A(n6739), .B(n6402), .X(\update_output_0/n2362 ) );
  nor_x1_sg U10866 ( .A(n6735), .B(n7209), .X(\update_output_0/n2358 ) );
  nor_x1_sg U10867 ( .A(n6732), .B(n6403), .X(\update_output_0/n2338 ) );
  nor_x1_sg U10868 ( .A(n6759), .B(n7206), .X(\update_output_0/n2334 ) );
  nor_x1_sg U10869 ( .A(n6751), .B(n6404), .X(\update_output_0/n2322 ) );
  nor_x1_sg U10870 ( .A(n6765), .B(n7206), .X(\update_output_0/n2318 ) );
  nor_x1_sg U10871 ( .A(n6756), .B(n6221), .X(\update_output_0/n2302 ) );
  nor_x1_sg U10872 ( .A(n6744), .B(n7206), .X(\update_output_0/n2294 ) );
  nor_x1_sg U10873 ( .A(n5933), .B(n7205), .X(\update_output_0/n2282 ) );
  nor_x1_sg U10874 ( .A(n6735), .B(n6222), .X(\update_output_0/n2278 ) );
  nor_x1_sg U10875 ( .A(n6729), .B(n6218), .X(\update_output_0/n2258 ) );
  nor_x1_sg U10876 ( .A(n6759), .B(n6058), .X(\update_output_0/n2254 ) );
  nor_x1_sg U10877 ( .A(n5936), .B(n7202), .X(\update_output_0/n2242 ) );
  nor_x1_sg U10878 ( .A(n6767), .B(n7200), .X(\update_output_0/n2238 ) );
  nor_x1_sg U10879 ( .A(n6756), .B(n6406), .X(\update_output_0/n2222 ) );
  nor_x1_sg U10880 ( .A(n6746), .B(n7200), .X(\update_output_0/n2214 ) );
  nor_x1_sg U10881 ( .A(n6740), .B(n7199), .X(\update_output_0/n2202 ) );
  nor_x1_sg U10882 ( .A(n6735), .B(n7200), .X(\update_output_0/n2198 ) );
  nor_x1_sg U10883 ( .A(n6732), .B(n6188), .X(\update_output_0/n2178 ) );
  nor_x1_sg U10884 ( .A(n6762), .B(n6188), .X(\update_output_0/n2174 ) );
  nor_x1_sg U10885 ( .A(n6749), .B(n6188), .X(\update_output_0/n2162 ) );
  nor_x1_sg U10886 ( .A(n6767), .B(n6428), .X(\update_output_0/n2158 ) );
  nor_x1_sg U10887 ( .A(n6757), .B(n7115), .X(\update_output_0/n2142 ) );
  nor_x1_sg U10888 ( .A(n6747), .B(n6428), .X(\update_output_0/n2134 ) );
  nor_x1_sg U10889 ( .A(n6741), .B(n6025), .X(\update_output_0/n2122 ) );
  nor_x1_sg U10890 ( .A(n6736), .B(n7114), .X(\update_output_0/n2118 ) );
  nor_x1_sg U10891 ( .A(n6730), .B(n6417), .X(\update_output_0/n2098 ) );
  nor_x1_sg U10892 ( .A(n6762), .B(n7171), .X(\update_output_0/n2094 ) );
  nor_x1_sg U10893 ( .A(n6750), .B(n6418), .X(\update_output_0/n2082 ) );
  nor_x1_sg U10894 ( .A(n6767), .B(n7171), .X(\update_output_0/n2078 ) );
  nor_x1_sg U10895 ( .A(n6754), .B(n6201), .X(\update_output_0/n2062 ) );
  nor_x1_sg U10896 ( .A(n6747), .B(n7171), .X(\update_output_0/n2054 ) );
  nor_x1_sg U10897 ( .A(n5933), .B(n7170), .X(\update_output_0/n2042 ) );
  nor_x1_sg U10898 ( .A(n6734), .B(n7172), .X(\update_output_0/n2038 ) );
  nor_x1_sg U10899 ( .A(n6730), .B(n6228), .X(\update_output_0/n2018 ) );
  nor_x1_sg U10900 ( .A(n6761), .B(n7214), .X(\update_output_0/n2014 ) );
  nor_x1_sg U10901 ( .A(n6752), .B(n6399), .X(\update_output_0/n2002 ) );
  nor_x1_sg U10902 ( .A(n6766), .B(n6400), .X(\update_output_0/n1998 ) );
  nor_x1_sg U10903 ( .A(n6756), .B(n6067), .X(\update_output_0/n1982 ) );
  nor_x1_sg U10904 ( .A(n6746), .B(n6068), .X(\update_output_0/n1974 ) );
  nor_x1_sg U10905 ( .A(n6742), .B(n6068), .X(\update_output_0/n1962 ) );
  nor_x1_sg U10906 ( .A(n5931), .B(n6227), .X(\update_output_0/n1958 ) );
  nor_x1_sg U10907 ( .A(n6731), .B(n6420), .X(\update_output_0/n1938 ) );
  nor_x1_sg U10908 ( .A(n6761), .B(n6037), .X(\update_output_0/n1934 ) );
  nor_x1_sg U10909 ( .A(n6750), .B(n6420), .X(\update_output_0/n1922 ) );
  nor_x1_sg U10910 ( .A(n6765), .B(n7167), .X(\update_output_0/n1918 ) );
  nor_x1_sg U10911 ( .A(n6755), .B(n6197), .X(\update_output_0/n1902 ) );
  nor_x1_sg U10912 ( .A(n6746), .B(n6420), .X(\update_output_0/n1894 ) );
  nor_x1_sg U10913 ( .A(n6742), .B(n7164), .X(\update_output_0/n1882 ) );
  nor_x1_sg U10914 ( .A(n6734), .B(n7166), .X(\update_output_0/n1878 ) );
  nor_x1_sg U10915 ( .A(n5929), .B(n6429), .X(\update_output_0/n1858 ) );
  nor_x1_sg U10916 ( .A(n6760), .B(n7110), .X(\update_output_0/n1854 ) );
  nor_x1_sg U10917 ( .A(n5936), .B(n6430), .X(\update_output_0/n1842 ) );
  nor_x1_sg U10918 ( .A(n6766), .B(n7110), .X(\update_output_0/n1838 ) );
  nor_x1_sg U10919 ( .A(n6756), .B(n6185), .X(\update_output_0/n1822 ) );
  nor_x1_sg U10920 ( .A(n6745), .B(n7110), .X(\update_output_0/n1814 ) );
  nor_x1_sg U10921 ( .A(n6742), .B(n7109), .X(\update_output_0/n1802 ) );
  nor_x1_sg U10922 ( .A(n6737), .B(n6186), .X(\update_output_0/n1798 ) );
  nor_x1_sg U10923 ( .A(n6732), .B(n7197), .X(\update_output_0/n1778 ) );
  nor_x1_sg U10924 ( .A(n6762), .B(n6407), .X(\update_output_0/n1774 ) );
  nor_x1_sg U10925 ( .A(n6752), .B(n6216), .X(\update_output_0/n1762 ) );
  nor_x1_sg U10926 ( .A(n6767), .B(n6056), .X(\update_output_0/n1758 ) );
  nor_x1_sg U10927 ( .A(n6757), .B(n6215), .X(\update_output_0/n1742 ) );
  nor_x1_sg U10928 ( .A(n6747), .B(n6408), .X(\update_output_0/n1734 ) );
  nor_x1_sg U10929 ( .A(n6741), .B(n7196), .X(\update_output_0/n1722 ) );
  nor_x1_sg U10930 ( .A(n6736), .B(n6216), .X(\update_output_0/n1718 ) );
  nor_x1_sg U10931 ( .A(n6729), .B(n6053), .X(\update_output_0/n1698 ) );
  nor_x1_sg U10932 ( .A(n6760), .B(n6409), .X(\update_output_0/n1694 ) );
  nor_x1_sg U10933 ( .A(n6752), .B(n7190), .X(\update_output_0/n1682 ) );
  nor_x1_sg U10934 ( .A(n6765), .B(n7191), .X(\update_output_0/n1678 ) );
  nor_x1_sg U10935 ( .A(n5938), .B(n7189), .X(\update_output_0/n1662 ) );
  nor_x1_sg U10936 ( .A(n6746), .B(n6052), .X(\update_output_0/n1654 ) );
  nor_x1_sg U10937 ( .A(n6740), .B(n6212), .X(\update_output_0/n1642 ) );
  nor_x1_sg U10938 ( .A(n6737), .B(n6410), .X(\update_output_0/n1638 ) );
  nor_x1_sg U10939 ( .A(n6731), .B(n6050), .X(\update_output_0/n1618 ) );
  nor_x1_sg U10940 ( .A(n5940), .B(n7185), .X(\update_output_0/n1614 ) );
  nor_x1_sg U10941 ( .A(n6752), .B(n7187), .X(\update_output_0/n1602 ) );
  nor_x1_sg U10942 ( .A(n6766), .B(n6411), .X(\update_output_0/n1598 ) );
  nor_x1_sg U10943 ( .A(n6755), .B(n7186), .X(\update_output_0/n1582 ) );
  nor_x1_sg U10944 ( .A(n5935), .B(n6210), .X(\update_output_0/n1574 ) );
  nor_x1_sg U10945 ( .A(n6741), .B(n6412), .X(\update_output_0/n1562 ) );
  nor_x1_sg U10946 ( .A(n6736), .B(n6209), .X(\update_output_0/n1558 ) );
  nor_x1_sg U10947 ( .A(n6542), .B(n6339), .X(\update_mask_0/n1053 ) );
  nor_x1_sg U10948 ( .A(n6542), .B(n6341), .X(\update_mask_0/n1021 ) );
  nor_x1_sg U10949 ( .A(n6540), .B(n6350), .X(\update_mask_0/n989 ) );
  nor_x1_sg U10950 ( .A(n6542), .B(n6345), .X(\update_mask_0/n957 ) );
  nor_x1_sg U10951 ( .A(n1452), .B(n6339), .X(\update_mask_0/n949 ) );
  nor_x1_sg U10952 ( .A(n1452), .B(n6342), .X(\update_mask_0/n1049 ) );
  nor_x1_sg U10953 ( .A(n6371), .B(n6351), .X(\update_mask_0/n1017 ) );
  nor_x1_sg U10954 ( .A(n6372), .B(n6345), .X(\update_mask_0/n985 ) );
  nand_x1_sg U10955 ( .A(n7016), .B(n1473), .X(\update_mask_0/n948 ) );
  nand_x1_sg U10956 ( .A(n6316), .B(n7457), .X(n1473) );
  nand_x1_sg U10957 ( .A(n6363), .B(n1474), .X(\update_mask_0/n1076 ) );
  nand_x1_sg U10958 ( .A(n7412), .B(n7456), .X(n1474) );
  nand_x1_sg U10959 ( .A(n7017), .B(n1475), .X(\update_mask_0/n1072 ) );
  nand_x1_sg U10960 ( .A(n6316), .B(n7441), .X(n1475) );
  nand_x1_sg U10961 ( .A(n6364), .B(n1476), .X(\update_mask_0/n1068 ) );
  nand_x1_sg U10962 ( .A(n7412), .B(n7413), .X(n1476) );
  nand_x1_sg U10963 ( .A(n7017), .B(n1477), .X(\update_mask_0/n1064 ) );
  nand_x1_sg U10964 ( .A(n7412), .B(n8897), .X(n1477) );
  nand_x1_sg U10965 ( .A(n7016), .B(n1478), .X(\update_mask_0/n1060 ) );
  nand_x1_sg U10966 ( .A(n6316), .B(n7392), .X(n1478) );
  nand_x1_sg U10967 ( .A(n7018), .B(n1479), .X(\update_mask_0/n1056 ) );
  nand_x1_sg U10968 ( .A(n7412), .B(n7393), .X(n1479) );
  nand_x1_sg U10969 ( .A(n6121), .B(n1481), .X(\update_mask_0/n1052 ) );
  nand_x1_sg U10970 ( .A(n6316), .B(n7390), .X(n1481) );
  nand_x1_sg U10971 ( .A(n7018), .B(n1484), .X(\update_mask_0/n1048 ) );
  nand_x1_sg U10972 ( .A(n7411), .B(n7457), .X(n1484) );
  nand_x1_sg U10973 ( .A(n5984), .B(n1485), .X(\update_mask_0/n1044 ) );
  nand_x1_sg U10974 ( .A(n6317), .B(n7456), .X(n1485) );
  nand_x1_sg U10975 ( .A(n6363), .B(n1486), .X(\update_mask_0/n1040 ) );
  nand_x1_sg U10976 ( .A(n7411), .B(n7441), .X(n1486) );
  nand_x1_sg U10977 ( .A(n7018), .B(n1487), .X(\update_mask_0/n1036 ) );
  nand_x1_sg U10978 ( .A(n6317), .B(n7413), .X(n1487) );
  nand_x1_sg U10979 ( .A(n6121), .B(n1488), .X(\update_mask_0/n1032 ) );
  nand_x1_sg U10980 ( .A(n7411), .B(n8897), .X(n1488) );
  nand_x1_sg U10981 ( .A(n7019), .B(n1489), .X(\update_mask_0/n1028 ) );
  nand_x1_sg U10982 ( .A(n6317), .B(n7392), .X(n1489) );
  nand_x1_sg U10983 ( .A(n7017), .B(n1490), .X(\update_mask_0/n1024 ) );
  nand_x1_sg U10984 ( .A(n7411), .B(n7393), .X(n1490) );
  nand_x1_sg U10985 ( .A(n7017), .B(n1492), .X(\update_mask_0/n1020 ) );
  nand_x1_sg U10986 ( .A(n6317), .B(n7390), .X(n1492) );
  nand_x1_sg U10987 ( .A(n6121), .B(n1494), .X(\update_mask_0/n1016 ) );
  nand_x1_sg U10988 ( .A(n7410), .B(n7457), .X(n1494) );
  nand_x1_sg U10989 ( .A(n6122), .B(n1495), .X(\update_mask_0/n1012 ) );
  nand_x1_sg U10990 ( .A(n6318), .B(n7456), .X(n1495) );
  nand_x1_sg U10991 ( .A(n7018), .B(n1496), .X(\update_mask_0/n1008 ) );
  nand_x1_sg U10992 ( .A(n7410), .B(n7441), .X(n1496) );
  nand_x1_sg U10993 ( .A(n6122), .B(n1497), .X(\update_mask_0/n1004 ) );
  nand_x1_sg U10994 ( .A(n6318), .B(n7413), .X(n1497) );
  nand_x1_sg U10995 ( .A(n7019), .B(n1499), .X(\update_mask_0/n1000 ) );
  nand_x1_sg U10996 ( .A(n7410), .B(n8897), .X(n1499) );
  nand_x1_sg U10997 ( .A(n6363), .B(n1448), .X(\update_mask_0/n996 ) );
  nand_x1_sg U10998 ( .A(n6318), .B(n7392), .X(n1448) );
  nand_x1_sg U10999 ( .A(n7019), .B(n1450), .X(\update_mask_0/n992 ) );
  nand_x1_sg U11000 ( .A(n7410), .B(n7393), .X(n1450) );
  nand_x1_sg U11001 ( .A(n6364), .B(n1451), .X(\update_mask_0/n988 ) );
  nand_x1_sg U11002 ( .A(n6318), .B(n7390), .X(n1451) );
  nand_x1_sg U11003 ( .A(n5984), .B(n1454), .X(\update_mask_0/n984 ) );
  nand_x1_sg U11004 ( .A(n7409), .B(n7457), .X(n1454) );
  nand_x1_sg U11005 ( .A(n6364), .B(n1456), .X(\update_mask_0/n980 ) );
  nand_x1_sg U11006 ( .A(n6319), .B(n7456), .X(n1456) );
  nand_x1_sg U11007 ( .A(n6121), .B(n1458), .X(\update_mask_0/n976 ) );
  nand_x1_sg U11008 ( .A(n7409), .B(n7441), .X(n1458) );
  nand_x1_sg U11009 ( .A(n6122), .B(n1460), .X(\update_mask_0/n972 ) );
  nand_x1_sg U11010 ( .A(n6319), .B(n7413), .X(n1460) );
  nand_x1_sg U11011 ( .A(n6363), .B(n1462), .X(\update_mask_0/n968 ) );
  nand_x1_sg U11012 ( .A(n7409), .B(n8897), .X(n1462) );
  nand_x1_sg U11013 ( .A(n6122), .B(n1463), .X(\update_mask_0/n964 ) );
  nand_x1_sg U11014 ( .A(n6319), .B(n6346), .X(n1463) );
  nand_x1_sg U11015 ( .A(n6364), .B(n1464), .X(\update_mask_0/n960 ) );
  nand_x1_sg U11016 ( .A(n7409), .B(n6352), .X(n1464) );
  nand_x1_sg U11017 ( .A(n7019), .B(n1467), .X(\update_mask_0/n956 ) );
  nand_x1_sg U11018 ( .A(n6319), .B(n7390), .X(n1467) );
  nor_x1_sg U11019 ( .A(n6508), .B(n7398), .X(n3696) );
  nand_x4_sg U11020 ( .A(n1305), .B(n1306), .X(n1301) );
  nand_x1_sg U11021 ( .A(n7144), .B(n9168), .X(n1303) );
  nand_x1_sg U11022 ( .A(n8968), .B(n1288), .X(n1287) );
  nor_x1_sg U11023 ( .A(n6362), .B(n1292), .X(n1290) );
  nand_x4_sg U11024 ( .A(n1009), .B(n1010), .X(n1005) );
  nand_x1_sg U11025 ( .A(n6240), .B(n1311), .X(n1310) );
  nand_x1_sg U11026 ( .A(n1312), .B(n9128), .X(n1309) );
  nand_x4_sg U11027 ( .A(n1273), .B(n1274), .X(n1269) );
  nand_x1_sg U11028 ( .A(n6323), .B(n9167), .X(n1271) );
  nand_x1_sg U11029 ( .A(n9003), .B(n1134), .X(n1130) );
  nand_x1_sg U11030 ( .A(n7260), .B(n9063), .X(n1133) );
  nand_x1_sg U11031 ( .A(n9007), .B(n1265), .X(n1261) );
  nand_x1_sg U11032 ( .A(n7268), .B(n9067), .X(n1264) );
  nand_x1_sg U11033 ( .A(n9017), .B(n805), .X(n800) );
  nand_x1_sg U11034 ( .A(n7271), .B(n9077), .X(n803) );
  nand_x1_sg U11035 ( .A(n7318), .B(n1015), .X(n1014) );
  nand_x1_sg U11036 ( .A(n7281), .B(n9212), .X(n1015) );
  nor_x1_sg U11037 ( .A(n1178), .B(n1179), .X(n1168) );
  nand_x1_sg U11038 ( .A(n5927), .B(n1148), .X(n1147) );
  nand_x1_sg U11039 ( .A(n1149), .B(n9123), .X(n1146) );
  nand_x1_sg U11040 ( .A(n6129), .B(n9203), .X(n1148) );
  nand_x1_sg U11041 ( .A(n6241), .B(n820), .X(n819) );
  nand_x1_sg U11042 ( .A(n821), .B(n9137), .X(n818) );
  nand_x1_sg U11043 ( .A(n6490), .B(n9217), .X(n820) );
  nand_x1_sg U11044 ( .A(n7319), .B(n983), .X(n982) );
  nand_x1_sg U11045 ( .A(n7280), .B(n9214), .X(n983) );
  nand_x1_sg U11046 ( .A(n9004), .B(n1166), .X(n1162) );
  nand_x1_sg U11047 ( .A(n7261), .B(n9064), .X(n1165) );
  nand_x1_sg U11048 ( .A(n9018), .B(n838), .X(n834) );
  nand_x1_sg U11049 ( .A(n7271), .B(n9078), .X(n837) );
  nand_x4_sg U11050 ( .A(n1258), .B(n8987), .X(n1254) );
  nand_x1_sg U11051 ( .A(n8967), .B(n1256), .X(n1255) );
  inv_x1_sg U11052 ( .A(n1259), .X(n8987) );
  nand_x4_sg U11053 ( .A(n1174), .B(n1175), .X(n1170) );
  nand_x1_sg U11054 ( .A(n6034), .B(n9164), .X(n1172) );
  nand_x1_sg U11055 ( .A(n7322), .B(n852), .X(n851) );
  nand_x1_sg U11056 ( .A(n853), .B(n9138), .X(n850) );
  nand_x1_sg U11057 ( .A(n7278), .B(n9218), .X(n852) );
  nand_x4_sg U11058 ( .A(n962), .B(n8994), .X(n958) );
  nand_x1_sg U11059 ( .A(n8974), .B(n960), .X(n959) );
  inv_x1_sg U11060 ( .A(n963), .X(n8994) );
  nand_x4_sg U11061 ( .A(n1159), .B(n8984), .X(n1155) );
  nand_x1_sg U11062 ( .A(n8964), .B(n1157), .X(n1156) );
  inv_x1_sg U11063 ( .A(n1160), .X(n8984) );
  nand_x4_sg U11064 ( .A(n1127), .B(n8983), .X(n1123) );
  nand_x1_sg U11065 ( .A(n8963), .B(n1125), .X(n1124) );
  inv_x1_sg U11066 ( .A(n1128), .X(n8983) );
  nand_x4_sg U11067 ( .A(n831), .B(n8998), .X(n827) );
  nand_x1_sg U11068 ( .A(n8978), .B(n829), .X(n828) );
  inv_x1_sg U11069 ( .A(n832), .X(n8998) );
  nand_x4_sg U11070 ( .A(n795), .B(n8997), .X(n789) );
  nand_x1_sg U11071 ( .A(n8977), .B(n791), .X(n790) );
  inv_x1_sg U11072 ( .A(n796), .X(n8997) );
  nand_x4_sg U11073 ( .A(n1401), .B(n1402), .X(n1397) );
  inv_x1_sg U11074 ( .A(n1400), .X(n9111) );
  nand_x1_sg U11075 ( .A(n8971), .B(n1384), .X(n1383) );
  nor_x1_sg U11076 ( .A(n7318), .B(n1388), .X(n1386) );
  nand_x4_sg U11077 ( .A(n1337), .B(n1338), .X(n1333) );
  nand_x1_sg U11078 ( .A(n6323), .B(n9169), .X(n1335) );
  nand_x1_sg U11079 ( .A(n7318), .B(n1407), .X(n1406) );
  nand_x1_sg U11080 ( .A(n1408), .B(n9131), .X(n1405) );
  nand_x1_sg U11081 ( .A(n3567), .B(n6315), .X(n3566) );
  nand_x1_sg U11082 ( .A(n8969), .B(n1320), .X(n1319) );
  nor_x1_sg U11083 ( .A(n7320), .B(n1324), .X(n1322) );
  nand_x4_sg U11084 ( .A(n1238), .B(n1239), .X(n1234) );
  nand_x1_sg U11085 ( .A(n7144), .B(n9165), .X(n1236) );
  nand_x4_sg U11086 ( .A(n1041), .B(n1042), .X(n1037) );
  nand_x1_sg U11087 ( .A(n6240), .B(n1343), .X(n1342) );
  nand_x1_sg U11088 ( .A(n1344), .B(n9129), .X(n1341) );
  nand_x1_sg U11089 ( .A(n6083), .B(n1111), .X(n1110) );
  nand_x1_sg U11090 ( .A(n1112), .B(n9136), .X(n1109) );
  nand_x1_sg U11091 ( .A(n6390), .B(n9216), .X(n1111) );
  nand_x4_sg U11092 ( .A(n1369), .B(n1370), .X(n1365) );
  nand_x1_sg U11093 ( .A(n7146), .B(n9170), .X(n1367) );
  nand_x1_sg U11094 ( .A(n8965), .B(n1221), .X(n1220) );
  nor_x1_sg U11095 ( .A(n6082), .B(n1225), .X(n1223) );
  nand_x1_sg U11096 ( .A(n8973), .B(n1024), .X(n1023) );
  nor_x1_sg U11097 ( .A(n7321), .B(n1028), .X(n1026) );
  nand_x1_sg U11098 ( .A(n7319), .B(n1047), .X(n1046) );
  nand_x1_sg U11099 ( .A(n6491), .B(n9213), .X(n1047) );
  nand_x4_sg U11100 ( .A(n942), .B(n943), .X(n938) );
  nand_x1_sg U11101 ( .A(n6241), .B(n1244), .X(n1243) );
  nand_x1_sg U11102 ( .A(n1245), .B(n9125), .X(n1242) );
  nand_x1_sg U11103 ( .A(n9010), .B(n1361), .X(n1357) );
  nand_x1_sg U11104 ( .A(n7261), .B(n9070), .X(n1360) );
  nand_x1_sg U11105 ( .A(n9016), .B(n1097), .X(n1093) );
  nand_x1_sg U11106 ( .A(n7262), .B(n9076), .X(n1096) );
  nand_x1_sg U11107 ( .A(n9015), .B(n1065), .X(n1061) );
  nand_x1_sg U11108 ( .A(n7271), .B(n9075), .X(n1064) );
  nand_x4_sg U11109 ( .A(n1206), .B(n1207), .X(n1202) );
  nand_x1_sg U11110 ( .A(n6034), .B(n9166), .X(n1204) );
  nand_x1_sg U11111 ( .A(n7320), .B(n1375), .X(n1374) );
  nand_x1_sg U11112 ( .A(n1376), .B(n9130), .X(n1373) );
  nand_x1_sg U11113 ( .A(n9006), .B(n1198), .X(n1194) );
  nand_x1_sg U11114 ( .A(n7270), .B(n9066), .X(n1197) );
  nand_x1_sg U11115 ( .A(n9002), .B(n1425), .X(n1421) );
  nand_x1_sg U11116 ( .A(n7261), .B(n9062), .X(n1424) );
  nand_x1_sg U11117 ( .A(n9019), .B(n870), .X(n866) );
  nand_x1_sg U11118 ( .A(n7266), .B(n9079), .X(n869) );
  nand_x1_sg U11119 ( .A(n9020), .B(n902), .X(n898) );
  nand_x1_sg U11120 ( .A(n7268), .B(n9080), .X(n901) );
  nand_x1_sg U11121 ( .A(n5927), .B(n1441), .X(n1440) );
  nand_x1_sg U11122 ( .A(n1443), .B(n9122), .X(n1439) );
  nand_x1_sg U11123 ( .A(n7322), .B(n1079), .X(n1078) );
  nand_x1_sg U11124 ( .A(n1080), .B(n9135), .X(n1077) );
  nand_x1_sg U11125 ( .A(n7280), .B(n9215), .X(n1079) );
  nand_x1_sg U11126 ( .A(n6083), .B(n884), .X(n883) );
  nand_x1_sg U11127 ( .A(n885), .B(n9139), .X(n882) );
  nand_x1_sg U11128 ( .A(n6492), .B(n9219), .X(n884) );
  nand_x1_sg U11129 ( .A(n7321), .B(n916), .X(n915) );
  nand_x1_sg U11130 ( .A(n917), .B(n9140), .X(n914) );
  nand_x1_sg U11131 ( .A(n6490), .B(n9220), .X(n916) );
  nor_x1_sg U11132 ( .A(n7459), .B(n6458), .X(n806) );
  nand_x4_sg U11133 ( .A(n1058), .B(n8995), .X(n1054) );
  nand_x1_sg U11134 ( .A(n8975), .B(n1056), .X(n1055) );
  inv_x1_sg U11135 ( .A(n1059), .X(n8995) );
  nand_x1_sg U11136 ( .A(n6362), .B(n948), .X(n947) );
  nand_x1_sg U11137 ( .A(n7278), .B(n9221), .X(n948) );
  nand_x1_sg U11138 ( .A(n7319), .B(n1212), .X(n1211) );
  nand_x1_sg U11139 ( .A(n1213), .B(n9126), .X(n1210) );
  nand_x1_sg U11140 ( .A(n6129), .B(n9206), .X(n1212) );
  nand_x4_sg U11141 ( .A(n863), .B(n8999), .X(n859) );
  nand_x1_sg U11142 ( .A(n8979), .B(n861), .X(n860) );
  inv_x1_sg U11143 ( .A(n864), .X(n8999) );
  nand_x4_sg U11144 ( .A(n1418), .B(n8982), .X(n1414) );
  nand_x1_sg U11145 ( .A(n8962), .B(n1416), .X(n1415) );
  inv_x1_sg U11146 ( .A(n1419), .X(n8982) );
  nand_x4_sg U11147 ( .A(n1105), .B(n1106), .X(n1101) );
  nand_x1_sg U11148 ( .A(n6035), .B(n9176), .X(n1103) );
  nand_x4_sg U11149 ( .A(n895), .B(n9000), .X(n891) );
  nand_x1_sg U11150 ( .A(n8980), .B(n893), .X(n892) );
  inv_x1_sg U11151 ( .A(n896), .X(n9000) );
  nand_x1_sg U11152 ( .A(n3567), .B(n6320), .X(n3911) );
  nand_x1_sg U11153 ( .A(n4040), .B(n7408), .X(n4039) );
  nor_x1_sg U11154 ( .A(n6510), .B(n3783), .X(n4040) );
  nand_x1_sg U11155 ( .A(n4125), .B(n6320), .X(n4124) );
  nor_x1_sg U11156 ( .A(n7414), .B(n3783), .X(n4125) );
  nand_x1_sg U11157 ( .A(n6472), .B(n777), .X(n4821) );
  inv_x1_sg U11158 ( .A(n3783), .X(n9226) );
  nand_x1_sg U11159 ( .A(n7400), .B(n6311), .X(n3954) );
  nand_x1_sg U11160 ( .A(n7005), .B(n4785), .X(n4784) );
  nand_x1_sg U11161 ( .A(n7005), .B(n4713), .X(n4712) );
  nand_x1_sg U11162 ( .A(n7000), .B(n4209), .X(n4208) );
  nand_x1_sg U11163 ( .A(n7001), .B(n4131), .X(n4130) );
  nand_x1_sg U11164 ( .A(n7002), .B(n4749), .X(n4748) );
  nand_x1_sg U11165 ( .A(n7004), .B(n4461), .X(n4460) );
  nand_x1_sg U11166 ( .A(n7315), .B(n4838), .X(n4837) );
  nand_x1_sg U11167 ( .A(n6470), .B(n4800), .X(n4799) );
  nand_x1_sg U11168 ( .A(n7314), .B(n4764), .X(n4763) );
  nand_x1_sg U11169 ( .A(n6141), .B(n4728), .X(n4727) );
  nand_x1_sg U11170 ( .A(n6141), .B(n4692), .X(n4691) );
  nand_x1_sg U11171 ( .A(n6469), .B(n4656), .X(n4655) );
  nand_x1_sg U11172 ( .A(n6469), .B(n4620), .X(n4619) );
  nand_x1_sg U11173 ( .A(n6472), .B(n4584), .X(n4583) );
  nand_x1_sg U11174 ( .A(n6474), .B(n4548), .X(n4547) );
  nand_x1_sg U11175 ( .A(n6140), .B(n4512), .X(n4511) );
  nand_x1_sg U11176 ( .A(n6474), .B(n4476), .X(n4475) );
  nand_x1_sg U11177 ( .A(n7316), .B(n4440), .X(n4439) );
  nand_x1_sg U11178 ( .A(n6141), .B(n4260), .X(n4259) );
  nand_x1_sg U11179 ( .A(n6473), .B(n4224), .X(n4223) );
  nand_x1_sg U11180 ( .A(n6080), .B(n4188), .X(n4187) );
  nand_x1_sg U11181 ( .A(n7316), .B(n4150), .X(n4149) );
  nor_x1_sg U11182 ( .A(n6311), .B(n6508), .X(n4849) );
  nor_x1_sg U11183 ( .A(n7404), .B(n3466), .X(n3826) );
  nor_x1_sg U11184 ( .A(n6097), .B(n7403), .X(n2262) );
  nor_x1_sg U11185 ( .A(n4883), .B(n4884), .X(n4878) );
  nand_x1_sg U11186 ( .A(n6159), .B(n9237), .X(n4883) );
  inv_x1_sg U11187 ( .A(n4879), .X(n9237) );
  nand_x1_sg U11188 ( .A(n7314), .B(n3463), .X(n3459) );
  nand_x1_sg U11189 ( .A(n3461), .B(n6495), .X(n3460) );
  nand_x1_sg U11190 ( .A(n3464), .B(n3465), .X(n3463) );
  nor_x1_sg U11191 ( .A(n7401), .B(n3471), .X(n3739) );
  nand_x1_sg U11192 ( .A(n7397), .B(n7401), .X(n3997) );
  nor_x1_sg U11193 ( .A(n6509), .B(n3869), .X(n3523) );
  nand_x1_sg U11194 ( .A(n6510), .B(n7400), .X(n3474) );
  nor_x1_sg U11195 ( .A(n3474), .B(n6311), .X(n4151) );
  nand_x1_sg U11196 ( .A(n3439), .B(n6491), .X(n3438) );
  nand_x1_sg U11197 ( .A(n6361), .B(n3440), .X(n3437) );
  nor_x1_sg U11198 ( .A(n7318), .B(n6263), .X(n3439) );
  nor_x1_sg U11199 ( .A(n6158), .B(n3464), .X(n3473) );
  nor_x1_sg U11200 ( .A(n5623), .B(n5624), .X(n5621) );
  nor_x1_sg U11201 ( .A(n7452), .B(n6482), .X(n5624) );
  nor_x1_sg U11202 ( .A(n5598), .B(n5602), .X(n5601) );
  nor_x1_sg U11203 ( .A(n4872), .B(n6366), .X(n5602) );
  nand_x1_sg U11204 ( .A(n4867), .B(n4865), .X(n5598) );
  nand_x1_sg U11205 ( .A(n7002), .B(n6458), .X(n3432) );
  nand_x1_sg U11206 ( .A(n4867), .B(n5606), .X(n4875) );
  nand_x1_sg U11207 ( .A(n6460), .B(n6541), .X(n5606) );
  nand_x1_sg U11208 ( .A(n6462), .B(n7405), .X(n4874) );
  nand_x1_sg U11209 ( .A(n6462), .B(n7424), .X(n5617) );
  nand_x1_sg U11210 ( .A(n6461), .B(n7389), .X(n4865) );
  nand_x1_sg U11211 ( .A(n5597), .B(n6460), .X(n5596) );
  nand_x1_sg U11212 ( .A(n6366), .B(n5598), .X(n5595) );
  nand_x1_sg U11213 ( .A(n6505), .B(n5612), .X(n5608) );
  nand_x1_sg U11214 ( .A(n7424), .B(n5614), .X(n5612) );
  nand_x1_sg U11215 ( .A(n7004), .B(n3479), .X(n3478) );
  nand_x1_sg U11216 ( .A(n7005), .B(n3466), .X(n3465) );
  nor_x1_sg U11217 ( .A(n7440), .B(n6099), .X(n2180) );
  nand_x1_sg U11218 ( .A(n5626), .B(n6461), .X(n5630) );
  nor_x1_sg U11219 ( .A(n6504), .B(n7309), .X(n5610) );
  nor_x1_sg U11220 ( .A(n3452), .B(n3453), .X(n3451) );
  nor_x1_sg U11221 ( .A(n6367), .B(n7389), .X(n5597) );
  nand_x1_sg U11222 ( .A(n9235), .B(n9236), .X(n5643) );
  nor_x1_sg U11223 ( .A(n8961), .B(n1470), .X(n1466) );
  nor_x1_sg U11224 ( .A(n1502), .B(n1471), .X(n1501) );
  nor_x1_sg U11225 ( .A(n1470), .B(n1466), .X(n1469) );
  nor_x1_sg U11226 ( .A(n765), .B(n7398), .X(n760) );
  nor_x1_sg U11227 ( .A(n765), .B(n4821), .X(n773) );
  nand_x1_sg U11228 ( .A(n1480), .B(n1469), .X(n1482) );
  nand_x1_sg U11229 ( .A(n1491), .B(n1469), .X(n1493) );
  nand_x1_sg U11230 ( .A(n1498), .B(n1469), .X(n1500) );
  nor_x1_sg U11231 ( .A(n7405), .B(n7407), .X(n1465) );
  inv_x1_sg U11232 ( .A(n6384), .X(n8897) );
  nand_x1_sg U11233 ( .A(n7373), .B(n6311), .X(n771) );
  nand_x1_sg U11234 ( .A(n760), .B(n761), .X(n759) );
  nand_x1_sg U11235 ( .A(n767), .B(n761), .X(n766) );
  nand_x1_sg U11236 ( .A(n773), .B(n761), .X(n772) );
  nand_x4_sg U11237 ( .A(n1553), .B(n1554), .X(n1552) );
  nor_x1_sg U11238 ( .A(n1564), .B(n1565), .X(n1559) );
  nand_x4_sg U11239 ( .A(n1570), .B(n1571), .X(n1569) );
  nor_x1_sg U11240 ( .A(n1581), .B(n1582), .X(n1576) );
  nand_x4_sg U11241 ( .A(n1636), .B(n1637), .X(n1635) );
  nor_x1_sg U11242 ( .A(n1647), .B(n1648), .X(n1641) );
  nand_x4_sg U11243 ( .A(n1653), .B(n1654), .X(n1652) );
  nor_x1_sg U11244 ( .A(n1664), .B(n1665), .X(n1658) );
  nand_x4_sg U11245 ( .A(n1721), .B(n1722), .X(n1720) );
  nor_x1_sg U11246 ( .A(n1732), .B(n1733), .X(n1727) );
  nand_x4_sg U11247 ( .A(n1738), .B(n1739), .X(n1737) );
  nor_x1_sg U11248 ( .A(n1749), .B(n1750), .X(n1744) );
  nand_x4_sg U11249 ( .A(n1891), .B(n1892), .X(n1890) );
  nor_x1_sg U11250 ( .A(n1902), .B(n1903), .X(n1897) );
  nand_x4_sg U11251 ( .A(n1908), .B(n1909), .X(n1907) );
  nor_x1_sg U11252 ( .A(n1919), .B(n1920), .X(n1914) );
  nand_x4_sg U11253 ( .A(n1974), .B(n1975), .X(n1973) );
  nor_x1_sg U11254 ( .A(n1985), .B(n1986), .X(n1979) );
  nand_x4_sg U11255 ( .A(n1991), .B(n1992), .X(n1990) );
  nor_x1_sg U11256 ( .A(n2002), .B(n2003), .X(n1996) );
  nand_x4_sg U11257 ( .A(n2059), .B(n2060), .X(n2058) );
  nor_x1_sg U11258 ( .A(n2070), .B(n2071), .X(n2065) );
  nand_x4_sg U11259 ( .A(n2076), .B(n2077), .X(n2075) );
  nor_x1_sg U11260 ( .A(n2087), .B(n2088), .X(n2082) );
  nand_x1_sg U11261 ( .A(n761), .B(n756), .X(n734) );
  nand_x1_sg U11262 ( .A(n2186), .B(n7394), .X(n1526) );
  nand_x1_sg U11263 ( .A(n5623), .B(n7394), .X(n1524) );
  nand_x1_sg U11264 ( .A(n5626), .B(n7396), .X(n1534) );
  nor_x1_sg U11265 ( .A(n3452), .B(n777), .X(\update_output_0/n1542 ) );
  nor_x1_sg U11266 ( .A(n1817), .B(n1818), .X(n1766) );
  nor_x1_sg U11267 ( .A(n2155), .B(n2156), .X(n2104) );
  nor_x1_sg U11268 ( .A(n2228), .B(n2229), .X(n2227) );
  nand_x4_sg U11269 ( .A(n2255), .B(n2256), .X(n2245) );
  nor_x1_sg U11270 ( .A(n2197), .B(n8901), .X(n2196) );
  nand_x4_sg U11271 ( .A(n2201), .B(n2202), .X(n2197) );
  nor_x1_sg U11272 ( .A(n2199), .B(n2200), .X(n2198) );
  nor_x1_sg U11273 ( .A(n1537), .B(n8924), .X(n1536) );
  nand_x4_sg U11274 ( .A(n1541), .B(n8915), .X(n1537) );
  nor_x1_sg U11275 ( .A(n1539), .B(n1540), .X(n1538) );
  nor_x1_sg U11276 ( .A(n1605), .B(n8925), .X(n1604) );
  nand_x4_sg U11277 ( .A(n1609), .B(n8916), .X(n1605) );
  nor_x1_sg U11278 ( .A(n1607), .B(n1608), .X(n1606) );
  nor_x1_sg U11279 ( .A(n1705), .B(n8928), .X(n1704) );
  nand_x4_sg U11280 ( .A(n1709), .B(n8917), .X(n1705) );
  nor_x1_sg U11281 ( .A(n1707), .B(n1708), .X(n1706) );
  nor_x1_sg U11282 ( .A(n1875), .B(n8932), .X(n1874) );
  nand_x4_sg U11283 ( .A(n1879), .B(n8919), .X(n1875) );
  nor_x1_sg U11284 ( .A(n1877), .B(n1878), .X(n1876) );
  nor_x1_sg U11285 ( .A(n1943), .B(n8933), .X(n1942) );
  nand_x4_sg U11286 ( .A(n1947), .B(n8920), .X(n1943) );
  nor_x1_sg U11287 ( .A(n1945), .B(n1946), .X(n1944) );
  nor_x1_sg U11288 ( .A(n2043), .B(n8936), .X(n2042) );
  nand_x4_sg U11289 ( .A(n2047), .B(n8921), .X(n2043) );
  nor_x1_sg U11290 ( .A(n2045), .B(n2046), .X(n2044) );
  nor_x1_sg U11291 ( .A(n1516), .B(n8923), .X(n1515) );
  nand_x4_sg U11292 ( .A(n1522), .B(n8939), .X(n1516) );
  nor_x1_sg U11293 ( .A(n1518), .B(n1519), .X(n1517) );
  nor_x1_sg U11294 ( .A(n1620), .B(n8926), .X(n1619) );
  nand_x4_sg U11295 ( .A(n1624), .B(n8941), .X(n1620) );
  nor_x1_sg U11296 ( .A(n1622), .B(n1623), .X(n1621) );
  nor_x1_sg U11297 ( .A(n1690), .B(n8927), .X(n1689) );
  nand_x4_sg U11298 ( .A(n1694), .B(n8944), .X(n1690) );
  nor_x1_sg U11299 ( .A(n1692), .B(n1693), .X(n1691) );
  nor_x1_sg U11300 ( .A(n1788), .B(n8930), .X(n1787) );
  nand_x4_sg U11301 ( .A(n1792), .B(n8946), .X(n1788) );
  nor_x1_sg U11302 ( .A(n1790), .B(n1791), .X(n1789) );
  nor_x1_sg U11303 ( .A(n1860), .B(n8931), .X(n1859) );
  nand_x4_sg U11304 ( .A(n1864), .B(n8949), .X(n1860) );
  nor_x1_sg U11305 ( .A(n1862), .B(n1863), .X(n1861) );
  nor_x1_sg U11306 ( .A(n1958), .B(n8934), .X(n1957) );
  nand_x4_sg U11307 ( .A(n1962), .B(n8951), .X(n1958) );
  nor_x1_sg U11308 ( .A(n1960), .B(n1961), .X(n1959) );
  nor_x1_sg U11309 ( .A(n2028), .B(n8935), .X(n2027) );
  nand_x4_sg U11310 ( .A(n2032), .B(n8954), .X(n2028) );
  nor_x1_sg U11311 ( .A(n2030), .B(n2031), .X(n2029) );
  nor_x1_sg U11312 ( .A(n2126), .B(n8938), .X(n2125) );
  nand_x4_sg U11313 ( .A(n2130), .B(n8956), .X(n2126) );
  nor_x1_sg U11314 ( .A(n2128), .B(n2129), .X(n2127) );
  nor_x1_sg U11315 ( .A(n6347), .B(n6338), .X(\update_mask_0/n1061 ) );
  nor_x1_sg U11316 ( .A(n6348), .B(n6341), .X(\update_mask_0/n1029 ) );
  nor_x1_sg U11317 ( .A(n6348), .B(n6351), .X(\update_mask_0/n997 ) );
  nor_x1_sg U11318 ( .A(n6347), .B(n6344), .X(\update_mask_0/n965 ) );
  nor_x1_sg U11319 ( .A(n7446), .B(n6338), .X(\update_mask_0/n1065 ) );
  nor_x1_sg U11320 ( .A(n6383), .B(n6342), .X(\update_mask_0/n1033 ) );
  nor_x1_sg U11321 ( .A(n7446), .B(n6350), .X(\update_mask_0/n1001 ) );
  nor_x1_sg U11322 ( .A(n6383), .B(n6344), .X(\update_mask_0/n969 ) );
  nor_x1_sg U11323 ( .A(n6374), .B(n6339), .X(\update_mask_0/n1077 ) );
  nor_x1_sg U11324 ( .A(n6374), .B(n6342), .X(\update_mask_0/n1045 ) );
  nor_x1_sg U11325 ( .A(n6375), .B(n6350), .X(\update_mask_0/n1013 ) );
  nor_x1_sg U11326 ( .A(n1455), .B(n6345), .X(\update_mask_0/n981 ) );
  nor_x1_sg U11327 ( .A(n6354), .B(n6338), .X(\update_mask_0/n1057 ) );
  nor_x1_sg U11328 ( .A(n6353), .B(n6342), .X(\update_mask_0/n1025 ) );
  nor_x1_sg U11329 ( .A(n1449), .B(n6350), .X(\update_mask_0/n993 ) );
  nor_x1_sg U11330 ( .A(n6354), .B(n6344), .X(\update_mask_0/n961 ) );
  nor_x1_sg U11331 ( .A(n9222), .B(n3452), .X(\update_output_0/n1543 ) );
  nor_x1_sg U11332 ( .A(n6380), .B(n6339), .X(\update_mask_0/n1073 ) );
  nor_x1_sg U11333 ( .A(n6377), .B(n6338), .X(\update_mask_0/n1069 ) );
  nor_x1_sg U11334 ( .A(n7442), .B(n6341), .X(\update_mask_0/n1041 ) );
  nor_x1_sg U11335 ( .A(n6378), .B(n6341), .X(\update_mask_0/n1037 ) );
  nor_x1_sg U11336 ( .A(n6380), .B(n6351), .X(\update_mask_0/n1009 ) );
  nor_x1_sg U11337 ( .A(n6377), .B(n6351), .X(\update_mask_0/n1005 ) );
  nor_x1_sg U11338 ( .A(n7442), .B(n6344), .X(\update_mask_0/n977 ) );
  nor_x1_sg U11339 ( .A(n6378), .B(n6345), .X(\update_mask_0/n973 ) );
  nor_x1_sg U11340 ( .A(n1566), .B(n1567), .X(n1509) );
  nor_x1_sg U11341 ( .A(n1649), .B(n1650), .X(n1598) );
  nor_x1_sg U11342 ( .A(n1734), .B(n1735), .X(n1683) );
  nor_x1_sg U11343 ( .A(n1904), .B(n1905), .X(n1853) );
  nor_x1_sg U11344 ( .A(n1987), .B(n1988), .X(n1936) );
  nor_x1_sg U11345 ( .A(n2072), .B(n2073), .X(n2021) );
  nor_x1_sg U11346 ( .A(n1471), .B(n1470), .X(n733) );
  nor_x1_sg U11347 ( .A(n8902), .B(n1470), .X(\update_mask_0/n952 ) );
  inv_x1_sg U11348 ( .A(n1471), .X(n8902) );
  nor_x1_sg U11349 ( .A(n1773), .B(n8929), .X(n1772) );
  nor_x1_sg U11350 ( .A(n2111), .B(n8937), .X(n2110) );
  nor_x1_sg U11351 ( .A(n1617), .B(n1618), .X(n1614) );
  nor_x1_sg U11352 ( .A(n6325), .B(n1616), .X(n1615) );
  nor_x1_sg U11353 ( .A(n1955), .B(n1956), .X(n1952) );
  nor_x1_sg U11354 ( .A(n6118), .B(n1954), .X(n1953) );
  nor_x1_sg U11355 ( .A(n2209), .B(n2210), .X(n2205) );
  nor_x1_sg U11356 ( .A(n2207), .B(n2208), .X(n2206) );
  nor_x1_sg U11357 ( .A(n1532), .B(n1533), .X(n1528) );
  nor_x1_sg U11358 ( .A(n1530), .B(n1531), .X(n1529) );
  nor_x1_sg U11359 ( .A(n1702), .B(n1703), .X(n1698) );
  nor_x1_sg U11360 ( .A(n1700), .B(n1701), .X(n1699) );
  nor_x1_sg U11361 ( .A(n1800), .B(n1801), .X(n1796) );
  nor_x1_sg U11362 ( .A(n1798), .B(n1799), .X(n1797) );
  nor_x1_sg U11363 ( .A(n1872), .B(n1873), .X(n1868) );
  nor_x1_sg U11364 ( .A(n1870), .B(n1871), .X(n1869) );
  nor_x1_sg U11365 ( .A(n2040), .B(n2041), .X(n2036) );
  nor_x1_sg U11366 ( .A(n2038), .B(n2039), .X(n2037) );
  nor_x1_sg U11367 ( .A(n2138), .B(n2139), .X(n2134) );
  nor_x1_sg U11368 ( .A(n2136), .B(n2137), .X(n2135) );
  nor_x1_sg U11369 ( .A(n7459), .B(n6369), .X(n792) );
  nand_x1_sg U11370 ( .A(n7084), .B(n9148), .X(n1306) );
  inv_x2_sg U11371 ( .A(\i_im[12][6] ), .X(n9148) );
  nand_x1_sg U11372 ( .A(n6653), .B(n6550), .X(n3775) );
  nand_x1_sg U11373 ( .A(\o_im[6][17] ), .B(n6513), .X(n3776) );
  nand_x1_sg U11374 ( .A(n6645), .B(n6550), .X(n3771) );
  nand_x1_sg U11375 ( .A(\o_im[6][15] ), .B(n6321), .X(n3772) );
  nand_x1_sg U11376 ( .A(n6563), .B(n6551), .X(n3767) );
  nand_x1_sg U11377 ( .A(\o_im[6][13] ), .B(n7406), .X(n3768) );
  nand_x1_sg U11378 ( .A(n6567), .B(n6549), .X(n3763) );
  nand_x1_sg U11379 ( .A(\o_im[6][11] ), .B(n6511), .X(n3764) );
  nand_x1_sg U11380 ( .A(n6633), .B(n6552), .X(n3759) );
  nand_x1_sg U11381 ( .A(\o_im[6][9] ), .B(n6513), .X(n3760) );
  nand_x1_sg U11382 ( .A(n6625), .B(n6552), .X(n3755) );
  nand_x1_sg U11383 ( .A(\o_im[6][7] ), .B(n6512), .X(n3756) );
  nand_x1_sg U11384 ( .A(n6621), .B(n6549), .X(n3751) );
  nand_x1_sg U11385 ( .A(\o_im[6][5] ), .B(n7406), .X(n3752) );
  nand_x1_sg U11386 ( .A(n6576), .B(n6549), .X(n3747) );
  nand_x1_sg U11387 ( .A(\o_im[6][3] ), .B(n7406), .X(n3748) );
  nand_x1_sg U11388 ( .A(n6613), .B(n6550), .X(n3743) );
  nand_x1_sg U11389 ( .A(\o_im[6][1] ), .B(n6511), .X(n3744) );
  nand_x1_sg U11390 ( .A(n6654), .B(n6116), .X(n3689) );
  nand_x1_sg U11391 ( .A(\o_im[4][17] ), .B(n6837), .X(n3690) );
  nand_x1_sg U11392 ( .A(n6646), .B(n6993), .X(n3685) );
  nand_x1_sg U11393 ( .A(\o_im[4][15] ), .B(n6836), .X(n3686) );
  nand_x1_sg U11394 ( .A(n6564), .B(n6995), .X(n3681) );
  nand_x1_sg U11395 ( .A(\o_im[4][13] ), .B(n6835), .X(n3682) );
  nand_x1_sg U11396 ( .A(n6568), .B(n6993), .X(n3677) );
  nand_x1_sg U11397 ( .A(\o_im[4][11] ), .B(n5968), .X(n3678) );
  nand_x1_sg U11398 ( .A(n6634), .B(n6993), .X(n3673) );
  nand_x1_sg U11399 ( .A(\o_im[4][9] ), .B(n6835), .X(n3674) );
  nand_x1_sg U11400 ( .A(n6626), .B(n6995), .X(n3669) );
  nand_x1_sg U11401 ( .A(\o_im[4][7] ), .B(n6835), .X(n3670) );
  nand_x1_sg U11402 ( .A(n6622), .B(n6994), .X(n3665) );
  nand_x1_sg U11403 ( .A(\o_im[4][5] ), .B(n6836), .X(n3666) );
  nand_x1_sg U11404 ( .A(n6577), .B(n6995), .X(n3661) );
  nand_x1_sg U11405 ( .A(\o_im[4][3] ), .B(n6835), .X(n3662) );
  nand_x1_sg U11406 ( .A(n6614), .B(n6995), .X(n3657) );
  nand_x1_sg U11407 ( .A(\o_im[4][1] ), .B(n6837), .X(n3658) );
  nand_x1_sg U11408 ( .A(n6661), .B(n6336), .X(n3779) );
  nand_x1_sg U11409 ( .A(\o_im[6][19] ), .B(n6512), .X(n3780) );
  nand_x1_sg U11410 ( .A(n6657), .B(n6335), .X(n3777) );
  nand_x1_sg U11411 ( .A(\o_im[6][18] ), .B(n6513), .X(n3778) );
  nand_x1_sg U11412 ( .A(n6649), .B(n6335), .X(n3773) );
  nand_x1_sg U11413 ( .A(\o_im[6][16] ), .B(n6512), .X(n3774) );
  nand_x1_sg U11414 ( .A(n6561), .B(n6336), .X(n3769) );
  nand_x1_sg U11415 ( .A(\o_im[6][14] ), .B(n6321), .X(n3770) );
  nand_x1_sg U11416 ( .A(n6641), .B(n6551), .X(n3765) );
  nand_x1_sg U11417 ( .A(\o_im[6][12] ), .B(n6513), .X(n3766) );
  nand_x1_sg U11418 ( .A(n6637), .B(n6336), .X(n3761) );
  nand_x1_sg U11419 ( .A(\o_im[6][10] ), .B(n6511), .X(n3762) );
  nand_x1_sg U11420 ( .A(n6629), .B(n6550), .X(n3757) );
  nand_x1_sg U11421 ( .A(\o_im[6][8] ), .B(n7406), .X(n3758) );
  nand_x1_sg U11422 ( .A(n6573), .B(n6335), .X(n3753) );
  nand_x1_sg U11423 ( .A(\o_im[6][6] ), .B(n6321), .X(n3754) );
  nand_x1_sg U11424 ( .A(n6617), .B(n6552), .X(n3749) );
  nand_x1_sg U11425 ( .A(\o_im[6][4] ), .B(n6321), .X(n3750) );
  nand_x1_sg U11426 ( .A(n6580), .B(n6336), .X(n3745) );
  nand_x1_sg U11427 ( .A(\o_im[6][2] ), .B(n6511), .X(n3746) );
  nand_x1_sg U11428 ( .A(n6609), .B(n6551), .X(n3740) );
  nand_x1_sg U11429 ( .A(\o_im[6][0] ), .B(n6512), .X(n3741) );
  nand_x1_sg U11430 ( .A(n6660), .B(n6994), .X(n3693) );
  nand_x1_sg U11431 ( .A(\o_im[4][19] ), .B(n6834), .X(n3694) );
  nand_x1_sg U11432 ( .A(n6658), .B(n6992), .X(n3691) );
  nand_x1_sg U11433 ( .A(\o_im[4][18] ), .B(n5968), .X(n3692) );
  nand_x1_sg U11434 ( .A(n6650), .B(n6992), .X(n3687) );
  nand_x1_sg U11435 ( .A(\o_im[4][16] ), .B(n5968), .X(n3688) );
  nand_x1_sg U11436 ( .A(n6560), .B(n6992), .X(n3683) );
  nand_x1_sg U11437 ( .A(\o_im[4][14] ), .B(n6836), .X(n3684) );
  nand_x1_sg U11438 ( .A(n6642), .B(n6994), .X(n3679) );
  nand_x1_sg U11439 ( .A(\o_im[4][12] ), .B(n6834), .X(n3680) );
  nand_x1_sg U11440 ( .A(n6638), .B(n6994), .X(n3675) );
  nand_x1_sg U11441 ( .A(\o_im[4][10] ), .B(n6834), .X(n3676) );
  nand_x1_sg U11442 ( .A(n6630), .B(n6116), .X(n3671) );
  nand_x1_sg U11443 ( .A(\o_im[4][8] ), .B(n6837), .X(n3672) );
  nand_x1_sg U11444 ( .A(n6572), .B(n6116), .X(n3667) );
  nand_x1_sg U11445 ( .A(\o_im[4][6] ), .B(n5968), .X(n3668) );
  nand_x1_sg U11446 ( .A(n6618), .B(n6116), .X(n3663) );
  nand_x1_sg U11447 ( .A(\o_im[4][4] ), .B(n6834), .X(n3664) );
  nand_x1_sg U11448 ( .A(n6581), .B(n6993), .X(n3659) );
  nand_x1_sg U11449 ( .A(\o_im[4][2] ), .B(n6836), .X(n3660) );
  nand_x1_sg U11450 ( .A(n6610), .B(n6992), .X(n3654) );
  nand_x1_sg U11451 ( .A(\o_im[4][0] ), .B(n6837), .X(n3655) );
  nor_x1_sg U11452 ( .A(n7395), .B(\update_output_0/N29 ), .X(n1438) );
  nor_x1_sg U11453 ( .A(n7299), .B(\i_im[3][12] ), .X(n970) );
  nand_x1_sg U11454 ( .A(n6440), .B(n9028), .X(n1288) );
  inv_x2_sg U11455 ( .A(\i_im[4][6] ), .X(n9028) );
  nand_x1_sg U11456 ( .A(n7083), .B(n9152), .X(n1010) );
  inv_x2_sg U11457 ( .A(\i_im[12][10] ), .X(n9152) );
  nor_x1_sg U11458 ( .A(n7289), .B(\i_im[11][6] ), .X(n1313) );
  nor_x1_sg U11459 ( .A(n7290), .B(\i_im[3][6] ), .X(n1298) );
  nor_x1_sg U11460 ( .A(n7301), .B(\i_im[3][1] ), .X(n1135) );
  nor_x1_sg U11461 ( .A(n7289), .B(\i_im[3][5] ), .X(n1266) );
  nor_x1_sg U11462 ( .A(n7294), .B(\i_im[3][10] ), .X(n1002) );
  nor_x1_sg U11463 ( .A(n7298), .B(\i_im[3][15] ), .X(n807) );
  nand_x1_sg U11464 ( .A(n6439), .B(n9147), .X(n1274) );
  inv_x2_sg U11465 ( .A(\i_im[12][5] ), .X(n9147) );
  nand_x1_sg U11466 ( .A(n7145), .B(n9048), .X(n1297) );
  inv_x2_sg U11467 ( .A(\i_im[5][6] ), .X(n9048) );
  nor_x1_sg U11468 ( .A(n7293), .B(\i_im[11][5] ), .X(n1281) );
  nor_x1_sg U11469 ( .A(n7295), .B(\i_im[11][1] ), .X(n1150) );
  nor_x1_sg U11470 ( .A(n7295), .B(\i_im[11][12] ), .X(n985) );
  nor_x1_sg U11471 ( .A(n7300), .B(\i_im[11][15] ), .X(n822) );
  nor_x1_sg U11472 ( .A(n7291), .B(\i_im[3][2] ), .X(n1167) );
  nor_x1_sg U11473 ( .A(n7301), .B(\i_im[3][16] ), .X(n839) );
  nand_x1_sg U11474 ( .A(n7086), .B(n9032), .X(n992) );
  nor_x1_sg U11475 ( .A(n7071), .B(\i_im[1][10] ), .X(n993) );
  nor_x1_sg U11476 ( .A(n7291), .B(\i_im[11][10] ), .X(n1017) );
  nand_x1_sg U11477 ( .A(n7267), .B(n9187), .X(n1280) );
  inv_x2_sg U11478 ( .A(\i_im[14][5] ), .X(n9187) );
  nor_x1_sg U11479 ( .A(n7294), .B(\i_im[11][2] ), .X(n1182) );
  nor_x1_sg U11480 ( .A(n7296), .B(\i_im[11][16] ), .X(n854) );
  nand_x1_sg U11481 ( .A(n6171), .B(n9144), .X(n1175) );
  inv_x2_sg U11482 ( .A(\i_im[12][2] ), .X(n9144) );
  nand_x1_sg U11483 ( .A(n6170), .B(n9027), .X(n1256) );
  inv_x2_sg U11484 ( .A(\i_im[4][5] ), .X(n9027) );
  nor_x1_sg U11485 ( .A(n979), .B(n980), .X(n977) );
  nand_x1_sg U11486 ( .A(n7085), .B(n9154), .X(n978) );
  nor_x1_sg U11487 ( .A(\i_im[10][12] ), .B(n7238), .X(n980) );
  nand_x1_sg U11488 ( .A(n7260), .B(n9184), .X(n1181) );
  inv_x2_sg U11489 ( .A(\i_im[14][2] ), .X(n9184) );
  nand_x1_sg U11490 ( .A(n6007), .B(n9024), .X(n1157) );
  inv_x2_sg U11491 ( .A(\i_im[4][2] ), .X(n9024) );
  nand_x1_sg U11492 ( .A(n6171), .B(n9034), .X(n960) );
  inv_x2_sg U11493 ( .A(\i_im[4][12] ), .X(n9034) );
  nor_x1_sg U11494 ( .A(n848), .B(n849), .X(n846) );
  nand_x1_sg U11495 ( .A(n7086), .B(n9158), .X(n847) );
  nor_x1_sg U11496 ( .A(\i_im[10][16] ), .B(n7238), .X(n849) );
  nand_x1_sg U11497 ( .A(n7083), .B(n9023), .X(n1125) );
  inv_x2_sg U11498 ( .A(\i_im[4][1] ), .X(n9023) );
  nand_x1_sg U11499 ( .A(n7084), .B(n9038), .X(n829) );
  inv_x2_sg U11500 ( .A(\i_im[4][16] ), .X(n9038) );
  nor_x1_sg U11501 ( .A(n816), .B(n817), .X(n814) );
  nand_x1_sg U11502 ( .A(n7085), .B(n9157), .X(n815) );
  nor_x1_sg U11503 ( .A(\i_im[10][15] ), .B(n7238), .X(n817) );
  nand_x1_sg U11504 ( .A(n6170), .B(n9037), .X(n791) );
  inv_x2_sg U11505 ( .A(\i_im[4][15] ), .X(n9037) );
  nor_x1_sg U11506 ( .A(\update_output_0/N28 ), .B(\update_output_0/N29 ), .X(
        n1433) );
  nor_x1_sg U11507 ( .A(\i_im[8][12] ), .B(n7152), .X(n979) );
  nor_x1_sg U11508 ( .A(\i_im[8][15] ), .B(n7157), .X(n816) );
  nor_x1_sg U11509 ( .A(n1275), .B(n1276), .X(n1273) );
  nor_x1_sg U11510 ( .A(\i_im[10][5] ), .B(n7229), .X(n1276) );
  nor_x1_sg U11511 ( .A(\i_im[8][5] ), .B(n7159), .X(n1275) );
  nor_x1_sg U11512 ( .A(n1011), .B(n1012), .X(n1009) );
  nor_x1_sg U11513 ( .A(\i_im[10][10] ), .B(n7232), .X(n1012) );
  nor_x1_sg U11514 ( .A(\i_im[8][10] ), .B(n7155), .X(n1011) );
  nor_x1_sg U11515 ( .A(\i_im[8][16] ), .B(n7156), .X(n848) );
  nor_x1_sg U11516 ( .A(n1176), .B(n1177), .X(n1174) );
  nor_x1_sg U11517 ( .A(\i_im[10][2] ), .B(n7230), .X(n1177) );
  nor_x1_sg U11518 ( .A(\i_im[8][2] ), .B(n7150), .X(n1176) );
  nor_x1_sg U11519 ( .A(n1307), .B(n1308), .X(n1305) );
  nor_x1_sg U11520 ( .A(\i_im[10][6] ), .B(n7236), .X(n1308) );
  nor_x1_sg U11521 ( .A(\i_im[8][6] ), .B(n7157), .X(n1307) );
  nor_x1_sg U11522 ( .A(n7078), .B(\i_im[1][5] ), .X(n1257) );
  nor_x1_sg U11523 ( .A(n7077), .B(\i_im[1][12] ), .X(n961) );
  nor_x1_sg U11524 ( .A(\i_im[10][1] ), .B(n7236), .X(n1145) );
  nand_x1_sg U11525 ( .A(n6008), .B(n9143), .X(n1143) );
  nor_x1_sg U11526 ( .A(n1144), .B(n1145), .X(n1142) );
  inv_x2_sg U11527 ( .A(\i_im[12][1] ), .X(n9143) );
  nor_x1_sg U11528 ( .A(n6457), .B(n7395), .X(n1442) );
  nor_x1_sg U11529 ( .A(n7070), .B(\i_im[1][1] ), .X(n1126) );
  nor_x1_sg U11530 ( .A(n7075), .B(\i_im[1][6] ), .X(n1289) );
  nor_x1_sg U11531 ( .A(n7081), .B(\i_im[1][15] ), .X(n793) );
  nor_x1_sg U11532 ( .A(n7081), .B(\i_im[1][16] ), .X(n830) );
  nor_x1_sg U11533 ( .A(n7322), .B(n964), .X(n962) );
  nor_x1_sg U11534 ( .A(\i_im[0][12] ), .B(n7159), .X(n964) );
  nand_x1_sg U11535 ( .A(n6490), .B(n9208), .X(n1311) );
  inv_x2_sg U11536 ( .A(\i_im[15][6] ), .X(n9208) );
  nor_x1_sg U11537 ( .A(n7231), .B(\i_im[2][6] ), .X(n1291) );
  nor_x1_sg U11538 ( .A(n7077), .B(\i_im[9][12] ), .X(n976) );
  nor_x1_sg U11539 ( .A(n7078), .B(\i_im[1][2] ), .X(n1158) );
  nor_x1_sg U11540 ( .A(\i_im[0][10] ), .B(n7153), .X(n996) );
  nor_x1_sg U11541 ( .A(n6361), .B(n1129), .X(n1127) );
  nor_x1_sg U11542 ( .A(\i_im[0][1] ), .B(n7150), .X(n1129) );
  nor_x1_sg U11543 ( .A(n7321), .B(n1260), .X(n1258) );
  nor_x1_sg U11544 ( .A(\i_im[0][5] ), .B(n7160), .X(n1260) );
  nor_x1_sg U11545 ( .A(n6082), .B(n798), .X(n795) );
  nor_x1_sg U11546 ( .A(\i_im[0][15] ), .B(n7161), .X(n798) );
  nor_x1_sg U11547 ( .A(n7320), .B(n996), .X(n994) );
  nor_x1_sg U11548 ( .A(n7231), .B(\i_im[2][10] ), .X(n995) );
  nand_x1_sg U11549 ( .A(n7262), .B(n9068), .X(n1296) );
  nand_x1_sg U11550 ( .A(n6390), .B(n9088), .X(n1295) );
  inv_x2_sg U11551 ( .A(\i_im[6][6] ), .X(n9068) );
  nor_x1_sg U11552 ( .A(n7070), .B(\i_im[9][1] ), .X(n1141) );
  nor_x1_sg U11553 ( .A(n7081), .B(\i_im[9][15] ), .X(n813) );
  nor_x1_sg U11554 ( .A(n7076), .B(\i_im[9][5] ), .X(n1272) );
  nor_x1_sg U11555 ( .A(n7073), .B(\i_im[9][6] ), .X(n1304) );
  nor_x1_sg U11556 ( .A(n7072), .B(\i_im[9][10] ), .X(n1008) );
  nor_x1_sg U11557 ( .A(\i_im[8][1] ), .B(n7160), .X(n1144) );
  nor_x1_sg U11558 ( .A(\i_im[0][6] ), .B(n7153), .X(n1292) );
  nor_x1_sg U11559 ( .A(n6362), .B(n1161), .X(n1159) );
  nor_x1_sg U11560 ( .A(\i_im[0][2] ), .B(n7151), .X(n1161) );
  nor_x1_sg U11561 ( .A(n6083), .B(n833), .X(n831) );
  nor_x1_sg U11562 ( .A(\i_im[0][16] ), .B(n7162), .X(n833) );
  nand_x1_sg U11563 ( .A(n6035), .B(n9163), .X(n1140) );
  inv_x2_sg U11564 ( .A(\i_im[13][1] ), .X(n9163) );
  nand_x1_sg U11565 ( .A(n7144), .B(n9177), .X(n812) );
  inv_x2_sg U11566 ( .A(\i_im[13][15] ), .X(n9177) );
  nor_x1_sg U11567 ( .A(n7080), .B(\i_im[9][16] ), .X(n845) );
  nor_x1_sg U11568 ( .A(n7070), .B(\i_im[9][2] ), .X(n1173) );
  nor_x1_sg U11569 ( .A(n7234), .B(\i_im[2][5] ), .X(n1259) );
  nand_x1_sg U11570 ( .A(n6389), .B(n9207), .X(n1279) );
  inv_x2_sg U11571 ( .A(\i_im[15][5] ), .X(n9207) );
  nand_x1_sg U11572 ( .A(n6421), .B(n9178), .X(n844) );
  inv_x2_sg U11573 ( .A(\i_im[13][16] ), .X(n9178) );
  nor_x1_sg U11574 ( .A(n7232), .B(\i_im[2][12] ), .X(n963) );
  nand_x1_sg U11575 ( .A(n6128), .B(n9087), .X(n1263) );
  inv_x2_sg U11576 ( .A(\i_im[7][5] ), .X(n9087) );
  nand_x1_sg U11577 ( .A(n7279), .B(n9092), .X(n999) );
  inv_x2_sg U11578 ( .A(\i_im[7][10] ), .X(n9092) );
  nor_x1_sg U11579 ( .A(n7239), .B(\i_im[2][1] ), .X(n1128) );
  nor_x1_sg U11580 ( .A(n7229), .B(\i_im[2][2] ), .X(n1160) );
  nor_x1_sg U11581 ( .A(n7240), .B(\i_im[2][15] ), .X(n796) );
  nand_x1_sg U11582 ( .A(n7319), .B(n1180), .X(n1179) );
  nand_x1_sg U11583 ( .A(n6492), .B(n9204), .X(n1180) );
  inv_x2_sg U11584 ( .A(\i_im[15][2] ), .X(n9204) );
  nor_x1_sg U11585 ( .A(n7235), .B(\i_im[2][16] ), .X(n832) );
  nand_x1_sg U11586 ( .A(n6389), .B(n9084), .X(n1164) );
  inv_x2_sg U11587 ( .A(\i_im[7][2] ), .X(n9084) );
  nand_x1_sg U11588 ( .A(n6491), .B(n9094), .X(n967) );
  inv_x2_sg U11589 ( .A(\i_im[7][12] ), .X(n9094) );
  nand_x1_sg U11590 ( .A(n6007), .B(n9151), .X(n1402) );
  inv_x2_sg U11591 ( .A(\i_im[12][9] ), .X(n9151) );
  nand_x1_sg U11592 ( .A(n7279), .B(n9098), .X(n836) );
  inv_x2_sg U11593 ( .A(\i_im[7][16] ), .X(n9098) );
  nand_x1_sg U11594 ( .A(n7281), .B(n9083), .X(n1132) );
  inv_x2_sg U11595 ( .A(\i_im[7][1] ), .X(n9083) );
  nand_x1_sg U11596 ( .A(n6422), .B(n9047), .X(n1265) );
  inv_x2_sg U11597 ( .A(\i_im[5][5] ), .X(n9047) );
  nand_x1_sg U11598 ( .A(n7083), .B(n9149), .X(n1338) );
  inv_x2_sg U11599 ( .A(\i_im[12][7] ), .X(n9149) );
  nand_x1_sg U11600 ( .A(n6439), .B(n9031), .X(n1384) );
  inv_x2_sg U11601 ( .A(\i_im[4][9] ), .X(n9031) );
  nor_x1_sg U11602 ( .A(n7290), .B(\i_im[11][9] ), .X(n1409) );
  nand_x1_sg U11603 ( .A(n7280), .B(n9097), .X(n802) );
  inv_x2_sg U11604 ( .A(\i_im[7][15] ), .X(n9097) );
  nand_x1_sg U11605 ( .A(n6324), .B(n9044), .X(n1166) );
  inv_x2_sg U11606 ( .A(\i_im[5][2] ), .X(n9044) );
  nor_x1_sg U11607 ( .A(n7294), .B(\i_im[3][9] ), .X(n1394) );
  nand_x1_sg U11608 ( .A(n7084), .B(n9029), .X(n1320) );
  inv_x2_sg U11609 ( .A(\i_im[4][7] ), .X(n9029) );
  nand_x1_sg U11610 ( .A(n7086), .B(n9145), .X(n1239) );
  inv_x2_sg U11611 ( .A(\i_im[12][3] ), .X(n9145) );
  nand_x1_sg U11612 ( .A(n7086), .B(n9153), .X(n1042) );
  inv_x2_sg U11613 ( .A(\i_im[12][11] ), .X(n9153) );
  nand_x1_sg U11614 ( .A(n7145), .B(n9051), .X(n1393) );
  inv_x2_sg U11615 ( .A(\i_im[5][9] ), .X(n9051) );
  nor_x1_sg U11616 ( .A(n7293), .B(\i_im[11][7] ), .X(n1345) );
  nor_x1_sg U11617 ( .A(n7289), .B(\i_im[11][14] ), .X(n1113) );
  nand_x1_sg U11618 ( .A(n6654), .B(n6954), .X(n3732) );
  nand_x1_sg U11619 ( .A(\o_im[5][17] ), .B(n6876), .X(n3733) );
  nand_x1_sg U11620 ( .A(n6643), .B(n6954), .X(n3728) );
  nand_x1_sg U11621 ( .A(\o_im[5][15] ), .B(n5976), .X(n3729) );
  nand_x1_sg U11622 ( .A(n6563), .B(n6954), .X(n3724) );
  nand_x1_sg U11623 ( .A(\o_im[5][13] ), .B(n5976), .X(n3725) );
  nand_x1_sg U11624 ( .A(n6569), .B(n6955), .X(n3720) );
  nand_x1_sg U11625 ( .A(\o_im[5][11] ), .B(n6874), .X(n3721) );
  nand_x1_sg U11626 ( .A(n6631), .B(n6953), .X(n3716) );
  nand_x1_sg U11627 ( .A(\o_im[5][9] ), .B(n6877), .X(n3717) );
  nand_x1_sg U11628 ( .A(n6624), .B(n6108), .X(n3712) );
  nand_x1_sg U11629 ( .A(\o_im[5][7] ), .B(n5976), .X(n3713) );
  nand_x1_sg U11630 ( .A(n6621), .B(n6953), .X(n3708) );
  nand_x1_sg U11631 ( .A(\o_im[5][5] ), .B(n6875), .X(n3709) );
  nand_x1_sg U11632 ( .A(n6574), .B(n6108), .X(n3704) );
  nand_x1_sg U11633 ( .A(\o_im[5][3] ), .B(n6874), .X(n3705) );
  nand_x1_sg U11634 ( .A(n6613), .B(n6952), .X(n3700) );
  nand_x1_sg U11635 ( .A(\o_im[5][1] ), .B(n6875), .X(n3701) );
  nand_x1_sg U11636 ( .A(n6651), .B(n6983), .X(n3516) );
  nand_x1_sg U11637 ( .A(\o_im[0][17] ), .B(n6891), .X(n3517) );
  nand_x1_sg U11638 ( .A(n6646), .B(n6982), .X(n3512) );
  nand_x1_sg U11639 ( .A(\o_im[0][15] ), .B(n6889), .X(n3513) );
  nand_x1_sg U11640 ( .A(n6563), .B(n6982), .X(n3508) );
  nand_x1_sg U11641 ( .A(\o_im[0][13] ), .B(n6891), .X(n3509) );
  nand_x1_sg U11642 ( .A(n6568), .B(n6983), .X(n3504) );
  nand_x1_sg U11643 ( .A(\o_im[0][11] ), .B(n5979), .X(n3505) );
  nand_x1_sg U11644 ( .A(n6633), .B(n6985), .X(n3500) );
  nand_x1_sg U11645 ( .A(\o_im[0][9] ), .B(n6892), .X(n3501) );
  nand_x1_sg U11646 ( .A(n6626), .B(n6114), .X(n3496) );
  nand_x1_sg U11647 ( .A(\o_im[0][7] ), .B(n6891), .X(n3497) );
  nand_x1_sg U11648 ( .A(n6622), .B(n6985), .X(n3492) );
  nand_x1_sg U11649 ( .A(\o_im[0][5] ), .B(n6890), .X(n3493) );
  nand_x1_sg U11650 ( .A(n6577), .B(n6114), .X(n3488) );
  nand_x1_sg U11651 ( .A(\o_im[0][3] ), .B(n6889), .X(n3489) );
  nand_x1_sg U11652 ( .A(n6614), .B(n6982), .X(n3484) );
  nand_x1_sg U11653 ( .A(\o_im[0][1] ), .B(n5979), .X(n3485) );
  nand_x1_sg U11654 ( .A(n6651), .B(n6969), .X(n3646) );
  nand_x1_sg U11655 ( .A(\o_im[3][17] ), .B(n6900), .X(n3647) );
  nand_x1_sg U11656 ( .A(n6643), .B(n6967), .X(n3642) );
  nand_x1_sg U11657 ( .A(\o_im[3][15] ), .B(n6898), .X(n3643) );
  nand_x1_sg U11658 ( .A(n6563), .B(n6968), .X(n3638) );
  nand_x1_sg U11659 ( .A(\o_im[3][13] ), .B(n6898), .X(n3639) );
  nand_x1_sg U11660 ( .A(n6567), .B(n6967), .X(n3634) );
  nand_x1_sg U11661 ( .A(\o_im[3][11] ), .B(n6900), .X(n3635) );
  nand_x1_sg U11662 ( .A(n6633), .B(n6968), .X(n3630) );
  nand_x1_sg U11663 ( .A(\o_im[3][9] ), .B(n6901), .X(n3631) );
  nand_x1_sg U11664 ( .A(n6624), .B(n6111), .X(n3626) );
  nand_x1_sg U11665 ( .A(\o_im[3][7] ), .B(n6899), .X(n3627) );
  nand_x1_sg U11666 ( .A(n6620), .B(n6969), .X(n3622) );
  nand_x1_sg U11667 ( .A(\o_im[3][5] ), .B(n6899), .X(n3623) );
  nand_x1_sg U11668 ( .A(n6576), .B(n6968), .X(n3618) );
  nand_x1_sg U11669 ( .A(\o_im[3][3] ), .B(n5981), .X(n3619) );
  nand_x1_sg U11670 ( .A(n6611), .B(n6111), .X(n3614) );
  nand_x1_sg U11671 ( .A(\o_im[3][1] ), .B(n6899), .X(n3615) );
  nand_x1_sg U11672 ( .A(n6651), .B(n6939), .X(n3819) );
  nand_x1_sg U11673 ( .A(\o_im[7][17] ), .B(n6871), .X(n3820) );
  nand_x1_sg U11674 ( .A(n6645), .B(n6105), .X(n3815) );
  nand_x1_sg U11675 ( .A(\o_im[7][15] ), .B(n6869), .X(n3816) );
  nand_x1_sg U11676 ( .A(n6565), .B(n6937), .X(n3811) );
  nand_x1_sg U11677 ( .A(\o_im[7][13] ), .B(n6869), .X(n3812) );
  nand_x1_sg U11678 ( .A(n6566), .B(n6937), .X(n3807) );
  nand_x1_sg U11679 ( .A(\o_im[7][11] ), .B(n5975), .X(n3808) );
  nand_x1_sg U11680 ( .A(n6634), .B(n6937), .X(n3803) );
  nand_x1_sg U11681 ( .A(\o_im[7][9] ), .B(n6872), .X(n3804) );
  nand_x1_sg U11682 ( .A(n6623), .B(n6940), .X(n3799) );
  nand_x1_sg U11683 ( .A(\o_im[7][7] ), .B(n6871), .X(n3800) );
  nand_x1_sg U11684 ( .A(n6619), .B(n6940), .X(n3795) );
  nand_x1_sg U11685 ( .A(\o_im[7][5] ), .B(n6871), .X(n3796) );
  nand_x1_sg U11686 ( .A(n6575), .B(n6938), .X(n3791) );
  nand_x1_sg U11687 ( .A(\o_im[7][3] ), .B(n5975), .X(n3792) );
  nand_x1_sg U11688 ( .A(n6611), .B(n6105), .X(n3787) );
  nand_x1_sg U11689 ( .A(\o_im[7][1] ), .B(n6870), .X(n3788) );
  nand_x1_sg U11690 ( .A(n6654), .B(n6975), .X(n3560) );
  nand_x1_sg U11691 ( .A(\o_im[1][17] ), .B(n6846), .X(n3561) );
  nand_x1_sg U11692 ( .A(n6644), .B(n6972), .X(n3556) );
  nand_x1_sg U11693 ( .A(\o_im[1][15] ), .B(n5970), .X(n3557) );
  nand_x1_sg U11694 ( .A(n6562), .B(n6974), .X(n3552) );
  nand_x1_sg U11695 ( .A(\o_im[1][13] ), .B(n5970), .X(n3553) );
  nand_x1_sg U11696 ( .A(n6566), .B(n6975), .X(n3548) );
  nand_x1_sg U11697 ( .A(\o_im[1][11] ), .B(n6844), .X(n3549) );
  nand_x1_sg U11698 ( .A(n6633), .B(n6974), .X(n3544) );
  nand_x1_sg U11699 ( .A(\o_im[1][9] ), .B(n6847), .X(n3545) );
  nand_x1_sg U11700 ( .A(n6623), .B(n6975), .X(n3540) );
  nand_x1_sg U11701 ( .A(\o_im[1][7] ), .B(n5970), .X(n3541) );
  nand_x1_sg U11702 ( .A(n6621), .B(n6972), .X(n3536) );
  nand_x1_sg U11703 ( .A(\o_im[1][5] ), .B(n6845), .X(n3537) );
  nand_x1_sg U11704 ( .A(n6575), .B(n6972), .X(n3532) );
  nand_x1_sg U11705 ( .A(\o_im[1][3] ), .B(n6846), .X(n3533) );
  nand_x1_sg U11706 ( .A(n6613), .B(n6112), .X(n3528) );
  nand_x1_sg U11707 ( .A(\o_im[1][1] ), .B(n6846), .X(n3529) );
  nand_x1_sg U11708 ( .A(n6662), .B(n6983), .X(n3520) );
  nand_x1_sg U11709 ( .A(\o_im[0][19] ), .B(n6891), .X(n3521) );
  nand_x1_sg U11710 ( .A(n6658), .B(n6984), .X(n3518) );
  nand_x1_sg U11711 ( .A(\o_im[0][18] ), .B(n6890), .X(n3519) );
  nand_x1_sg U11712 ( .A(n6649), .B(n6982), .X(n3514) );
  nand_x1_sg U11713 ( .A(\o_im[0][16] ), .B(n6892), .X(n3515) );
  nand_x1_sg U11714 ( .A(n6558), .B(n6984), .X(n3510) );
  nand_x1_sg U11715 ( .A(\o_im[0][14] ), .B(n6892), .X(n3511) );
  nand_x1_sg U11716 ( .A(n6641), .B(n6114), .X(n3506) );
  nand_x1_sg U11717 ( .A(\o_im[0][12] ), .B(n5979), .X(n3507) );
  nand_x1_sg U11718 ( .A(n6636), .B(n6985), .X(n3502) );
  nand_x1_sg U11719 ( .A(\o_im[0][10] ), .B(n6889), .X(n3503) );
  nand_x1_sg U11720 ( .A(n6627), .B(n6984), .X(n3498) );
  nand_x1_sg U11721 ( .A(\o_im[0][8] ), .B(n5979), .X(n3499) );
  nand_x1_sg U11722 ( .A(n6571), .B(n6983), .X(n3494) );
  nand_x1_sg U11723 ( .A(\o_im[0][6] ), .B(n6890), .X(n3495) );
  nand_x1_sg U11724 ( .A(n6615), .B(n6985), .X(n3490) );
  nand_x1_sg U11725 ( .A(\o_im[0][4] ), .B(n6890), .X(n3491) );
  nand_x1_sg U11726 ( .A(n6580), .B(n6114), .X(n3486) );
  nand_x1_sg U11727 ( .A(\o_im[0][2] ), .B(n6892), .X(n3487) );
  nand_x1_sg U11728 ( .A(n6610), .B(n6984), .X(n3481) );
  nand_x1_sg U11729 ( .A(\o_im[0][0] ), .B(n6889), .X(n3482) );
  nand_x1_sg U11730 ( .A(n6661), .B(n6967), .X(n3650) );
  nand_x1_sg U11731 ( .A(\o_im[3][19] ), .B(n5981), .X(n3651) );
  nand_x1_sg U11732 ( .A(n6657), .B(n6970), .X(n3648) );
  nand_x1_sg U11733 ( .A(\o_im[3][18] ), .B(n6901), .X(n3649) );
  nand_x1_sg U11734 ( .A(n6647), .B(n6967), .X(n3644) );
  nand_x1_sg U11735 ( .A(\o_im[3][16] ), .B(n6900), .X(n3645) );
  nand_x1_sg U11736 ( .A(n6559), .B(n6970), .X(n3640) );
  nand_x1_sg U11737 ( .A(\o_im[3][14] ), .B(n6898), .X(n3641) );
  nand_x1_sg U11738 ( .A(n6639), .B(n6968), .X(n3636) );
  nand_x1_sg U11739 ( .A(\o_im[3][12] ), .B(n5981), .X(n3637) );
  nand_x1_sg U11740 ( .A(n6638), .B(n6969), .X(n3632) );
  nand_x1_sg U11741 ( .A(\o_im[3][10] ), .B(n6900), .X(n3633) );
  nand_x1_sg U11742 ( .A(n6628), .B(n6970), .X(n3628) );
  nand_x1_sg U11743 ( .A(\o_im[3][8] ), .B(n6898), .X(n3629) );
  nand_x1_sg U11744 ( .A(n6570), .B(n6111), .X(n3624) );
  nand_x1_sg U11745 ( .A(\o_im[3][6] ), .B(n6899), .X(n3625) );
  nand_x1_sg U11746 ( .A(n6616), .B(n6970), .X(n3620) );
  nand_x1_sg U11747 ( .A(\o_im[3][4] ), .B(n5981), .X(n3621) );
  nand_x1_sg U11748 ( .A(n6581), .B(n6111), .X(n3616) );
  nand_x1_sg U11749 ( .A(\o_im[3][2] ), .B(n6901), .X(n3617) );
  nand_x1_sg U11750 ( .A(n6607), .B(n6969), .X(n3611) );
  nand_x1_sg U11751 ( .A(\o_im[3][0] ), .B(n6901), .X(n3612) );
  nand_x1_sg U11752 ( .A(n6661), .B(n6938), .X(n3823) );
  nand_x1_sg U11753 ( .A(\o_im[7][19] ), .B(n5975), .X(n3824) );
  nand_x1_sg U11754 ( .A(n6658), .B(n6940), .X(n3821) );
  nand_x1_sg U11755 ( .A(\o_im[7][18] ), .B(n6872), .X(n3822) );
  nand_x1_sg U11756 ( .A(n6650), .B(n6937), .X(n3817) );
  nand_x1_sg U11757 ( .A(\o_im[7][16] ), .B(n6872), .X(n3818) );
  nand_x1_sg U11758 ( .A(n6560), .B(n6939), .X(n3813) );
  nand_x1_sg U11759 ( .A(\o_im[7][14] ), .B(n6871), .X(n3814) );
  nand_x1_sg U11760 ( .A(n6641), .B(n6938), .X(n3809) );
  nand_x1_sg U11761 ( .A(\o_im[7][12] ), .B(n6869), .X(n3810) );
  nand_x1_sg U11762 ( .A(n6638), .B(n6105), .X(n3805) );
  nand_x1_sg U11763 ( .A(\o_im[7][10] ), .B(n5975), .X(n3806) );
  nand_x1_sg U11764 ( .A(n6628), .B(n6939), .X(n3801) );
  nand_x1_sg U11765 ( .A(\o_im[7][8] ), .B(n6870), .X(n3802) );
  nand_x1_sg U11766 ( .A(n6572), .B(n6939), .X(n3797) );
  nand_x1_sg U11767 ( .A(\o_im[7][6] ), .B(n6870), .X(n3798) );
  nand_x1_sg U11768 ( .A(n6617), .B(n6105), .X(n3793) );
  nand_x1_sg U11769 ( .A(\o_im[7][4] ), .B(n6870), .X(n3794) );
  nand_x1_sg U11770 ( .A(n6578), .B(n6938), .X(n3789) );
  nand_x1_sg U11771 ( .A(\o_im[7][2] ), .B(n6872), .X(n3790) );
  nand_x1_sg U11772 ( .A(n6609), .B(n6940), .X(n3784) );
  nand_x1_sg U11773 ( .A(\o_im[7][0] ), .B(n6869), .X(n3785) );
  nand_x1_sg U11774 ( .A(n6659), .B(n6975), .X(n3564) );
  nand_x1_sg U11775 ( .A(\o_im[1][19] ), .B(n6844), .X(n3565) );
  nand_x1_sg U11776 ( .A(n6658), .B(n6112), .X(n3562) );
  nand_x1_sg U11777 ( .A(\o_im[1][18] ), .B(n6847), .X(n3563) );
  nand_x1_sg U11778 ( .A(n6650), .B(n6973), .X(n3558) );
  nand_x1_sg U11779 ( .A(\o_im[1][16] ), .B(n6845), .X(n3559) );
  nand_x1_sg U11780 ( .A(n6559), .B(n6974), .X(n3554) );
  nand_x1_sg U11781 ( .A(\o_im[1][14] ), .B(n6847), .X(n3555) );
  nand_x1_sg U11782 ( .A(n6642), .B(n6974), .X(n3550) );
  nand_x1_sg U11783 ( .A(\o_im[1][12] ), .B(n6845), .X(n3551) );
  nand_x1_sg U11784 ( .A(n6635), .B(n6112), .X(n3546) );
  nand_x1_sg U11785 ( .A(\o_im[1][10] ), .B(n6844), .X(n3547) );
  nand_x1_sg U11786 ( .A(n6627), .B(n6112), .X(n3542) );
  nand_x1_sg U11787 ( .A(\o_im[1][8] ), .B(n5970), .X(n3543) );
  nand_x1_sg U11788 ( .A(n6573), .B(n6973), .X(n3538) );
  nand_x1_sg U11789 ( .A(\o_im[1][6] ), .B(n6845), .X(n3539) );
  nand_x1_sg U11790 ( .A(n6616), .B(n6972), .X(n3534) );
  nand_x1_sg U11791 ( .A(\o_im[1][4] ), .B(n6846), .X(n3535) );
  nand_x1_sg U11792 ( .A(n6581), .B(n6973), .X(n3530) );
  nand_x1_sg U11793 ( .A(\o_im[1][2] ), .B(n6844), .X(n3531) );
  nand_x1_sg U11794 ( .A(n6608), .B(n6973), .X(n3525) );
  nand_x1_sg U11795 ( .A(\o_im[1][0] ), .B(n6847), .X(n3526) );
  nand_x1_sg U11796 ( .A(n6659), .B(n6953), .X(n3736) );
  nand_x1_sg U11797 ( .A(\o_im[5][19] ), .B(n6876), .X(n3737) );
  nand_x1_sg U11798 ( .A(n6655), .B(n6955), .X(n3734) );
  nand_x1_sg U11799 ( .A(\o_im[5][18] ), .B(n6876), .X(n3735) );
  nand_x1_sg U11800 ( .A(n6648), .B(n6955), .X(n3730) );
  nand_x1_sg U11801 ( .A(\o_im[5][16] ), .B(n6877), .X(n3731) );
  nand_x1_sg U11802 ( .A(n6561), .B(n6108), .X(n3726) );
  nand_x1_sg U11803 ( .A(\o_im[5][14] ), .B(n6874), .X(n3727) );
  nand_x1_sg U11804 ( .A(n6639), .B(n6955), .X(n3722) );
  nand_x1_sg U11805 ( .A(\o_im[5][12] ), .B(n6874), .X(n3723) );
  nand_x1_sg U11806 ( .A(n6636), .B(n6953), .X(n3718) );
  nand_x1_sg U11807 ( .A(\o_im[5][10] ), .B(n5976), .X(n3719) );
  nand_x1_sg U11808 ( .A(n6630), .B(n6952), .X(n3714) );
  nand_x1_sg U11809 ( .A(\o_im[5][8] ), .B(n6875), .X(n3715) );
  nand_x1_sg U11810 ( .A(n6570), .B(n6108), .X(n3710) );
  nand_x1_sg U11811 ( .A(\o_im[5][6] ), .B(n6875), .X(n3711) );
  nand_x1_sg U11812 ( .A(n6618), .B(n6952), .X(n3706) );
  nand_x1_sg U11813 ( .A(\o_im[5][4] ), .B(n6876), .X(n3707) );
  nand_x1_sg U11814 ( .A(n6578), .B(n6952), .X(n3702) );
  nand_x1_sg U11815 ( .A(\o_im[5][2] ), .B(n6877), .X(n3703) );
  nand_x1_sg U11816 ( .A(n6609), .B(n6954), .X(n3697) );
  nand_x1_sg U11817 ( .A(\o_im[5][0] ), .B(n6877), .X(n3698) );
  nand_x1_sg U11818 ( .A(n6457), .B(\update_output_0/N28 ), .X(n1445) );
  nand_x1_sg U11819 ( .A(n7083), .B(n9150), .X(n1370) );
  inv_x2_sg U11820 ( .A(\i_im[12][8] ), .X(n9150) );
  nand_x1_sg U11821 ( .A(n6659), .B(n6933), .X(n3608) );
  nand_x1_sg U11822 ( .A(\o_im[2][19] ), .B(n6886), .X(n3607) );
  nand_x1_sg U11823 ( .A(n6656), .B(n6934), .X(n3606) );
  nand_x1_sg U11824 ( .A(\o_im[2][18] ), .B(n6887), .X(n3605) );
  nand_x1_sg U11825 ( .A(n6652), .B(n6935), .X(n3604) );
  nand_x1_sg U11826 ( .A(\o_im[2][17] ), .B(n6887), .X(n3603) );
  nand_x1_sg U11827 ( .A(n6647), .B(n6932), .X(n3602) );
  nand_x1_sg U11828 ( .A(\o_im[2][16] ), .B(n6887), .X(n3601) );
  nand_x1_sg U11829 ( .A(n6644), .B(n6933), .X(n3600) );
  nand_x1_sg U11830 ( .A(\o_im[2][15] ), .B(n6886), .X(n3599) );
  nand_x1_sg U11831 ( .A(n6559), .B(n6933), .X(n3598) );
  nand_x1_sg U11832 ( .A(\o_im[2][14] ), .B(n6887), .X(n3597) );
  nand_x1_sg U11833 ( .A(n6562), .B(n6104), .X(n3596) );
  nand_x1_sg U11834 ( .A(\o_im[2][13] ), .B(n5978), .X(n3595) );
  nand_x1_sg U11835 ( .A(n6640), .B(n6933), .X(n3594) );
  nand_x1_sg U11836 ( .A(\o_im[2][12] ), .B(n6884), .X(n3593) );
  nand_x1_sg U11837 ( .A(n6566), .B(n6932), .X(n3592) );
  nand_x1_sg U11838 ( .A(\o_im[2][11] ), .B(n6885), .X(n3591) );
  nand_x1_sg U11839 ( .A(n6636), .B(n6104), .X(n3590) );
  nand_x1_sg U11840 ( .A(\o_im[2][10] ), .B(n6885), .X(n3589) );
  nand_x1_sg U11841 ( .A(n6631), .B(n6935), .X(n3588) );
  nand_x1_sg U11842 ( .A(\o_im[2][9] ), .B(n6886), .X(n3587) );
  nand_x1_sg U11843 ( .A(n6628), .B(n6104), .X(n3586) );
  nand_x1_sg U11844 ( .A(\o_im[2][8] ), .B(n5978), .X(n3585) );
  nand_x1_sg U11845 ( .A(n6624), .B(n6935), .X(n3584) );
  nand_x1_sg U11846 ( .A(\o_im[2][7] ), .B(n5978), .X(n3583) );
  nand_x1_sg U11847 ( .A(n6571), .B(n6932), .X(n3582) );
  nand_x1_sg U11848 ( .A(\o_im[2][6] ), .B(n6884), .X(n3581) );
  nand_x1_sg U11849 ( .A(n6620), .B(n6934), .X(n3580) );
  nand_x1_sg U11850 ( .A(\o_im[2][5] ), .B(n5978), .X(n3579) );
  nand_x1_sg U11851 ( .A(n6615), .B(n6932), .X(n3578) );
  nand_x1_sg U11852 ( .A(\o_im[2][4] ), .B(n6884), .X(n3577) );
  nand_x1_sg U11853 ( .A(n6575), .B(n6934), .X(n3576) );
  nand_x1_sg U11854 ( .A(\o_im[2][3] ), .B(n6885), .X(n3575) );
  nand_x1_sg U11855 ( .A(n6579), .B(n6935), .X(n3574) );
  nand_x1_sg U11856 ( .A(\o_im[2][2] ), .B(n6886), .X(n3573) );
  nand_x1_sg U11857 ( .A(n6612), .B(n6934), .X(n3572) );
  nand_x1_sg U11858 ( .A(\o_im[2][1] ), .B(n6885), .X(n3571) );
  nand_x1_sg U11859 ( .A(n6608), .B(n6104), .X(n3569) );
  nand_x1_sg U11860 ( .A(\o_im[2][0] ), .B(n6884), .X(n3568) );
  nand_x1_sg U11861 ( .A(n7271), .B(n9197), .X(n821) );
  inv_x2_sg U11862 ( .A(\i_im[14][15] ), .X(n9197) );
  nand_x1_sg U11863 ( .A(n7147), .B(n9043), .X(n1134) );
  inv_x2_sg U11864 ( .A(\i_im[5][1] ), .X(n9043) );
  nand_x1_sg U11865 ( .A(n7145), .B(n9058), .X(n838) );
  inv_x2_sg U11866 ( .A(\i_im[5][16] ), .X(n9058) );
  nor_x1_sg U11867 ( .A(n7295), .B(\i_im[3][8] ), .X(n1362) );
  nor_x1_sg U11868 ( .A(n7290), .B(\i_im[3][14] ), .X(n1098) );
  nor_x1_sg U11869 ( .A(n7291), .B(\i_im[3][13] ), .X(n1066) );
  nand_x1_sg U11870 ( .A(n6440), .B(n9025), .X(n1221) );
  inv_x2_sg U11871 ( .A(\i_im[4][3] ), .X(n9025) );
  nand_x1_sg U11872 ( .A(n6008), .B(n9033), .X(n1024) );
  inv_x2_sg U11873 ( .A(\i_im[4][11] ), .X(n9033) );
  nand_x1_sg U11874 ( .A(n6171), .B(n9161), .X(n943) );
  inv_x2_sg U11875 ( .A(\i_im[12][19] ), .X(n9161) );
  nand_x1_sg U11876 ( .A(n7462), .B(n9183), .X(n1149) );
  inv_x2_sg U11877 ( .A(\i_im[14][1] ), .X(n9183) );
  nand_x1_sg U11878 ( .A(n7264), .B(n9188), .X(n1312) );
  inv_x2_sg U11879 ( .A(\i_im[14][6] ), .X(n9188) );
  nand_x1_sg U11880 ( .A(n7269), .B(n9198), .X(n853) );
  inv_x2_sg U11881 ( .A(\i_im[14][16] ), .X(n9198) );
  nor_x1_sg U11882 ( .A(n7296), .B(\i_im[11][3] ), .X(n1246) );
  nor_x1_sg U11883 ( .A(n7301), .B(\i_im[11][11] ), .X(n1049) );
  nor_x1_sg U11884 ( .A(n7300), .B(\i_im[3][7] ), .X(n1330) );
  nor_x1_sg U11885 ( .A(n7291), .B(\i_im[3][11] ), .X(n1034) );
  nor_x1_sg U11886 ( .A(n7298), .B(\i_im[3][4] ), .X(n1199) );
  nor_x1_sg U11887 ( .A(n7294), .B(\i_im[3][0] ), .X(n1426) );
  nor_x1_sg U11888 ( .A(n7299), .B(\i_im[3][17] ), .X(n871) );
  nor_x1_sg U11889 ( .A(n7293), .B(\i_im[3][19] ), .X(n935) );
  nor_x1_sg U11890 ( .A(n7296), .B(\i_im[3][18] ), .X(n903) );
  nand_x1_sg U11891 ( .A(n6440), .B(n9146), .X(n1207) );
  inv_x2_sg U11892 ( .A(\i_im[12][4] ), .X(n9146) );
  nand_x1_sg U11893 ( .A(n6422), .B(n9049), .X(n1329) );
  inv_x2_sg U11894 ( .A(\i_im[5][7] ), .X(n9049) );
  nand_x1_sg U11895 ( .A(n6170), .B(n9030), .X(n1352) );
  nor_x1_sg U11896 ( .A(n7076), .B(\i_im[1][8] ), .X(n1353) );
  nor_x1_sg U11897 ( .A(n7300), .B(\i_im[11][8] ), .X(n1377) );
  nor_x1_sg U11898 ( .A(n7301), .B(\i_im[11][0] ), .X(n1444) );
  nor_x1_sg U11899 ( .A(n7295), .B(\i_im[11][13] ), .X(n1081) );
  nor_x1_sg U11900 ( .A(n7299), .B(\i_im[11][17] ), .X(n886) );
  nor_x1_sg U11901 ( .A(n7293), .B(\i_im[11][18] ), .X(n918) );
  nor_x1_sg U11902 ( .A(n7290), .B(\i_im[3][3] ), .X(n1231) );
  nand_x1_sg U11903 ( .A(n6323), .B(n9057), .X(n805) );
  inv_x2_sg U11904 ( .A(\i_im[5][15] ), .X(n9057) );
  nand_x1_sg U11905 ( .A(n6007), .B(n9041), .X(n925) );
  nor_x1_sg U11906 ( .A(n7080), .B(\i_im[1][19] ), .X(n926) );
  nand_x1_sg U11907 ( .A(n6324), .B(n9045), .X(n1230) );
  inv_x2_sg U11908 ( .A(\i_im[5][3] ), .X(n9045) );
  nor_x1_sg U11909 ( .A(n7298), .B(\i_im[11][4] ), .X(n1214) );
  nand_x1_sg U11910 ( .A(n6008), .B(n9035), .X(n1056) );
  inv_x2_sg U11911 ( .A(\i_im[4][13] ), .X(n9035) );
  nor_x1_sg U11912 ( .A(n880), .B(n881), .X(n878) );
  nand_x1_sg U11913 ( .A(n7084), .B(n9159), .X(n879) );
  nor_x1_sg U11914 ( .A(\i_im[10][17] ), .B(n7229), .X(n881) );
  nand_x1_sg U11915 ( .A(n6439), .B(n9026), .X(n1189) );
  nor_x1_sg U11916 ( .A(n7080), .B(\i_im[1][4] ), .X(n1190) );
  nor_x1_sg U11917 ( .A(n7289), .B(\i_im[11][19] ), .X(n950) );
  nor_x1_sg U11918 ( .A(n1436), .B(n1437), .X(n1434) );
  nand_x1_sg U11919 ( .A(n7085), .B(n9142), .X(n1435) );
  nor_x1_sg U11920 ( .A(\i_im[10][0] ), .B(n7239), .X(n1437) );
  nand_x1_sg U11921 ( .A(n6170), .B(n9039), .X(n861) );
  inv_x2_sg U11922 ( .A(\i_im[4][17] ), .X(n9039) );
  nand_x1_sg U11923 ( .A(n6439), .B(n9022), .X(n1416) );
  inv_x2_sg U11924 ( .A(\i_im[4][0] ), .X(n9022) );
  nand_x1_sg U11925 ( .A(n7085), .B(n9156), .X(n1106) );
  inv_x2_sg U11926 ( .A(\i_im[12][14] ), .X(n9156) );
  nor_x1_sg U11927 ( .A(n912), .B(n913), .X(n910) );
  nand_x1_sg U11928 ( .A(n6008), .B(n9160), .X(n911) );
  nor_x1_sg U11929 ( .A(\i_im[10][18] ), .B(n7240), .X(n913) );
  nand_x1_sg U11930 ( .A(n6007), .B(n9040), .X(n893) );
  inv_x2_sg U11931 ( .A(\i_im[4][18] ), .X(n9040) );
  nor_x1_sg U11932 ( .A(n7071), .B(\i_im[1][14] ), .X(n1089) );
  nor_x1_sg U11933 ( .A(n1403), .B(n1404), .X(n1401) );
  nor_x1_sg U11934 ( .A(\i_im[8][9] ), .B(n7152), .X(n1403) );
  nor_x1_sg U11935 ( .A(\i_im[10][9] ), .B(n7232), .X(n1404) );
  nand_x1_sg U11936 ( .A(n6129), .B(n9211), .X(n1407) );
  inv_x2_sg U11937 ( .A(\i_im[15][9] ), .X(n9211) );
  nor_x1_sg U11938 ( .A(n7231), .B(\i_im[2][9] ), .X(n1387) );
  nor_x1_sg U11939 ( .A(\i_im[8][0] ), .B(n7155), .X(n1436) );
  nor_x1_sg U11940 ( .A(\i_im[8][17] ), .B(n7161), .X(n880) );
  nor_x1_sg U11941 ( .A(\i_im[8][18] ), .B(n7156), .X(n912) );
  nor_x1_sg U11942 ( .A(n1339), .B(n1340), .X(n1337) );
  nor_x1_sg U11943 ( .A(\i_im[10][7] ), .B(n7236), .X(n1340) );
  nor_x1_sg U11944 ( .A(\i_im[8][7] ), .B(n7155), .X(n1339) );
  nor_x1_sg U11945 ( .A(n1371), .B(n1372), .X(n1369) );
  nor_x1_sg U11946 ( .A(\i_im[10][8] ), .B(n7234), .X(n1372) );
  nor_x1_sg U11947 ( .A(\i_im[8][8] ), .B(n7162), .X(n1371) );
  nor_x1_sg U11948 ( .A(n1208), .B(n1209), .X(n1206) );
  nor_x1_sg U11949 ( .A(\i_im[10][4] ), .B(n7240), .X(n1209) );
  nor_x1_sg U11950 ( .A(\i_im[8][4] ), .B(n7150), .X(n1208) );
  nor_x1_sg U11951 ( .A(n1043), .B(n1044), .X(n1041) );
  nor_x1_sg U11952 ( .A(\i_im[10][11] ), .B(n7239), .X(n1044) );
  nor_x1_sg U11953 ( .A(\i_im[8][11] ), .B(n7152), .X(n1043) );
  nor_x1_sg U11954 ( .A(n1075), .B(n1076), .X(n1073) );
  nor_x1_sg U11955 ( .A(\i_im[10][13] ), .B(n7235), .X(n1076) );
  nand_x1_sg U11956 ( .A(n7267), .B(n9071), .X(n1392) );
  nand_x1_sg U11957 ( .A(n7278), .B(n9091), .X(n1391) );
  inv_x2_sg U11958 ( .A(\i_im[6][9] ), .X(n9071) );
  nor_x1_sg U11959 ( .A(n1240), .B(n1241), .X(n1238) );
  nor_x1_sg U11960 ( .A(\i_im[10][3] ), .B(n7240), .X(n1241) );
  nor_x1_sg U11961 ( .A(\i_im[8][3] ), .B(n7156), .X(n1240) );
  nor_x1_sg U11962 ( .A(n944), .B(n945), .X(n942) );
  nor_x1_sg U11963 ( .A(\i_im[10][19] ), .B(n7235), .X(n945) );
  nor_x1_sg U11964 ( .A(\i_im[8][19] ), .B(n7151), .X(n944) );
  nor_x1_sg U11965 ( .A(n1107), .B(n1108), .X(n1105) );
  nor_x1_sg U11966 ( .A(\i_im[8][14] ), .B(n7157), .X(n1107) );
  nor_x1_sg U11967 ( .A(\i_im[10][14] ), .B(n7231), .X(n1108) );
  nand_x1_sg U11968 ( .A(n7281), .B(n9209), .X(n1343) );
  inv_x2_sg U11969 ( .A(\i_im[15][7] ), .X(n9209) );
  nor_x1_sg U11970 ( .A(n7232), .B(\i_im[2][7] ), .X(n1323) );
  nor_x1_sg U11971 ( .A(n7076), .B(\i_im[1][11] ), .X(n1025) );
  nor_x1_sg U11972 ( .A(n7075), .B(\i_im[1][13] ), .X(n1057) );
  nand_x1_sg U11973 ( .A(n6128), .B(n9096), .X(n1095) );
  inv_x2_sg U11974 ( .A(\i_im[7][14] ), .X(n9096) );
  nand_x1_sg U11975 ( .A(n7269), .B(n9069), .X(n1328) );
  nand_x1_sg U11976 ( .A(n7279), .B(n9089), .X(n1327) );
  inv_x2_sg U11977 ( .A(\i_im[6][7] ), .X(n9069) );
  nor_x1_sg U11978 ( .A(n7071), .B(\i_im[1][7] ), .X(n1321) );
  nor_x1_sg U11979 ( .A(n7076), .B(\i_im[1][9] ), .X(n1385) );
  nor_x1_sg U11980 ( .A(n7075), .B(\i_im[1][0] ), .X(n1417) );
  nor_x1_sg U11981 ( .A(n7072), .B(\i_im[1][17] ), .X(n862) );
  nor_x1_sg U11982 ( .A(n7078), .B(\i_im[1][18] ), .X(n894) );
  nor_x1_sg U11983 ( .A(\i_im[0][8] ), .B(n7159), .X(n1356) );
  nor_x1_sg U11984 ( .A(n6362), .B(n1060), .X(n1058) );
  nor_x1_sg U11985 ( .A(\i_im[0][13] ), .B(n7161), .X(n1060) );
  nor_x1_sg U11986 ( .A(n6361), .B(n1356), .X(n1354) );
  nor_x1_sg U11987 ( .A(n7234), .B(\i_im[2][8] ), .X(n1355) );
  nor_x1_sg U11988 ( .A(n7234), .B(\i_im[2][3] ), .X(n1224) );
  nor_x1_sg U11989 ( .A(n7230), .B(\i_im[2][11] ), .X(n1027) );
  nand_x1_sg U11990 ( .A(n6654), .B(n6959), .X(n3862) );
  nand_x1_sg U11991 ( .A(\o_im[8][17] ), .B(n6906), .X(n3863) );
  nand_x1_sg U11992 ( .A(n6646), .B(n6959), .X(n3858) );
  nand_x1_sg U11993 ( .A(\o_im[8][15] ), .B(n5982), .X(n3859) );
  nand_x1_sg U11994 ( .A(n6565), .B(n6960), .X(n3854) );
  nand_x1_sg U11995 ( .A(\o_im[8][13] ), .B(n6905), .X(n3855) );
  nand_x1_sg U11996 ( .A(n6569), .B(n6959), .X(n3850) );
  nand_x1_sg U11997 ( .A(\o_im[8][11] ), .B(n6904), .X(n3851) );
  nand_x1_sg U11998 ( .A(n6631), .B(n6960), .X(n3846) );
  nand_x1_sg U11999 ( .A(\o_im[8][9] ), .B(n6906), .X(n3847) );
  nand_x1_sg U12000 ( .A(n6625), .B(n6957), .X(n3842) );
  nand_x1_sg U12001 ( .A(\o_im[8][7] ), .B(n6904), .X(n3843) );
  nand_x1_sg U12002 ( .A(n6620), .B(n6958), .X(n3838) );
  nand_x1_sg U12003 ( .A(\o_im[8][5] ), .B(n6905), .X(n3839) );
  nand_x1_sg U12004 ( .A(n6577), .B(n6960), .X(n3834) );
  nand_x1_sg U12005 ( .A(\o_im[8][3] ), .B(n6903), .X(n3835) );
  nand_x1_sg U12006 ( .A(n6612), .B(n6109), .X(n3830) );
  nand_x1_sg U12007 ( .A(\o_im[8][1] ), .B(n6904), .X(n3831) );
  nand_x1_sg U12008 ( .A(n6653), .B(n6963), .X(n4118) );
  nand_x1_sg U12009 ( .A(\o_im[14][17] ), .B(n6881), .X(n4119) );
  nand_x1_sg U12010 ( .A(n6645), .B(n6963), .X(n4114) );
  nand_x1_sg U12011 ( .A(\o_im[14][15] ), .B(n6880), .X(n4115) );
  nand_x1_sg U12012 ( .A(n6564), .B(n6964), .X(n4110) );
  nand_x1_sg U12013 ( .A(\o_im[14][13] ), .B(n6879), .X(n4111) );
  nand_x1_sg U12014 ( .A(n6566), .B(n6110), .X(n4106) );
  nand_x1_sg U12015 ( .A(\o_im[14][11] ), .B(n5977), .X(n4107) );
  nand_x1_sg U12016 ( .A(n6634), .B(n6965), .X(n4102) );
  nand_x1_sg U12017 ( .A(\o_im[14][9] ), .B(n6882), .X(n4103) );
  nand_x1_sg U12018 ( .A(n6625), .B(n6965), .X(n4098) );
  nand_x1_sg U12019 ( .A(\o_im[14][7] ), .B(n6880), .X(n4099) );
  nand_x1_sg U12020 ( .A(n6621), .B(n6962), .X(n4094) );
  nand_x1_sg U12021 ( .A(\o_im[14][5] ), .B(n6879), .X(n4095) );
  nand_x1_sg U12022 ( .A(n6577), .B(n6110), .X(n4090) );
  nand_x1_sg U12023 ( .A(\o_im[14][3] ), .B(n5977), .X(n4091) );
  nand_x1_sg U12024 ( .A(n6614), .B(n6110), .X(n4086) );
  nand_x1_sg U12025 ( .A(\o_im[14][1] ), .B(n6880), .X(n4087) );
  nand_x1_sg U12026 ( .A(n6653), .B(n6113), .X(n3990) );
  nand_x1_sg U12027 ( .A(\o_im[11][17] ), .B(n6866), .X(n3991) );
  nand_x1_sg U12028 ( .A(n6646), .B(n6980), .X(n3986) );
  nand_x1_sg U12029 ( .A(\o_im[11][15] ), .B(n6865), .X(n3987) );
  nand_x1_sg U12030 ( .A(n6562), .B(n6113), .X(n3982) );
  nand_x1_sg U12031 ( .A(\o_im[11][13] ), .B(n5974), .X(n3983) );
  nand_x1_sg U12032 ( .A(n6567), .B(n6979), .X(n3978) );
  nand_x1_sg U12033 ( .A(\o_im[11][11] ), .B(n6866), .X(n3979) );
  nand_x1_sg U12034 ( .A(n6632), .B(n6977), .X(n3974) );
  nand_x1_sg U12035 ( .A(\o_im[11][9] ), .B(n6867), .X(n3975) );
  nand_x1_sg U12036 ( .A(n6625), .B(n6978), .X(n3970) );
  nand_x1_sg U12037 ( .A(\o_im[11][7] ), .B(n5974), .X(n3971) );
  nand_x1_sg U12038 ( .A(n6622), .B(n6977), .X(n3966) );
  nand_x1_sg U12039 ( .A(\o_im[11][5] ), .B(n6866), .X(n3967) );
  nand_x1_sg U12040 ( .A(n6574), .B(n6979), .X(n3962) );
  nand_x1_sg U12041 ( .A(\o_im[11][3] ), .B(n5974), .X(n3963) );
  nand_x1_sg U12042 ( .A(n6612), .B(n6113), .X(n3958) );
  nand_x1_sg U12043 ( .A(\o_im[11][1] ), .B(n5974), .X(n3959) );
  nand_x1_sg U12044 ( .A(n6652), .B(n6927), .X(n3905) );
  nand_x1_sg U12045 ( .A(\o_im[9][17] ), .B(n6855), .X(n3906) );
  nand_x1_sg U12046 ( .A(n6644), .B(n6927), .X(n3901) );
  nand_x1_sg U12047 ( .A(\o_im[9][15] ), .B(n6856), .X(n3902) );
  nand_x1_sg U12048 ( .A(n6564), .B(n6930), .X(n3897) );
  nand_x1_sg U12049 ( .A(\o_im[9][13] ), .B(n6855), .X(n3898) );
  nand_x1_sg U12050 ( .A(n6568), .B(n6928), .X(n3893) );
  nand_x1_sg U12051 ( .A(\o_im[9][11] ), .B(n5972), .X(n3894) );
  nand_x1_sg U12052 ( .A(n6632), .B(n6927), .X(n3889) );
  nand_x1_sg U12053 ( .A(\o_im[9][9] ), .B(n6857), .X(n3890) );
  nand_x1_sg U12054 ( .A(n6626), .B(n6103), .X(n3885) );
  nand_x1_sg U12055 ( .A(\o_im[9][7] ), .B(n6854), .X(n3886) );
  nand_x1_sg U12056 ( .A(n6619), .B(n6929), .X(n3881) );
  nand_x1_sg U12057 ( .A(\o_im[9][5] ), .B(n5972), .X(n3882) );
  nand_x1_sg U12058 ( .A(n6575), .B(n6929), .X(n3877) );
  nand_x1_sg U12059 ( .A(\o_im[9][3] ), .B(n5972), .X(n3878) );
  nand_x1_sg U12060 ( .A(n6613), .B(n6929), .X(n3873) );
  nand_x1_sg U12061 ( .A(\o_im[9][1] ), .B(n6854), .X(n3874) );
  nand_x1_sg U12062 ( .A(n6652), .B(n6102), .X(n4033) );
  nand_x1_sg U12063 ( .A(\o_im[12][17] ), .B(n6862), .X(n4034) );
  nand_x1_sg U12064 ( .A(n6643), .B(n6102), .X(n4029) );
  nand_x1_sg U12065 ( .A(\o_im[12][15] ), .B(n6860), .X(n4030) );
  nand_x1_sg U12066 ( .A(n6565), .B(n6923), .X(n4025) );
  nand_x1_sg U12067 ( .A(\o_im[12][13] ), .B(n5973), .X(n4026) );
  nand_x1_sg U12068 ( .A(n6569), .B(n6922), .X(n4021) );
  nand_x1_sg U12069 ( .A(\o_im[12][11] ), .B(n6859), .X(n4022) );
  nand_x1_sg U12070 ( .A(n6632), .B(n6923), .X(n4017) );
  nand_x1_sg U12071 ( .A(\o_im[12][9] ), .B(n6861), .X(n4018) );
  nand_x1_sg U12072 ( .A(n6623), .B(n6924), .X(n4013) );
  nand_x1_sg U12073 ( .A(\o_im[12][7] ), .B(n6861), .X(n4014) );
  nand_x1_sg U12074 ( .A(n6619), .B(n6925), .X(n4009) );
  nand_x1_sg U12075 ( .A(\o_im[12][5] ), .B(n6859), .X(n4010) );
  nand_x1_sg U12076 ( .A(n6576), .B(n6922), .X(n4005) );
  nand_x1_sg U12077 ( .A(\o_im[12][3] ), .B(n6861), .X(n4006) );
  nand_x1_sg U12078 ( .A(n6611), .B(n6925), .X(n4001) );
  nand_x1_sg U12079 ( .A(\o_im[12][1] ), .B(n5973), .X(n4002) );
  nand_x1_sg U12080 ( .A(n6653), .B(n6945), .X(n4076) );
  nand_x1_sg U12081 ( .A(\o_im[13][17] ), .B(n6850), .X(n4077) );
  nand_x1_sg U12082 ( .A(n6645), .B(n6944), .X(n4072) );
  nand_x1_sg U12083 ( .A(\o_im[13][15] ), .B(n5971), .X(n4073) );
  nand_x1_sg U12084 ( .A(n6562), .B(n6945), .X(n4068) );
  nand_x1_sg U12085 ( .A(\o_im[13][13] ), .B(n6851), .X(n4069) );
  nand_x1_sg U12086 ( .A(n6568), .B(n6106), .X(n4064) );
  nand_x1_sg U12087 ( .A(\o_im[13][11] ), .B(n6850), .X(n4065) );
  nand_x1_sg U12088 ( .A(n6634), .B(n6942), .X(n4060) );
  nand_x1_sg U12089 ( .A(\o_im[13][9] ), .B(n6852), .X(n4061) );
  nand_x1_sg U12090 ( .A(n6626), .B(n6106), .X(n4056) );
  nand_x1_sg U12091 ( .A(\o_im[13][7] ), .B(n5971), .X(n4057) );
  nand_x1_sg U12092 ( .A(n6622), .B(n6106), .X(n4052) );
  nand_x1_sg U12093 ( .A(\o_im[13][5] ), .B(n6849), .X(n4053) );
  nand_x1_sg U12094 ( .A(n6574), .B(n6945), .X(n4048) );
  nand_x1_sg U12095 ( .A(\o_im[13][3] ), .B(n6850), .X(n4049) );
  nand_x1_sg U12096 ( .A(n6614), .B(n6942), .X(n4044) );
  nand_x1_sg U12097 ( .A(\o_im[13][1] ), .B(n6849), .X(n4045) );
  nand_x1_sg U12098 ( .A(n6652), .B(n6949), .X(n3947) );
  nand_x1_sg U12099 ( .A(\o_im[10][17] ), .B(n6911), .X(n3948) );
  nand_x1_sg U12100 ( .A(n6644), .B(n6948), .X(n3943) );
  nand_x1_sg U12101 ( .A(\o_im[10][15] ), .B(n5983), .X(n3944) );
  nand_x1_sg U12102 ( .A(n6564), .B(n6107), .X(n3939) );
  nand_x1_sg U12103 ( .A(\o_im[10][13] ), .B(n6909), .X(n3940) );
  nand_x1_sg U12104 ( .A(n6567), .B(n6107), .X(n3935) );
  nand_x1_sg U12105 ( .A(\o_im[10][11] ), .B(n6909), .X(n3936) );
  nand_x1_sg U12106 ( .A(n6631), .B(n6948), .X(n3931) );
  nand_x1_sg U12107 ( .A(\o_im[10][9] ), .B(n6911), .X(n3932) );
  nand_x1_sg U12108 ( .A(n6624), .B(n6950), .X(n3927) );
  nand_x1_sg U12109 ( .A(\o_im[10][7] ), .B(n6908), .X(n3928) );
  nand_x1_sg U12110 ( .A(n6620), .B(n6950), .X(n3923) );
  nand_x1_sg U12111 ( .A(\o_im[10][5] ), .B(n5983), .X(n3924) );
  nand_x1_sg U12112 ( .A(n6576), .B(n6948), .X(n3919) );
  nand_x1_sg U12113 ( .A(\o_im[10][3] ), .B(n6909), .X(n3920) );
  nand_x1_sg U12114 ( .A(n6612), .B(n6949), .X(n3915) );
  nand_x1_sg U12115 ( .A(\o_im[10][1] ), .B(n6909), .X(n3916) );
  nand_x1_sg U12116 ( .A(n6660), .B(n6930), .X(n3909) );
  nand_x1_sg U12117 ( .A(\o_im[9][19] ), .B(n6854), .X(n3910) );
  nand_x1_sg U12118 ( .A(n6656), .B(n6103), .X(n3907) );
  nand_x1_sg U12119 ( .A(\o_im[9][18] ), .B(n6857), .X(n3908) );
  nand_x1_sg U12120 ( .A(n6648), .B(n6928), .X(n3903) );
  nand_x1_sg U12121 ( .A(\o_im[9][16] ), .B(n6855), .X(n3904) );
  nand_x1_sg U12122 ( .A(n6558), .B(n6930), .X(n3899) );
  nand_x1_sg U12123 ( .A(\o_im[9][14] ), .B(n6856), .X(n3900) );
  nand_x1_sg U12124 ( .A(n6640), .B(n6927), .X(n3895) );
  nand_x1_sg U12125 ( .A(\o_im[9][12] ), .B(n6856), .X(n3896) );
  nand_x1_sg U12126 ( .A(n6637), .B(n6103), .X(n3891) );
  nand_x1_sg U12127 ( .A(\o_im[9][10] ), .B(n6854), .X(n3892) );
  nand_x1_sg U12128 ( .A(n6627), .B(n6103), .X(n3887) );
  nand_x1_sg U12129 ( .A(\o_im[9][8] ), .B(n6856), .X(n3888) );
  nand_x1_sg U12130 ( .A(n6571), .B(n6930), .X(n3883) );
  nand_x1_sg U12131 ( .A(\o_im[9][6] ), .B(n6855), .X(n3884) );
  nand_x1_sg U12132 ( .A(n6618), .B(n6929), .X(n3879) );
  nand_x1_sg U12133 ( .A(\o_im[9][4] ), .B(n5972), .X(n3880) );
  nand_x1_sg U12134 ( .A(n6580), .B(n6928), .X(n3875) );
  nand_x1_sg U12135 ( .A(\o_im[9][2] ), .B(n6857), .X(n3876) );
  nand_x1_sg U12136 ( .A(n6607), .B(n6928), .X(n3870) );
  nand_x1_sg U12137 ( .A(\o_im[9][0] ), .B(n6857), .X(n3871) );
  nand_x1_sg U12138 ( .A(n6661), .B(n6923), .X(n4037) );
  nand_x1_sg U12139 ( .A(\o_im[12][19] ), .B(n5973), .X(n4038) );
  nand_x1_sg U12140 ( .A(n6655), .B(n6923), .X(n4035) );
  nand_x1_sg U12141 ( .A(\o_im[12][18] ), .B(n6860), .X(n4036) );
  nand_x1_sg U12142 ( .A(n6649), .B(n6922), .X(n4031) );
  nand_x1_sg U12143 ( .A(\o_im[12][16] ), .B(n6862), .X(n4032) );
  nand_x1_sg U12144 ( .A(n6561), .B(n6925), .X(n4027) );
  nand_x1_sg U12145 ( .A(\o_im[12][14] ), .B(n6859), .X(n4028) );
  nand_x1_sg U12146 ( .A(n6642), .B(n6925), .X(n4023) );
  nand_x1_sg U12147 ( .A(\o_im[12][12] ), .B(n5973), .X(n4024) );
  nand_x1_sg U12148 ( .A(n6638), .B(n6924), .X(n4019) );
  nand_x1_sg U12149 ( .A(\o_im[12][10] ), .B(n6860), .X(n4020) );
  nand_x1_sg U12150 ( .A(n6629), .B(n6102), .X(n4015) );
  nand_x1_sg U12151 ( .A(\o_im[12][8] ), .B(n6861), .X(n4016) );
  nand_x1_sg U12152 ( .A(n6570), .B(n6102), .X(n4011) );
  nand_x1_sg U12153 ( .A(\o_im[12][6] ), .B(n6859), .X(n4012) );
  nand_x1_sg U12154 ( .A(n6615), .B(n6922), .X(n4007) );
  nand_x1_sg U12155 ( .A(\o_im[12][4] ), .B(n6860), .X(n4008) );
  nand_x1_sg U12156 ( .A(n6579), .B(n6924), .X(n4003) );
  nand_x1_sg U12157 ( .A(\o_im[12][2] ), .B(n6862), .X(n4004) );
  nand_x1_sg U12158 ( .A(n6610), .B(n6924), .X(n3998) );
  nand_x1_sg U12159 ( .A(\o_im[12][0] ), .B(n6862), .X(n3999) );
  nand_x1_sg U12160 ( .A(n6662), .B(n6990), .X(n4818) );
  nand_x1_sg U12161 ( .A(\o_im[15][19] ), .B(n6839), .X(n4819) );
  nand_x1_sg U12162 ( .A(n6659), .B(n6944), .X(n4080) );
  nand_x1_sg U12163 ( .A(\o_im[13][19] ), .B(n6849), .X(n4081) );
  nand_x1_sg U12164 ( .A(n6656), .B(n6944), .X(n4078) );
  nand_x1_sg U12165 ( .A(\o_im[13][18] ), .B(n6852), .X(n4079) );
  nand_x1_sg U12166 ( .A(n6649), .B(n6945), .X(n4074) );
  nand_x1_sg U12167 ( .A(\o_im[13][16] ), .B(n6852), .X(n4075) );
  nand_x1_sg U12168 ( .A(n6560), .B(n6106), .X(n4070) );
  nand_x1_sg U12169 ( .A(\o_im[13][14] ), .B(n6851), .X(n4071) );
  nand_x1_sg U12170 ( .A(n6641), .B(n6943), .X(n4066) );
  nand_x1_sg U12171 ( .A(\o_im[13][12] ), .B(n6849), .X(n4067) );
  nand_x1_sg U12172 ( .A(n6637), .B(n6942), .X(n4062) );
  nand_x1_sg U12173 ( .A(\o_im[13][10] ), .B(n5971), .X(n4063) );
  nand_x1_sg U12174 ( .A(n6630), .B(n6943), .X(n4058) );
  nand_x1_sg U12175 ( .A(\o_im[13][8] ), .B(n5971), .X(n4059) );
  nand_x1_sg U12176 ( .A(n6572), .B(n6942), .X(n4054) );
  nand_x1_sg U12177 ( .A(\o_im[13][6] ), .B(n6851), .X(n4055) );
  nand_x1_sg U12178 ( .A(n6615), .B(n6943), .X(n4050) );
  nand_x1_sg U12179 ( .A(\o_im[13][4] ), .B(n6851), .X(n4051) );
  nand_x1_sg U12180 ( .A(n6579), .B(n6944), .X(n4046) );
  nand_x1_sg U12181 ( .A(\o_im[13][2] ), .B(n6852), .X(n4047) );
  nand_x1_sg U12182 ( .A(n6608), .B(n6943), .X(n4041) );
  nand_x1_sg U12183 ( .A(\o_im[13][0] ), .B(n6850), .X(n4042) );
  nand_x1_sg U12184 ( .A(n6660), .B(n6107), .X(n3951) );
  nand_x1_sg U12185 ( .A(\o_im[10][19] ), .B(n5983), .X(n3952) );
  nand_x1_sg U12186 ( .A(n6656), .B(n6947), .X(n3949) );
  nand_x1_sg U12187 ( .A(\o_im[10][18] ), .B(n6911), .X(n3950) );
  nand_x1_sg U12188 ( .A(n6647), .B(n6949), .X(n3945) );
  nand_x1_sg U12189 ( .A(\o_im[10][16] ), .B(n6910), .X(n3946) );
  nand_x1_sg U12190 ( .A(n6559), .B(n6950), .X(n3941) );
  nand_x1_sg U12191 ( .A(\o_im[10][14] ), .B(n6911), .X(n3942) );
  nand_x1_sg U12192 ( .A(n6640), .B(n6949), .X(n3937) );
  nand_x1_sg U12193 ( .A(\o_im[10][12] ), .B(n6908), .X(n3938) );
  nand_x1_sg U12194 ( .A(n6635), .B(n6950), .X(n3933) );
  nand_x1_sg U12195 ( .A(\o_im[10][10] ), .B(n6910), .X(n3934) );
  nand_x1_sg U12196 ( .A(n6628), .B(n6948), .X(n3929) );
  nand_x1_sg U12197 ( .A(\o_im[10][8] ), .B(n5983), .X(n3930) );
  nand_x1_sg U12198 ( .A(n6571), .B(n6947), .X(n3925) );
  nand_x1_sg U12199 ( .A(\o_im[10][6] ), .B(n6908), .X(n3926) );
  nand_x1_sg U12200 ( .A(n6617), .B(n6947), .X(n3921) );
  nand_x1_sg U12201 ( .A(\o_im[10][4] ), .B(n6910), .X(n3922) );
  nand_x1_sg U12202 ( .A(n6579), .B(n6947), .X(n3917) );
  nand_x1_sg U12203 ( .A(\o_im[10][2] ), .B(n6910), .X(n3918) );
  nand_x1_sg U12204 ( .A(n6608), .B(n6107), .X(n3912) );
  nand_x1_sg U12205 ( .A(\o_im[10][0] ), .B(n6908), .X(n3913) );
  nand_x1_sg U12206 ( .A(n6662), .B(n6109), .X(n3866) );
  nand_x1_sg U12207 ( .A(\o_im[8][19] ), .B(n6903), .X(n3867) );
  nand_x1_sg U12208 ( .A(n6655), .B(n6109), .X(n3864) );
  nand_x1_sg U12209 ( .A(\o_im[8][18] ), .B(n6906), .X(n3865) );
  nand_x1_sg U12210 ( .A(n6647), .B(n6960), .X(n3860) );
  nand_x1_sg U12211 ( .A(\o_im[8][16] ), .B(n6903), .X(n3861) );
  nand_x1_sg U12212 ( .A(n6561), .B(n6109), .X(n3856) );
  nand_x1_sg U12213 ( .A(\o_im[8][14] ), .B(n6903), .X(n3857) );
  nand_x1_sg U12214 ( .A(n6642), .B(n6957), .X(n3852) );
  nand_x1_sg U12215 ( .A(\o_im[8][12] ), .B(n6905), .X(n3853) );
  nand_x1_sg U12216 ( .A(n6636), .B(n6958), .X(n3848) );
  nand_x1_sg U12217 ( .A(\o_im[8][10] ), .B(n6905), .X(n3849) );
  nand_x1_sg U12218 ( .A(n6629), .B(n6958), .X(n3844) );
  nand_x1_sg U12219 ( .A(\o_im[8][8] ), .B(n5982), .X(n3845) );
  nand_x1_sg U12220 ( .A(n6572), .B(n6957), .X(n3840) );
  nand_x1_sg U12221 ( .A(\o_im[8][6] ), .B(n5982), .X(n3841) );
  nand_x1_sg U12222 ( .A(n6618), .B(n6958), .X(n3836) );
  nand_x1_sg U12223 ( .A(\o_im[8][4] ), .B(n5982), .X(n3837) );
  nand_x1_sg U12224 ( .A(n6578), .B(n6957), .X(n3832) );
  nand_x1_sg U12225 ( .A(\o_im[8][2] ), .B(n6904), .X(n3833) );
  nand_x1_sg U12226 ( .A(n6609), .B(n6959), .X(n3827) );
  nand_x1_sg U12227 ( .A(\o_im[8][0] ), .B(n6906), .X(n3828) );
  nand_x1_sg U12228 ( .A(n6662), .B(n6964), .X(n4122) );
  nand_x1_sg U12229 ( .A(\o_im[14][19] ), .B(n5977), .X(n4123) );
  nand_x1_sg U12230 ( .A(n6657), .B(n6962), .X(n4120) );
  nand_x1_sg U12231 ( .A(\o_im[14][18] ), .B(n6882), .X(n4121) );
  nand_x1_sg U12232 ( .A(n6650), .B(n6110), .X(n4116) );
  nand_x1_sg U12233 ( .A(\o_im[14][16] ), .B(n6881), .X(n4117) );
  nand_x1_sg U12234 ( .A(n6560), .B(n6962), .X(n4112) );
  nand_x1_sg U12235 ( .A(\o_im[14][14] ), .B(n6882), .X(n4113) );
  nand_x1_sg U12236 ( .A(n6639), .B(n6965), .X(n4108) );
  nand_x1_sg U12237 ( .A(\o_im[14][12] ), .B(n6880), .X(n4109) );
  nand_x1_sg U12238 ( .A(n6637), .B(n6963), .X(n4104) );
  nand_x1_sg U12239 ( .A(\o_im[14][10] ), .B(n5977), .X(n4105) );
  nand_x1_sg U12240 ( .A(n6629), .B(n6962), .X(n4100) );
  nand_x1_sg U12241 ( .A(\o_im[14][8] ), .B(n6881), .X(n4101) );
  nand_x1_sg U12242 ( .A(n6573), .B(n6964), .X(n4096) );
  nand_x1_sg U12243 ( .A(\o_im[14][6] ), .B(n6881), .X(n4097) );
  nand_x1_sg U12244 ( .A(n6617), .B(n6964), .X(n4092) );
  nand_x1_sg U12245 ( .A(\o_im[14][4] ), .B(n6879), .X(n4093) );
  nand_x1_sg U12246 ( .A(n6581), .B(n6965), .X(n4088) );
  nand_x1_sg U12247 ( .A(\o_im[14][2] ), .B(n6882), .X(n4089) );
  nand_x1_sg U12248 ( .A(n6607), .B(n6963), .X(n4083) );
  nand_x1_sg U12249 ( .A(\o_im[14][0] ), .B(n6879), .X(n4084) );
  nand_x1_sg U12250 ( .A(n6660), .B(n6977), .X(n3994) );
  nand_x1_sg U12251 ( .A(\o_im[11][19] ), .B(n6866), .X(n3995) );
  nand_x1_sg U12252 ( .A(n6657), .B(n6978), .X(n3992) );
  nand_x1_sg U12253 ( .A(\o_im[11][18] ), .B(n6865), .X(n3993) );
  nand_x1_sg U12254 ( .A(n6648), .B(n6980), .X(n3988) );
  nand_x1_sg U12255 ( .A(\o_im[11][16] ), .B(n6867), .X(n3989) );
  nand_x1_sg U12256 ( .A(n6558), .B(n6978), .X(n3984) );
  nand_x1_sg U12257 ( .A(\o_im[11][14] ), .B(n6864), .X(n3985) );
  nand_x1_sg U12258 ( .A(n6640), .B(n6979), .X(n3980) );
  nand_x1_sg U12259 ( .A(\o_im[11][12] ), .B(n6864), .X(n3981) );
  nand_x1_sg U12260 ( .A(n6635), .B(n6980), .X(n3976) );
  nand_x1_sg U12261 ( .A(\o_im[11][10] ), .B(n6864), .X(n3977) );
  nand_x1_sg U12262 ( .A(n6630), .B(n6113), .X(n3972) );
  nand_x1_sg U12263 ( .A(\o_im[11][8] ), .B(n6865), .X(n3973) );
  nand_x1_sg U12264 ( .A(n6573), .B(n6978), .X(n3968) );
  nand_x1_sg U12265 ( .A(\o_im[11][6] ), .B(n6865), .X(n3969) );
  nand_x1_sg U12266 ( .A(n6616), .B(n6980), .X(n3964) );
  nand_x1_sg U12267 ( .A(\o_im[11][4] ), .B(n6864), .X(n3965) );
  nand_x1_sg U12268 ( .A(n6580), .B(n6977), .X(n3960) );
  nand_x1_sg U12269 ( .A(\o_im[11][2] ), .B(n6867), .X(n3961) );
  nand_x1_sg U12270 ( .A(n6610), .B(n6979), .X(n3955) );
  nand_x1_sg U12271 ( .A(\o_im[11][0] ), .B(n6867), .X(n3956) );
  nor_x1_sg U12272 ( .A(n7077), .B(\i_im[9][13] ), .X(n1072) );
  nor_x1_sg U12273 ( .A(n7077), .B(\i_im[9][8] ), .X(n1368) );
  nor_x1_sg U12274 ( .A(n7073), .B(\i_im[1][3] ), .X(n1222) );
  nor_x1_sg U12275 ( .A(\i_im[0][7] ), .B(n7162), .X(n1324) );
  nor_x1_sg U12276 ( .A(\i_im[0][9] ), .B(n7161), .X(n1388) );
  nor_x1_sg U12277 ( .A(\i_im[0][4] ), .B(n7162), .X(n1193) );
  nor_x1_sg U12278 ( .A(\i_im[0][11] ), .B(n7153), .X(n1028) );
  nor_x1_sg U12279 ( .A(\i_im[8][13] ), .B(n7150), .X(n1075) );
  nor_x1_sg U12280 ( .A(n7322), .B(n1420), .X(n1418) );
  nor_x1_sg U12281 ( .A(\i_im[0][0] ), .B(n7151), .X(n1420) );
  nor_x1_sg U12282 ( .A(n6082), .B(n865), .X(n863) );
  nor_x1_sg U12283 ( .A(\i_im[0][17] ), .B(n7156), .X(n865) );
  nor_x1_sg U12284 ( .A(n6361), .B(n897), .X(n895) );
  nor_x1_sg U12285 ( .A(\i_im[0][18] ), .B(n7157), .X(n897) );
  nand_x1_sg U12286 ( .A(n6655), .B(n6989), .X(n4783) );
  nand_x1_sg U12287 ( .A(\o_im[15][18] ), .B(n6840), .X(n4782) );
  nand_x1_sg U12288 ( .A(n6651), .B(n6987), .X(n4747) );
  nand_x1_sg U12289 ( .A(\o_im[15][17] ), .B(n5969), .X(n4746) );
  nand_x1_sg U12290 ( .A(n6648), .B(n6988), .X(n4711) );
  nand_x1_sg U12291 ( .A(\o_im[15][16] ), .B(n6841), .X(n4710) );
  nand_x1_sg U12292 ( .A(n6643), .B(n6115), .X(n4675) );
  nand_x1_sg U12293 ( .A(\o_im[15][15] ), .B(n6839), .X(n4674) );
  nand_x1_sg U12294 ( .A(n6558), .B(n6988), .X(n4639) );
  nand_x1_sg U12295 ( .A(\o_im[15][14] ), .B(n6842), .X(n4638) );
  nand_x1_sg U12296 ( .A(n6565), .B(n6989), .X(n4603) );
  nand_x1_sg U12297 ( .A(\o_im[15][13] ), .B(n6840), .X(n4602) );
  nand_x1_sg U12298 ( .A(n6639), .B(n6987), .X(n4567) );
  nand_x1_sg U12299 ( .A(\o_im[15][12] ), .B(n5969), .X(n4566) );
  nand_x1_sg U12300 ( .A(n6569), .B(n6987), .X(n4531) );
  nand_x1_sg U12301 ( .A(\o_im[15][11] ), .B(n5969), .X(n4530) );
  nand_x1_sg U12302 ( .A(n6635), .B(n6989), .X(n4495) );
  nand_x1_sg U12303 ( .A(\o_im[15][10] ), .B(n6841), .X(n4494) );
  nand_x1_sg U12304 ( .A(n6632), .B(n6990), .X(n4459) );
  nand_x1_sg U12305 ( .A(\o_im[15][9] ), .B(n6840), .X(n4458) );
  nand_x1_sg U12306 ( .A(n6627), .B(n6990), .X(n4423) );
  nand_x1_sg U12307 ( .A(\o_im[15][8] ), .B(n6842), .X(n4422) );
  nand_x1_sg U12308 ( .A(n6623), .B(n6989), .X(n4387) );
  nand_x1_sg U12309 ( .A(\o_im[15][7] ), .B(n6839), .X(n4386) );
  nand_x1_sg U12310 ( .A(n6570), .B(n6988), .X(n4351) );
  nand_x1_sg U12311 ( .A(\o_im[15][6] ), .B(n6840), .X(n4350) );
  nand_x1_sg U12312 ( .A(n6619), .B(n6988), .X(n4315) );
  nand_x1_sg U12313 ( .A(\o_im[15][5] ), .B(n6839), .X(n4314) );
  nand_x1_sg U12314 ( .A(n6616), .B(n6115), .X(n4279) );
  nand_x1_sg U12315 ( .A(\o_im[15][4] ), .B(n6841), .X(n4278) );
  nand_x1_sg U12316 ( .A(n6574), .B(n6115), .X(n4243) );
  nand_x1_sg U12317 ( .A(\o_im[15][3] ), .B(n6842), .X(n4242) );
  nand_x1_sg U12318 ( .A(n6578), .B(n6990), .X(n4207) );
  nand_x1_sg U12319 ( .A(\o_im[15][2] ), .B(n6842), .X(n4206) );
  nand_x1_sg U12320 ( .A(n6611), .B(n6987), .X(n4171) );
  nand_x1_sg U12321 ( .A(\o_im[15][1] ), .B(n6841), .X(n4170) );
  nand_x1_sg U12322 ( .A(n6607), .B(n6115), .X(n4128) );
  nand_x1_sg U12323 ( .A(\o_im[15][0] ), .B(n5969), .X(n4127) );
  nor_x1_sg U12324 ( .A(n6241), .B(n1193), .X(n1191) );
  nor_x1_sg U12325 ( .A(n7229), .B(\i_im[2][4] ), .X(n1192) );
  nand_x1_sg U12326 ( .A(n6128), .B(n9210), .X(n1375) );
  inv_x2_sg U12327 ( .A(\i_im[15][8] ), .X(n9210) );
  nand_x1_sg U12328 ( .A(n6490), .B(n9205), .X(n1244) );
  inv_x2_sg U12329 ( .A(\i_im[15][3] ), .X(n9205) );
  nand_x1_sg U12330 ( .A(n7146), .B(n9171), .X(n1399) );
  inv_x2_sg U12331 ( .A(\i_im[13][9] ), .X(n9171) );
  nand_x1_sg U12332 ( .A(n7270), .B(n9065), .X(n1229) );
  nand_x1_sg U12333 ( .A(n6389), .B(n9085), .X(n1228) );
  inv_x2_sg U12334 ( .A(\i_im[6][3] ), .X(n9065) );
  nand_x1_sg U12335 ( .A(n7147), .B(n9175), .X(n1071) );
  inv_x2_sg U12336 ( .A(\i_im[13][13] ), .X(n9175) );
  nor_x1_sg U12337 ( .A(n7073), .B(\i_im[9][9] ), .X(n1400) );
  nor_x1_sg U12338 ( .A(n7070), .B(\i_im[9][0] ), .X(n1432) );
  nor_x1_sg U12339 ( .A(n7080), .B(\i_im[9][17] ), .X(n877) );
  nor_x1_sg U12340 ( .A(n7072), .B(\i_im[9][18] ), .X(n909) );
  nor_x1_sg U12341 ( .A(n7075), .B(\i_im[9][7] ), .X(n1336) );
  nor_x1_sg U12342 ( .A(n7081), .B(\i_im[9][4] ), .X(n1205) );
  nor_x1_sg U12343 ( .A(n7073), .B(\i_im[9][11] ), .X(n1040) );
  nor_x1_sg U12344 ( .A(n7072), .B(\i_im[9][14] ), .X(n1104) );
  nor_x1_sg U12345 ( .A(n7068), .B(\i_im[9][19] ), .X(n941) );
  nor_x1_sg U12346 ( .A(\i_im[0][3] ), .B(n7153), .X(n1225) );
  nor_x1_sg U12347 ( .A(\i_im[0][19] ), .B(n7160), .X(n929) );
  nor_x1_sg U12348 ( .A(n5927), .B(n929), .X(n927) );
  nor_x1_sg U12349 ( .A(n7235), .B(\i_im[2][19] ), .X(n928) );
  nand_x1_sg U12350 ( .A(n6390), .B(n9090), .X(n1359) );
  inv_x2_sg U12351 ( .A(\i_im[7][8] ), .X(n9090) );
  nand_x1_sg U12352 ( .A(n6492), .B(n9093), .X(n1031) );
  nand_x1_sg U12353 ( .A(n6422), .B(n9162), .X(n1431) );
  inv_x2_sg U12354 ( .A(\i_im[13][0] ), .X(n9162) );
  nand_x1_sg U12355 ( .A(n7144), .B(n9179), .X(n876) );
  inv_x2_sg U12356 ( .A(\i_im[13][17] ), .X(n9179) );
  nand_x1_sg U12357 ( .A(n7145), .B(n9180), .X(n908) );
  inv_x2_sg U12358 ( .A(\i_im[13][18] ), .X(n9180) );
  nor_x1_sg U12359 ( .A(n7078), .B(\i_im[9][3] ), .X(n1237) );
  nor_x1_sg U12360 ( .A(n7236), .B(\i_im[2][13] ), .X(n1059) );
  nand_x1_sg U12361 ( .A(n7281), .B(n9086), .X(n1196) );
  inv_x2_sg U12362 ( .A(\i_im[7][4] ), .X(n9086) );
  nand_x1_sg U12363 ( .A(n6491), .B(n9095), .X(n1063) );
  inv_x2_sg U12364 ( .A(\i_im[7][13] ), .X(n9095) );
  nand_x1_sg U12365 ( .A(n7280), .B(n9101), .X(n932) );
  inv_x2_sg U12366 ( .A(\i_im[7][19] ), .X(n9101) );
  nand_x1_sg U12367 ( .A(n6421), .B(n9056), .X(n1097) );
  inv_x2_sg U12368 ( .A(\i_im[5][14] ), .X(n9056) );
  nor_x1_sg U12369 ( .A(n7239), .B(\i_im[2][0] ), .X(n1419) );
  nor_x1_sg U12370 ( .A(n7238), .B(\i_im[2][17] ), .X(n864) );
  nor_x1_sg U12371 ( .A(n7230), .B(\i_im[2][18] ), .X(n896) );
  nor_x1_sg U12372 ( .A(\i_im[0][14] ), .B(n7151), .X(n1092) );
  nor_x1_sg U12373 ( .A(n6240), .B(n1092), .X(n1090) );
  nor_x1_sg U12374 ( .A(n7230), .B(\i_im[2][14] ), .X(n1091) );
  nand_x1_sg U12375 ( .A(n6389), .B(n9099), .X(n868) );
  inv_x2_sg U12376 ( .A(\i_im[7][17] ), .X(n9099) );
  nand_x1_sg U12377 ( .A(n7279), .B(n9202), .X(n1441) );
  inv_x2_sg U12378 ( .A(\i_im[15][0] ), .X(n9202) );
  nand_x1_sg U12379 ( .A(n6128), .B(n9082), .X(n1423) );
  inv_x2_sg U12380 ( .A(\i_im[7][0] ), .X(n9082) );
  nand_x1_sg U12381 ( .A(n6421), .B(n9050), .X(n1361) );
  inv_x2_sg U12382 ( .A(\i_im[5][8] ), .X(n9050) );
  nand_x1_sg U12383 ( .A(n6390), .B(n9100), .X(n900) );
  inv_x2_sg U12384 ( .A(\i_im[7][18] ), .X(n9100) );
  nand_x1_sg U12385 ( .A(n6323), .B(n9046), .X(n1198) );
  inv_x2_sg U12386 ( .A(\i_im[5][4] ), .X(n9046) );
  nand_x1_sg U12387 ( .A(n6035), .B(n9055), .X(n1065) );
  inv_x2_sg U12388 ( .A(\i_im[5][13] ), .X(n9055) );
  nand_x1_sg U12389 ( .A(n6035), .B(n9059), .X(n870) );
  inv_x2_sg U12390 ( .A(\i_im[5][17] ), .X(n9059) );
  nand_x1_sg U12391 ( .A(n7146), .B(n9042), .X(n1425) );
  inv_x2_sg U12392 ( .A(\i_im[5][0] ), .X(n9042) );
  nand_x1_sg U12393 ( .A(n7267), .B(n9189), .X(n1344) );
  inv_x2_sg U12394 ( .A(\i_im[14][7] ), .X(n9189) );
  nand_x1_sg U12395 ( .A(n7260), .B(n9190), .X(n1376) );
  inv_x2_sg U12396 ( .A(\i_im[14][8] ), .X(n9190) );
  nand_x1_sg U12397 ( .A(n7268), .B(n9195), .X(n1080) );
  inv_x2_sg U12398 ( .A(\i_im[14][13] ), .X(n9195) );
  nand_x1_sg U12399 ( .A(n7267), .B(n9200), .X(n917) );
  inv_x2_sg U12400 ( .A(\i_im[14][18] ), .X(n9200) );
  nand_x1_sg U12401 ( .A(n7261), .B(n9191), .X(n1408) );
  inv_x2_sg U12402 ( .A(\i_im[14][9] ), .X(n9191) );
  nand_x1_sg U12403 ( .A(n7262), .B(n9186), .X(n1213) );
  inv_x2_sg U12404 ( .A(\i_im[14][4] ), .X(n9186) );
  nand_x1_sg U12405 ( .A(n7266), .B(n9185), .X(n1245) );
  inv_x2_sg U12406 ( .A(\i_im[14][3] ), .X(n9185) );
  nand_x1_sg U12407 ( .A(n7264), .B(n9182), .X(n1443) );
  inv_x2_sg U12408 ( .A(\i_im[14][0] ), .X(n9182) );
  nand_x1_sg U12409 ( .A(n7263), .B(n9196), .X(n1112) );
  inv_x2_sg U12410 ( .A(\i_im[14][14] ), .X(n9196) );
  nand_x1_sg U12411 ( .A(n7263), .B(n9199), .X(n885) );
  inv_x2_sg U12412 ( .A(\i_im[14][17] ), .X(n9199) );
  nand_x1_sg U12413 ( .A(n6324), .B(n9060), .X(n902) );
  inv_x2_sg U12414 ( .A(\i_im[5][18] ), .X(n9060) );
  nor_x1_sg U12415 ( .A(n6329), .B(\mask_state[0] ), .X(n5633) );
  nand_x1_sg U12416 ( .A(i_mask[21]), .B(n7341), .X(n4933) );
  nand_x1_sg U12417 ( .A(\update_mask_0/reg_i_mask[21] ), .B(n5992), .X(n4934)
         );
  nand_x1_sg U12418 ( .A(i_mask[6]), .B(n6260), .X(n4903) );
  nand_x1_sg U12419 ( .A(\update_mask_0/reg_i_mask[6] ), .B(n5997), .X(n4904)
         );
  nand_x1_sg U12420 ( .A(\i_im[15][19] ), .B(n7363), .X(n5593) );
  nand_x1_sg U12421 ( .A(\update_mask_0/reg_out[15][19] ), .B(n6445), .X(n5594) );
  nand_x1_sg U12422 ( .A(\i_im[15][18] ), .B(n6261), .X(n5591) );
  nand_x1_sg U12423 ( .A(\update_mask_0/reg_out[15][18] ), .B(n7044), .X(n5592) );
  nand_x1_sg U12424 ( .A(\i_im[15][17] ), .B(n7367), .X(n5589) );
  nand_x1_sg U12425 ( .A(\update_mask_0/reg_out[15][17] ), .B(n7043), .X(n5590) );
  nand_x1_sg U12426 ( .A(\i_im[15][16] ), .B(n6522), .X(n5587) );
  nand_x1_sg U12427 ( .A(\update_mask_0/reg_out[15][16] ), .B(n5996), .X(n5588) );
  nand_x1_sg U12428 ( .A(\i_im[15][15] ), .B(n6258), .X(n5585) );
  nand_x1_sg U12429 ( .A(\update_mask_0/reg_out[15][15] ), .B(n6268), .X(n5586) );
  nand_x1_sg U12430 ( .A(\i_im[15][14] ), .B(n6259), .X(n5583) );
  nand_x1_sg U12431 ( .A(\update_mask_0/reg_out[15][14] ), .B(n6268), .X(n5584) );
  nand_x1_sg U12432 ( .A(\i_im[15][13] ), .B(n6534), .X(n5581) );
  nand_x1_sg U12433 ( .A(\update_mask_0/reg_out[15][13] ), .B(n6452), .X(n5582) );
  nand_x1_sg U12434 ( .A(\i_im[15][12] ), .B(n7366), .X(n5579) );
  nand_x1_sg U12435 ( .A(\update_mask_0/reg_out[15][12] ), .B(n7029), .X(n5580) );
  nand_x1_sg U12436 ( .A(\i_im[15][11] ), .B(n7349), .X(n5577) );
  nand_x1_sg U12437 ( .A(\update_mask_0/reg_out[15][11] ), .B(n7335), .X(n5578) );
  nand_x1_sg U12438 ( .A(\i_im[15][10] ), .B(n6544), .X(n5575) );
  nand_x1_sg U12439 ( .A(\update_mask_0/reg_out[15][10] ), .B(n6286), .X(n5576) );
  nand_x1_sg U12440 ( .A(\i_im[15][9] ), .B(n6259), .X(n5573) );
  nand_x1_sg U12441 ( .A(\update_mask_0/reg_out[15][9] ), .B(n7325), .X(n5574)
         );
  nand_x1_sg U12442 ( .A(\i_im[15][8] ), .B(n7354), .X(n5571) );
  nand_x1_sg U12443 ( .A(\update_mask_0/reg_out[15][8] ), .B(n6454), .X(n5572)
         );
  nand_x1_sg U12444 ( .A(\i_im[15][7] ), .B(n6546), .X(n5569) );
  nand_x1_sg U12445 ( .A(\update_mask_0/reg_out[15][7] ), .B(n7029), .X(n5570)
         );
  nand_x1_sg U12446 ( .A(\i_im[15][6] ), .B(n6515), .X(n5567) );
  nand_x1_sg U12447 ( .A(\update_mask_0/reg_out[15][6] ), .B(n6271), .X(n5568)
         );
  nand_x1_sg U12448 ( .A(\i_im[15][5] ), .B(n6532), .X(n5565) );
  nand_x1_sg U12449 ( .A(\update_mask_0/reg_out[15][5] ), .B(n7047), .X(n5566)
         );
  nand_x1_sg U12450 ( .A(\i_im[15][4] ), .B(n6547), .X(n5563) );
  nand_x1_sg U12451 ( .A(\update_mask_0/reg_out[15][4] ), .B(n5989), .X(n5564)
         );
  nand_x1_sg U12452 ( .A(\i_im[15][3] ), .B(n6305), .X(n5561) );
  nand_x1_sg U12453 ( .A(\update_mask_0/reg_out[15][3] ), .B(n7021), .X(n5562)
         );
  nand_x1_sg U12454 ( .A(\i_im[15][2] ), .B(n6090), .X(n5559) );
  nand_x1_sg U12455 ( .A(\update_mask_0/reg_out[15][2] ), .B(n7046), .X(n5560)
         );
  nand_x1_sg U12456 ( .A(\i_im[15][1] ), .B(n7365), .X(n5557) );
  nand_x1_sg U12457 ( .A(\update_mask_0/reg_out[15][1] ), .B(n7331), .X(n5558)
         );
  nand_x1_sg U12458 ( .A(\i_im[15][0] ), .B(n6306), .X(n5555) );
  nand_x1_sg U12459 ( .A(\update_mask_0/reg_out[15][0] ), .B(n5997), .X(n5556)
         );
  nand_x1_sg U12460 ( .A(\i_im[14][19] ), .B(n6257), .X(n5553) );
  nand_x1_sg U12461 ( .A(\update_mask_0/reg_out[14][19] ), .B(n7028), .X(n5554) );
  nand_x1_sg U12462 ( .A(\i_im[14][18] ), .B(n6254), .X(n5551) );
  nand_x1_sg U12463 ( .A(\update_mask_0/reg_out[14][18] ), .B(n7049), .X(n5552) );
  nand_x1_sg U12464 ( .A(\i_im[14][17] ), .B(n6517), .X(n5549) );
  nand_x1_sg U12465 ( .A(\update_mask_0/reg_out[14][17] ), .B(n5995), .X(n5550) );
  nand_x1_sg U12466 ( .A(\i_im[14][16] ), .B(n6518), .X(n5547) );
  nand_x1_sg U12467 ( .A(\update_mask_0/reg_out[14][16] ), .B(n6453), .X(n5548) );
  nand_x1_sg U12468 ( .A(\i_im[14][15] ), .B(n6519), .X(n5545) );
  nand_x1_sg U12469 ( .A(\update_mask_0/reg_out[14][15] ), .B(n6292), .X(n5546) );
  nand_x1_sg U12470 ( .A(\i_im[14][14] ), .B(n6525), .X(n5543) );
  nand_x1_sg U12471 ( .A(\update_mask_0/reg_out[14][14] ), .B(n7029), .X(n5544) );
  nand_x1_sg U12472 ( .A(\i_im[14][13] ), .B(n7340), .X(n5541) );
  nand_x1_sg U12473 ( .A(\update_mask_0/reg_out[14][13] ), .B(n7027), .X(n5542) );
  nand_x1_sg U12474 ( .A(\i_im[14][12] ), .B(n6520), .X(n5539) );
  nand_x1_sg U12475 ( .A(\update_mask_0/reg_out[14][12] ), .B(n7333), .X(n5540) );
  nand_x1_sg U12476 ( .A(\i_im[14][11] ), .B(n6085), .X(n5537) );
  nand_x1_sg U12477 ( .A(\update_mask_0/reg_out[14][11] ), .B(n7045), .X(n5538) );
  nand_x1_sg U12478 ( .A(\i_im[14][10] ), .B(n7351), .X(n5535) );
  nand_x1_sg U12479 ( .A(\update_mask_0/reg_out[14][10] ), .B(n6449), .X(n5536) );
  nand_x1_sg U12480 ( .A(\i_im[14][9] ), .B(n7367), .X(n5533) );
  nand_x1_sg U12481 ( .A(\update_mask_0/reg_out[14][9] ), .B(n7047), .X(n5534)
         );
  nand_x1_sg U12482 ( .A(\i_im[14][8] ), .B(n6466), .X(n5531) );
  nand_x1_sg U12483 ( .A(\update_mask_0/reg_out[14][8] ), .B(n6282), .X(n5532)
         );
  nand_x1_sg U12484 ( .A(\i_im[14][7] ), .B(n7372), .X(n5529) );
  nand_x1_sg U12485 ( .A(\update_mask_0/reg_out[14][7] ), .B(n6292), .X(n5530)
         );
  nand_x1_sg U12486 ( .A(\i_im[14][6] ), .B(n6247), .X(n5527) );
  nand_x1_sg U12487 ( .A(\update_mask_0/reg_out[14][6] ), .B(n6456), .X(n5528)
         );
  nand_x1_sg U12488 ( .A(\i_im[14][5] ), .B(n6529), .X(n5525) );
  nand_x1_sg U12489 ( .A(\update_mask_0/reg_out[14][5] ), .B(n6445), .X(n5526)
         );
  nand_x1_sg U12490 ( .A(\i_im[14][4] ), .B(n6085), .X(n5523) );
  nand_x1_sg U12491 ( .A(\update_mask_0/reg_out[14][4] ), .B(n6447), .X(n5524)
         );
  nand_x1_sg U12492 ( .A(\i_im[14][3] ), .B(n6525), .X(n5521) );
  nand_x1_sg U12493 ( .A(\update_mask_0/reg_out[14][3] ), .B(n5993), .X(n5522)
         );
  nand_x1_sg U12494 ( .A(\i_im[14][2] ), .B(n7345), .X(n5519) );
  nand_x1_sg U12495 ( .A(\update_mask_0/reg_out[14][2] ), .B(n7021), .X(n5520)
         );
  nand_x1_sg U12496 ( .A(\i_im[14][1] ), .B(n7354), .X(n5517) );
  nand_x1_sg U12497 ( .A(\update_mask_0/reg_out[14][1] ), .B(n5986), .X(n5518)
         );
  nand_x1_sg U12498 ( .A(\i_im[14][0] ), .B(n7362), .X(n5515) );
  nand_x1_sg U12499 ( .A(\update_mask_0/reg_out[14][0] ), .B(n7042), .X(n5516)
         );
  nand_x1_sg U12500 ( .A(\i_im[13][19] ), .B(n6092), .X(n5513) );
  nand_x1_sg U12501 ( .A(\update_mask_0/reg_out[13][19] ), .B(n5994), .X(n5514) );
  nand_x1_sg U12502 ( .A(\i_im[13][18] ), .B(n6253), .X(n5511) );
  nand_x1_sg U12503 ( .A(\update_mask_0/reg_out[13][18] ), .B(n7045), .X(n5512) );
  nand_x1_sg U12504 ( .A(\i_im[13][17] ), .B(n6518), .X(n5509) );
  nand_x1_sg U12505 ( .A(\update_mask_0/reg_out[13][17] ), .B(n6448), .X(n5510) );
  nand_x1_sg U12506 ( .A(\i_im[13][16] ), .B(n7347), .X(n5507) );
  nand_x1_sg U12507 ( .A(\update_mask_0/reg_out[13][16] ), .B(n5993), .X(n5508) );
  nand_x1_sg U12508 ( .A(\i_im[13][15] ), .B(n6301), .X(n5505) );
  nand_x1_sg U12509 ( .A(\update_mask_0/reg_out[13][15] ), .B(n7330), .X(n5506) );
  nand_x1_sg U12510 ( .A(\i_im[13][14] ), .B(n7350), .X(n5503) );
  nand_x1_sg U12511 ( .A(\update_mask_0/reg_out[13][14] ), .B(n7043), .X(n5504) );
  nand_x1_sg U12512 ( .A(\i_im[13][13] ), .B(n6535), .X(n5501) );
  nand_x1_sg U12513 ( .A(\update_mask_0/reg_out[13][13] ), .B(n7030), .X(n5502) );
  nand_x1_sg U12514 ( .A(\i_im[13][12] ), .B(n7344), .X(n5499) );
  nand_x1_sg U12515 ( .A(\update_mask_0/reg_out[13][12] ), .B(n6154), .X(n5500) );
  nand_x1_sg U12516 ( .A(\i_im[13][11] ), .B(n7354), .X(n5497) );
  nand_x1_sg U12517 ( .A(\update_mask_0/reg_out[13][11] ), .B(n7041), .X(n5498) );
  nand_x1_sg U12518 ( .A(\i_im[13][10] ), .B(n6523), .X(n5495) );
  nand_x1_sg U12519 ( .A(\update_mask_0/reg_out[13][10] ), .B(n7035), .X(n5496) );
  nand_x1_sg U12520 ( .A(\i_im[13][9] ), .B(n6528), .X(n5493) );
  nand_x1_sg U12521 ( .A(\update_mask_0/reg_out[13][9] ), .B(n6281), .X(n5494)
         );
  nand_x1_sg U12522 ( .A(\i_im[13][8] ), .B(n6092), .X(n5491) );
  nand_x1_sg U12523 ( .A(\update_mask_0/reg_out[13][8] ), .B(n6291), .X(n5492)
         );
  nand_x1_sg U12524 ( .A(\i_im[13][7] ), .B(n6295), .X(n5489) );
  nand_x1_sg U12525 ( .A(\update_mask_0/reg_out[13][7] ), .B(n6143), .X(n5490)
         );
  nand_x1_sg U12526 ( .A(\i_im[13][6] ), .B(n6466), .X(n5487) );
  nand_x1_sg U12527 ( .A(\update_mask_0/reg_out[13][6] ), .B(n7326), .X(n5488)
         );
  nand_x1_sg U12528 ( .A(\i_im[13][5] ), .B(n6545), .X(n5485) );
  nand_x1_sg U12529 ( .A(\update_mask_0/reg_out[13][5] ), .B(n7021), .X(n5486)
         );
  nand_x1_sg U12530 ( .A(\i_im[13][4] ), .B(n7344), .X(n5483) );
  nand_x1_sg U12531 ( .A(\update_mask_0/reg_out[13][4] ), .B(n7050), .X(n5484)
         );
  nand_x1_sg U12532 ( .A(\i_im[13][3] ), .B(n7347), .X(n5481) );
  nand_x1_sg U12533 ( .A(\update_mask_0/reg_out[13][3] ), .B(n7022), .X(n5482)
         );
  nand_x1_sg U12534 ( .A(\i_im[13][2] ), .B(n7352), .X(n5479) );
  nand_x1_sg U12535 ( .A(\update_mask_0/reg_out[13][2] ), .B(n6445), .X(n5480)
         );
  nand_x1_sg U12536 ( .A(\i_im[13][1] ), .B(n6515), .X(n5477) );
  nand_x1_sg U12537 ( .A(\update_mask_0/reg_out[13][1] ), .B(n7334), .X(n5478)
         );
  nand_x1_sg U12538 ( .A(\i_im[13][0] ), .B(n6467), .X(n5475) );
  nand_x1_sg U12539 ( .A(\update_mask_0/reg_out[13][0] ), .B(n6267), .X(n5476)
         );
  nand_x1_sg U12540 ( .A(\i_im[12][19] ), .B(n6538), .X(n5473) );
  nand_x1_sg U12541 ( .A(\update_mask_0/reg_out[12][19] ), .B(n6358), .X(n5474) );
  nand_x1_sg U12542 ( .A(\i_im[12][18] ), .B(n7345), .X(n5471) );
  nand_x1_sg U12543 ( .A(\update_mask_0/reg_out[12][18] ), .B(n6286), .X(n5472) );
  nand_x1_sg U12544 ( .A(\i_im[12][17] ), .B(n6467), .X(n5469) );
  nand_x1_sg U12545 ( .A(\update_mask_0/reg_out[12][17] ), .B(n7038), .X(n5470) );
  nand_x1_sg U12546 ( .A(\i_im[12][16] ), .B(n7369), .X(n5467) );
  nand_x1_sg U12547 ( .A(\update_mask_0/reg_out[12][16] ), .B(n5990), .X(n5468) );
  nand_x1_sg U12548 ( .A(\i_im[12][15] ), .B(n6523), .X(n5465) );
  nand_x1_sg U12549 ( .A(\update_mask_0/reg_out[12][15] ), .B(n6281), .X(n5466) );
  nand_x1_sg U12550 ( .A(\i_im[12][14] ), .B(n7368), .X(n5463) );
  nand_x1_sg U12551 ( .A(\update_mask_0/reg_out[12][14] ), .B(n6451), .X(n5464) );
  nand_x1_sg U12552 ( .A(\i_im[12][13] ), .B(n7341), .X(n5461) );
  nand_x1_sg U12553 ( .A(\update_mask_0/reg_out[12][13] ), .B(n6145), .X(n5462) );
  nand_x1_sg U12554 ( .A(\i_im[12][12] ), .B(n7372), .X(n5459) );
  nand_x1_sg U12555 ( .A(\update_mask_0/reg_out[12][12] ), .B(n6446), .X(n5460) );
  nand_x1_sg U12556 ( .A(\i_im[12][11] ), .B(n7371), .X(n5457) );
  nand_x1_sg U12557 ( .A(\update_mask_0/reg_out[12][11] ), .B(n7033), .X(n5458) );
  nand_x1_sg U12558 ( .A(\i_im[12][10] ), .B(n6085), .X(n5455) );
  nand_x1_sg U12559 ( .A(\update_mask_0/reg_out[12][10] ), .B(n7046), .X(n5456) );
  nand_x1_sg U12560 ( .A(\i_im[12][9] ), .B(n6536), .X(n5453) );
  nand_x1_sg U12561 ( .A(\update_mask_0/reg_out[12][9] ), .B(n7024), .X(n5454)
         );
  nand_x1_sg U12562 ( .A(\i_im[12][8] ), .B(n7371), .X(n5451) );
  nand_x1_sg U12563 ( .A(\update_mask_0/reg_out[12][8] ), .B(n7034), .X(n5452)
         );
  nand_x1_sg U12564 ( .A(\i_im[12][7] ), .B(n6294), .X(n5449) );
  nand_x1_sg U12565 ( .A(\update_mask_0/reg_out[12][7] ), .B(n7026), .X(n5450)
         );
  nand_x1_sg U12566 ( .A(\i_im[12][6] ), .B(n7343), .X(n5447) );
  nand_x1_sg U12567 ( .A(\update_mask_0/reg_out[12][6] ), .B(n7028), .X(n5448)
         );
  nand_x1_sg U12568 ( .A(\i_im[12][5] ), .B(n7370), .X(n5445) );
  nand_x1_sg U12569 ( .A(\update_mask_0/reg_out[12][5] ), .B(n6358), .X(n5446)
         );
  nand_x1_sg U12570 ( .A(\i_im[12][4] ), .B(n7366), .X(n5443) );
  nand_x1_sg U12571 ( .A(\update_mask_0/reg_out[12][4] ), .B(n7050), .X(n5444)
         );
  nand_x1_sg U12572 ( .A(\i_im[12][3] ), .B(n6255), .X(n5441) );
  nand_x1_sg U12573 ( .A(\update_mask_0/reg_out[12][3] ), .B(n7039), .X(n5442)
         );
  nand_x1_sg U12574 ( .A(\i_im[12][2] ), .B(n6298), .X(n5439) );
  nand_x1_sg U12575 ( .A(\update_mask_0/reg_out[12][2] ), .B(n7331), .X(n5440)
         );
  nand_x1_sg U12576 ( .A(\i_im[12][1] ), .B(n7367), .X(n5437) );
  nand_x1_sg U12577 ( .A(\update_mask_0/reg_out[12][1] ), .B(n7051), .X(n5438)
         );
  nand_x1_sg U12578 ( .A(\i_im[12][0] ), .B(n6301), .X(n5435) );
  nand_x1_sg U12579 ( .A(\update_mask_0/reg_out[12][0] ), .B(n6146), .X(n5436)
         );
  nand_x1_sg U12580 ( .A(\i_im[11][19] ), .B(n6247), .X(n5433) );
  nand_x1_sg U12581 ( .A(\update_mask_0/reg_out[11][19] ), .B(n7040), .X(n5434) );
  nand_x1_sg U12582 ( .A(\i_im[11][18] ), .B(n7358), .X(n5431) );
  nand_x1_sg U12583 ( .A(\update_mask_0/reg_out[11][18] ), .B(n6151), .X(n5432) );
  nand_x1_sg U12584 ( .A(\i_im[11][17] ), .B(n7362), .X(n5429) );
  nand_x1_sg U12585 ( .A(\update_mask_0/reg_out[11][17] ), .B(n6282), .X(n5430) );
  nand_x1_sg U12586 ( .A(\i_im[11][16] ), .B(n6256), .X(n5427) );
  nand_x1_sg U12587 ( .A(\update_mask_0/reg_out[11][16] ), .B(n7329), .X(n5428) );
  nand_x1_sg U12588 ( .A(\i_im[11][15] ), .B(n7346), .X(n5425) );
  nand_x1_sg U12589 ( .A(\update_mask_0/reg_out[11][15] ), .B(n5997), .X(n5426) );
  nand_x1_sg U12590 ( .A(\i_im[11][14] ), .B(n7370), .X(n5423) );
  nand_x1_sg U12591 ( .A(\update_mask_0/reg_out[11][14] ), .B(n7031), .X(n5424) );
  nand_x1_sg U12592 ( .A(\i_im[11][13] ), .B(n6297), .X(n5421) );
  nand_x1_sg U12593 ( .A(\update_mask_0/reg_out[11][13] ), .B(n6156), .X(n5422) );
  nand_x1_sg U12594 ( .A(\i_im[11][12] ), .B(n6088), .X(n5419) );
  nand_x1_sg U12595 ( .A(\update_mask_0/reg_out[11][12] ), .B(n6447), .X(n5420) );
  nand_x1_sg U12596 ( .A(\i_im[11][11] ), .B(n6466), .X(n5417) );
  nand_x1_sg U12597 ( .A(\update_mask_0/reg_out[11][11] ), .B(n6453), .X(n5418) );
  nand_x1_sg U12598 ( .A(\i_im[11][10] ), .B(n6522), .X(n5415) );
  nand_x1_sg U12599 ( .A(\update_mask_0/reg_out[11][10] ), .B(n7045), .X(n5416) );
  nand_x1_sg U12600 ( .A(\i_im[11][1] ), .B(n6537), .X(n5397) );
  nand_x1_sg U12601 ( .A(\update_mask_0/reg_out[11][1] ), .B(n7022), .X(n5398)
         );
  nand_x1_sg U12602 ( .A(\i_im[11][0] ), .B(n7365), .X(n5395) );
  nand_x1_sg U12603 ( .A(\update_mask_0/reg_out[11][0] ), .B(n6451), .X(n5396)
         );
  nand_x1_sg U12604 ( .A(\i_im[10][19] ), .B(n6092), .X(n5393) );
  nand_x1_sg U12605 ( .A(\update_mask_0/reg_out[10][19] ), .B(n6445), .X(n5394) );
  nand_x1_sg U12606 ( .A(\i_im[10][18] ), .B(n7372), .X(n5391) );
  nand_x1_sg U12607 ( .A(\update_mask_0/reg_out[10][18] ), .B(n7046), .X(n5392) );
  nand_x1_sg U12608 ( .A(\i_im[10][17] ), .B(n6248), .X(n5389) );
  nand_x1_sg U12609 ( .A(\update_mask_0/reg_out[10][17] ), .B(n7020), .X(n5390) );
  nand_x1_sg U12610 ( .A(\i_im[10][16] ), .B(n6524), .X(n5387) );
  nand_x1_sg U12611 ( .A(\update_mask_0/reg_out[10][16] ), .B(n6277), .X(n5388) );
  nand_x1_sg U12612 ( .A(\i_im[10][15] ), .B(n6463), .X(n5385) );
  nand_x1_sg U12613 ( .A(\update_mask_0/reg_out[10][15] ), .B(n7034), .X(n5386) );
  nand_x1_sg U12614 ( .A(\i_im[10][14] ), .B(n6536), .X(n5383) );
  nand_x1_sg U12615 ( .A(\update_mask_0/reg_out[10][14] ), .B(n6358), .X(n5384) );
  nand_x1_sg U12616 ( .A(\i_im[10][13] ), .B(n6537), .X(n5381) );
  nand_x1_sg U12617 ( .A(\update_mask_0/reg_out[10][13] ), .B(n6455), .X(n5382) );
  nand_x1_sg U12618 ( .A(\i_im[10][12] ), .B(n6297), .X(n5379) );
  nand_x1_sg U12619 ( .A(\update_mask_0/reg_out[10][12] ), .B(n6449), .X(n5380) );
  nand_x1_sg U12620 ( .A(\i_im[10][11] ), .B(n7360), .X(n5377) );
  nand_x1_sg U12621 ( .A(\update_mask_0/reg_out[10][11] ), .B(n6272), .X(n5378) );
  nand_x1_sg U12622 ( .A(\i_im[10][10] ), .B(n7366), .X(n5375) );
  nand_x1_sg U12623 ( .A(\update_mask_0/reg_out[10][10] ), .B(n6148), .X(n5376) );
  nand_x1_sg U12624 ( .A(\i_im[10][9] ), .B(n6517), .X(n5373) );
  nand_x1_sg U12625 ( .A(\update_mask_0/reg_out[10][9] ), .B(n6148), .X(n5374)
         );
  nand_x1_sg U12626 ( .A(\i_im[10][8] ), .B(n6088), .X(n5371) );
  nand_x1_sg U12627 ( .A(\update_mask_0/reg_out[10][8] ), .B(n7041), .X(n5372)
         );
  nand_x1_sg U12628 ( .A(\i_im[10][7] ), .B(n6293), .X(n5369) );
  nand_x1_sg U12629 ( .A(\update_mask_0/reg_out[10][7] ), .B(n6355), .X(n5370)
         );
  nand_x1_sg U12630 ( .A(\i_im[10][6] ), .B(n6522), .X(n5367) );
  nand_x1_sg U12631 ( .A(\update_mask_0/reg_out[10][6] ), .B(n6156), .X(n5368)
         );
  nand_x1_sg U12632 ( .A(\i_im[10][5] ), .B(n7349), .X(n5365) );
  nand_x1_sg U12633 ( .A(\update_mask_0/reg_out[10][5] ), .B(n6358), .X(n5366)
         );
  nand_x1_sg U12634 ( .A(\i_im[10][4] ), .B(n6305), .X(n5363) );
  nand_x1_sg U12635 ( .A(\update_mask_0/reg_out[10][4] ), .B(n6452), .X(n5364)
         );
  nand_x1_sg U12636 ( .A(\i_im[10][3] ), .B(n6529), .X(n5361) );
  nand_x1_sg U12637 ( .A(\update_mask_0/reg_out[10][3] ), .B(n6271), .X(n5362)
         );
  nand_x1_sg U12638 ( .A(\i_im[10][2] ), .B(n6529), .X(n5359) );
  nand_x1_sg U12639 ( .A(\update_mask_0/reg_out[10][2] ), .B(n6357), .X(n5360)
         );
  nand_x1_sg U12640 ( .A(\i_im[10][1] ), .B(n6306), .X(n5357) );
  nand_x1_sg U12641 ( .A(\update_mask_0/reg_out[10][1] ), .B(n7051), .X(n5358)
         );
  nand_x1_sg U12642 ( .A(\i_im[10][0] ), .B(n6519), .X(n5355) );
  nand_x1_sg U12643 ( .A(\update_mask_0/reg_out[10][0] ), .B(n7030), .X(n5356)
         );
  nand_x1_sg U12644 ( .A(\i_im[9][19] ), .B(n7342), .X(n5353) );
  nand_x1_sg U12645 ( .A(\update_mask_0/reg_out[9][19] ), .B(n6148), .X(n5354)
         );
  nand_x1_sg U12646 ( .A(\i_im[9][18] ), .B(n6530), .X(n5351) );
  nand_x1_sg U12647 ( .A(\update_mask_0/reg_out[9][18] ), .B(n6268), .X(n5352)
         );
  nand_x1_sg U12648 ( .A(\i_im[9][17] ), .B(n6538), .X(n5349) );
  nand_x1_sg U12649 ( .A(\update_mask_0/reg_out[9][17] ), .B(n7029), .X(n5350)
         );
  nand_x1_sg U12650 ( .A(\i_im[9][16] ), .B(n6467), .X(n5347) );
  nand_x1_sg U12651 ( .A(\update_mask_0/reg_out[9][16] ), .B(n5988), .X(n5348)
         );
  nand_x1_sg U12652 ( .A(\i_im[9][15] ), .B(n6536), .X(n5345) );
  nand_x1_sg U12653 ( .A(\update_mask_0/reg_out[9][15] ), .B(n7325), .X(n5346)
         );
  nand_x1_sg U12654 ( .A(\i_im[9][14] ), .B(n7349), .X(n5343) );
  nand_x1_sg U12655 ( .A(\update_mask_0/reg_out[9][14] ), .B(n6272), .X(n5344)
         );
  nand_x1_sg U12656 ( .A(\i_im[9][13] ), .B(n6306), .X(n5341) );
  nand_x1_sg U12657 ( .A(\update_mask_0/reg_out[9][13] ), .B(n6357), .X(n5342)
         );
  nand_x1_sg U12658 ( .A(\i_im[9][12] ), .B(n7346), .X(n5339) );
  nand_x1_sg U12659 ( .A(\update_mask_0/reg_out[9][12] ), .B(n6456), .X(n5340)
         );
  nand_x1_sg U12660 ( .A(\i_im[9][11] ), .B(n6521), .X(n5337) );
  nand_x1_sg U12661 ( .A(\update_mask_0/reg_out[9][11] ), .B(n6360), .X(n5338)
         );
  nand_x1_sg U12662 ( .A(\i_im[9][10] ), .B(n6464), .X(n5335) );
  nand_x1_sg U12663 ( .A(\update_mask_0/reg_out[9][10] ), .B(n6359), .X(n5336)
         );
  nand_x1_sg U12664 ( .A(\i_im[9][9] ), .B(n6260), .X(n5333) );
  nand_x1_sg U12665 ( .A(\update_mask_0/reg_out[9][9] ), .B(n6150), .X(n5334)
         );
  nand_x1_sg U12666 ( .A(\i_im[9][8] ), .B(n7346), .X(n5331) );
  nand_x1_sg U12667 ( .A(\update_mask_0/reg_out[9][8] ), .B(n5988), .X(n5332)
         );
  nand_x1_sg U12668 ( .A(\i_im[9][7] ), .B(n6538), .X(n5329) );
  nand_x1_sg U12669 ( .A(\update_mask_0/reg_out[9][7] ), .B(n6357), .X(n5330)
         );
  nand_x1_sg U12670 ( .A(\i_im[9][6] ), .B(n7359), .X(n5327) );
  nand_x1_sg U12671 ( .A(\update_mask_0/reg_out[9][6] ), .B(n6145), .X(n5328)
         );
  nand_x1_sg U12672 ( .A(\i_im[9][5] ), .B(n6296), .X(n5325) );
  nand_x1_sg U12673 ( .A(\update_mask_0/reg_out[9][5] ), .B(n6356), .X(n5326)
         );
  nand_x1_sg U12674 ( .A(\i_im[9][4] ), .B(n6524), .X(n5323) );
  nand_x1_sg U12675 ( .A(\update_mask_0/reg_out[9][4] ), .B(n7333), .X(n5324)
         );
  nand_x1_sg U12676 ( .A(\i_im[9][3] ), .B(n7365), .X(n5321) );
  nand_x1_sg U12677 ( .A(\update_mask_0/reg_out[9][3] ), .B(n5992), .X(n5322)
         );
  nand_x1_sg U12678 ( .A(\i_im[9][2] ), .B(n7342), .X(n5319) );
  nand_x1_sg U12679 ( .A(\update_mask_0/reg_out[9][2] ), .B(n5991), .X(n5320)
         );
  nand_x1_sg U12680 ( .A(\i_im[9][1] ), .B(n6085), .X(n5317) );
  nand_x1_sg U12681 ( .A(\update_mask_0/reg_out[9][1] ), .B(n7023), .X(n5318)
         );
  nand_x1_sg U12682 ( .A(\i_im[9][0] ), .B(n7352), .X(n5315) );
  nand_x1_sg U12683 ( .A(\update_mask_0/reg_out[9][0] ), .B(n6143), .X(n5316)
         );
  nand_x1_sg U12684 ( .A(\i_im[8][19] ), .B(n7360), .X(n5313) );
  nand_x1_sg U12685 ( .A(\update_mask_0/reg_out[8][19] ), .B(n6452), .X(n5314)
         );
  nand_x1_sg U12686 ( .A(\i_im[8][18] ), .B(n6521), .X(n5311) );
  nand_x1_sg U12687 ( .A(\update_mask_0/reg_out[8][18] ), .B(n6451), .X(n5312)
         );
  nand_x1_sg U12688 ( .A(\i_im[8][17] ), .B(n6547), .X(n5309) );
  nand_x1_sg U12689 ( .A(\update_mask_0/reg_out[8][17] ), .B(n5995), .X(n5310)
         );
  nand_x1_sg U12690 ( .A(\i_im[8][16] ), .B(n6254), .X(n5307) );
  nand_x1_sg U12691 ( .A(\update_mask_0/reg_out[8][16] ), .B(n7020), .X(n5308)
         );
  nand_x1_sg U12692 ( .A(\i_im[8][15] ), .B(n6295), .X(n5305) );
  nand_x1_sg U12693 ( .A(\update_mask_0/reg_out[8][15] ), .B(n7020), .X(n5306)
         );
  nand_x1_sg U12694 ( .A(\i_im[8][14] ), .B(n7352), .X(n5303) );
  nand_x1_sg U12695 ( .A(\update_mask_0/reg_out[8][14] ), .B(n6276), .X(n5304)
         );
  nand_x1_sg U12696 ( .A(\i_im[8][13] ), .B(n6294), .X(n5301) );
  nand_x1_sg U12697 ( .A(\update_mask_0/reg_out[8][13] ), .B(n7329), .X(n5302)
         );
  nand_x1_sg U12698 ( .A(\i_im[8][12] ), .B(n6538), .X(n5299) );
  nand_x1_sg U12699 ( .A(\update_mask_0/reg_out[8][12] ), .B(n6272), .X(n5300)
         );
  nand_x1_sg U12700 ( .A(\i_im[8][11] ), .B(n7370), .X(n5297) );
  nand_x1_sg U12701 ( .A(\update_mask_0/reg_out[8][11] ), .B(n7050), .X(n5298)
         );
  nand_x1_sg U12702 ( .A(\i_im[8][10] ), .B(n6528), .X(n5295) );
  nand_x1_sg U12703 ( .A(\update_mask_0/reg_out[8][10] ), .B(n7033), .X(n5296)
         );
  nand_x1_sg U12704 ( .A(\i_im[8][9] ), .B(n6305), .X(n5293) );
  nand_x1_sg U12705 ( .A(\update_mask_0/reg_out[8][9] ), .B(n5996), .X(n5294)
         );
  nand_x1_sg U12706 ( .A(\i_im[8][8] ), .B(n7362), .X(n5291) );
  nand_x1_sg U12707 ( .A(\update_mask_0/reg_out[8][8] ), .B(n6153), .X(n5292)
         );
  nand_x1_sg U12708 ( .A(\i_im[8][7] ), .B(n6301), .X(n5289) );
  nand_x1_sg U12709 ( .A(\update_mask_0/reg_out[8][7] ), .B(n7035), .X(n5290)
         );
  nand_x1_sg U12710 ( .A(\i_im[8][6] ), .B(n6293), .X(n5287) );
  nand_x1_sg U12711 ( .A(\update_mask_0/reg_out[8][6] ), .B(n5990), .X(n5288)
         );
  nand_x1_sg U12712 ( .A(\i_im[8][5] ), .B(n6248), .X(n5285) );
  nand_x1_sg U12713 ( .A(\update_mask_0/reg_out[8][5] ), .B(n7041), .X(n5286)
         );
  nand_x1_sg U12714 ( .A(\i_im[8][4] ), .B(n6258), .X(n5283) );
  nand_x1_sg U12715 ( .A(\update_mask_0/reg_out[8][4] ), .B(n7024), .X(n5284)
         );
  nand_x1_sg U12716 ( .A(\i_im[8][3] ), .B(n6248), .X(n5281) );
  nand_x1_sg U12717 ( .A(\update_mask_0/reg_out[8][3] ), .B(n5994), .X(n5282)
         );
  nand_x1_sg U12718 ( .A(\i_im[8][2] ), .B(n7370), .X(n5279) );
  nand_x1_sg U12719 ( .A(\update_mask_0/reg_out[8][2] ), .B(n6448), .X(n5280)
         );
  nand_x1_sg U12720 ( .A(\i_im[8][1] ), .B(n6526), .X(n5277) );
  nand_x1_sg U12721 ( .A(\update_mask_0/reg_out[8][1] ), .B(n5988), .X(n5278)
         );
  nand_x1_sg U12722 ( .A(\i_im[8][0] ), .B(n6298), .X(n5275) );
  nand_x1_sg U12723 ( .A(\update_mask_0/reg_out[8][0] ), .B(n6153), .X(n5276)
         );
  nand_x1_sg U12724 ( .A(\i_im[7][19] ), .B(n6521), .X(n5273) );
  nand_x1_sg U12725 ( .A(\update_mask_0/reg_out[7][19] ), .B(n7042), .X(n5274)
         );
  nand_x1_sg U12726 ( .A(\i_im[7][18] ), .B(n6293), .X(n5271) );
  nand_x1_sg U12727 ( .A(\update_mask_0/reg_out[7][18] ), .B(n5989), .X(n5272)
         );
  nand_x1_sg U12728 ( .A(\i_im[7][17] ), .B(n7371), .X(n5269) );
  nand_x1_sg U12729 ( .A(\update_mask_0/reg_out[7][17] ), .B(n6144), .X(n5270)
         );
  nand_x1_sg U12730 ( .A(\i_im[7][16] ), .B(n6464), .X(n5267) );
  nand_x1_sg U12731 ( .A(\update_mask_0/reg_out[7][16] ), .B(n6155), .X(n5268)
         );
  nand_x1_sg U12732 ( .A(\i_im[7][15] ), .B(n6468), .X(n5265) );
  nand_x1_sg U12733 ( .A(\update_mask_0/reg_out[7][15] ), .B(n7043), .X(n5266)
         );
  nand_x1_sg U12734 ( .A(\i_im[7][14] ), .B(n6530), .X(n5263) );
  nand_x1_sg U12735 ( .A(\update_mask_0/reg_out[7][14] ), .B(n5992), .X(n5264)
         );
  nand_x1_sg U12736 ( .A(\i_im[7][13] ), .B(n6514), .X(n5261) );
  nand_x1_sg U12737 ( .A(\update_mask_0/reg_out[7][13] ), .B(n6146), .X(n5262)
         );
  nand_x1_sg U12738 ( .A(\i_im[7][12] ), .B(n6249), .X(n5259) );
  nand_x1_sg U12739 ( .A(\update_mask_0/reg_out[7][12] ), .B(n5990), .X(n5260)
         );
  nand_x1_sg U12740 ( .A(\i_im[7][11] ), .B(n7364), .X(n5257) );
  nand_x1_sg U12741 ( .A(\update_mask_0/reg_out[7][11] ), .B(n6277), .X(n5258)
         );
  nand_x1_sg U12742 ( .A(\i_im[7][10] ), .B(n6262), .X(n5255) );
  nand_x1_sg U12743 ( .A(\update_mask_0/reg_out[7][10] ), .B(n6451), .X(n5256)
         );
  nand_x1_sg U12744 ( .A(\i_im[7][9] ), .B(n6515), .X(n5253) );
  nand_x1_sg U12745 ( .A(\update_mask_0/reg_out[7][9] ), .B(n6446), .X(n5254)
         );
  nand_x1_sg U12746 ( .A(\i_im[7][8] ), .B(n6544), .X(n5251) );
  nand_x1_sg U12747 ( .A(\update_mask_0/reg_out[7][8] ), .B(n7038), .X(n5252)
         );
  nand_x1_sg U12748 ( .A(\i_im[7][7] ), .B(n7343), .X(n5249) );
  nand_x1_sg U12749 ( .A(\update_mask_0/reg_out[7][7] ), .B(n7327), .X(n5250)
         );
  nand_x1_sg U12750 ( .A(\i_im[7][6] ), .B(n6260), .X(n5247) );
  nand_x1_sg U12751 ( .A(\update_mask_0/reg_out[7][6] ), .B(n6448), .X(n5248)
         );
  nand_x1_sg U12752 ( .A(\i_im[7][5] ), .B(n6259), .X(n5245) );
  nand_x1_sg U12753 ( .A(\update_mask_0/reg_out[7][5] ), .B(n6455), .X(n5246)
         );
  nand_x1_sg U12754 ( .A(\i_im[7][4] ), .B(n7345), .X(n5243) );
  nand_x1_sg U12755 ( .A(\update_mask_0/reg_out[7][4] ), .B(n7047), .X(n5244)
         );
  nand_x1_sg U12756 ( .A(\i_im[7][3] ), .B(n6247), .X(n5241) );
  nand_x1_sg U12757 ( .A(\update_mask_0/reg_out[7][3] ), .B(n7052), .X(n5242)
         );
  nand_x1_sg U12758 ( .A(\i_im[7][2] ), .B(n7348), .X(n5239) );
  nand_x1_sg U12759 ( .A(\update_mask_0/reg_out[7][2] ), .B(n6455), .X(n5240)
         );
  nand_x1_sg U12760 ( .A(\i_im[7][1] ), .B(n6254), .X(n5237) );
  nand_x1_sg U12761 ( .A(\update_mask_0/reg_out[7][1] ), .B(n6144), .X(n5238)
         );
  nand_x1_sg U12762 ( .A(\i_im[7][0] ), .B(n6531), .X(n5235) );
  nand_x1_sg U12763 ( .A(\update_mask_0/reg_out[7][0] ), .B(n7052), .X(n5236)
         );
  nand_x1_sg U12764 ( .A(\i_im[6][19] ), .B(n7361), .X(n5233) );
  nand_x1_sg U12765 ( .A(\update_mask_0/reg_out[6][19] ), .B(n6452), .X(n5234)
         );
  nand_x1_sg U12766 ( .A(\i_im[6][18] ), .B(n6250), .X(n5231) );
  nand_x1_sg U12767 ( .A(\update_mask_0/reg_out[6][18] ), .B(n7036), .X(n5232)
         );
  nand_x1_sg U12768 ( .A(\i_im[6][17] ), .B(n6256), .X(n5229) );
  nand_x1_sg U12769 ( .A(\update_mask_0/reg_out[6][17] ), .B(n6360), .X(n5230)
         );
  nand_x1_sg U12770 ( .A(\i_im[6][16] ), .B(n6531), .X(n5227) );
  nand_x1_sg U12771 ( .A(\update_mask_0/reg_out[6][16] ), .B(n7034), .X(n5228)
         );
  nand_x1_sg U12772 ( .A(\i_im[6][15] ), .B(n6544), .X(n5225) );
  nand_x1_sg U12773 ( .A(\update_mask_0/reg_out[6][15] ), .B(n7326), .X(n5226)
         );
  nand_x1_sg U12774 ( .A(\i_im[6][14] ), .B(n7358), .X(n5223) );
  nand_x1_sg U12775 ( .A(\update_mask_0/reg_out[6][14] ), .B(n7035), .X(n5224)
         );
  nand_x1_sg U12776 ( .A(\i_im[6][13] ), .B(n6306), .X(n5221) );
  nand_x1_sg U12777 ( .A(\update_mask_0/reg_out[6][13] ), .B(n7036), .X(n5222)
         );
  nand_x1_sg U12778 ( .A(\i_im[6][12] ), .B(n6248), .X(n5219) );
  nand_x1_sg U12779 ( .A(\update_mask_0/reg_out[6][12] ), .B(n6292), .X(n5220)
         );
  nand_x1_sg U12780 ( .A(\i_im[6][3] ), .B(n6531), .X(n5201) );
  nand_x1_sg U12781 ( .A(\update_mask_0/reg_out[6][3] ), .B(n7036), .X(n5202)
         );
  nand_x1_sg U12782 ( .A(\i_im[6][2] ), .B(n6298), .X(n5199) );
  nand_x1_sg U12783 ( .A(\update_mask_0/reg_out[6][2] ), .B(n5997), .X(n5200)
         );
  nand_x1_sg U12784 ( .A(\i_im[6][1] ), .B(n7345), .X(n5197) );
  nand_x1_sg U12785 ( .A(\update_mask_0/reg_out[6][1] ), .B(n7031), .X(n5198)
         );
  nand_x1_sg U12786 ( .A(\i_im[6][0] ), .B(n7341), .X(n5195) );
  nand_x1_sg U12787 ( .A(\update_mask_0/reg_out[6][0] ), .B(n6449), .X(n5196)
         );
  nand_x1_sg U12788 ( .A(\i_im[5][19] ), .B(n6514), .X(n5193) );
  nand_x1_sg U12789 ( .A(\update_mask_0/reg_out[5][19] ), .B(n6448), .X(n5194)
         );
  nand_x1_sg U12790 ( .A(\i_im[5][18] ), .B(n6520), .X(n5191) );
  nand_x1_sg U12791 ( .A(\update_mask_0/reg_out[5][18] ), .B(n7039), .X(n5192)
         );
  nand_x1_sg U12792 ( .A(\i_im[5][17] ), .B(n6521), .X(n5189) );
  nand_x1_sg U12793 ( .A(\update_mask_0/reg_out[5][17] ), .B(n6149), .X(n5190)
         );
  nand_x1_sg U12794 ( .A(\i_im[5][16] ), .B(n6528), .X(n5187) );
  nand_x1_sg U12795 ( .A(\update_mask_0/reg_out[5][16] ), .B(n5996), .X(n5188)
         );
  nand_x1_sg U12796 ( .A(\i_im[5][15] ), .B(n7353), .X(n5185) );
  nand_x1_sg U12797 ( .A(\update_mask_0/reg_out[5][15] ), .B(n7020), .X(n5186)
         );
  nand_x1_sg U12798 ( .A(\i_im[5][14] ), .B(n6253), .X(n5183) );
  nand_x1_sg U12799 ( .A(\update_mask_0/reg_out[5][14] ), .B(n6151), .X(n5184)
         );
  nand_x1_sg U12800 ( .A(\i_im[5][13] ), .B(n6302), .X(n5181) );
  nand_x1_sg U12801 ( .A(\update_mask_0/reg_out[5][13] ), .B(n5991), .X(n5182)
         );
  nand_x1_sg U12802 ( .A(\i_im[5][12] ), .B(n6519), .X(n5179) );
  nand_x1_sg U12803 ( .A(\update_mask_0/reg_out[5][12] ), .B(n6446), .X(n5180)
         );
  nand_x1_sg U12804 ( .A(\i_im[5][11] ), .B(n6296), .X(n5177) );
  nand_x1_sg U12805 ( .A(\update_mask_0/reg_out[5][11] ), .B(n6276), .X(n5178)
         );
  nand_x1_sg U12806 ( .A(\i_im[5][10] ), .B(n6532), .X(n5175) );
  nand_x1_sg U12807 ( .A(\update_mask_0/reg_out[5][10] ), .B(n6143), .X(n5176)
         );
  nand_x1_sg U12808 ( .A(\i_im[5][9] ), .B(n6520), .X(n5173) );
  nand_x1_sg U12809 ( .A(\update_mask_0/reg_out[5][9] ), .B(n6356), .X(n5174)
         );
  nand_x1_sg U12810 ( .A(\i_im[5][8] ), .B(n6468), .X(n5171) );
  nand_x1_sg U12811 ( .A(\update_mask_0/reg_out[5][8] ), .B(n6271), .X(n5172)
         );
  nand_x1_sg U12812 ( .A(\i_im[5][7] ), .B(n7369), .X(n5169) );
  nand_x1_sg U12813 ( .A(\update_mask_0/reg_out[5][7] ), .B(n7333), .X(n5170)
         );
  nand_x1_sg U12814 ( .A(\i_im[5][6] ), .B(n6466), .X(n5167) );
  nand_x1_sg U12815 ( .A(\update_mask_0/reg_out[5][6] ), .B(n6154), .X(n5168)
         );
  nand_x1_sg U12816 ( .A(\i_im[5][5] ), .B(n6532), .X(n5165) );
  nand_x1_sg U12817 ( .A(\update_mask_0/reg_out[5][5] ), .B(n6267), .X(n5166)
         );
  nand_x1_sg U12818 ( .A(\i_im[5][4] ), .B(n7342), .X(n5163) );
  nand_x1_sg U12819 ( .A(\update_mask_0/reg_out[5][4] ), .B(n7044), .X(n5164)
         );
  nand_x1_sg U12820 ( .A(\i_im[5][3] ), .B(n6524), .X(n5161) );
  nand_x1_sg U12821 ( .A(\update_mask_0/reg_out[5][3] ), .B(n6450), .X(n5162)
         );
  nand_x1_sg U12822 ( .A(\i_im[5][2] ), .B(n6293), .X(n5159) );
  nand_x1_sg U12823 ( .A(\update_mask_0/reg_out[5][2] ), .B(n7327), .X(n5160)
         );
  nand_x1_sg U12824 ( .A(\i_im[5][1] ), .B(n7371), .X(n5157) );
  nand_x1_sg U12825 ( .A(\update_mask_0/reg_out[5][1] ), .B(n6150), .X(n5158)
         );
  nand_x1_sg U12826 ( .A(\i_im[5][0] ), .B(n7344), .X(n5155) );
  nand_x1_sg U12827 ( .A(\update_mask_0/reg_out[5][0] ), .B(n6282), .X(n5156)
         );
  nand_x1_sg U12828 ( .A(\i_im[4][19] ), .B(n6253), .X(n5153) );
  nand_x1_sg U12829 ( .A(\update_mask_0/reg_out[4][19] ), .B(n6155), .X(n5154)
         );
  nand_x1_sg U12830 ( .A(\i_im[4][18] ), .B(n6257), .X(n5151) );
  nand_x1_sg U12831 ( .A(\update_mask_0/reg_out[4][18] ), .B(n6149), .X(n5152)
         );
  nand_x1_sg U12832 ( .A(\i_im[4][17] ), .B(n6530), .X(n5149) );
  nand_x1_sg U12833 ( .A(\update_mask_0/reg_out[4][17] ), .B(n7050), .X(n5150)
         );
  nand_x1_sg U12834 ( .A(\i_im[4][16] ), .B(n6090), .X(n5147) );
  nand_x1_sg U12835 ( .A(\update_mask_0/reg_out[4][16] ), .B(n6360), .X(n5148)
         );
  nand_x1_sg U12836 ( .A(\i_im[4][15] ), .B(n7363), .X(n5145) );
  nand_x1_sg U12837 ( .A(\update_mask_0/reg_out[4][15] ), .B(n5986), .X(n5146)
         );
  nand_x1_sg U12838 ( .A(\i_im[4][14] ), .B(n6302), .X(n5143) );
  nand_x1_sg U12839 ( .A(\update_mask_0/reg_out[4][14] ), .B(n7030), .X(n5144)
         );
  nand_x1_sg U12840 ( .A(\i_im[4][13] ), .B(n6255), .X(n5141) );
  nand_x1_sg U12841 ( .A(\update_mask_0/reg_out[4][13] ), .B(n7049), .X(n5142)
         );
  nand_x1_sg U12842 ( .A(\i_im[4][12] ), .B(n7365), .X(n5139) );
  nand_x1_sg U12843 ( .A(\update_mask_0/reg_out[4][12] ), .B(n7038), .X(n5140)
         );
  nand_x1_sg U12844 ( .A(\i_im[4][11] ), .B(n6255), .X(n5137) );
  nand_x1_sg U12845 ( .A(\update_mask_0/reg_out[4][11] ), .B(n7028), .X(n5138)
         );
  nand_x1_sg U12846 ( .A(\i_im[4][10] ), .B(n6545), .X(n5135) );
  nand_x1_sg U12847 ( .A(\update_mask_0/reg_out[4][10] ), .B(n7022), .X(n5136)
         );
  nand_x1_sg U12848 ( .A(\i_im[4][9] ), .B(n6463), .X(n5133) );
  nand_x1_sg U12849 ( .A(\update_mask_0/reg_out[4][9] ), .B(n7024), .X(n5134)
         );
  nand_x1_sg U12850 ( .A(\i_im[4][8] ), .B(n6305), .X(n5131) );
  nand_x1_sg U12851 ( .A(\update_mask_0/reg_out[4][8] ), .B(n6154), .X(n5132)
         );
  nand_x1_sg U12852 ( .A(\i_im[4][7] ), .B(n7350), .X(n5129) );
  nand_x1_sg U12853 ( .A(\update_mask_0/reg_out[4][7] ), .B(n7335), .X(n5130)
         );
  nand_x1_sg U12854 ( .A(\i_im[4][6] ), .B(n6464), .X(n5127) );
  nand_x1_sg U12855 ( .A(\update_mask_0/reg_out[4][6] ), .B(n6447), .X(n5128)
         );
  nand_x1_sg U12856 ( .A(\i_im[4][5] ), .B(n6259), .X(n5125) );
  nand_x1_sg U12857 ( .A(\update_mask_0/reg_out[4][5] ), .B(n6150), .X(n5126)
         );
  nand_x1_sg U12858 ( .A(\i_im[4][4] ), .B(n7340), .X(n5123) );
  nand_x1_sg U12859 ( .A(\update_mask_0/reg_out[4][4] ), .B(n7042), .X(n5124)
         );
  nand_x1_sg U12860 ( .A(\i_im[4][3] ), .B(n6295), .X(n5121) );
  nand_x1_sg U12861 ( .A(\update_mask_0/reg_out[4][3] ), .B(n6155), .X(n5122)
         );
  nand_x1_sg U12862 ( .A(\i_im[4][2] ), .B(n7351), .X(n5119) );
  nand_x1_sg U12863 ( .A(\update_mask_0/reg_out[4][2] ), .B(n7023), .X(n5120)
         );
  nand_x1_sg U12864 ( .A(\i_im[4][1] ), .B(n6535), .X(n5117) );
  nand_x1_sg U12865 ( .A(\update_mask_0/reg_out[4][1] ), .B(n6277), .X(n5118)
         );
  nand_x1_sg U12866 ( .A(\i_im[4][0] ), .B(n6250), .X(n5115) );
  nand_x1_sg U12867 ( .A(\update_mask_0/reg_out[4][0] ), .B(n7042), .X(n5116)
         );
  nand_x1_sg U12868 ( .A(\i_im[3][19] ), .B(n6528), .X(n5113) );
  nand_x1_sg U12869 ( .A(\update_mask_0/reg_out[3][19] ), .B(n6356), .X(n5114)
         );
  nand_x1_sg U12870 ( .A(\i_im[3][18] ), .B(n6257), .X(n5111) );
  nand_x1_sg U12871 ( .A(\update_mask_0/reg_out[3][18] ), .B(n6146), .X(n5112)
         );
  nand_x1_sg U12872 ( .A(\i_im[3][17] ), .B(n7341), .X(n5109) );
  nand_x1_sg U12873 ( .A(\update_mask_0/reg_out[3][17] ), .B(n6450), .X(n5110)
         );
  nand_x1_sg U12874 ( .A(\i_im[3][16] ), .B(n6515), .X(n5107) );
  nand_x1_sg U12875 ( .A(\update_mask_0/reg_out[3][16] ), .B(n6281), .X(n5108)
         );
  nand_x1_sg U12876 ( .A(\i_im[3][15] ), .B(n6463), .X(n5105) );
  nand_x1_sg U12877 ( .A(\update_mask_0/reg_out[3][15] ), .B(n7022), .X(n5106)
         );
  nand_x1_sg U12878 ( .A(\i_im[3][14] ), .B(n6302), .X(n5103) );
  nand_x1_sg U12879 ( .A(\update_mask_0/reg_out[3][14] ), .B(n7052), .X(n5104)
         );
  nand_x1_sg U12880 ( .A(\i_im[3][13] ), .B(n6468), .X(n5101) );
  nand_x1_sg U12881 ( .A(\update_mask_0/reg_out[3][13] ), .B(n6455), .X(n5102)
         );
  nand_x1_sg U12882 ( .A(\i_im[3][12] ), .B(n7369), .X(n5099) );
  nand_x1_sg U12883 ( .A(\update_mask_0/reg_out[3][12] ), .B(n7047), .X(n5100)
         );
  nand_x1_sg U12884 ( .A(\i_im[3][11] ), .B(n7361), .X(n5097) );
  nand_x1_sg U12885 ( .A(\update_mask_0/reg_out[3][11] ), .B(n6144), .X(n5098)
         );
  nand_x1_sg U12886 ( .A(\i_im[3][10] ), .B(n7343), .X(n5095) );
  nand_x1_sg U12887 ( .A(\update_mask_0/reg_out[3][10] ), .B(n6286), .X(n5096)
         );
  nand_x1_sg U12888 ( .A(\i_im[3][9] ), .B(n6534), .X(n5093) );
  nand_x1_sg U12889 ( .A(\update_mask_0/reg_out[3][9] ), .B(n6272), .X(n5094)
         );
  nand_x1_sg U12890 ( .A(\i_im[3][8] ), .B(n6298), .X(n5091) );
  nand_x1_sg U12891 ( .A(\update_mask_0/reg_out[3][8] ), .B(n7329), .X(n5092)
         );
  nand_x1_sg U12892 ( .A(\i_im[3][7] ), .B(n7351), .X(n5089) );
  nand_x1_sg U12893 ( .A(\update_mask_0/reg_out[3][7] ), .B(n6446), .X(n5090)
         );
  nand_x1_sg U12894 ( .A(\i_im[3][6] ), .B(n7348), .X(n5087) );
  nand_x1_sg U12895 ( .A(\update_mask_0/reg_out[3][6] ), .B(n6359), .X(n5088)
         );
  nand_x1_sg U12896 ( .A(\i_im[3][5] ), .B(n7350), .X(n5085) );
  nand_x1_sg U12897 ( .A(\update_mask_0/reg_out[3][5] ), .B(n7031), .X(n5086)
         );
  nand_x1_sg U12898 ( .A(\i_im[3][4] ), .B(n6523), .X(n5083) );
  nand_x1_sg U12899 ( .A(\update_mask_0/reg_out[3][4] ), .B(n5991), .X(n5084)
         );
  nand_x1_sg U12900 ( .A(\i_im[3][3] ), .B(n7353), .X(n5081) );
  nand_x1_sg U12901 ( .A(\update_mask_0/reg_out[3][3] ), .B(n7025), .X(n5082)
         );
  nand_x1_sg U12902 ( .A(\i_im[3][2] ), .B(n7363), .X(n5079) );
  nand_x1_sg U12903 ( .A(\update_mask_0/reg_out[3][2] ), .B(n7335), .X(n5080)
         );
  nand_x1_sg U12904 ( .A(\i_im[3][1] ), .B(n6302), .X(n5077) );
  nand_x1_sg U12905 ( .A(\update_mask_0/reg_out[3][1] ), .B(n6454), .X(n5078)
         );
  nand_x1_sg U12906 ( .A(\i_im[3][0] ), .B(n6518), .X(n5075) );
  nand_x1_sg U12907 ( .A(\update_mask_0/reg_out[3][0] ), .B(n6153), .X(n5076)
         );
  nand_x1_sg U12908 ( .A(\i_im[2][19] ), .B(n6297), .X(n5073) );
  nand_x1_sg U12909 ( .A(\update_mask_0/reg_out[2][19] ), .B(n7026), .X(n5074)
         );
  nand_x1_sg U12910 ( .A(\i_im[2][18] ), .B(n6258), .X(n5071) );
  nand_x1_sg U12911 ( .A(\update_mask_0/reg_out[2][18] ), .B(n6453), .X(n5072)
         );
  nand_x1_sg U12912 ( .A(\i_im[2][17] ), .B(n7359), .X(n5069) );
  nand_x1_sg U12913 ( .A(\update_mask_0/reg_out[2][17] ), .B(n7027), .X(n5070)
         );
  nand_x1_sg U12914 ( .A(\i_im[2][16] ), .B(n7360), .X(n5067) );
  nand_x1_sg U12915 ( .A(\update_mask_0/reg_out[2][16] ), .B(n6291), .X(n5068)
         );
  nand_x1_sg U12916 ( .A(\i_im[2][15] ), .B(n6247), .X(n5065) );
  nand_x1_sg U12917 ( .A(\update_mask_0/reg_out[2][15] ), .B(n6276), .X(n5066)
         );
  nand_x1_sg U12918 ( .A(\i_im[2][14] ), .B(n6520), .X(n5063) );
  nand_x1_sg U12919 ( .A(\update_mask_0/reg_out[2][14] ), .B(n6151), .X(n5064)
         );
  nand_x1_sg U12920 ( .A(\i_im[2][13] ), .B(n6249), .X(n5061) );
  nand_x1_sg U12921 ( .A(\update_mask_0/reg_out[2][13] ), .B(n6156), .X(n5062)
         );
  nand_x1_sg U12922 ( .A(\i_im[2][12] ), .B(n6517), .X(n5059) );
  nand_x1_sg U12923 ( .A(\update_mask_0/reg_out[2][12] ), .B(n7030), .X(n5060)
         );
  nand_x1_sg U12924 ( .A(\i_im[2][11] ), .B(n7340), .X(n5057) );
  nand_x1_sg U12925 ( .A(\update_mask_0/reg_out[2][11] ), .B(n7051), .X(n5058)
         );
  nand_x1_sg U12926 ( .A(\i_im[2][10] ), .B(n6256), .X(n5055) );
  nand_x1_sg U12927 ( .A(\update_mask_0/reg_out[2][10] ), .B(n6292), .X(n5056)
         );
  nand_x1_sg U12928 ( .A(\i_im[2][9] ), .B(n6261), .X(n5053) );
  nand_x1_sg U12929 ( .A(\update_mask_0/reg_out[2][9] ), .B(n7046), .X(n5054)
         );
  nand_x1_sg U12930 ( .A(\i_im[2][8] ), .B(n7360), .X(n5051) );
  nand_x1_sg U12931 ( .A(\update_mask_0/reg_out[2][8] ), .B(n5986), .X(n5052)
         );
  nand_x1_sg U12932 ( .A(\i_im[2][7] ), .B(n6260), .X(n5049) );
  nand_x1_sg U12933 ( .A(\update_mask_0/reg_out[2][7] ), .B(n7052), .X(n5050)
         );
  nand_x1_sg U12934 ( .A(\i_im[2][6] ), .B(n7359), .X(n5047) );
  nand_x1_sg U12935 ( .A(\update_mask_0/reg_out[2][6] ), .B(n5986), .X(n5048)
         );
  nand_x1_sg U12936 ( .A(\i_im[2][5] ), .B(n6088), .X(n5045) );
  nand_x1_sg U12937 ( .A(\update_mask_0/reg_out[2][5] ), .B(n7034), .X(n5046)
         );
  nand_x1_sg U12938 ( .A(\i_im[2][4] ), .B(n6535), .X(n5043) );
  nand_x1_sg U12939 ( .A(\update_mask_0/reg_out[2][4] ), .B(n6355), .X(n5044)
         );
  nand_x1_sg U12940 ( .A(\i_im[2][3] ), .B(n6464), .X(n5041) );
  nand_x1_sg U12941 ( .A(\update_mask_0/reg_out[2][3] ), .B(n6287), .X(n5042)
         );
  nand_x1_sg U12942 ( .A(\i_im[2][2] ), .B(n7350), .X(n5039) );
  nand_x1_sg U12943 ( .A(\update_mask_0/reg_out[2][2] ), .B(n7331), .X(n5040)
         );
  nand_x1_sg U12944 ( .A(\i_im[2][1] ), .B(n6518), .X(n5037) );
  nand_x1_sg U12945 ( .A(\update_mask_0/reg_out[2][1] ), .B(n7040), .X(n5038)
         );
  nand_x1_sg U12946 ( .A(\i_im[2][0] ), .B(n7344), .X(n5035) );
  nand_x1_sg U12947 ( .A(\update_mask_0/reg_out[2][0] ), .B(n5987), .X(n5036)
         );
  nand_x1_sg U12948 ( .A(\i_im[1][19] ), .B(n6262), .X(n5033) );
  nand_x1_sg U12949 ( .A(\update_mask_0/reg_out[1][19] ), .B(n7049), .X(n5034)
         );
  nand_x1_sg U12950 ( .A(\i_im[1][18] ), .B(n6294), .X(n5031) );
  nand_x1_sg U12951 ( .A(\update_mask_0/reg_out[1][18] ), .B(n7335), .X(n5032)
         );
  nand_x1_sg U12952 ( .A(\update_mask_0/reg_out[1][17] ), .B(n6287), .X(n5030)
         );
  nand_x1_sg U12953 ( .A(\i_im[1][16] ), .B(n7347), .X(n5027) );
  nand_x1_sg U12954 ( .A(\update_mask_0/reg_out[1][16] ), .B(n6454), .X(n5028)
         );
  nand_x1_sg U12955 ( .A(\i_im[1][15] ), .B(n7342), .X(n5025) );
  nand_x1_sg U12956 ( .A(\update_mask_0/reg_out[1][15] ), .B(n7026), .X(n5026)
         );
  nand_x1_sg U12957 ( .A(\i_im[1][14] ), .B(n6296), .X(n5023) );
  nand_x1_sg U12958 ( .A(\update_mask_0/reg_out[1][14] ), .B(n6355), .X(n5024)
         );
  nand_x1_sg U12959 ( .A(\i_im[1][5] ), .B(n6258), .X(n5005) );
  nand_x1_sg U12960 ( .A(\update_mask_0/reg_out[1][5] ), .B(n7035), .X(n5006)
         );
  nand_x1_sg U12961 ( .A(\i_im[1][4] ), .B(n7348), .X(n5003) );
  nand_x1_sg U12962 ( .A(\update_mask_0/reg_out[1][4] ), .B(n7027), .X(n5004)
         );
  nand_x1_sg U12963 ( .A(\i_im[1][3] ), .B(n7364), .X(n5001) );
  nand_x1_sg U12964 ( .A(\update_mask_0/reg_out[1][3] ), .B(n7044), .X(n5002)
         );
  nand_x1_sg U12965 ( .A(\i_im[1][2] ), .B(n6526), .X(n4999) );
  nand_x1_sg U12966 ( .A(\update_mask_0/reg_out[1][2] ), .B(n7021), .X(n5000)
         );
  nand_x1_sg U12967 ( .A(\i_im[1][1] ), .B(n7352), .X(n4997) );
  nand_x1_sg U12968 ( .A(\update_mask_0/reg_out[1][1] ), .B(n5995), .X(n4998)
         );
  nand_x1_sg U12969 ( .A(\i_im[1][0] ), .B(n6301), .X(n4995) );
  nand_x1_sg U12970 ( .A(\update_mask_0/reg_out[1][0] ), .B(n6267), .X(n4996)
         );
  nand_x1_sg U12971 ( .A(\i_im[0][19] ), .B(n7354), .X(n4993) );
  nand_x1_sg U12972 ( .A(\update_mask_0/reg_out[0][19] ), .B(n7027), .X(n4994)
         );
  nand_x1_sg U12973 ( .A(\i_im[0][18] ), .B(n6249), .X(n4991) );
  nand_x1_sg U12974 ( .A(\update_mask_0/reg_out[0][18] ), .B(n6360), .X(n4992)
         );
  nand_x1_sg U12975 ( .A(\i_im[0][17] ), .B(n6255), .X(n4989) );
  nand_x1_sg U12976 ( .A(\update_mask_0/reg_out[0][17] ), .B(n5988), .X(n4990)
         );
  nand_x1_sg U12977 ( .A(\i_im[0][16] ), .B(n6547), .X(n4987) );
  nand_x1_sg U12978 ( .A(\update_mask_0/reg_out[0][16] ), .B(n6447), .X(n4988)
         );
  nand_x1_sg U12979 ( .A(\i_im[0][15] ), .B(n6250), .X(n4985) );
  nand_x1_sg U12980 ( .A(\update_mask_0/reg_out[0][15] ), .B(n5994), .X(n4986)
         );
  nand_x1_sg U12981 ( .A(\i_im[0][14] ), .B(n6519), .X(n4983) );
  nand_x1_sg U12982 ( .A(\update_mask_0/reg_out[0][14] ), .B(n6456), .X(n4984)
         );
  nand_x1_sg U12983 ( .A(\i_im[0][13] ), .B(n6514), .X(n4981) );
  nand_x1_sg U12984 ( .A(\update_mask_0/reg_out[0][13] ), .B(n7327), .X(n4982)
         );
  nand_x1_sg U12985 ( .A(\i_im[0][12] ), .B(n7367), .X(n4979) );
  nand_x1_sg U12986 ( .A(\update_mask_0/reg_out[0][12] ), .B(n6450), .X(n4980)
         );
  nand_x1_sg U12987 ( .A(\i_im[0][11] ), .B(n7343), .X(n4977) );
  nand_x1_sg U12988 ( .A(\update_mask_0/reg_out[0][11] ), .B(n7038), .X(n4978)
         );
  nand_x1_sg U12989 ( .A(\i_im[0][10] ), .B(n7358), .X(n4975) );
  nand_x1_sg U12990 ( .A(\update_mask_0/reg_out[0][10] ), .B(n6287), .X(n4976)
         );
  nand_x1_sg U12991 ( .A(\i_im[0][9] ), .B(n6261), .X(n4973) );
  nand_x1_sg U12992 ( .A(\update_mask_0/reg_out[0][9] ), .B(n7028), .X(n4974)
         );
  nand_x1_sg U12993 ( .A(\i_im[0][8] ), .B(n6467), .X(n4971) );
  nand_x1_sg U12994 ( .A(\update_mask_0/reg_out[0][8] ), .B(n6450), .X(n4972)
         );
  nand_x1_sg U12995 ( .A(\i_im[0][7] ), .B(n7368), .X(n4969) );
  nand_x1_sg U12996 ( .A(\update_mask_0/reg_out[0][7] ), .B(n6268), .X(n4970)
         );
  nand_x1_sg U12997 ( .A(\i_im[0][6] ), .B(n6535), .X(n4967) );
  nand_x1_sg U12998 ( .A(\update_mask_0/reg_out[0][6] ), .B(n7023), .X(n4968)
         );
  nand_x1_sg U12999 ( .A(\i_im[0][5] ), .B(n6262), .X(n4965) );
  nand_x1_sg U13000 ( .A(\update_mask_0/reg_out[0][5] ), .B(n6355), .X(n4966)
         );
  nand_x1_sg U13001 ( .A(\i_im[0][4] ), .B(n6468), .X(n4963) );
  nand_x1_sg U13002 ( .A(\update_mask_0/reg_out[0][4] ), .B(n6359), .X(n4964)
         );
  nand_x1_sg U13003 ( .A(\i_im[0][3] ), .B(n6537), .X(n4961) );
  nand_x1_sg U13004 ( .A(\update_mask_0/reg_out[0][3] ), .B(n5994), .X(n4962)
         );
  nand_x1_sg U13005 ( .A(\i_im[0][2] ), .B(n6463), .X(n4959) );
  nand_x1_sg U13006 ( .A(\update_mask_0/reg_out[0][2] ), .B(n7040), .X(n4960)
         );
  nand_x1_sg U13007 ( .A(\i_im[0][1] ), .B(n6256), .X(n4957) );
  nand_x1_sg U13008 ( .A(\update_mask_0/reg_out[0][1] ), .B(n7043), .X(n4958)
         );
  nand_x1_sg U13009 ( .A(\i_im[0][0] ), .B(n6545), .X(n4955) );
  nand_x1_sg U13010 ( .A(\update_mask_0/reg_out[0][0] ), .B(n7334), .X(n4956)
         );
  nand_x1_sg U13011 ( .A(i_mask[31]), .B(n6526), .X(n4953) );
  nand_x1_sg U13012 ( .A(\update_mask_0/reg_i_mask[31] ), .B(n7025), .X(n4954)
         );
  nand_x1_sg U13013 ( .A(i_mask[30]), .B(n6261), .X(n4951) );
  nand_x1_sg U13014 ( .A(\update_mask_0/reg_i_mask[30] ), .B(n5996), .X(n4952)
         );
  nand_x1_sg U13015 ( .A(i_mask[29]), .B(n6546), .X(n4949) );
  nand_x1_sg U13016 ( .A(\update_mask_0/reg_i_mask[29] ), .B(n7033), .X(n4950)
         );
  nand_x1_sg U13017 ( .A(i_mask[28]), .B(n7348), .X(n4947) );
  nand_x1_sg U13018 ( .A(\update_mask_0/reg_i_mask[28] ), .B(n6287), .X(n4948)
         );
  nand_x1_sg U13019 ( .A(i_mask[27]), .B(n6537), .X(n4945) );
  nand_x1_sg U13020 ( .A(\update_mask_0/reg_i_mask[27] ), .B(n6359), .X(n4946)
         );
  nand_x1_sg U13021 ( .A(i_mask[26]), .B(n7366), .X(n4943) );
  nand_x1_sg U13022 ( .A(\update_mask_0/reg_i_mask[26] ), .B(n7039), .X(n4944)
         );
  nand_x1_sg U13023 ( .A(i_mask[25]), .B(n6087), .X(n4941) );
  nand_x1_sg U13024 ( .A(\update_mask_0/reg_i_mask[25] ), .B(n6357), .X(n4942)
         );
  nand_x1_sg U13025 ( .A(i_mask[24]), .B(n7363), .X(n4939) );
  nand_x1_sg U13026 ( .A(\update_mask_0/reg_i_mask[24] ), .B(n7041), .X(n4940)
         );
  nand_x1_sg U13027 ( .A(i_mask[23]), .B(n6534), .X(n4937) );
  nand_x1_sg U13028 ( .A(\update_mask_0/reg_i_mask[23] ), .B(n7330), .X(n4938)
         );
  nand_x1_sg U13029 ( .A(i_mask[22]), .B(n6296), .X(n4935) );
  nand_x1_sg U13030 ( .A(\update_mask_0/reg_i_mask[22] ), .B(n7051), .X(n4936)
         );
  nand_x1_sg U13031 ( .A(i_mask[20]), .B(n6297), .X(n4931) );
  nand_x1_sg U13032 ( .A(\update_mask_0/reg_i_mask[20] ), .B(n5987), .X(n4932)
         );
  nand_x1_sg U13033 ( .A(i_mask[19]), .B(n7347), .X(n4929) );
  nand_x1_sg U13034 ( .A(\update_mask_0/reg_i_mask[19] ), .B(n5987), .X(n4930)
         );
  nand_x1_sg U13035 ( .A(i_mask[18]), .B(n6294), .X(n4927) );
  nand_x1_sg U13036 ( .A(\update_mask_0/reg_i_mask[18] ), .B(n6277), .X(n4928)
         );
  nand_x1_sg U13037 ( .A(i_mask[17]), .B(n6295), .X(n4925) );
  nand_x1_sg U13038 ( .A(\update_mask_0/reg_i_mask[17] ), .B(n7049), .X(n4926)
         );
  nand_x1_sg U13039 ( .A(i_mask[16]), .B(n6087), .X(n4923) );
  nand_x1_sg U13040 ( .A(\update_mask_0/reg_i_mask[16] ), .B(n7036), .X(n4924)
         );
  nand_x1_sg U13041 ( .A(i_mask[15]), .B(n7351), .X(n4921) );
  nand_x1_sg U13042 ( .A(\update_mask_0/reg_i_mask[15] ), .B(n7325), .X(n4922)
         );
  nand_x1_sg U13043 ( .A(i_mask[14]), .B(n7353), .X(n4919) );
  nand_x1_sg U13044 ( .A(\update_mask_0/reg_i_mask[14] ), .B(n5989), .X(n4920)
         );
  nand_x1_sg U13045 ( .A(i_mask[13]), .B(n6087), .X(n4917) );
  nand_x1_sg U13046 ( .A(\update_mask_0/reg_i_mask[13] ), .B(n7023), .X(n4918)
         );
  nand_x1_sg U13047 ( .A(i_mask[12]), .B(n7353), .X(n4915) );
  nand_x1_sg U13048 ( .A(\update_mask_0/reg_i_mask[12] ), .B(n6145), .X(n4916)
         );
  nand_x1_sg U13049 ( .A(i_mask[11]), .B(n6529), .X(n4913) );
  nand_x1_sg U13050 ( .A(\update_mask_0/reg_i_mask[11] ), .B(n6153), .X(n4914)
         );
  nand_x1_sg U13051 ( .A(i_mask[10]), .B(n6092), .X(n4911) );
  nand_x1_sg U13052 ( .A(\update_mask_0/reg_i_mask[10] ), .B(n7040), .X(n4912)
         );
  nand_x1_sg U13053 ( .A(i_mask[9]), .B(n6250), .X(n4909) );
  nand_x1_sg U13054 ( .A(\update_mask_0/reg_i_mask[9] ), .B(n6286), .X(n4910)
         );
  nand_x1_sg U13055 ( .A(i_mask[8]), .B(n7349), .X(n4907) );
  nand_x1_sg U13056 ( .A(\update_mask_0/reg_i_mask[8] ), .B(n7033), .X(n4908)
         );
  nand_x1_sg U13057 ( .A(i_mask[7]), .B(n6088), .X(n4905) );
  nand_x1_sg U13058 ( .A(\update_mask_0/reg_i_mask[7] ), .B(n7025), .X(n4906)
         );
  nand_x1_sg U13059 ( .A(i_mask[5]), .B(n7364), .X(n4901) );
  nand_x1_sg U13060 ( .A(\update_mask_0/reg_i_mask[5] ), .B(n6453), .X(n4902)
         );
  nand_x1_sg U13061 ( .A(i_mask[4]), .B(n6517), .X(n4899) );
  nand_x1_sg U13062 ( .A(\update_mask_0/reg_i_mask[4] ), .B(n7031), .X(n4900)
         );
  nand_x1_sg U13063 ( .A(i_mask[3]), .B(n6547), .X(n4897) );
  nand_x1_sg U13064 ( .A(\update_mask_0/reg_i_mask[3] ), .B(n7330), .X(n4898)
         );
  nand_x1_sg U13065 ( .A(i_mask[2]), .B(n6524), .X(n4895) );
  nand_x1_sg U13066 ( .A(\update_mask_0/reg_i_mask[2] ), .B(n7025), .X(n4896)
         );
  nand_x1_sg U13067 ( .A(i_mask[1]), .B(n7362), .X(n4893) );
  nand_x1_sg U13068 ( .A(\update_mask_0/reg_i_mask[1] ), .B(n7326), .X(n4894)
         );
  nand_x1_sg U13069 ( .A(i_mask[0]), .B(n6257), .X(n4889) );
  nand_x1_sg U13070 ( .A(\update_mask_0/reg_i_mask[0] ), .B(n6281), .X(n4890)
         );
  nand_x1_sg U13071 ( .A(\i_im[11][9] ), .B(n7364), .X(n5413) );
  nand_x1_sg U13072 ( .A(\update_mask_0/reg_out[11][9] ), .B(n6148), .X(n5414)
         );
  nand_x1_sg U13073 ( .A(\i_im[11][8] ), .B(n7359), .X(n5411) );
  nand_x1_sg U13074 ( .A(\update_mask_0/reg_out[11][8] ), .B(n6149), .X(n5412)
         );
  nand_x1_sg U13075 ( .A(\i_im[11][7] ), .B(n6249), .X(n5409) );
  nand_x1_sg U13076 ( .A(\update_mask_0/reg_out[11][7] ), .B(n7024), .X(n5410)
         );
  nand_x1_sg U13077 ( .A(\i_im[11][6] ), .B(n7368), .X(n5407) );
  nand_x1_sg U13078 ( .A(\update_mask_0/reg_out[11][6] ), .B(n7026), .X(n5408)
         );
  nand_x1_sg U13079 ( .A(\i_im[11][5] ), .B(n6514), .X(n5405) );
  nand_x1_sg U13080 ( .A(\update_mask_0/reg_out[11][5] ), .B(n6356), .X(n5406)
         );
  nand_x1_sg U13081 ( .A(\i_im[11][4] ), .B(n6523), .X(n5403) );
  nand_x1_sg U13082 ( .A(\update_mask_0/reg_out[11][4] ), .B(n6456), .X(n5404)
         );
  nand_x1_sg U13083 ( .A(\i_im[11][3] ), .B(n6254), .X(n5401) );
  nand_x1_sg U13084 ( .A(\update_mask_0/reg_out[11][3] ), .B(n5993), .X(n5402)
         );
  nand_x1_sg U13085 ( .A(\i_im[11][2] ), .B(n6522), .X(n5399) );
  nand_x1_sg U13086 ( .A(\update_mask_0/reg_out[11][2] ), .B(n7334), .X(n5400)
         );
  nand_x1_sg U13087 ( .A(\i_im[6][11] ), .B(n6532), .X(n5217) );
  nand_x1_sg U13088 ( .A(\update_mask_0/reg_out[6][11] ), .B(n6276), .X(n5218)
         );
  nand_x1_sg U13089 ( .A(\i_im[6][10] ), .B(n7368), .X(n5215) );
  nand_x1_sg U13090 ( .A(\update_mask_0/reg_out[6][10] ), .B(n7045), .X(n5216)
         );
  nand_x1_sg U13091 ( .A(\i_im[6][9] ), .B(n6536), .X(n5213) );
  nand_x1_sg U13092 ( .A(\update_mask_0/reg_out[6][9] ), .B(n7044), .X(n5214)
         );
  nand_x1_sg U13093 ( .A(\i_im[6][8] ), .B(n7361), .X(n5211) );
  nand_x1_sg U13094 ( .A(\update_mask_0/reg_out[6][8] ), .B(n6282), .X(n5212)
         );
  nand_x1_sg U13095 ( .A(\i_im[6][7] ), .B(n6253), .X(n5209) );
  nand_x1_sg U13096 ( .A(\update_mask_0/reg_out[6][7] ), .B(n6291), .X(n5210)
         );
  nand_x1_sg U13097 ( .A(\i_im[6][6] ), .B(n7361), .X(n5207) );
  nand_x1_sg U13098 ( .A(\update_mask_0/reg_out[6][6] ), .B(n6454), .X(n5208)
         );
  nand_x1_sg U13099 ( .A(\i_im[6][5] ), .B(n7372), .X(n5205) );
  nand_x1_sg U13100 ( .A(\update_mask_0/reg_out[6][5] ), .B(n6291), .X(n5206)
         );
  nand_x1_sg U13101 ( .A(\i_im[6][4] ), .B(n6530), .X(n5203) );
  nand_x1_sg U13102 ( .A(\update_mask_0/reg_out[6][4] ), .B(n7039), .X(n5204)
         );
  nand_x1_sg U13103 ( .A(\i_im[1][13] ), .B(n6534), .X(n5021) );
  nand_x1_sg U13104 ( .A(\update_mask_0/reg_out[1][13] ), .B(n7331), .X(n5022)
         );
  nand_x1_sg U13105 ( .A(\i_im[1][12] ), .B(n6531), .X(n5019) );
  nand_x1_sg U13106 ( .A(\update_mask_0/reg_out[1][12] ), .B(n6449), .X(n5020)
         );
  nand_x1_sg U13107 ( .A(\i_im[1][11] ), .B(n6526), .X(n5017) );
  nand_x1_sg U13108 ( .A(\update_mask_0/reg_out[1][11] ), .B(n6271), .X(n5018)
         );
  nand_x1_sg U13109 ( .A(\i_im[1][10] ), .B(n6525), .X(n5015) );
  nand_x1_sg U13110 ( .A(\update_mask_0/reg_out[1][10] ), .B(n6143), .X(n5016)
         );
  nand_x1_sg U13111 ( .A(\i_im[1][9] ), .B(n6262), .X(n5013) );
  nand_x1_sg U13112 ( .A(\update_mask_0/reg_out[1][9] ), .B(n5992), .X(n5014)
         );
  nand_x1_sg U13113 ( .A(\i_im[1][8] ), .B(n6090), .X(n5011) );
  nand_x1_sg U13114 ( .A(\update_mask_0/reg_out[1][8] ), .B(n6267), .X(n5012)
         );
  nand_x1_sg U13115 ( .A(\i_im[1][7] ), .B(n7346), .X(n5009) );
  nand_x1_sg U13116 ( .A(\update_mask_0/reg_out[1][7] ), .B(n7327), .X(n5010)
         );
  nand_x1_sg U13117 ( .A(\i_im[1][6] ), .B(n6525), .X(n5007) );
  nand_x1_sg U13118 ( .A(\update_mask_0/reg_out[1][6] ), .B(n5990), .X(n5008)
         );
  nand_x1_sg U13119 ( .A(n4126), .B(n6312), .X(n3783) );
  nor_x1_sg U13120 ( .A(n6333), .B(n7404), .X(n4126) );
  nor_x1_sg U13121 ( .A(n5921), .B(\output_state[0] ), .X(n4863) );
  nor_x1_sg U13122 ( .A(n4834), .B(n4835), .X(n4832) );
  nand_x1_sg U13123 ( .A(n7132), .B(n5897), .X(n4833) );
  nor_x1_sg U13124 ( .A(\update_output_0/pre_o_im[13][19] ), .B(n6915), .X(
        n4835) );
  nor_x1_sg U13125 ( .A(n4760), .B(n4761), .X(n4758) );
  nand_x1_sg U13126 ( .A(n7134), .B(n5717), .X(n4759) );
  nor_x1_sg U13127 ( .A(\update_output_0/pre_o_im[13][17] ), .B(n6917), .X(
        n4761) );
  nor_x1_sg U13128 ( .A(n4688), .B(n4689), .X(n4686) );
  nand_x1_sg U13129 ( .A(n7135), .B(n5908), .X(n4687) );
  nor_x1_sg U13130 ( .A(\update_output_0/pre_o_im[13][15] ), .B(n6920), .X(
        n4689) );
  nor_x1_sg U13131 ( .A(n4616), .B(n4617), .X(n4614) );
  nand_x1_sg U13132 ( .A(n7130), .B(n5866), .X(n4615) );
  nor_x1_sg U13133 ( .A(\update_output_0/pre_o_im[13][13] ), .B(n6920), .X(
        n4617) );
  nor_x1_sg U13134 ( .A(n4544), .B(n4545), .X(n4542) );
  nand_x1_sg U13135 ( .A(n7141), .B(n5729), .X(n4543) );
  nor_x1_sg U13136 ( .A(\update_output_0/pre_o_im[13][11] ), .B(n6915), .X(
        n4545) );
  nor_x1_sg U13137 ( .A(n4472), .B(n4473), .X(n4470) );
  nand_x1_sg U13138 ( .A(n7136), .B(n5906), .X(n4471) );
  nor_x1_sg U13139 ( .A(\update_output_0/pre_o_im[13][9] ), .B(n6914), .X(
        n4473) );
  nor_x1_sg U13140 ( .A(n4256), .B(n4257), .X(n4254) );
  nand_x1_sg U13141 ( .A(n7134), .B(n5861), .X(n4255) );
  nor_x1_sg U13142 ( .A(\update_output_0/pre_o_im[13][3] ), .B(n6919), .X(
        n4257) );
  nor_x1_sg U13143 ( .A(n4184), .B(n4185), .X(n4182) );
  nand_x1_sg U13144 ( .A(n7129), .B(n5836), .X(n4183) );
  nor_x1_sg U13145 ( .A(\update_output_0/pre_o_im[13][1] ), .B(n6919), .X(
        n4185) );
  nor_x1_sg U13146 ( .A(n4796), .B(n4797), .X(n4794) );
  nand_x1_sg U13147 ( .A(n7134), .B(n5863), .X(n4795) );
  nor_x1_sg U13148 ( .A(\update_output_0/pre_o_im[13][18] ), .B(n6917), .X(
        n4797) );
  nor_x1_sg U13149 ( .A(n4724), .B(n4725), .X(n4722) );
  nand_x1_sg U13150 ( .A(n7137), .B(n5894), .X(n4723) );
  nor_x1_sg U13151 ( .A(\update_output_0/pre_o_im[13][16] ), .B(n6918), .X(
        n4725) );
  nor_x1_sg U13152 ( .A(n4652), .B(n4653), .X(n4650) );
  nand_x1_sg U13153 ( .A(n7130), .B(n5723), .X(n4651) );
  nor_x1_sg U13154 ( .A(\update_output_0/pre_o_im[13][14] ), .B(n6914), .X(
        n4653) );
  nor_x1_sg U13155 ( .A(n4580), .B(n4581), .X(n4578) );
  nand_x1_sg U13156 ( .A(n7141), .B(n5907), .X(n4579) );
  nor_x1_sg U13157 ( .A(\update_output_0/pre_o_im[13][12] ), .B(n6919), .X(
        n4581) );
  nor_x1_sg U13158 ( .A(n4508), .B(n4509), .X(n4506) );
  nand_x1_sg U13159 ( .A(n7142), .B(n5843), .X(n4507) );
  nor_x1_sg U13160 ( .A(\update_output_0/pre_o_im[13][10] ), .B(n6915), .X(
        n4509) );
  nor_x1_sg U13161 ( .A(n4436), .B(n4437), .X(n4434) );
  nand_x1_sg U13162 ( .A(n7131), .B(n5733), .X(n4435) );
  nor_x1_sg U13163 ( .A(\update_output_0/pre_o_im[13][8] ), .B(n6914), .X(
        n4437) );
  nor_x1_sg U13164 ( .A(n4220), .B(n4221), .X(n4218) );
  nand_x1_sg U13165 ( .A(n7135), .B(n5741), .X(n4219) );
  nor_x1_sg U13166 ( .A(\update_output_0/pre_o_im[13][2] ), .B(n6917), .X(
        n4221) );
  nor_x1_sg U13167 ( .A(n4144), .B(n4145), .X(n4141) );
  nand_x1_sg U13168 ( .A(n7129), .B(n5711), .X(n4142) );
  nor_x1_sg U13169 ( .A(\update_output_0/pre_o_im[13][0] ), .B(n6920), .X(
        n4145) );
  nand_x1_sg U13170 ( .A(n4849), .B(n6333), .X(n4146) );
  nand_x4_sg U13171 ( .A(n4847), .B(n4848), .X(n4843) );
  nand_x1_sg U13172 ( .A(n6237), .B(n5849), .X(n4845) );
  nand_x4_sg U13173 ( .A(n4809), .B(n4810), .X(n4805) );
  nand_x1_sg U13174 ( .A(n6236), .B(n5745), .X(n4807) );
  nand_x4_sg U13175 ( .A(n4269), .B(n4270), .X(n4265) );
  nand_x1_sg U13176 ( .A(n6236), .B(n5761), .X(n4267) );
  nand_x4_sg U13177 ( .A(n4233), .B(n4234), .X(n4229) );
  nand_x1_sg U13178 ( .A(n7258), .B(n5762), .X(n4231) );
  nand_x4_sg U13179 ( .A(n4773), .B(n4774), .X(n4769) );
  nand_x1_sg U13180 ( .A(n7255), .B(n5718), .X(n4771) );
  nand_x4_sg U13181 ( .A(n4737), .B(n4738), .X(n4733) );
  nand_x1_sg U13182 ( .A(n6393), .B(n5878), .X(n4735) );
  nand_x4_sg U13183 ( .A(n4701), .B(n4702), .X(n4697) );
  nand_x1_sg U13184 ( .A(n6077), .B(n5747), .X(n4699) );
  nand_x4_sg U13185 ( .A(n4665), .B(n4666), .X(n4661) );
  nand_x1_sg U13186 ( .A(n7256), .B(n5724), .X(n4663) );
  nand_x4_sg U13187 ( .A(n4629), .B(n4630), .X(n4625) );
  nand_x1_sg U13188 ( .A(n6236), .B(n5837), .X(n4627) );
  nand_x4_sg U13189 ( .A(n4593), .B(n4594), .X(n4589) );
  nand_x1_sg U13190 ( .A(n7255), .B(n5749), .X(n4591) );
  nand_x4_sg U13191 ( .A(n4557), .B(n4558), .X(n4553) );
  nand_x1_sg U13192 ( .A(n6237), .B(n5750), .X(n4555) );
  nand_x4_sg U13193 ( .A(n4521), .B(n4522), .X(n4517) );
  nand_x1_sg U13194 ( .A(n7256), .B(n5891), .X(n4519) );
  nand_x4_sg U13195 ( .A(n4485), .B(n4486), .X(n4481) );
  nand_x1_sg U13196 ( .A(n7257), .B(n5753), .X(n4483) );
  nand_x4_sg U13197 ( .A(n4449), .B(n4450), .X(n4445) );
  nand_x1_sg U13198 ( .A(n7257), .B(n5754), .X(n4447) );
  nand_x4_sg U13199 ( .A(n4197), .B(n4198), .X(n4193) );
  nand_x1_sg U13200 ( .A(n7255), .B(n5880), .X(n4195) );
  nand_x4_sg U13201 ( .A(n4161), .B(n4162), .X(n4157) );
  nand_x1_sg U13202 ( .A(n6394), .B(n5713), .X(n4159) );
  nor_x1_sg U13203 ( .A(n6473), .B(n4307), .X(n4305) );
  nand_x1_sg U13204 ( .A(n6893), .B(n5782), .X(n4306) );
  nor_x1_sg U13205 ( .A(\update_output_0/pre_o_im[4][4] ), .B(n7242), .X(n4307) );
  nor_x1_sg U13206 ( .A(n6469), .B(n4415), .X(n4413) );
  nand_x1_sg U13207 ( .A(n6894), .B(n5787), .X(n4414) );
  nor_x1_sg U13208 ( .A(\update_output_0/pre_o_im[4][7] ), .B(n7247), .X(n4415) );
  nor_x1_sg U13209 ( .A(n7315), .B(n4379), .X(n4377) );
  nand_x1_sg U13210 ( .A(n6895), .B(n5676), .X(n4378) );
  nor_x1_sg U13211 ( .A(\update_output_0/pre_o_im[4][6] ), .B(n7251), .X(n4379) );
  nor_x1_sg U13212 ( .A(n7316), .B(n4343), .X(n4341) );
  nand_x1_sg U13213 ( .A(n6896), .B(n5790), .X(n4342) );
  nor_x1_sg U13214 ( .A(\update_output_0/pre_o_im[4][5] ), .B(n7249), .X(n4343) );
  nor_x1_sg U13215 ( .A(n6474), .B(n4811), .X(n4809) );
  nor_x1_sg U13216 ( .A(\update_output_0/pre_o_im[4][18] ), .B(n7249), .X(
        n4811) );
  nor_x1_sg U13217 ( .A(n7313), .B(n4775), .X(n4773) );
  nor_x1_sg U13218 ( .A(\update_output_0/pre_o_im[4][17] ), .B(n7247), .X(
        n4775) );
  nor_x1_sg U13219 ( .A(n6140), .B(n4739), .X(n4737) );
  nor_x1_sg U13220 ( .A(\update_output_0/pre_o_im[4][16] ), .B(n7245), .X(
        n4739) );
  nor_x1_sg U13221 ( .A(n7315), .B(n4703), .X(n4701) );
  nor_x1_sg U13222 ( .A(\update_output_0/pre_o_im[4][15] ), .B(n7251), .X(
        n4703) );
  nor_x1_sg U13223 ( .A(n7314), .B(n4667), .X(n4665) );
  nor_x1_sg U13224 ( .A(\update_output_0/pre_o_im[4][14] ), .B(n7244), .X(
        n4667) );
  nor_x1_sg U13225 ( .A(n7315), .B(n4631), .X(n4629) );
  nor_x1_sg U13226 ( .A(\update_output_0/pre_o_im[4][13] ), .B(n7245), .X(
        n4631) );
  nor_x1_sg U13227 ( .A(n7313), .B(n4595), .X(n4593) );
  nor_x1_sg U13228 ( .A(\update_output_0/pre_o_im[4][12] ), .B(n7252), .X(
        n4595) );
  nor_x1_sg U13229 ( .A(n6469), .B(n4559), .X(n4557) );
  nor_x1_sg U13230 ( .A(\update_output_0/pre_o_im[4][11] ), .B(n7250), .X(
        n4559) );
  nor_x1_sg U13231 ( .A(n6472), .B(n4523), .X(n4521) );
  nor_x1_sg U13232 ( .A(\update_output_0/pre_o_im[4][10] ), .B(n7242), .X(
        n4523) );
  nor_x1_sg U13233 ( .A(n6141), .B(n4487), .X(n4485) );
  nor_x1_sg U13234 ( .A(\update_output_0/pre_o_im[4][9] ), .B(n7244), .X(n4487) );
  nor_x1_sg U13235 ( .A(n6470), .B(n4451), .X(n4449) );
  nor_x1_sg U13236 ( .A(\update_output_0/pre_o_im[4][8] ), .B(n7250), .X(n4451) );
  nor_x1_sg U13237 ( .A(n6140), .B(n4271), .X(n4269) );
  nor_x1_sg U13238 ( .A(\update_output_0/pre_o_im[4][3] ), .B(n7253), .X(n4271) );
  nor_x1_sg U13239 ( .A(n6470), .B(n4235), .X(n4233) );
  nor_x1_sg U13240 ( .A(\update_output_0/pre_o_im[4][2] ), .B(n7246), .X(n4235) );
  nor_x1_sg U13241 ( .A(n7316), .B(n4199), .X(n4197) );
  nor_x1_sg U13242 ( .A(\update_output_0/pre_o_im[4][1] ), .B(n7253), .X(n4199) );
  nor_x1_sg U13243 ( .A(n6472), .B(n4163), .X(n4161) );
  nor_x1_sg U13244 ( .A(\update_output_0/pre_o_im[4][0] ), .B(n7247), .X(n4163) );
  nor_x1_sg U13245 ( .A(n6473), .B(n4850), .X(n4847) );
  nor_x1_sg U13246 ( .A(\update_output_0/pre_o_im[4][19] ), .B(n7253), .X(
        n4850) );
  nand_x1_sg U13247 ( .A(n7132), .B(n5744), .X(n4846) );
  nand_x1_sg U13248 ( .A(n7135), .B(n5819), .X(n4808) );
  nand_x1_sg U13249 ( .A(n7142), .B(n5900), .X(n4772) );
  nand_x1_sg U13250 ( .A(n7140), .B(n5746), .X(n4736) );
  nand_x1_sg U13251 ( .A(n7134), .B(n5893), .X(n4700) );
  nand_x1_sg U13252 ( .A(n7140), .B(n5850), .X(n4664) );
  nand_x1_sg U13253 ( .A(n7131), .B(n5748), .X(n4628) );
  nand_x1_sg U13254 ( .A(n7142), .B(n5848), .X(n4592) );
  nand_x1_sg U13255 ( .A(n7140), .B(n5855), .X(n4556) );
  nand_x1_sg U13256 ( .A(n7139), .B(n5752), .X(n4520) );
  nand_x1_sg U13257 ( .A(n7137), .B(n5856), .X(n4484) );
  nand_x1_sg U13258 ( .A(n7130), .B(n5838), .X(n4448) );
  nand_x1_sg U13259 ( .A(n7141), .B(n5874), .X(n4268) );
  nand_x1_sg U13260 ( .A(n7136), .B(n5853), .X(n4232) );
  nand_x1_sg U13261 ( .A(n7132), .B(n5764), .X(n4196) );
  nand_x1_sg U13262 ( .A(n7139), .B(n5822), .X(n4160) );
  nor_x1_sg U13263 ( .A(\update_output_0/pre_o_im[12][19] ), .B(n7245), .X(
        n4834) );
  nor_x1_sg U13264 ( .A(\update_output_0/pre_o_im[12][18] ), .B(n7242), .X(
        n4796) );
  nor_x1_sg U13265 ( .A(\update_output_0/pre_o_im[12][17] ), .B(n7251), .X(
        n4760) );
  nor_x1_sg U13266 ( .A(\update_output_0/pre_o_im[12][16] ), .B(n7242), .X(
        n4724) );
  nor_x1_sg U13267 ( .A(\update_output_0/pre_o_im[12][15] ), .B(n7249), .X(
        n4688) );
  nor_x1_sg U13268 ( .A(\update_output_0/pre_o_im[12][14] ), .B(n7246), .X(
        n4652) );
  nor_x1_sg U13269 ( .A(\update_output_0/pre_o_im[12][13] ), .B(n7246), .X(
        n4616) );
  nor_x1_sg U13270 ( .A(\update_output_0/pre_o_im[12][12] ), .B(n7244), .X(
        n4580) );
  nor_x1_sg U13271 ( .A(\update_output_0/pre_o_im[12][11] ), .B(n7246), .X(
        n4544) );
  nor_x1_sg U13272 ( .A(\update_output_0/pre_o_im[12][10] ), .B(n7247), .X(
        n4508) );
  nor_x1_sg U13273 ( .A(\update_output_0/pre_o_im[12][9] ), .B(n7244), .X(
        n4472) );
  nor_x1_sg U13274 ( .A(\update_output_0/pre_o_im[12][8] ), .B(n7252), .X(
        n4436) );
  nor_x1_sg U13275 ( .A(\update_output_0/pre_o_im[12][3] ), .B(n7250), .X(
        n4256) );
  nor_x1_sg U13276 ( .A(\update_output_0/pre_o_im[12][2] ), .B(n7249), .X(
        n4220) );
  nor_x1_sg U13277 ( .A(\update_output_0/pre_o_im[12][1] ), .B(n7245), .X(
        n4184) );
  nor_x1_sg U13278 ( .A(\update_output_0/pre_o_im[12][0] ), .B(n7252), .X(
        n4144) );
  nor_x1_sg U13279 ( .A(n4400), .B(n4401), .X(n4398) );
  nor_x1_sg U13280 ( .A(\update_output_0/pre_o_im[13][7] ), .B(n6919), .X(
        n4401) );
  nor_x1_sg U13281 ( .A(\update_output_0/pre_o_im[12][7] ), .B(n7250), .X(
        n4400) );
  nor_x1_sg U13282 ( .A(n4364), .B(n4365), .X(n4362) );
  nor_x1_sg U13283 ( .A(\update_output_0/pre_o_im[13][6] ), .B(n6915), .X(
        n4365) );
  nor_x1_sg U13284 ( .A(\update_output_0/pre_o_im[12][6] ), .B(n7251), .X(
        n4364) );
  nor_x1_sg U13285 ( .A(n4328), .B(n4329), .X(n4326) );
  nor_x1_sg U13286 ( .A(\update_output_0/pre_o_im[13][5] ), .B(n6918), .X(
        n4329) );
  nor_x1_sg U13287 ( .A(\update_output_0/pre_o_im[12][5] ), .B(n7253), .X(
        n4328) );
  nor_x1_sg U13288 ( .A(n4292), .B(n4293), .X(n4290) );
  nor_x1_sg U13289 ( .A(\update_output_0/pre_o_im[13][4] ), .B(n6917), .X(
        n4293) );
  nor_x1_sg U13290 ( .A(\update_output_0/pre_o_im[12][4] ), .B(n7252), .X(
        n4292) );
  nand_x1_sg U13291 ( .A(n7283), .B(n5694), .X(n4396) );
  nand_x1_sg U13292 ( .A(n6387), .B(n5903), .X(n4360) );
  nand_x1_sg U13293 ( .A(n6388), .B(n5777), .X(n4324) );
  nand_x1_sg U13294 ( .A(n6486), .B(n5696), .X(n4288) );
  nand_x1_sg U13295 ( .A(n6131), .B(n5686), .X(n4830) );
  nand_x1_sg U13296 ( .A(n6076), .B(n5714), .X(n4831) );
  nand_x1_sg U13297 ( .A(n6488), .B(n5794), .X(n4792) );
  nand_x1_sg U13298 ( .A(n6394), .B(n5905), .X(n4793) );
  nand_x1_sg U13299 ( .A(n7283), .B(n5769), .X(n4756) );
  nand_x1_sg U13300 ( .A(n7256), .B(n5821), .X(n4757) );
  nand_x1_sg U13301 ( .A(n7284), .B(n5688), .X(n4720) );
  nand_x1_sg U13302 ( .A(n6393), .B(n5720), .X(n4721) );
  nand_x1_sg U13303 ( .A(n6132), .B(n5786), .X(n4684) );
  nand_x1_sg U13304 ( .A(n7258), .B(n5875), .X(n4685) );
  nand_x1_sg U13305 ( .A(n6388), .B(n5808), .X(n4648) );
  nand_x1_sg U13306 ( .A(n6077), .B(n5859), .X(n4649) );
  nand_x1_sg U13307 ( .A(n7286), .B(n5690), .X(n4612) );
  nand_x1_sg U13308 ( .A(n7257), .B(n5726), .X(n4613) );
  nand_x1_sg U13309 ( .A(n7284), .B(n5795), .X(n4576) );
  nand_x1_sg U13310 ( .A(n6237), .B(n5869), .X(n4577) );
  nand_x1_sg U13311 ( .A(n6487), .B(n5812), .X(n4540) );
  nand_x1_sg U13312 ( .A(n6077), .B(n5867), .X(n4541) );
  nand_x1_sg U13313 ( .A(n7286), .B(n5692), .X(n4504) );
  nand_x1_sg U13314 ( .A(n7257), .B(n5730), .X(n4505) );
  nand_x1_sg U13315 ( .A(n6486), .B(n5876), .X(n4468) );
  nand_x1_sg U13316 ( .A(n7258), .B(n5857), .X(n4469) );
  nand_x1_sg U13317 ( .A(n7285), .B(n5771), .X(n4432) );
  nand_x1_sg U13318 ( .A(n6236), .B(n5890), .X(n4433) );
  nand_x1_sg U13319 ( .A(n6131), .B(n5873), .X(n4252) );
  nand_x1_sg U13320 ( .A(n6077), .B(n5901), .X(n4253) );
  nand_x1_sg U13321 ( .A(n6131), .B(n5815), .X(n4216) );
  nand_x1_sg U13322 ( .A(n6076), .B(n5881), .X(n4217) );
  nand_x1_sg U13323 ( .A(n6488), .B(n5698), .X(n4180) );
  nand_x1_sg U13324 ( .A(n6076), .B(n5742), .X(n4181) );
  nand_x1_sg U13325 ( .A(n6132), .B(n5766), .X(n4138) );
  nand_x1_sg U13326 ( .A(n6237), .B(n5851), .X(n4139) );
  nand_x1_sg U13327 ( .A(\update_mask_0/N26 ), .B(\update_mask_0/N27 ), .X(
        n4886) );
  nand_x1_sg U13328 ( .A(n6539), .B(n4888), .X(n4887) );
  nor_x1_sg U13329 ( .A(n7402), .B(n6329), .X(n4888) );
  nand_x1_sg U13330 ( .A(n4878), .B(n6310), .X(n4880) );
  nand_x1_sg U13331 ( .A(n4882), .B(n7016), .X(n4881) );
  nor_x1_sg U13332 ( .A(n4878), .B(n4879), .X(n4882) );
  nor_x1_sg U13333 ( .A(n6312), .B(n3471), .X(n3567) );
  nand_x1_sg U13334 ( .A(n6829), .B(n3480), .X(n3464) );
  nand_x1_sg U13335 ( .A(\update_output_0/n2821 ), .B(n6999), .X(n3480) );
  nand_x1_sg U13336 ( .A(\update_output_0/N33 ), .B(n7397), .X(n3466) );
  nand_x1_sg U13337 ( .A(n6509), .B(n6332), .X(n3479) );
  nand_x1_sg U13338 ( .A(n4856), .B(n4857), .X(n4851) );
  nand_x1_sg U13339 ( .A(n6194), .B(n5715), .X(n4853) );
  nand_x1_sg U13340 ( .A(n4816), .B(n4817), .X(n4812) );
  nand_x1_sg U13341 ( .A(n6423), .B(n5896), .X(n4814) );
  nand_x1_sg U13342 ( .A(n4780), .B(n4781), .X(n4776) );
  nand_x1_sg U13343 ( .A(n7124), .B(n5719), .X(n4778) );
  nand_x1_sg U13344 ( .A(n4744), .B(n4745), .X(n4740) );
  nand_x1_sg U13345 ( .A(n7123), .B(n5721), .X(n4742) );
  nand_x1_sg U13346 ( .A(n4708), .B(n4709), .X(n4704) );
  nand_x1_sg U13347 ( .A(n7125), .B(n5860), .X(n4706) );
  nand_x1_sg U13348 ( .A(n4672), .B(n4673), .X(n4668) );
  nand_x1_sg U13349 ( .A(n7126), .B(n5725), .X(n4670) );
  nand_x1_sg U13350 ( .A(n4636), .B(n4637), .X(n4632) );
  nand_x1_sg U13351 ( .A(n6195), .B(n5727), .X(n4634) );
  nand_x1_sg U13352 ( .A(n4600), .B(n4601), .X(n4596) );
  nand_x1_sg U13353 ( .A(n7124), .B(n5839), .X(n4598) );
  nand_x1_sg U13354 ( .A(n4564), .B(n4565), .X(n4560) );
  nand_x1_sg U13355 ( .A(n6032), .B(n5751), .X(n4562) );
  nand_x1_sg U13356 ( .A(n4528), .B(n4529), .X(n4524) );
  nand_x1_sg U13357 ( .A(n6502), .B(n5670), .X(n4527) );
  nand_x1_sg U13358 ( .A(n4492), .B(n4493), .X(n4488) );
  nand_x1_sg U13359 ( .A(n7065), .B(n5807), .X(n4491) );
  nand_x1_sg U13360 ( .A(n4456), .B(n4457), .X(n4452) );
  nand_x1_sg U13361 ( .A(n4276), .B(n4277), .X(n4272) );
  nand_x1_sg U13362 ( .A(n6194), .B(n5887), .X(n4274) );
  nand_x1_sg U13363 ( .A(n4240), .B(n4241), .X(n4236) );
  nand_x1_sg U13364 ( .A(n7125), .B(n5763), .X(n4238) );
  nand_x1_sg U13365 ( .A(n4204), .B(n4205), .X(n4200) );
  nand_x1_sg U13366 ( .A(n7123), .B(n5743), .X(n4202) );
  nand_x1_sg U13367 ( .A(n4168), .B(n4169), .X(n4164) );
  nand_x1_sg U13368 ( .A(n6424), .B(n5909), .X(n4166) );
  nand_x1_sg U13369 ( .A(n7275), .B(n5654), .X(n4856) );
  nand_x1_sg U13370 ( .A(n6391), .B(n5774), .X(n4816) );
  nand_x1_sg U13371 ( .A(n7276), .B(n5700), .X(n4780) );
  nand_x1_sg U13372 ( .A(n7275), .B(n5659), .X(n4744) );
  nand_x1_sg U13373 ( .A(n6494), .B(n5829), .X(n4708) );
  nand_x1_sg U13374 ( .A(n6494), .B(n5702), .X(n4672) );
  nand_x1_sg U13375 ( .A(n6391), .B(n5664), .X(n4636) );
  nand_x1_sg U13376 ( .A(n6392), .B(n5767), .X(n4600) );
  nand_x1_sg U13377 ( .A(n6495), .B(n5704), .X(n4564) );
  nand_x1_sg U13378 ( .A(n7276), .B(n5669), .X(n4528) );
  nand_x1_sg U13379 ( .A(n6392), .B(n5788), .X(n4492) );
  nand_x1_sg U13380 ( .A(n7276), .B(n5706), .X(n4456) );
  nand_x1_sg U13381 ( .A(n7275), .B(n5801), .X(n4276) );
  nand_x1_sg U13382 ( .A(n7274), .B(n5710), .X(n4240) );
  nand_x1_sg U13383 ( .A(n6125), .B(n5684), .X(n4204) );
  nand_x1_sg U13384 ( .A(n6495), .B(n5772), .X(n4168) );
  nand_x1_sg U13385 ( .A(n7285), .B(n5773), .X(n4857) );
  nand_x1_sg U13386 ( .A(n7286), .B(n5699), .X(n4817) );
  nand_x1_sg U13387 ( .A(n6487), .B(n5658), .X(n4781) );
  nand_x1_sg U13388 ( .A(n7285), .B(n5870), .X(n4745) );
  nand_x1_sg U13389 ( .A(n6387), .B(n5701), .X(n4709) );
  nand_x1_sg U13390 ( .A(n6388), .B(n5663), .X(n4673) );
  nand_x1_sg U13391 ( .A(n6487), .B(n5784), .X(n4637) );
  nand_x1_sg U13392 ( .A(n6486), .B(n5703), .X(n4601) );
  nand_x1_sg U13393 ( .A(n6131), .B(n5668), .X(n4565) );
  nand_x1_sg U13394 ( .A(n6388), .B(n5775), .X(n4529) );
  nand_x1_sg U13395 ( .A(n6387), .B(n5705), .X(n4493) );
  nand_x1_sg U13396 ( .A(n6488), .B(n5673), .X(n4457) );
  nand_x1_sg U13397 ( .A(n6387), .B(n5709), .X(n4277) );
  nand_x1_sg U13398 ( .A(n7284), .B(n5683), .X(n4241) );
  nand_x1_sg U13399 ( .A(n7286), .B(n5823), .X(n4205) );
  nand_x1_sg U13400 ( .A(n6486), .B(n5653), .X(n4169) );
  nand_x1_sg U13401 ( .A(n6132), .B(n5810), .X(n4421) );
  nand_x1_sg U13402 ( .A(n7274), .B(n5674), .X(n4420) );
  nand_x1_sg U13403 ( .A(n7285), .B(n5707), .X(n4385) );
  nand_x1_sg U13404 ( .A(n6496), .B(n5828), .X(n4384) );
  nand_x1_sg U13405 ( .A(n7283), .B(n5678), .X(n4349) );
  nand_x1_sg U13406 ( .A(n7273), .B(n5708), .X(n4348) );
  nand_x1_sg U13407 ( .A(n7284), .B(n5888), .X(n4313) );
  nand_x1_sg U13408 ( .A(n6126), .B(n5679), .X(n4312) );
  nor_x1_sg U13409 ( .A(n4855), .B(\update_output_0/N33 ), .X(n4154) );
  nand_x1_sg U13410 ( .A(n6332), .B(n7414), .X(n4855) );
  nand_x1_sg U13411 ( .A(n6500), .B(n5779), .X(n4405) );
  nand_x1_sg U13412 ( .A(n6498), .B(n5792), .X(n4369) );
  nand_x1_sg U13413 ( .A(n7065), .B(n5677), .X(n4333) );
  nand_x1_sg U13414 ( .A(n7067), .B(n5835), .X(n4297) );
  nand_x1_sg U13415 ( .A(n6494), .B(n5884), .X(n4406) );
  nand_x1_sg U13416 ( .A(n6391), .B(n5695), .X(n4370) );
  nand_x1_sg U13417 ( .A(n7275), .B(n5827), .X(n4334) );
  nand_x1_sg U13418 ( .A(n6392), .B(n5785), .X(n4298) );
  nand_x1_sg U13419 ( .A(n6392), .B(n5693), .X(n4478) );
  nand_x1_sg U13420 ( .A(n6125), .B(n5816), .X(n4840) );
  nand_x1_sg U13421 ( .A(n6501), .B(n5791), .X(n4839) );
  nand_x1_sg U13422 ( .A(n7274), .B(n5687), .X(n4802) );
  nand_x1_sg U13423 ( .A(n6004), .B(n5781), .X(n4801) );
  nand_x1_sg U13424 ( .A(n6494), .B(n5783), .X(n4766) );
  nand_x1_sg U13425 ( .A(n6497), .B(n5657), .X(n4765) );
  nand_x1_sg U13426 ( .A(n6496), .B(n5826), .X(n4730) );
  nand_x1_sg U13427 ( .A(n6498), .B(n5802), .X(n4729) );
  nand_x1_sg U13428 ( .A(n7276), .B(n5689), .X(n4694) );
  nand_x1_sg U13429 ( .A(n6497), .B(n5871), .X(n4693) );
  nand_x1_sg U13430 ( .A(n6126), .B(n5798), .X(n4658) );
  nand_x1_sg U13431 ( .A(n7064), .B(n5662), .X(n4657) );
  nand_x1_sg U13432 ( .A(n6126), .B(n5832), .X(n4622) );
  nand_x1_sg U13433 ( .A(n6498), .B(n5824), .X(n4621) );
  nand_x1_sg U13434 ( .A(n6496), .B(n5691), .X(n4586) );
  nand_x1_sg U13435 ( .A(n7064), .B(n5776), .X(n4585) );
  nand_x1_sg U13436 ( .A(n7273), .B(n5803), .X(n4550) );
  nand_x1_sg U13437 ( .A(n7066), .B(n5667), .X(n4549) );
  nand_x1_sg U13438 ( .A(n6125), .B(n5804), .X(n4514) );
  nand_x1_sg U13439 ( .A(n6500), .B(n5834), .X(n4513) );
  nand_x1_sg U13440 ( .A(n7274), .B(n5833), .X(n4442) );
  nand_x1_sg U13441 ( .A(n6004), .B(n5672), .X(n4441) );
  nand_x1_sg U13442 ( .A(n6391), .B(n5697), .X(n4262) );
  nand_x1_sg U13443 ( .A(n6005), .B(n5817), .X(n4261) );
  nand_x1_sg U13444 ( .A(n6125), .B(n5799), .X(n4226) );
  nand_x1_sg U13445 ( .A(n7067), .B(n5682), .X(n4225) );
  nand_x1_sg U13446 ( .A(n6495), .B(n5797), .X(n4190) );
  nand_x1_sg U13447 ( .A(n6502), .B(n5811), .X(n4189) );
  nand_x1_sg U13448 ( .A(n7273), .B(n5652), .X(n4153) );
  nand_x1_sg U13449 ( .A(n7065), .B(n5910), .X(n4152) );
  nand_x1_sg U13450 ( .A(n6473), .B(n4404), .X(n4403) );
  nand_x1_sg U13451 ( .A(n6194), .B(n5847), .X(n4404) );
  nand_x1_sg U13452 ( .A(n6470), .B(n4368), .X(n4367) );
  nand_x1_sg U13453 ( .A(n6424), .B(n5736), .X(n4368) );
  nand_x1_sg U13454 ( .A(n6140), .B(n4332), .X(n4331) );
  nand_x1_sg U13455 ( .A(n7126), .B(n5902), .X(n4332) );
  nand_x1_sg U13456 ( .A(n7314), .B(n4296), .X(n4295) );
  nand_x1_sg U13457 ( .A(n6195), .B(n5883), .X(n4296) );
  nand_x1_sg U13458 ( .A(n4879), .B(n5985), .X(n4876) );
  nand_x1_sg U13459 ( .A(n4878), .B(n6329), .X(n4877) );
  nand_x1_sg U13460 ( .A(n7067), .B(n5655), .X(n4854) );
  nand_x1_sg U13461 ( .A(n7066), .B(n5872), .X(n4815) );
  nand_x1_sg U13462 ( .A(n6497), .B(n5899), .X(n4779) );
  nand_x1_sg U13463 ( .A(n6501), .B(n5660), .X(n4743) );
  nand_x1_sg U13464 ( .A(n6500), .B(n5770), .X(n4707) );
  nand_x1_sg U13465 ( .A(n6500), .B(n5765), .X(n4671) );
  nand_x1_sg U13466 ( .A(n6501), .B(n5665), .X(n4635) );
  nand_x1_sg U13467 ( .A(n6005), .B(n5825), .X(n4599) );
  nand_x1_sg U13468 ( .A(n6004), .B(n5778), .X(n4563) );
  nand_x1_sg U13469 ( .A(n7065), .B(n5675), .X(n4419) );
  nand_x1_sg U13470 ( .A(n7064), .B(n5889), .X(n4383) );
  nand_x1_sg U13471 ( .A(n6501), .B(n5830), .X(n4347) );
  nand_x1_sg U13472 ( .A(n6497), .B(n5768), .X(n4275) );
  nand_x1_sg U13473 ( .A(n7064), .B(n5813), .X(n4239) );
  nand_x1_sg U13474 ( .A(n6502), .B(n5685), .X(n4203) );
  nand_x1_sg U13475 ( .A(n7067), .B(n5831), .X(n4167) );
  nand_x1_sg U13476 ( .A(n6423), .B(n5731), .X(n4526) );
  nand_x1_sg U13477 ( .A(n6194), .B(n5840), .X(n4490) );
  nand_x1_sg U13478 ( .A(n6424), .B(n5755), .X(n4454) );
  nand_x1_sg U13479 ( .A(n6312), .B(n3477), .X(n3476) );
  nand_x1_sg U13480 ( .A(n6487), .B(n3462), .X(n3475) );
  nand_x1_sg U13481 ( .A(n3464), .B(n3478), .X(n3477) );
  nand_x1_sg U13482 ( .A(n6031), .B(n5886), .X(n4838) );
  nand_x1_sg U13483 ( .A(n6423), .B(n5716), .X(n4800) );
  nand_x1_sg U13484 ( .A(n7125), .B(n5862), .X(n4764) );
  nand_x1_sg U13485 ( .A(n6195), .B(n5879), .X(n4728) );
  nand_x1_sg U13486 ( .A(n7123), .B(n5722), .X(n4692) );
  nand_x1_sg U13487 ( .A(n7126), .B(n5841), .X(n4656) );
  nand_x1_sg U13488 ( .A(n7123), .B(n5885), .X(n4620) );
  nand_x1_sg U13489 ( .A(n6423), .B(n5728), .X(n4584) );
  nand_x1_sg U13490 ( .A(n7125), .B(n5868), .X(n4548) );
  nand_x1_sg U13491 ( .A(n6195), .B(n5844), .X(n4512) );
  nand_x1_sg U13492 ( .A(n7124), .B(n5732), .X(n4476) );
  nand_x1_sg U13493 ( .A(n6032), .B(n5904), .X(n4440) );
  nand_x1_sg U13494 ( .A(n6032), .B(n5740), .X(n4260) );
  nand_x1_sg U13495 ( .A(n6031), .B(n5842), .X(n4224) );
  nand_x1_sg U13496 ( .A(n7124), .B(n5882), .X(n4188) );
  nand_x1_sg U13497 ( .A(n6032), .B(n5712), .X(n4150) );
  nand_x1_sg U13498 ( .A(n7439), .B(n6332), .X(n3467) );
  nand_x1_sg U13499 ( .A(n3462), .B(n7400), .X(n3468) );
  nand_x1_sg U13500 ( .A(n7006), .B(n3442), .X(n3441) );
  nand_x1_sg U13501 ( .A(n6313), .B(\update_output_0/N28 ), .X(n3442) );
  nand_x1_sg U13502 ( .A(n7007), .B(n3456), .X(n3455) );
  nand_x1_sg U13503 ( .A(n6313), .B(n3443), .X(n3454) );
  nand_x1_sg U13504 ( .A(n7459), .B(n7300), .X(n3456) );
  nand_x1_sg U13505 ( .A(n4860), .B(n7008), .X(n4859) );
  nand_x1_sg U13506 ( .A(n6096), .B(n3443), .X(n4858) );
  nor_x1_sg U13507 ( .A(n6096), .B(n6457), .X(n4860) );
  nor_x1_sg U13508 ( .A(n6330), .B(reset), .X(n5635) );
  nor_x1_sg U13509 ( .A(reset), .B(n5634), .X(n5632) );
  nor_x1_sg U13510 ( .A(\update_mask_0/n1835 ), .B(n4872), .X(n5634) );
  nand_x1_sg U13511 ( .A(n7452), .B(\update_mask_0/N30 ), .X(n5618) );
  nand_x1_sg U13512 ( .A(n6461), .B(n5620), .X(n5619) );
  nand_x1_sg U13513 ( .A(n5621), .B(n5622), .X(n5620) );
  nor_x1_sg U13514 ( .A(reset), .B(n6460), .X(n5607) );
  nand_x1_sg U13515 ( .A(n6462), .B(n6376), .X(n5599) );
  nand_x1_sg U13516 ( .A(\update_mask_0/N25 ), .B(n9229), .X(n5600) );
  nand_x1_sg U13517 ( .A(\update_mask_0/N27 ), .B(n4873), .X(n4868) );
  nor_x1_sg U13518 ( .A(n6307), .B(n4872), .X(n4870) );
  nor_x1_sg U13519 ( .A(n5617), .B(n5631), .X(n5629) );
  nand_x1_sg U13520 ( .A(\update_mask_0/N28 ), .B(n7440), .X(n5631) );
  nand_x1_sg U13521 ( .A(n7452), .B(\update_mask_0/N29 ), .X(n5628) );
  nor_x1_sg U13522 ( .A(n5629), .B(n9230), .X(n5627) );
  nand_x1_sg U13523 ( .A(n5605), .B(n6461), .X(n5604) );
  nand_x1_sg U13524 ( .A(n6308), .B(n4875), .X(n5603) );
  nor_x1_sg U13525 ( .A(\update_mask_0/N26 ), .B(n7460), .X(n5605) );
  nand_x1_sg U13526 ( .A(n9228), .B(n7394), .X(n5616) );
  nand_x1_sg U13527 ( .A(n7452), .B(n6100), .X(n5615) );
  nand_x1_sg U13528 ( .A(n4865), .B(n4866), .X(\update_mask_0/n1442 ) );
  nand_x1_sg U13529 ( .A(n9232), .B(\update_mask_0/N23 ), .X(n4866) );
  inv_x1_sg U13530 ( .A(n4867), .X(n9232) );
  nor_x1_sg U13531 ( .A(\update_mask_0/N25 ), .B(n7389), .X(n2251) );
  nand_x1_sg U13532 ( .A(n3432), .B(n3433), .X(\update_output_0/n3151 ) );
  nand_x1_sg U13533 ( .A(n3434), .B(n6369), .X(n3433) );
  nor_x1_sg U13534 ( .A(n7006), .B(n3436), .X(n3434) );
  nor_x1_sg U13535 ( .A(\update_mask_0/N27 ), .B(n6540), .X(n4871) );
  nor_x1_sg U13536 ( .A(\mask_state[0] ), .B(n7447), .X(n2191) );
  nand_x1_sg U13537 ( .A(n2180), .B(\update_mask_0/N30 ), .X(n5611) );
  nand_x1_sg U13538 ( .A(n3446), .B(\update_output_0/n6096 ), .X(n3445) );
  nand_x1_sg U13539 ( .A(n9239), .B(n9227), .X(n3444) );
  nor_x1_sg U13540 ( .A(n3447), .B(n3436), .X(n3446) );
  nor_x1_sg U13541 ( .A(n3449), .B(n3450), .X(\update_output_0/n3148 ) );
  nor_x1_sg U13542 ( .A(n6095), .B(n3436), .X(n3449) );
  nand_x1_sg U13543 ( .A(n3448), .B(n9227), .X(n3450) );
  nand_x1_sg U13544 ( .A(n5642), .B(n7402), .X(n5640) );
  nand_x1_sg U13545 ( .A(n6329), .B(\update_output_0/n6096 ), .X(n5641) );
  nor_x1_sg U13546 ( .A(state[1]), .B(\output_state[0] ), .X(n5642) );
  nor_x1_sg U13547 ( .A(reset), .B(n5636), .X(n20) );
  nor_x1_sg U13548 ( .A(n5637), .B(n5638), .X(n5636) );
  nor_x1_sg U13549 ( .A(n9233), .B(n5643), .X(n5637) );
  nor_x1_sg U13550 ( .A(n5639), .B(n9235), .X(n5638) );
  nand_x1_sg U13551 ( .A(state[0]), .B(n6330), .X(n5649) );
  nor_x1_sg U13552 ( .A(reset), .B(n5644), .X(n19) );
  nor_x1_sg U13553 ( .A(n5645), .B(n5646), .X(n5644) );
  nor_x1_sg U13554 ( .A(n5647), .B(n9236), .X(n5646) );
  nor_x1_sg U13555 ( .A(n5648), .B(n5649), .X(n5645) );
  nand_x1_sg U13556 ( .A(n5650), .B(\update_output_0/n6096 ), .X(n5648) );
  nor_x1_sg U13557 ( .A(n6095), .B(n6310), .X(n5650) );
  nor_x1_sg U13558 ( .A(n7396), .B(\update_mask_0/N29 ), .X(n5623) );
  nor_x1_sg U13559 ( .A(n7440), .B(\update_mask_0/N28 ), .X(n5626) );
  nor_x1_sg U13560 ( .A(n6095), .B(n9234), .X(n3447) );
  nand_x1_sg U13561 ( .A(\update_mask_0/N30 ), .B(n7394), .X(n5622) );
  inv_x1_sg U13562 ( .A(state[0]), .X(n9235) );
  nor_x1_sg U13563 ( .A(state[0]), .B(n9234), .X(n5647) );
  inv_x1_sg U13564 ( .A(state[1]), .X(n9236) );
  nor_x1_sg U13565 ( .A(n6309), .B(n6366), .X(n2265) );
  nor_x1_sg U13566 ( .A(n6509), .B(n6333), .X(n761) );
  nor_x1_sg U13567 ( .A(n6367), .B(n6098), .X(n2254) );
  nor_x1_sg U13568 ( .A(n6327), .B(n6308), .X(n1480) );
  nor_x1_sg U13569 ( .A(n6327), .B(n6307), .X(n1491) );
  nor_x1_sg U13570 ( .A(n6330), .B(n4884), .X(n2189) );
  nor_x1_sg U13571 ( .A(n6308), .B(n7407), .X(n1498) );
  nor_x1_sg U13572 ( .A(n6098), .B(n7403), .X(n2261) );
  nor_x1_sg U13573 ( .A(\update_mask_0/N29 ), .B(n6101), .X(n2186) );
  nor_x1_sg U13574 ( .A(n6327), .B(n2211), .X(n2194) );
  nand_x4_sg U13575 ( .A(n2219), .B(n2220), .X(n2212) );
  nand_x4_sg U13576 ( .A(n2214), .B(n2215), .X(n2213) );
  nand_x1_sg U13577 ( .A(n6312), .B(n7373), .X(n765) );
  nor_x1_sg U13578 ( .A(n6308), .B(n2203), .X(n2201) );
  nor_x1_sg U13579 ( .A(\update_mask_0/reg_i_mask[5] ), .B(n6348), .X(n2203)
         );
  nor_x1_sg U13580 ( .A(\update_mask_0/N25 ), .B(\update_mask_0/N23 ), .X(
        n2252) );
  nor_x1_sg U13581 ( .A(n6347), .B(\update_mask_0/reg_i_mask[29] ), .X(n2260)
         );
  nor_x1_sg U13582 ( .A(n6347), .B(\update_mask_0/reg_i_mask[13] ), .X(n2224)
         );
  nor_x1_sg U13583 ( .A(n6433), .B(\update_mask_0/reg_out[0][0] ), .X(n1563)
         );
  nor_x1_sg U13584 ( .A(n6179), .B(\update_mask_0/reg_out[0][1] ), .X(n1580)
         );
  nor_x1_sg U13585 ( .A(n7099), .B(\update_mask_0/reg_out[0][5] ), .X(n1731)
         );
  nor_x1_sg U13586 ( .A(n6016), .B(\update_mask_0/reg_out[0][6] ), .X(n1748)
         );
  nor_x1_sg U13587 ( .A(n7099), .B(\update_mask_0/reg_out[0][9] ), .X(n1846)
         );
  nor_x1_sg U13588 ( .A(n6180), .B(\update_mask_0/reg_out[0][10] ), .X(n1901)
         );
  nor_x1_sg U13589 ( .A(n7098), .B(\update_mask_0/reg_out[0][11] ), .X(n1918)
         );
  nor_x1_sg U13590 ( .A(n6179), .B(\update_mask_0/reg_out[0][15] ), .X(n2069)
         );
  nor_x1_sg U13591 ( .A(n6017), .B(\update_mask_0/reg_out[0][16] ), .X(n2086)
         );
  nor_x1_sg U13592 ( .A(n7101), .B(\update_mask_0/reg_out[0][19] ), .X(n2185)
         );
  nor_x1_sg U13593 ( .A(n6384), .B(\update_mask_0/reg_i_mask[4] ), .X(n2207)
         );
  nand_x1_sg U13594 ( .A(n2227), .B(n6327), .X(n2192) );
  nor_x1_sg U13595 ( .A(n6374), .B(\update_mask_0/reg_i_mask[1] ), .X(n2210)
         );
  nor_x1_sg U13596 ( .A(\update_mask_0/reg_out[12][8] ), .B(n6435), .X(n1780)
         );
  nor_x1_sg U13597 ( .A(\update_mask_0/reg_out[8][8] ), .B(n6180), .X(n1779)
         );
  nor_x1_sg U13598 ( .A(\update_mask_0/reg_out[12][18] ), .B(n6013), .X(n2118)
         );
  nor_x1_sg U13599 ( .A(\update_mask_0/reg_out[8][18] ), .B(n6433), .X(n2117)
         );
  nor_x1_sg U13600 ( .A(\update_mask_0/reg_out[5][0] ), .B(n7055), .X(n1565)
         );
  nor_x1_sg U13601 ( .A(\update_mask_0/reg_out[1][0] ), .B(n6167), .X(n1564)
         );
  nor_x1_sg U13602 ( .A(\update_mask_0/reg_out[5][1] ), .B(n7054), .X(n1582)
         );
  nor_x1_sg U13603 ( .A(\update_mask_0/reg_out[1][1] ), .B(n6167), .X(n1581)
         );
  nor_x1_sg U13604 ( .A(\update_mask_0/reg_out[15][1] ), .B(n6479), .X(n1589)
         );
  nor_x1_sg U13605 ( .A(\update_mask_0/reg_out[11][1] ), .B(n6385), .X(n1588)
         );
  nor_x1_sg U13606 ( .A(\update_mask_0/reg_out[9][1] ), .B(n6167), .X(n1592)
         );
  nor_x1_sg U13607 ( .A(\update_mask_0/reg_out[10][1] ), .B(n7089), .X(n1597)
         );
  nor_x1_sg U13608 ( .A(\update_mask_0/reg_out[10][4] ), .B(n7090), .X(n1648)
         );
  nor_x1_sg U13609 ( .A(\update_mask_0/reg_out[13][4] ), .B(n7055), .X(n1647)
         );
  nor_x1_sg U13610 ( .A(\update_mask_0/reg_out[10][2] ), .B(n6011), .X(n1665)
         );
  nor_x1_sg U13611 ( .A(\update_mask_0/reg_out[13][2] ), .B(n6164), .X(n1664)
         );
  nor_x1_sg U13612 ( .A(\update_mask_0/reg_out[6][4] ), .B(n6074), .X(n1671)
         );
  nor_x1_sg U13613 ( .A(\update_mask_0/reg_out[2][4] ), .B(n6010), .X(n1670)
         );
  nor_x1_sg U13614 ( .A(\update_mask_0/reg_out[7][4] ), .B(n6476), .X(n1673)
         );
  nor_x1_sg U13615 ( .A(\update_mask_0/reg_out[4][4] ), .B(n7094), .X(n1676)
         );
  nor_x1_sg U13616 ( .A(\update_mask_0/reg_out[5][4] ), .B(n7054), .X(n1680)
         );
  nor_x1_sg U13617 ( .A(\update_mask_0/reg_out[5][5] ), .B(n7057), .X(n1733)
         );
  nor_x1_sg U13618 ( .A(\update_mask_0/reg_out[1][5] ), .B(n6002), .X(n1732)
         );
  nor_x1_sg U13619 ( .A(\update_mask_0/reg_out[5][6] ), .B(n6444), .X(n1750)
         );
  nor_x1_sg U13620 ( .A(\update_mask_0/reg_out[1][6] ), .B(n7061), .X(n1749)
         );
  nor_x1_sg U13621 ( .A(\update_mask_0/reg_out[15][6] ), .B(n6137), .X(n1757)
         );
  nor_x1_sg U13622 ( .A(\update_mask_0/reg_out[11][6] ), .B(n7306), .X(n1756)
         );
  nor_x1_sg U13623 ( .A(\update_mask_0/reg_out[9][6] ), .B(n7061), .X(n1760)
         );
  nor_x1_sg U13624 ( .A(\update_mask_0/reg_out[10][6] ), .B(n6438), .X(n1765)
         );
  nor_x1_sg U13625 ( .A(\update_mask_0/reg_out[15][9] ), .B(n6475), .X(n1808)
         );
  nor_x1_sg U13626 ( .A(\update_mask_0/reg_out[11][9] ), .B(n7305), .X(n1807)
         );
  nor_x1_sg U13627 ( .A(\update_mask_0/reg_out[9][9] ), .B(n7062), .X(n1811)
         );
  nor_x1_sg U13628 ( .A(\update_mask_0/reg_out[10][9] ), .B(n6011), .X(n1816)
         );
  nor_x1_sg U13629 ( .A(\update_mask_0/reg_out[15][7] ), .B(n6480), .X(n1825)
         );
  nor_x1_sg U13630 ( .A(\update_mask_0/reg_out[11][7] ), .B(n6483), .X(n1824)
         );
  nor_x1_sg U13631 ( .A(\update_mask_0/reg_out[9][7] ), .B(n7059), .X(n1828)
         );
  nor_x1_sg U13632 ( .A(\update_mask_0/reg_out[10][7] ), .B(n7089), .X(n1833)
         );
  nor_x1_sg U13633 ( .A(\update_mask_0/reg_out[6][9] ), .B(n6395), .X(n1839)
         );
  nor_x1_sg U13634 ( .A(\update_mask_0/reg_out[2][9] ), .B(n6174), .X(n1838)
         );
  nor_x1_sg U13635 ( .A(\update_mask_0/reg_out[7][9] ), .B(n7311), .X(n1841)
         );
  nor_x1_sg U13636 ( .A(\update_mask_0/reg_out[5][10] ), .B(n7056), .X(n1903)
         );
  nor_x1_sg U13637 ( .A(\update_mask_0/reg_out[1][10] ), .B(n7061), .X(n1902)
         );
  nor_x1_sg U13638 ( .A(\update_mask_0/reg_out[5][11] ), .B(n6443), .X(n1920)
         );
  nor_x1_sg U13639 ( .A(\update_mask_0/reg_out[1][11] ), .B(n7062), .X(n1919)
         );
  nor_x1_sg U13640 ( .A(\update_mask_0/reg_out[15][11] ), .B(n6478), .X(n1927)
         );
  nor_x1_sg U13641 ( .A(\update_mask_0/reg_out[11][11] ), .B(n7303), .X(n1926)
         );
  nor_x1_sg U13642 ( .A(\update_mask_0/reg_out[9][11] ), .B(n6441), .X(n1930)
         );
  nor_x1_sg U13643 ( .A(\update_mask_0/reg_out[10][11] ), .B(n6010), .X(n1935)
         );
  nor_x1_sg U13644 ( .A(\update_mask_0/reg_out[10][14] ), .B(n6011), .X(n1986)
         );
  nor_x1_sg U13645 ( .A(\update_mask_0/reg_out[13][14] ), .B(n7056), .X(n1985)
         );
  nor_x1_sg U13646 ( .A(\update_mask_0/reg_out[10][12] ), .B(n6438), .X(n2003)
         );
  nor_x1_sg U13647 ( .A(\update_mask_0/reg_out[13][12] ), .B(n5999), .X(n2002)
         );
  nor_x1_sg U13648 ( .A(\update_mask_0/reg_out[6][14] ), .B(n7226), .X(n2009)
         );
  nor_x1_sg U13649 ( .A(\update_mask_0/reg_out[2][14] ), .B(n6173), .X(n2008)
         );
  nor_x1_sg U13650 ( .A(\update_mask_0/reg_out[7][14] ), .B(n7308), .X(n2011)
         );
  nor_x1_sg U13651 ( .A(\update_mask_0/reg_out[4][14] ), .B(n6436), .X(n2014)
         );
  nor_x1_sg U13652 ( .A(\update_mask_0/reg_out[5][14] ), .B(n6164), .X(n2018)
         );
  nor_x1_sg U13653 ( .A(\update_mask_0/reg_out[5][15] ), .B(n6443), .X(n2071)
         );
  nor_x1_sg U13654 ( .A(\update_mask_0/reg_out[1][15] ), .B(n6168), .X(n2070)
         );
  nor_x1_sg U13655 ( .A(\update_mask_0/reg_out[5][16] ), .B(n6444), .X(n2088)
         );
  nor_x1_sg U13656 ( .A(\update_mask_0/reg_out[1][16] ), .B(n6003), .X(n2087)
         );
  nor_x1_sg U13657 ( .A(\update_mask_0/reg_out[15][16] ), .B(n7311), .X(n2095)
         );
  nor_x1_sg U13658 ( .A(\update_mask_0/reg_out[11][16] ), .B(n6484), .X(n2094)
         );
  nor_x1_sg U13659 ( .A(\update_mask_0/reg_out[9][16] ), .B(n6442), .X(n2098)
         );
  nor_x1_sg U13660 ( .A(\update_mask_0/reg_out[10][16] ), .B(n6011), .X(n2103)
         );
  nor_x1_sg U13661 ( .A(\update_mask_0/reg_out[15][19] ), .B(n6479), .X(n2146)
         );
  nor_x1_sg U13662 ( .A(\update_mask_0/reg_out[11][19] ), .B(n6482), .X(n2145)
         );
  nor_x1_sg U13663 ( .A(\update_mask_0/reg_out[9][19] ), .B(n6002), .X(n2149)
         );
  nor_x1_sg U13664 ( .A(\update_mask_0/reg_out[10][19] ), .B(n6173), .X(n2154)
         );
  nor_x1_sg U13665 ( .A(\update_mask_0/reg_out[15][17] ), .B(n7308), .X(n2163)
         );
  nor_x1_sg U13666 ( .A(\update_mask_0/reg_out[11][17] ), .B(n6134), .X(n2162)
         );
  nor_x1_sg U13667 ( .A(\update_mask_0/reg_out[9][17] ), .B(n6003), .X(n2166)
         );
  nor_x1_sg U13668 ( .A(\update_mask_0/reg_out[10][17] ), .B(n6173), .X(n2171)
         );
  nor_x1_sg U13669 ( .A(\update_mask_0/reg_out[6][19] ), .B(n6396), .X(n2177)
         );
  nor_x1_sg U13670 ( .A(\update_mask_0/reg_out[2][19] ), .B(n6438), .X(n2176)
         );
  nor_x1_sg U13671 ( .A(\update_mask_0/reg_out[7][19] ), .B(n6138), .X(n2179)
         );
  nor_x1_sg U13672 ( .A(\update_mask_0/reg_i_mask[18] ), .B(n7442), .X(n2235)
         );
  nor_x1_sg U13673 ( .A(\update_mask_0/reg_i_mask[17] ), .B(n1455), .X(n2234)
         );
  nor_x1_sg U13674 ( .A(\update_mask_0/reg_i_mask[20] ), .B(n6383), .X(n2237)
         );
  nor_x1_sg U13675 ( .A(\update_mask_0/reg_i_mask[22] ), .B(n6353), .X(n2240)
         );
  nor_x1_sg U13676 ( .A(\update_mask_0/reg_i_mask[16] ), .B(n6371), .X(n2244)
         );
  nor_x1_sg U13677 ( .A(\update_mask_0/reg_i_mask[28] ), .B(n7446), .X(n2253)
         );
  nor_x1_sg U13678 ( .A(\update_mask_0/reg_i_mask[27] ), .B(n6377), .X(n2250)
         );
  nor_x1_sg U13679 ( .A(n6354), .B(\update_mask_0/reg_i_mask[30] ), .X(n2259)
         );
  nor_x1_sg U13680 ( .A(n6353), .B(\update_mask_0/reg_i_mask[14] ), .X(n2223)
         );
  nor_x1_sg U13681 ( .A(n7062), .B(\update_mask_0/reg_out[1][2] ), .X(n1519)
         );
  nor_x1_sg U13682 ( .A(n6443), .B(\update_mask_0/reg_out[5][2] ), .X(n1518)
         );
  nor_x1_sg U13683 ( .A(n6386), .B(\update_mask_0/reg_out[3][2] ), .X(n1531)
         );
  nor_x1_sg U13684 ( .A(n7308), .B(\update_mask_0/reg_out[7][2] ), .X(n1530)
         );
  nor_x1_sg U13685 ( .A(n6437), .B(\update_mask_0/reg_out[2][2] ), .X(n1533)
         );
  nor_x1_sg U13686 ( .A(n7224), .B(\update_mask_0/reg_out[6][2] ), .X(n1532)
         );
  nor_x1_sg U13687 ( .A(n7056), .B(\update_mask_0/reg_out[13][0] ), .X(n1540)
         );
  nor_x1_sg U13688 ( .A(n7091), .B(\update_mask_0/reg_out[10][0] ), .X(n1539)
         );
  nor_x1_sg U13689 ( .A(n6475), .B(\update_mask_0/reg_out[15][0] ), .X(n1548)
         );
  nor_x1_sg U13690 ( .A(n6073), .B(\update_mask_0/reg_out[14][0] ), .X(n1550)
         );
  nor_x1_sg U13691 ( .A(n7098), .B(\update_mask_0/reg_out[8][4] ), .X(n1646)
         );
  nor_x1_sg U13692 ( .A(n7093), .B(\update_mask_0/reg_out[12][4] ), .X(n1645)
         );
  nor_x1_sg U13693 ( .A(n6443), .B(\update_mask_0/reg_out[13][3] ), .X(n1608)
         );
  nor_x1_sg U13694 ( .A(n7088), .B(\update_mask_0/reg_out[10][3] ), .X(n1607)
         );
  nor_x1_sg U13695 ( .A(n6138), .B(\update_mask_0/reg_out[15][3] ), .X(n1616)
         );
  nor_x1_sg U13696 ( .A(n6074), .B(\update_mask_0/reg_out[14][3] ), .X(n1618)
         );
  nor_x1_sg U13697 ( .A(n7306), .B(\update_mask_0/reg_out[11][3] ), .X(n1617)
         );
  nor_x1_sg U13698 ( .A(n6168), .B(\update_mask_0/reg_out[1][3] ), .X(n1623)
         );
  nor_x1_sg U13699 ( .A(n6165), .B(\update_mask_0/reg_out[5][3] ), .X(n1622)
         );
  nor_x1_sg U13700 ( .A(n6385), .B(\update_mask_0/reg_out[3][3] ), .X(n1631)
         );
  nor_x1_sg U13701 ( .A(n6138), .B(\update_mask_0/reg_out[7][3] ), .X(n1630)
         );
  nor_x1_sg U13702 ( .A(n7090), .B(\update_mask_0/reg_out[2][3] ), .X(n1633)
         );
  nor_x1_sg U13703 ( .A(n6180), .B(\update_mask_0/reg_out[8][2] ), .X(n1663)
         );
  nor_x1_sg U13704 ( .A(n6176), .B(\update_mask_0/reg_out[12][2] ), .X(n1662)
         );
  nor_x1_sg U13705 ( .A(n7062), .B(\update_mask_0/reg_out[1][7] ), .X(n1693)
         );
  nor_x1_sg U13706 ( .A(n7054), .B(\update_mask_0/reg_out[5][7] ), .X(n1692)
         );
  nor_x1_sg U13707 ( .A(n7304), .B(\update_mask_0/reg_out[3][7] ), .X(n1701)
         );
  nor_x1_sg U13708 ( .A(n6137), .B(\update_mask_0/reg_out[7][7] ), .X(n1700)
         );
  nor_x1_sg U13709 ( .A(n6174), .B(\update_mask_0/reg_out[2][7] ), .X(n1703)
         );
  nor_x1_sg U13710 ( .A(n6395), .B(\update_mask_0/reg_out[6][7] ), .X(n1702)
         );
  nor_x1_sg U13711 ( .A(n6165), .B(\update_mask_0/reg_out[13][5] ), .X(n1708)
         );
  nor_x1_sg U13712 ( .A(n6437), .B(\update_mask_0/reg_out[10][5] ), .X(n1707)
         );
  nor_x1_sg U13713 ( .A(n7309), .B(\update_mask_0/reg_out[15][5] ), .X(n1716)
         );
  nor_x1_sg U13714 ( .A(n7226), .B(\update_mask_0/reg_out[14][5] ), .X(n1718)
         );
  nor_x1_sg U13715 ( .A(n6167), .B(\update_mask_0/reg_out[1][8] ), .X(n1791)
         );
  nor_x1_sg U13716 ( .A(n5999), .B(\update_mask_0/reg_out[5][8] ), .X(n1790)
         );
  nor_x1_sg U13717 ( .A(n6135), .B(\update_mask_0/reg_out[3][8] ), .X(n1799)
         );
  nor_x1_sg U13718 ( .A(n6478), .B(\update_mask_0/reg_out[7][8] ), .X(n1798)
         );
  nor_x1_sg U13719 ( .A(n6010), .B(\update_mask_0/reg_out[2][8] ), .X(n1801)
         );
  nor_x1_sg U13720 ( .A(n6233), .B(\update_mask_0/reg_out[6][8] ), .X(n1800)
         );
  nor_x1_sg U13721 ( .A(n7059), .B(\update_mask_0/reg_out[1][12] ), .X(n1863)
         );
  nor_x1_sg U13722 ( .A(n6444), .B(\update_mask_0/reg_out[5][12] ), .X(n1862)
         );
  nor_x1_sg U13723 ( .A(n7306), .B(\update_mask_0/reg_out[3][12] ), .X(n1871)
         );
  nor_x1_sg U13724 ( .A(n7310), .B(\update_mask_0/reg_out[7][12] ), .X(n1870)
         );
  nor_x1_sg U13725 ( .A(n7088), .B(\update_mask_0/reg_out[2][12] ), .X(n1873)
         );
  nor_x1_sg U13726 ( .A(n6395), .B(\update_mask_0/reg_out[6][12] ), .X(n1872)
         );
  nor_x1_sg U13727 ( .A(n6000), .B(\update_mask_0/reg_out[13][10] ), .X(n1878)
         );
  nor_x1_sg U13728 ( .A(n6437), .B(\update_mask_0/reg_out[10][10] ), .X(n1877)
         );
  nor_x1_sg U13729 ( .A(n7310), .B(\update_mask_0/reg_out[15][10] ), .X(n1886)
         );
  nor_x1_sg U13730 ( .A(n6395), .B(\update_mask_0/reg_out[14][10] ), .X(n1888)
         );
  nor_x1_sg U13731 ( .A(n6434), .B(\update_mask_0/reg_out[8][14] ), .X(n1984)
         );
  nor_x1_sg U13732 ( .A(n7093), .B(\update_mask_0/reg_out[12][14] ), .X(n1983)
         );
  nor_x1_sg U13733 ( .A(n7057), .B(\update_mask_0/reg_out[13][13] ), .X(n1946)
         );
  nor_x1_sg U13734 ( .A(n7089), .B(\update_mask_0/reg_out[10][13] ), .X(n1945)
         );
  nor_x1_sg U13735 ( .A(n7309), .B(\update_mask_0/reg_out[15][13] ), .X(n1954)
         );
  nor_x1_sg U13736 ( .A(n7225), .B(\update_mask_0/reg_out[14][13] ), .X(n1956)
         );
  nor_x1_sg U13737 ( .A(n6483), .B(\update_mask_0/reg_out[11][13] ), .X(n1955)
         );
  nor_x1_sg U13738 ( .A(n6003), .B(\update_mask_0/reg_out[1][13] ), .X(n1961)
         );
  nor_x1_sg U13739 ( .A(n7055), .B(\update_mask_0/reg_out[5][13] ), .X(n1960)
         );
  nor_x1_sg U13740 ( .A(n6134), .B(\update_mask_0/reg_out[3][13] ), .X(n1969)
         );
  nor_x1_sg U13741 ( .A(n6475), .B(\update_mask_0/reg_out[7][13] ), .X(n1968)
         );
  nor_x1_sg U13742 ( .A(n7089), .B(\update_mask_0/reg_out[2][13] ), .X(n1971)
         );
  nor_x1_sg U13743 ( .A(n7101), .B(\update_mask_0/reg_out[8][12] ), .X(n2001)
         );
  nor_x1_sg U13744 ( .A(n6176), .B(\update_mask_0/reg_out[12][12] ), .X(n2000)
         );
  nor_x1_sg U13745 ( .A(n6441), .B(\update_mask_0/reg_out[1][17] ), .X(n2031)
         );
  nor_x1_sg U13746 ( .A(n6000), .B(\update_mask_0/reg_out[5][17] ), .X(n2030)
         );
  nor_x1_sg U13747 ( .A(n6483), .B(\update_mask_0/reg_out[3][17] ), .X(n2039)
         );
  nor_x1_sg U13748 ( .A(n6137), .B(\update_mask_0/reg_out[7][17] ), .X(n2038)
         );
  nor_x1_sg U13749 ( .A(n7090), .B(\update_mask_0/reg_out[2][17] ), .X(n2041)
         );
  nor_x1_sg U13750 ( .A(n6234), .B(\update_mask_0/reg_out[6][17] ), .X(n2040)
         );
  nor_x1_sg U13751 ( .A(n6165), .B(\update_mask_0/reg_out[13][15] ), .X(n2046)
         );
  nor_x1_sg U13752 ( .A(n7090), .B(\update_mask_0/reg_out[10][15] ), .X(n2045)
         );
  nor_x1_sg U13753 ( .A(n7310), .B(\update_mask_0/reg_out[15][15] ), .X(n2054)
         );
  nor_x1_sg U13754 ( .A(n6234), .B(\update_mask_0/reg_out[14][15] ), .X(n2056)
         );
  nor_x1_sg U13755 ( .A(n7060), .B(\update_mask_0/reg_out[1][18] ), .X(n2129)
         );
  nor_x1_sg U13756 ( .A(n6165), .B(\update_mask_0/reg_out[5][18] ), .X(n2128)
         );
  nor_x1_sg U13757 ( .A(n6386), .B(\update_mask_0/reg_out[3][18] ), .X(n2137)
         );
  nor_x1_sg U13758 ( .A(n6138), .B(\update_mask_0/reg_out[7][18] ), .X(n2136)
         );
  nor_x1_sg U13759 ( .A(n6010), .B(\update_mask_0/reg_out[2][18] ), .X(n2139)
         );
  nor_x1_sg U13760 ( .A(n6233), .B(\update_mask_0/reg_out[6][18] ), .X(n2138)
         );
  nor_x1_sg U13761 ( .A(n6541), .B(\update_mask_0/reg_i_mask[7] ), .X(n2200)
         );
  nor_x1_sg U13762 ( .A(n1452), .B(\update_mask_0/reg_i_mask[0] ), .X(n2199)
         );
  nor_x1_sg U13763 ( .A(n6378), .B(\update_mask_0/reg_i_mask[3] ), .X(n2208)
         );
  nor_x1_sg U13764 ( .A(n6380), .B(\update_mask_0/reg_i_mask[2] ), .X(n2209)
         );
  nor_x1_sg U13765 ( .A(n2218), .B(n6307), .X(n2214) );
  nor_x1_sg U13766 ( .A(\update_mask_0/reg_i_mask[12] ), .B(n6384), .X(n2218)
         );
  nand_x1_sg U13767 ( .A(n6100), .B(n2186), .X(n1520) );
  nand_x1_sg U13768 ( .A(n6100), .B(n5623), .X(n1521) );
  nor_x1_sg U13769 ( .A(n6325), .B(n1784), .X(n1783) );
  nor_x1_sg U13770 ( .A(n6476), .B(\update_mask_0/reg_out[15][8] ), .X(n1784)
         );
  nor_x1_sg U13771 ( .A(n6118), .B(n2122), .X(n2121) );
  nor_x1_sg U13772 ( .A(n6479), .B(\update_mask_0/reg_out[15][18] ), .X(n2122)
         );
  nor_x1_sg U13773 ( .A(n1640), .B(n7013), .X(n1636) );
  nor_x1_sg U13774 ( .A(\update_mask_0/reg_out[15][4] ), .B(n6476), .X(n1640)
         );
  nor_x1_sg U13775 ( .A(n1657), .B(n7011), .X(n1653) );
  nor_x1_sg U13776 ( .A(\update_mask_0/reg_out[15][2] ), .B(n7311), .X(n1657)
         );
  nor_x1_sg U13777 ( .A(n1978), .B(n6325), .X(n1974) );
  nor_x1_sg U13778 ( .A(\update_mask_0/reg_out[15][14] ), .B(n6478), .X(n1978)
         );
  nor_x1_sg U13779 ( .A(n1995), .B(n7014), .X(n1991) );
  nor_x1_sg U13780 ( .A(\update_mask_0/reg_out[15][12] ), .B(n6479), .X(n1995)
         );
  nor_x1_sg U13781 ( .A(n1785), .B(n1786), .X(n1782) );
  nor_x1_sg U13782 ( .A(n6385), .B(\update_mask_0/reg_out[11][8] ), .X(n1785)
         );
  nor_x1_sg U13783 ( .A(n7225), .B(\update_mask_0/reg_out[14][8] ), .X(n1786)
         );
  nor_x1_sg U13784 ( .A(n2123), .B(n2124), .X(n2120) );
  nor_x1_sg U13785 ( .A(n7305), .B(\update_mask_0/reg_out[11][18] ), .X(n2123)
         );
  nor_x1_sg U13786 ( .A(n7227), .B(\update_mask_0/reg_out[14][18] ), .X(n2124)
         );
  nor_x1_sg U13787 ( .A(n1543), .B(n1544), .X(n1541) );
  nor_x1_sg U13788 ( .A(\update_mask_0/reg_out[8][0] ), .B(n6016), .X(n1543)
         );
  nor_x1_sg U13789 ( .A(\update_mask_0/reg_out[12][0] ), .B(n6436), .X(n1544)
         );
  nor_x1_sg U13790 ( .A(n1611), .B(n1612), .X(n1609) );
  nor_x1_sg U13791 ( .A(\update_mask_0/reg_out[8][3] ), .B(n6017), .X(n1611)
         );
  nor_x1_sg U13792 ( .A(\update_mask_0/reg_out[12][3] ), .B(n6177), .X(n1612)
         );
  nor_x1_sg U13793 ( .A(n1711), .B(n1712), .X(n1709) );
  nor_x1_sg U13794 ( .A(\update_mask_0/reg_out[8][5] ), .B(n7099), .X(n1711)
         );
  nor_x1_sg U13795 ( .A(\update_mask_0/reg_out[12][5] ), .B(n7093), .X(n1712)
         );
  nor_x1_sg U13796 ( .A(n1881), .B(n1882), .X(n1879) );
  nor_x1_sg U13797 ( .A(\update_mask_0/reg_out[8][10] ), .B(n6017), .X(n1881)
         );
  nor_x1_sg U13798 ( .A(\update_mask_0/reg_out[12][10] ), .B(n6435), .X(n1882)
         );
  nor_x1_sg U13799 ( .A(n1949), .B(n1950), .X(n1947) );
  nor_x1_sg U13800 ( .A(\update_mask_0/reg_out[8][13] ), .B(n6179), .X(n1949)
         );
  nor_x1_sg U13801 ( .A(\update_mask_0/reg_out[12][13] ), .B(n6436), .X(n1950)
         );
  nor_x1_sg U13802 ( .A(n2049), .B(n2050), .X(n2047) );
  nor_x1_sg U13803 ( .A(\update_mask_0/reg_out[8][15] ), .B(n6016), .X(n2049)
         );
  nor_x1_sg U13804 ( .A(\update_mask_0/reg_out[12][15] ), .B(n6014), .X(n2050)
         );
  nor_x1_sg U13805 ( .A(n1555), .B(n1556), .X(n1554) );
  nor_x1_sg U13806 ( .A(\update_mask_0/reg_out[2][0] ), .B(n6438), .X(n1555)
         );
  nor_x1_sg U13807 ( .A(\update_mask_0/reg_out[6][0] ), .B(n6233), .X(n1556)
         );
  nor_x1_sg U13808 ( .A(n1557), .B(n1558), .X(n1553) );
  nor_x1_sg U13809 ( .A(\update_mask_0/reg_out[3][0] ), .B(n6385), .X(n1557)
         );
  nor_x1_sg U13810 ( .A(\update_mask_0/reg_out[7][0] ), .B(n7311), .X(n1558)
         );
  nand_x1_sg U13811 ( .A(n8903), .B(n7013), .X(n1562) );
  nor_x1_sg U13812 ( .A(\update_mask_0/reg_out[4][0] ), .B(n7096), .X(n1561)
         );
  nor_x1_sg U13813 ( .A(n1572), .B(n1573), .X(n1571) );
  nor_x1_sg U13814 ( .A(\update_mask_0/reg_out[2][1] ), .B(n6174), .X(n1572)
         );
  nor_x1_sg U13815 ( .A(\update_mask_0/reg_out[6][1] ), .B(n6234), .X(n1573)
         );
  nor_x1_sg U13816 ( .A(n1574), .B(n1575), .X(n1570) );
  nor_x1_sg U13817 ( .A(\update_mask_0/reg_out[3][1] ), .B(n6134), .X(n1574)
         );
  nor_x1_sg U13818 ( .A(\update_mask_0/reg_out[7][1] ), .B(n7310), .X(n1575)
         );
  nand_x1_sg U13819 ( .A(n8904), .B(n6119), .X(n1579) );
  nor_x1_sg U13820 ( .A(\update_mask_0/reg_out[4][1] ), .B(n6176), .X(n1578)
         );
  nor_x1_sg U13821 ( .A(n1638), .B(n1639), .X(n1637) );
  nor_x1_sg U13822 ( .A(\update_mask_0/reg_out[14][4] ), .B(n7226), .X(n1638)
         );
  nor_x1_sg U13823 ( .A(\update_mask_0/reg_out[11][4] ), .B(n7304), .X(n1639)
         );
  nor_x1_sg U13824 ( .A(n1643), .B(n8942), .X(n1642) );
  nor_x1_sg U13825 ( .A(\update_mask_0/reg_out[9][4] ), .B(n7059), .X(n1643)
         );
  nor_x1_sg U13826 ( .A(n1645), .B(n1646), .X(n1644) );
  nor_x1_sg U13827 ( .A(n1655), .B(n1656), .X(n1654) );
  nor_x1_sg U13828 ( .A(\update_mask_0/reg_out[14][2] ), .B(n7224), .X(n1655)
         );
  nor_x1_sg U13829 ( .A(\update_mask_0/reg_out[11][2] ), .B(n6484), .X(n1656)
         );
  nor_x1_sg U13830 ( .A(n1660), .B(n8943), .X(n1659) );
  nor_x1_sg U13831 ( .A(\update_mask_0/reg_out[9][2] ), .B(n6168), .X(n1660)
         );
  nor_x1_sg U13832 ( .A(n1662), .B(n1663), .X(n1661) );
  nor_x1_sg U13833 ( .A(n1723), .B(n1724), .X(n1722) );
  nor_x1_sg U13834 ( .A(\update_mask_0/reg_out[2][5] ), .B(n6173), .X(n1723)
         );
  nor_x1_sg U13835 ( .A(\update_mask_0/reg_out[6][5] ), .B(n6233), .X(n1724)
         );
  nor_x1_sg U13836 ( .A(n1725), .B(n1726), .X(n1721) );
  nor_x1_sg U13837 ( .A(\update_mask_0/reg_out[3][5] ), .B(n6134), .X(n1725)
         );
  nor_x1_sg U13838 ( .A(\update_mask_0/reg_out[7][5] ), .B(n6480), .X(n1726)
         );
  nand_x1_sg U13839 ( .A(n8906), .B(n6118), .X(n1730) );
  nor_x1_sg U13840 ( .A(\update_mask_0/reg_out[4][5] ), .B(n6013), .X(n1729)
         );
  nor_x1_sg U13841 ( .A(n1740), .B(n1741), .X(n1739) );
  nor_x1_sg U13842 ( .A(\update_mask_0/reg_out[2][6] ), .B(n6174), .X(n1740)
         );
  nor_x1_sg U13843 ( .A(\update_mask_0/reg_out[6][6] ), .B(n7227), .X(n1741)
         );
  nor_x1_sg U13844 ( .A(n1742), .B(n1743), .X(n1738) );
  nor_x1_sg U13845 ( .A(\update_mask_0/reg_out[3][6] ), .B(n7304), .X(n1742)
         );
  nor_x1_sg U13846 ( .A(\update_mask_0/reg_out[7][6] ), .B(n7309), .X(n1743)
         );
  nand_x1_sg U13847 ( .A(n8907), .B(n6326), .X(n1747) );
  nor_x1_sg U13848 ( .A(\update_mask_0/reg_out[4][6] ), .B(n7096), .X(n1746)
         );
  nand_x1_sg U13849 ( .A(n8908), .B(n7012), .X(n1845) );
  nor_x1_sg U13850 ( .A(\update_mask_0/reg_out[4][9] ), .B(n7096), .X(n1844)
         );
  nor_x1_sg U13851 ( .A(n1847), .B(n1848), .X(n1842) );
  nor_x1_sg U13852 ( .A(\update_mask_0/reg_out[1][9] ), .B(n7059), .X(n1847)
         );
  nor_x1_sg U13853 ( .A(\update_mask_0/reg_out[5][9] ), .B(n6000), .X(n1848)
         );
  nor_x1_sg U13854 ( .A(n1893), .B(n1894), .X(n1892) );
  nor_x1_sg U13855 ( .A(\update_mask_0/reg_out[2][10] ), .B(n7091), .X(n1893)
         );
  nor_x1_sg U13856 ( .A(\update_mask_0/reg_out[6][10] ), .B(n7225), .X(n1894)
         );
  nor_x1_sg U13857 ( .A(n1895), .B(n1896), .X(n1891) );
  nor_x1_sg U13858 ( .A(\update_mask_0/reg_out[3][10] ), .B(n6482), .X(n1895)
         );
  nor_x1_sg U13859 ( .A(\update_mask_0/reg_out[7][10] ), .B(n6137), .X(n1896)
         );
  nand_x1_sg U13860 ( .A(n8909), .B(n7012), .X(n1900) );
  nor_x1_sg U13861 ( .A(\update_mask_0/reg_out[4][10] ), .B(n6013), .X(n1899)
         );
  nor_x1_sg U13862 ( .A(n1910), .B(n1911), .X(n1909) );
  nor_x1_sg U13863 ( .A(\update_mask_0/reg_out[2][11] ), .B(n7091), .X(n1910)
         );
  nor_x1_sg U13864 ( .A(\update_mask_0/reg_out[6][11] ), .B(n6396), .X(n1911)
         );
  nor_x1_sg U13865 ( .A(n1912), .B(n1913), .X(n1908) );
  nor_x1_sg U13866 ( .A(\update_mask_0/reg_out[3][11] ), .B(n6386), .X(n1912)
         );
  nor_x1_sg U13867 ( .A(\update_mask_0/reg_out[7][11] ), .B(n6475), .X(n1913)
         );
  nand_x1_sg U13868 ( .A(n8910), .B(n6118), .X(n1917) );
  nor_x1_sg U13869 ( .A(\update_mask_0/reg_out[4][11] ), .B(n6014), .X(n1916)
         );
  nor_x1_sg U13870 ( .A(n1976), .B(n1977), .X(n1975) );
  nor_x1_sg U13871 ( .A(\update_mask_0/reg_out[14][14] ), .B(n7227), .X(n1976)
         );
  nor_x1_sg U13872 ( .A(\update_mask_0/reg_out[11][14] ), .B(n7303), .X(n1977)
         );
  nor_x1_sg U13873 ( .A(n1981), .B(n8952), .X(n1980) );
  nor_x1_sg U13874 ( .A(\update_mask_0/reg_out[9][14] ), .B(n6002), .X(n1981)
         );
  nor_x1_sg U13875 ( .A(n1983), .B(n1984), .X(n1982) );
  nor_x1_sg U13876 ( .A(n1993), .B(n1994), .X(n1992) );
  nor_x1_sg U13877 ( .A(\update_mask_0/reg_out[14][12] ), .B(n6074), .X(n1993)
         );
  nor_x1_sg U13878 ( .A(\update_mask_0/reg_out[11][12] ), .B(n7305), .X(n1994)
         );
  nor_x1_sg U13879 ( .A(n1998), .B(n8953), .X(n1997) );
  nor_x1_sg U13880 ( .A(\update_mask_0/reg_out[9][12] ), .B(n6442), .X(n1998)
         );
  nor_x1_sg U13881 ( .A(n2000), .B(n2001), .X(n1999) );
  nor_x1_sg U13882 ( .A(n2061), .B(n2062), .X(n2060) );
  nor_x1_sg U13883 ( .A(\update_mask_0/reg_out[2][15] ), .B(n7088), .X(n2061)
         );
  nor_x1_sg U13884 ( .A(\update_mask_0/reg_out[6][15] ), .B(n7227), .X(n2062)
         );
  nor_x1_sg U13885 ( .A(n2063), .B(n2064), .X(n2059) );
  nor_x1_sg U13886 ( .A(\update_mask_0/reg_out[3][15] ), .B(n6386), .X(n2063)
         );
  nor_x1_sg U13887 ( .A(\update_mask_0/reg_out[7][15] ), .B(n6480), .X(n2064)
         );
  nand_x1_sg U13888 ( .A(n8912), .B(n7011), .X(n2068) );
  nor_x1_sg U13889 ( .A(\update_mask_0/reg_out[4][15] ), .B(n6435), .X(n2067)
         );
  nor_x1_sg U13890 ( .A(n2078), .B(n2079), .X(n2077) );
  nor_x1_sg U13891 ( .A(\update_mask_0/reg_out[2][16] ), .B(n7088), .X(n2078)
         );
  nor_x1_sg U13892 ( .A(\update_mask_0/reg_out[6][16] ), .B(n7224), .X(n2079)
         );
  nor_x1_sg U13893 ( .A(n2080), .B(n2081), .X(n2076) );
  nor_x1_sg U13894 ( .A(\update_mask_0/reg_out[3][16] ), .B(n6135), .X(n2080)
         );
  nor_x1_sg U13895 ( .A(\update_mask_0/reg_out[7][16] ), .B(n6476), .X(n2081)
         );
  nand_x1_sg U13896 ( .A(n8913), .B(n7014), .X(n2085) );
  nor_x1_sg U13897 ( .A(\update_mask_0/reg_out[4][16] ), .B(n7095), .X(n2084)
         );
  nand_x1_sg U13898 ( .A(n8914), .B(n6119), .X(n2184) );
  nor_x1_sg U13899 ( .A(\update_mask_0/reg_out[4][19] ), .B(n6177), .X(n2183)
         );
  nor_x1_sg U13900 ( .A(n2187), .B(n2188), .X(n2181) );
  nor_x1_sg U13901 ( .A(\update_mask_0/reg_out[1][19] ), .B(n7060), .X(n2187)
         );
  nor_x1_sg U13902 ( .A(\update_mask_0/reg_out[5][19] ), .B(n7056), .X(n2188)
         );
  nor_x1_sg U13903 ( .A(n2257), .B(n8900), .X(n2256) );
  nor_x1_sg U13904 ( .A(\update_mask_0/reg_i_mask[31] ), .B(n6540), .X(n2257)
         );
  nor_x1_sg U13905 ( .A(n2259), .B(n2260), .X(n2258) );
  nor_x1_sg U13906 ( .A(n2263), .B(n2264), .X(n2255) );
  nor_x1_sg U13907 ( .A(\update_mask_0/reg_i_mask[24] ), .B(n6371), .X(n2263)
         );
  nor_x1_sg U13908 ( .A(\update_mask_0/reg_i_mask[25] ), .B(n6375), .X(n2264)
         );
  nor_x1_sg U13909 ( .A(n2216), .B(n2217), .X(n2215) );
  nor_x1_sg U13910 ( .A(\update_mask_0/reg_i_mask[10] ), .B(n6381), .X(n2216)
         );
  nor_x1_sg U13911 ( .A(\update_mask_0/reg_i_mask[11] ), .B(n6378), .X(n2217)
         );
  nor_x1_sg U13912 ( .A(n2221), .B(n8899), .X(n2220) );
  nor_x1_sg U13913 ( .A(\update_mask_0/reg_i_mask[15] ), .B(n6541), .X(n2221)
         );
  nor_x1_sg U13914 ( .A(n2223), .B(n2224), .X(n2222) );
  nor_x1_sg U13915 ( .A(n2225), .B(n2226), .X(n2219) );
  nor_x1_sg U13916 ( .A(\update_mask_0/reg_i_mask[8] ), .B(n6372), .X(n2225)
         );
  nor_x1_sg U13917 ( .A(\update_mask_0/reg_i_mask[9] ), .B(n1455), .X(n2226)
         );
  nor_x1_sg U13918 ( .A(n6506), .B(n1525), .X(n1522) );
  nor_x1_sg U13919 ( .A(\update_mask_0/reg_out[0][2] ), .B(n6180), .X(n1525)
         );
  nor_x1_sg U13920 ( .A(n6506), .B(n1626), .X(n1624) );
  nor_x1_sg U13921 ( .A(\update_mask_0/reg_out[0][3] ), .B(n7101), .X(n1626)
         );
  nor_x1_sg U13922 ( .A(n6506), .B(n1696), .X(n1694) );
  nor_x1_sg U13923 ( .A(\update_mask_0/reg_out[0][7] ), .B(n7100), .X(n1696)
         );
  nor_x1_sg U13924 ( .A(n6504), .B(n1794), .X(n1792) );
  nor_x1_sg U13925 ( .A(\update_mask_0/reg_out[0][8] ), .B(n6016), .X(n1794)
         );
  nor_x1_sg U13926 ( .A(n6504), .B(n1866), .X(n1864) );
  nor_x1_sg U13927 ( .A(\update_mask_0/reg_out[0][12] ), .B(n6433), .X(n1866)
         );
  nor_x1_sg U13928 ( .A(n6505), .B(n1964), .X(n1962) );
  nor_x1_sg U13929 ( .A(\update_mask_0/reg_out[0][13] ), .B(n6434), .X(n1964)
         );
  nor_x1_sg U13930 ( .A(n6504), .B(n2034), .X(n2032) );
  nor_x1_sg U13931 ( .A(\update_mask_0/reg_out[0][17] ), .B(n7098), .X(n2034)
         );
  nor_x1_sg U13932 ( .A(n6505), .B(n2132), .X(n2130) );
  nor_x1_sg U13933 ( .A(\update_mask_0/reg_out[0][18] ), .B(n6434), .X(n2132)
         );
  nand_x1_sg U13934 ( .A(n2242), .B(n7405), .X(n2241) );
  nand_x1_sg U13935 ( .A(n7392), .B(n8895), .X(n2242) );
  inv_x1_sg U13936 ( .A(\update_mask_0/reg_i_mask[21] ), .X(n8895) );
  nand_x1_sg U13937 ( .A(n8905), .B(n6325), .X(n1677) );
  nor_x1_sg U13938 ( .A(n6017), .B(\update_mask_0/reg_out[0][4] ), .X(n1678)
         );
  nand_x1_sg U13939 ( .A(n8911), .B(n7011), .X(n2015) );
  nor_x1_sg U13940 ( .A(n7099), .B(\update_mask_0/reg_out[0][14] ), .X(n2016)
         );
  nand_x1_sg U13941 ( .A(n7393), .B(n8896), .X(n2202) );
  inv_x1_sg U13942 ( .A(\update_mask_0/reg_i_mask[6] ), .X(n8896) );
  nor_x1_sg U13943 ( .A(n1549), .B(n1550), .X(n1546) );
  nor_x1_sg U13944 ( .A(n6326), .B(n1548), .X(n1547) );
  nor_x1_sg U13945 ( .A(n6483), .B(\update_mask_0/reg_out[11][0] ), .X(n1549)
         );
  nor_x1_sg U13946 ( .A(n1632), .B(n1633), .X(n1628) );
  nor_x1_sg U13947 ( .A(n1630), .B(n1631), .X(n1629) );
  nor_x1_sg U13948 ( .A(n6396), .B(\update_mask_0/reg_out[6][3] ), .X(n1632)
         );
  nor_x1_sg U13949 ( .A(n1717), .B(n1718), .X(n1714) );
  nor_x1_sg U13950 ( .A(n7011), .B(n1716), .X(n1715) );
  nor_x1_sg U13951 ( .A(n7303), .B(\update_mask_0/reg_out[11][5] ), .X(n1717)
         );
  nor_x1_sg U13952 ( .A(n1887), .B(n1888), .X(n1884) );
  nor_x1_sg U13953 ( .A(n7014), .B(n1886), .X(n1885) );
  nor_x1_sg U13954 ( .A(n6484), .B(\update_mask_0/reg_out[11][10] ), .X(n1887)
         );
  nor_x1_sg U13955 ( .A(n1970), .B(n1971), .X(n1966) );
  nor_x1_sg U13956 ( .A(n1968), .B(n1969), .X(n1967) );
  nor_x1_sg U13957 ( .A(n7224), .B(\update_mask_0/reg_out[6][13] ), .X(n1970)
         );
  nor_x1_sg U13958 ( .A(n2055), .B(n2056), .X(n2052) );
  nor_x1_sg U13959 ( .A(n7012), .B(n2054), .X(n2053) );
  nor_x1_sg U13960 ( .A(n7305), .B(\update_mask_0/reg_out[11][15] ), .X(n2055)
         );
  nor_x1_sg U13961 ( .A(n2249), .B(n2250), .X(n2248) );
  nor_x1_sg U13962 ( .A(n2253), .B(n7405), .X(n2247) );
  nor_x1_sg U13963 ( .A(\update_mask_0/reg_i_mask[26] ), .B(n6381), .X(n2249)
         );
  nor_x1_sg U13964 ( .A(n1779), .B(n1780), .X(n1777) );
  nor_x1_sg U13965 ( .A(n6441), .B(\update_mask_0/reg_out[9][8] ), .X(n1778)
         );
  nor_x1_sg U13966 ( .A(n2117), .B(n2118), .X(n2115) );
  nor_x1_sg U13967 ( .A(n6168), .B(\update_mask_0/reg_out[9][18] ), .X(n2116)
         );
  nor_x1_sg U13968 ( .A(n1587), .B(n1588), .X(n1586) );
  nor_x1_sg U13969 ( .A(n1589), .B(n7014), .X(n1585) );
  nor_x1_sg U13970 ( .A(\update_mask_0/reg_out[14][1] ), .B(n6073), .X(n1587)
         );
  nor_x1_sg U13971 ( .A(n1596), .B(n1597), .X(n1590) );
  nor_x1_sg U13972 ( .A(n1592), .B(n8940), .X(n1591) );
  nor_x1_sg U13973 ( .A(\update_mask_0/reg_out[13][1] ), .B(n5999), .X(n1596)
         );
  nor_x1_sg U13974 ( .A(n1672), .B(n1673), .X(n1668) );
  nor_x1_sg U13975 ( .A(n1670), .B(n1671), .X(n1669) );
  nor_x1_sg U13976 ( .A(\update_mask_0/reg_out[3][4] ), .B(n6135), .X(n1672)
         );
  nor_x1_sg U13977 ( .A(n1679), .B(n1680), .X(n1674) );
  nor_x1_sg U13978 ( .A(\update_mask_0/reg_out[1][4] ), .B(n6003), .X(n1679)
         );
  nor_x1_sg U13979 ( .A(n1755), .B(n1756), .X(n1754) );
  nor_x1_sg U13980 ( .A(n1757), .B(n6119), .X(n1753) );
  nor_x1_sg U13981 ( .A(\update_mask_0/reg_out[14][6] ), .B(n7225), .X(n1755)
         );
  nor_x1_sg U13982 ( .A(n1764), .B(n1765), .X(n1758) );
  nor_x1_sg U13983 ( .A(n1760), .B(n8945), .X(n1759) );
  nor_x1_sg U13984 ( .A(\update_mask_0/reg_out[13][6] ), .B(n6164), .X(n1764)
         );
  nor_x1_sg U13985 ( .A(n1806), .B(n1807), .X(n1805) );
  nor_x1_sg U13986 ( .A(n1808), .B(n7012), .X(n1804) );
  nor_x1_sg U13987 ( .A(\update_mask_0/reg_out[14][9] ), .B(n6396), .X(n1806)
         );
  nor_x1_sg U13988 ( .A(n1815), .B(n1816), .X(n1809) );
  nor_x1_sg U13989 ( .A(n1811), .B(n8947), .X(n1810) );
  nor_x1_sg U13990 ( .A(\update_mask_0/reg_out[13][9] ), .B(n5999), .X(n1815)
         );
  nor_x1_sg U13991 ( .A(n1823), .B(n1824), .X(n1822) );
  nor_x1_sg U13992 ( .A(n1825), .B(n7013), .X(n1821) );
  nor_x1_sg U13993 ( .A(\update_mask_0/reg_out[14][7] ), .B(n6074), .X(n1823)
         );
  nor_x1_sg U13994 ( .A(n1832), .B(n1833), .X(n1826) );
  nor_x1_sg U13995 ( .A(n1828), .B(n8948), .X(n1827) );
  nor_x1_sg U13996 ( .A(\update_mask_0/reg_out[13][7] ), .B(n6444), .X(n1832)
         );
  nor_x1_sg U13997 ( .A(n1840), .B(n1841), .X(n1836) );
  nor_x1_sg U13998 ( .A(n1838), .B(n1839), .X(n1837) );
  nor_x1_sg U13999 ( .A(\update_mask_0/reg_out[3][9] ), .B(n7306), .X(n1840)
         );
  nor_x1_sg U14000 ( .A(n1925), .B(n1926), .X(n1924) );
  nor_x1_sg U14001 ( .A(n1927), .B(n7013), .X(n1923) );
  nor_x1_sg U14002 ( .A(\update_mask_0/reg_out[14][11] ), .B(n6073), .X(n1925)
         );
  nor_x1_sg U14003 ( .A(n1934), .B(n1935), .X(n1928) );
  nor_x1_sg U14004 ( .A(n1930), .B(n8950), .X(n1929) );
  nor_x1_sg U14005 ( .A(\update_mask_0/reg_out[13][11] ), .B(n7057), .X(n1934)
         );
  nor_x1_sg U14006 ( .A(n2010), .B(n2011), .X(n2006) );
  nor_x1_sg U14007 ( .A(n2008), .B(n2009), .X(n2007) );
  nor_x1_sg U14008 ( .A(\update_mask_0/reg_out[3][14] ), .B(n7304), .X(n2010)
         );
  nor_x1_sg U14009 ( .A(n2017), .B(n2018), .X(n2012) );
  nor_x1_sg U14010 ( .A(\update_mask_0/reg_out[1][14] ), .B(n6441), .X(n2017)
         );
  nor_x1_sg U14011 ( .A(n2093), .B(n2094), .X(n2092) );
  nor_x1_sg U14012 ( .A(n2095), .B(n6119), .X(n2091) );
  nor_x1_sg U14013 ( .A(\update_mask_0/reg_out[14][16] ), .B(n6234), .X(n2093)
         );
  nor_x1_sg U14014 ( .A(n2102), .B(n2103), .X(n2096) );
  nor_x1_sg U14015 ( .A(n2098), .B(n8955), .X(n2097) );
  nor_x1_sg U14016 ( .A(\update_mask_0/reg_out[13][16] ), .B(n7054), .X(n2102)
         );
  nor_x1_sg U14017 ( .A(n2144), .B(n2145), .X(n2143) );
  nor_x1_sg U14018 ( .A(n2146), .B(n6326), .X(n2142) );
  nor_x1_sg U14019 ( .A(\update_mask_0/reg_out[14][19] ), .B(n7226), .X(n2144)
         );
  nor_x1_sg U14020 ( .A(n2153), .B(n2154), .X(n2147) );
  nor_x1_sg U14021 ( .A(n2149), .B(n8957), .X(n2148) );
  nor_x1_sg U14022 ( .A(\update_mask_0/reg_out[13][19] ), .B(n7057), .X(n2153)
         );
  nor_x1_sg U14023 ( .A(n2161), .B(n2162), .X(n2160) );
  nor_x1_sg U14024 ( .A(n2163), .B(n6326), .X(n2159) );
  nor_x1_sg U14025 ( .A(\update_mask_0/reg_out[14][17] ), .B(n6073), .X(n2161)
         );
  nor_x1_sg U14026 ( .A(n2170), .B(n2171), .X(n2164) );
  nor_x1_sg U14027 ( .A(n2166), .B(n8958), .X(n2165) );
  nor_x1_sg U14028 ( .A(\update_mask_0/reg_out[13][17] ), .B(n6164), .X(n2170)
         );
  nor_x1_sg U14029 ( .A(n2178), .B(n2179), .X(n2174) );
  nor_x1_sg U14030 ( .A(n2176), .B(n2177), .X(n2175) );
  nor_x1_sg U14031 ( .A(\update_mask_0/reg_out[3][19] ), .B(n6482), .X(n2178)
         );
  nor_x1_sg U14032 ( .A(n2236), .B(n2237), .X(n2232) );
  nor_x1_sg U14033 ( .A(n2234), .B(n2235), .X(n2233) );
  nor_x1_sg U14034 ( .A(\update_mask_0/reg_i_mask[19] ), .B(n1459), .X(n2236)
         );
  nor_x1_sg U14035 ( .A(n2243), .B(n2244), .X(n2238) );
  nor_x1_sg U14036 ( .A(\update_mask_0/reg_i_mask[23] ), .B(n6541), .X(n2243)
         );
  nor_x1_sg U14037 ( .A(n1594), .B(n1595), .X(n1593) );
  nor_x1_sg U14038 ( .A(n6014), .B(\update_mask_0/reg_out[12][1] ), .X(n1594)
         );
  nor_x1_sg U14039 ( .A(n7098), .B(\update_mask_0/reg_out[8][1] ), .X(n1595)
         );
  nor_x1_sg U14040 ( .A(n1762), .B(n1763), .X(n1761) );
  nor_x1_sg U14041 ( .A(n6014), .B(\update_mask_0/reg_out[12][6] ), .X(n1762)
         );
  nor_x1_sg U14042 ( .A(n6434), .B(\update_mask_0/reg_out[8][6] ), .X(n1763)
         );
  nor_x1_sg U14043 ( .A(n1813), .B(n1814), .X(n1812) );
  nor_x1_sg U14044 ( .A(n7095), .B(\update_mask_0/reg_out[12][9] ), .X(n1813)
         );
  nor_x1_sg U14045 ( .A(n6179), .B(\update_mask_0/reg_out[8][9] ), .X(n1814)
         );
  nor_x1_sg U14046 ( .A(n1775), .B(n1776), .X(n1774) );
  nor_x1_sg U14047 ( .A(n6437), .B(\update_mask_0/reg_out[10][8] ), .X(n1775)
         );
  nor_x1_sg U14048 ( .A(n7055), .B(\update_mask_0/reg_out[13][8] ), .X(n1776)
         );
  nor_x1_sg U14049 ( .A(n1830), .B(n1831), .X(n1829) );
  nor_x1_sg U14050 ( .A(n7095), .B(\update_mask_0/reg_out[12][7] ), .X(n1830)
         );
  nor_x1_sg U14051 ( .A(n7100), .B(\update_mask_0/reg_out[8][7] ), .X(n1831)
         );
  nor_x1_sg U14052 ( .A(n1932), .B(n1933), .X(n1931) );
  nor_x1_sg U14053 ( .A(n6435), .B(\update_mask_0/reg_out[12][11] ), .X(n1932)
         );
  nor_x1_sg U14054 ( .A(n7101), .B(\update_mask_0/reg_out[8][11] ), .X(n1933)
         );
  nor_x1_sg U14055 ( .A(n2100), .B(n2101), .X(n2099) );
  nor_x1_sg U14056 ( .A(n7095), .B(\update_mask_0/reg_out[12][16] ), .X(n2100)
         );
  nor_x1_sg U14057 ( .A(n7100), .B(\update_mask_0/reg_out[8][16] ), .X(n2101)
         );
  nor_x1_sg U14058 ( .A(n2151), .B(n2152), .X(n2150) );
  nor_x1_sg U14059 ( .A(n7094), .B(\update_mask_0/reg_out[12][19] ), .X(n2151)
         );
  nor_x1_sg U14060 ( .A(n7100), .B(\update_mask_0/reg_out[8][19] ), .X(n2152)
         );
  nor_x1_sg U14061 ( .A(n2113), .B(n2114), .X(n2112) );
  nor_x1_sg U14062 ( .A(n7091), .B(\update_mask_0/reg_out[10][18] ), .X(n2113)
         );
  nor_x1_sg U14063 ( .A(n6000), .B(\update_mask_0/reg_out[13][18] ), .X(n2114)
         );
  nor_x1_sg U14064 ( .A(n2168), .B(n2169), .X(n2167) );
  nor_x1_sg U14065 ( .A(n7096), .B(\update_mask_0/reg_out[12][17] ), .X(n2168)
         );
  nor_x1_sg U14066 ( .A(n6433), .B(\update_mask_0/reg_out[8][17] ), .X(n2169)
         );
  nor_x1_sg U14067 ( .A(n6442), .B(\update_mask_0/reg_out[9][0] ), .X(n1542)
         );
  nor_x1_sg U14068 ( .A(n7060), .B(\update_mask_0/reg_out[9][3] ), .X(n1610)
         );
  nor_x1_sg U14069 ( .A(n6002), .B(\update_mask_0/reg_out[9][5] ), .X(n1710)
         );
  nor_x1_sg U14070 ( .A(n7061), .B(\update_mask_0/reg_out[9][10] ), .X(n1880)
         );
  nor_x1_sg U14071 ( .A(n6442), .B(\update_mask_0/reg_out[9][13] ), .X(n1948)
         );
  nor_x1_sg U14072 ( .A(n7060), .B(\update_mask_0/reg_out[9][15] ), .X(n2048)
         );
  nor_x1_sg U14073 ( .A(n7094), .B(\update_mask_0/reg_out[4][2] ), .X(n1523)
         );
  nor_x1_sg U14074 ( .A(n6436), .B(\update_mask_0/reg_out[4][3] ), .X(n1625)
         );
  nor_x1_sg U14075 ( .A(n7094), .B(\update_mask_0/reg_out[4][7] ), .X(n1695)
         );
  nor_x1_sg U14076 ( .A(n6176), .B(\update_mask_0/reg_out[4][8] ), .X(n1793)
         );
  nor_x1_sg U14077 ( .A(n6177), .B(\update_mask_0/reg_out[4][12] ), .X(n1865)
         );
  nor_x1_sg U14078 ( .A(n7093), .B(\update_mask_0/reg_out[4][13] ), .X(n1963)
         );
  nor_x1_sg U14079 ( .A(n6177), .B(\update_mask_0/reg_out[4][17] ), .X(n2033)
         );
  nor_x1_sg U14080 ( .A(n6013), .B(\update_mask_0/reg_out[4][18] ), .X(n2131)
         );
endmodule

