
module sparsity ( clk, reset, i_0, i_1, i_2, i_3, i_4, i_5, i_6, i_7, i_8, i_9, 
        i_10, i_11, i_12, i_13, i_14, i_15, w_0, w_1, w_2, w_3, w_4, w_5, w_6, 
        w_7, w_8, w_9, w_10, w_11, w_12, w_13, w_14, w_15, i_mask, w_mask, 
        input_ready, output_taken, oi_0, oi_1, oi_2, oi_3, oi_4, oi_5, oi_6, 
        oi_7, oi_8, oi_9, oi_10, oi_11, oi_12, oi_13, oi_14, oi_15, ow_0, ow_1, 
        ow_2, ow_3, ow_4, ow_5, ow_6, ow_7, ow_8, ow_9, ow_10, ow_11, ow_12, 
        ow_13, ow_14, ow_15, o_mask, state, input_taken );
  input [19:0] i_0;
  input [19:0] i_1;
  input [19:0] i_2;
  input [19:0] i_3;
  input [19:0] i_4;
  input [19:0] i_5;
  input [19:0] i_6;
  input [19:0] i_7;
  input [19:0] i_8;
  input [19:0] i_9;
  input [19:0] i_10;
  input [19:0] i_11;
  input [19:0] i_12;
  input [19:0] i_13;
  input [19:0] i_14;
  input [19:0] i_15;
  input [19:0] w_0;
  input [19:0] w_1;
  input [19:0] w_2;
  input [19:0] w_3;
  input [19:0] w_4;
  input [19:0] w_5;
  input [19:0] w_6;
  input [19:0] w_7;
  input [19:0] w_8;
  input [19:0] w_9;
  input [19:0] w_10;
  input [19:0] w_11;
  input [19:0] w_12;
  input [19:0] w_13;
  input [19:0] w_14;
  input [19:0] w_15;
  input [31:0] i_mask;
  input [31:0] w_mask;
  output [19:0] oi_0;
  output [19:0] oi_1;
  output [19:0] oi_2;
  output [19:0] oi_3;
  output [19:0] oi_4;
  output [19:0] oi_5;
  output [19:0] oi_6;
  output [19:0] oi_7;
  output [19:0] oi_8;
  output [19:0] oi_9;
  output [19:0] oi_10;
  output [19:0] oi_11;
  output [19:0] oi_12;
  output [19:0] oi_13;
  output [19:0] oi_14;
  output [19:0] oi_15;
  output [19:0] ow_0;
  output [19:0] ow_1;
  output [19:0] ow_2;
  output [19:0] ow_3;
  output [19:0] ow_4;
  output [19:0] ow_5;
  output [19:0] ow_6;
  output [19:0] ow_7;
  output [19:0] ow_8;
  output [19:0] ow_9;
  output [19:0] ow_10;
  output [19:0] ow_11;
  output [19:0] ow_12;
  output [19:0] ow_13;
  output [19:0] ow_14;
  output [19:0] ow_15;
  output [31:0] o_mask;
  output [1:0] state;
  input clk, reset, input_ready, output_taken;
  output input_taken;
  wire   n68592, n68593, n68594, n68595, n68596, n68597, n68598, n68599,
         n68600, n68601, n68602, n68603, n68604, n68605, n68606, n68607,
         n68608, n68609, n68610, n68611, n68612, n68613, n68614, n68615,
         n68616, n68617, n68618, n68619, n68620, n68621, n68622, n68623,
         n68624, n68625, n68626, n68627, n68628, n68629, n68630, n68631,
         n68632, n68633, n68634, n68635, n68636, n68637, n68638, n68639,
         n68640, n68641, n68642, n68643, n68644, n68645, n68646, n68647,
         n68648, n68649, n68650, n68651, n68652, n68653, n68654, n68655,
         n68656, n68657, n68658, n68659, n68660, n68661, n68662, n68663,
         n68664, n68665, n68666, n68667, n68668, n68669, n68670, n68671,
         n68672, n68673, n68674, n68675, n68676, n68677, n68678, n68679,
         n68680, n68681, n68682, n68683, n68684, n68685, n68686, n68687,
         n68688, n68689, n68690, n68691, n68692, n68693, n68694, n68695,
         n68696, n68697, n68698, n68699, n68700, n68701, n68702, n68703,
         n68704, n68705, n68706, n68707, n68708, n68709, n68710, n68711,
         n68712, n68713, n68714, n68715, n68716, n68717, n68718, n68719,
         n68720, n68721, n68722, n68723, n68724, n68725, n68726, n68727,
         n68728, n68729, n68730, n68731, n68732, n68733, n68734, n68735,
         n68736, n68737, n68738, n68739, n68740, n68741, n68742, n68743,
         n68744, n68745, n68746, n68747, n68748, n68749, n68750, n68751,
         n68752, n68753, n68754, n68755, n68756, n68757, n68758, n68759,
         n68760, n68761, n68762, n68763, n68764, n68765, n68766, n68767,
         n68768, n68769, n68770, n68771, n68772, n68773, n68774, n68775,
         n68776, n68777, n68778, n68779, n68780, n68781, n68782, n68783,
         n68784, n68785, n68786, n68787, n68788, n68789, n68790, n68791,
         n68792, n68793, n68794, n68795, n68796, n68797, n68798, n68799,
         n68800, n68801, n68802, n68803, n68804, n68805, n68806, n68807,
         n68808, n68809, n68810, n68811, n68812, n68813, n68814, n68815,
         n68816, n68817, n68818, n68819, n68820, n68821, n68822, n68823,
         n68824, n68825, n68826, n68827, n68828, n68829, n68830, n68831,
         n68832, n68833, n68834, n68835, n68836, n68837, n68838, n68839,
         n68840, n68841, n68842, n68843, n68844, n68845, n68846, n68847,
         n68848, n68849, n68850, n68851, n68852, n68853, n68854, n68855,
         n68856, n68857, n68858, n68859, n68860, n68861, n68862, n68863,
         n68864, n68865, n68866, n68867, n68868, n68869, n68870, n68871,
         n68872, n68873, n68874, n68875, n68876, n68877, n68878, n68879,
         n68880, n68881, n68882, n68883, n68884, n68885, n68886, n68887,
         n68888, n68889, n68890, n68891, n68892, n68893, n68894, n68895,
         n68896, n68897, n68898, n68899, n68900, n68901, n68902, n68903,
         n68904, n68905, n68906, n68907, n68908, n68909, n68910, n68911,
         n68912, n68913, n68914, n68915, n68916, n68917, n68918, n68919,
         n68920, n68921, n68922, n68923, n68924, n68925, n68926, n68927,
         n68928, n68929, n68930, n68931, n68932, n68933, n68934, n68935,
         n68936, n68937, n68938, n68939, n68940, n68941, n68942, n68943,
         n68944, n68945, n68946, n68947, n68948, n68949, n68950, n68951,
         n68952, n68953, n68954, n68955, n68956, n68957, n68958, n68959,
         n68960, n68961, n68962, n68963, n68964, n68965, n68966, n68967,
         n68968, n68969, n68970, n68971, n68972, n68973, n68974, n68975,
         n68976, n68977, n68978, n68979, n68980, n68981, n68982, n68983,
         n68984, n68985, n68986, n68987, n68988, n68989, n68990, n68991,
         n68992, n68993, n68994, n68995, n68996, n68997, n68998, n68999,
         n69000, n69001, n69002, n69003, n69004, n69005, n69006, n69007,
         n69008, n69009, n69010, n69011, n69012, n69013, n69014, n69015,
         n69016, n69017, n69018, n69019, n69020, n69021, n69022, n69023,
         n69024, n69025, n69026, n69027, n69028, n69029, n69030, n69031,
         n69032, n69033, n69034, n69035, n69036, n69037, n69038, n69039,
         n69040, n69041, n69042, n69043, n69044, n69045, n69046, n69047,
         n69048, n69049, n69050, n69051, n69052, n69053, n69054, n69055,
         n69056, n69057, n69058, n69059, n69060, n69061, n69062, n69063,
         n69064, n69065, n69066, n69067, n69068, n69069, n69070, n69071,
         n69072, n69073, n69074, n69075, n69076, n69077, n69078, n69079,
         n69080, n69081, n69082, n69083, n69084, n69085, n69086, n69087,
         n69088, n69089, n69090, n69091, n69092, n69093, n69094, n69095,
         n69096, n69097, n69098, n69099, n69100, n69101, n69102, n69103,
         n69104, n69105, n69106, n69107, n69108, n69109, n69110, n69111,
         n69112, n69113, n69114, n69115, n69116, n69117, n69118, n69119,
         n69120, n69121, n69122, n69123, n69124, n69125, n69126, n69127,
         n69128, n69129, n69130, n69131, n69132, n69133, n69134, n69135,
         n69136, n69137, n69138, n69139, n69140, n69141, n69142, n69143,
         n69144, n69145, n69146, n69147, n69148, n69149, n69150, n69151,
         n69152, n69153, n69154, n69155, n69156, n69157, n69158, n69159,
         n69160, n69161, n69162, n69163, n69164, n69165, n69166, n69167,
         n69168, n69169, n69170, n69171, n69172, n69173, n69174, n69175,
         n69176, n69177, n69178, n69179, n69180, n69181, n69182, n69183,
         n69184, n69185, n69186, n69187, n69188, n69189, n69190, n69191,
         n69192, n69193, n69194, n69195, n69196, n69197, n69198, n69199,
         n69200, n69201, n69202, n69203, n69204, n69205, n69206, n69207,
         n69208, n69209, n69210, n69211, n69212, n69213, n69214, n69215,
         n69216, n69217, n69218, n69219, n69220, n69221, n69222, n69223,
         n69224, n69225, n69226, n69227, n69228, n69229, n69230, n69231,
         n69232, n69233, n69234, n69235, n69236, n69237, n69238, n69239,
         n69240, n69241, n69242, n69243, n69244, n69245, n69246, n69247,
         n69248, n69249, n69250, n69251, n69252, n69253, n69254, n69255,
         n69256, n69257, n69258, n69259, n69260, n69261, n69262, n69263,
         mask_input_ready, delayed_input_ready, filter_input_ready, n10398,
         n10399, n10400, n10401, n10402, n10403, n10404, n10405, n10406,
         n10407, n10408, n10409, n10410, n10411, n10412, n10413, n10414,
         n10415, n10416, n10417, n10418, n10419, n10420, n10421, n10422,
         n10423, n10424, n10425, n10426, n10427, n10428, n10429, n10430,
         n10431, n10432, n10433, n10434, n10435, n10436, n10437, n10438,
         n10439, n10440, n10441, n10442, n10443, n10444, n10445, n10446,
         n10447, n10448, n10449, n10450, n10451, n10452, n10453, n10454,
         n10455, n10456, n10457, n10458, n10459, n10460, n10461, n10462,
         n69264, n69265, n69266, \mask_0/n1655 , \mask_0/n1654 ,
         \filter_0/n12237 , \filter_0/n11596 , \filter_0/n11595 ,
         \filter_0/n11594 , \filter_0/n11593 , \filter_0/n11592 ,
         \filter_0/n11591 , \filter_0/n11590 , \filter_0/n11589 ,
         \filter_0/n11588 , \filter_0/n11587 , \filter_0/n11586 ,
         \filter_0/n11585 , \filter_0/n11584 , \filter_0/n11583 ,
         \filter_0/n11582 , \filter_0/n11581 , \filter_0/n11580 ,
         \filter_0/n11579 , \filter_0/n11578 , \filter_0/n11577 ,
         \filter_0/n11576 , \filter_0/n11575 , \filter_0/n11574 ,
         \filter_0/n11573 , \filter_0/n11572 , \filter_0/n11571 ,
         \filter_0/n11570 , \filter_0/n11569 , \filter_0/n11568 ,
         \filter_0/n11567 , \filter_0/n11566 , \filter_0/n11565 ,
         \filter_0/n11564 , \filter_0/n11563 , \filter_0/n11562 ,
         \filter_0/n11561 , \filter_0/n11560 , \filter_0/n11559 ,
         \filter_0/n11558 , \filter_0/n11557 , \filter_0/n11556 ,
         \filter_0/n11555 , \filter_0/n11554 , \filter_0/n11553 ,
         \filter_0/n11552 , \filter_0/n11551 , \filter_0/n11550 ,
         \filter_0/n11549 , \filter_0/n11548 , \filter_0/n11547 ,
         \filter_0/n11546 , \filter_0/n11545 , \filter_0/n11544 ,
         \filter_0/n11543 , \filter_0/n11542 , \filter_0/n11541 ,
         \filter_0/n11540 , \filter_0/n11539 , \filter_0/n11538 ,
         \filter_0/n11537 , \filter_0/n11536 , \filter_0/n11535 ,
         \filter_0/n11534 , \filter_0/n11533 , \filter_0/n11532 ,
         \filter_0/n11531 , \filter_0/n11530 , \filter_0/n11529 ,
         \filter_0/n11528 , \filter_0/n11527 , \filter_0/n11526 ,
         \filter_0/n11525 , \filter_0/n11524 , \filter_0/n11523 ,
         \filter_0/n11522 , \filter_0/n11521 , \filter_0/n11520 ,
         \filter_0/n11519 , \filter_0/n11518 , \filter_0/n11517 ,
         \filter_0/n11516 , \filter_0/n11515 , \filter_0/n11514 ,
         \filter_0/n11513 , \filter_0/n11512 , \filter_0/n11511 ,
         \filter_0/n11510 , \filter_0/n11509 , \filter_0/n11508 ,
         \filter_0/n11507 , \filter_0/n11506 , \filter_0/n11505 ,
         \filter_0/n11504 , \filter_0/n11503 , \filter_0/n11502 ,
         \filter_0/n11501 , \filter_0/N1845 , \filter_0/done ,
         \filter_0/n17951 , \filter_0/n17950 , \filter_0/n17949 ,
         \filter_0/n17948 , \filter_0/n17947 , \filter_0/n17946 ,
         \filter_0/n17945 , \filter_0/n17944 , \filter_0/n17943 ,
         \filter_0/n17942 , \filter_0/n17941 , \filter_0/n17940 ,
         \filter_0/n17939 , \filter_0/n17938 , \filter_0/n17937 ,
         \filter_0/n17936 , \filter_0/n17935 , \filter_0/n17934 ,
         \filter_0/n17933 , \filter_0/n17932 , \filter_0/n17931 ,
         \filter_0/n17930 , \filter_0/n17929 , \filter_0/n17928 ,
         \filter_0/n17927 , \filter_0/n17926 , \filter_0/n17925 ,
         \filter_0/n17924 , \filter_0/n17923 , \filter_0/n17922 ,
         \filter_0/n17921 , \filter_0/n17920 , \filter_0/n17919 ,
         \filter_0/n17918 , \filter_0/n17917 , \filter_0/n17916 ,
         \filter_0/n17915 , \filter_0/n17914 , \filter_0/n17913 ,
         \filter_0/n17912 , \filter_0/n17911 , \filter_0/n17910 ,
         \filter_0/n17909 , \filter_0/n17908 , \filter_0/n17907 ,
         \filter_0/n17906 , \filter_0/n17905 , \filter_0/n17904 ,
         \filter_0/n17903 , \filter_0/n17902 , \filter_0/n17901 ,
         \filter_0/n17900 , \filter_0/n17899 , \filter_0/n17898 ,
         \filter_0/n17897 , \filter_0/n17896 , \filter_0/n17895 ,
         \filter_0/n17894 , \filter_0/n17893 , \filter_0/n17892 ,
         \filter_0/n17891 , \filter_0/n17890 , \filter_0/n17889 ,
         \filter_0/n17888 , \filter_0/n17887 , \filter_0/n17886 ,
         \filter_0/n17885 , \filter_0/n17884 , \filter_0/n17883 ,
         \filter_0/n17882 , \filter_0/n17881 , \filter_0/n17880 ,
         \filter_0/n17879 , \filter_0/n17878 , \filter_0/n17877 ,
         \filter_0/n17876 , \filter_0/n17875 , \filter_0/n17874 ,
         \filter_0/n17873 , \filter_0/n17872 , \filter_0/n17871 ,
         \filter_0/n17870 , \filter_0/n17869 , \filter_0/n17868 ,
         \filter_0/n17867 , \filter_0/n17866 , \filter_0/n17865 ,
         \filter_0/n17864 , \filter_0/n17863 , \filter_0/n17862 ,
         \filter_0/n17861 , \filter_0/n17860 , \filter_0/n17859 ,
         \filter_0/n17858 , \filter_0/n17857 , \filter_0/n17856 ,
         \filter_0/n17855 , \filter_0/n17854 , \filter_0/n17853 ,
         \filter_0/n17852 , \filter_0/n17851 , \filter_0/n17850 ,
         \filter_0/n17849 , \filter_0/n17848 , \filter_0/n17847 ,
         \filter_0/n17846 , \filter_0/n17845 , \filter_0/n17844 ,
         \filter_0/n17843 , \filter_0/n17842 , \filter_0/n17841 ,
         \filter_0/n17840 , \filter_0/n17839 , \filter_0/n17838 ,
         \filter_0/n17837 , \filter_0/n17836 , \filter_0/n17835 ,
         \filter_0/n17834 , \filter_0/n17833 , \filter_0/n17832 ,
         \filter_0/n17831 , \filter_0/n17830 , \filter_0/n17829 ,
         \filter_0/n17828 , \filter_0/n17827 , \filter_0/n17826 ,
         \filter_0/n17825 , \filter_0/n17824 , \filter_0/n17823 ,
         \filter_0/n17822 , \filter_0/n17821 , \filter_0/n17820 ,
         \filter_0/n17819 , \filter_0/n17818 , \filter_0/n17817 ,
         \filter_0/n17816 , \filter_0/n17815 , \filter_0/n17814 ,
         \filter_0/n17813 , \filter_0/n17812 , \filter_0/n17811 ,
         \filter_0/n17810 , \filter_0/n17809 , \filter_0/n17808 ,
         \filter_0/n17807 , \filter_0/n17806 , \filter_0/n17805 ,
         \filter_0/n17804 , \filter_0/n17803 , \filter_0/n17802 ,
         \filter_0/n17801 , \filter_0/n17800 , \filter_0/n17799 ,
         \filter_0/n17798 , \filter_0/n17797 , \filter_0/n17796 ,
         \filter_0/n17795 , \filter_0/n17794 , \filter_0/n17793 ,
         \filter_0/n17792 , \filter_0/n17791 , \filter_0/n17790 ,
         \filter_0/n17789 , \filter_0/n17788 , \filter_0/n17787 ,
         \filter_0/n17786 , \filter_0/n17785 , \filter_0/n17784 ,
         \filter_0/n17783 , \filter_0/n17782 , \filter_0/n17781 ,
         \filter_0/n17780 , \filter_0/n17779 , \filter_0/n17778 ,
         \filter_0/n17777 , \filter_0/n17776 , \filter_0/n17775 ,
         \filter_0/n17774 , \filter_0/n17773 , \filter_0/n17772 ,
         \filter_0/n17771 , \filter_0/n17770 , \filter_0/n17769 ,
         \filter_0/n17768 , \filter_0/n17767 , \filter_0/n17766 ,
         \filter_0/n17765 , \filter_0/n17764 , \filter_0/n17763 ,
         \filter_0/n17762 , \filter_0/n17761 , \filter_0/n17760 ,
         \filter_0/n17759 , \filter_0/n17758 , \filter_0/n17757 ,
         \filter_0/n17756 , \filter_0/n17755 , \filter_0/n17754 ,
         \filter_0/n17753 , \filter_0/n17752 , \filter_0/n17751 ,
         \filter_0/n17750 , \filter_0/n17749 , \filter_0/n17748 ,
         \filter_0/n17747 , \filter_0/n17746 , \filter_0/n17745 ,
         \filter_0/n17744 , \filter_0/n17743 , \filter_0/n17742 ,
         \filter_0/n17741 , \filter_0/n17740 , \filter_0/n17739 ,
         \filter_0/n17738 , \filter_0/n17737 , \filter_0/n17736 ,
         \filter_0/n17735 , \filter_0/n17734 , \filter_0/n17733 ,
         \filter_0/n17732 , \filter_0/n17731 , \filter_0/n17730 ,
         \filter_0/n17729 , \filter_0/n17728 , \filter_0/n17727 ,
         \filter_0/n17726 , \filter_0/n17725 , \filter_0/n17724 ,
         \filter_0/n17723 , \filter_0/n17722 , \filter_0/n17721 ,
         \filter_0/n17720 , \filter_0/n17719 , \filter_0/n17718 ,
         \filter_0/n17717 , \filter_0/n17716 , \filter_0/n17715 ,
         \filter_0/n17714 , \filter_0/n17713 , \filter_0/n17712 ,
         \filter_0/n17711 , \filter_0/n17710 , \filter_0/n17709 ,
         \filter_0/n17708 , \filter_0/n17707 , \filter_0/n17706 ,
         \filter_0/n17705 , \filter_0/n17704 , \filter_0/n17703 ,
         \filter_0/n17702 , \filter_0/n17701 , \filter_0/n17700 ,
         \filter_0/n17699 , \filter_0/n17698 , \filter_0/n17697 ,
         \filter_0/n17696 , \filter_0/n17695 , \filter_0/n17694 ,
         \filter_0/n17693 , \filter_0/n17692 , \filter_0/n17691 ,
         \filter_0/n17690 , \filter_0/n17689 , \filter_0/n17688 ,
         \filter_0/n17687 , \filter_0/n17686 , \filter_0/n17685 ,
         \filter_0/n17684 , \filter_0/n17683 , \filter_0/n17682 ,
         \filter_0/n17681 , \filter_0/n17680 , \filter_0/n17679 ,
         \filter_0/n17678 , \filter_0/n17677 , \filter_0/n17676 ,
         \filter_0/n17675 , \filter_0/n17674 , \filter_0/n17673 ,
         \filter_0/n17672 , \filter_0/n17671 , \filter_0/n17670 ,
         \filter_0/n17669 , \filter_0/n17668 , \filter_0/n17667 ,
         \filter_0/n17666 , \filter_0/n17665 , \filter_0/n17664 ,
         \filter_0/n17663 , \filter_0/n17662 , \filter_0/n17661 ,
         \filter_0/n17660 , \filter_0/n17659 , \filter_0/n17658 ,
         \filter_0/n17657 , \filter_0/n17656 , \filter_0/n17655 ,
         \filter_0/n17654 , \filter_0/n17653 , \filter_0/n17652 ,
         \filter_0/n17651 , \filter_0/n17650 , \filter_0/n17649 ,
         \filter_0/n17648 , \filter_0/n17647 , \filter_0/n17646 ,
         \filter_0/n17645 , \filter_0/n17644 , \filter_0/n17643 ,
         \filter_0/n17642 , \filter_0/n17641 , \filter_0/n17640 ,
         \filter_0/n17639 , \filter_0/n17638 , \filter_0/n17637 ,
         \filter_0/n17636 , \filter_0/n17635 , \filter_0/n17634 ,
         \filter_0/n17633 , \filter_0/n17632 , \filter_0/n17631 ,
         \filter_0/n17630 , \filter_0/n17629 , \filter_0/n17628 ,
         \filter_0/n17627 , \filter_0/n17626 , \filter_0/n17625 ,
         \filter_0/n17624 , \filter_0/n17623 , \filter_0/n17622 ,
         \filter_0/n17621 , \filter_0/n17620 , \filter_0/n17619 ,
         \filter_0/n17618 , \filter_0/n17617 , \filter_0/n17616 ,
         \filter_0/n17615 , \filter_0/n17614 , \filter_0/n17613 ,
         \filter_0/n17612 , \filter_0/n17611 , \filter_0/n17610 ,
         \filter_0/n17609 , \filter_0/n17608 , \filter_0/n17607 ,
         \filter_0/n17606 , \filter_0/n17605 , \filter_0/n17604 ,
         \filter_0/n17603 , \filter_0/n17602 , \filter_0/n17601 ,
         \filter_0/n17600 , \filter_0/n17599 , \filter_0/n17598 ,
         \filter_0/n17597 , \filter_0/n17596 , \filter_0/n17595 ,
         \filter_0/n17594 , \filter_0/n17593 , \filter_0/n17592 ,
         \filter_0/n17591 , \filter_0/n17590 , \filter_0/n17589 ,
         \filter_0/n17588 , \filter_0/n17587 , \filter_0/n17586 ,
         \filter_0/n17585 , \filter_0/n17584 , \filter_0/n17583 ,
         \filter_0/n17582 , \filter_0/n17581 , \filter_0/n17580 ,
         \filter_0/n17579 , \filter_0/n17578 , \filter_0/n17577 ,
         \filter_0/n17576 , \filter_0/n17575 , \filter_0/n17574 ,
         \filter_0/n17573 , \filter_0/n17572 , \filter_0/n17571 ,
         \filter_0/n17570 , \filter_0/n17569 , \filter_0/n17568 ,
         \filter_0/n17567 , \filter_0/n17566 , \filter_0/n17565 ,
         \filter_0/n17564 , \filter_0/n17563 , \filter_0/n17562 ,
         \filter_0/n17561 , \filter_0/n17560 , \filter_0/n17559 ,
         \filter_0/n17558 , \filter_0/n17557 , \filter_0/n17556 ,
         \filter_0/n17555 , \filter_0/n17554 , \filter_0/n17553 ,
         \filter_0/n17552 , \filter_0/n17551 , \filter_0/n17550 ,
         \filter_0/n17549 , \filter_0/n17548 , \filter_0/n17547 ,
         \filter_0/n17546 , \filter_0/n17545 , \filter_0/n17544 ,
         \filter_0/n17543 , \filter_0/n17542 , \filter_0/n17541 ,
         \filter_0/n17540 , \filter_0/n17539 , \filter_0/n17538 ,
         \filter_0/n17537 , \filter_0/n17536 , \filter_0/n17535 ,
         \filter_0/n17534 , \filter_0/n17533 , \filter_0/n17532 ,
         \filter_0/n17531 , \filter_0/n17530 , \filter_0/n17529 ,
         \filter_0/n17528 , \filter_0/n17527 , \filter_0/n17526 ,
         \filter_0/n17525 , \filter_0/n17524 , \filter_0/n17523 ,
         \filter_0/n17522 , \filter_0/n17521 , \filter_0/n17520 ,
         \filter_0/n17519 , \filter_0/n17518 , \filter_0/n17517 ,
         \filter_0/n17516 , \filter_0/n17515 , \filter_0/n17514 ,
         \filter_0/n17513 , \filter_0/n17512 , \filter_0/n17511 ,
         \filter_0/n17510 , \filter_0/n17509 , \filter_0/n17508 ,
         \filter_0/n17507 , \filter_0/n17506 , \filter_0/n17505 ,
         \filter_0/n17504 , \filter_0/n17503 , \filter_0/n17502 ,
         \filter_0/n17501 , \filter_0/n17500 , \filter_0/n17499 ,
         \filter_0/n17498 , \filter_0/n17497 , \filter_0/n17496 ,
         \filter_0/n17495 , \filter_0/n17494 , \filter_0/n17493 ,
         \filter_0/n17492 , \filter_0/n17491 , \filter_0/n17490 ,
         \filter_0/n17489 , \filter_0/n17488 , \filter_0/n17487 ,
         \filter_0/n17486 , \filter_0/n17485 , \filter_0/n17484 ,
         \filter_0/n17483 , \filter_0/n17482 , \filter_0/n17481 ,
         \filter_0/n17480 , \filter_0/n17479 , \filter_0/n17478 ,
         \filter_0/n17477 , \filter_0/n17476 , \filter_0/n17475 ,
         \filter_0/n17474 , \filter_0/n17473 , \filter_0/n17472 ,
         \filter_0/n17471 , \filter_0/n17470 , \filter_0/n17469 ,
         \filter_0/n17468 , \filter_0/n17467 , \filter_0/n17466 ,
         \filter_0/n17465 , \filter_0/n17464 , \filter_0/n17463 ,
         \filter_0/n17462 , \filter_0/n17461 , \filter_0/n17460 ,
         \filter_0/n17459 , \filter_0/n17458 , \filter_0/n17457 ,
         \filter_0/n17456 , \filter_0/n17455 , \filter_0/n17454 ,
         \filter_0/n17453 , \filter_0/n17452 , \filter_0/n17451 ,
         \filter_0/n17450 , \filter_0/n17449 , \filter_0/n17448 ,
         \filter_0/n17447 , \filter_0/n17446 , \filter_0/n17445 ,
         \filter_0/n17444 , \filter_0/n17443 , \filter_0/n17442 ,
         \filter_0/n17441 , \filter_0/n17440 , \filter_0/n17439 ,
         \filter_0/n17438 , \filter_0/n17437 , \filter_0/n17436 ,
         \filter_0/n17435 , \filter_0/n17434 , \filter_0/n17433 ,
         \filter_0/n17432 , \filter_0/n17431 , \filter_0/n17430 ,
         \filter_0/n17429 , \filter_0/n17428 , \filter_0/n17427 ,
         \filter_0/n17426 , \filter_0/n17425 , \filter_0/n17424 ,
         \filter_0/n17423 , \filter_0/n17422 , \filter_0/n17421 ,
         \filter_0/n17420 , \filter_0/n17419 , \filter_0/n17418 ,
         \filter_0/n17417 , \filter_0/n17416 , \filter_0/n17415 ,
         \filter_0/n17414 , \filter_0/n17413 , \filter_0/n17412 ,
         \filter_0/n17411 , \filter_0/n17410 , \filter_0/n17409 ,
         \filter_0/n17408 , \filter_0/n17407 , \filter_0/n17406 ,
         \filter_0/n17405 , \filter_0/n17404 , \filter_0/n17403 ,
         \filter_0/n17402 , \filter_0/n17401 , \filter_0/n17400 ,
         \filter_0/n17399 , \filter_0/n17398 , \filter_0/n17397 ,
         \filter_0/n17396 , \filter_0/n17395 , \filter_0/n17394 ,
         \filter_0/n17393 , \filter_0/n17392 , \filter_0/n17391 ,
         \filter_0/n17390 , \filter_0/n17389 , \filter_0/n17388 ,
         \filter_0/n17387 , \filter_0/n17386 , \filter_0/n17385 ,
         \filter_0/n17384 , \filter_0/n17383 , \filter_0/n17382 ,
         \filter_0/n17381 , \filter_0/n17380 , \filter_0/n17379 ,
         \filter_0/n17378 , \filter_0/n17377 , \filter_0/n17376 ,
         \filter_0/n17375 , \filter_0/n17374 , \filter_0/n17373 ,
         \filter_0/n17372 , \filter_0/n17371 , \filter_0/n17370 ,
         \filter_0/n17369 , \filter_0/n17368 , \filter_0/n17367 ,
         \filter_0/n17366 , \filter_0/n17365 , \filter_0/n17364 ,
         \filter_0/n17363 , \filter_0/n17362 , \filter_0/n17361 ,
         \filter_0/n17360 , \filter_0/n17359 , \filter_0/n17358 ,
         \filter_0/n17357 , \filter_0/n17356 , \filter_0/n17355 ,
         \filter_0/n17354 , \filter_0/n17353 , \filter_0/n17352 ,
         \filter_0/n17351 , \filter_0/n17350 , \filter_0/n17349 ,
         \filter_0/n17348 , \filter_0/n17347 , \filter_0/n17346 ,
         \filter_0/n17345 , \filter_0/n17344 , \filter_0/n17343 ,
         \filter_0/n17342 , \filter_0/n17341 , \filter_0/n17340 ,
         \filter_0/n17339 , \filter_0/n17338 , \filter_0/n17337 ,
         \filter_0/n17336 , \filter_0/n17335 , \filter_0/n17334 ,
         \filter_0/n17333 , \filter_0/n17332 , \filter_0/n17331 ,
         \filter_0/n17330 , \filter_0/n17329 , \filter_0/n17328 ,
         \filter_0/n17327 , \filter_0/n17326 , \filter_0/n17325 ,
         \filter_0/n17324 , \filter_0/n17323 , \filter_0/n17322 ,
         \filter_0/n17321 , \filter_0/n17320 , \filter_0/n17319 ,
         \filter_0/n17318 , \filter_0/n17317 , \filter_0/n17316 ,
         \filter_0/n17315 , \filter_0/n17314 , \filter_0/n17313 ,
         \filter_0/n17312 , \filter_0/n17311 , \filter_0/n17310 ,
         \filter_0/n17309 , \filter_0/N16 , \filter_0/N15 , \filter_0/N14 ,
         \filter_0/N13 , \filter_0/N12 , \shifter_0/n14056 ,
         \shifter_0/n27116 , \shifter_0/n27115 , \shifter_0/n27114 , n29326,
         n29327, n29328, n29329, n29332, n29333, n29336, n29337, n29338,
         n29339, n29344, n29345, n29346, n29347, n29348, n29349, n29350,
         n29351, n29352, n29353, n29354, n29355, n29356, n29357, n29358,
         n29359, n29360, n29361, n29362, n29363, n29364, n29365, n29366,
         n29367, n29368, n29369, n29370, n29371, n29372, n29373, n29374,
         n29375, n29376, n29377, n29378, n29379, n29380, n29381, n29382,
         n29383, n29384, n29385, n29386, n29387, n29388, n29389, n29390,
         n29391, n29392, n29393, n29394, n29395, n29396, n29397, n29398,
         n29399, n29400, n29401, n29402, n29403, n29404, n29405, n29406,
         n29407, n29408, n29409, n29410, n29411, n29412, n29413, n29414,
         n29415, n29416, n29417, n29418, n29419, n29420, n29421, n29422,
         n29423, n29424, n29425, n29426, n29427, n29428, n29429, n29430,
         n29431, n29432, n29433, n29434, n29435, n29436, n29437, n29438,
         n29439, n29440, n29441, n29442, n29443, n29444, n29445, n29446,
         n29447, n29448, n29449, n29450, n29451, n29452, n29453, n29454,
         n29455, n29456, n29457, n29458, n29459, n29460, n29461, n29462,
         n29463, n29464, n29465, n29466, n29467, n29468, n29469, n29470,
         n29471, n29472, n29473, n29474, n29475, n29476, n29477, n29478,
         n29479, n29480, n29481, n29482, n29483, n29484, n29485, n29486,
         n29487, n29488, n29489, n29490, n29491, n29492, n29493, n29494,
         n29495, n29496, n29497, n29498, n29499, n29500, n29501, n29502,
         n29503, n29504, n29505, n29506, n29507, n29508, n29509, n29510,
         n29511, n29512, n29513, n29514, n29515, n29516, n29517, n29518,
         n29519, n29520, n29521, n29522, n29523, n29524, n29525, n29526,
         n29527, n29528, n29529, n29530, n29531, n29532, n29533, n29534,
         n29535, n29536, n29537, n29538, n29539, n29540, n29541, n29542,
         n29543, n29544, n29545, n29546, n29547, n29548, n29549, n29550,
         n29551, n29552, n29553, n29554, n29555, n29556, n29557, n29558,
         n29559, n29560, n29561, n29562, n29563, n29564, n29565, n29566,
         n29567, n29568, n29569, n29570, n29571, n29572, n29573, n29574,
         n29575, n29576, n29577, n29578, n29579, n29580, n29581, n29582,
         n29583, n29584, n29585, n29586, n29587, n29588, n29589, n29590,
         n29591, n29592, n29593, n29594, n29595, n29596, n29597, n29598,
         n29599, n29600, n29601, n29602, n29603, n29604, n29605, n29606,
         n29607, n29608, n29609, n29610, n29611, n29612, n29613, n29614,
         n29615, n29616, n29617, n29618, n29619, n29620, n29621, n29622,
         n29623, n29624, n29625, n29626, n29627, n29628, n29629, n29630,
         n29631, n29632, n29633, n29634, n29635, n29636, n29637, n29638,
         n29639, n29640, n29641, n29642, n29643, n29644, n29645, n29646,
         n29647, n29648, n29649, n29650, n29651, n29652, n29653, n29654,
         n29655, n29656, n29657, n29658, n29659, n29660, n29661, n29662,
         n29663, n29664, n29665, n29666, n29667, n29668, n29669, n29670,
         n29671, n29672, n29673, n29674, n29675, n29676, n29677, n29678,
         n29679, n29680, n29681, n29682, n29683, n29684, n29685, n29686,
         n29687, n29688, n29689, n29690, n29691, n29692, n29693, n29694,
         n29695, n29696, n29697, n29698, n29699, n29700, n29701, n29702,
         n29703, n29704, n29705, n29706, n29707, n29708, n29709, n29710,
         n29711, n29712, n29713, n29714, n29715, n29716, n29717, n29718,
         n29719, n29720, n29721, n29722, n29723, n29724, n29725, n29726,
         n29727, n29728, n29729, n29730, n29731, n29732, n29733, n29734,
         n29735, n29736, n29737, n29738, n29739, n29740, n29741, n29742,
         n29743, n29744, n29745, n29746, n29747, n29748, n29749, n29750,
         n29751, n29752, n29753, n29754, n29755, n29756, n29757, n29758,
         n29759, n29760, n29761, n29762, n29763, n29764, n29765, n29766,
         n29767, n29768, n29769, n29770, n29771, n29772, n29773, n29774,
         n29775, n29776, n29777, n29778, n29779, n29780, n29781, n29782,
         n29783, n29784, n29785, n29786, n29787, n29788, n29789, n29790,
         n29791, n29792, n29793, n29794, n29795, n29796, n29797, n29798,
         n29799, n29800, n29801, n29802, n29803, n29804, n29805, n29806,
         n29807, n29808, n29809, n29810, n29811, n29812, n29813, n29814,
         n29815, n29816, n29817, n29818, n29819, n29820, n29821, n29822,
         n29823, n29824, n29825, n29826, n29827, n29828, n29829, n29830,
         n29831, n29832, n29833, n29834, n29835, n29836, n29837, n29838,
         n29839, n29840, n29841, n29842, n29843, n29844, n29845, n29846,
         n29847, n29848, n29849, n29850, n29851, n29852, n29853, n29854,
         n29855, n29856, n29857, n29858, n29859, n29860, n29861, n29862,
         n29863, n29864, n29865, n29866, n29867, n29868, n29869, n29870,
         n29871, n29872, n29873, n29874, n29875, n29876, n29877, n29878,
         n29879, n29880, n29881, n29882, n29883, n29884, n29885, n29886,
         n29887, n29888, n29889, n29890, n29891, n29892, n29893, n29894,
         n29895, n29896, n29897, n29898, n29899, n29900, n29901, n29902,
         n29903, n29904, n29905, n29906, n29907, n29908, n29909, n29910,
         n29911, n29912, n29913, n29914, n29915, n29916, n29917, n29918,
         n29919, n29920, n29921, n29922, n29923, n29924, n29925, n29926,
         n29927, n29928, n29929, n29930, n29931, n29932, n29933, n29934,
         n29935, n29936, n29937, n29938, n29939, n29940, n29941, n29942,
         n29943, n29944, n29945, n29946, n29947, n29948, n29949, n29950,
         n29951, n29952, n29953, n29954, n29955, n29956, n29957, n29958,
         n29959, n29960, n29961, n29962, n29963, n29964, n29965, n29966,
         n29967, n29968, n29969, n29970, n29971, n29972, n29973, n29974,
         n29975, n29976, n29977, n29978, n29979, n29980, n29981, n29982,
         n29983, n29984, n29985, n29986, n29987, n29988, n29989, n29990,
         n29991, n29992, n29993, n29994, n29995, n29996, n29997, n29998,
         n29999, n30000, n30001, n30002, n30003, n30004, n30005, n30006,
         n30007, n30008, n30009, n30010, n30011, n30012, n30013, n30014,
         n30015, n30016, n30017, n30018, n30019, n30020, n30021, n30022,
         n30023, n30024, n30025, n30026, n30027, n30028, n30029, n30030,
         n30031, n30032, n30033, n30034, n30035, n30036, n30037, n30038,
         n30039, n30040, n30041, n30042, n30043, n30044, n30045, n30046,
         n30047, n30048, n30049, n30050, n30051, n30052, n30053, n30054,
         n30055, n30056, n30057, n30058, n30059, n30060, n30061, n30062,
         n30063, n30064, n30065, n30066, n30067, n30068, n30069, n30070,
         n30071, n30072, n30073, n30074, n30075, n30076, n30077, n30078,
         n30079, n30080, n30081, n30082, n30083, n30084, n30085, n30086,
         n30087, n30088, n30089, n30090, n30091, n30092, n30093, n30094,
         n30095, n30096, n30097, n30098, n30099, n30100, n30101, n30102,
         n30103, n30104, n30105, n30106, n30107, n30108, n30109, n30110,
         n30111, n30112, n30113, n30114, n30115, n30116, n30117, n30118,
         n30119, n30120, n30121, n30122, n30123, n30124, n30125, n30126,
         n30127, n30128, n30129, n30130, n30131, n30132, n30133, n30134,
         n30135, n30136, n30137, n30138, n30139, n30140, n30141, n30142,
         n30143, n30144, n30145, n30146, n30147, n30148, n30149, n30150,
         n30151, n30152, n30153, n30154, n30155, n30156, n30157, n30158,
         n30159, n30160, n30161, n30162, n30163, n30164, n30165, n30166,
         n30167, n30168, n30169, n30170, n30171, n30172, n30173, n30174,
         n30175, n30176, n30177, n30178, n30179, n30180, n30181, n30182,
         n30183, n30184, n30185, n30186, n30187, n30188, n30189, n30190,
         n30191, n30192, n30193, n30194, n30195, n30196, n30197, n30198,
         n30199, n30200, n30201, n30202, n30203, n30204, n30205, n30206,
         n30207, n30208, n30209, n30210, n30211, n30212, n30213, n30214,
         n30215, n30216, n30217, n30218, n30219, n30220, n30221, n30222,
         n30223, n30224, n30225, n30226, n30227, n30228, n30229, n30230,
         n30231, n30232, n30233, n30234, n30235, n30236, n30237, n30238,
         n30239, n30240, n30241, n30242, n30243, n30244, n30245, n30246,
         n30247, n30248, n30249, n30250, n30251, n30252, n30253, n30254,
         n30255, n30256, n30257, n30258, n30259, n30260, n30261, n30262,
         n30263, n30264, n30265, n30266, n30267, n30268, n30269, n30270,
         n30271, n30272, n30273, n30274, n30275, n30276, n30277, n30278,
         n30279, n30280, n30281, n30282, n30283, n30284, n30285, n30286,
         n30287, n30288, n30289, n30290, n30291, n30292, n30293, n30294,
         n30295, n30296, n30297, n30298, n30299, n30300, n30301, n30302,
         n30303, n30304, n30305, n30306, n30307, n30308, n30309, n30310,
         n30311, n30312, n30313, n30314, n30315, n30316, n30317, n30318,
         n30319, n30320, n30321, n30322, n30323, n30324, n30325, n30326,
         n30327, n30328, n30329, n30330, n30331, n30332, n30333, n30334,
         n30335, n30336, n30337, n30338, n30339, n30340, n30341, n30342,
         n30343, n30344, n30345, n30346, n30347, n30348, n30349, n30350,
         n30351, n30352, n30353, n30354, n30355, n30356, n30357, n30358,
         n30359, n30360, n30361, n30362, n30363, n30364, n30365, n30366,
         n30367, n30368, n30369, n30370, n30371, n30372, n30373, n30374,
         n30375, n30376, n30377, n30378, n30379, n30380, n30381, n30382,
         n30383, n30384, n30385, n30386, n30387, n30388, n30389, n30390,
         n30391, n30392, n30393, n30394, n30395, n30396, n30397, n30398,
         n30399, n30400, n30401, n30402, n30403, n30404, n30405, n30406,
         n30407, n30408, n30409, n30410, n30411, n30412, n30413, n30414,
         n30415, n30416, n30417, n30418, n30419, n30420, n30421, n30422,
         n30423, n30424, n30425, n30426, n30427, n30428, n30429, n30430,
         n30431, n30432, n30433, n30434, n30435, n30436, n30437, n30438,
         n30439, n30440, n30441, n30442, n30443, n30444, n30445, n30446,
         n30447, n30448, n30449, n30450, n30451, n30452, n30453, n30454,
         n30455, n30456, n30457, n30458, n30459, n30460, n30461, n30462,
         n30463, n30464, n30465, n30466, n30467, n30468, n30469, n30470,
         n30471, n30472, n30473, n30474, n30475, n30476, n30477, n30478,
         n30479, n30480, n30481, n30482, n30483, n30484, n30485, n30486,
         n30487, n30488, n30489, n30490, n30491, n30492, n30493, n30494,
         n30495, n30496, n30497, n30498, n30499, n30500, n30501, n30502,
         n30503, n30504, n30505, n30506, n30507, n30508, n30509, n30510,
         n30511, n30512, n30513, n30514, n30515, n30516, n30517, n30518,
         n30519, n30520, n30521, n30522, n30523, n30524, n30525, n30526,
         n30527, n30528, n30529, n30530, n30531, n30532, n30533, n30534,
         n30535, n30536, n30537, n30538, n30539, n30540, n30541, n30542,
         n30543, n30544, n30545, n30546, n30547, n30548, n30549, n30550,
         n30551, n30552, n30553, n30554, n30555, n30556, n30557, n30558,
         n30559, n30560, n30561, n30562, n30563, n30564, n30565, n30566,
         n30567, n30568, n30569, n30570, n30571, n30572, n30573, n30574,
         n30575, n30576, n30577, n30578, n30579, n30580, n30581, n30582,
         n30583, n30584, n30585, n30586, n30587, n30588, n30589, n30590,
         n30591, n30592, n30593, n30594, n30595, n30596, n30597, n30598,
         n30599, n30600, n30601, n30602, n30603, n30604, n30605, n30606,
         n30607, n30608, n30609, n30610, n30611, n30612, n30613, n30614,
         n30615, n30616, n30617, n30618, n30619, n30620, n30621, n30622,
         n30623, n30624, n30625, n30626, n30627, n31921, n31922, n31923,
         n31924, n31925, n31926, n31927, n31928, n31931, n31932, n31933,
         n31934, n31935, n31936, n31937, n31938, n31939, n31940, n31941,
         n31942, n31943, n31944, n31945, n31946, n31947, n31948, n31949,
         n31950, n31951, n31952, n31953, n31954, n31955, n31957, n31958,
         n31959, n31960, n31961, n31962, n31963, n31964, n31966, n31967,
         n31968, n31969, n31970, n31971, n31972, n31973, n31974, n31975,
         n31976, n31977, n31978, n31979, n31980, n31981, n31982, n31983,
         n31984, n31985, n31986, n31987, n31988, n31989, n31990, n31991,
         n31992, n31993, n31994, n31995, n31996, n31997, n31998, n32001,
         n32002, n32003, n32004, n32005, n32006, n32007, n32008, n32009,
         n32010, n32011, n32012, n32013, n32014, n32015, n32016, n32017,
         n32018, n32019, n32020, n32021, n32022, n32023, n32024, n32025,
         n32026, n32027, n32028, n32029, n32030, n32031, n32032, n32033,
         n32034, n32035, n32036, n32037, n32038, n32039, n32041, n32042,
         n32043, n32044, n32045, n32046, n32047, n32048, n32049, n32050,
         n32051, n32052, n32053, n32054, n32056, n32057, n32058, n32059,
         n32060, n32061, n32062, n32063, n32064, n32065, n32066, n32067,
         n32068, n32072, n32073, n32074, n32075, n32076, n32077, n32078,
         n32079, n32080, n32081, n32082, n32083, n32084, n32085, n32086,
         n32087, n32088, n32089, n32090, n32091, n32092, n32093, n32094,
         n32095, n32098, n32099, n32100, n32101, n32102, n32103, n32104,
         n32105, n32106, n32107, n32108, n32109, n32110, n32111, n32112,
         n32113, n32114, n32115, n32116, n32117, n32118, n32119, n32120,
         n32121, n32122, n32123, n32124, n32125, n32126, n32127, n32128,
         n32129, n32130, n32131, n32132, n32133, n32134, n32135, n32136,
         n32137, n32138, n32139, n32140, n32141, n32142, n32143, n32144,
         n32145, n32146, n32147, n32148, n32149, n32150, n32151, n32152,
         n32153, n32154, n32155, n32156, n32157, n32158, n32159, n32160,
         n32161, n32162, n32163, n32164, n32165, n32166, n32167, n32168,
         n32169, n32170, n32171, n32172, n32175, n32176, n32177, n32178,
         n32179, n32180, n32181, n32182, n32183, n32184, n32185, n32186,
         n32187, n32188, n32189, n32190, n32191, n32192, n32193, n32194,
         n32195, n32196, n32197, n32198, n32199, n32200, n32201, n32202,
         n32203, n32204, n32205, n32206, n32207, n32208, n32209, n32210,
         n32211, n32212, n32222, n32223, n32224, n32225, n32226, n32227,
         n32228, n32229, n32230, n32231, n32232, n32233, n32234, n32235,
         n32236, n32237, n32238, n32239, n32240, n32241, n32242, n32243,
         n32244, n32245, n32246, n32247, n32248, n32249, n32250, n32251,
         n32252, n32253, n32254, n32255, n32256, n32257, n32258, n32259,
         n32260, n32261, n32262, n32263, n32264, n32265, n32266, n32267,
         n32268, n32269, n32270, n32271, n32272, n32273, n32274, n32275,
         n32276, n32277, n32278, n32279, n32280, n32281, n32282, n32283,
         n32284, n32285, n32286, n32287, n32288, n32289, n32290, n32291,
         n32292, n32293, n32294, n32295, n32296, n32297, n32298, n32299,
         n32300, n32301, n32302, n32303, n32304, n32305, n32306, n32307,
         n32308, n32309, n32310, n32311, n32312, n32313, n32314, n32315,
         n32316, n32317, n32318, n32319, n32320, n32321, n32322, n32323,
         n32324, n32325, n32326, n32327, n32328, n32329, n32330, n32331,
         n32332, n32333, n32334, n32335, n32336, n32337, n32338, n32339,
         n32340, n32341, n32342, n32343, n32344, n32345, n32346, n32347,
         n32348, n32349, n32350, n32351, n32352, n32353, n32354, n32366,
         n32367, n32368, n32369, n32370, n32371, n32372, n32373, n32374,
         n32375, n32376, n32377, n32378, n32379, n32380, n32381, n32382,
         n32383, n32384, n32385, n32386, n32387, n32388, n32389, n32390,
         n32391, n32392, n32393, n32394, n32395, n32396, n32399, n32400,
         n32401, n32402, n32403, n32404, n32405, n32406, n32407, n32408,
         n32409, n32410, n32411, n32412, n32413, n32414, n32415, n32416,
         n32417, n32418, n32419, n32420, n32421, n32422, n32423, n32424,
         n32425, n32426, n32427, n32428, n32429, n32430, n32431, n32433,
         n32434, n32435, n32436, n32437, n32438, n32439, n32440, n32443,
         n32444, n32445, n32446, n32447, n32448, n32449, n32450, n32451,
         n32452, n32453, n32454, n32455, n32456, n32457, n32458, n32459,
         n32460, n32461, n32462, n32463, n32464, n32465, n32466, n32467,
         n32468, n32469, n32470, n32471, n32472, n32473, n32474, n32475,
         n32476, n32477, n32478, n32479, n32480, n32481, n32482, n32483,
         n32484, n32485, n32486, n32487, n32488, n32489, n32490, n32491,
         n32492, n32493, n32494, n32495, n32496, n32497, n32499, n32500,
         n32504, n32505, n32506, n32507, n32508, n32509, n32510, n32511,
         n32512, n32513, n32514, n32517, n32518, n32519, n32520, n32521,
         n32522, n32523, n32524, n32525, n32526, n32527, n32528, n32529,
         n32530, n32531, n32532, n32533, n32534, n32535, n32536, n32537,
         n32538, n32539, n32540, n32543, n32544, n32545, n32546, n32547,
         n32548, n32549, n32550, n32551, n32552, n32553, n32554, n32555,
         n32556, n32557, n32558, n32559, n32560, n32561, n32562, n32563,
         n32564, n32565, n32566, n32567, n32568, n32569, n32570, n32571,
         n32572, n32573, n32574, n32575, n32576, n32577, n32578, n32579,
         n32580, n32581, n32582, n32583, n32584, n32585, n32586, n32587,
         n32588, n32589, n32590, n32591, n32592, n32593, n32594, n32595,
         n32596, n32597, n32598, n32599, n32600, n32601, n32602, n32603,
         n32604, n32605, n32606, n32607, n32608, n32609, n32610, n32611,
         n32612, n32613, n32614, n32615, n32616, n32617, n32620, n32621,
         n32622, n32623, n32624, n32625, n32626, n32627, n32628, n32629,
         n32630, n32631, n32632, n32633, n32634, n32635, n32636, n32637,
         n32638, n32639, n32640, n32641, n32642, n32643, n32644, n32645,
         n32646, n32647, n32648, n32649, n32650, n32651, n32652, n32653,
         n32654, n32655, n32656, n32657, n32667, n32668, n32669, n32670,
         n32671, n32672, n32673, n32674, n32675, n32676, n32677, n32678,
         n32679, n32680, n32681, n32682, n32683, n32684, n32685, n32686,
         n32687, n32688, n32689, n32690, n32691, n32692, n32693, n32694,
         n32695, n32696, n32697, n32698, n32699, n32700, n32701, n32702,
         n32703, n32704, n32705, n32706, n32707, n32708, n32709, n32710,
         n32711, n32712, n32713, n32714, n32715, n32716, n32717, n32718,
         n32719, n32720, n32721, n32722, n32723, n32724, n32725, n32726,
         n32727, n32728, n32729, n32730, n32731, n32732, n32733, n32734,
         n32735, n32736, n32737, n32738, n32739, n32740, n32741, n32742,
         n32743, n32744, n32745, n32746, n32747, n32748, n32749, n32750,
         n32751, n32752, n32753, n32754, n32755, n32756, n32757, n32758,
         n32759, n32760, n32761, n32762, n32763, n32764, n32765, n32766,
         n32767, n32768, n32769, n32770, n32771, n32772, n32773, n32774,
         n32775, n32776, n32777, n32778, n32779, n32780, n32781, n32782,
         n32783, n32784, n32785, n32786, n32787, n32788, n32789, n32790,
         n32791, n32792, n32793, n32794, n32795, n32796, n32797, n32798,
         n32799, n32800, n32801, n32802, n32803, n32804, n32805, n32806,
         n32807, n32808, n32809, n32810, n32811, n32812, n32813, n32814,
         n32815, n32816, n32817, n32818, n32819, n32820, n32821, n32822,
         n32823, n32824, n32825, n32826, n32827, n32828, n32829, n32830,
         n32831, n32832, n32833, n32834, n32835, n32836, n32837, n32838,
         n32839, n32840, n32841, n32842, n32843, n32844, n32845, n32846,
         n32847, n32848, n32849, n32850, n32851, n32852, n32853, n32854,
         n32855, n32856, n32857, n32858, n32859, n32860, n32861, n32862,
         n32863, n32864, n32865, n32866, n32867, n32868, n32869, n32870,
         n32871, n32872, n32873, n32874, n32875, n32876, n32877, n32878,
         n32879, n32880, n32881, n32882, n32883, n32884, n32885, n32886,
         n32887, n32888, n32889, n32890, n32891, n32892, n32893, n32894,
         n32895, n32896, n32897, n32898, n32899, n32900, n32901, n32902,
         n32903, n32904, n32905, n32906, n32907, n32908, n32909, n32910,
         n32911, n32912, n32913, n32914, n32915, n32916, n32917, n32918,
         n32919, n32920, n32921, n32922, n32923, n32924, n32925, n32926,
         n32927, n32928, n32929, n32930, n32931, n32932, n32933, n32934,
         n32935, n32936, n32937, n32938, n32939, n32940, n32941, n32942,
         n32943, n32944, n32945, n32946, n32947, n32948, n32949, n32950,
         n32951, n32952, n32953, n32954, n32955, n32956, n32957, n32958,
         n32959, n32960, n32961, n32962, n32963, n32964, n32965, n32966,
         n32967, n32968, n32969, n32970, n32971, n32972, n32973, n32974,
         n32975, n32976, n32977, n32978, n32979, n32980, n32981, n32982,
         n32983, n32984, n32985, n32986, n32987, n32988, n32989, n32990,
         n32991, n32992, n32993, n32994, n32995, n32996, n32997, n32998,
         n32999, n33000, n33001, n33002, n33003, n33004, n33005, n33006,
         n33007, n33008, n33009, n33010, n33011, n33012, n33013, n33014,
         n33015, n33016, n33017, n33018, n33019, n33020, n33021, n33022,
         n33023, n33024, n33025, n33026, n33027, n33028, n33029, n33030,
         n33031, n33032, n33033, n33034, n33035, n33036, n33037, n33038,
         n33039, n33040, n33041, n33042, n33043, n33044, n33045, n33046,
         n33047, n33048, n33049, n33050, n33051, n33052, n33053, n33054,
         n33055, n33056, n33057, n33058, n33059, n33060, n33061, n33062,
         n33063, n33064, n33065, n33066, n33067, n33068, n33069, n33070,
         n33071, n33072, n33073, n33074, n33075, n33076, n33077, n33078,
         n33079, n33080, n33081, n33082, n33083, n33084, n33085, n33086,
         n33087, n33088, n33089, n33090, n33091, n33092, n33093, n33094,
         n33095, n33096, n33097, n33098, n33099, n33100, n33101, n33102,
         n33103, n33104, n33105, n33106, n33107, n33108, n33109, n33110,
         n33111, n33112, n33113, n33114, n33115, n33116, n33117, n33118,
         n33119, n33120, n33121, n33122, n33123, n33124, n33125, n33126,
         n33127, n33128, n33129, n33130, n33131, n33132, n33133, n33134,
         n33135, n33136, n33137, n33138, n33139, n33140, n33141, n33142,
         n33143, n33144, n33145, n33146, n33147, n33148, n33149, n33150,
         n33151, n33152, n33153, n33154, n33155, n33156, n33157, n33158,
         n33159, n33160, n33161, n33162, n33163, n33164, n33165, n33166,
         n33167, n33168, n33169, n33170, n33171, n33172, n33173, n33174,
         n33175, n33176, n33177, n33178, n33179, n33180, n33181, n33182,
         n33183, n33184, n33185, n33186, n33187, n33188, n33189, n33190,
         n33191, n33192, n33193, n33194, n33195, n33196, n33197, n33198,
         n33199, n33200, n33201, n33202, n33203, n33204, n33205, n33206,
         n33207, n33208, n33209, n33210, n33211, n33212, n33213, n33214,
         n33215, n33216, n33217, n33218, n33219, n33220, n33221, n33222,
         n33223, n33224, n33225, n33226, n33227, n33228, n33229, n33230,
         n33231, n33232, n33233, n33234, n33235, n33236, n33237, n33238,
         n33239, n33240, n33241, n33242, n33243, n33244, n33245, n33246,
         n33247, n33248, n33249, n33250, n33251, n33252, n33253, n33254,
         n33255, n33256, n33257, n33258, n33259, n33260, n33261, n33262,
         n33263, n33264, n33265, n33266, n33267, n33268, n33269, n33270,
         n33271, n33272, n33273, n33274, n33275, n33276, n33277, n33278,
         n33279, n33280, n33281, n33282, n33283, n33284, n33285, n33286,
         n33287, n33288, n33289, n33290, n33291, n33292, n33293, n33294,
         n33295, n33296, n33297, n33298, n33299, n33300, n33301, n33302,
         n33303, n33304, n33305, n33306, n33307, n33308, n33309, n33310,
         n33311, n33312, n33313, n33314, n33315, n33316, n33317, n33318,
         n33319, n33320, n33321, n33322, n33323, n33324, n33325, n33326,
         n33327, n33328, n33329, n33330, n33331, n33332, n33333, n33334,
         n33335, n33336, n33337, n33338, n33339, n33340, n33341, n33342,
         n33343, n33344, n33345, n33346, n33347, n33348, n33349, n33350,
         n33351, n33352, n33353, n33354, n33355, n33356, n33357, n33358,
         n33359, n33360, n33361, n33362, n33363, n33364, n33365, n33366,
         n33367, n33368, n33369, n33370, n33371, n33372, n33373, n33374,
         n33375, n33376, n33377, n33378, n33379, n33380, n33381, n33382,
         n33383, n33384, n33385, n33386, n33387, n33388, n33389, n33390,
         n33391, n33392, n33393, n33394, n33395, n33396, n33397, n33398,
         n33399, n33400, n33401, n33402, n33403, n33404, n33405, n33406,
         n33407, n33408, n33409, n33410, n33411, n33412, n33413, n33414,
         n33415, n33416, n33417, n33418, n33419, n33420, n33421, n33422,
         n33423, n33424, n33425, n33426, n33427, n33428, n33429, n33430,
         n33431, n33432, n33433, n33434, n33435, n33436, n33437, n33438,
         n33439, n33440, n33441, n33442, n33443, n33444, n33445, n33446,
         n33447, n33448, n33449, n33450, n33451, n33452, n33453, n33454,
         n33455, n33456, n33457, n33458, n33459, n33460, n33461, n33462,
         n33463, n33464, n33465, n33466, n33467, n33468, n33469, n33470,
         n33471, n33472, n33473, n33474, n33475, n33476, n33477, n33478,
         n33479, n33480, n33481, n33482, n33483, n33484, n33485, n33486,
         n33487, n33488, n33489, n33490, n33491, n33492, n33493, n33494,
         n33495, n33496, n33497, n33498, n33499, n33500, n33501, n33502,
         n33503, n33504, n33505, n33506, n33507, n33508, n33509, n33510,
         n33511, n33512, n33513, n33514, n33515, n33516, n33517, n33518,
         n33519, n33520, n33521, n33522, n33523, n33524, n33525, n33526,
         n33527, n33528, n33529, n33530, n33531, n33532, n33533, n33534,
         n33535, n33536, n33537, n33538, n33539, n33540, n33541, n33542,
         n33543, n33544, n33545, n33546, n33547, n33548, n33549, n33550,
         n33551, n33552, n33553, n33554, n33555, n33556, n33557, n33558,
         n33559, n33560, n33561, n33562, n33563, n33564, n33565, n33566,
         n33567, n33568, n33569, n33570, n33571, n33572, n33573, n33574,
         n33575, n33576, n33577, n33578, n33579, n33580, n33581, n33582,
         n33583, n33584, n33585, n33586, n33587, n33588, n33589, n33590,
         n33591, n33592, n33593, n33594, n33595, n33596, n33597, n33598,
         n33599, n33600, n33601, n33602, n33603, n33604, n33605, n33606,
         n33607, n33608, n33609, n33610, n33611, n33612, n33613, n33614,
         n33615, n33616, n33617, n33618, n33619, n33620, n33621, n33622,
         n33623, n33624, n33625, n33626, n33627, n33628, n33629, n33630,
         n33631, n33632, n33633, n33634, n33635, n33636, n33637, n33638,
         n33639, n33640, n33641, n33642, n33643, n33644, n33645, n33646,
         n33647, n33648, n33649, n33650, n33651, n33652, n33653, n33654,
         n33655, n33656, n33657, n33658, n33659, n33660, n33661, n33662,
         n33663, n33664, n33665, n33666, n33667, n33668, n33669, n33670,
         n33671, n33672, n33673, n33674, n33675, n33676, n33677, n33678,
         n33679, n33680, n33681, n33682, n33683, n33684, n33685, n33686,
         n33687, n33688, n33689, n33690, n33691, n33692, n33693, n33694,
         n33695, n33696, n33697, n33698, n33699, n33700, n33701, n33702,
         n33703, n33704, n33705, n33706, n33707, n33708, n33709, n33710,
         n33711, n33712, n33713, n33714, n33715, n33716, n33717, n33718,
         n33719, n33720, n33721, n33722, n33723, n33724, n33725, n33726,
         n33727, n33728, n33729, n33730, n33731, n33732, n33733, n33734,
         n33735, n33736, n33737, n33738, n33739, n33740, n33741, n33742,
         n33743, n33744, n33745, n33746, n33747, n33748, n33749, n33750,
         n33751, n33752, n33753, n33754, n33755, n33756, n33757, n33758,
         n33759, n33760, n33761, n33762, n33763, n33764, n33765, n33766,
         n33767, n33768, n33769, n33770, n33771, n33772, n33773, n33774,
         n33775, n33776, n33777, n33778, n33779, n33780, n33781, n33782,
         n33783, n33784, n33785, n33786, n33787, n33788, n33789, n33790,
         n33791, n33792, n33793, n33794, n33795, n33796, n33797, n33798,
         n33799, n33800, n33801, n33802, n33803, n33804, n33805, n33806,
         n33807, n33808, n33809, n33810, n33811, n33812, n33813, n33814,
         n33815, n33816, n33817, n33818, n33819, n33820, n33821, n33822,
         n33823, n33824, n33825, n33826, n33827, n33828, n33829, n33830,
         n33831, n33832, n33833, n33834, n33835, n33836, n33837, n33838,
         n33839, n33840, n33841, n33842, n33843, n33844, n33845, n33846,
         n33847, n33848, n33849, n33850, n33851, n33852, n33853, n33854,
         n33855, n33856, n33857, n33858, n33859, n33860, n33861, n33862,
         n33863, n33864, n33865, n33866, n33867, n33868, n33869, n33870,
         n33871, n33872, n33873, n33874, n33875, n33876, n33877, n33878,
         n33879, n33880, n33881, n33882, n33883, n33884, n33885, n33886,
         n33887, n33888, n33889, n33890, n33891, n33892, n33893, n33894,
         n33895, n33896, n33897, n33898, n33899, n33900, n33901, n33902,
         n33903, n33904, n33905, n33906, n33907, n33908, n33909, n33910,
         n33911, n33912, n33913, n33914, n33915, n33916, n33917, n33918,
         n33919, n33920, n33921, n33922, n33923, n33924, n33925, n33926,
         n33927, n33928, n33929, n33930, n33931, n33932, n33933, n33934,
         n33935, n33936, n33937, n33938, n33939, n33940, n33941, n33942,
         n33943, n33944, n33945, n33946, n33947, n33948, n33949, n33950,
         n33951, n33952, n33953, n33954, n33955, n33956, n33957, n33958,
         n33959, n33960, n33961, n33962, n33963, n33964, n33965, n33966,
         n33967, n33968, n33969, n33970, n33971, n33972, n33973, n33974,
         n33975, n33976, n33977, n33978, n33979, n33980, n33981, n33982,
         n33983, n33984, n33985, n33986, n33987, n33988, n33989, n33990,
         n33991, n33992, n33993, n33994, n33995, n33996, n33997, n33998,
         n33999, n34000, n34001, n34002, n34003, n34004, n34005, n34006,
         n34007, n34008, n34009, n34010, n34011, n34012, n34013, n34014,
         n34015, n34016, n34017, n34018, n34019, n34020, n34021, n34022,
         n34023, n34024, n34025, n34026, n34027, n34028, n34029, n34030,
         n34031, n34032, n34033, n34034, n34035, n34036, n34037, n34038,
         n34039, n34040, n34041, n34042, n34043, n34044, n34045, n34046,
         n34047, n34048, n34049, n34050, n34051, n34052, n34053, n34054,
         n34055, n34056, n34057, n34058, n34059, n34060, n34061, n34062,
         n34063, n34064, n34065, n34066, n34067, n34068, n34069, n34070,
         n34071, n34072, n34073, n34074, n34075, n34076, n34077, n34078,
         n34079, n34080, n34081, n34082, n34083, n34084, n34085, n34086,
         n34087, n34088, n34089, n34090, n34091, n34092, n34093, n34094,
         n34095, n34096, n34097, n34098, n34099, n34100, n34101, n34102,
         n34103, n34104, n34105, n34106, n34107, n34108, n34109, n34110,
         n34111, n34112, n34113, n34114, n34115, n34116, n34117, n34118,
         n34119, n34120, n34121, n34122, n34123, n34124, n34125, n34126,
         n34127, n34128, n34129, n34130, n34131, n34132, n34133, n34134,
         n34135, n34136, n34137, n34138, n34139, n34140, n34141, n34142,
         n34143, n34144, n34145, n34146, n34147, n34148, n34149, n34150,
         n34151, n34152, n34153, n34154, n34155, n34156, n34157, n34158,
         n34159, n34160, n34161, n34162, n34163, n34164, n34165, n34166,
         n34167, n34168, n34169, n34170, n34171, n34172, n34173, n34174,
         n34175, n34176, n34177, n34178, n34179, n34180, n34181, n34182,
         n34183, n34184, n34185, n34186, n34187, n34188, n34189, n34190,
         n34191, n34192, n34193, n34194, n34195, n34196, n34197, n34198,
         n34199, n34200, n34201, n34202, n34203, n34204, n34205, n34206,
         n34207, n34208, n34209, n34210, n34211, n34212, n34213, n34214,
         n34215, n34216, n34217, n34218, n34219, n34220, n34221, n34222,
         n34223, n34224, n34225, n34226, n34227, n34228, n34229, n34230,
         n34231, n34232, n34233, n34234, n34235, n34236, n34237, n34238,
         n34239, n34240, n34241, n34242, n34243, n34244, n34245, n34246,
         n34247, n34248, n34249, n34250, n34251, n34252, n34253, n34254,
         n34255, n34256, n34257, n34258, n34259, n34260, n34261, n34262,
         n34263, n34264, n34265, n34266, n34267, n34268, n34269, n34270,
         n34271, n34272, n34273, n34274, n34275, n34276, n34277, n34278,
         n34279, n34280, n34281, n34282, n34283, n34284, n34285, n34286,
         n34287, n34288, n34289, n34290, n34291, n34292, n34293, n34294,
         n34295, n34296, n34297, n34298, n34299, n34300, n34301, n34302,
         n34303, n34304, n34305, n34306, n34307, n34308, n34309, n34310,
         n34311, n34312, n34313, n34314, n34315, n34316, n34317, n34318,
         n34319, n34320, n34321, n34322, n34323, n34324, n34325, n34326,
         n34327, n34328, n34329, n34330, n34331, n34332, n34333, n34334,
         n34335, n34336, n34337, n34338, n34339, n34340, n34341, n34342,
         n34343, n34344, n34345, n34346, n34347, n34348, n34349, n34350,
         n34351, n34352, n34353, n34354, n34355, n34356, n34357, n34358,
         n34359, n34360, n34361, n34362, n34363, n34364, n34365, n34366,
         n34367, n34368, n34369, n34370, n34371, n34372, n34373, n34374,
         n34375, n34376, n34377, n34378, n34379, n34380, n34381, n34382,
         n34383, n34384, n34385, n34386, n34387, n34388, n34389, n34390,
         n34391, n34392, n34393, n34394, n34395, n34396, n34397, n34398,
         n34399, n34400, n34401, n34402, n34403, n34404, n34405, n34406,
         n34407, n34408, n34409, n34410, n34411, n34412, n34413, n34414,
         n34415, n34416, n34417, n34418, n34419, n34420, n34421, n34422,
         n34423, n34424, n34425, n34426, n34427, n34428, n34429, n34430,
         n34431, n34432, n34433, n34434, n34435, n34436, n34437, n34438,
         n34439, n34440, n34441, n34442, n34443, n34444, n34445, n34446,
         n34447, n34448, n34449, n34450, n34451, n34452, n34453, n34454,
         n34455, n34456, n34457, n34458, n34459, n34460, n34461, n34462,
         n34463, n34464, n34465, n34466, n34467, n34468, n34469, n34470,
         n34471, n34472, n34473, n34474, n34475, n34476, n34477, n34478,
         n34479, n34480, n34481, n34482, n34483, n34484, n34485, n34486,
         n34487, n34488, n34489, n34490, n34491, n34492, n34493, n34494,
         n34495, n34496, n34497, n34498, n34499, n34500, n34501, n34502,
         n34503, n34504, n34505, n34506, n34507, n34508, n34509, n34510,
         n34511, n34512, n34513, n34514, n34515, n34516, n34517, n34518,
         n34519, n34520, n34521, n34522, n34523, n34524, n34525, n34526,
         n34527, n34528, n34529, n34530, n34531, n34532, n34533, n34534,
         n34535, n34536, n34537, n34538, n34539, n34540, n34541, n34542,
         n34543, n34544, n34545, n34546, n34547, n34548, n34549, n34550,
         n34551, n34552, n34553, n34554, n34555, n34556, n34557, n34558,
         n34559, n34560, n34561, n34562, n34563, n34564, n34565, n34566,
         n34567, n34568, n34569, n34570, n34571, n34572, n34573, n34574,
         n34575, n34576, n34577, n34578, n34579, n34580, n34581, n34582,
         n34583, n34584, n34585, n34586, n34587, n34588, n34589, n34590,
         n34591, n34592, n34593, n34594, n34595, n34596, n34597, n34598,
         n34599, n34600, n34601, n34602, n34603, n34604, n34605, n34606,
         n34607, n34608, n34609, n34610, n34611, n34612, n34613, n34614,
         n34615, n34616, n34617, n34618, n34619, n34620, n34621, n34622,
         n34623, n34624, n34625, n34626, n34627, n34628, n34629, n34630,
         n34631, n34632, n34633, n34634, n34635, n34636, n34637, n34638,
         n34639, n34640, n34641, n34642, n34643, n34644, n34645, n34646,
         n34647, n34648, n34649, n34650, n34651, n34652, n34653, n34654,
         n34655, n34656, n34657, n34658, n34659, n34660, n34661, n34662,
         n34663, n34664, n34665, n34666, n34667, n34668, n34669, n34670,
         n34671, n34672, n34673, n34674, n34675, n34676, n34677, n34678,
         n34679, n34680, n34681, n34682, n34683, n34684, n34685, n34686,
         n34687, n34688, n34689, n34690, n34691, n34692, n34693, n34694,
         n34695, n34696, n34697, n34698, n34699, n34700, n34701, n34702,
         n34703, n34704, n34705, n34706, n34707, n34708, n34709, n34710,
         n34711, n34712, n34713, n34714, n34715, n34716, n34717, n34718,
         n34719, n34720, n34721, n34722, n34723, n34724, n34725, n34726,
         n34727, n34728, n34729, n34730, n34731, n34732, n34733, n34734,
         n34735, n34736, n34737, n34738, n34739, n34740, n34741, n34742,
         n34743, n34744, n34745, n34746, n34747, n34748, n34749, n34750,
         n34751, n34752, n34753, n34754, n34755, n34756, n34757, n34758,
         n34759, n34760, n34761, n34762, n34763, n34764, n34765, n34766,
         n34767, n34768, n34769, n34770, n34771, n34772, n34773, n34774,
         n34775, n34776, n34777, n34778, n34779, n34780, n34781, n34782,
         n34783, n34784, n34785, n34786, n34787, n34788, n34789, n34790,
         n34791, n34792, n34793, n34794, n34795, n34796, n34797, n34798,
         n34799, n34800, n34801, n34802, n34803, n34804, n34805, n34806,
         n34807, n34808, n34809, n34810, n34811, n34812, n34813, n34814,
         n34815, n34816, n34817, n34818, n34819, n34820, n34821, n34822,
         n34823, n34824, n34825, n34826, n34827, n34828, n34829, n34830,
         n34831, n34832, n34833, n34834, n34835, n34836, n34837, n34838,
         n34839, n34840, n34841, n34842, n34843, n34844, n34845, n34846,
         n34847, n34848, n34849, n34850, n34851, n34852, n34853, n34854,
         n34855, n34856, n34857, n34858, n34859, n34860, n34861, n34862,
         n34863, n34864, n34865, n34866, n34867, n34868, n34869, n34870,
         n34871, n34872, n34873, n34874, n34875, n34876, n34877, n34878,
         n34879, n34880, n34881, n34882, n34883, n34884, n34885, n34886,
         n34887, n34888, n34889, n34890, n34891, n34892, n34893, n34894,
         n34895, n34896, n34897, n34898, n34899, n34900, n34901, n34902,
         n34903, n34904, n34905, n34906, n34907, n34908, n34909, n34910,
         n34911, n34912, n34913, n34914, n34915, n34916, n34917, n34918,
         n34919, n34920, n34921, n34922, n34923, n34924, n34925, n34926,
         n34927, n34928, n34929, n34930, n34931, n34932, n34933, n34934,
         n34935, n34936, n34937, n34938, n34939, n34940, n34941, n34942,
         n34943, n34944, n34945, n34946, n34947, n34948, n34949, n34950,
         n34951, n34952, n34953, n34954, n34955, n34956, n34957, n34958,
         n34959, n34960, n34961, n34962, n34963, n34964, n34965, n34966,
         n34967, n34968, n34969, n34970, n34971, n34972, n34973, n34974,
         n34975, n34976, n34977, n34978, n34979, n34980, n34981, n34982,
         n34983, n34984, n34985, n34986, n34987, n34988, n34989, n34990,
         n34991, n34992, n34993, n34994, n34995, n34996, n34997, n34998,
         n34999, n35000, n35001, n35002, n35003, n35004, n35005, n35006,
         n35007, n35008, n35009, n35010, n35011, n35012, n35013, n35014,
         n35015, n35016, n35017, n35018, n35019, n35020, n35021, n35022,
         n35023, n35024, n35025, n35026, n35027, n35028, n35029, n35030,
         n35031, n35032, n35033, n35034, n35035, n35036, n35037, n35038,
         n35039, n35040, n35041, n35042, n35043, n35044, n35045, n35046,
         n35047, n35048, n35049, n35050, n35051, n35052, n35053, n35054,
         n35055, n35056, n35057, n35058, n35059, n35060, n35061, n35062,
         n35063, n35064, n35065, n35066, n35067, n35068, n35069, n35070,
         n35071, n35072, n35073, n35074, n35075, n35076, n35077, n35078,
         n35079, n35080, n35081, n35082, n35083, n35084, n35085, n35086,
         n35087, n35088, n35089, n35090, n35091, n35092, n35093, n35094,
         n35095, n35096, n35097, n35098, n35099, n35100, n35101, n35102,
         n35103, n35104, n35105, n35106, n35107, n35108, n35109, n35110,
         n35111, n35112, n35113, n35114, n35115, n35116, n35117, n35118,
         n35119, n35120, n35121, n35122, n35123, n35124, n35125, n35126,
         n35127, n35128, n35129, n35130, n35131, n35132, n35133, n35134,
         n35135, n35136, n35137, n35138, n35139, n35140, n35141, n35142,
         n35143, n35144, n35145, n35146, n35147, n35148, n35149, n35150,
         n35151, n35152, n35153, n35154, n35155, n35156, n35157, n35158,
         n35159, n35160, n35161, n35162, n35163, n35164, n35165, n35166,
         n35167, n35168, n35169, n35170, n35171, n35172, n35173, n35174,
         n35175, n35176, n35177, n35178, n35179, n35180, n35181, n35182,
         n35183, n35184, n35185, n35186, n35187, n35188, n35189, n35190,
         n35191, n35192, n35193, n35194, n35195, n35196, n35197, n35198,
         n35199, n35200, n35201, n35202, n35203, n35204, n35205, n35206,
         n35207, n35208, n35209, n35210, n35211, n35212, n35213, n35214,
         n35215, n35216, n35217, n35218, n35219, n35220, n35221, n35222,
         n35223, n35224, n35225, n35226, n35227, n35228, n35229, n35230,
         n35231, n35232, n35233, n35234, n35235, n35236, n35237, n35238,
         n35239, n35240, n35241, n35242, n35243, n35244, n35245, n35246,
         n35247, n35248, n35249, n35250, n35251, n35252, n35253, n35254,
         n35255, n35256, n35257, n35258, n35259, n35260, n35261, n35262,
         n35263, n35264, n35265, n35266, n35267, n35268, n35269, n35270,
         n35271, n35272, n35273, n35274, n35275, n35276, n35277, n35278,
         n35279, n35280, n35281, n35282, n35283, n35284, n35285, n35286,
         n35287, n35288, n35289, n35290, n35291, n35292, n35293, n35294,
         n35295, n35296, n35297, n35298, n35299, n35300, n35301, n35302,
         n35303, n35304, n35305, n35306, n35307, n35308, n35309, n35310,
         n35311, n35312, n35313, n35314, n35315, n35316, n35317, n35318,
         n35319, n35320, n35321, n35322, n35323, n35324, n35325, n35326,
         n35327, n35328, n35329, n35330, n35331, n35332, n35333, n35334,
         n35335, n35336, n35337, n35338, n35339, n35340, n35341, n35342,
         n35343, n35344, n35345, n35346, n35347, n35348, n35349, n35350,
         n35351, n35352, n35353, n35354, n35355, n35356, n35357, n35358,
         n35359, n35360, n35361, n35362, n35363, n35364, n35365, n35366,
         n35367, n35368, n35369, n35370, n35371, n35372, n35373, n35374,
         n35375, n35376, n35377, n35378, n35379, n35380, n35381, n35382,
         n35383, n35384, n35385, n35386, n35387, n35388, n35389, n35390,
         n35391, n35392, n35393, n35394, n35395, n35396, n35397, n35398,
         n35399, n35400, n35401, n35402, n35403, n35404, n35405, n35406,
         n35407, n35408, n35409, n35410, n35411, n35412, n35413, n35414,
         n35415, n35416, n35417, n35418, n35419, n35420, n35421, n35422,
         n35423, n35424, n35425, n35426, n35427, n35428, n35429, n35430,
         n35431, n35432, n35433, n35434, n35435, n35436, n35437, n35438,
         n35439, n35440, n35441, n35442, n35443, n35444, n35445, n35446,
         n35447, n35448, n35449, n35450, n35451, n35452, n35453, n35454,
         n35455, n35456, n35457, n35458, n35459, n35460, n35461, n35462,
         n35463, n35464, n35465, n35466, n35467, n35468, n35469, n35470,
         n35471, n35472, n35473, n35474, n35475, n35476, n35477, n35478,
         n35479, n35480, n35481, n35482, n35483, n35484, n35485, n35486,
         n35487, n35488, n35489, n35490, n35491, n35492, n35493, n35494,
         n35495, n35496, n35497, n35498, n35499, n35500, n35501, n35502,
         n35503, n35504, n35505, n35506, n35507, n35508, n35509, n35510,
         n35511, n35512, n35513, n35514, n35515, n35516, n35517, n35518,
         n35519, n35520, n35521, n35522, n35523, n35524, n35525, n35526,
         n35527, n35528, n35529, n35530, n35531, n35532, n35533, n35534,
         n35535, n35536, n35537, n35538, n35539, n35540, n35541, n35542,
         n35543, n35544, n35545, n35546, n35547, n35548, n35549, n35550,
         n35551, n35552, n35553, n35554, n35555, n35556, n35557, n35558,
         n35559, n35560, n35561, n35562, n35563, n35564, n35565, n35566,
         n35567, n35568, n35569, n35570, n35571, n35572, n35573, n35574,
         n35575, n35576, n35577, n35578, n35579, n35580, n35581, n35582,
         n35583, n35584, n35585, n35586, n35587, n35588, n35589, n35590,
         n35591, n35592, n35593, n35594, n35595, n35596, n35597, n35598,
         n35599, n35600, n35601, n35602, n35603, n35604, n35605, n35606,
         n35607, n35608, n35609, n35610, n35611, n35612, n35613, n35614,
         n35615, n35616, n35617, n35618, n35619, n35620, n35621, n35622,
         n35623, n35624, n35625, n35626, n35627, n35628, n35629, n35630,
         n35631, n35632, n35633, n35634, n35635, n35636, n35637, n35638,
         n35639, n35640, n35641, n35642, n35643, n35644, n35645, n35646,
         n35647, n35648, n35649, n35650, n35651, n35652, n35653, n35654,
         n35655, n35656, n35657, n35658, n35659, n35660, n35661, n35662,
         n35663, n35664, n35665, n35666, n35667, n35668, n35669, n35670,
         n35671, n35672, n35673, n35674, n35675, n35676, n35677, n35678,
         n35679, n35680, n35681, n35682, n35683, n35684, n35685, n35686,
         n35687, n35688, n35689, n35690, n35691, n35692, n35693, n35694,
         n35695, n35696, n35697, n35698, n35699, n35700, n35701, n35702,
         n35703, n35704, n35705, n35706, n35707, n35708, n35709, n35710,
         n35711, n35712, n35713, n35714, n35715, n35716, n35717, n35718,
         n35719, n35720, n35721, n35722, n35723, n35724, n35725, n35726,
         n35727, n35728, n35729, n35730, n35731, n35732, n35733, n35734,
         n35735, n35736, n35737, n35738, n35739, n35740, n35741, n35742,
         n35743, n35744, n35745, n35746, n35747, n35748, n35749, n35750,
         n35751, n35752, n35753, n35754, n35755, n35756, n35757, n35758,
         n35759, n35760, n35761, n35762, n35763, n35764, n35765, n35766,
         n35767, n35768, n35769, n35770, n35771, n35772, n35773, n35774,
         n35775, n35776, n35777, n35778, n35779, n35780, n35781, n35782,
         n35783, n35784, n35785, n35786, n35787, n35788, n35789, n35790,
         n35791, n35792, n35793, n35794, n35795, n35796, n35797, n35798,
         n35799, n35800, n35801, n35802, n35803, n35804, n35805, n35806,
         n35807, n35808, n35809, n35810, n35811, n35812, n35813, n35814,
         n35815, n35816, n35817, n35818, n35819, n35820, n35821, n35822,
         n35823, n35824, n35825, n35826, n35827, n35828, n35829, n35830,
         n35831, n35832, n35833, n35834, n35835, n35836, n35837, n35838,
         n35839, n35840, n35841, n35842, n35843, n35844, n35845, n35846,
         n35847, n35848, n35849, n35850, n35851, n35852, n35853, n35854,
         n35855, n35856, n35857, n35858, n35859, n35860, n35861, n35862,
         n35863, n35864, n35865, n35866, n35867, n35868, n35869, n35870,
         n35871, n35872, n35873, n35874, n35875, n35876, n35877, n35878,
         n35879, n35880, n35881, n35882, n35883, n35884, n35885, n35886,
         n35887, n35888, n35889, n35890, n35891, n35892, n35893, n35894,
         n35895, n35896, n35897, n35898, n35899, n35900, n35901, n35902,
         n35903, n35904, n35905, n35906, n35907, n35908, n35909, n35910,
         n35911, n35912, n35913, n35914, n35915, n35916, n35917, n35918,
         n35919, n35920, n35921, n35922, n35923, n35924, n35925, n35926,
         n35927, n35928, n35929, n35930, n35931, n35932, n35933, n35934,
         n35935, n35936, n35937, n35938, n35939, n35940, n35941, n35942,
         n35943, n35944, n35945, n35946, n35947, n35948, n35949, n35950,
         n35951, n35952, n35953, n35954, n35955, n35956, n35957, n35958,
         n35959, n35960, n35961, n35962, n35963, n35964, n35965, n35966,
         n35967, n35968, n35969, n35970, n35971, n35972, n35973, n35974,
         n35975, n35976, n35977, n35978, n35979, n35980, n35981, n35982,
         n35983, n35984, n35985, n35986, n35987, n35988, n35989, n35990,
         n35991, n35992, n35993, n35994, n35995, n35996, n35997, n35998,
         n35999, n36000, n36001, n36002, n36003, n36004, n36005, n36006,
         n36007, n36008, n36009, n36010, n36011, n36012, n36013, n36014,
         n36015, n36016, n36017, n36018, n36019, n36020, n36021, n36022,
         n36023, n36024, n36025, n36026, n36027, n36028, n36029, n36030,
         n36031, n36032, n36033, n36034, n36035, n36036, n36037, n36038,
         n36039, n36040, n36041, n36042, n36043, n36044, n36045, n36046,
         n36047, n36048, n36049, n36050, n36051, n36052, n36053, n36054,
         n36055, n36056, n36057, n36058, n36059, n36060, n36061, n36062,
         n36063, n36064, n36065, n36066, n36067, n36068, n36069, n36070,
         n36071, n36072, n36073, n36074, n36075, n36076, n36077, n36078,
         n36079, n36080, n36081, n36082, n36083, n36084, n36085, n36086,
         n36087, n36088, n36089, n36090, n36091, n36092, n36093, n36094,
         n36095, n36096, n36097, n36098, n36099, n36100, n36101, n36102,
         n36103, n36104, n36105, n36106, n36107, n36108, n36109, n36110,
         n36111, n36112, n36113, n36114, n36115, n36116, n36117, n36118,
         n36119, n36120, n36121, n36122, n36123, n36124, n36125, n36126,
         n36127, n36128, n36129, n36130, n36131, n36132, n36133, n36134,
         n36135, n36136, n36137, n36138, n36139, n36140, n36141, n36142,
         n36143, n36144, n36145, n36146, n36147, n36148, n36149, n36150,
         n36151, n36152, n36153, n36154, n36155, n36156, n36157, n36158,
         n36159, n36160, n36161, n36162, n36163, n36164, n36165, n36166,
         n36167, n36168, n36169, n36170, n36171, n36172, n36173, n36174,
         n36175, n36176, n36177, n36178, n36179, n36180, n36181, n36182,
         n36183, n36184, n36185, n36186, n36187, n36188, n36189, n36190,
         n36191, n36192, n36193, n36194, n36195, n36196, n36197, n36198,
         n36199, n36200, n36201, n36202, n36203, n36204, n36205, n36206,
         n36207, n36208, n36209, n36210, n36211, n36212, n36213, n36214,
         n36215, n36216, n36217, n36218, n36219, n36220, n36221, n36222,
         n36223, n36224, n36225, n36226, n36227, n36228, n36229, n36230,
         n36231, n36232, n36233, n36234, n36235, n36236, n36237, n36238,
         n36239, n36240, n36241, n36242, n36243, n36244, n36245, n36246,
         n36247, n36248, n36249, n36250, n36251, n36252, n36253, n36254,
         n36255, n36256, n36257, n36258, n36259, n36260, n36261, n36262,
         n36263, n36264, n36265, n36266, n36267, n36268, n36269, n36270,
         n36271, n36272, n36273, n36274, n36275, n36276, n36277, n36278,
         n36279, n36280, n36281, n36282, n36283, n36284, n36285, n36286,
         n36287, n36288, n36289, n36290, n36291, n36292, n36293, n36294,
         n36295, n36296, n36297, n36298, n36299, n36300, n36301, n36302,
         n36303, n36304, n36305, n36306, n36307, n36308, n36309, n36310,
         n36311, n36312, n36313, n36314, n36315, n36316, n36317, n36318,
         n36319, n36320, n36321, n36322, n36323, n36324, n36325, n36326,
         n36327, n36328, n36329, n36330, n36331, n36332, n36333, n36334,
         n36335, n36336, n36337, n36338, n36339, n36340, n36341, n36342,
         n36343, n36344, n36345, n36346, n36347, n36348, n36349, n36350,
         n36351, n36352, n36353, n36354, n36355, n36356, n36357, n36358,
         n36359, n36360, n36361, n36362, n36363, n36364, n36365, n36366,
         n36367, n36368, n36369, n36370, n36371, n36372, n36373, n36374,
         n36375, n36376, n36377, n36378, n36379, n36380, n36381, n36382,
         n36383, n36384, n36385, n36386, n36387, n36388, n36389, n36390,
         n36391, n36392, n36393, n36394, n36395, n36396, n36397, n36398,
         n36399, n36400, n36401, n36402, n36403, n36404, n36405, n36406,
         n36407, n36408, n36409, n36410, n36411, n36412, n36413, n36414,
         n36415, n36416, n36417, n36418, n36419, n36420, n36421, n36422,
         n36423, n36424, n36425, n36426, n36427, n36428, n36429, n36430,
         n36431, n36432, n36433, n36434, n36435, n36436, n36437, n36438,
         n36439, n36440, n36441, n36442, n36443, n36444, n36445, n36446,
         n36447, n36448, n36449, n36450, n36451, n36452, n36453, n36454,
         n36455, n36456, n36457, n36458, n36459, n36460, n36461, n36462,
         n36463, n36464, n36465, n36466, n36467, n36468, n36469, n36470,
         n36471, n36472, n36473, n36474, n36475, n36476, n36477, n36478,
         n36479, n36480, n36481, n36482, n36483, n36484, n36485, n36486,
         n36487, n36488, n36489, n36490, n36491, n36492, n36493, n36494,
         n36495, n36496, n36497, n36498, n36499, n36500, n36501, n36502,
         n36503, n36504, n36505, n36506, n36507, n36508, n36509, n36510,
         n36511, n36512, n36513, n36514, n36515, n36516, n36517, n36518,
         n36519, n36520, n36521, n36522, n36523, n36524, n36525, n36526,
         n36527, n36528, n36529, n36530, n36531, n36532, n36533, n36534,
         n36535, n36536, n36537, n36538, n36539, n36540, n36541, n36542,
         n36543, n36544, n36545, n36546, n36547, n36548, n36549, n36550,
         n36551, n36552, n36553, n36554, n36555, n36556, n36557, n36558,
         n36559, n36560, n36561, n36562, n36563, n36564, n36565, n36566,
         n36567, n36568, n36569, n36570, n36571, n36572, n36573, n36574,
         n36575, n36576, n36577, n36578, n36579, n36580, n36581, n36582,
         n36583, n36584, n36585, n36586, n36587, n36588, n36589, n36590,
         n36591, n36592, n36593, n36594, n36595, n36596, n36597, n36598,
         n36599, n36600, n36601, n36602, n36603, n36604, n36605, n36606,
         n36607, n36608, n36609, n36610, n36611, n36612, n36613, n36614,
         n36615, n36616, n36617, n36618, n36619, n36620, n36621, n36622,
         n36623, n36624, n36625, n36626, n36627, n36628, n36629, n36630,
         n36631, n36632, n36633, n36634, n36635, n36636, n36637, n36638,
         n36639, n36640, n36641, n36642, n36643, n36644, n36645, n36646,
         n36647, n36648, n36649, n36650, n36651, n36652, n36653, n36654,
         n36655, n36656, n36657, n36658, n36659, n36660, n36661, n36662,
         n36663, n36664, n36665, n36666, n36667, n36668, n36669, n36670,
         n36671, n36672, n36673, n36674, n36675, n36676, n36677, n36678,
         n36679, n36680, n36681, n36682, n36683, n36684, n36685, n36686,
         n36687, n36688, n36689, n36690, n36691, n36692, n36693, n36694,
         n36695, n36696, n36697, n36698, n36699, n36700, n36701, n36702,
         n36703, n36704, n36705, n36706, n36707, n36708, n36709, n36710,
         n36711, n36712, n36713, n36714, n36715, n36716, n36717, n36718,
         n36719, n36720, n36721, n36722, n36723, n36724, n36725, n36726,
         n36727, n36728, n36729, n36730, n36731, n36732, n36733, n36734,
         n36735, n36736, n36737, n36738, n36739, n36740, n36741, n36742,
         n36743, n36744, n36745, n36746, n36747, n36748, n36749, n36750,
         n36751, n36752, n36753, n36754, n36755, n36756, n36757, n36758,
         n36759, n36760, n36761, n36762, n36763, n36764, n36765, n36766,
         n36767, n36768, n36769, n36770, n36771, n36772, n36773, n36774,
         n36775, n36776, n36777, n36778, n36779, n36780, n36781, n36782,
         n36783, n36784, n36785, n36786, n36787, n36788, n36789, n36790,
         n36791, n36792, n36793, n36794, n36795, n36796, n36797, n36798,
         n36799, n36800, n36801, n36802, n36803, n36804, n36805, n36806,
         n36807, n36808, n36809, n36810, n36811, n36812, n36813, n36814,
         n36815, n36816, n36817, n36818, n36819, n36820, n36821, n36822,
         n36823, n36824, n36825, n36826, n36827, n36828, n36829, n36830,
         n36831, n36832, n36833, n36834, n36835, n36836, n36837, n36838,
         n36839, n36840, n36841, n36842, n36843, n36844, n36845, n36846,
         n36847, n36848, n36849, n36850, n36851, n36852, n36853, n36854,
         n36855, n36856, n36857, n36858, n36859, n36860, n36861, n36862,
         n36863, n36864, n36865, n36866, n36867, n36868, n36869, n36870,
         n36871, n36872, n36873, n36874, n36875, n36876, n36877, n36878,
         n36879, n36880, n36881, n36882, n36883, n36884, n36885, n36886,
         n36887, n36888, n36889, n36890, n36891, n36892, n36893, n36894,
         n36895, n36896, n36897, n36898, n36899, n36900, n36901, n36902,
         n36903, n36904, n36905, n36906, n36907, n36908, n36909, n36910,
         n36911, n36912, n36913, n36914, n36915, n36916, n36917, n36918,
         n36919, n36920, n36921, n36922, n36923, n36924, n36925, n36926,
         n36927, n36928, n36929, n36930, n36931, n36932, n36933, n36934,
         n36935, n36936, n36937, n36938, n36939, n36940, n36941, n36942,
         n36943, n36944, n36945, n36946, n36947, n36948, n36949, n36950,
         n36951, n36952, n36953, n36954, n36955, n36956, n36957, n36958,
         n36959, n36960, n36961, n36962, n36963, n36964, n36965, n36966,
         n36967, n36968, n36969, n36970, n36971, n36972, n36973, n36974,
         n36975, n36976, n36977, n36978, n36979, n36980, n36981, n36982,
         n36983, n36984, n36985, n36986, n36987, n36988, n36989, n36990,
         n36991, n36992, n36993, n36994, n36995, n36996, n36997, n36998,
         n36999, n37000, n37001, n37002, n37003, n37004, n37005, n37006,
         n37007, n37008, n37009, n37010, n37011, n37012, n37013, n37014,
         n37015, n37016, n37017, n37018, n37019, n37020, n37021, n37022,
         n37023, n37024, n37025, n37026, n37027, n37028, n37029, n37030,
         n37031, n37032, n37033, n37034, n37035, n37036, n37037, n37038,
         n37039, n37040, n37041, n37042, n37043, n37044, n37045, n37046,
         n37047, n37048, n37049, n37050, n37051, n37052, n37053, n37054,
         n37055, n37056, n37057, n37058, n37059, n37060, n37061, n37062,
         n37063, n37064, n37065, n37066, n37067, n37068, n37069, n37070,
         n37071, n37072, n37073, n37074, n37075, n37076, n37077, n37078,
         n37079, n37080, n37081, n37082, n37083, n37084, n37085, n37086,
         n37087, n37088, n37089, n37090, n37091, n37092, n37093, n37094,
         n37095, n37096, n37097, n37098, n37099, n37100, n37101, n37102,
         n37103, n37104, n37105, n37106, n37107, n37108, n37109, n37110,
         n37111, n37112, n37113, n37114, n37115, n37116, n37117, n37118,
         n37119, n37120, n37121, n37122, n37123, n37124, n37125, n37126,
         n37127, n37128, n37129, n37130, n37131, n37132, n37133, n37134,
         n37135, n37136, n37137, n37138, n37139, n37140, n37141, n37142,
         n37143, n37144, n37145, n37146, n37147, n37148, n37149, n37150,
         n37151, n37152, n37153, n37154, n37155, n37156, n37157, n37158,
         n37159, n37160, n37161, n37162, n37163, n37164, n37165, n37166,
         n37167, n37168, n37169, n37170, n37171, n37172, n37173, n37174,
         n37175, n37176, n37177, n37178, n37179, n37180, n37181, n37182,
         n37183, n37184, n37185, n37186, n37187, n37188, n37189, n37190,
         n37191, n37192, n37193, n37194, n37195, n37196, n37197, n37198,
         n37199, n37200, n37201, n37202, n37203, n37204, n37205, n37206,
         n37207, n37208, n37209, n37210, n37211, n37212, n37213, n37214,
         n37215, n37216, n37217, n37218, n37219, n37220, n37221, n37222,
         n37223, n37224, n37225, n37226, n37227, n37228, n37229, n37230,
         n37231, n37232, n37233, n37234, n37235, n37236, n37237, n37238,
         n37239, n37240, n37241, n37242, n37243, n37244, n37245, n37246,
         n37247, n37248, n37249, n37250, n37251, n37252, n37253, n37254,
         n37255, n37256, n37257, n37258, n37259, n37260, n37261, n37262,
         n37263, n37264, n37265, n37266, n37267, n37268, n37269, n37270,
         n37271, n37272, n37273, n37274, n37275, n37276, n37277, n37278,
         n37279, n37280, n37281, n37282, n37283, n37284, n37285, n37286,
         n37287, n37288, n37289, n37290, n37291, n37292, n37293, n37294,
         n37295, n37296, n37297, n37298, n37299, n37300, n37301, n37302,
         n37303, n37304, n37305, n37306, n37307, n37308, n37309, n37310,
         n37311, n37312, n37313, n37314, n37315, n37316, n37317, n37318,
         n37319, n37320, n37321, n37322, n37323, n37324, n37325, n37326,
         n37327, n37328, n37329, n37330, n37331, n37332, n37333, n37334,
         n37335, n37336, n37337, n37338, n37339, n37340, n37341, n37342,
         n37343, n37344, n37345, n37346, n37347, n37348, n37349, n37350,
         n37351, n37352, n37353, n37354, n37355, n37356, n37357, n37358,
         n37359, n37360, n37361, n37362, n37363, n37364, n37365, n37366,
         n37367, n37368, n37369, n37370, n37371, n37372, n37373, n37374,
         n37375, n37376, n37377, n37378, n37379, n37380, n37381, n37382,
         n37383, n37384, n37385, n37386, n37387, n37388, n37389, n37390,
         n37391, n37392, n37393, n37394, n37395, n37396, n37397, n37398,
         n37399, n37400, n37401, n37402, n37403, n37404, n37405, n37406,
         n37407, n37408, n37409, n37410, n37411, n37412, n37413, n37414,
         n37415, n37416, n37417, n37418, n37419, n37420, n37421, n37422,
         n37423, n37424, n37425, n37426, n37427, n37428, n37429, n37430,
         n37431, n37432, n37433, n37434, n37435, n37436, n37437, n37438,
         n37439, n37440, n37441, n37442, n37443, n37444, n37445, n37446,
         n37447, n37448, n37449, n37450, n37451, n37452, n37453, n37454,
         n37455, n37456, n37457, n37458, n37459, n37460, n37461, n37462,
         n37463, n37464, n37465, n37466, n37467, n37468, n37469, n37470,
         n37471, n37472, n37473, n37474, n37475, n37476, n37477, n37478,
         n37479, n37480, n37481, n37482, n37483, n37484, n37485, n37486,
         n37487, n37488, n37489, n37490, n37491, n37492, n37493, n37494,
         n37495, n37496, n37497, n37498, n37499, n37500, n37501, n37502,
         n37503, n37504, n37505, n37506, n37507, n37508, n37509, n37510,
         n37511, n37512, n37513, n37514, n37515, n37516, n37517, n37518,
         n37519, n37520, n37521, n37522, n37523, n37524, n37525, n37526,
         n37527, n37528, n37529, n37530, n37531, n37532, n37533, n37534,
         n37535, n37536, n37537, n37538, n37539, n37540, n37541, n37542,
         n37543, n37544, n37545, n37546, n37547, n37548, n37549, n37550,
         n37551, n37552, n37553, n37554, n37555, n37556, n37557, n37558,
         n37559, n37560, n37561, n37562, n37563, n37564, n37565, n37566,
         n37567, n37568, n37569, n37570, n37571, n37572, n37573, n37574,
         n37575, n37576, n37577, n37578, n37579, n37580, n37581, n37582,
         n37583, n37584, n37585, n37586, n37587, n37588, n37589, n37590,
         n37591, n37592, n37593, n37594, n37595, n37596, n37597, n37598,
         n37599, n37600, n37601, n37602, n37603, n37604, n37605, n37606,
         n37607, n37608, n37609, n37610, n37611, n37612, n37613, n37614,
         n37615, n37616, n37617, n37618, n37619, n37620, n37621, n37622,
         n37623, n37624, n37625, n37626, n37627, n37628, n37629, n37630,
         n37631, n37632, n37633, n37634, n37635, n37636, n37637, n37638,
         n37639, n37640, n37641, n37642, n37643, n37644, n37645, n37646,
         n37647, n37648, n37649, n37650, n37651, n37652, n37653, n37654,
         n37655, n37656, n37657, n37658, n37659, n37660, n37661, n37662,
         n37663, n37664, n37665, n37666, n37667, n37668, n37669, n37670,
         n37671, n37672, n37673, n37674, n37675, n37676, n37677, n37678,
         n37679, n37680, n37681, n37682, n37683, n37684, n37685, n37686,
         n37687, n37688, n37689, n37690, n37691, n37692, n37693, n37694,
         n37695, n37696, n37697, n37698, n37699, n37700, n37701, n37702,
         n37703, n37704, n37705, n37706, n37707, n37708, n37709, n37710,
         n37711, n37712, n37713, n37714, n37715, n37716, n37717, n37718,
         n37719, n37720, n37721, n37722, n37723, n37724, n37725, n37726,
         n37727, n37728, n37729, n37730, n37731, n37732, n37733, n37734,
         n37735, n37736, n37737, n37738, n37739, n37740, n37741, n37742,
         n37743, n37744, n37745, n37746, n37747, n37748, n37749, n37750,
         n37751, n37752, n37753, n37754, n37755, n37756, n37757, n37758,
         n37759, n37760, n37761, n37762, n37763, n37764, n37765, n37766,
         n37767, n37768, n37769, n37770, n37771, n37772, n37773, n37774,
         n37775, n37776, n37777, n37778, n37779, n37780, n37781, n37782,
         n37783, n37784, n37785, n37786, n37787, n37788, n37789, n37790,
         n37791, n37792, n37793, n37794, n37795, n37796, n37797, n37798,
         n37799, n37800, n37801, n37802, n37803, n37804, n37805, n37806,
         n37807, n37808, n37809, n37810, n37811, n37812, n37813, n37814,
         n37815, n37816, n37817, n37818, n37819, n37820, n37821, n37822,
         n37823, n37824, n37825, n37826, n37827, n37828, n37829, n37830,
         n37831, n37832, n37833, n37834, n37835, n37836, n37837, n37838,
         n37839, n37840, n37841, n37842, n37843, n37844, n37845, n37846,
         n37847, n37848, n37849, n37850, n37851, n37852, n37853, n37854,
         n37855, n37856, n37857, n37858, n37859, n37860, n37861, n37862,
         n37863, n37864, n37865, n37866, n37867, n37868, n37869, n37870,
         n37871, n37872, n37873, n37874, n37875, n37876, n37877, n37878,
         n37879, n37880, n37881, n37882, n37883, n37884, n37885, n37886,
         n37887, n37888, n37889, n37890, n37891, n37892, n37893, n37894,
         n37895, n37896, n37897, n37898, n37899, n37900, n37901, n37902,
         n37903, n37904, n37905, n37906, n37907, n37908, n37909, n37910,
         n37911, n37912, n37913, n37914, n37915, n37916, n37917, n37918,
         n37919, n37920, n37921, n37922, n37923, n37924, n37925, n37926,
         n37927, n37928, n37929, n37930, n37931, n37932, n37933, n37934,
         n37935, n37936, n37937, n37938, n37939, n37940, n37941, n37942,
         n37943, n37944, n37945, n37946, n37947, n37948, n37949, n37950,
         n37951, n37952, n37953, n37954, n37955, n37956, n37957, n37958,
         n37959, n37960, n37961, n37962, n37963, n37964, n37965, n37966,
         n37967, n37968, n37969, n37970, n37971, n37972, n37973, n37974,
         n37975, n37976, n37977, n37978, n37979, n37980, n37981, n37982,
         n37983, n37984, n37985, n37986, n37987, n37988, n37989, n37990,
         n37991, n37992, n37993, n37994, n37995, n37996, n37997, n37998,
         n37999, n38000, n38001, n38002, n38003, n38004, n38005, n38006,
         n38007, n38008, n38009, n38010, n38011, n38012, n38013, n38014,
         n38015, n38016, n38017, n38018, n38019, n38020, n38021, n38022,
         n38023, n38024, n38025, n38026, n38027, n38028, n38029, n38030,
         n38031, n38032, n38033, n38034, n38035, n38036, n38037, n38038,
         n38039, n38040, n38041, n38042, n38043, n38044, n38045, n38046,
         n38047, n38048, n38049, n38050, n38051, n38052, n38053, n38054,
         n38055, n38056, n38057, n38058, n38059, n38060, n38061, n38062,
         n38063, n38064, n38065, n38066, n38067, n38068, n38069, n38070,
         n38071, n38072, n38073, n38074, n38075, n38076, n38077, n38078,
         n38079, n38080, n38081, n38082, n38083, n38084, n38085, n38086,
         n38087, n38088, n38089, n38090, n38091, n38092, n38093, n38094,
         n38095, n38096, n38097, n38098, n38099, n38100, n38101, n38102,
         n38103, n38104, n38105, n38106, n38107, n38108, n38109, n38110,
         n38111, n38112, n38113, n38114, n38115, n38116, n38117, n38118,
         n38119, n38120, n38121, n38122, n38123, n38124, n38125, n38126,
         n38127, n38128, n38129, n38130, n38131, n38132, n38133, n38134,
         n38135, n38136, n38137, n38138, n38139, n38140, n38141, n38142,
         n38143, n38144, n38145, n38146, n38147, n38148, n38149, n38150,
         n38151, n38152, n38153, n38154, n38155, n38156, n38157, n38158,
         n38159, n38160, n38161, n38162, n38163, n38164, n38165, n38166,
         n38167, n38168, n38169, n38170, n38171, n38172, n38173, n38174,
         n38175, n38176, n38177, n38178, n38179, n38180, n38181, n38182,
         n38183, n38184, n38185, n38186, n38187, n38188, n38189, n38190,
         n38191, n38192, n38193, n38194, n38195, n38196, n38197, n38198,
         n38199, n38200, n38201, n38202, n38203, n38204, n38205, n38206,
         n38207, n38208, n38209, n38210, n38211, n38212, n38213, n38214,
         n38215, n38216, n38217, n38218, n38219, n38220, n38221, n38222,
         n38223, n38224, n38225, n38226, n38227, n38228, n38229, n38230,
         n38231, n38232, n38233, n38234, n38235, n38236, n38237, n38238,
         n38239, n38240, n38241, n38242, n38243, n38244, n38245, n38246,
         n38247, n38248, n38249, n38250, n38251, n38252, n38253, n38254,
         n38255, n38256, n38257, n38258, n38259, n38260, n38261, n38262,
         n38263, n38264, n38265, n38266, n38267, n38268, n38269, n38270,
         n38271, n38272, n38273, n38274, n38275, n38276, n38277, n38278,
         n38279, n38280, n38281, n38282, n38283, n38284, n38285, n38286,
         n38287, n38288, n38289, n38290, n38291, n38292, n38293, n38294,
         n38295, n38296, n38297, n38298, n38299, n38300, n38301, n38302,
         n38303, n38304, n38305, n38306, n38307, n38308, n38309, n38310,
         n38311, n38312, n38313, n38314, n38315, n38316, n38317, n38318,
         n38319, n38320, n38321, n38322, n38323, n38324, n38325, n38326,
         n38327, n38328, n38329, n38330, n38331, n38332, n38333, n38334,
         n38335, n38336, n38337, n38338, n38339, n38340, n38341, n38342,
         n38343, n38344, n38345, n38346, n38347, n38348, n38349, n38350,
         n38351, n38352, n38353, n38354, n38355, n38356, n38357, n38358,
         n38359, n38360, n38361, n38362, n38363, n38364, n38365, n38366,
         n38367, n38368, n38369, n38370, n38371, n38372, n38373, n38374,
         n38375, n38376, n38377, n38378, n38379, n38380, n38381, n38382,
         n38383, n38384, n38385, n38386, n38387, n38388, n38389, n38390,
         n38391, n38392, n38393, n38394, n38395, n38396, n38397, n38398,
         n38399, n38400, n38401, n38402, n38403, n38404, n38405, n38406,
         n38407, n38408, n38409, n38410, n38411, n38412, n38413, n38414,
         n38415, n38416, n38417, n38418, n38419, n38420, n38421, n38422,
         n38423, n38424, n38425, n38426, n38427, n38428, n38429, n38430,
         n38431, n38432, n38433, n38434, n38435, n38436, n38437, n38438,
         n38439, n38440, n38441, n38442, n38443, n38444, n38445, n38446,
         n38447, n38448, n38449, n38450, n38451, n38452, n38453, n38454,
         n38455, n38456, n38457, n38458, n38459, n38460, n38461, n38462,
         n38463, n38464, n38465, n38466, n38467, n38468, n38469, n38470,
         n38471, n38472, n38473, n38474, n38475, n38476, n38477, n38478,
         n38479, n38480, n38481, n38482, n38483, n38484, n38485, n38486,
         n38487, n38488, n38489, n38490, n38491, n38492, n38493, n38494,
         n38495, n38496, n38497, n38498, n38499, n38500, n38501, n38502,
         n38503, n38504, n38505, n38506, n38507, n38508, n38509, n38510,
         n38511, n38512, n38513, n38514, n38515, n38516, n38517, n38518,
         n38519, n38520, n38521, n38522, n38523, n38524, n38525, n38526,
         n38527, n38528, n38529, n38530, n38531, n38532, n38533, n38534,
         n38535, n38536, n38537, n38538, n38539, n38540, n38541, n38542,
         n38543, n38544, n38545, n38546, n38547, n38548, n38549, n38550,
         n38551, n38552, n38553, n38554, n38555, n38556, n38557, n38558,
         n38559, n38560, n38561, n38562, n38563, n38564, n38565, n38566,
         n38567, n38568, n38569, n38570, n38571, n38572, n38573, n38574,
         n38575, n38576, n38577, n38578, n38579, n38580, n38581, n38582,
         n38583, n38584, n38585, n38586, n38587, n38588, n38589, n38590,
         n38591, n38592, n38593, n38594, n38595, n38596, n38597, n38598,
         n38599, n38600, n38601, n38602, n38603, n38604, n38605, n38606,
         n38607, n38608, n38609, n38610, n38611, n38612, n38613, n38614,
         n38615, n38616, n38617, n38618, n38619, n38620, n38621, n38622,
         n38623, n38624, n38625, n38626, n38627, n38628, n38629, n38630,
         n38631, n38632, n38633, n38634, n38635, n38636, n38637, n38638,
         n38639, n38640, n38641, n38642, n38643, n38644, n38645, n38646,
         n38647, n38648, n38649, n38650, n38651, n38652, n38653, n38654,
         n38655, n38656, n38657, n38658, n38659, n38660, n38661, n38662,
         n38663, n38664, n38665, n38666, n38667, n38668, n38669, n38670,
         n38671, n38672, n38673, n38674, n38675, n38676, n38677, n38678,
         n38679, n38680, n38681, n38682, n38683, n38684, n38685, n38686,
         n38687, n38688, n38689, n38690, n38691, n38692, n38693, n38694,
         n38695, n38696, n38697, n38698, n38699, n38700, n38701, n38702,
         n38703, n38704, n38705, n38706, n38707, n38708, n38709, n38710,
         n38711, n38712, n38713, n38714, n38715, n38716, n38717, n38718,
         n38719, n38720, n38721, n38722, n38723, n38724, n38725, n38726,
         n38727, n38728, n38729, n38730, n38731, n38732, n38733, n38734,
         n38735, n38736, n38737, n38738, n38739, n38740, n38741, n38742,
         n38743, n38744, n38745, n38746, n38747, n38748, n38749, n38750,
         n38751, n38752, n38753, n38754, n38755, n38756, n38757, n38758,
         n38759, n38760, n38761, n38762, n38763, n38764, n38765, n38766,
         n38767, n38768, n38769, n38770, n38771, n38772, n38773, n38774,
         n38775, n38776, n38777, n38778, n38779, n38780, n38781, n38782,
         n38783, n38784, n38785, n38786, n38787, n38788, n38789, n38790,
         n38791, n38792, n38793, n38794, n38795, n38796, n38797, n38798,
         n38799, n38800, n38801, n38802, n38803, n38804, n38805, n38806,
         n38807, n38808, n38809, n38810, n38811, n38812, n38813, n38814,
         n38815, n38816, n38817, n38818, n38819, n38820, n38821, n38822,
         n38823, n38824, n38825, n38826, n38827, n38828, n38829, n38830,
         n38831, n38832, n38833, n38834, n38835, n38836, n38837, n38838,
         n38839, n38840, n38841, n38842, n38843, n38844, n38845, n38846,
         n38847, n38848, n38849, n38850, n38851, n38852, n38853, n38854,
         n38855, n38856, n38857, n38858, n38859, n38860, n38861, n38862,
         n38863, n38864, n38865, n38866, n38867, n38868, n38869, n38870,
         n38871, n38872, n38873, n38874, n38875, n38876, n38877, n38878,
         n38879, n38880, n38881, n38882, n38883, n38884, n38885, n38886,
         n38887, n38888, n38889, n38890, n38891, n38892, n38893, n38894,
         n38895, n38896, n38897, n38898, n38899, n38900, n38901, n38902,
         n38903, n38904, n38905, n38906, n38907, n38908, n38909, n38910,
         n38911, n38912, n38913, n38914, n38915, n38916, n38917, n38918,
         n38919, n38920, n38921, n38922, n38923, n38924, n38925, n38926,
         n38927, n38928, n38929, n38930, n38931, n38932, n38933, n38934,
         n38935, n38936, n38937, n38938, n38939, n38940, n38941, n38942,
         n38943, n38944, n38945, n38946, n38947, n38948, n38949, n38950,
         n38951, n38952, n38953, n38954, n38955, n38956, n38957, n38958,
         n38959, n38960, n38961, n38962, n38963, n38964, n38965, n38966,
         n38967, n38968, n38969, n38970, n38971, n38972, n38973, n38974,
         n38975, n38976, n38977, n38978, n38979, n38980, n38981, n38982,
         n38983, n38984, n38985, n38986, n38987, n38988, n38989, n38990,
         n38991, n38992, n38993, n38994, n38995, n38996, n38997, n38998,
         n38999, n39000, n39001, n39002, n39003, n39004, n39005, n39006,
         n39007, n39008, n39009, n39010, n39011, n39012, n39013, n39014,
         n39015, n39016, n39017, n39018, n39019, n39020, n39021, n39022,
         n39023, n39024, n39025, n39026, n39027, n39028, n39029, n39030,
         n39031, n39032, n39033, n39034, n39035, n39036, n39037, n39038,
         n39039, n39040, n39041, n39042, n39043, n39044, n39045, n39046,
         n39047, n39048, n39049, n39050, n39051, n39052, n39053, n39054,
         n39055, n39056, n39057, n39058, n39059, n39060, n39061, n39062,
         n39063, n39064, n39065, n39066, n39067, n39068, n39069, n39070,
         n39071, n39072, n39073, n39074, n39075, n39076, n39077, n39078,
         n39079, n39080, n39081, n39082, n39083, n39084, n39085, n39086,
         n39087, n39088, n39089, n39090, n39091, n39092, n39093, n39094,
         n39095, n39096, n39097, n39098, n39099, n39100, n39101, n39102,
         n39103, n39104, n39105, n39106, n39107, n39108, n39109, n39110,
         n39111, n39112, n39113, n39114, n39115, n39116, n39117, n39118,
         n39119, n39120, n39121, n39122, n39123, n39124, n39125, n39126,
         n39127, n39128, n39129, n39130, n39131, n39132, n39133, n39134,
         n39135, n39136, n39137, n39138, n39139, n39140, n39141, n39142,
         n39143, n39144, n39145, n39146, n39147, n39148, n39149, n39150,
         n39151, n39152, n39153, n39154, n39155, n39156, n39157, n39158,
         n39159, n39160, n39161, n39162, n39163, n39164, n39165, n39166,
         n39167, n39168, n39169, n39170, n39171, n39172, n39173, n39174,
         n39175, n39176, n39177, n39178, n39179, n39180, n39181, n39182,
         n39183, n39184, n39185, n39186, n39187, n39188, n39189, n39190,
         n39191, n39192, n39193, n39194, n39195, n39196, n39197, n39198,
         n39199, n39200, n39201, n39202, n39203, n39204, n39205, n39206,
         n39207, n39208, n39209, n39210, n39211, n39212, n39213, n39214,
         n39215, n39216, n39217, n39218, n39219, n39220, n39221, n39222,
         n39223, n39224, n39225, n39226, n39227, n39228, n39229, n39230,
         n39231, n39232, n39233, n39234, n39235, n39236, n39237, n39238,
         n39239, n39240, n39241, n39242, n39243, n39244, n39245, n39246,
         n39247, n39248, n39249, n39250, n39251, n39252, n39253, n39254,
         n39255, n39256, n39257, n39258, n39259, n39260, n39261, n39262,
         n39263, n39264, n39265, n39266, n39267, n39268, n39269, n39270,
         n39271, n39272, n39273, n39274, n39275, n39276, n39277, n39278,
         n39279, n39280, n39281, n39282, n39283, n39284, n39285, n39286,
         n39287, n39288, n39289, n39290, n39291, n39292, n39293, n39294,
         n39295, n39296, n39297, n39298, n39299, n39300, n39301, n39302,
         n39303, n39304, n39305, n39306, n39307, n39308, n39309, n39310,
         n39311, n39312, n39313, n39314, n39315, n39316, n39317, n39318,
         n39319, n39320, n39321, n39322, n39323, n39324, n39325, n39326,
         n39327, n39328, n39329, n39330, n39331, n39332, n39333, n39334,
         n39335, n39336, n39337, n39338, n39339, n39340, n39341, n39342,
         n39343, n39344, n39345, n39346, n39347, n39348, n39349, n39350,
         n39351, n39352, n39353, n39354, n39355, n39356, n39357, n39358,
         n39359, n39360, n39361, n39362, n39363, n39364, n39365, n39366,
         n39367, n39368, n39369, n39370, n39371, n39372, n39373, n39374,
         n39375, n39376, n39377, n39378, n39379, n39380, n39381, n39382,
         n39383, n39384, n39385, n39386, n39387, n39388, n39389, n39390,
         n39391, n39392, n39393, n39394, n39395, n39396, n39397, n39398,
         n39399, n39400, n39401, n39402, n39403, n39404, n39405, n39406,
         n39407, n39408, n39409, n39410, n39411, n39412, n39413, n39414,
         n39415, n39416, n39417, n39418, n39419, n39420, n39421, n39422,
         n39423, n39424, n39425, n39426, n39427, n39428, n39429, n39430,
         n39431, n39432, n39433, n39434, n39435, n39436, n39437, n39438,
         n39439, n39440, n39441, n39442, n39443, n39444, n39445, n39446,
         n39447, n39448, n39449, n39450, n39451, n39452, n39453, n39454,
         n39455, n39456, n39457, n39458, n39459, n39460, n39461, n39462,
         n39463, n39464, n39465, n39466, n39467, n39468, n39469, n39470,
         n39471, n39472, n39473, n39474, n39475, n39476, n39477, n39478,
         n39479, n39480, n39481, n39482, n39483, n39484, n39485, n39486,
         n39487, n39488, n39489, n39490, n39491, n39492, n39493, n39494,
         n39495, n39496, n39497, n39498, n39499, n39500, n39501, n39502,
         n39503, n39504, n39505, n39506, n39507, n39508, n39509, n39510,
         n39511, n39512, n39513, n39514, n39515, n39516, n39517, n39518,
         n39519, n39520, n39521, n39522, n39523, n39524, n39525, n39526,
         n39527, n39528, n39529, n39530, n39531, n39532, n39533, n39534,
         n39535, n39536, n39537, n39538, n39539, n39540, n39541, n39542,
         n39543, n39544, n39545, n39546, n39547, n39548, n39549, n39550,
         n39551, n39552, n39553, n39554, n39555, n39556, n39557, n39558,
         n39559, n39560, n39561, n39562, n39563, n39564, n39565, n39566,
         n39567, n39568, n39569, n39570, n39571, n39572, n39573, n39574,
         n39575, n39576, n39577, n39578, n39579, n39580, n39581, n39582,
         n39583, n39584, n39585, n39586, n39587, n39588, n39589, n39590,
         n39591, n39592, n39593, n39594, n39595, n39596, n39597, n39598,
         n39599, n39600, n39601, n39602, n39603, n39604, n39605, n39606,
         n39607, n39608, n39609, n39610, n39611, n39612, n39613, n39614,
         n39615, n39616, n39617, n39618, n39619, n39620, n39621, n39622,
         n39623, n39624, n39625, n39626, n39627, n39628, n39629, n39630,
         n39631, n39632, n39633, n39634, n39635, n39636, n39637, n39638,
         n39639, n39640, n39641, n39642, n39643, n39644, n39645, n39646,
         n39647, n39648, n39649, n39650, n39651, n39652, n39653, n39654,
         n39655, n39656, n39657, n39658, n39659, n39660, n39661, n39662,
         n39663, n39664, n39665, n39666, n39667, n39668, n39669, n39670,
         n39671, n39672, n39673, n39674, n39675, n39676, n39677, n39678,
         n39679, n39680, n39681, n39682, n39683, n39684, n39685, n39686,
         n39687, n39688, n39689, n39690, n39691, n39692, n39693, n39694,
         n39695, n39696, n39697, n39698, n39699, n39700, n39701, n39702,
         n39703, n39704, n39705, n39706, n39707, n39708, n39709, n39710,
         n39711, n39712, n39713, n39714, n39715, n39716, n39717, n39718,
         n39719, n39720, n39721, n39722, n39723, n39724, n39725, n39726,
         n39727, n39728, n39729, n39730, n39731, n39732, n39733, n39734,
         n39735, n39736, n39737, n39738, n39739, n39740, n39741, n39742,
         n39743, n39744, n39745, n39746, n39747, n39748, n39749, n39750,
         n39751, n39752, n39753, n39754, n39755, n39756, n39757, n39758,
         n39759, n39760, n39761, n39762, n39763, n39764, n39765, n39766,
         n39767, n39768, n39769, n39770, n39771, n39772, n39773, n39774,
         n39775, n39776, n39777, n39778, n39779, n39780, n39781, n39782,
         n39783, n39784, n39785, n39786, n39787, n39788, n39789, n39790,
         n39791, n39792, n39793, n39794, n39795, n39796, n39797, n39798,
         n39799, n39800, n39801, n39802, n39803, n39804, n39805, n39806,
         n39807, n39808, n39809, n39810, n39811, n39812, n39813, n39814,
         n39815, n39816, n39817, n39818, n39819, n39820, n39821, n39822,
         n39823, n39824, n39825, n39826, n39827, n39828, n39829, n39830,
         n39831, n39832, n39833, n39834, n39835, n39836, n39837, n39838,
         n39839, n39840, n39841, n39842, n39843, n39844, n39845, n39846,
         n39847, n39848, n39849, n39850, n39851, n39852, n39853, n39854,
         n39855, n39856, n39857, n39858, n39859, n39860, n39861, n39862,
         n39863, n39864, n39865, n39866, n39867, n39868, n39869, n39870,
         n39871, n39872, n39873, n39874, n39875, n39876, n39877, n39878,
         n39879, n39880, n39881, n39882, n39883, n39884, n39885, n39886,
         n39887, n39888, n39889, n39890, n39891, n39892, n39893, n39894,
         n39895, n39896, n39897, n39898, n39899, n39900, n39901, n39902,
         n39903, n39904, n39905, n39906, n39907, n39908, n39909, n39910,
         n39911, n39912, n39913, n39914, n39915, n39916, n39917, n39918,
         n39919, n39920, n39921, n39922, n39923, n39924, n39925, n39926,
         n39927, n39928, n39929, n39930, n39931, n39932, n39933, n39934,
         n39935, n39936, n39937, n39938, n39939, n39940, n39941, n39942,
         n39943, n39944, n39945, n39946, n39947, n39948, n39949, n39950,
         n39951, n39952, n39953, n39954, n39955, n39956, n39957, n39958,
         n39959, n39960, n39961, n39962, n39963, n39964, n39965, n39966,
         n39967, n39968, n39969, n39970, n39971, n39972, n39973, n39974,
         n39975, n39976, n39977, n39978, n39979, n39980, n39981, n39982,
         n39983, n39984, n39985, n39986, n39987, n39988, n39989, n39990,
         n39991, n39992, n39993, n39994, n39995, n39996, n39997, n39998,
         n39999, n40000, n40001, n40002, n40003, n40004, n40005, n40006,
         n40007, n40008, n40009, n40010, n40011, n40012, n40013, n40014,
         n40015, n40016, n40017, n40018, n40019, n40020, n40021, n40022,
         n40023, n40024, n40025, n40026, n40027, n40028, n40029, n40030,
         n40031, n40032, n40033, n40034, n40035, n40036, n40037, n40038,
         n40039, n40040, n40041, n40042, n40043, n40044, n40045, n40046,
         n40047, n40048, n40049, n40050, n40051, n40052, n40053, n40054,
         n40055, n40056, n40057, n40058, n40059, n40060, n40061, n40062,
         n40063, n40064, n40065, n40066, n40067, n40068, n40069, n40070,
         n40071, n40072, n40073, n40074, n40075, n40076, n40077, n40078,
         n40079, n40080, n40081, n40082, n40083, n40084, n40085, n40086,
         n40087, n40088, n40089, n40090, n40091, n40092, n40093, n40094,
         n40095, n40096, n40097, n40098, n40099, n40100, n40101, n40102,
         n40103, n40104, n40105, n40106, n40107, n40108, n40109, n40110,
         n40111, n40112, n40113, n40114, n40115, n40116, n40117, n40118,
         n40119, n40120, n40121, n40122, n40123, n40124, n40125, n40126,
         n40127, n40128, n40129, n40130, n40131, n40132, n40133, n40134,
         n40135, n40136, n40137, n40138, n40139, n40140, n40141, n40142,
         n40143, n40144, n40145, n40146, n40147, n40148, n40149, n40150,
         n40151, n40152, n40153, n40154, n40155, n40156, n40157, n40158,
         n40159, n40160, n40161, n40162, n40163, n40164, n40165, n40166,
         n40167, n40168, n40169, n40170, n40171, n40172, n40173, n40174,
         n40175, n40176, n40177, n40178, n40179, n40180, n40181, n40182,
         n40183, n40184, n40185, n40186, n40187, n40188, n40189, n40190,
         n40191, n40192, n40193, n40194, n40195, n40196, n40197, n40198,
         n40199, n40200, n40201, n40202, n40203, n40204, n40205, n40206,
         n40207, n40208, n40209, n40210, n40211, n40212, n40213, n40214,
         n40215, n40216, n40217, n40218, n40219, n40220, n40221, n40222,
         n40223, n40224, n40225, n40226, n40227, n40228, n40229, n40230,
         n40231, n40232, n40233, n40234, n40235, n40236, n40237, n40238,
         n40239, n40240, n40241, n40242, n40243, n40244, n40245, n40246,
         n40247, n40248, n40249, n40250, n40251, n40252, n40253, n40254,
         n40255, n40256, n40257, n40258, n40259, n40260, n40261, n40262,
         n40263, n40264, n40265, n40266, n40267, n40268, n40269, n40270,
         n40271, n40272, n40273, n40274, n40275, n40276, n40277, n40278,
         n40279, n40280, n40281, n40282, n40283, n40284, n40285, n40286,
         n40287, n40288, n40289, n40290, n40291, n40292, n40293, n40294,
         n40295, n40296, n40297, n40298, n40299, n40300, n40301, n40302,
         n40303, n40304, n40305, n40306, n40307, n40308, n40309, n40310,
         n40311, n40312, n40313, n40314, n40315, n40316, n40317, n40318,
         n40319, n40320, n40321, n40322, n40323, n40324, n40325, n40326,
         n40327, n40328, n40329, n40330, n40331, n40332, n40333, n40334,
         n40335, n40336, n40337, n40338, n40339, n40340, n40341, n40342,
         n40343, n40344, n40345, n40346, n40347, n40348, n40349, n40350,
         n40351, n40352, n40353, n40354, n40355, n40356, n40357, n40358,
         n40359, n40360, n40361, n40362, n40363, n40364, n40365, n40366,
         n40367, n40368, n40369, n40370, n40371, n40372, n40373, n40374,
         n40375, n40376, n40377, n40378, n40379, n40380, n40381, n40382,
         n40383, n40384, n40385, n40386, n40387, n40388, n40389, n40390,
         n40391, n40392, n40393, n40394, n40395, n40396, n40397, n40398,
         n40399, n40400, n40401, n40402, n40403, n40404, n40405, n40406,
         n40407, n40408, n40409, n40410, n40411, n40412, n40413, n40414,
         n40415, n40416, n40417, n40418, n40419, n40420, n40421, n40422,
         n40423, n40424, n40425, n40426, n40427, n40428, n40429, n40430,
         n40431, n40432, n40433, n40434, n40435, n40436, n40437, n40438,
         n40439, n40440, n40441, n40442, n40443, n40444, n40445, n40446,
         n40447, n40448, n40449, n40450, n40451, n40452, n40453, n40454,
         n40455, n40456, n40457, n40458, n40459, n40460, n40461, n40462,
         n40463, n40464, n40465, n40466, n40467, n40468, n40469, n40470,
         n40471, n40472, n40473, n40474, n40475, n40476, n40477, n40478,
         n40479, n40480, n40481, n40482, n40483, n40484, n40485, n40486,
         n40487, n40488, n40489, n40490, n40491, n40492, n40493, n40494,
         n40495, n40496, n40497, n40498, n40499, n40500, n40501, n40502,
         n40503, n40504, n40505, n40506, n40507, n40508, n40509, n40510,
         n40511, n40512, n40513, n40514, n40515, n40516, n40517, n40518,
         n40519, n40520, n40521, n40522, n40523, n40524, n40525, n40526,
         n40527, n40528, n40529, n40530, n40531, n40532, n40533, n40534,
         n40535, n40536, n40537, n40538, n40539, n40540, n40541, n40542,
         n40543, n40544, n40545, n40546, n40547, n40548, n40549, n40550,
         n40551, n40552, n40553, n40554, n40555, n40556, n40557, n40558,
         n40559, n40560, n40561, n40562, n40563, n40564, n40565, n40566,
         n40567, n40568, n40569, n40570, n40571, n40572, n40573, n40574,
         n40575, n40576, n40577, n40578, n40579, n40580, n40581, n40582,
         n40583, n40584, n40585, n40586, n40587, n40588, n40589, n40590,
         n40591, n40592, n40593, n40594, n40595, n40596, n40597, n40598,
         n40599, n40600, n40601, n40602, n40603, n40604, n40605, n40606,
         n40607, n40608, n40609, n40610, n40611, n40612, n40613, n40614,
         n40615, n40616, n40617, n40618, n40619, n40620, n40621, n40622,
         n40623, n40624, n40625, n40626, n40627, n40628, n40629, n40630,
         n40631, n40632, n40633, n40634, n40635, n40636, n40637, n40638,
         n40639, n40640, n40641, n40642, n40643, n40644, n40645, n40646,
         n40647, n40648, n40649, n40650, n40651, n40652, n40653, n40654,
         n40655, n40656, n40657, n40658, n40659, n40660, n40661, n40662,
         n40663, n40664, n40665, n40666, n40667, n40668, n40669, n40670,
         n40671, n40672, n40673, n40674, n40675, n40676, n40677, n40678,
         n40679, n40680, n40681, n40682, n40683, n40684, n40685, n40686,
         n40687, n40688, n40689, n40690, n40691, n40692, n40693, n40694,
         n40695, n40696, n40697, n40698, n40699, n40700, n40701, n40702,
         n40703, n40704, n40705, n40706, n40707, n40708, n40709, n40710,
         n40711, n40712, n40713, n40714, n40715, n40716, n40717, n40718,
         n40719, n40720, n40721, n40722, n40723, n40724, n40725, n40726,
         n40727, n40728, n40729, n40730, n40731, n40732, n40733, n40734,
         n40735, n40736, n40737, n40738, n40739, n40740, n40741, n40742,
         n40743, n40744, n40745, n40746, n40747, n40748, n40749, n40750,
         n40751, n40752, n40753, n40754, n40755, n40756, n40757, n40758,
         n40759, n40760, n40761, n40762, n40763, n40764, n40765, n40766,
         n40767, n40768, n40769, n40770, n40771, n40772, n40773, n40774,
         n40775, n40776, n40777, n40778, n40779, n40780, n40781, n40782,
         n40783, n40784, n40785, n40786, n40787, n40788, n40789, n40790,
         n40791, n40792, n40793, n40794, n40795, n40796, n40797, n40798,
         n40799, n40800, n40801, n40802, n40803, n40804, n40805, n40806,
         n40807, n40808, n40809, n40810, n40811, n40812, n40813, n40814,
         n40815, n40816, n40817, n40818, n40819, n40820, n40821, n40822,
         n40823, n40824, n40825, n40826, n40827, n40828, n40829, n40830,
         n40831, n40832, n40833, n40834, n40835, n40836, n40837, n40838,
         n40839, n40840, n40841, n40842, n40843, n40844, n40845, n40846,
         n40847, n40848, n40849, n40850, n40851, n40852, n40853, n40854,
         n40855, n40856, n40857, n40858, n40859, n40860, n40861, n40862,
         n40863, n40864, n40865, n40866, n40867, n40868, n40869, n40870,
         n40871, n40872, n40873, n40874, n40875, n40876, n40877, n40878,
         n40879, n40880, n41521, n41522, n41523, n41524, n41525, n41526,
         n41527, n41528, n41529, n41530, n41531, n41532, n41533, n41534,
         n41535, n41536, n41537, n41538, n41539, n41540, n41541, n41542,
         n41543, n41544, n41545, n41546, n41547, n41548, n41549, n41550,
         n41551, n41552, n41553, n41554, n41555, n41556, n41557, n41558,
         n41559, n41560, n41561, n41562, n41563, n41564, n41565, n41566,
         n41567, n41568, n41569, n41570, n41571, n41572, n41573, n41574,
         n41575, n41576, n41577, n41578, n41579, n41580, n41581, n41582,
         n41583, n41584, n41585, n41586, n41587, n41588, n41589, n41590,
         n41591, n41592, n41593, n41594, n41595, n41596, n41597, n41598,
         n41599, n41600, n41601, n41602, n41603, n41604, n41605, n41606,
         n41607, n41608, n41609, n41610, n41611, n41612, n41613, n41614,
         n41615, n41616, n41617, n41618, n41619, n41620, n41621, n41622,
         n41623, n41624, n41625, n41626, n41627, n41628, n41629, n41630,
         n41631, n41632, n41633, n41634, n41635, n41636, n41637, n41638,
         n41639, n41640, n41641, n41642, n41643, n41644, n41645, n41646,
         n41647, n41648, n41649, n41650, n41651, n41652, n41653, n41654,
         n41655, n41656, n41657, n41658, n41659, n41660, n41661, n41662,
         n41663, n41664, n41665, n41666, n41667, n41668, n41669, n41670,
         n41671, n41672, n41673, n41674, n41675, n41676, n41677, n41678,
         n41679, n41680, n41681, n41682, n41683, n41684, n41685, n41686,
         n41687, n41688, n41689, n41690, n41691, n41692, n41693, n41694,
         n41695, n41696, n41697, n41698, n41699, n41700, n41701, n41702,
         n41703, n41704, n41705, n41706, n41707, n41708, n41709, n41710,
         n41711, n41712, n41713, n41714, n41715, n41716, n41717, n41718,
         n41719, n41720, n41721, n41722, n41723, n41724, n41725, n41726,
         n41727, n41728, n41729, n41730, n41731, n41732, n41733, n41734,
         n41735, n41736, n41737, n41738, n41739, n41740, n41741, n41742,
         n41743, n41744, n41745, n41746, n41747, n41748, n41749, n41750,
         n41751, n41752, n41753, n41754, n41755, n41756, n41757, n41758,
         n41759, n41760, n41761, n41762, n41763, n41764, n41765, n41766,
         n41767, n41768, n41769, n41770, n41771, n41772, n41773, n41774,
         n41775, n41776, n41777, n41778, n41779, n41780, n41781, n41782,
         n41783, n41784, n41785, n41786, n41787, n41788, n41789, n41790,
         n41791, n41792, n41793, n41794, n41795, n41796, n41797, n41798,
         n41799, n41800, n41801, n41802, n41803, n41804, n41805, n41806,
         n41807, n41808, n41809, n41810, n41811, n41812, n41813, n41814,
         n41815, n41816, n41817, n41818, n41819, n41820, n41821, n41822,
         n41823, n41824, n41825, n41826, n41827, n41828, n41829, n41830,
         n41831, n41832, n41833, n41834, n41835, n41836, n41837, n41838,
         n41839, n41840, n41841, n41842, n41843, n41844, n41845, n41846,
         n41847, n41848, n41849, n41850, n41851, n41852, n41853, n41854,
         n41855, n41856, n41857, n41858, n41859, n41860, n41861, n41862,
         n41863, n41864, n41865, n41866, n41867, n41868, n41869, n41870,
         n41871, n41872, n41873, n41874, n41875, n41876, n41877, n41878,
         n41879, n41880, n41881, n41882, n41883, n41884, n41885, n41886,
         n41887, n41888, n41889, n41890, n41891, n41892, n41893, n41894,
         n41895, n41896, n41897, n41898, n41899, n41900, n41901, n41902,
         n41903, n41904, n41905, n41906, n41907, n41908, n41909, n41910,
         n41911, n41912, n41913, n41914, n41915, n41916, n41917, n41918,
         n41919, n41920, n41921, n41922, n41923, n41924, n41925, n41926,
         n41927, n41928, n41929, n41930, n41931, n41932, n41933, n41934,
         n41935, n41936, n41937, n41938, n41939, n41940, n41941, n41942,
         n41943, n41944, n41945, n41946, n41947, n41948, n41949, n41950,
         n41951, n41952, n41953, n41954, n41955, n41956, n41957, n41958,
         n41959, n41960, n41961, n41962, n41963, n41964, n41965, n41966,
         n41967, n41968, n41969, n41970, n41971, n41972, n41973, n41974,
         n41975, n41976, n41977, n41978, n41979, n41980, n41981, n41982,
         n41983, n41984, n41985, n41986, n41987, n41988, n41989, n41990,
         n41991, n41992, n41993, n41994, n41995, n41996, n41997, n41998,
         n41999, n42000, n42001, n42002, n42003, n42004, n42005, n42006,
         n42007, n42008, n42009, n42010, n42011, n42012, n42013, n42014,
         n42015, n42016, n42017, n42018, n42019, n42020, n42021, n42022,
         n42023, n42024, n42025, n42026, n42027, n42028, n42029, n42030,
         n42031, n42032, n42033, n42034, n42035, n42036, n42037, n42038,
         n42039, n42040, n42041, n42042, n42043, n42044, n42045, n42046,
         n42047, n42048, n42049, n42050, n42051, n42052, n42053, n42054,
         n42055, n42056, n42057, n42058, n42059, n42060, n42061, n42062,
         n42063, n42064, n42065, n42066, n42067, n42068, n42069, n42070,
         n42071, n42072, n42073, n42074, n42075, n42076, n42077, n42078,
         n42079, n42080, n42081, n42082, n42083, n42084, n42085, n42086,
         n42087, n42088, n42089, n42090, n42091, n42092, n42093, n42094,
         n42095, n42096, n42097, n42098, n42099, n42100, n42101, n42102,
         n42103, n42104, n42105, n42106, n42107, n42108, n42109, n42110,
         n42111, n42112, n42113, n42114, n42115, n42116, n42117, n42118,
         n42119, n42120, n42121, n42122, n42123, n42124, n42125, n42126,
         n42127, n42128, n42129, n42130, n42131, n42132, n42133, n42134,
         n42135, n42136, n42137, n42138, n42139, n42140, n42141, n42142,
         n42143, n42144, n42145, n42146, n42147, n42148, n42149, n42150,
         n42151, n42152, n42153, n42154, n42155, n42156, n42157, n42158,
         n42159, n42160, n42161, n42162, n42163, n42164, n42165, n42166,
         n42167, n42168, n42169, n42170, n42171, n42172, n42173, n42174,
         n42175, n42176, n42177, n42178, n42179, n42180, n42181, n42182,
         n42183, n42184, n42185, n42186, n42187, n42188, n42189, n42190,
         n42191, n42192, n42193, n42194, n42195, n42196, n42197, n42198,
         n42199, n42200, n42201, n42202, n42203, n42204, n42205, n42206,
         n42207, n42208, n42209, n42210, n42211, n42212, n42213, n42214,
         n42215, n42216, n42217, n42218, n42219, n42220, n42221, n42222,
         n42223, n42224, n42225, n42226, n42227, n42228, n42229, n42230,
         n42231, n42232, n42233, n42234, n42235, n42236, n42237, n42238,
         n42239, n42240, n42241, n42242, n42243, n42244, n42245, n42246,
         n42247, n42248, n42249, n42250, n42251, n42252, n42253, n42254,
         n42255, n42256, n42257, n42258, n42259, n42260, n42261, n42262,
         n42263, n42264, n42265, n42266, n42267, n42268, n42269, n42270,
         n42271, n42272, n42273, n42274, n42275, n42276, n42277, n42278,
         n42279, n42280, n42281, n42282, n42283, n42284, n42285, n42286,
         n42287, n42288, n42289, n42290, n42291, n42292, n42293, n42294,
         n42295, n42296, n42297, n42298, n42299, n42300, n42301, n42302,
         n42303, n42304, n42305, n42306, n42307, n42308, n42309, n42310,
         n42311, n42312, n42313, n42314, n42315, n42316, n42317, n42318,
         n42319, n42320, n42321, n42322, n42323, n42324, n42325, n42326,
         n42327, n42328, n42329, n42330, n42331, n42332, n42333, n42334,
         n42335, n42336, n42337, n42338, n42339, n42340, n42341, n42342,
         n42343, n42344, n42345, n42346, n42347, n42348, n42349, n42350,
         n42351, n42352, n42353, n42354, n42355, n42356, n42357, n42358,
         n42359, n42360, n42361, n42362, n42363, n42364, n42365, n42366,
         n42367, n42368, n42369, n42370, n42371, n42372, n42373, n42374,
         n42375, n42376, n42377, n42378, n42379, n42380, n42381, n42382,
         n42383, n42384, n42385, n42386, n42387, n42388, n42389, n42390,
         n42391, n42392, n42393, n42394, n42395, n42396, n42397, n42398,
         n42399, n42400, n42401, n42402, n42403, n42404, n42405, n42406,
         n42407, n42408, n42409, n42410, n42411, n42412, n42413, n42414,
         n42415, n42416, n42417, n42418, n42419, n42420, n42421, n42422,
         n42423, n42424, n42425, n42426, n42427, n42428, n42429, n42430,
         n42431, n42432, n42433, n42434, n42435, n42436, n42437, n42438,
         n42439, n42440, n42441, n42442, n42443, n42444, n42445, n42446,
         n42447, n42448, n42449, n42450, n42451, n42452, n42453, n42454,
         n42455, n42456, n42457, n42458, n42459, n42460, n42461, n42462,
         n42463, n42464, n42465, n42466, n42467, n42468, n42469, n42470,
         n42471, n42472, n42473, n42474, n42475, n42476, n42477, n42478,
         n42479, n42480, n42481, n42482, n42483, n42484, n42485, n42486,
         n42487, n42488, n42489, n42490, n42491, n42492, n42493, n42494,
         n42495, n42496, n42497, n42498, n42499, n42500, n42501, n42502,
         n42503, n42504, n42505, n42506, n42507, n42508, n42509, n42510,
         n42511, n42512, n42513, n42514, n42515, n42516, n42517, n42518,
         n42519, n42520, n42521, n42522, n42523, n42524, n42525, n42526,
         n42527, n42528, n42529, n42530, n42531, n42532, n42533, n42534,
         n42535, n42536, n42537, n42538, n42539, n42540, n42541, n42542,
         n42543, n42544, n42545, n42546, n42547, n42548, n42549, n42550,
         n42551, n42552, n42553, n42554, n42555, n42556, n42557, n42558,
         n42559, n42560, n42561, n42562, n42563, n42564, n42565, n42566,
         n42567, n42568, n42569, n42570, n42571, n42572, n42573, n42574,
         n42575, n42576, n42577, n42578, n42579, n42580, n42581, n42582,
         n42583, n42584, n42585, n42586, n42587, n42588, n42589, n42590,
         n42591, n42592, n42593, n42594, n42595, n42596, n42597, n42598,
         n42599, n42600, n42601, n42602, n42603, n42604, n42605, n42606,
         n42607, n42608, n42609, n42610, n42611, n42612, n42613, n42614,
         n42615, n42616, n42617, n42618, n42619, n42620, n42621, n42622,
         n42623, n42624, n42625, n42626, n42627, n42628, n42629, n42630,
         n42631, n42632, n42633, n42634, n42635, n42636, n42637, n42638,
         n42639, n42640, n42641, n42642, n42643, n42644, n42645, n42646,
         n42647, n42648, n42649, n42650, n42651, n42652, n42653, n42654,
         n42655, n42656, n42657, n42658, n42659, n42660, n42661, n42662,
         n42663, n42664, n42665, n42666, n42667, n42668, n42669, n42670,
         n42671, n42672, n42673, n42674, n42675, n42676, n42677, n42678,
         n42679, n42680, n42681, n42682, n42683, n42684, n42685, n42686,
         n42687, n42688, n42689, n42690, n42691, n42692, n42693, n42694,
         n42695, n42696, n42697, n42698, n42699, n42700, n42701, n42702,
         n42703, n42704, n42705, n42706, n42707, n42708, n42709, n42710,
         n42711, n42712, n42713, n42714, n42715, n42716, n42717, n42718,
         n42719, n42720, n42721, n42722, n42723, n42724, n42725, n42726,
         n42727, n42728, n42729, n42730, n42731, n42732, n42733, n42734,
         n42735, n42736, n42737, n42738, n42739, n42740, n42741, n42742,
         n42743, n42744, n42745, n42746, n42747, n42748, n42749, n42750,
         n42751, n42752, n42753, n42754, n42755, n42756, n42757, n42758,
         n42759, n42760, n42761, n42762, n42763, n42764, n42765, n42766,
         n42767, n42768, n42769, n42770, n42771, n42772, n42773, n42774,
         n42775, n42776, n42777, n42778, n42779, n42780, n42781, n42782,
         n42783, n42784, n42785, n42786, n42787, n42788, n42789, n42790,
         n42791, n42792, n42793, n42794, n42795, n42796, n42797, n42798,
         n42799, n42800, n42801, n42802, n42803, n42804, n42805, n42806,
         n42807, n42808, n42809, n42810, n42811, n42812, n42813, n42814,
         n42815, n42816, n42817, n42818, n42819, n42820, n42821, n42822,
         n42823, n42824, n42825, n42826, n42827, n42828, n42829, n42830,
         n42831, n42832, n42833, n42834, n42835, n42836, n42837, n42838,
         n42839, n42840, n42841, n42842, n42843, n42844, n42845, n42846,
         n42847, n42848, n42849, n42850, n42851, n42852, n42853, n42854,
         n42855, n42856, n42857, n42858, n42859, n42860, n42861, n42862,
         n42863, n42864, n42865, n42866, n42867, n42868, n42869, n42870,
         n42871, n42872, n42873, n42874, n42875, n42876, n42877, n42878,
         n42879, n42880, n42881, n42882, n42883, n42884, n42885, n42886,
         n42887, n42888, n42889, n42890, n42891, n42892, n42893, n42894,
         n42895, n42896, n42897, n42898, n42899, n42900, n42901, n42902,
         n42903, n42904, n42905, n42906, n42907, n42908, n42909, n42910,
         n42911, n42912, n42913, n42914, n42915, n42916, n42917, n42918,
         n42919, n42920, n42921, n42922, n42923, n42924, n42925, n42926,
         n42927, n42928, n42929, n42930, n42931, n42932, n42933, n42934,
         n42935, n42936, n42937, n42938, n42939, n42940, n42941, n42942,
         n42943, n42944, n42945, n42946, n42947, n42948, n42949, n42950,
         n42951, n42952, n42953, n42954, n42955, n42956, n42957, n42958,
         n42959, n42960, n42961, n42962, n42963, n42964, n42965, n42966,
         n42967, n42968, n42969, n42970, n42971, n42972, n42973, n42974,
         n42975, n42976, n42977, n42978, n42979, n42980, n42981, n42982,
         n42983, n42984, n42985, n42986, n42987, n42988, n42989, n42990,
         n42991, n42992, n42993, n42994, n42995, n42996, n42997, n42998,
         n42999, n43000, n43001, n43002, n43003, n43004, n43005, n43006,
         n43007, n43008, n43009, n43010, n43011, n43012, n43013, n43014,
         n43015, n43016, n43017, n43018, n43019, n43020, n43021, n43022,
         n43023, n43024, n43025, n43026, n43027, n43028, n43029, n43030,
         n43031, n43032, n43033, n43034, n43035, n43036, n43037, n43038,
         n43039, n43040, n43041, n43042, n43043, n43044, n43045, n43046,
         n43047, n43048, n43049, n43050, n43051, n43052, n43053, n43054,
         n43055, n43056, n43057, n43058, n43059, n43060, n43061, n43062,
         n43063, n43064, n43065, n43066, n43067, n43068, n43069, n43070,
         n43071, n43072, n43073, n43074, n43075, n43076, n43077, n43078,
         n43079, n43080, n43081, n43082, n43083, n43084, n43085, n43086,
         n43087, n43088, n43089, n43090, n43091, n43092, n43093, n43094,
         n43095, n43096, n43097, n43098, n43099, n43100, n43101, n43102,
         n43103, n43104, n43105, n43106, n43107, n43108, n43109, n43110,
         n43111, n43112, n43113, n43114, n43115, n43116, n43117, n43118,
         n43119, n43120, n43121, n43122, n43123, n43124, n43125, n43126,
         n43127, n43128, n43129, n43130, n43131, n43132, n43133, n43134,
         n43135, n43136, n43137, n43138, n43139, n43140, n43141, n43142,
         n43143, n43144, n43145, n43146, n43147, n43148, n43149, n43150,
         n43151, n43152, n43153, n43154, n43155, n43156, n43157, n43158,
         n43159, n43160, n43161, n43162, n43163, n43164, n43165, n43166,
         n43167, n43168, n43169, n43170, n43171, n43172, n43173, n43174,
         n43175, n43176, n43177, n43178, n43179, n43180, n43181, n43182,
         n43183, n43184, n43185, n43186, n43187, n43188, n43189, n43190,
         n43191, n43192, n43193, n43194, n43195, n43196, n43197, n43198,
         n43199, n43200, n43201, n43202, n43203, n43204, n43205, n43206,
         n43207, n43208, n43209, n43210, n43211, n43212, n43213, n43214,
         n43215, n43216, n43217, n43218, n43219, n43220, n43221, n43222,
         n43223, n43224, n43225, n43226, n43227, n43228, n43229, n43230,
         n43231, n43232, n43233, n43234, n43235, n43236, n43237, n43238,
         n43239, n43240, n43241, n43242, n43243, n43244, n43245, n43246,
         n43247, n43248, n43249, n43250, n43251, n43252, n43253, n43254,
         n43255, n43256, n43257, n43258, n43259, n43260, n43261, n43262,
         n43263, n43264, n43265, n43266, n43267, n43268, n43269, n43270,
         n43271, n43272, n43273, n43274, n43275, n43276, n43277, n43278,
         n43279, n43280, n43281, n43282, n43283, n43284, n43285, n43286,
         n43287, n43288, n43289, n43290, n43291, n43292, n43293, n43294,
         n43295, n43296, n43297, n43298, n43299, n43300, n43301, n43302,
         n43303, n43304, n43305, n43306, n43307, n43308, n43309, n43310,
         n43311, n43312, n43313, n43314, n43315, n43316, n43317, n43318,
         n43319, n43320, n43321, n43322, n43323, n43324, n43325, n43326,
         n43327, n43328, n43329, n43330, n43331, n43332, n43333, n43334,
         n43335, n43336, n43337, n43338, n43339, n43340, n43341, n43342,
         n43343, n43344, n43345, n43346, n43347, n43348, n43349, n43350,
         n43351, n43352, n43353, n43354, n43355, n43356, n43357, n43358,
         n43359, n43360, n43361, n43362, n43363, n43364, n43365, n43366,
         n43367, n43368, n43369, n43370, n43371, n43372, n43373, n43374,
         n43375, n43376, n43377, n43378, n43379, n43380, n43381, n43382,
         n43383, n43384, n43385, n43386, n43387, n43388, n43389, n43390,
         n43391, n43392, n43393, n43394, n43395, n43396, n43397, n43398,
         n43399, n43400, n43401, n43402, n43403, n43404, n43405, n43406,
         n43407, n43408, n43409, n43410, n43411, n43412, n43413, n43414,
         n43415, n43416, n43417, n43418, n43419, n43420, n43421, n43422,
         n43423, n43424, n43425, n43426, n43427, n43428, n43429, n43430,
         n43431, n43432, n43433, n43434, n43435, n43436, n43437, n43438,
         n43439, n43440, n43441, n43442, n43443, n43444, n43445, n43446,
         n43447, n43448, n43449, n43450, n43451, n43452, n43453, n43454,
         n43455, n43456, n43457, n43458, n43459, n43460, n43461, n43462,
         n43463, n43464, n43465, n43466, n43467, n43468, n43469, n43470,
         n43471, n43472, n43473, n43474, n43475, n43476, n43477, n43478,
         n43479, n43480, n43481, n43482, n43483, n43484, n43485, n43486,
         n43487, n43488, n43489, n43490, n43491, n43492, n43493, n43494,
         n43495, n43496, n43497, n43498, n43499, n43500, n43501, n43502,
         n43503, n43504, n43505, n43506, n43507, n43508, n43509, n43510,
         n43511, n43512, n43513, n43514, n43515, n43516, n43517, n43518,
         n43519, n43520, n43521, n43522, n43523, n43524, n43525, n43526,
         n43527, n43528, n43529, n43530, n43531, n43532, n43533, n43534,
         n43535, n43536, n43537, n43538, n43539, n43540, n43541, n43542,
         n43543, n43544, n43545, n43546, n43547, n43548, n43549, n43550,
         n43551, n43552, n43553, n43554, n43555, n43556, n43557, n43558,
         n43559, n43560, n43561, n43562, n43563, n43564, n43565, n43566,
         n43567, n43568, n43569, n43570, n43571, n43572, n43573, n43574,
         n43575, n43576, n43577, n43578, n43579, n43580, n43581, n43582,
         n43583, n43584, n43585, n43586, n43587, n43588, n43589, n43590,
         n43591, n43592, n43593, n43594, n43595, n43596, n43597, n43598,
         n43599, n43600, n43601, n43602, n43603, n43604, n43605, n43606,
         n43607, n43608, n43609, n43610, n43611, n43612, n43613, n43614,
         n43615, n43616, n43617, n43618, n43619, n43620, n43621, n43622,
         n43623, n43624, n43625, n43626, n43627, n43628, n43629, n43630,
         n43631, n43632, n43633, n43634, n43635, n43636, n43637, n43638,
         n43639, n43640, n43641, n43642, n43643, n43644, n43645, n43646,
         n43647, n43648, n43649, n43650, n43651, n43652, n43653, n43654,
         n43655, n43656, n43657, n43658, n43659, n43660, n43661, n43662,
         n43663, n43664, n43665, n43666, n43667, n43668, n43669, n43670,
         n43671, n43672, n43673, n43674, n43675, n43676, n43677, n43678,
         n43679, n43680, n43681, n43682, n43683, n43684, n43685, n43686,
         n43687, n43688, n43689, n43690, n43691, n43692, n43693, n43694,
         n43695, n43696, n43697, n43698, n43699, n43700, n43701, n43702,
         n43703, n43704, n43705, n43706, n43707, n43708, n43709, n43710,
         n43711, n43712, n43713, n43714, n43715, n43716, n43717, n43718,
         n43719, n43720, n43721, n43722, n43723, n43724, n43725, n43726,
         n43727, n43728, n43729, n43730, n43731, n43732, n43733, n43734,
         n43735, n43736, n43737, n43738, n43739, n43740, n43741, n43742,
         n43743, n43744, n43745, n43746, n43747, n43748, n43749, n43750,
         n43751, n43752, n43753, n43754, n43755, n43756, n43757, n43758,
         n43759, n43760, n43761, n43762, n43763, n43764, n43765, n43766,
         n43767, n43768, n43769, n43770, n43771, n43772, n43773, n43774,
         n43775, n43776, n43777, n43778, n43779, n43780, n43781, n43782,
         n43783, n43784, n43785, n43786, n43787, n43788, n43789, n43790,
         n43791, n43792, n43793, n43794, n43795, n43796, n43797, n43798,
         n43799, n43800, n43801, n43802, n43803, n43804, n43805, n43806,
         n43807, n43808, n43809, n43810, n43811, n43812, n43813, n43814,
         n43815, n43816, n43817, n43818, n43819, n43820, n43821, n43822,
         n43823, n43824, n43825, n43826, n43827, n43828, n43829, n43830,
         n43831, n43832, n43833, n43834, n43835, n43836, n43837, n43838,
         n43839, n43840, n43841, n43842, n43843, n43844, n43845, n43846,
         n43847, n43848, n43849, n43850, n43851, n43852, n43853, n43854,
         n43855, n43856, n43857, n43858, n43859, n43860, n43861, n43862,
         n43863, n43864, n43865, n43866, n43867, n43868, n43869, n43870,
         n43871, n43872, n43873, n43874, n43875, n43876, n43877, n43878,
         n43879, n43880, n43881, n43882, n43883, n43884, n43885, n43886,
         n43887, n43888, n43889, n43890, n43891, n43892, n43893, n43894,
         n43895, n43896, n43897, n43898, n43899, n43900, n43901, n43902,
         n43903, n43904, n43905, n43906, n43907, n43908, n43909, n43910,
         n43911, n43912, n43913, n43914, n43915, n43916, n43917, n43918,
         n43919, n43920, n43921, n43922, n43923, n43924, n43925, n43926,
         n43927, n43928, n43929, n43930, n43931, n43932, n43933, n43934,
         n43935, n43936, n43937, n43938, n43939, n43940, n43941, n43942,
         n43943, n43944, n43945, n43946, n43947, n43948, n43949, n43950,
         n43951, n43952, n43953, n43954, n43955, n43956, n43957, n43958,
         n43959, n43960, n43961, n43962, n43963, n43964, n43965, n43966,
         n43967, n43968, n43969, n43970, n43971, n43972, n43973, n43974,
         n43975, n43976, n43977, n43978, n43979, n43980, n43981, n43982,
         n43983, n43984, n43985, n43986, n43987, n43988, n43989, n43990,
         n43991, n43992, n43993, n43994, n43995, n43996, n43997, n43998,
         n43999, n44000, n44001, n44002, n44003, n44004, n44005, n44006,
         n44007, n44008, n44009, n44010, n44011, n44012, n44013, n44014,
         n44015, n44016, n44017, n44018, n44019, n44020, n44021, n44022,
         n44023, n44024, n44025, n44026, n44027, n44028, n44029, n44030,
         n44031, n44032, n44033, n44034, n44035, n44036, n44037, n44038,
         n44039, n44040, n44041, n44042, n44043, n44044, n44045, n44046,
         n44047, n44048, n44049, n44050, n44051, n44052, n44053, n44054,
         n44055, n44056, n44057, n44058, n44059, n44060, n44061, n44062,
         n44063, n44064, n44065, n44066, n44067, n44068, n44069, n44070,
         n44071, n44072, n44073, n44074, n44075, n44076, n44077, n44078,
         n44079, n44080, n44081, n44082, n44083, n44084, n44085, n44086,
         n44087, n44088, n44089, n44090, n44091, n44092, n44093, n44094,
         n44095, n44096, n44097, n44098, n44099, n44100, n44101, n44102,
         n44103, n44104, n44105, n44106, n44107, n44108, n44109, n44110,
         n44111, n44112, n44113, n44114, n44115, n44116, n44117, n44118,
         n44119, n44120, n44121, n44122, n44123, n44124, n44125, n44126,
         n44127, n44128, n44129, n44130, n44131, n44132, n44133, n44134,
         n44135, n44136, n44137, n44138, n44139, n44140, n44141, n44142,
         n44143, n44144, n44145, n44146, n44147, n44148, n44149, n44150,
         n44151, n44152, n44153, n44154, n44155, n44156, n44157, n44158,
         n44159, n44160, n44161, n44162, n44163, n44164, n44165, n44166,
         n44167, n44168, n44169, n44170, n44171, n44172, n44173, n44174,
         n44175, n44176, n44177, n44178, n44179, n44180, n44181, n44182,
         n44183, n44184, n44185, n44186, n44187, n44188, n44189, n44190,
         n44191, n44192, n44193, n44194, n44195, n44196, n44197, n44198,
         n44199, n44200, n44201, n44202, n44203, n44204, n44205, n44206,
         n44207, n44208, n44209, n44210, n44211, n44212, n44213, n44214,
         n44215, n44216, n44217, n44218, n44219, n44220, n44221, n44222,
         n44223, n44224, n44225, n44226, n44227, n44228, n44229, n44230,
         n44231, n44232, n44233, n44234, n44235, n44236, n44237, n44238,
         n44239, n44240, n44241, n44242, n44243, n44244, n44245, n44246,
         n44247, n44248, n44249, n44250, n44251, n44252, n44253, n44254,
         n44255, n44256, n44257, n44258, n44259, n44260, n44261, n44262,
         n44263, n44264, n44265, n44266, n44267, n44268, n44269, n44270,
         n44271, n44272, n44273, n44274, n44275, n44276, n44277, n44278,
         n44279, n44280, n44281, n44282, n44283, n44284, n44285, n44286,
         n44287, n44288, n44289, n44290, n44291, n44292, n44293, n44294,
         n44295, n44296, n44297, n44298, n44299, n44300, n44301, n44302,
         n44303, n44304, n44305, n44306, n44307, n44308, n44309, n44310,
         n44311, n44312, n44313, n44314, n44315, n44316, n44317, n44318,
         n44319, n44320, n44321, n44322, n44323, n44324, n44325, n44326,
         n44327, n44328, n44329, n44330, n44331, n44332, n44333, n44334,
         n44335, n44336, n44337, n44338, n44339, n44340, n44341, n44342,
         n44343, n44344, n44345, n44346, n44347, n44348, n44349, n44350,
         n44351, n44352, n44353, n44354, n44355, n44356, n44357, n44358,
         n44359, n44360, n44361, n44362, n44363, n44364, n44365, n44366,
         n44367, n44368, n44369, n44370, n44371, n44372, n44373, n44374,
         n44375, n44376, n44377, n44378, n44379, n44380, n44381, n44382,
         n44383, n44384, n44385, n44386, n44387, n44388, n44389, n44390,
         n44391, n44392, n44393, n44394, n44395, n44396, n44397, n44398,
         n44399, n44400, n44401, n44402, n44403, n44404, n44405, n44406,
         n44407, n44408, n44409, n44410, n44411, n44412, n44413, n44414,
         n44415, n44416, n44417, n44418, n44419, n44420, n44421, n44422,
         n44423, n44424, n44425, n44426, n44427, n44428, n44429, n44430,
         n44431, n44432, n44433, n44434, n44435, n44436, n44437, n44438,
         n44439, n44440, n44441, n44442, n44443, n44444, n44445, n44446,
         n44447, n44448, n44449, n44450, n44451, n44452, n44453, n44454,
         n44455, n44456, n44457, n44458, n44459, n44460, n44461, n44462,
         n44463, n44464, n44465, n44466, n44467, n44468, n44469, n44470,
         n44471, n44472, n44473, n44474, n44475, n44476, n44477, n44478,
         n44479, n44480, n44481, n44482, n44483, n44484, n44485, n44486,
         n44487, n44488, n44489, n44490, n44491, n44492, n44493, n44494,
         n44495, n44496, n44497, n44498, n44499, n44500, n44501, n44502,
         n44503, n44504, n44505, n44506, n44507, n44508, n44509, n44510,
         n44511, n44512, n44513, n44514, n44515, n44516, n44517, n44518,
         n44519, n44520, n44521, n44522, n44523, n44524, n44525, n44526,
         n44527, n44528, n44529, n44530, n44531, n44532, n44533, n44534,
         n44535, n44536, n44537, n44538, n44539, n44540, n44541, n44542,
         n44543, n44544, n44545, n44546, n44547, n44548, n44549, n44550,
         n44551, n44552, n44553, n44554, n44555, n44556, n44557, n44558,
         n44559, n44560, n44561, n44562, n44563, n44564, n44565, n44566,
         n44567, n44568, n44569, n44570, n44571, n44572, n44573, n44574,
         n44575, n44576, n44577, n44578, n44579, n44580, n44581, n44582,
         n44583, n44584, n44585, n44586, n44587, n44588, n44589, n44590,
         n44591, n44592, n44593, n44594, n44595, n44596, n44597, n44598,
         n44599, n44600, n44601, n44602, n44603, n44604, n44605, n44606,
         n44607, n44608, n44609, n44610, n44611, n44612, n44613, n44614,
         n44615, n44616, n44617, n44618, n44619, n44620, n44621, n44622,
         n44623, n44624, n44625, n44626, n44627, n44628, n44629, n44630,
         n44631, n44632, n44633, n44634, n44635, n44636, n44637, n44638,
         n44639, n44640, n44641, n44642, n44643, n44644, n44645, n44646,
         n44647, n44648, n44649, n44650, n44651, n44652, n44653, n44654,
         n44655, n44656, n44657, n44658, n44659, n44660, n44661, n44662,
         n44663, n44664, n44665, n44666, n44667, n44668, n44669, n44670,
         n44671, n44672, n44673, n44674, n44675, n44676, n44677, n44678,
         n44679, n44680, n44681, n44682, n44683, n44684, n44685, n44686,
         n44687, n44688, n44689, n44690, n44691, n44692, n44693, n44694,
         n44695, n44696, n44697, n44698, n44699, n44700, n44701, n44702,
         n44703, n44704, n44705, n44706, n44707, n44708, n44709, n44710,
         n44711, n44712, n44713, n44714, n44715, n44716, n44717, n44718,
         n44719, n44720, n44721, n44722, n44723, n44724, n44725, n44726,
         n44727, n44728, n44729, n44730, n44731, n44732, n44733, n44734,
         n44735, n44736, n44737, n44738, n44739, n44740, n44741, n44742,
         n44743, n44744, n44745, n44746, n44747, n44748, n44749, n44750,
         n44751, n44752, n44753, n44754, n44755, n44756, n44757, n44758,
         n44759, n44760, n44761, n44762, n44763, n44764, n44765, n44766,
         n44767, n44768, n44769, n44770, n44771, n44772, n44773, n44774,
         n44775, n44776, n44777, n44778, n44779, n44780, n44781, n44782,
         n44783, n44784, n44785, n44786, n44787, n44788, n44789, n44790,
         n44791, n44792, n44793, n44794, n44795, n44796, n44797, n44798,
         n44799, n44800, n44801, n44802, n44803, n44804, n44805, n44806,
         n44807, n44808, n44809, n44810, n44811, n44812, n44813, n44814,
         n44815, n44816, n44817, n44818, n44819, n44820, n44821, n44822,
         n44823, n44824, n44825, n44826, n44827, n44828, n44829, n44830,
         n44831, n44832, n44833, n44834, n44835, n44836, n44837, n44838,
         n44839, n44840, n44841, n44842, n44843, n44844, n44845, n44846,
         n44847, n44848, n44849, n44850, n44851, n44852, n44853, n44854,
         n44855, n44856, n44857, n44858, n44859, n44860, n44861, n44862,
         n44863, n44864, n44865, n44866, n44867, n44868, n44869, n44870,
         n44871, n44872, n44873, n44874, n44875, n44876, n44877, n44878,
         n44879, n44880, n44881, n44882, n44883, n44884, n44885, n44886,
         n44887, n44888, n44889, n44890, n44891, n44892, n44893, n44894,
         n44895, n44896, n44897, n44898, n44899, n44900, n44901, n44902,
         n44903, n44904, n44905, n44906, n44907, n44908, n44909, n44910,
         n44911, n44912, n44913, n44914, n44915, n44916, n44917, n44918,
         n44919, n44920, n44921, n44922, n44923, n44924, n44925, n44926,
         n44927, n44928, n44929, n44930, n44931, n44932, n44933, n44934,
         n44935, n44936, n44937, n44938, n44939, n44940, n44941, n44942,
         n44943, n44944, n44945, n44946, n44947, n44948, n44949, n44950,
         n44951, n44952, n44953, n44954, n44955, n44956, n44957, n44958,
         n44959, n44960, n44961, n44962, n44963, n44964, n44965, n44966,
         n44967, n44968, n44969, n44970, n44971, n44972, n44973, n44974,
         n44975, n44976, n44977, n44978, n44979, n44980, n44981, n44982,
         n44983, n44984, n44985, n44986, n44987, n44988, n44989, n44990,
         n44991, n44992, n44993, n44994, n44995, n44996, n44997, n44998,
         n44999, n45000, n45001, n45002, n45003, n45004, n45005, n45006,
         n45007, n45008, n45009, n45010, n45011, n45012, n45013, n45014,
         n45015, n45016, n45017, n45018, n45019, n45020, n45021, n45022,
         n45023, n45024, n45025, n45026, n45027, n45028, n45029, n45030,
         n45031, n45032, n45033, n45034, n45035, n45036, n45037, n45038,
         n45039, n45040, n45041, n45042, n45043, n45044, n45045, n45046,
         n45047, n45048, n45049, n45050, n45051, n45052, n45053, n45054,
         n45055, n45056, n45057, n45058, n45059, n45060, n45061, n45062,
         n45063, n45064, n45065, n45066, n45067, n45068, n45069, n45070,
         n45071, n45072, n45073, n45074, n45075, n45076, n45077, n45078,
         n45079, n45080, n45081, n45082, n45083, n45084, n45085, n45086,
         n45087, n45088, n45089, n45090, n45091, n45092, n45093, n45094,
         n45095, n45096, n45097, n45098, n45099, n45100, n45101, n45102,
         n45103, n45104, n45105, n45106, n45107, n45108, n45109, n45110,
         n45111, n45112, n45113, n45114, n45115, n45116, n45117, n45118,
         n45119, n45120, n45121, n45122, n45123, n45124, n45125, n45126,
         n45127, n45128, n45129, n45130, n45131, n45132, n45133, n45134,
         n45135, n45136, n45137, n45138, n45139, n45140, n45141, n45142,
         n45143, n45144, n45145, n45146, n45147, n45148, n45149, n45150,
         n45151, n45152, n45153, n45154, n45155, n45156, n45157, n45158,
         n45159, n45160, n45161, n45162, n45163, n45164, n45165, n45166,
         n45167, n45168, n45169, n45170, n45171, n45172, n45173, n45174,
         n45175, n45176, n45177, n45178, n45179, n45180, n45181, n45182,
         n45183, n45184, n45185, n45186, n45187, n45188, n45189, n45190,
         n45191, n45192, n45193, n45194, n45195, n45196, n45197, n45198,
         n45199, n45200, n45201, n45202, n45203, n45204, n45205, n45206,
         n45207, n45208, n45209, n45210, n45211, n45212, n45213, n45214,
         n45215, n45216, n45217, n45218, n45219, n45220, n45221, n45222,
         n45223, n45224, n45225, n45226, n45227, n45228, n45229, n45230,
         n45231, n45232, n45233, n45234, n45235, n45236, n45237, n45238,
         n45239, n45240, n45241, n45242, n45243, n45244, n45245, n45246,
         n45247, n45248, n45249, n45250, n45251, n45252, n45253, n45254,
         n45255, n45256, n45257, n45258, n45259, n45260, n45261, n45262,
         n45263, n45264, n45265, n45266, n45267, n45268, n45269, n45270,
         n45271, n45272, n45273, n45274, n45275, n45276, n45277, n45278,
         n45279, n45280, n45281, n45282, n45283, n45284, n45285, n45286,
         n45287, n45288, n45289, n45290, n45291, n45292, n45293, n45294,
         n45295, n45296, n45297, n45298, n45299, n45300, n45301, n45302,
         n45303, n45304, n45305, n45306, n45307, n45308, n45309, n45310,
         n45311, n45312, n45313, n45314, n45315, n45316, n45317, n45318,
         n45319, n45320, n45321, n45322, n45323, n45324, n45325, n45326,
         n45327, n45328, n45329, n45330, n45331, n45332, n45333, n45334,
         n45335, n45336, n45337, n45338, n45339, n45340, n45341, n45342,
         n45343, n45344, n45345, n45346, n45347, n45348, n45349, n45350,
         n45351, n45352, n45353, n45354, n45355, n45356, n45357, n45358,
         n45359, n45360, n45361, n45362, n45363, n45364, n45365, n45366,
         n45367, n45368, n45369, n45370, n45371, n45372, n45373, n45374,
         n45375, n45376, n45377, n45378, n45379, n45380, n45381, n45382,
         n45383, n45384, n45385, n45386, n45387, n45388, n45389, n45390,
         n45391, n45392, n45393, n45394, n45395, n45396, n45397, n45398,
         n45399, n45400, n45401, n45402, n45403, n45404, n45405, n45406,
         n45407, n45408, n45409, n45410, n45411, n45412, n45413, n45414,
         n45415, n45416, n45417, n45418, n45419, n45420, n45421, n45422,
         n45423, n45424, n45425, n45426, n45427, n45428, n45429, n45430,
         n45431, n45432, n45433, n45434, n45435, n45436, n45437, n45438,
         n45439, n45440, n45441, n45442, n45443, n45444, n45445, n45446,
         n45447, n45448, n45449, n45450, n45451, n45452, n45453, n45454,
         n45455, n45456, n45457, n45458, n45459, n45460, n45461, n45462,
         n45463, n45464, n45465, n45466, n45467, n45468, n45469, n45470,
         n45471, n45472, n45473, n45474, n45475, n45476, n45477, n45478,
         n45479, n45480, n45481, n45482, n45483, n45484, n45485, n45486,
         n45487, n45488, n45489, n45490, n45491, n45492, n45493, n45494,
         n45495, n45496, n45497, n45498, n45499, n45500, n45501, n45502,
         n45503, n45504, n45505, n45506, n45507, n45508, n45509, n45510,
         n45511, n45512, n45513, n45514, n45515, n45516, n45517, n45518,
         n45519, n45520, n45521, n45522, n45523, n45524, n45525, n45526,
         n45527, n45528, n45529, n45530, n45531, n45532, n45533, n45534,
         n45535, n45536, n45537, n45538, n45539, n45540, n45541, n45542,
         n45543, n45544, n45545, n45546, n45547, n45548, n45549, n45550,
         n45551, n45552, n45553, n45554, n45555, n45556, n45557, n45558,
         n45559, n45560, n45561, n45562, n45563, n45564, n45565, n45566,
         n45567, n45568, n45569, n45570, n45571, n45572, n45573, n45574,
         n45575, n45576, n45577, n45578, n45579, n45580, n45581, n45582,
         n45583, n45584, n45585, n45586, n45587, n45588, n45589, n45590,
         n45591, n45592, n45593, n45594, n45595, n45596, n45597, n45598,
         n45599, n45600, n45601, n45602, n45603, n45604, n45605, n45606,
         n45607, n45608, n45609, n45610, n45611, n45612, n45613, n45614,
         n45615, n45616, n45617, n45618, n45619, n45620, n45621, n45622,
         n45623, n45624, n45625, n45626, n45627, n45628, n45629, n45630,
         n45631, n45632, n45633, n45634, n45635, n45636, n45637, n45638,
         n45639, n45640, n45641, n45642, n45643, n45644, n45645, n45646,
         n45647, n45648, n45649, n45650, n45651, n45652, n45653, n45654,
         n45655, n45656, n45657, n45658, n45659, n45660, n45661, n45662,
         n45663, n45664, n45665, n45666, n45667, n45668, n45669, n45670,
         n45671, n45672, n45673, n45674, n45675, n45676, n45677, n45678,
         n45679, n45680, n45681, n45682, n45683, n45684, n45685, n45686,
         n45687, n45688, n45689, n45690, n45691, n45692, n45693, n45694,
         n45695, n45696, n45697, n45698, n45699, n45700, n45701, n45702,
         n45703, n45704, n45705, n45706, n45707, n45708, n45709, n45710,
         n45711, n45712, n45713, n45714, n45715, n45716, n45717, n45718,
         n45719, n45720, n45721, n45722, n45723, n45724, n45725, n45726,
         n45727, n45728, n45729, n45730, n45731, n45732, n45733, n45734,
         n45735, n45736, n45737, n45738, n45739, n45740, n45741, n45742,
         n45743, n45744, n45745, n45746, n45747, n45748, n45749, n45750,
         n45751, n45752, n45753, n45754, n45755, n45756, n45757, n45758,
         n45759, n45760, n45761, n45762, n45763, n45764, n45765, n45766,
         n45767, n45768, n45769, n45770, n45771, n45772, n45773, n45774,
         n45775, n45776, n45777, n45778, n45779, n45780, n45781, n45782,
         n45783, n45784, n45785, n45786, n45787, n45788, n45789, n45790,
         n45791, n45792, n45793, n45794, n45795, n45796, n45797, n45798,
         n45799, n45800, n45801, n45802, n45803, n45804, n45805, n45806,
         n45807, n45808, n45809, n45810, n45811, n45812, n45813, n45814,
         n45815, n45816, n45817, n45818, n45819, n45820, n45821, n45822,
         n45823, n45824, n45825, n45826, n45827, n45828, n45829, n45830,
         n45831, n45832, n45833, n45834, n45835, n45836, n45837, n45838,
         n45839, n45840, n45841, n45842, n45843, n45844, n45845, n45846,
         n45847, n45848, n45849, n45850, n45851, n45852, n45853, n45854,
         n45855, n45856, n45857, n45858, n45859, n45860, n45861, n45862,
         n45863, n45864, n45865, n45866, n45867, n45868, n45869, n45870,
         n45871, n45872, n45873, n45874, n45875, n45876, n45877, n45878,
         n45879, n45880, n45881, n45882, n45883, n45884, n45885, n45886,
         n45887, n45888, n45889, n45890, n45891, n45892, n45893, n45894,
         n45895, n45896, n45897, n45898, n45899, n45900, n45901, n45902,
         n45903, n45904, n45905, n45906, n45907, n45908, n45909, n45910,
         n45911, n45912, n45913, n45914, n45915, n45916, n45917, n45918,
         n45919, n45920, n45921, n45922, n45923, n45924, n45925, n45926,
         n45927, n45928, n45929, n45930, n45931, n45932, n45933, n45934,
         n45935, n45936, n45937, n45938, n45939, n45940, n45941, n45942,
         n45943, n45944, n45945, n45946, n45947, n45948, n45949, n45950,
         n45951, n45952, n45953, n45954, n45955, n45956, n45957, n45958,
         n45959, n45960, n45961, n45962, n45963, n45964, n45965, n45966,
         n45967, n45968, n45969, n45970, n45971, n45972, n45973, n45974,
         n45975, n45976, n45977, n45978, n45979, n45980, n45981, n45982,
         n45983, n45984, n45985, n45986, n45987, n45988, n45989, n45990,
         n45991, n45992, n45993, n45994, n45995, n45996, n45997, n45998,
         n45999, n46000, n46001, n46002, n46003, n46004, n46005, n46006,
         n46007, n46008, n46009, n46010, n46011, n46012, n46013, n46014,
         n46015, n46016, n46017, n46018, n46019, n46020, n46021, n46022,
         n46023, n46024, n46025, n46026, n46027, n46028, n46029, n46030,
         n46031, n46032, n46033, n46034, n46035, n46036, n46037, n46038,
         n46039, n46040, n46041, n46042, n46043, n46044, n46045, n46046,
         n46047, n46048, n46049, n46050, n46051, n46052, n46053, n46054,
         n46055, n46056, n46057, n46058, n46059, n46060, n46061, n46062,
         n46063, n46064, n46065, n46066, n46067, n46068, n46069, n46070,
         n46071, n46072, n46073, n46074, n46075, n46076, n46077, n46078,
         n46079, n46080, n46081, n46082, n46083, n46084, n46085, n46086,
         n46087, n46088, n46089, n46090, n46091, n46092, n46093, n46094,
         n46095, n46096, n46097, n46098, n46099, n46100, n46101, n46102,
         n46103, n46104, n46105, n46106, n46107, n46108, n46109, n46110,
         n46111, n46112, n46113, n46114, n46115, n46116, n46117, n46118,
         n46119, n46120, n46121, n46122, n46123, n46124, n46125, n46126,
         n46127, n46128, n46129, n46130, n46131, n46132, n46133, n46134,
         n46135, n46136, n46137, n46138, n46139, n46140, n46141, n46142,
         n46143, n46144, n46145, n46146, n46147, n46148, n46149, n46150,
         n46151, n46152, n46153, n46154, n46155, n46156, n46157, n46158,
         n46159, n46160, n46161, n46162, n46163, n46164, n46165, n46166,
         n46167, n46168, n46169, n46170, n46171, n46172, n46173, n46174,
         n46175, n46176, n46177, n46178, n46179, n46180, n46181, n46182,
         n46183, n46184, n46185, n46186, n46187, n46188, n46189, n46190,
         n46191, n46192, n46193, n46194, n46195, \shifter_0/n12761 ,
         \shifter_0/n12760 , \shifter_0/n12757 , \shifter_0/n12756 ,
         \shifter_0/n12753 , \shifter_0/n12752 , \shifter_0/n12749 ,
         \shifter_0/n12748 , \shifter_0/n12745 , \shifter_0/n12744 ,
         \shifter_0/n12741 , \shifter_0/n12740 , \shifter_0/n12737 ,
         \shifter_0/n12736 , \shifter_0/n12733 , \shifter_0/n12732 ,
         \shifter_0/n12729 , \shifter_0/n12728 , \shifter_0/n12725 ,
         \shifter_0/n12724 , \shifter_0/n12721 , \shifter_0/n12720 ,
         \shifter_0/n12717 , \shifter_0/n12716 , \shifter_0/n12713 ,
         \shifter_0/n12712 , \shifter_0/n12709 , \shifter_0/n12708 ,
         \shifter_0/n12705 , \shifter_0/n12704 , \shifter_0/n12701 ,
         \shifter_0/n12700 , \shifter_0/n12697 , \shifter_0/n12696 ,
         \shifter_0/n12693 , \shifter_0/n12692 , \shifter_0/n12689 ,
         \shifter_0/n12688 , \shifter_0/n12685 , \shifter_0/n12684 ,
         \shifter_0/n12681 , \shifter_0/n12680 , \shifter_0/n12677 ,
         \shifter_0/n12676 , \shifter_0/n12673 , \shifter_0/n12672 ,
         \shifter_0/n12669 , \shifter_0/n12668 , \shifter_0/n12665 ,
         \shifter_0/n12664 , \shifter_0/n12661 , \shifter_0/n12660 ,
         \shifter_0/n12657 , \shifter_0/n12656 , \shifter_0/n12653 ,
         \shifter_0/n12652 , \shifter_0/n12649 , \shifter_0/n12648 ,
         \shifter_0/n12645 , \shifter_0/n12644 , \shifter_0/n12641 ,
         \shifter_0/n12640 , \shifter_0/n12637 , \shifter_0/n12636 ,
         \shifter_0/n12633 , \shifter_0/n12632 , \shifter_0/n12629 ,
         \shifter_0/n12628 , \shifter_0/n12625 , \shifter_0/n12624 ,
         \shifter_0/n12621 , \shifter_0/n12620 , \shifter_0/n12617 ,
         \shifter_0/n12616 , \shifter_0/n12613 , \shifter_0/n12612 ,
         \shifter_0/n12609 , \shifter_0/n12608 , \shifter_0/n12605 ,
         \shifter_0/n12604 , \shifter_0/n12601 , \shifter_0/n12600 ,
         \shifter_0/n12597 , \shifter_0/n12596 , \shifter_0/n12593 ,
         \shifter_0/n12592 , \shifter_0/n12589 , \shifter_0/n12588 ,
         \shifter_0/n12585 , \shifter_0/n12584 , \shifter_0/n12581 ,
         \shifter_0/n12580 , \shifter_0/n12577 , \shifter_0/n12576 ,
         \shifter_0/n12573 , \shifter_0/n12572 , \shifter_0/n12569 ,
         \shifter_0/n12568 , \shifter_0/n12565 , \shifter_0/n12564 ,
         \shifter_0/n12561 , \shifter_0/n12560 , \shifter_0/n12557 ,
         \shifter_0/n12556 , \shifter_0/n12553 , \shifter_0/n12552 ,
         \shifter_0/n12549 , \shifter_0/n12548 , \shifter_0/n12545 ,
         \shifter_0/n12544 , \shifter_0/n12541 , \shifter_0/n12540 ,
         \shifter_0/n12537 , \shifter_0/n12536 , \shifter_0/n12533 ,
         \shifter_0/n12532 , \shifter_0/n12529 , \shifter_0/n12528 ,
         \shifter_0/n12525 , \shifter_0/n12524 , \shifter_0/n12521 ,
         \shifter_0/n12520 , \shifter_0/n12517 , \shifter_0/n12516 ,
         \shifter_0/n12513 , \shifter_0/n12512 , \shifter_0/n12509 ,
         \shifter_0/n12508 , \shifter_0/n12505 , \shifter_0/n12504 ,
         \shifter_0/n12501 , \shifter_0/n12500 , \shifter_0/n12497 ,
         \shifter_0/n12496 , \shifter_0/n12493 , \shifter_0/n12492 ,
         \shifter_0/n12489 , \shifter_0/n12488 , \shifter_0/n12485 ,
         \shifter_0/n12484 , \shifter_0/n12481 , \shifter_0/n12480 ,
         \shifter_0/n12477 , \shifter_0/n12476 , \shifter_0/n12473 ,
         \shifter_0/n12472 , \shifter_0/n12469 , \shifter_0/n12468 ,
         \shifter_0/n12465 , \shifter_0/n12464 , \shifter_0/n12461 ,
         \shifter_0/n12460 , \shifter_0/n12457 , \shifter_0/n12456 ,
         \shifter_0/n12453 , \shifter_0/n12452 , \shifter_0/n12449 ,
         \shifter_0/n12448 , \shifter_0/n12445 , \shifter_0/n12444 ,
         \shifter_0/n12441 , \shifter_0/n12440 , \shifter_0/n12437 ,
         \shifter_0/n12436 , \shifter_0/n12433 , \shifter_0/n12432 ,
         \shifter_0/n12429 , \shifter_0/n12428 , \shifter_0/n12425 ,
         \shifter_0/n12424 , \shifter_0/n12421 , \shifter_0/n12420 ,
         \shifter_0/n12417 , \shifter_0/n12416 , \shifter_0/n12413 ,
         \shifter_0/n12412 , \shifter_0/n12409 , \shifter_0/n12408 ,
         \shifter_0/n12405 , \shifter_0/n12404 , \shifter_0/n12401 ,
         \shifter_0/n12400 , \shifter_0/n12397 , \shifter_0/n12396 ,
         \shifter_0/n12393 , \shifter_0/n12392 , \shifter_0/n12389 ,
         \shifter_0/n12388 , \shifter_0/n12385 , \shifter_0/n12384 ,
         \shifter_0/n12381 , \shifter_0/n12380 , \shifter_0/n12377 ,
         \shifter_0/n12376 , \shifter_0/n12373 , \shifter_0/n12372 ,
         \shifter_0/n12369 , \shifter_0/n12368 , \shifter_0/n12365 ,
         \shifter_0/n12364 , \shifter_0/n12361 , \shifter_0/n12360 ,
         \shifter_0/n12357 , \shifter_0/n12356 , \shifter_0/n12353 ,
         \shifter_0/n12352 , \shifter_0/n12349 , \shifter_0/n12348 ,
         \shifter_0/n12345 , \shifter_0/n12344 , \shifter_0/n12341 ,
         \shifter_0/n12340 , \shifter_0/n12337 , \shifter_0/n12336 ,
         \shifter_0/n12333 , \shifter_0/n12332 , \shifter_0/n12329 ,
         \shifter_0/n12328 , \shifter_0/n12325 , \shifter_0/n12324 ,
         \shifter_0/n12321 , \shifter_0/n12320 , \shifter_0/n12317 ,
         \shifter_0/n12316 , \shifter_0/n12313 , \shifter_0/n12312 ,
         \shifter_0/n12309 , \shifter_0/n12308 , \shifter_0/n12305 ,
         \shifter_0/n12304 , \shifter_0/n12301 , \shifter_0/n12300 ,
         \shifter_0/n12297 , \shifter_0/n12296 , \shifter_0/n12293 ,
         \shifter_0/n12292 , \shifter_0/n12289 , \shifter_0/n12288 ,
         \shifter_0/n12285 , \shifter_0/n12284 , \shifter_0/n12281 ,
         \shifter_0/n12280 , \shifter_0/n12277 , \shifter_0/n12276 ,
         \shifter_0/n12273 , \shifter_0/n12272 , \shifter_0/n12269 ,
         \shifter_0/n12268 , \shifter_0/n12265 , \shifter_0/n12264 ,
         \shifter_0/n12261 , \shifter_0/n12260 , \shifter_0/n12257 ,
         \shifter_0/n12256 , \shifter_0/n12253 , \shifter_0/n12252 ,
         \shifter_0/n12249 , \shifter_0/n12248 , \shifter_0/n12245 ,
         \shifter_0/n12244 , \shifter_0/n12241 , \shifter_0/n12240 ,
         \shifter_0/n12237 , \shifter_0/n12236 , \shifter_0/n12233 ,
         \shifter_0/n12232 , \shifter_0/n12229 , \shifter_0/n12228 ,
         \shifter_0/n12225 , \shifter_0/n12224 , \shifter_0/n12221 ,
         \shifter_0/n12220 , \shifter_0/n12217 , \shifter_0/n12216 ,
         \shifter_0/n12213 , \shifter_0/n12212 , \shifter_0/n12209 ,
         \shifter_0/n12208 , \shifter_0/n12205 , \shifter_0/n12204 ,
         \shifter_0/n12201 , \shifter_0/n12200 , \shifter_0/n12197 ,
         \shifter_0/n12196 , \shifter_0/n12193 , \shifter_0/n12192 ,
         \shifter_0/n12189 , \shifter_0/n12188 , \shifter_0/n12185 ,
         \shifter_0/n12184 , \shifter_0/n12181 , \shifter_0/n12180 ,
         \shifter_0/n12177 , \shifter_0/n12176 , \shifter_0/n12173 ,
         \shifter_0/n12172 , \shifter_0/n12169 , \shifter_0/n12168 ,
         \shifter_0/n12165 , \shifter_0/n12164 , \shifter_0/n12161 ,
         \shifter_0/n12160 , \shifter_0/n12157 , \shifter_0/n12156 ,
         \shifter_0/n12153 , \shifter_0/n12152 , \shifter_0/n12149 ,
         \shifter_0/n12148 , \shifter_0/n12145 , \shifter_0/n12144 ,
         \shifter_0/n12141 , \shifter_0/n12140 , \shifter_0/n12137 ,
         \shifter_0/n12136 , \shifter_0/n12133 , \shifter_0/n12132 ,
         \shifter_0/n12129 , \shifter_0/n12128 , \shifter_0/n12125 ,
         \shifter_0/n12124 , \shifter_0/n12121 , \shifter_0/n12120 ,
         \shifter_0/n12117 , \shifter_0/n12116 , \shifter_0/n12113 ,
         \shifter_0/n12112 , \shifter_0/n12109 , \shifter_0/n12108 ,
         \shifter_0/n12105 , \shifter_0/n12104 , \shifter_0/n12101 ,
         \shifter_0/n12100 , \shifter_0/n12097 , \shifter_0/n12096 ,
         \shifter_0/n12093 , \shifter_0/n12092 , \shifter_0/n12089 ,
         \shifter_0/n12088 , \shifter_0/n12085 , \shifter_0/n12084 ,
         \shifter_0/n12081 , \shifter_0/n12080 , \shifter_0/n12077 ,
         \shifter_0/n12076 , \shifter_0/n12073 , \shifter_0/n12072 ,
         \shifter_0/n12069 , \shifter_0/n12068 , \shifter_0/n12065 ,
         \shifter_0/n12064 , \shifter_0/n12061 , \shifter_0/n12060 ,
         \shifter_0/n12057 , \shifter_0/n12056 , \shifter_0/n12053 ,
         \shifter_0/n12052 , \shifter_0/n12049 , \shifter_0/n12048 ,
         \shifter_0/n12045 , \shifter_0/n12044 , \shifter_0/n12041 ,
         \shifter_0/n12040 , \shifter_0/n12037 , \shifter_0/n12036 ,
         \shifter_0/n12033 , \shifter_0/n12032 , \shifter_0/n12029 ,
         \shifter_0/n12028 , \shifter_0/n12025 , \shifter_0/n12024 ,
         \shifter_0/n12021 , \shifter_0/n12020 , \shifter_0/n12017 ,
         \shifter_0/n12016 , \shifter_0/n12013 , \shifter_0/n12012 ,
         \shifter_0/n12009 , \shifter_0/n12008 , \shifter_0/n12005 ,
         \shifter_0/n12004 , \shifter_0/n12001 , \shifter_0/n12000 ,
         \shifter_0/n11997 , \shifter_0/n11996 , \shifter_0/n11993 ,
         \shifter_0/n11992 , \shifter_0/n11989 , \shifter_0/n11988 ,
         \shifter_0/n11985 , \shifter_0/n11984 , \shifter_0/n11981 ,
         \shifter_0/n11980 , \shifter_0/n11977 , \shifter_0/n11976 ,
         \shifter_0/n11973 , \shifter_0/n11972 , \shifter_0/n11969 ,
         \shifter_0/n11968 , \shifter_0/n11965 , \shifter_0/n11964 ,
         \shifter_0/n11961 , \shifter_0/n11960 , \shifter_0/n11957 ,
         \shifter_0/n11956 , \shifter_0/n11953 , \shifter_0/n11952 ,
         \shifter_0/n11949 , \shifter_0/n11948 , \shifter_0/n11945 ,
         \shifter_0/n11944 , \shifter_0/n11941 , \shifter_0/n11940 ,
         \shifter_0/n11937 , \shifter_0/n11936 , \shifter_0/n11933 ,
         \shifter_0/n11932 , \shifter_0/n11929 , \shifter_0/n11928 ,
         \shifter_0/n11925 , \shifter_0/n11924 , \shifter_0/n11921 ,
         \shifter_0/n11920 , \shifter_0/n11917 , \shifter_0/n11916 ,
         \shifter_0/n11913 , \shifter_0/n11912 , \shifter_0/n11909 ,
         \shifter_0/n11908 , \shifter_0/n11905 , \shifter_0/n11904 ,
         \shifter_0/n11901 , \shifter_0/n11900 , \shifter_0/n11897 ,
         \shifter_0/n11896 , \shifter_0/n11893 , \shifter_0/n11892 ,
         \shifter_0/n11889 , \shifter_0/n11888 , \shifter_0/n11884 ,
         \shifter_0/n11880 , \shifter_0/n11876 , \shifter_0/n11872 ,
         \shifter_0/n11868 , \shifter_0/n11864 , \shifter_0/n11860 ,
         \shifter_0/n11856 , \shifter_0/n11852 , \shifter_0/n11848 ,
         \shifter_0/n11844 , \shifter_0/n11840 , \shifter_0/n11836 ,
         \shifter_0/n11832 , \shifter_0/n11828 , \shifter_0/n11824 ,
         \shifter_0/n11820 , \shifter_0/n11816 , \shifter_0/n11812 ,
         \shifter_0/n11808 , \shifter_0/n11804 , \shifter_0/n11800 ,
         \shifter_0/n11796 , \shifter_0/n11792 , \shifter_0/n11788 ,
         \shifter_0/n11784 , \shifter_0/n11780 , \shifter_0/n11776 ,
         \shifter_0/n11772 , \shifter_0/n11768 , \shifter_0/n11764 ,
         \shifter_0/n11760 , \shifter_0/n11756 , \shifter_0/n11752 ,
         \shifter_0/n11748 , \shifter_0/n11744 , \shifter_0/n11740 ,
         \shifter_0/n11736 , \shifter_0/n11732 , \shifter_0/n11728 ,
         \shifter_0/n11725 , \shifter_0/n11724 , \shifter_0/n11721 ,
         \shifter_0/n11720 , \shifter_0/n11717 , \shifter_0/n11716 ,
         \shifter_0/n11713 , \shifter_0/n11712 , \shifter_0/n11709 ,
         \shifter_0/n11708 , \shifter_0/n11705 , \shifter_0/n11704 ,
         \shifter_0/n11701 , \shifter_0/n11700 , \shifter_0/n11697 ,
         \shifter_0/n11696 , \shifter_0/n11693 , \shifter_0/n11692 ,
         \shifter_0/n11689 , \shifter_0/n11688 , \shifter_0/n11685 ,
         \shifter_0/n11684 , \shifter_0/n11681 , \shifter_0/n11680 ,
         \shifter_0/n11677 , \shifter_0/n11676 , \shifter_0/n11673 ,
         \shifter_0/n11672 , \shifter_0/n11669 , \shifter_0/n11668 ,
         \shifter_0/n11665 , \shifter_0/n11664 , \shifter_0/n11661 ,
         \shifter_0/n11660 , \shifter_0/n11657 , \shifter_0/n11656 ,
         \shifter_0/n11653 , \shifter_0/n11652 , \shifter_0/n11649 ,
         \shifter_0/n11648 , \shifter_0/n11645 , \shifter_0/n11644 ,
         \shifter_0/n11641 , \shifter_0/n11640 , \shifter_0/n11637 ,
         \shifter_0/n11636 , \shifter_0/n11633 , \shifter_0/n11632 ,
         \shifter_0/n11629 , \shifter_0/n11628 , \shifter_0/n11625 ,
         \shifter_0/n11624 , \shifter_0/n11621 , \shifter_0/n11620 ,
         \shifter_0/n11617 , \shifter_0/n11616 , \shifter_0/n11613 ,
         \shifter_0/n11612 , \shifter_0/n11609 , \shifter_0/n11608 ,
         \shifter_0/n11605 , \shifter_0/n11604 , \shifter_0/n11601 ,
         \shifter_0/n11600 , \shifter_0/n11597 , \shifter_0/n11596 ,
         \shifter_0/n11593 , \shifter_0/n11592 , \shifter_0/n11589 ,
         \shifter_0/n11588 , \shifter_0/n11585 , \shifter_0/n11584 ,
         \shifter_0/n11581 , \shifter_0/n11580 , \shifter_0/n11577 ,
         \shifter_0/n11576 , \shifter_0/n11573 , \shifter_0/n11572 ,
         \shifter_0/n11569 , \shifter_0/n11568 , \shifter_0/n11565 ,
         \shifter_0/n11564 , \shifter_0/n11561 , \shifter_0/n11560 ,
         \shifter_0/n11557 , \shifter_0/n11556 , \shifter_0/n11553 ,
         \shifter_0/n11552 , \shifter_0/n11549 , \shifter_0/n11548 ,
         \shifter_0/n11545 , \shifter_0/n11544 , \shifter_0/n11541 ,
         \shifter_0/n11540 , \shifter_0/n11537 , \shifter_0/n11536 ,
         \shifter_0/n11533 , \shifter_0/n11532 , \shifter_0/n11529 ,
         \shifter_0/n11528 , \shifter_0/n11525 , \shifter_0/n11524 ,
         \shifter_0/n11521 , \shifter_0/n11520 , \shifter_0/n11517 ,
         \shifter_0/n11516 , \shifter_0/n11513 , \shifter_0/n11512 ,
         \shifter_0/n11509 , \shifter_0/n11508 , \shifter_0/n11505 ,
         \shifter_0/n11504 , \shifter_0/n11501 , \shifter_0/n11500 ,
         \shifter_0/n11497 , \shifter_0/n11496 , \shifter_0/n11493 ,
         \shifter_0/n11492 , \shifter_0/n11489 , \shifter_0/n11488 ,
         \shifter_0/n11485 , \shifter_0/n11484 , \shifter_0/n11481 ,
         \shifter_0/n11480 , \shifter_0/n11477 , \shifter_0/n11476 ,
         \shifter_0/n11473 , \shifter_0/n11472 , \shifter_0/n11469 ,
         \shifter_0/n11468 , \shifter_0/n11465 , \shifter_0/n11464 ,
         \shifter_0/n11461 , \shifter_0/n11460 , \shifter_0/n11457 ,
         \shifter_0/n11456 , \shifter_0/n11453 , \shifter_0/n11452 ,
         \shifter_0/n11449 , \shifter_0/n11448 , \shifter_0/n11445 ,
         \shifter_0/n11444 , \shifter_0/n11441 , \shifter_0/n11440 ,
         \shifter_0/n11437 , \shifter_0/n11436 , \shifter_0/n11433 ,
         \shifter_0/n11432 , \shifter_0/n11429 , \shifter_0/n11428 ,
         \shifter_0/n11425 , \shifter_0/n11424 , \shifter_0/n11421 ,
         \shifter_0/n11420 , \shifter_0/n11417 , \shifter_0/n11416 ,
         \shifter_0/n11413 , \shifter_0/n11412 , \shifter_0/n11409 ,
         \shifter_0/n11408 , \shifter_0/n11405 , \shifter_0/n11404 ,
         \shifter_0/n11401 , \shifter_0/n11400 , \shifter_0/n11397 ,
         \shifter_0/n11396 , \shifter_0/n11393 , \shifter_0/n11392 ,
         \shifter_0/n11389 , \shifter_0/n11388 , \shifter_0/n11385 ,
         \shifter_0/n11384 , \shifter_0/n11381 , \shifter_0/n11380 ,
         \shifter_0/n11377 , \shifter_0/n11376 , \shifter_0/n11373 ,
         \shifter_0/n11372 , \shifter_0/n11369 , \shifter_0/n11368 ,
         \shifter_0/n11365 , \shifter_0/n11364 , \shifter_0/n11361 ,
         \shifter_0/n11360 , \shifter_0/n11357 , \shifter_0/n11356 ,
         \shifter_0/n11353 , \shifter_0/n11352 , \shifter_0/n11349 ,
         \shifter_0/n11348 , \shifter_0/n11345 , \shifter_0/n11344 ,
         \shifter_0/n11341 , \shifter_0/n11340 , \shifter_0/n11337 ,
         \shifter_0/n11336 , \shifter_0/n11333 , \shifter_0/n11332 ,
         \shifter_0/n11329 , \shifter_0/n11328 , \shifter_0/n11325 ,
         \shifter_0/n11324 , \shifter_0/n11321 , \shifter_0/n11320 ,
         \shifter_0/n11317 , \shifter_0/n11316 , \shifter_0/n11313 ,
         \shifter_0/n11312 , \shifter_0/n11309 , \shifter_0/n11308 ,
         \shifter_0/n11305 , \shifter_0/n11304 , \shifter_0/n11301 ,
         \shifter_0/n11300 , \shifter_0/n11297 , \shifter_0/n11296 ,
         \shifter_0/n11293 , \shifter_0/n11292 , \shifter_0/n11289 ,
         \shifter_0/n11288 , \shifter_0/n11285 , \shifter_0/n11284 ,
         \shifter_0/n11281 , \shifter_0/n11280 , \shifter_0/n11277 ,
         \shifter_0/n11276 , \shifter_0/n11273 , \shifter_0/n11272 ,
         \shifter_0/n11269 , \shifter_0/n11268 , \shifter_0/n11265 ,
         \shifter_0/n11264 , \shifter_0/n11261 , \shifter_0/n11260 ,
         \shifter_0/n11257 , \shifter_0/n11256 , \shifter_0/n11253 ,
         \shifter_0/n11252 , \shifter_0/n11249 , \shifter_0/n11248 ,
         \shifter_0/n11245 , \shifter_0/n11244 , \shifter_0/n11241 ,
         \shifter_0/n11240 , \shifter_0/n11237 , \shifter_0/n11236 ,
         \shifter_0/n11233 , \shifter_0/n11232 , \shifter_0/n11229 ,
         \shifter_0/n11228 , \shifter_0/n11225 , \shifter_0/n11224 ,
         \shifter_0/n11221 , \shifter_0/n11220 , \shifter_0/n11217 ,
         \shifter_0/n11216 , \shifter_0/n11213 , \shifter_0/n11212 ,
         \shifter_0/n11209 , \shifter_0/n11208 , \shifter_0/n11205 ,
         \shifter_0/n11204 , \shifter_0/n11201 , \shifter_0/n11200 ,
         \shifter_0/n11197 , \shifter_0/n11196 , \shifter_0/n11193 ,
         \shifter_0/n11192 , \shifter_0/n11189 , \shifter_0/n11188 ,
         \shifter_0/n11185 , \shifter_0/n11184 , \shifter_0/n11181 ,
         \shifter_0/n11180 , \shifter_0/n11177 , \shifter_0/n11176 ,
         \shifter_0/n11173 , \shifter_0/n11172 , \shifter_0/n11169 ,
         \shifter_0/n11168 , \shifter_0/n11165 , \shifter_0/n11164 ,
         \shifter_0/n11161 , \shifter_0/n11160 , \shifter_0/n11157 ,
         \shifter_0/n11156 , \shifter_0/n11153 , \shifter_0/n11152 ,
         \shifter_0/n11149 , \shifter_0/n11148 , \shifter_0/n11145 ,
         \shifter_0/n11144 , \shifter_0/n11141 , \shifter_0/n11140 ,
         \shifter_0/n11137 , \shifter_0/n11136 , \shifter_0/n11133 ,
         \shifter_0/n11132 , \shifter_0/n11129 , \shifter_0/n11128 ,
         \shifter_0/n11125 , \shifter_0/n11124 , \shifter_0/n11121 ,
         \shifter_0/n11120 , \shifter_0/n11117 , \shifter_0/n11116 ,
         \shifter_0/n11113 , \shifter_0/n11112 , \shifter_0/n11109 ,
         \shifter_0/n11108 , \shifter_0/n11105 , \shifter_0/n11104 ,
         \shifter_0/n11101 , \shifter_0/n11100 , \shifter_0/n11097 ,
         \shifter_0/n11096 , \shifter_0/n11093 , \shifter_0/n11092 ,
         \shifter_0/n11089 , \shifter_0/n11088 , \shifter_0/n11085 ,
         \shifter_0/n11084 , \shifter_0/n11081 , \shifter_0/n11080 ,
         \shifter_0/n11077 , \shifter_0/n11076 , \shifter_0/n11073 ,
         \shifter_0/n11072 , \shifter_0/n11069 , \shifter_0/n11068 ,
         \shifter_0/n11065 , \shifter_0/n11064 , \shifter_0/n11061 ,
         \shifter_0/n11060 , \shifter_0/n11057 , \shifter_0/n11056 ,
         \shifter_0/n11053 , \shifter_0/n11052 , \shifter_0/n11049 ,
         \shifter_0/n11048 , \shifter_0/n11045 , \shifter_0/n11044 ,
         \shifter_0/n11041 , \shifter_0/n11040 , \shifter_0/n11037 ,
         \shifter_0/n11036 , \shifter_0/n11033 , \shifter_0/n11032 ,
         \shifter_0/n11029 , \shifter_0/n11028 , \shifter_0/n11025 ,
         \shifter_0/n11024 , \shifter_0/n11021 , \shifter_0/n11020 ,
         \shifter_0/n11017 , \shifter_0/n11016 , \shifter_0/n11013 ,
         \shifter_0/n11012 , \shifter_0/n11009 , \shifter_0/n11008 ,
         \shifter_0/n11005 , \shifter_0/n11004 , \shifter_0/n11001 ,
         \shifter_0/n11000 , \shifter_0/n10997 , \shifter_0/n10996 ,
         \shifter_0/n10993 , \shifter_0/n10992 , \shifter_0/n10989 ,
         \shifter_0/n10988 , \shifter_0/n10985 , \shifter_0/n10984 ,
         \shifter_0/n10981 , \shifter_0/n10980 , \shifter_0/n10977 ,
         \shifter_0/n10976 , \shifter_0/n10973 , \shifter_0/n10972 ,
         \shifter_0/n10969 , \shifter_0/n10968 , \shifter_0/n10965 ,
         \shifter_0/n10964 , \shifter_0/n10961 , \shifter_0/n10960 ,
         \shifter_0/n10957 , \shifter_0/n10956 , \shifter_0/n10953 ,
         \shifter_0/n10952 , \shifter_0/n10949 , \shifter_0/n10948 ,
         \shifter_0/n10945 , \shifter_0/n10944 , \shifter_0/n10941 ,
         \shifter_0/n10940 , \shifter_0/n10937 , \shifter_0/n10936 ,
         \shifter_0/n10933 , \shifter_0/n10932 , \shifter_0/n10929 ,
         \shifter_0/n10928 , \shifter_0/n10925 , \shifter_0/n10924 ,
         \shifter_0/n10921 , \shifter_0/n10920 , \shifter_0/n10917 ,
         \shifter_0/n10916 , \shifter_0/n10913 , \shifter_0/n10912 ,
         \shifter_0/n10909 , \shifter_0/n10908 , \shifter_0/n10905 ,
         \shifter_0/n10904 , \shifter_0/n10901 , \shifter_0/n10900 ,
         \shifter_0/n10897 , \shifter_0/n10896 , \shifter_0/n10893 ,
         \shifter_0/n10892 , \shifter_0/n10889 , \shifter_0/n10888 ,
         \shifter_0/n10885 , \shifter_0/n10884 , \shifter_0/n10881 ,
         \shifter_0/n10880 , \shifter_0/n10877 , \shifter_0/n10876 ,
         \shifter_0/n10873 , \shifter_0/n10872 , \shifter_0/n10869 ,
         \shifter_0/n10868 , \shifter_0/n10865 , \shifter_0/n10864 ,
         \shifter_0/n10861 , \shifter_0/n10860 , \shifter_0/n10857 ,
         \shifter_0/n10856 , \shifter_0/n10853 , \shifter_0/n10852 ,
         \shifter_0/n10849 , \shifter_0/n10848 , \shifter_0/n10845 ,
         \shifter_0/n10844 , \shifter_0/n10841 , \shifter_0/n10840 ,
         \shifter_0/n10837 , \shifter_0/n10836 , \shifter_0/n10833 ,
         \shifter_0/n10832 , \shifter_0/n10829 , \shifter_0/n10828 ,
         \shifter_0/n10825 , \shifter_0/n10824 , \shifter_0/n10821 ,
         \shifter_0/n10820 , \shifter_0/n10817 , \shifter_0/n10816 ,
         \shifter_0/n10813 , \shifter_0/n10812 , \shifter_0/n10809 ,
         \shifter_0/n10808 , \shifter_0/n10805 , \shifter_0/n10804 ,
         \shifter_0/n10801 , \shifter_0/n10800 , \shifter_0/n10797 ,
         \shifter_0/n10796 , \shifter_0/n10793 , \shifter_0/n10792 ,
         \shifter_0/n10789 , \shifter_0/n10788 , \shifter_0/n10785 ,
         \shifter_0/n10784 , \shifter_0/n10781 , \shifter_0/n10780 ,
         \shifter_0/n10777 , \shifter_0/n10776 , \shifter_0/n10773 ,
         \shifter_0/n10772 , \shifter_0/n10769 , \shifter_0/n10768 ,
         \shifter_0/n10765 , \shifter_0/n10764 , \shifter_0/n10761 ,
         \shifter_0/n10760 , \shifter_0/n10757 , \shifter_0/n10756 ,
         \shifter_0/n10753 , \shifter_0/n10752 , \shifter_0/n10749 ,
         \shifter_0/n10748 , \shifter_0/n10745 , \shifter_0/n10744 ,
         \shifter_0/n10741 , \shifter_0/n10740 , \shifter_0/n10737 ,
         \shifter_0/n10736 , \shifter_0/n10733 , \shifter_0/n10732 ,
         \shifter_0/n10729 , \shifter_0/n10728 , \shifter_0/n10725 ,
         \shifter_0/n10724 , \shifter_0/n10721 , \shifter_0/n10720 ,
         \shifter_0/n10717 , \shifter_0/n10716 , \shifter_0/n10713 ,
         \shifter_0/n10712 , \shifter_0/n10709 , \shifter_0/n10708 ,
         \shifter_0/n10705 , \shifter_0/n10704 , \shifter_0/n10701 ,
         \shifter_0/n10700 , \shifter_0/n10697 , \shifter_0/n10696 ,
         \shifter_0/n10693 , \shifter_0/n10692 , \shifter_0/n10689 ,
         \shifter_0/n10688 , \shifter_0/n10685 , \shifter_0/n10684 ,
         \shifter_0/n10681 , \shifter_0/n10680 , \shifter_0/n10677 ,
         \shifter_0/n10676 , \shifter_0/n10673 , \shifter_0/n10672 ,
         \shifter_0/n10669 , \shifter_0/n10668 , \shifter_0/n10665 ,
         \shifter_0/n10664 , \shifter_0/n10661 , \shifter_0/n10660 ,
         \shifter_0/n10657 , \shifter_0/n10656 , \shifter_0/n10653 ,
         \shifter_0/n10652 , \shifter_0/n10649 , \shifter_0/n10648 ,
         \shifter_0/n10645 , \shifter_0/n10644 , \shifter_0/n10641 ,
         \shifter_0/n10640 , \shifter_0/n10637 , \shifter_0/n10636 ,
         \shifter_0/n10633 , \shifter_0/n10632 , \shifter_0/n10629 ,
         \shifter_0/n10628 , \shifter_0/n10625 , \shifter_0/n10624 ,
         \shifter_0/n10621 , \shifter_0/n10620 , \shifter_0/n10617 ,
         \shifter_0/n10616 , \shifter_0/n10613 , \shifter_0/n10612 ,
         \shifter_0/n10609 , \shifter_0/n10608 , \shifter_0/n10605 ,
         \shifter_0/n10604 , \shifter_0/n10601 , \shifter_0/n10600 ,
         \shifter_0/n10597 , \shifter_0/n10596 , \shifter_0/n10593 ,
         \shifter_0/n10592 , \shifter_0/n10589 , \shifter_0/n10588 ,
         \shifter_0/n10585 , \shifter_0/n10584 , \shifter_0/n10581 ,
         \shifter_0/n10580 , \shifter_0/n10577 , \shifter_0/n10576 ,
         \shifter_0/n10573 , \shifter_0/n10572 , \shifter_0/n10569 ,
         \shifter_0/n10568 , \shifter_0/n10565 , \shifter_0/n10564 ,
         \shifter_0/n10561 , \shifter_0/n10560 , \shifter_0/n10557 ,
         \shifter_0/n10556 , \shifter_0/n10553 , \shifter_0/n10552 ,
         \shifter_0/n10549 , \shifter_0/n10548 , \shifter_0/n10545 ,
         \shifter_0/n10544 , \shifter_0/n10541 , \shifter_0/n10540 ,
         \shifter_0/n10537 , \shifter_0/n10536 , \shifter_0/n10533 ,
         \shifter_0/n10532 , \shifter_0/n10529 , \shifter_0/n10528 ,
         \shifter_0/n10525 , \shifter_0/n10524 , \shifter_0/n10521 ,
         \shifter_0/n10520 , \shifter_0/n10517 , \shifter_0/n10516 ,
         \shifter_0/n10513 , \shifter_0/n10512 , \shifter_0/n10509 ,
         \shifter_0/n10508 , \shifter_0/n10505 , \shifter_0/n10504 ,
         \shifter_0/n10501 , \shifter_0/n10500 , \shifter_0/n10497 ,
         \shifter_0/n10496 , \shifter_0/n10493 , \shifter_0/n10492 ,
         \shifter_0/n10489 , \shifter_0/n10488 , \shifter_0/n10485 ,
         \shifter_0/n10484 , \shifter_0/n10481 , \shifter_0/n10480 ,
         \shifter_0/n10477 , \shifter_0/n10476 , \shifter_0/n10473 ,
         \shifter_0/n10472 , \shifter_0/n10469 , \shifter_0/n10468 ,
         \shifter_0/n10465 , \shifter_0/n10464 , \shifter_0/n10461 ,
         \shifter_0/n10460 , \shifter_0/n10457 , \shifter_0/n10456 ,
         \shifter_0/n10453 , \shifter_0/n10452 , \shifter_0/n10449 ,
         \shifter_0/n10448 , \shifter_0/n10445 , \shifter_0/n10444 ,
         \shifter_0/n10441 , \shifter_0/n10440 , \shifter_0/n10437 ,
         \shifter_0/n10436 , \shifter_0/n10433 , \shifter_0/n10432 ,
         \shifter_0/n10429 , \shifter_0/n10428 , \shifter_0/n10425 ,
         \shifter_0/n10424 , \shifter_0/n10421 , \shifter_0/n10420 ,
         \shifter_0/n10417 , \shifter_0/n10416 , \shifter_0/n10413 ,
         \shifter_0/n10412 , \shifter_0/n10409 , \shifter_0/n10408 ,
         \shifter_0/n10405 , \shifter_0/n10404 , \shifter_0/n10401 ,
         \shifter_0/n10400 , \shifter_0/n10397 , \shifter_0/n10396 ,
         \shifter_0/n10393 , \shifter_0/n10392 , \shifter_0/n10389 ,
         \shifter_0/n10388 , \shifter_0/n10385 , \shifter_0/n10384 ,
         \shifter_0/n10381 , \shifter_0/n10380 , \shifter_0/n10377 ,
         \shifter_0/n10376 , \shifter_0/n10373 , \shifter_0/n10372 ,
         \shifter_0/n10369 , \shifter_0/n10368 , \shifter_0/n10365 ,
         \shifter_0/n10364 , \shifter_0/n10361 , \shifter_0/n10360 ,
         \shifter_0/n10357 , \shifter_0/n10356 , \shifter_0/n10353 ,
         \shifter_0/n10352 , \shifter_0/n10349 , \shifter_0/n10348 ,
         \shifter_0/n10345 , \shifter_0/n10344 , \shifter_0/n10341 ,
         \shifter_0/n10340 , \shifter_0/n10337 , \shifter_0/n10336 ,
         \shifter_0/n10333 , \shifter_0/n10332 , \shifter_0/n10329 ,
         \shifter_0/n10328 , \shifter_0/n10325 , \shifter_0/n10324 ,
         \shifter_0/n10321 , \shifter_0/n10320 , \shifter_0/n10317 ,
         \shifter_0/n10316 , \shifter_0/n10313 , \shifter_0/n10312 ,
         \shifter_0/n10309 , \shifter_0/n10308 , \shifter_0/n10305 ,
         \shifter_0/n10304 , \shifter_0/n10301 , \shifter_0/n10300 ,
         \shifter_0/n10297 , \shifter_0/n10296 , \shifter_0/n10293 ,
         \shifter_0/n10292 , \shifter_0/n10289 , \shifter_0/n10288 ,
         \shifter_0/n10285 , \shifter_0/n10284 , \shifter_0/n10281 ,
         \shifter_0/n10280 , \shifter_0/n10277 , \shifter_0/n10276 ,
         \shifter_0/n10273 , \shifter_0/n10272 , \shifter_0/n10269 ,
         \shifter_0/n10268 , \shifter_0/n10265 , \shifter_0/n10264 ,
         \shifter_0/n10261 , \shifter_0/n10260 , \shifter_0/n10257 ,
         \shifter_0/n10256 , \shifter_0/n10253 , \shifter_0/n10252 ,
         \shifter_0/n10249 , \shifter_0/n10248 , \shifter_0/n10245 ,
         \shifter_0/n10244 , \shifter_0/n10241 , \shifter_0/n10240 ,
         \shifter_0/n10237 , \shifter_0/n10236 , \shifter_0/n10233 ,
         \shifter_0/n10232 , \shifter_0/n10229 , \shifter_0/n10228 ,
         \shifter_0/n10225 , \shifter_0/n10224 , \shifter_0/n10221 ,
         \shifter_0/n10220 , \shifter_0/n10217 , \shifter_0/n10216 ,
         \shifter_0/n10213 , \shifter_0/n10212 , \shifter_0/n10209 ,
         \shifter_0/n10208 , \shifter_0/n10205 , \shifter_0/n10204 , n26335,
         n26334, n26333, n26332, n26331, n26330, n26329, n26328, n26327,
         n26326, n26325, n26324, n26323, n26322, n26321, n26320, n26319,
         n26318, n26317, n26316, n26315, n26314, n26313, n26312, n26311,
         n26310, n26309, n26308, n26307, n26306, n26305, n26304, n26303,
         n26302, n26301, n26300, n26299, n26298, n26297, n26296, n26295,
         n26294, n26293, n26292, n26291, n26290, n26289, n26288, n26287,
         n26286, n26285, n26284, n26283, n26282, n26281, n26280, n26279,
         n26278, n26277, n26276, n26275, n26274, n26273, n26272, n26271,
         n26270, n26269, n26268, n26267, n26266, n26265, n26264, n26263,
         n26262, n26261, n26260, n26259, n26258, n26257, n26256, n26255,
         n26254, n26253, n26252, n26251, n26250, n26249, n26248, n26247,
         n26246, n26245, n26244, n26243, n26242, n26241, n26240, n26239,
         n26238, n26237, n26236, n26235, n26234, n26233, n26232, n26231,
         n26230, n26229, n26228, n26227, n26226, n26225, n26224, n26223,
         n26222, n26221, n26220, n26219, n26218, n26217, n26216, n26215,
         n26214, n26213, n26212, n26211, n26210, n26209, n26208, n26207,
         n26206, n26205, n26204, n26203, n26202, n26201, n26200, n26199,
         n26198, n26197, n26196, n26195, n26194, n26193, n26192, n26191,
         n26190, n26189, n26188, n26187, n26186, n26185, n26184, n26183,
         n26182, n26181, n26180, n26179, n26178, n26177, n26176, n26175,
         n26174, n26173, n26172, n26171, n26170, n26169, n26168, n26167,
         n26166, n26165, n26164, n26163, n26162, n26161, n26160, n26159,
         n26158, n26157, n26156, n26155, n26154, n26153, n26152, n26151,
         n26150, n26149, n26148, n26147, n26146, n26145, n26144, n26143,
         n26142, n26141, n26140, n26139, n26138, n26137, n26136, n26135,
         n26134, n26133, n26132, n26131, n26130, n26129, n26128, n26127,
         n26126, n26125, n26124, n26123, n26122, n26121, n26120, n26119,
         n26118, n26117, n26116, n26115, n26114, n26113, n26112, n26111,
         n26110, n26109, n26108, n26107, n26106, n26105, n26104, n26103,
         n26102, n26101, n26100, n26099, n26098, n26097, n26096, n26095,
         n26094, n26093, n26092, n26091, n26090, n26089, n26088, n26087,
         n26086, n26085, n26084, n26083, n26082, n26081, n26080, n26079,
         n26078, n26077, n26076, n26075, n26074, n26073, n26072, n26071,
         n26070, n26069, n26068, n26067, n26066, n26065, n26064, n26063,
         n26062, n26061, n26060, n26059, n26058, n26057, n26056, n26055,
         n26054, n26053, n26052, n26051, n26050, n26049, n26048, n26047,
         n26046, n26045, n26044, n26043, n26042, n26041, n26040, n26039,
         n26038, n26037, n26036, n26035, n26034, n26033, n26032, n26031,
         n26030, n26029, n26028, n26027, n26026, n26025, n26024, n26023,
         n26022, n26021, n26020, n26019, n26018, n26017, n26016, n26015,
         n26014, n26013, n26012, n26011, n26010, n26009, n26008, n26007,
         n26006, n26003, n26002, n26001, n25996, n25995, n25992, n25991,
         n25990, n25987, n25986, n25985, n25984, n25983, n25982, n25981,
         n25980, n25979, n25978, n25977, n25976, n25974, n25973, n25972,
         n25971, n25970, n25965, n25964, n25961, n25960, n25959, n25956,
         n25955, n25954, n25953, n25952, n25951, n25950, n25949, n25948,
         n25947, n25946, n25945, n25944, n25943, n25942, n25941, n25940,
         n25935, n25934, n25931, n25930, n25929, n25926, n25925, n25924,
         n25923, n25922, n25921, n25920, n25919, n25918, n25917, n25916,
         n25915, n25914, n25913, n25912, n25911, n25910, n25905, n25904,
         n25901, n25900, n25899, n25896, n25895, n25894, n25893, n25892,
         n25891, n25890, n25889, n25888, n25887, n25886, n25885, n25884,
         n25883, n25882, n25881, n25880, n25875, n25874, n25871, n25870,
         n25869, n25866, n25865, n25864, n25863, n25862, n25861, n25860,
         n25859, n25858, n25857, n25856, n25855, n25854, n25853, n25852,
         n25851, n25850, n25845, n25844, n25841, n25840, n25839, n25836,
         n25835, n25834, n25833, n25832, n25831, n25830, n25829, n25828,
         n25827, n25826, n25825, n25824, n25823, n25822, n25821, n25820,
         n25815, n25814, n25811, n25810, n25809, n25806, n25805, n25804,
         n25803, n25802, n25801, n25800, n25799, n25798, n25797, n25796,
         n25795, n25794, n25793, n25792, n25791, n25790, n25785, n25784,
         n25781, n25780, n25779, n25776, n25775, n25774, n25773, n25772,
         n25771, n25770, n25769, n25768, n25767, n25766, n25765, n25764,
         n25763, n25762, n25761, n25760, n25755, n25754, n25751, n25750,
         n25749, n25746, n25745, n25744, n25743, n25742, n25741, n25740,
         n25739, n25738, n25737, n25736, n25735, n25734, n25733, n25732,
         n25731, n25730, n25725, n25724, n25721, n25720, n25719, n25716,
         n25715, n25714, n25713, n25712, n25711, n25710, n25709, n25708,
         n25707, n25706, n25705, n25704, n25703, n25702, n25701, n25700,
         n25695, n25694, n25691, n25690, n25689, n25686, n25685, n25684,
         n25683, n25682, n25681, n25680, n25679, n25678, n25677, n25676,
         n25675, n25674, n25673, n25672, n25671, n25670, n25665, n25664,
         n25661, n25660, n25659, n25656, n25655, n25654, n25653, n25652,
         n25651, n25650, n25649, n25648, n25647, n25646, n25645, n25644,
         n25643, n25642, n25641, n25640, n25635, n25634, n25631, n25630,
         n25629, n25626, n25625, n25624, n25623, n25622, n25621, n25620,
         n25619, n25618, n25617, n25616, n25615, n25614, n25613, n25612,
         n25611, n25610, n25605, n25604, n25601, n25600, n25599, n25596,
         n25595, n25594, n25593, n25592, n25591, n25590, n25589, n25588,
         n25587, n25586, n25585, n25584, n25583, n25582, n25581, n25580,
         n25575, n25574, n25571, n25570, n25569, n25566, n25565, n25564,
         n25563, n25562, n25561, n25560, n25559, n25558, n25557, n25556,
         n25555, n25554, n25553, n25552, n25551, n25550, n25545, n25544,
         n25541, n25540, n25539, n25536, n25535, n25534, n25533, n25532,
         n25531, n25530, n25529, n25528, n25527, n25526, n25525, n25524,
         n25523, n25522, n25521, n25520, n25515, n25514, n25511, n25510,
         n25509, n25506, n25505, n25504, n25503, n25502, n25501, n25500,
         n25499, n25498, n25497, n25496, n25495, n25494, n25493, n25492,
         n25491, n25490, n25485, n25484, n25481, n25480, n25479, n25476,
         n25475, n25474, n25473, n25472, n25471, n25470, n25469, n25468,
         n25467, n25466, n25465, n25464, n25463, n25462, n25461, n25460,
         n25455, n25454, n25451, n25450, n25449, n25446, n25445, n25444,
         n25443, n25442, n25441, n25440, n25439, n25438, n25437, n25436,
         n25435, n25434, n25433, n25432, n25431, n25430, n25425, n25424,
         n25421, n25420, n25419, n25416, n25415, n25414, n25413, n25412,
         n25411, n25410, n25409, n25408, n25407, n25406, n25405, n25404,
         n25403, n25402, n25401, n25400, n25399, n25394, n25393, n25390,
         n25389, n25388, n25385, n25384, n25383, n25382, n25381, n25380,
         n25379, n25378, n25377, n25376, n25375, n25374, n25372, n25371,
         n25370, n25369, n25368, n25363, n25362, n25359, n25358, n25357,
         n25354, n25353, n25352, n25351, n25350, n25349, n25348, n25347,
         n25346, n25345, n25344, n25343, n25342, n25341, n25340, n25339,
         n25338, n25333, n25332, n25329, n25328, n25327, n25324, n25323,
         n25322, n25321, n25320, n25319, n25318, n25317, n25316, n25315,
         n25314, n25313, n25312, n25311, n25310, n25309, n25308, n25303,
         n25302, n25299, n25298, n25297, n25294, n25293, n25292, n25291,
         n25290, n25289, n25288, n25287, n25286, n25285, n25284, n25283,
         n25282, n25281, n25280, n25279, n25278, n25273, n25272, n25269,
         n25268, n25267, n25264, n25263, n25262, n25261, n25260, n25259,
         n25258, n25257, n25256, n25255, n25254, n25253, n25252, n25251,
         n25250, n25249, n25248, n25243, n25242, n25239, n25238, n25237,
         n25234, n25233, n25232, n25231, n25230, n25229, n25228, n25227,
         n25226, n25225, n25224, n25223, n25222, n25221, n25220, n25219,
         n25218, n25213, n25212, n25209, n25208, n25207, n25204, n25203,
         n25202, n25201, n25200, n25199, n25198, n25197, n25196, n25195,
         n25194, n25193, n25192, n25191, n25190, n25189, n25188, n25183,
         n25182, n25179, n25178, n25177, n25174, n25173, n25172, n25171,
         n25170, n25169, n25168, n25167, n25166, n25165, n25164, n25163,
         n25162, n25161, n25160, n25159, n25158, n25153, n25152, n25149,
         n25148, n25147, n25144, n25143, n25142, n25141, n25140, n25139,
         n25138, n25137, n25136, n25135, n25134, n25133, n25132, n25131,
         n25130, n25129, n25128, n25123, n25122, n25119, n25118, n25117,
         n25114, n25113, n25112, n25111, n25110, n25109, n25108, n25107,
         n25106, n25105, n25104, n25103, n25102, n25101, n25100, n25099,
         n25098, n25093, n25092, n25089, n25088, n25087, n25084, n25083,
         n25082, n25081, n25080, n25079, n25078, n25077, n25076, n25075,
         n25074, n25073, n25072, n25071, n25070, n25069, n25068, n25063,
         n25062, n25059, n25058, n25057, n25054, n25053, n25052, n25051,
         n25050, n25049, n25048, n25047, n25046, n25045, n25044, n25043,
         n25042, n25041, n25040, n25039, n25038, n25033, n25032, n25029,
         n25028, n25027, n25024, n25023, n25022, n25021, n25020, n25019,
         n25018, n25017, n25016, n25015, n25014, n25013, n25012, n25011,
         n25010, n25009, n25008, n25003, n25002, n24999, n24998, n24997,
         n24994, n24993, n24992, n24991, n24990, n24989, n24988, n24987,
         n24986, n24985, n24984, n24983, n24982, n24981, n24980, n24979,
         n24978, n24973, n24972, n24969, n24968, n24967, n24964, n24963,
         n24962, n24961, n24960, n24959, n24958, n24957, n24956, n24955,
         n24954, n24953, n24952, n24951, n24950, n24949, n24948, n24943,
         n24942, n24939, n24938, n24937, n24934, n24933, n24932, n24931,
         n24930, n24929, n24928, n24927, n24926, n24925, n24924, n24923,
         n24922, n24921, n24920, n24919, n24918, n24913, n24912, n24909,
         n24908, n24907, n24904, n24903, n24902, n24901, n24900, n24899,
         n24898, n24897, n24896, n24895, n24894, n24893, n24892, n24891,
         n24890, n24889, n24888, n24883, n24882, n24879, n24878, n24877,
         n24874, n24873, n24872, n24871, n24870, n24869, n24868, n24867,
         n24866, n24865, n24864, n24863, n24862, n24861, n24860, n24859,
         n24858, n24853, n24852, n24849, n24848, n24847, n24844, n24843,
         n24842, n24841, n24840, n24839, n24838, n24837, n24836, n24835,
         n24834, n24833, n24832, n24831, n24830, n24829, n24828, n24827,
         n24822, n24821, n24817, n24816, n24815, n24808, n24807, n24806,
         n24805, n24802, n24801, n24799, n24798, n24797, n24796, n24795,
         n24794, n24793, n24792, n24791, n24790, n24789, n24788, n24785,
         n24784, n24783, n24782, n24781, n24780, n24779, n24778, n24777,
         n24776, n24775, n24774, n24773, n24772, n24771, n24770, n24769,
         n24768, n24767, n24766, n24765, n24764, n24763, n24762, n24761,
         n24760, n24759, n24758, n24757, n24756, n24755, n24754, n24753,
         n24752, n24751, n24750, n24749, n24748, n24747, n24746, n24745,
         n24744, n24743, n24742, n24741, n24740, n24739, n24738, n24737,
         n24736, n24735, n24734, n24733, n24732, n24731, n24730, n24729,
         n24728, n24727, n24726, n24725, n24724, n24723, n24722, n24721,
         n24720, n24719, n24718, n24717, n24716, n24715, n24714, n24713,
         n24712, n24711, n24710, n24709, n24708, n24707, n24706, n24705,
         n24704, n24703, n24702, n24701, n24700, n24699, n24698, n24697,
         n24696, n24695, n24692, n24690, n24689, n24688, n24687, n24686,
         n24685, n24684, n24683, n24682, n24681, n24680, n24679, n24678,
         n24677, n24676, n24675, n24674, n24673, n24672, n24671, n24670,
         n24669, n24668, n24667, n24666, n24665, n24664, n24663, n24662,
         n24661, n24660, n24659, n24658, n24657, n24656, n24655, n24654,
         n24653, n24652, n24651, n24650, n24649, n24648, n24647, n24646,
         n24645, n24644, n24643, n24642, n24641, n24640, n24639, n24638,
         n24637, n24636, n24635, n24634, n24633, n24632, n24631, n24630,
         n24629, n24628, n24627, n24626, n24625, n24624, n24623, n24622,
         n24621, n24620, n24619, n24618, n24617, n24616, n24615, n24614,
         n24613, n24612, n24611, n24610, n24609, n24608, n24606, n24605,
         n24604, n24603, n24602, n24601, n24600, n24599, n24597, n24594,
         n24593, n24592, n24591, n24590, n24589, n24588, n24587, n24586,
         n24585, n24584, n24583, n24582, n24581, n24580, n24579, n24578,
         n24577, n24576, n24575, n24574, n24573, n24572, n24571, n24570,
         n24569, n24568, n24567, n24566, n24565, n24564, n24563, n24562,
         n24561, n24560, n24559, n24558, n24557, n24556, n24555, n24554,
         n24553, n24552, n24551, n24550, n24549, n24548, n24547, n24546,
         n24545, n24544, n24543, n24542, n24541, n24540, n24539, n24538,
         n24537, n24536, n24535, n24534, n24533, n24532, n24531, n24530,
         n24529, n24528, n24527, n24526, n24525, n24524, n24523, n24522,
         n24521, n24520, n24519, n24518, n24517, n24516, n24515, n24514,
         n24513, n24512, n24511, n24510, n24509, n24508, n24507, n24506,
         n24505, n24504, n24503, n24502, n24501, n24500, n24499, n24498,
         n24497, n24496, n24495, n24494, n24493, n24492, n24491, n24490,
         n24489, n24488, n24487, n24485, n24482, n24481, n24480, n24479,
         n24478, n24477, n24476, n24475, n24474, n24473, n24472, n24471,
         n24470, n24469, n24468, n24467, n24466, n24465, n24464, n24463,
         n24462, n24461, n24460, n24459, n24458, n24457, n24456, n24455,
         n24454, n24453, n24452, n24451, n24450, n24449, n24448, n24447,
         n24446, n24445, n24444, n24443, n24442, n24441, n24440, n24439,
         n24438, n24437, n24436, n24435, n24434, n24433, n24432, n24431,
         n24430, n24429, n24428, n24427, n24426, n24425, n24424, n24423,
         n24422, n24421, n24420, n24419, n24418, n24417, n24416, n24415,
         n24414, n24413, n24412, n24411, n24410, n24409, n24408, n24407,
         n24406, n24405, n24404, n24403, n24402, n24401, n24400, n24399,
         n24398, n24397, n24396, n24395, n24394, n24393, n24392, n24391,
         n24390, n24389, n24388, n24387, n24386, n24385, n24384, n24383,
         n24382, n24381, n24380, n24379, n24378, n24377, n24376, n24375,
         n24374, n24373, n24372, n24371, n24370, n24369, n24368, n24367,
         n24366, n24365, n24364, n24363, n24362, n24361, n24360, n24359,
         n24358, n24357, n24356, n24355, n24354, n24353, n24352, n24351,
         n24350, n24349, n24348, n24347, n24346, n24345, n24344, n24343,
         n24342, n24341, n24340, n24339, n24338, n24337, n24336, n24335,
         n24334, n24333, n24332, n24331, n24330, n24329, n24328, n24327,
         n24326, n24325, n24324, n24323, n24322, n24321, n24320, n24319,
         n24318, n24317, n24316, n24315, n24314, n24313, n24312, n24311,
         n24310, n24309, n24308, n24307, n24306, n24305, n24304, n24303,
         n24302, n24301, n24300, n24299, n24298, n24297, n24296, n24295,
         n24294, n24293, n24292, n24291, n24290, n24289, n24288, n24287,
         n24286, n24285, n24284, n24283, n24282, n24281, n24280, n24279,
         n24278, n24277, n24276, n24275, n24274, n24273, n24272, n24271,
         n24270, n24269, n24268, n24267, n24266, n24265, n24264, n24263,
         n24262, n24261, n24260, n24259, n24258, n24257, n24256, n24255,
         n24254, n24253, n24252, n24251, n24250, n24249, n24248, n24247,
         n24246, n24245, n24244, n24243, n24242, n24241, n24240, n24239,
         n24238, n24237, n24236, n24235, n24234, n24233, n24232, n24231,
         n24230, n24229, n24228, n24227, n24226, n24225, n24224, n24223,
         n24222, n24221, n24220, n24219, n24218, n24217, n24216, n24215,
         n24214, n24213, n24212, n24211, n24210, n24209, n24208, n24207,
         n24206, n24205, n24204, n24203, n24202, n24201, n24200, n24199,
         n24198, n24197, n24196, n24195, n24194, n24193, n24192, n24191,
         n24190, n24189, n24188, n24187, n24186, n24185, n24184, n24183,
         n24182, n24181, n24180, n24179, n24178, n24177, n24176, n24175,
         n24174, n24173, n24172, n24171, n24170, n24169, n24168, n24167,
         n24166, n24165, n24164, n24163, n24162, n24161, n24160, n24159,
         n24158, n24157, n24156, n24155, n24154, n24153, n24152, n24151,
         n24150, n24149, n24148, n24147, n24146, n24145, n24144, n24143,
         n24142, n24141, n24140, n24139, n24138, n24137, n24136, n24135,
         n24134, n24133, n24132, n24131, n24130, n24129, n24128, n24127,
         n24126, n24125, n24124, n24123, n24122, n24121, n24120, n24119,
         n24118, n24117, n24116, n24115, n24114, n24113, n24112, n24111,
         n24110, n24109, n24108, n24107, n24106, n24105, n24104, n24103,
         n24102, n24101, n24100, n24099, n24098, n24097, n24096, n24095,
         n24094, n24093, n24092, n24091, n24090, n24089, n24088, n24087,
         n24086, n24085, n24084, n24083, n24082, n24081, n24080, n24079,
         n24078, n24077, n24076, n24075, n24074, n24073, n24072, n24071,
         n24070, n24069, n24068, n24067, n24066, n24065, n24064, n24063,
         n24062, n24061, n24060, n24059, n24058, n24057, n24056, n24055,
         n24054, n24053, n24052, n24050, n24049, n24047, n24046, n24045,
         n24044, n24043, n24042, n24041, n24040, n24039, n24038, n24037,
         n24036, n24035, n24034, n24033, n24032, n24031, n24030, n24029,
         n24028, n24027, n24026, n24025, n24024, n24023, n24022, n24021,
         n24020, n24019, n24018, n24017, n24016, n24015, n24014, n24013,
         n24012, n24011, n24010, n24009, n24008, n24007, n24006, n24005,
         n24004, n24003, n24002, n24001, n24000, n23999, n23998, n23997,
         n23996, n23995, n23994, n23993, n23992, n23991, n23990, n23989,
         n23988, n23987, n23986, n23985, n23984, n23983, n23982, n23981,
         n23980, n23979, n23978, n23977, n23976, n23975, n23974, n23973,
         n23972, n23971, n23970, n23969, n23968, n23967, n23966, n23965,
         n23964, n23963, n23962, n23961, n23960, n23959, n23958, n23957,
         n23956, n23955, n23954, n23953, n23952, n23951, n23950, n23949,
         n23948, n23947, n23946, n23945, n23944, n23943, n23942, n23940,
         n23939, n23938, n23936, n23935, n23934, n23933, n23932, n23931,
         n23930, n23929, n23928, n23926, n23925, n23924, n23923, n23922,
         n23920, n23919, n23918, n23917, n23916, n23914, n23913, n23912,
         n23911, n23910, n23908, n23907, n23906, n23905, n23904, n23902,
         n23901, n23900, n23899, n23898, n23896, n23895, n23894, n23893,
         n23892, n23890, n23889, n23888, n23887, n23886, n23884, n23883,
         n23882, n23881, n23880, n23878, n23877, n23876, n23875, n23874,
         n23872, n23871, n23870, n23869, n23868, n23866, n23865, n23864,
         n23863, n23862, n23860, n23859, n23858, n23857, n23856, n23854,
         n23853, n23852, n23851, n23850, n23848, n23847, n23846, n23845,
         n23844, n23842, n23841, n23840, n23839, n23838, n23836, n23835,
         n23834, n23833, n23832, n23830, n23829, n23828, n23827, n23826,
         n23824, n23823, n23822, n23821, n23820, n23818, n23817, n23816,
         n23815, n23814, n23813, n23811, n23810, n23809, n23807, n23806,
         n23805, n23804, n23803, n23802, n23801, n23800, n23799, n23797,
         n23796, n23795, n23794, n23793, n23791, n23790, n23789, n23788,
         n23787, n23785, n23784, n23783, n23782, n23781, n23779, n23778,
         n23777, n23776, n23775, n23773, n23772, n23771, n23770, n23769,
         n23767, n23766, n23765, n23764, n23763, n23761, n23760, n23759,
         n23758, n23757, n23755, n23754, n23753, n23752, n23751, n23749,
         n23748, n23747, n23746, n23745, n23743, n23742, n23741, n23740,
         n23739, n23737, n23736, n23735, n23734, n23733, n23731, n23730,
         n23729, n23728, n23727, n23725, n23724, n23723, n23722, n23721,
         n23719, n23718, n23717, n23716, n23715, n23713, n23712, n23711,
         n23710, n23709, n23707, n23706, n23705, n23704, n23703, n23701,
         n23700, n23699, n23698, n23697, n23695, n23694, n23693, n23692,
         n23691, n23688, n23687, n23686, n23685, n23684, n23683, n23682,
         n23681, n23680, n23677, n23675, n23674, n23673, n23672, n23671,
         n23670, n23669, n23668, n23667, n23666, n23665, n23664, n23663,
         n23662, n23661, n23660, n23659, n23658, n23657, n23656, n23655,
         n23654, n23653, n23652, n23651, n23650, n23649, n23648, n23647,
         n23646, n23645, n23644, n23643, n23642, n23641, n23640, n23639,
         n23638, n23637, n23636, n23635, n23634, n23633, n23632, n23631,
         n23630, n23629, n23628, n23627, n23626, n23625, n23624, n23623,
         n23622, n23621, n23620, n23619, n23618, n23617, n23616, n23615,
         n23614, n23613, n23612, n23611, n23610, n23609, n23608, n23607,
         n23606, n23605, n23604, n23603, n23602, n23601, n23600, n23599,
         n23598, n23597, n23596, n23595, n23594, n23593, n23592, n23591,
         n23590, n23589, n23588, n23587, n23586, n23585, n23584, n23583,
         n23582, n23581, n23580, n23579, n23578, n23577, n23576, n23575,
         n23574, n23573, n23572, n23571, n23570, n23569, n23568, n23567,
         n23566, n23565, n23564, n23563, n23562, n23561, n23560, n23559,
         n23558, n23557, n23556, n23555, n23554, n23553, n23552, n23551,
         n23550, n23549, n23546, n23543, n23542, n23541, n23540, n23539,
         n23538, n23537, n23536, n23535, n23534, n23533, n23532, n23531,
         n23530, n23529, n23528, n23527, n23526, n23525, n23524, n23523,
         n23522, n23521, n23520, n23519, n23518, n23517, n23516, n23515,
         n23514, n23513, n23512, n23511, n23510, n23509, n23508, n23507,
         n23506, n23505, n23504, n23503, n23502, n23501, n23500, n23499,
         n23498, n23497, n23496, n23495, n23494, n23493, n23492, n23491,
         n23490, n23489, n23488, n23487, n23486, n23485, n23484, n23483,
         n23482, n23481, n23480, n23479, n23478, n23477, n23476, n23475,
         n23474, n23473, n23472, n23471, n23470, n23469, n23468, n23467,
         n23466, n23465, n23464, n23463, n23462, n23461, n23460, n23459,
         n23458, n23457, n23456, n23455, n23454, n23453, n23452, n23451,
         n23450, n23449, n23448, n23447, n23446, n23445, n23444, n23443,
         n23442, n23441, n23440, n23439, n23438, n23437, n23436, n23435,
         n23434, n23433, n23432, n23431, n23430, n23429, n23428, n23427,
         n23424, n23423, n23422, n23421, n23420, n23419, n23418, n23417,
         n23416, n23415, n23414, n23413, n23412, n23411, n23410, n23409,
         n23408, n23407, n23406, n23405, n23404, n23403, n23402, n23401,
         n23400, n23399, n23398, n23397, n23396, n23395, n23394, n23393,
         n23392, n23391, n23390, n23389, n23388, n23387, n23386, n23385,
         n23384, n23383, n23382, n23381, n23380, n23379, n23378, n23377,
         n23376, n23375, n23374, n23373, n23372, n23371, n23370, n23369,
         n23368, n23367, n23366, n23365, n23364, n23363, n23362, n23361,
         n23360, n23359, n23358, n23357, n23356, n23355, n23354, n23353,
         n23352, n23351, n23350, n23349, n23348, n23347, n23346, n23345,
         n23344, n23343, n23342, n23341, n23340, n23339, n23338, n23337,
         n23336, n23335, n23334, n23333, n23332, n23331, n23330, n23329,
         n23328, n23327, n23326, n23325, n23324, n23323, n23322, n23321,
         n23320, n23319, n23318, n23317, n23316, n23315, n23314, n23313,
         n23312, n23311, n23310, n23309, n23308, n23307, n23306, n23305,
         n23304, n23303, n23302, n23301, n23300, n23299, n23298, n23297,
         n23296, n23295, n23294, n23293, n23292, n23291, n23290, n23289,
         n23288, n23287, n23286, n23285, n23284, n23283, n23282, n23281,
         n23280, n23279, n23278, n23277, n23276, n23275, n23274, n23273,
         n23272, n23271, n23270, n23269, n23268, n23267, n23266, n23265,
         n23264, n23263, n23262, n23261, n23260, n23259, n23258, n23257,
         n23256, n23255, n23254, n23253, n23252, n23251, n23250, n23249,
         n23248, n23247, n23246, n23245, n23244, n23243, n23242, n23241,
         n23240, n23239, n23238, n23237, n23236, n23235, n23234, n23233,
         n23232, n23231, n23230, n23229, n23228, n23227, n23226, n23225,
         n23224, n23223, n23222, n23221, n23220, n23219, n23218, n23217,
         n23216, n23215, n23214, n23213, n23212, n23211, n23210, n23209,
         n23208, n23207, n23206, n23205, n23204, n23203, n23202, n23200,
         n23199, n23198, n23197, n23196, n23194, n23193, n23192, n23191,
         n23190, n23189, n23188, n23187, n23186, n23185, n23183, n23182,
         n23181, n23180, n23179, n23178, n23177, n23176, n23175, n23174,
         n23172, n23171, n23170, n23169, n23168, n23167, n23166, n23165,
         n23164, n23163, n23161, n23160, n23159, n23158, n23157, n23156,
         n23155, n23154, n23153, n23152, n23150, n23149, n23148, n23147,
         n23146, n23145, n23144, n23143, n23142, n23141, n23139, n23138,
         n23137, n23136, n23135, n23134, n23133, n23132, n23131, n23130,
         n23128, n23127, n23126, n23125, n23124, n23123, n23122, n23121,
         n23120, n23119, n23117, n23116, n23115, n23114, n23113, n23112,
         n23111, n23110, n23109, n23108, n23106, n23105, n23104, n23103,
         n23102, n23101, n23100, n23099, n23098, n23097, n23095, n23094,
         n23093, n23092, n23091, n23090, n23089, n23088, n23087, n23086,
         n23084, n23083, n23082, n23081, n23080, n23079, n23078, n23077,
         n23076, n23075, n23073, n23072, n23071, n23070, n23069, n23068,
         n23067, n23066, n23065, n23064, n23062, n23061, n23060, n23059,
         n23058, n23057, n23056, n23055, n23054, n23053, n23051, n23050,
         n23049, n23048, n23047, n23046, n23045, n23044, n23043, n23042,
         n23040, n23039, n23038, n23037, n23036, n23035, n23034, n23033,
         n23032, n23031, n23029, n23028, n23027, n23026, n23025, n23024,
         n23023, n23022, n23021, n23020, n23018, n23017, n23016, n23015,
         n23014, n23013, n23012, n23011, n23010, n23009, n23007, n23006,
         n23005, n23004, n23003, n23002, n23001, n23000, n22999, n22998,
         n22996, n22995, n22994, n22993, n22992, n22991, n22990, n22989,
         n22988, n22987, n22986, n22985, n22983, n22982, n22981, n22980,
         n22979, n22978, n22977, n22976, n22975, n22974, n22973, n22972,
         n22971, n22970, n22969, n22967, n22966, n22965, n22964, n22963,
         n22962, n22961, n22960, n22959, n22958, n22956, n22955, n22954,
         n22953, n22952, n22951, n22950, n22949, n22948, n22947, n22945,
         n22944, n22943, n22942, n22941, n22940, n22939, n22938, n22937,
         n22936, n22934, n22933, n22932, n22931, n22930, n22929, n22928,
         n22927, n22926, n22925, n22923, n22922, n22921, n22920, n22919,
         n22918, n22917, n22916, n22915, n22914, n22912, n22911, n22910,
         n22909, n22908, n22907, n22906, n22905, n22904, n22903, n22901,
         n22900, n22899, n22898, n22897, n22896, n22895, n22894, n22893,
         n22892, n22890, n22889, n22888, n22887, n22886, n22885, n22884,
         n22883, n22882, n22881, n22879, n22878, n22877, n22876, n22875,
         n22874, n22873, n22872, n22871, n22870, n22868, n22867, n22866,
         n22865, n22864, n22863, n22862, n22861, n22860, n22859, n22857,
         n22856, n22855, n22854, n22853, n22852, n22851, n22850, n22849,
         n22848, n22846, n22845, n22844, n22843, n22842, n22841, n22840,
         n22839, n22838, n22837, n22835, n22834, n22833, n22832, n22831,
         n22830, n22829, n22828, n22827, n22826, n22824, n22823, n22822,
         n22821, n22820, n22819, n22818, n22817, n22816, n22815, n22813,
         n22812, n22811, n22810, n22809, n22808, n22807, n22806, n22805,
         n22804, n22802, n22801, n22800, n22799, n22798, n22797, n22796,
         n22795, n22794, n22793, n22791, n22790, n22789, n22788, n22787,
         n22786, n22785, n22784, n22783, n22782, n22780, n22779, n22778,
         n22777, n22776, n22775, n22774, n22773, n22772, n22771, n22769,
         n22768, n22767, n22766, n22765, n22764, n22763, n22762, n22761,
         n22760, n22759, n22757, n22755, n22754, n22753, n22752, n22751,
         n22750, n22749, n22748, n22747, n22746, n22745, n22744, n22743,
         n22742, n22741, n22740, n22739, n22738, n22737, n22736, n22735,
         n22734, n22733, n22732, n22731, n22730, n22729, n22728, n22727,
         n22726, n22725, n22724, n22723, n22722, n22721, n22720, n22719,
         n22718, n22717, n22716, n22715, n22714, n22713, n22712, n22711,
         n22710, n22709, n22708, n22707, n22706, n22705, n22704, n22703,
         n22702, n22701, n22700, n22699, n22698, n22697, n22696, n22695,
         n22694, n22693, n22692, n22691, n22690, n22689, n22688, n22687,
         n22686, n22685, n22684, n22683, n22682, n22681, n22680, n22679,
         n22678, n22677, n22676, n22675, n22674, n22673, n22672, n22671,
         n22670, n22669, n22668, n22667, n22666, n22665, n22664, n22663,
         n22662, n22661, n22660, n22659, n22658, n22657, n22656, n22655,
         n22654, n22653, n22652, n22651, n22650, n22649, n22648, n22647,
         n22646, n22645, n22644, n22643, n22642, n22641, n22640, n22639,
         n22638, n22637, n22636, n22635, n22634, n22633, n22632, n22631,
         n22630, n22629, n22628, n22627, n22626, n22625, n22624, n22623,
         n22622, n22621, n22620, n22619, n22618, n22617, n22616, n22615,
         n22614, n22613, n22612, n22611, n22610, n22609, n22608, n22607,
         n22606, n22605, n22604, n22603, n22602, n22601, n22600, n22599,
         n22598, n22597, n22596, n22595, n22594, n22593, n22592, n22591,
         n22590, n22589, n22588, n22587, n22586, n22585, n22584, n22583,
         n22582, n22581, n22580, n22579, n22578, n22577, n22576, n22575,
         n22574, n22573, n22572, n22571, n22570, n22569, n22568, n22567,
         n22566, n22565, n22564, n22563, n22562, n22561, n22560, n22559,
         n22558, n22557, n22556, n22555, n22554, n22553, n22552, n22551,
         n22550, n22549, n22548, n22547, n22546, n22545, n22544, n22543,
         n22542, n22541, n22540, n22539, n22538, n22537, n22536, n22535,
         n22534, n22533, n22532, n22531, n22530, n22529, n22528, n22527,
         n22526, n22525, n22524, n22523, n22522, n22521, n22520, n22519,
         n22518, n22517, n22516, n22515, n22514, n22513, n22512, n22511,
         n22510, n22509, n22508, n22507, n22506, n22505, n22504, n22503,
         n22502, n22501, n22500, n22499, n22498, n22497, n22496, n22495,
         n22494, n22493, n22492, n22491, n22490, n22489, n22488, n22487,
         n22486, n22485, n22484, n22483, n22482, n22481, n22480, n22479,
         n22478, n22477, n22476, n22475, n22474, n22473, n22471, n22470,
         n22469, n22468, n22467, n22466, n22465, n22464, n22463, n22462,
         n22461, n22460, n22459, n22458, n22457, n22456, n22455, n22454,
         n22453, n22452, n22451, n22450, n22449, n22448, n22447, n22446,
         n22445, n22444, n22443, n22442, n22441, n22440, n22439, n22438,
         n22437, n22436, n22435, n22434, n22433, n22432, n22431, n22430,
         n22429, n22428, n22427, n22426, n22425, n22424, n22423, n22422,
         n22421, n22420, n22418, n22417, n22416, n22415, n22414, n22413,
         n22412, n22411, n22410, n22409, n22408, n22407, n22406, n22405,
         n22404, n22403, n22402, n22401, n22400, n22399, n22398, n22397,
         n22396, n22395, \filter_0/n9999 , \filter_0/n9996 , \filter_0/n9995 ,
         \filter_0/n9992 , \filter_0/n9991 , \filter_0/n9988 ,
         \filter_0/n9987 , \filter_0/n9984 , \filter_0/n9983 ,
         \filter_0/n9980 , \filter_0/n9979 , \filter_0/n9976 ,
         \filter_0/n9975 , \filter_0/n9972 , \filter_0/n9971 ,
         \filter_0/n9968 , \filter_0/n9967 , \filter_0/n9964 ,
         \filter_0/n9963 , \filter_0/n9960 , \filter_0/n9959 ,
         \filter_0/n9956 , \filter_0/n9955 , \filter_0/n9952 ,
         \filter_0/n9951 , \filter_0/n9948 , \filter_0/n9947 ,
         \filter_0/n9944 , \filter_0/n9943 , \filter_0/n9940 ,
         \filter_0/n9939 , \filter_0/n9936 , \filter_0/n9935 ,
         \filter_0/n9932 , \filter_0/n9931 , \filter_0/n9928 ,
         \filter_0/n9927 , \filter_0/n9924 , \filter_0/n9923 ,
         \filter_0/n9920 , \filter_0/n9919 , \filter_0/n9916 ,
         \filter_0/n9915 , \filter_0/n9912 , \filter_0/n9911 ,
         \filter_0/n9908 , \filter_0/n9907 , \filter_0/n9904 ,
         \filter_0/n9903 , \filter_0/n9900 , \filter_0/n9899 ,
         \filter_0/n9896 , \filter_0/n9895 , \filter_0/n9892 ,
         \filter_0/n9891 , \filter_0/n9888 , \filter_0/n9887 ,
         \filter_0/n9884 , \filter_0/n9883 , \filter_0/n9880 ,
         \filter_0/n9879 , \filter_0/n9876 , \filter_0/n9875 ,
         \filter_0/n9872 , \filter_0/n9871 , \filter_0/n9868 ,
         \filter_0/n9867 , \filter_0/n9864 , \filter_0/n9863 ,
         \filter_0/n9860 , \filter_0/n9859 , \filter_0/n9856 ,
         \filter_0/n9855 , \filter_0/n9852 , \filter_0/n9851 ,
         \filter_0/n9848 , \filter_0/n9847 , \filter_0/n9844 ,
         \filter_0/n9843 , \filter_0/n9840 , \filter_0/n9839 ,
         \filter_0/n9836 , \filter_0/n9835 , \filter_0/n9832 ,
         \filter_0/n9831 , \filter_0/n9828 , \filter_0/n9827 ,
         \filter_0/n9824 , \filter_0/n9823 , \filter_0/n9820 ,
         \filter_0/n9819 , \filter_0/n9816 , \filter_0/n9815 ,
         \filter_0/n9812 , \filter_0/n9811 , \filter_0/n9808 ,
         \filter_0/n9807 , \filter_0/n9804 , \filter_0/n9803 ,
         \filter_0/n9800 , \filter_0/n9799 , \filter_0/n9796 ,
         \filter_0/n9795 , \filter_0/n9792 , \filter_0/n9791 ,
         \filter_0/n9788 , \filter_0/n9787 , \filter_0/n9784 ,
         \filter_0/n9783 , \filter_0/n9780 , \filter_0/n9779 ,
         \filter_0/n9776 , \filter_0/n9775 , \filter_0/n9772 ,
         \filter_0/n9771 , \filter_0/n9768 , \filter_0/n9767 ,
         \filter_0/n9764 , \filter_0/n9763 , \filter_0/n9760 ,
         \filter_0/n9759 , \filter_0/n9756 , \filter_0/n9755 ,
         \filter_0/n9752 , \filter_0/n9751 , \filter_0/n9748 ,
         \filter_0/n9747 , \filter_0/n9744 , \filter_0/n9743 ,
         \filter_0/n9740 , \filter_0/n9739 , \filter_0/n9736 ,
         \filter_0/n9735 , \filter_0/n9732 , \filter_0/n9731 ,
         \filter_0/n9728 , \filter_0/n9727 , \filter_0/n9724 ,
         \filter_0/n9723 , \filter_0/n9720 , \filter_0/n9719 ,
         \filter_0/n9716 , \filter_0/n9715 , \filter_0/n9712 ,
         \filter_0/n9711 , \filter_0/n9708 , \filter_0/n9707 ,
         \filter_0/n9704 , \filter_0/n9703 , \filter_0/n9700 ,
         \filter_0/n9699 , \filter_0/n9696 , \filter_0/n9695 ,
         \filter_0/n9692 , \filter_0/n9691 , \filter_0/n9688 ,
         \filter_0/n9687 , \filter_0/n9684 , \filter_0/n9683 ,
         \filter_0/n9680 , \filter_0/n9679 , \filter_0/n9676 ,
         \filter_0/n9675 , \filter_0/n9672 , \filter_0/n9671 ,
         \filter_0/n9668 , \filter_0/n9667 , \filter_0/n9664 ,
         \filter_0/n9663 , \filter_0/n9660 , \filter_0/n9659 ,
         \filter_0/n9656 , \filter_0/n9655 , \filter_0/n9652 ,
         \filter_0/n9651 , \filter_0/n9648 , \filter_0/n9647 ,
         \filter_0/n9644 , \filter_0/n9643 , \filter_0/n9640 ,
         \filter_0/n9639 , \filter_0/n9636 , \filter_0/n9635 ,
         \filter_0/n9632 , \filter_0/n9631 , \filter_0/n9628 ,
         \filter_0/n9627 , \filter_0/n9624 , \filter_0/n9623 ,
         \filter_0/n9620 , \filter_0/n9619 , \filter_0/n9616 ,
         \filter_0/n9615 , \filter_0/n9612 , \filter_0/n9611 ,
         \filter_0/n9608 , \filter_0/n9607 , \filter_0/n9604 ,
         \filter_0/n9603 , \filter_0/n9600 , \filter_0/n9599 ,
         \filter_0/n9596 , \filter_0/n9595 , \filter_0/n9592 ,
         \filter_0/n9591 , \filter_0/n9588 , \filter_0/n9587 ,
         \filter_0/n9584 , \filter_0/n9583 , \filter_0/n9580 ,
         \filter_0/n9579 , \filter_0/n9576 , \filter_0/n9575 ,
         \filter_0/n9572 , \filter_0/n9571 , \filter_0/n9568 ,
         \filter_0/n9567 , \filter_0/n9564 , \filter_0/n9563 ,
         \filter_0/n9560 , \filter_0/n9559 , \filter_0/n9556 ,
         \filter_0/n9555 , \filter_0/n9552 , \filter_0/n9551 ,
         \filter_0/n9548 , \filter_0/n9547 , \filter_0/n9544 ,
         \filter_0/n9543 , \filter_0/n9540 , \filter_0/n9539 ,
         \filter_0/n9536 , \filter_0/n9535 , \filter_0/n9532 ,
         \filter_0/n9531 , \filter_0/n9528 , \filter_0/n9527 ,
         \filter_0/n9524 , \filter_0/n9523 , \filter_0/n9520 ,
         \filter_0/n9519 , \filter_0/n9516 , \filter_0/n9515 ,
         \filter_0/n9512 , \filter_0/n9511 , \filter_0/n9508 ,
         \filter_0/n9507 , \filter_0/n9504 , \filter_0/n9503 ,
         \filter_0/n9500 , \filter_0/n9499 , \filter_0/n9496 ,
         \filter_0/n9495 , \filter_0/n9492 , \filter_0/n9491 ,
         \filter_0/n9488 , \filter_0/n9487 , \filter_0/n9484 ,
         \filter_0/n9483 , \filter_0/n9480 , \filter_0/n9479 ,
         \filter_0/n9476 , \filter_0/n9475 , \filter_0/n9472 ,
         \filter_0/n9471 , \filter_0/n9468 , \filter_0/n9467 ,
         \filter_0/n9464 , \filter_0/n9463 , \filter_0/n9460 ,
         \filter_0/n9459 , \filter_0/n9456 , \filter_0/n9455 ,
         \filter_0/n9452 , \filter_0/n9451 , \filter_0/n9448 ,
         \filter_0/n9447 , \filter_0/n9444 , \filter_0/n9443 ,
         \filter_0/n9440 , \filter_0/n9439 , \filter_0/n9436 ,
         \filter_0/n9435 , \filter_0/n9432 , \filter_0/n9431 ,
         \filter_0/n9428 , \filter_0/n9427 , \filter_0/n9424 ,
         \filter_0/n9423 , \filter_0/n9420 , \filter_0/n9419 ,
         \filter_0/n9416 , \filter_0/n9415 , \filter_0/n9412 ,
         \filter_0/n9411 , \filter_0/n9408 , \filter_0/n9407 ,
         \filter_0/n9404 , \filter_0/n9403 , \filter_0/n9400 ,
         \filter_0/n9399 , \filter_0/n9396 , \filter_0/n9395 ,
         \filter_0/n9392 , \filter_0/n9391 , \filter_0/n9388 ,
         \filter_0/n9387 , \filter_0/n9384 , \filter_0/n9383 ,
         \filter_0/n9380 , \filter_0/n9379 , \filter_0/n9376 ,
         \filter_0/n9375 , \filter_0/n9372 , \filter_0/n9371 ,
         \filter_0/n9368 , \filter_0/n9367 , \filter_0/n9364 ,
         \filter_0/n9363 , \filter_0/n9360 , \filter_0/n9359 ,
         \filter_0/n9356 , \filter_0/n9355 , \filter_0/n9352 ,
         \filter_0/n9351 , \filter_0/n9348 , \filter_0/n9347 ,
         \filter_0/n9344 , \filter_0/n9343 , \filter_0/n9340 ,
         \filter_0/n9339 , \filter_0/n9336 , \filter_0/n9335 ,
         \filter_0/n9332 , \filter_0/n9331 , \filter_0/n9328 ,
         \filter_0/n9327 , \filter_0/n9324 , \filter_0/n9323 ,
         \filter_0/n9320 , \filter_0/n9319 , \filter_0/n9316 ,
         \filter_0/n9315 , \filter_0/n9312 , \filter_0/n9311 ,
         \filter_0/n9308 , \filter_0/n9307 , \filter_0/n9304 ,
         \filter_0/n9303 , \filter_0/n9300 , \filter_0/n9299 ,
         \filter_0/n9296 , \filter_0/n9295 , \filter_0/n9292 ,
         \filter_0/n9291 , \filter_0/n9288 , \filter_0/n9287 ,
         \filter_0/n9284 , \filter_0/n9283 , \filter_0/n9280 ,
         \filter_0/n9279 , \filter_0/n9276 , \filter_0/n9275 ,
         \filter_0/n9272 , \filter_0/n9271 , \filter_0/n9268 ,
         \filter_0/n9267 , \filter_0/n9264 , \filter_0/n9263 ,
         \filter_0/n9260 , \filter_0/n9259 , \filter_0/n9256 ,
         \filter_0/n9255 , \filter_0/n9252 , \filter_0/n9251 ,
         \filter_0/n9248 , \filter_0/n9247 , \filter_0/n9244 ,
         \filter_0/n9243 , \filter_0/n9240 , \filter_0/n9239 ,
         \filter_0/n9236 , \filter_0/n9235 , \filter_0/n9232 ,
         \filter_0/n9231 , \filter_0/n9228 , \filter_0/n9227 ,
         \filter_0/n9224 , \filter_0/n9223 , \filter_0/n9220 ,
         \filter_0/n9219 , \filter_0/n9216 , \filter_0/n9215 ,
         \filter_0/n9212 , \filter_0/n9211 , \filter_0/n9208 ,
         \filter_0/n9207 , \filter_0/n9204 , \filter_0/n9203 ,
         \filter_0/n9200 , \filter_0/n9199 , \filter_0/n9196 ,
         \filter_0/n9195 , \filter_0/n9192 , \filter_0/n9191 ,
         \filter_0/n9188 , \filter_0/n9187 , \filter_0/n9184 ,
         \filter_0/n9183 , \filter_0/n9180 , \filter_0/n9179 ,
         \filter_0/n9176 , \filter_0/n9175 , \filter_0/n9172 ,
         \filter_0/n9171 , \filter_0/n9168 , \filter_0/n9167 ,
         \filter_0/n9164 , \filter_0/n9163 , \filter_0/n9160 ,
         \filter_0/n9159 , \filter_0/n9156 , \filter_0/n9155 ,
         \filter_0/n9152 , \filter_0/n9151 , \filter_0/n9148 ,
         \filter_0/n9147 , \filter_0/n9144 , \filter_0/n9143 ,
         \filter_0/n9140 , \filter_0/n9139 , \filter_0/n9136 ,
         \filter_0/n9135 , \filter_0/n9132 , \filter_0/n9131 ,
         \filter_0/n9128 , \filter_0/n9127 , \filter_0/n9124 ,
         \filter_0/n9123 , \filter_0/n9120 , \filter_0/n9119 ,
         \filter_0/n9116 , \filter_0/n9115 , \filter_0/n9112 ,
         \filter_0/n9111 , \filter_0/n9108 , \filter_0/n9107 ,
         \filter_0/n9104 , \filter_0/n9103 , \filter_0/n9100 ,
         \filter_0/n9099 , \filter_0/n9096 , \filter_0/n9095 ,
         \filter_0/n9092 , \filter_0/n9091 , \filter_0/n9088 ,
         \filter_0/n9087 , \filter_0/n9084 , \filter_0/n9083 ,
         \filter_0/n9080 , \filter_0/n9079 , \filter_0/n9076 ,
         \filter_0/n9075 , \filter_0/n9072 , \filter_0/n9071 ,
         \filter_0/n9068 , \filter_0/n9067 , \filter_0/n9064 ,
         \filter_0/n9063 , \filter_0/n9060 , \filter_0/n9059 ,
         \filter_0/n9056 , \filter_0/n9055 , \filter_0/n9052 ,
         \filter_0/n9051 , \filter_0/n9048 , \filter_0/n9047 ,
         \filter_0/n9044 , \filter_0/n9043 , \filter_0/n9040 ,
         \filter_0/n9039 , \filter_0/n9036 , \filter_0/n9035 ,
         \filter_0/n9032 , \filter_0/n9031 , \filter_0/n9028 ,
         \filter_0/n9027 , \filter_0/n9024 , \filter_0/n9023 ,
         \filter_0/n9020 , \filter_0/n9019 , \filter_0/n9016 ,
         \filter_0/n9015 , \filter_0/n9012 , \filter_0/n9011 ,
         \filter_0/n9008 , \filter_0/n9007 , \filter_0/n9004 ,
         \filter_0/n9003 , \filter_0/n9000 , \filter_0/n8999 ,
         \filter_0/n8996 , \filter_0/n8995 , \filter_0/n8992 ,
         \filter_0/n8991 , \filter_0/n8988 , \filter_0/n8987 ,
         \filter_0/n8984 , \filter_0/n8983 , \filter_0/n8980 ,
         \filter_0/n8979 , \filter_0/n8976 , \filter_0/n8975 ,
         \filter_0/n8972 , \filter_0/n8971 , \filter_0/n8968 ,
         \filter_0/n8967 , \filter_0/n8964 , \filter_0/n8963 ,
         \filter_0/n8960 , \filter_0/n8959 , \filter_0/n8956 ,
         \filter_0/n8955 , \filter_0/n8952 , \filter_0/n8951 ,
         \filter_0/n8948 , \filter_0/n8947 , \filter_0/n8944 ,
         \filter_0/n8943 , \filter_0/n8940 , \filter_0/n8939 ,
         \filter_0/n8936 , \filter_0/n8935 , \filter_0/n8932 ,
         \filter_0/n8931 , \filter_0/n8928 , \filter_0/n8927 ,
         \filter_0/n8924 , \filter_0/n8923 , \filter_0/n8920 ,
         \filter_0/n8919 , \filter_0/n8916 , \filter_0/n8915 ,
         \filter_0/n8912 , \filter_0/n8911 , \filter_0/n8908 ,
         \filter_0/n8907 , \filter_0/n8904 , \filter_0/n8903 ,
         \filter_0/n8900 , \filter_0/n8899 , \filter_0/n8896 ,
         \filter_0/n8895 , \filter_0/n8892 , \filter_0/n8891 ,
         \filter_0/n8888 , \filter_0/n8887 , \filter_0/n8884 ,
         \filter_0/n8883 , \filter_0/n8880 , \filter_0/n8879 ,
         \filter_0/n8876 , \filter_0/n8875 , \filter_0/n8872 ,
         \filter_0/n8871 , \filter_0/n8868 , \filter_0/n8867 ,
         \filter_0/n8864 , \filter_0/n8863 , \filter_0/n8860 ,
         \filter_0/n8859 , \filter_0/n8856 , \filter_0/n8855 ,
         \filter_0/n8852 , \filter_0/n8851 , \filter_0/n8848 ,
         \filter_0/n8847 , \filter_0/n8844 , \filter_0/n8843 ,
         \filter_0/n8840 , \filter_0/n8839 , \filter_0/n8836 ,
         \filter_0/n8835 , \filter_0/n8832 , \filter_0/n8831 ,
         \filter_0/n8828 , \filter_0/n8827 , \filter_0/n8824 ,
         \filter_0/n8823 , \filter_0/n8820 , \filter_0/n8819 ,
         \filter_0/n8816 , \filter_0/n8815 , \filter_0/n8812 ,
         \filter_0/n8811 , \filter_0/n8808 , \filter_0/n8807 ,
         \filter_0/n8804 , \filter_0/n8803 , \filter_0/n8800 ,
         \filter_0/n8799 , \filter_0/n8796 , \filter_0/n8795 ,
         \filter_0/n8792 , \filter_0/n8791 , \filter_0/n8788 ,
         \filter_0/n8787 , \filter_0/n8784 , \filter_0/n8783 ,
         \filter_0/n8780 , \filter_0/n8779 , \filter_0/n8776 ,
         \filter_0/n8775 , \filter_0/n8772 , \filter_0/n8771 ,
         \filter_0/n8768 , \filter_0/n8767 , \filter_0/n8764 ,
         \filter_0/n8763 , \filter_0/n8760 , \filter_0/n8759 ,
         \filter_0/n8756 , \filter_0/n8755 , \filter_0/n8752 ,
         \filter_0/n8751 , \filter_0/n8748 , \filter_0/n8747 ,
         \filter_0/n8744 , \filter_0/n8743 , \filter_0/n8740 ,
         \filter_0/n8739 , \filter_0/n8736 , \filter_0/n8735 ,
         \filter_0/n8732 , \filter_0/n8731 , \filter_0/n8728 ,
         \filter_0/n8727 , \filter_0/n8724 , \filter_0/n8723 ,
         \filter_0/n8720 , \filter_0/n8719 , \filter_0/n8716 ,
         \filter_0/n8715 , \filter_0/n8712 , \filter_0/n8711 ,
         \filter_0/n8708 , \filter_0/n8707 , \filter_0/n8704 ,
         \filter_0/n8703 , \filter_0/n8700 , \filter_0/n8699 ,
         \filter_0/n8696 , \filter_0/n8695 , \filter_0/n8692 ,
         \filter_0/n8691 , \filter_0/n8688 , \filter_0/n8687 ,
         \filter_0/n8684 , \filter_0/n8683 , \filter_0/n8680 ,
         \filter_0/n8679 , \filter_0/n8676 , \filter_0/n8675 ,
         \filter_0/n8672 , \filter_0/n8671 , \filter_0/n8668 ,
         \filter_0/n8667 , \filter_0/n8664 , \filter_0/n8663 ,
         \filter_0/n8660 , \filter_0/n8659 , \filter_0/n8656 ,
         \filter_0/n8655 , \filter_0/n8652 , \filter_0/n8651 ,
         \filter_0/n8648 , \filter_0/n8647 , \filter_0/n8644 ,
         \filter_0/n8643 , \filter_0/n8640 , \filter_0/n8639 ,
         \filter_0/n8636 , \filter_0/n8635 , \filter_0/n8632 ,
         \filter_0/n8631 , \filter_0/n8628 , \filter_0/n8627 ,
         \filter_0/n8624 , \filter_0/n8623 , \filter_0/n8620 ,
         \filter_0/n8619 , \filter_0/n8616 , \filter_0/n8615 ,
         \filter_0/n8612 , \filter_0/n8611 , \filter_0/n8608 ,
         \filter_0/n8607 , \filter_0/n8604 , \filter_0/n8603 ,
         \filter_0/n8600 , \filter_0/n8599 , \filter_0/n8596 ,
         \filter_0/n8595 , \filter_0/n8592 , \filter_0/n8591 ,
         \filter_0/n8588 , \filter_0/n8587 , \filter_0/n8584 ,
         \filter_0/n8583 , \filter_0/n8580 , \filter_0/n8579 ,
         \filter_0/n8576 , \filter_0/n8575 , \filter_0/n8572 ,
         \filter_0/n8571 , \filter_0/n8568 , \filter_0/n8567 ,
         \filter_0/n8564 , \filter_0/n8563 , \filter_0/n8560 ,
         \filter_0/n8559 , \filter_0/n8556 , \filter_0/n8555 ,
         \filter_0/n8552 , \filter_0/n8551 , \filter_0/n8548 ,
         \filter_0/n8547 , \filter_0/n8544 , \filter_0/n8543 ,
         \filter_0/n8540 , \filter_0/n8539 , \filter_0/n8536 ,
         \filter_0/n8535 , \filter_0/n8532 , \filter_0/n8531 ,
         \filter_0/n8528 , \filter_0/n8527 , \filter_0/n8524 ,
         \filter_0/n8523 , \filter_0/n8520 , \filter_0/n8519 ,
         \filter_0/n8516 , \filter_0/n8515 , \filter_0/n8512 ,
         \filter_0/n8511 , \filter_0/n8508 , \filter_0/n8507 ,
         \filter_0/n8504 , \filter_0/n8503 , \filter_0/n8500 ,
         \filter_0/n8499 , \filter_0/n8496 , \filter_0/n8495 ,
         \filter_0/n8492 , \filter_0/n8491 , \filter_0/n8488 ,
         \filter_0/n8487 , \filter_0/n8484 , \filter_0/n8483 ,
         \filter_0/n8480 , \filter_0/n8479 , \filter_0/n8476 ,
         \filter_0/n8475 , \filter_0/n8472 , \filter_0/n8471 ,
         \filter_0/n8468 , \filter_0/n8467 , \filter_0/n8464 ,
         \filter_0/n8463 , \filter_0/n8460 , \filter_0/n8459 ,
         \filter_0/n8456 , \filter_0/n8455 , \filter_0/n8452 ,
         \filter_0/n8451 , \filter_0/n8448 , \filter_0/n8447 ,
         \filter_0/n8444 , \filter_0/n8443 , \filter_0/n8440 ,
         \filter_0/n8439 , \filter_0/n8436 , \filter_0/n8435 ,
         \filter_0/n8432 , \filter_0/n8431 , \filter_0/n8428 ,
         \filter_0/n8427 , \filter_0/n8424 , \filter_0/n8423 ,
         \filter_0/n8420 , \filter_0/n8419 , \filter_0/n8416 ,
         \filter_0/n8415 , \filter_0/n8412 , \filter_0/n8411 ,
         \filter_0/n8408 , \filter_0/n8407 , \filter_0/n8404 ,
         \filter_0/n8403 , \filter_0/n8400 , \filter_0/n8399 ,
         \filter_0/n8396 , \filter_0/n8395 , \filter_0/n8392 ,
         \filter_0/n8391 , \filter_0/n8388 , \filter_0/n8387 ,
         \filter_0/n8384 , \filter_0/n8383 , \filter_0/n8380 ,
         \filter_0/n8379 , \filter_0/n8376 , \filter_0/n8375 ,
         \filter_0/n8372 , \filter_0/n8371 , \filter_0/n8368 ,
         \filter_0/n8367 , \filter_0/n8364 , \filter_0/n8363 ,
         \filter_0/n8360 , \filter_0/n8359 , \filter_0/n8356 ,
         \filter_0/n8355 , \filter_0/n8352 , \filter_0/n8351 ,
         \filter_0/n8348 , \filter_0/n8347 , \filter_0/n8344 ,
         \filter_0/n8343 , \filter_0/n8340 , \filter_0/n8339 ,
         \filter_0/n8336 , \filter_0/n8335 , \filter_0/n8332 ,
         \filter_0/n8331 , \filter_0/n8328 , \filter_0/n8327 ,
         \filter_0/n8324 , \filter_0/n8323 , \filter_0/n8320 ,
         \filter_0/n8319 , \filter_0/n8316 , \filter_0/n8315 ,
         \filter_0/n8312 , \filter_0/n8311 , \filter_0/n8308 ,
         \filter_0/n8307 , \filter_0/n8304 , \filter_0/n8303 ,
         \filter_0/n8300 , \filter_0/n8299 , \filter_0/n8296 ,
         \filter_0/n8295 , \filter_0/n8292 , \filter_0/n8291 ,
         \filter_0/n8287 , \filter_0/n8284 , \filter_0/n8279 ,
         \filter_0/n8276 , \filter_0/n8272 , \filter_0/n8271 ,
         \filter_0/n8268 , \filter_0/n8264 , \filter_0/n8259 ,
         \filter_0/n8255 , \filter_0/n8252 , \filter_0/n8247 ,
         \filter_0/n8243 , \filter_0/n8240 , \filter_0/n8236 ,
         \filter_0/n8235 , \filter_0/n10844 , \filter_0/n10843 ,
         \filter_0/n10840 , \filter_0/n10839 , \filter_0/n10836 ,
         \filter_0/n10835 , \filter_0/n10832 , \filter_0/n10831 ,
         \filter_0/n10828 , \filter_0/n10827 , \filter_0/n10824 ,
         \filter_0/n10823 , \filter_0/n10820 , \filter_0/n10819 ,
         \filter_0/n10816 , \filter_0/n10815 , \filter_0/n10812 ,
         \filter_0/n10811 , \filter_0/n10808 , \filter_0/n10807 ,
         \filter_0/n10804 , \filter_0/n10803 , \filter_0/n10800 ,
         \filter_0/n10799 , \filter_0/n10796 , \filter_0/n10795 ,
         \filter_0/n10792 , \filter_0/n10791 , \filter_0/n10788 ,
         \filter_0/n10787 , \filter_0/n10784 , \filter_0/n10783 ,
         \filter_0/n10780 , \filter_0/n10779 , \filter_0/n10776 ,
         \filter_0/n10775 , \filter_0/n10772 , \filter_0/n10771 ,
         \filter_0/n10768 , \filter_0/n10767 , \filter_0/n10764 ,
         \filter_0/n10763 , \filter_0/n10760 , \filter_0/n10759 ,
         \filter_0/n10756 , \filter_0/n10755 , \filter_0/n10752 ,
         \filter_0/n10751 , \filter_0/n10748 , \filter_0/n10747 ,
         \filter_0/n10744 , \filter_0/n10743 , \filter_0/n10740 ,
         \filter_0/n10739 , \filter_0/n10736 , \filter_0/n10735 ,
         \filter_0/n10732 , \filter_0/n10731 , \filter_0/n10728 ,
         \filter_0/n10727 , \filter_0/n10724 , \filter_0/n10723 ,
         \filter_0/n10720 , \filter_0/n10719 , \filter_0/n10716 ,
         \filter_0/n10715 , \filter_0/n10712 , \filter_0/n10711 ,
         \filter_0/n10708 , \filter_0/n10707 , \filter_0/n10704 ,
         \filter_0/n10703 , \filter_0/n10700 , \filter_0/n10699 ,
         \filter_0/n10696 , \filter_0/n10695 , \filter_0/n10692 ,
         \filter_0/n10691 , \filter_0/n10688 , \filter_0/n10687 ,
         \filter_0/n10684 , \filter_0/n10683 , \filter_0/n10680 ,
         \filter_0/n10679 , \filter_0/n10676 , \filter_0/n10675 ,
         \filter_0/n10672 , \filter_0/n10671 , \filter_0/n10668 ,
         \filter_0/n10667 , \filter_0/n10664 , \filter_0/n10663 ,
         \filter_0/n10660 , \filter_0/n10659 , \filter_0/n10656 ,
         \filter_0/n10655 , \filter_0/n10652 , \filter_0/n10651 ,
         \filter_0/n10648 , \filter_0/n10647 , \filter_0/n10644 ,
         \filter_0/n10643 , \filter_0/n10640 , \filter_0/n10639 ,
         \filter_0/n10636 , \filter_0/n10635 , \filter_0/n10632 ,
         \filter_0/n10631 , \filter_0/n10628 , \filter_0/n10627 ,
         \filter_0/n10624 , \filter_0/n10623 , \filter_0/n10620 ,
         \filter_0/n10619 , \filter_0/n10616 , \filter_0/n10615 ,
         \filter_0/n10612 , \filter_0/n10611 , \filter_0/n10608 ,
         \filter_0/n10607 , \filter_0/n10604 , \filter_0/n10603 ,
         \filter_0/n10600 , \filter_0/n10599 , \filter_0/n10596 ,
         \filter_0/n10595 , \filter_0/n10592 , \filter_0/n10591 ,
         \filter_0/n10588 , \filter_0/n10587 , \filter_0/n10584 ,
         \filter_0/n10583 , \filter_0/n10580 , \filter_0/n10579 ,
         \filter_0/n10576 , \filter_0/n10575 , \filter_0/n10572 ,
         \filter_0/n10571 , \filter_0/n10568 , \filter_0/n10567 ,
         \filter_0/n10564 , \filter_0/n10563 , \filter_0/n10560 ,
         \filter_0/n10559 , \filter_0/n10556 , \filter_0/n10555 ,
         \filter_0/n10552 , \filter_0/n10551 , \filter_0/n10548 ,
         \filter_0/n10547 , \filter_0/n10544 , \filter_0/n10543 ,
         \filter_0/n10540 , \filter_0/n10539 , \filter_0/n10536 ,
         \filter_0/n10535 , \filter_0/n10532 , \filter_0/n10531 ,
         \filter_0/n10528 , \filter_0/n10527 , \filter_0/n10524 ,
         \filter_0/n10523 , \filter_0/n10520 , \filter_0/n10519 ,
         \filter_0/n10516 , \filter_0/n10515 , \filter_0/n10512 ,
         \filter_0/n10511 , \filter_0/n10508 , \filter_0/n10507 ,
         \filter_0/n10504 , \filter_0/n10503 , \filter_0/n10500 ,
         \filter_0/n10499 , \filter_0/n10496 , \filter_0/n10495 ,
         \filter_0/n10492 , \filter_0/n10491 , \filter_0/n10488 ,
         \filter_0/n10487 , \filter_0/n10484 , \filter_0/n10483 ,
         \filter_0/n10480 , \filter_0/n10479 , \filter_0/n10476 ,
         \filter_0/n10475 , \filter_0/n10472 , \filter_0/n10471 ,
         \filter_0/n10468 , \filter_0/n10467 , \filter_0/n10464 ,
         \filter_0/n10463 , \filter_0/n10460 , \filter_0/n10459 ,
         \filter_0/n10456 , \filter_0/n10455 , \filter_0/n10452 ,
         \filter_0/n10451 , \filter_0/n10448 , \filter_0/n10447 ,
         \filter_0/n10444 , \filter_0/n10443 , \filter_0/n10440 ,
         \filter_0/n10439 , \filter_0/n10436 , \filter_0/n10435 ,
         \filter_0/n10432 , \filter_0/n10431 , \filter_0/n10428 ,
         \filter_0/n10427 , \filter_0/n10424 , \filter_0/n10423 ,
         \filter_0/n10420 , \filter_0/n10419 , \filter_0/n10416 ,
         \filter_0/n10415 , \filter_0/n10412 , \filter_0/n10411 ,
         \filter_0/n10408 , \filter_0/n10407 , \filter_0/n10404 ,
         \filter_0/n10403 , \filter_0/n10400 , \filter_0/n10399 ,
         \filter_0/n10396 , \filter_0/n10395 , \filter_0/n10392 ,
         \filter_0/n10391 , \filter_0/n10388 , \filter_0/n10387 ,
         \filter_0/n10384 , \filter_0/n10383 , \filter_0/n10380 ,
         \filter_0/n10379 , \filter_0/n10376 , \filter_0/n10375 ,
         \filter_0/n10372 , \filter_0/n10371 , \filter_0/n10368 ,
         \filter_0/n10367 , \filter_0/n10364 , \filter_0/n10363 ,
         \filter_0/n10360 , \filter_0/n10359 , \filter_0/n10356 ,
         \filter_0/n10355 , \filter_0/n10352 , \filter_0/n10351 ,
         \filter_0/n10348 , \filter_0/n10347 , \filter_0/n10344 ,
         \filter_0/n10343 , \filter_0/n10340 , \filter_0/n10339 ,
         \filter_0/n10336 , \filter_0/n10335 , \filter_0/n10332 ,
         \filter_0/n10331 , \filter_0/n10328 , \filter_0/n10327 ,
         \filter_0/n10324 , \filter_0/n10323 , \filter_0/n10320 ,
         \filter_0/n10319 , \filter_0/n10316 , \filter_0/n10315 ,
         \filter_0/n10312 , \filter_0/n10311 , \filter_0/n10308 ,
         \filter_0/n10307 , \filter_0/n10304 , \filter_0/n10303 ,
         \filter_0/n10300 , \filter_0/n10299 , \filter_0/n10296 ,
         \filter_0/n10295 , \filter_0/n10292 , \filter_0/n10291 ,
         \filter_0/n10288 , \filter_0/n10287 , \filter_0/n10284 ,
         \filter_0/n10283 , \filter_0/n10280 , \filter_0/n10279 ,
         \filter_0/n10276 , \filter_0/n10275 , \filter_0/n10272 ,
         \filter_0/n10271 , \filter_0/n10268 , \filter_0/n10267 ,
         \filter_0/n10264 , \filter_0/n10263 , \filter_0/n10260 ,
         \filter_0/n10259 , \filter_0/n10256 , \filter_0/n10255 ,
         \filter_0/n10252 , \filter_0/n10251 , \filter_0/n10248 ,
         \filter_0/n10247 , \filter_0/n10244 , \filter_0/n10243 ,
         \filter_0/n10240 , \filter_0/n10239 , \filter_0/n10236 ,
         \filter_0/n10235 , \filter_0/n10232 , \filter_0/n10231 ,
         \filter_0/n10228 , \filter_0/n10227 , \filter_0/n10224 ,
         \filter_0/n10223 , \filter_0/n10220 , \filter_0/n10219 ,
         \filter_0/n10216 , \filter_0/n10215 , \filter_0/n10212 ,
         \filter_0/n10211 , \filter_0/n10208 , \filter_0/n10207 ,
         \filter_0/n10204 , \filter_0/n10203 , \filter_0/n10200 ,
         \filter_0/n10199 , \filter_0/n10196 , \filter_0/n10195 ,
         \filter_0/n10192 , \filter_0/n10191 , \filter_0/n10188 ,
         \filter_0/n10187 , \filter_0/n10184 , \filter_0/n10183 ,
         \filter_0/n10180 , \filter_0/n10179 , \filter_0/n10176 ,
         \filter_0/n10175 , \filter_0/n10172 , \filter_0/n10171 ,
         \filter_0/n10168 , \filter_0/n10167 , \filter_0/n10164 ,
         \filter_0/n10163 , \filter_0/n10160 , \filter_0/n10159 ,
         \filter_0/n10156 , \filter_0/n10155 , \filter_0/n10152 ,
         \filter_0/n10151 , \filter_0/n10148 , \filter_0/n10147 ,
         \filter_0/n10144 , \filter_0/n10143 , \filter_0/n10140 ,
         \filter_0/n10139 , \filter_0/n10136 , \filter_0/n10135 ,
         \filter_0/n10132 , \filter_0/n10131 , \filter_0/n10128 ,
         \filter_0/n10127 , \filter_0/n10124 , \filter_0/n10123 ,
         \filter_0/n10120 , \filter_0/n10119 , \filter_0/n10116 ,
         \filter_0/n10115 , \filter_0/n10112 , \filter_0/n10111 ,
         \filter_0/n10108 , \filter_0/n10107 , \filter_0/n10104 ,
         \filter_0/n10103 , \filter_0/n10100 , \filter_0/n10099 ,
         \filter_0/n10096 , \filter_0/n10095 , \filter_0/n10092 ,
         \filter_0/n10091 , \filter_0/n10088 , \filter_0/n10087 ,
         \filter_0/n10084 , \filter_0/n10083 , \filter_0/n10080 ,
         \filter_0/n10079 , \filter_0/n10076 , \filter_0/n10075 ,
         \filter_0/n10072 , \filter_0/n10071 , \filter_0/n10068 ,
         \filter_0/n10067 , \filter_0/n10064 , \filter_0/n10063 ,
         \filter_0/n10060 , \filter_0/n10059 , \filter_0/n10056 ,
         \filter_0/n10055 , \filter_0/n10052 , \filter_0/n10051 ,
         \filter_0/n10048 , \filter_0/n10047 , \filter_0/n10044 ,
         \filter_0/n10043 , \filter_0/n10040 , \filter_0/n10039 ,
         \filter_0/n10036 , \filter_0/n10035 , \filter_0/n10032 ,
         \filter_0/n10031 , \filter_0/n10028 , \filter_0/n10027 ,
         \filter_0/n10024 , \filter_0/n10023 , \filter_0/n10020 ,
         \filter_0/n10019 , \filter_0/n10016 , \filter_0/n10015 ,
         \filter_0/n10012 , \filter_0/n10011 , \filter_0/n10008 ,
         \filter_0/n10007 , \filter_0/n10004 , \filter_0/n10003 ,
         \filter_0/n10000 , n46196, n46197, n46198, n46199, n46200, n46201,
         n46202, n46203, n46204, n46205, n46206, n46207, n46208, n46209,
         n46210, n46211, n46212, n46213, n46214, n46215, n46216, n46217,
         n46218, n46219, n46220, n46221, n46222, n46223, n46224, n46225,
         n46226, n46227, n46228, n46229, n46230, n46231, n46232, n46233,
         n46234, n46235, n46236, n46237, n46238, n46239, n46240, n46241,
         n46242, n46243, n46244, n46245, n46246, n46247, n46248, n46249,
         n46250, n46251, n46252, n46253, n46254, n46255, n46256, n46257,
         n46258, n46259, n46260, n46261, n46262, n46263, n46264, n46265,
         n46266, n46267, n46268, n46269, n46270, n46271, n46272, n46273,
         n46274, n46275, n46276, n46277, n46278, n46279, n46280, n46281,
         n46282, n46283, n46284, n46285, n46286, n46287, n46288, n46289,
         n46290, n46291, n46292, n46293, n46294, n46295, n46296, n46297,
         n46298, n46299, n46300, n46301, n46302, n46303, n46304, n46305,
         n46306, n46307, n46308, n46309, n46310, n46311, n46312, n46313,
         n46314, n46315, n46316, n46317, n46318, n46319, n46320, n46321,
         n46322, n46323, n46324, n46325, n46326, n46327, n46328, n46329,
         n46330, n46331, n46332, n46333, n46334, n46335, n46336, n46337,
         n46338, n46339, n46340, n46341, n46342, n46343, n46344, n46345,
         n46346, n46347, n46348, n46349, n46350, n46351, n46352, n46353,
         n46354, n46355, n46356, n46357, n46358, n46359, n46360, n46361,
         n46362, n46363, n46364, n46365, n46366, n46367, n46368, n46369,
         n46370, n46371, n46372, n46373, n46374, n46375, n46376, n46377,
         n46378, n46379, n46380, n46381, n46382, n46383, n46384, n46385,
         n46386, n46387, n46388, n46389, n46390, n46391, n46392, n46393,
         n46394, n46395, n46396, n46397, n46398, n46399, n46400, n46401,
         n46402, n46403, n46404, n46405, n46406, n46407, n46408, n46409,
         n46410, n46411, n46412, n46413, n46414, n46415, n46416, n46417,
         n46418, n46419, n46420, n46421, n46422, n46423, n46424, n46425,
         n46426, n46427, n46428, n46429, n46430, n46431, n46432, n46433,
         n46434, n46435, n46436, n46437, n46438, n46439, n46440, n46441,
         n46442, n46443, n46444, n46445, n46446, n46447, n46448, n46449,
         n46450, n46451, n46452, n46453, n46454, n46455, n46456, n46457,
         n46458, n46459, n46460, n46461, n46462, n46463, n46464, n46465,
         n46466, n46467, n46468, n46469, n46470, n46471, n46472, n46473,
         n46474, n46475, n46476, n46477, n46478, n46479, n46480, n46481,
         n46482, n46483, n46484, n46485, n46486, n46487, n46488, n46489,
         n46490, n46491, n46492, n46493, n46494, n46495, n46496, n46497,
         n46498, n46499, n46500, n46501, n46502, n46503, n46504, n46505,
         n46506, n46507, n46508, n46509, n46510, n46511, n46512, n46513,
         n46514, n46515, n46516, n46517, n46518, n46519, n46520, n46521,
         n46522, n46523, n46524, n46525, n46526, n46527, n46528, n46529,
         n46530, n46531, n46532, n46533, n46534, n46535, n46536, n46537,
         n46538, n46539, n46540, n46541, n46542, n46543, n46544, n46545,
         n46546, n46547, n46548, n46549, n46550, n46551, n46552, n46553,
         n46554, n46555, n46556, n46557, n46558, n46559, n46560, n46561,
         n46562, n46563, n46564, n46565, n46566, n46567, n46568, n46569,
         n46570, n46571, n46572, n46573, n46574, n46575, n46576, n46577,
         n46578, n46579, n46580, n46581, n46582, n46583, n46584, n46585,
         n46586, n46587, n46588, n46589, n46590, n46591, n46592, n46593,
         n46594, n46595, n46596, n46597, n46598, n46599, n46600, n46601,
         n46602, n46603, n46604, n46605, n46606, n46607, n46608, n46609,
         n46610, n46611, n46612, n46613, n46614, n46615, n46616, n46617,
         n46618, n46619, n46620, n46621, n46622, n46623, n46624, n46625,
         n46626, n46627, n46628, n46629, n46630, n46631, n46632, n46633,
         n46634, n46635, n46636, n46637, n46638, n46639, n46640, n46641,
         n46642, n46643, n46644, n46645, n46646, n46647, n46648, n46649,
         n46650, n46651, n46652, n46653, n46654, n46655, n46656, n46657,
         n46658, n46659, n46660, n46661, n46662, n46663, n46664, n46665,
         n46666, n46667, n46668, n46669, n46670, n46671, n46672, n46673,
         n46674, n46675, n46676, n46677, n46678, n46679, n46680, n46681,
         n46682, n46683, n46684, n46685, n46686, n46687, n46688, n46689,
         n46690, n46691, n46692, n46693, n46694, n46695, n46696, n46697,
         n46698, n46699, n46700, n46701, n46702, n46703, n46704, n46705,
         n46706, n46707, n46708, n46709, n46710, n46711, n46712, n46713,
         n46714, n46715, n46716, n46717, n46718, n46719, n46720, n46721,
         n46722, n46723, n46724, n46725, n46726, n46727, n46728, n46729,
         n46730, n46731, n46732, n46733, n46734, n46735, n46736, n46737,
         n46738, n46739, n46740, n46741, n46742, n46743, n46744, n46745,
         n46746, n46747, n46748, n46749, n46750, n46751, n46752, n46753,
         n46754, n46755, n46756, n46757, n46758, n46759, n46760, n46761,
         n46762, n46763, n46764, n46765, n46766, n46767, n46768, n46769,
         n46770, n46771, n46772, n46773, n46774, n46775, n46776, n46777,
         n46778, n46779, n46780, n46781, n46782, n46783, n46784, n46785,
         n46786, n46787, n46788, n46789, n46790, n46791, n46792, n46793,
         n46794, n46795, n46796, n46797, n46798, n46799, n46800, n46801,
         n46802, n46803, n46804, n46805, n46806, n46807, n46808, n46809,
         n46810, n46811, n46812, n46813, n46814, n46815, n46816, n46817,
         n46818, n46819, n46820, n46821, n46822, n46823, n46824, n46825,
         n46826, n46827, n46828, n46829, n46830, n46831, n46832, n46833,
         n46834, n46835, n46836, n46837, n46838, n46839, n46840, n46841,
         n46842, n46843, n46844, n46845, n46846, n46847, n46848, n46849,
         n46850, n46851, n46852, n46853, n46854, n46855, n46856, n46857,
         n46858, n46859, n46860, n46861, n46862, n46863, n46864, n46865,
         n46866, n46867, n46868, n46869, n46870, n46871, n46872, n46873,
         n46874, n46875, n46876, n46877, n46878, n46879, n46880, n46881,
         n46882, n46883, n46884, n46885, n46886, n46887, n46888, n46889,
         n46890, n46891, n46892, n46893, n46894, n46895, n46896, n46897,
         n46898, n46899, n46900, n46901, n46902, n46903, n46904, n46905,
         n46906, n46907, n46908, n46909, n46910, n46911, n46912, n46913,
         n46914, n46915, n46916, n46917, n46918, n46919, n46920, n46921,
         n46922, n46923, n46924, n46925, n46926, n46927, n46928, n46929,
         n46930, n46931, n46932, n46933, n46934, n46935, n46936, n46937,
         n46938, n46939, n46940, n46941, n46942, n46943, n46944, n46945,
         n46946, n46947, n46948, n46949, n46950, n46951, n46952, n46953,
         n46954, n46955, n46956, n46957, n46958, n46959, n46960, n46961,
         n46962, n46963, n46964, n46965, n46966, n46967, n46968, n46969,
         n46970, n46971, n46972, n46973, n46974, n46975, n46976, n46977,
         n46978, n46979, n46980, n46981, n46982, n46983, n46984, n46985,
         n46986, n46987, n46988, n46989, n46990, n46991, n46992, n46993,
         n46994, n46995, n46996, n46997, n46998, n46999, n47000, n47001,
         n47002, n47003, n47004, n47005, n47006, n47007, n47008, n47009,
         n47010, n47011, n47012, n47013, n47014, n47015, n47016, n47017,
         n47018, n47019, n47020, n47021, n47022, n47023, n47024, n47025,
         n47026, n47027, n47028, n47029, n47030, n47031, n47032, n47033,
         n47034, n47035, n47036, n47037, n47038, n47039, n47040, n47041,
         n47042, n47043, n47044, n47045, n47046, n47047, n47048, n47049,
         n47050, n47051, n47052, n47053, n47054, n47055, n47056, n47057,
         n47058, n47059, n47060, n47061, n47062, n47063, n47064, n47065,
         n47066, n47067, n47068, n47069, n47070, n47071, n47072, n47073,
         n47074, n47075, n47076, n47077, n47078, n47079, n47080, n47081,
         n47082, n47083, n47084, n47085, n47086, n47087, n47088, n47089,
         n47090, n47091, n47092, n47093, n47094, n47095, n47096, n47097,
         n47098, n47099, n47100, n47101, n47102, n47103, n47104, n47105,
         n47106, n47107, n47108, n47109, n47110, n47111, n47112, n47113,
         n47114, n47115, n47116, n47117, n47118, n47119, n47120, n47121,
         n47122, n47123, n47124, n47125, n47126, n47127, n47128, n47129,
         n47130, n47131, n47132, n47133, n47134, n47135, n47136, n47137,
         n47138, n47139, n47140, n47141, n47142, n47143, n47144, n47145,
         n47146, n47147, n47148, n47149, n47150, n47151, n47152, n47153,
         n47154, n47155, n47156, n47157, n47158, n47159, n47160, n47161,
         n47162, n47163, n47164, n47165, n47166, n47167, n47168, n47169,
         n47170, n47171, n47172, n47173, n47174, n47175, n47176, n47177,
         n47178, n47179, n47180, n47181, n47182, n47183, n47184, n47185,
         n47186, n47187, n47188, n47189, n47190, n47191, n47192, n47193,
         n47194, n47195, n47196, n47197, n47198, n47199, n47200, n47201,
         n47202, n47203, n47204, n47205, n47206, n47207, n47208, n47209,
         n47210, n47211, n47212, n47213, n47214, n47215, n47216, n47217,
         n47218, n47219, n47220, n47221, n47222, n47223, n47224, n47225,
         n47226, n47227, n47228, n47229, n47230, n47231, n47232, n47233,
         n47234, n47235, n47236, n47237, n47238, n47239, n47240, n47241,
         n47242, n47243, n47244, n47245, n47246, n47247, n47248, n47249,
         n47250, n47251, n47252, n47253, n47254, n47255, n47256, n47257,
         n47258, n47259, n47260, n47261, n47262, n47263, n47264, n47265,
         n47266, n47267, n47268, n47269, n47270, n47271, n47272, n47273,
         n47274, n47275, n47276, n47277, n47278, n47279, n47280, n47281,
         n47282, n47283, n47284, n47285, n47286, n47287, n47288, n47289,
         n47290, n47291, n47292, n47293, n47294, n47295, n47296, n47297,
         n47298, n47299, n47300, n47301, n47302, n47303, n47304, n47305,
         n47306, n47307, n47308, n47309, n47310, n47311, n47312, n47313,
         n47314, n47315, n47316, n47317, n47318, n47319, n47320, n47321,
         n47322, n47323, n47324, n47325, n47326, n47327, n47328, n47329,
         n47330, n47331, n47332, n47333, n47334, n47335, n47336, n47337,
         n47338, n47339, n47340, n47341, n47342, n47343, n47344, n47345,
         n47346, n47347, n47348, n47349, n47350, n47351, n47352, n47353,
         n47354, n47355, n47356, n47357, n47358, n47359, n47360, n47361,
         n47362, n47363, n47364, n47365, n47366, n47367, n47368, n47369,
         n47370, n47371, n47372, n47373, n47374, n47375, n47376, n47377,
         n47378, n47379, n47380, n47381, n47382, n47383, n47384, n47385,
         n47386, n47387, n47388, n47389, n47390, n47391, n47392, n47393,
         n47394, n47395, n47396, n47397, n47398, n47399, n47400, n47401,
         n47402, n47403, n47404, n47405, n47406, n47407, n47408, n47409,
         n47410, n47411, n47412, n47413, n47414, n47415, n47416, n47417,
         n47418, n47419, n47420, n47421, n47422, n47423, n47424, n47425,
         n47426, n47427, n47428, n47429, n47430, n47431, n47432, n47433,
         n47434, n47435, n47436, n47437, n47438, n47439, n47440, n47441,
         n47442, n47443, n47444, n47445, n47446, n47447, n47448, n47449,
         n47450, n47451, n47452, n47453, n47454, n47455, n47456, n47457,
         n47458, n47459, n47460, n47461, n47462, n47463, n47464, n47465,
         n47466, n47467, n47468, n47469, n47470, n47471, n47472, n47473,
         n47474, n47475, n47476, n47477, n47478, n47479, n47480, n47481,
         n47482, n47483, n47484, n47485, n47486, n47487, n47488, n47489,
         n47490, n47491, n47492, n47493, n47494, n47495, n47496, n47497,
         n47498, n47499, n47500, n47501, n47502, n47503, n47504, n47505,
         n47506, n47507, n47508, n47509, n47510, n47511, n47512, n47513,
         n47514, n47515, n47516, n47517, n47518, n47519, n47520, n47521,
         n47522, n47523, n47524, n47525, n47526, n47527, n47528, n47529,
         n47530, n47531, n47532, n47533, n47534, n47535, n47536, n47537,
         n47538, n47539, n47540, n47541, n47542, n47543, n47544, n47545,
         n47546, n47547, n47548, n47549, n47550, n47551, n47552, n47553,
         n47554, n47555, n47556, n47557, n47558, n47559, n47560, n47561,
         n47562, n47563, n47564, n47565, n47566, n47567, n47568, n47569,
         n47570, n47571, n47572, n47573, n47574, n47575, n47576, n47577,
         n47578, n47579, n47580, n47581, n47582, n47583, n47584, n47585,
         n47586, n47587, n47588, n47589, n47590, n47591, n47592, n47593,
         n47594, n47595, n47596, n47597, n47598, n47599, n47600, n47601,
         n47602, n47603, n47604, n47605, n47606, n47607, n47608, n47609,
         n47610, n47611, n47612, n47613, n47614, n47615, n47616, n47617,
         n47618, n47619, n47620, n47621, n47622, n47623, n47624, n47625,
         n47626, n47627, n47628, n47629, n47630, n47631, n47632, n47633,
         n47634, n47635, n47636, n47637, n47638, n47639, n47640, n47641,
         n47642, n47643, n47644, n47645, n47646, n47647, n47648, n47649,
         n47650, n47651, n47652, n47653, n47654, n47655, n47656, n47657,
         n47658, n47659, n47660, n47661, n47662, n47663, n47664, n47665,
         n47666, n47667, n47668, n47669, n47670, n47671, n47672, n47673,
         n47674, n47675, n47676, n47677, n47678, n47679, n47680, n47681,
         n47682, n47683, n47684, n47685, n47686, n47687, n47688, n47689,
         n47690, n47691, n47692, n47693, n47694, n47695, n47696, n47697,
         n47698, n47699, n47700, n47701, n47702, n47703, n47704, n47705,
         n47706, n47707, n47708, n47709, n47710, n47711, n47712, n47713,
         n47714, n47715, n47716, n47717, n47718, n47719, n47720, n47721,
         n47722, n47723, n47724, n47725, n47726, n47727, n47728, n47729,
         n47730, n47731, n47732, n47733, n47734, n47735, n47736, n47737,
         n47738, n47739, n47740, n47742, n47743, n47744, n47745, n47746,
         n47747, n47748, n47749, n47750, n47751, n47752, n47753, n47754,
         n47755, n47756, n47757, n47758, n47759, n47760, n47761, n47762,
         n47763, n47764, n47765, n47766, n47767, n47768, n47769, n47770,
         n47771, n47772, n47773, n47774, n47775, n47776, n47777, n47778,
         n47779, n47780, n47781, n47782, n47783, n47784, n47785, n47786,
         n47787, n47788, n47789, n47790, n47791, n47792, n47793, n47794,
         n47795, n47796, n47797, n47798, n47799, n47800, n47801, n47802,
         n47803, n47804, n47805, n47806, n47807, n47808, n47809, n47810,
         n47811, n47812, n47813, n47814, n47815, n47816, n47817, n47818,
         n47819, n47820, n47821, n47822, n47823, n47824, n47825, n47826,
         n47827, n47828, n47829, n47830, n47831, n47832, n47833, n47834,
         n47835, n47836, n47837, n47838, n47839, n47840, n47841, n47842,
         n47843, n47844, n47845, n47846, n47847, n47848, n47849, n47850,
         n47851, n47852, n47853, n47854, n47855, n47856, n47857, n47858,
         n47859, n47860, n47861, n47862, n47863, n47864, n47865, n47866,
         n47867, n47868, n47869, n47870, n47871, n47872, n47873, n47874,
         n47875, n47876, n47877, n47878, n47879, n47880, n47881, n47882,
         n47883, n47884, n47885, n47886, n47887, n47888, n47889, n47890,
         n47891, n47892, n47893, n47894, n47895, n47896, n47897, n47898,
         n47899, n47900, n47901, n47902, n47903, n47904, n47905, n47906,
         n47907, n47908, n47909, n47910, n47911, n47912, n47913, n47914,
         n47915, n47916, n47917, n47918, n47919, n47920, n47921, n47922,
         n47923, n47924, n47925, n47926, n47927, n47928, n47929, n47930,
         n47931, n47932, n47933, n47934, n47935, n47936, n47937, n47938,
         n47939, n47940, n47941, n47942, n47943, n47944, n47945, n47946,
         n47947, n47948, n47949, n47950, n47951, n47952, n47953, n47954,
         n47955, n47956, n47957, n47958, n47959, n47960, n47961, n47962,
         n47963, n47964, n47965, n47966, n47967, n47968, n47969, n47970,
         n47971, n47972, n47973, n47974, n47975, n47976, n47977, n47978,
         n47979, n47980, n47981, n47982, n47983, n47984, n47985, n47986,
         n47987, n47988, n47989, n47990, n47991, n47992, n47993, n47994,
         n47995, n47996, n47997, n47998, n47999, n48000, n48001, n48002,
         n48003, n48004, n48005, n48006, n48007, n48008, n48009, n48010,
         n48011, n48012, n48013, n48014, n48015, n48016, n48017, n48018,
         n48019, n48020, n48021, n48022, n48023, n48024, n48025, n48026,
         n48027, n48028, n48029, n48030, n48031, n48032, n48033, n48034,
         n48035, n48036, n48037, n48038, n48039, n48040, n48041, n48042,
         n48043, n48044, n48045, n48046, n48047, n48048, n48049, n48050,
         n48051, n48052, n48053, n48054, n48055, n48056, n48057, n48058,
         n48059, n48060, n48061, n48062, n48063, n48064, n48065, n48066,
         n48067, n48068, n48069, n48070, n48071, n48072, n48073, n48074,
         n48075, n48076, n48077, n48078, n48079, n48080, n48081, n48082,
         n48083, n48084, n48085, n48086, n48087, n48088, n48089, n48090,
         n48091, n48092, n48093, n48094, n48095, n48096, n48097, n48098,
         n48099, n48100, n48101, n48102, n48103, n48104, n48105, n48106,
         n48107, n48108, n48109, n48110, n48111, n48112, n48113, n48114,
         n48115, n48116, n48117, n48118, n48119, n48120, n48121, n48122,
         n48123, n48124, n48125, n48126, n48127, n48128, n48129, n48130,
         n48131, n48132, n48133, n48134, n48135, n48136, n48137, n48138,
         n48139, n48140, n48141, n48142, n48143, n48144, n48145, n48146,
         n48147, n48148, n48149, n48150, n48151, n48152, n48153, n48154,
         n48155, n48156, n48157, n48158, n48159, n48160, n48161, n48162,
         n48163, n48164, n48165, n48166, n48167, n48168, n48169, n48170,
         n48171, n48172, n48173, n48174, n48175, n48176, n48177, n48178,
         n48179, n48180, n48181, n48182, n48183, n48184, n48185, n48186,
         n48187, n48188, n48189, n48190, n48191, n48192, n48193, n48194,
         n48195, n48196, n48197, n48198, n48199, n48200, n48201, n48202,
         n48203, n48204, n48205, n48206, n48207, n48208, n48209, n48210,
         n48211, n48212, n48213, n48214, n48215, n48216, n48217, n48218,
         n48219, n48220, n48221, n48222, n48223, n48224, n48225, n48226,
         n48227, n48228, n48229, n48230, n48231, n48232, n48233, n48234,
         n48235, n48236, n48237, n48238, n48239, n48240, n48241, n48242,
         n48243, n48244, n48245, n48246, n48247, n48248, n48249, n48250,
         n48251, n48252, n48253, n48254, n48255, n48256, n48257, n48258,
         n48259, n48260, n48261, n48262, n48263, n48264, n48265, n48266,
         n48267, n48268, n48269, n48270, n48271, n48272, n48273, n48274,
         n48275, n48276, n48277, n48278, n48279, n48280, n48281, n48282,
         n48283, n48284, n48285, n48286, n48287, n48288, n48289, n48290,
         n48291, n48292, n48293, n48294, n48295, n48296, n48297, n48298,
         n48299, n48300, n48301, n48302, n48303, n48304, n48305, n48306,
         n48307, n48308, n48309, n48310, n48311, n48312, n48313, n48314,
         n48315, n48316, n48317, n48318, n48319, n48320, n48321, n48322,
         n48323, n48324, n48325, n48326, n48327, n48328, n48329, n48330,
         n48331, n48332, n48333, n48334, n48335, n48336, n48337, n48338,
         n48339, n48340, n48341, n48342, n48343, n48344, n48345, n48346,
         n48347, n48348, n48349, n48350, n48351, n48352, n48353, n48354,
         n48355, n48356, n48357, n48358, n48359, n48360, n48361, n48362,
         n48363, n48364, n48365, n48366, n48367, n48368, n48369, n48370,
         n48371, n48372, n48373, n48374, n48375, n48376, n48377, n48378,
         n48379, n48380, n48381, n48382, n48383, n48384, n48385, n48386,
         n48387, n48388, n48389, n48390, n48391, n48392, n48393, n48394,
         n48395, n48396, n48397, n48398, n48399, n48400, n48401, n48402,
         n48403, n48404, n48405, n48406, n48407, n48408, n48409, n48410,
         n48411, n48412, n48413, n48414, n48415, n48416, n48417, n48418,
         n48419, n48420, n48421, n48422, n48423, n48424, n48425, n48426,
         n48427, n48428, n48429, n48430, n48431, n48432, n48433, n48434,
         n48435, n48436, n48437, n48438, n48439, n48440, n48441, n48442,
         n48443, n48444, n48445, n48446, n48447, n48448, n48449, n48450,
         n48451, n48452, n48453, n48454, n48455, n48456, n48457, n48458,
         n48459, n48460, n48461, n48462, n48463, n48464, n48465, n48466,
         n48467, n48468, n48469, n48470, n48471, n48472, n48473, n48474,
         n48475, n48476, n48477, n48478, n48479, n48480, n48481, n48482,
         n48483, n48484, n48485, n48486, n48487, n48488, n48489, n48490,
         n48491, n48492, n48493, n48494, n48495, n48496, n48497, n48498,
         n48499, n48500, n48501, n48502, n48503, n48504, n48505, n48506,
         n48507, n48508, n48509, n48510, n48511, n48512, n48513, n48514,
         n48515, n48516, n48517, n48518, n48519, n48520, n48521, n48522,
         n48523, n48524, n48525, n48526, n48527, n48528, n48529, n48530,
         n48531, n48532, n48533, n48534, n48535, n48536, n48537, n48538,
         n48539, n48540, n48541, n48542, n48543, n48544, n48545, n48546,
         n48547, n48548, n48549, n48550, n48551, n48552, n48553, n48554,
         n48555, n48556, n48557, n48558, n48559, n48560, n48561, n48562,
         n48563, n48564, n48565, n48566, n48567, n48568, n48569, n48570,
         n48571, n48572, n48573, n48574, n48575, n48576, n48577, n48578,
         n48579, n48580, n48581, n48582, n48583, n48584, n48585, n48586,
         n48587, n48588, n48589, n48590, n48591, n48592, n48593, n48594,
         n48595, n48596, n48597, n48598, n48599, n48600, n48601, n48602,
         n48603, n48604, n48605, n48606, n48607, n48608, n48609, n48610,
         n48611, n48612, n48613, n48614, n48615, n48616, n48617, n48618,
         n48619, n48620, n48621, n48622, n48623, n48624, n48625, n48626,
         n48627, n48628, n48629, n48630, n48631, n48632, n48633, n48634,
         n48635, n48636, n48637, n48638, n48639, n48640, n48641, n48642,
         n48643, n48644, n48645, n48646, n48647, n48648, n48649, n48650,
         n48651, n48652, n48653, n48654, n48655, n48656, n48657, n48658,
         n48659, n48660, n48661, n48662, n48663, n48664, n48665, n48666,
         n48667, n48668, n48669, n48670, n48671, n48672, n48673, n48674,
         n48675, n48676, n48677, n48678, n48679, n48680, n48681, n48682,
         n48683, n48684, n48685, n48686, n48687, n48688, n48689, n48690,
         n48691, n48692, n48693, n48694, n48695, n48696, n48697, n48698,
         n48699, n48700, n48701, n48702, n48703, n48704, n48705, n48706,
         n48707, n48708, n48709, n48710, n48711, n48712, n48713, n48714,
         n48715, n48716, n48717, n48718, n48719, n48720, n48721, n48722,
         n48723, n48724, n48725, n48726, n48727, n48728, n48729, n48730,
         n48731, n48732, n48733, n48734, n48735, n48736, n48737, n48738,
         n48739, n48740, n48741, n48742, n48743, n48744, n48745, n48746,
         n48747, n48748, n48749, n48750, n48751, n48752, n48753, n48754,
         n48755, n48756, n48757, n48758, n48759, n48760, n48761, n48762,
         n48763, n48764, n48765, n48766, n48767, n48768, n48769, n48770,
         n48771, n48772, n48773, n48774, n48775, n48776, n48777, n48778,
         n48779, n48780, n48781, n48782, n48783, n48784, n48785, n48786,
         n48787, n48788, n48789, n48790, n48791, n48792, n48793, n48794,
         n48795, n48796, n48797, n48798, n48799, n48800, n48801, n48802,
         n48803, n48804, n48805, n48806, n48807, n48808, n48809, n48810,
         n48811, n48812, n48813, n48814, n48815, n48816, n48817, n48818,
         n48819, n48820, n48821, n48822, n48823, n48824, n48825, n48826,
         n48827, n48828, n48829, n48830, n48831, n48832, n48833, n48834,
         n48835, n48836, n48837, n48838, n48839, n48840, n48841, n48842,
         n48843, n48844, n48845, n48846, n48847, n48848, n48849, n48850,
         n48851, n48852, n48853, n48854, n48855, n48856, n48857, n48858,
         n48859, n48860, n48861, n48862, n48863, n48864, n48865, n48866,
         n48867, n48868, n48869, n48870, n48871, n48872, n48873, n48874,
         n48875, n48876, n48877, n48878, n48879, n48880, n48881, n48882,
         n48883, n48884, n48885, n48886, n48887, n48888, n48889, n48890,
         n48891, n48892, n48893, n48894, n48895, n48896, n48897, n48898,
         n48899, n48900, n48901, n48902, n48903, n48904, n48905, n48906,
         n48907, n48908, n48909, n48910, n48911, n48912, n48913, n48914,
         n48915, n48916, n48917, n48918, n48919, n48920, n48921, n48922,
         n48923, n48924, n48925, n48926, n48927, n48928, n48929, n48930,
         n48931, n48932, n48933, n48934, n48935, n48936, n48937, n48938,
         n48939, n48940, n48941, n48942, n48943, n48944, n48945, n48946,
         n48947, n48948, n48949, n48950, n48951, n48952, n48953, n48954,
         n48955, n48956, n48957, n48958, n48959, n48960, n48961, n48962,
         n48963, n48964, n48965, n48966, n48967, n48968, n48969, n48970,
         n48971, n48972, n48973, n48974, n48975, n48976, n48977, n48978,
         n48979, n48980, n48981, n48982, n48983, n48984, n48985, n48986,
         n48987, n48988, n48989, n48990, n48991, n48992, n48993, n48994,
         n48995, n48996, n48997, n48998, n48999, n49000, n49001, n49002,
         n49003, n49004, n49005, n49006, n49007, n49008, n49009, n49010,
         n49011, n49012, n49013, n49014, n49015, n49016, n49017, n49018,
         n49019, n49020, n49021, n49022, n49023, n49024, n49025, n49026,
         n49027, n49028, n49029, n49030, n49031, n49032, n49033, n49034,
         n49035, n49036, n49037, n49038, n49039, n49040, n49041, n49042,
         n49043, n49044, n49045, n49046, n49047, n49048, n49049, n49050,
         n49051, n49052, n49053, n49054, n49055, n49056, n49057, n49058,
         n49059, n49060, n49061, n49062, n49063, n49064, n49065, n49066,
         n49067, n49068, n49069, n49070, n49071, n49072, n49073, n49074,
         n49075, n49076, n49077, n49078, n49079, n49080, n49081, n49082,
         n49083, n49084, n49085, n49086, n49087, n49088, n49089, n49090,
         n49091, n49092, n49093, n49094, n49095, n49096, n49097, n49098,
         n49099, n49100, n49101, n49102, n49103, n49104, n49105, n49106,
         n49107, n49108, n49109, n49110, n49111, n49112, n49113, n49114,
         n49115, n49116, n49117, n49118, n49119, n49120, n49121, n49122,
         n49123, n49124, n49125, n49126, n49127, n49128, n49129, n49130,
         n49131, n49132, n49133, n49134, n49135, n49136, n49137, n49138,
         n49139, n49140, n49141, n49142, n49143, n49144, n49145, n49146,
         n49147, n49148, n49149, n49150, n49151, n49152, n49153, n49154,
         n49155, n49156, n49157, n49158, n49159, n49160, n49161, n49162,
         n49163, n49164, n49165, n49166, n49167, n49168, n49169, n49170,
         n49171, n49172, n49173, n49174, n49175, n49176, n49177, n49178,
         n49179, n49180, n49181, n49182, n49183, n49184, n49185, n49186,
         n49187, n49188, n49189, n49190, n49191, n49192, n49193, n49194,
         n49195, n49196, n49197, n49198, n49199, n49200, n49201, n49202,
         n49203, n49204, n49205, n49206, n49207, n49208, n49209, n49210,
         n49211, n49212, n49213, n49214, n49215, n49216, n49217, n49218,
         n49219, n49220, n49221, n49222, n49223, n49224, n49225, n49226,
         n49227, n49228, n49229, n49230, n49231, n49232, n49233, n49234,
         n49235, n49236, n49237, n49238, n49239, n49240, n49241, n49242,
         n49243, n49244, n49245, n49246, n49247, n49248, n49249, n49250,
         n49251, n49252, n49253, n49254, n49255, n49256, n49257, n49258,
         n49259, n49260, n49261, n49262, n49263, n49264, n49265, n49266,
         n49267, n49268, n49269, n49270, n49271, n49272, n49273, n49274,
         n49275, n49276, n49277, n49278, n49279, n49280, n49281, n49282,
         n49283, n49284, n49285, n49286, n49287, n49288, n49289, n49290,
         n49291, n49292, n49293, n49294, n49295, n49296, n49297, n49298,
         n49299, n49300, n49301, n49302, n49303, n49304, n49305, n49306,
         n49307, n49308, n49309, n49310, n49311, n49312, n49313, n49314,
         n49315, n49316, n49317, n49318, n49319, n49320, n49321, n49322,
         n49323, n49324, n49325, n49326, n49327, n49328, n49329, n49330,
         n49331, n49332, n49333, n49334, n49335, n49336, n49337, n49338,
         n49339, n49340, n49341, n49342, n49343, n49344, n49345, n49346,
         n49347, n49348, n49349, n49350, n49351, n49352, n49353, n49354,
         n49355, n49356, n49357, n49358, n49359, n49360, n49361, n49362,
         n49363, n49364, n49365, n49366, n49367, n49368, n49369, n49370,
         n49371, n49372, n49373, n49374, n49375, n49376, n49377, n49378,
         n49379, n49380, n49381, n49382, n49383, n49384, n49385, n49386,
         n49387, n49388, n49389, n49390, n49391, n49392, n49393, n49394,
         n49395, n49396, n49397, n49398, n49399, n49400, n49401, n49402,
         n49403, n49404, n49405, n49406, n49407, n49408, n49409, n49410,
         n49411, n49412, n49413, n49414, n49415, n49416, n49417, n49418,
         n49419, n49420, n49421, n49422, n49423, n49424, n49425, n49426,
         n49427, n49428, n49429, n49430, n49431, n49432, n49433, n49434,
         n49435, n49436, n49437, n49438, n49439, n49440, n49441, n49442,
         n49443, n49444, n49445, n49446, n49447, n49448, n49449, n49450,
         n49451, n49452, n49453, n49454, n49455, n49456, n49457, n49458,
         n49459, n49460, n49461, n49462, n49463, n49464, n49465, n49466,
         n49467, n49468, n49469, n49470, n49471, n49472, n49473, n49474,
         n49475, n49476, n49477, n49478, n49479, n49480, n49481, n49482,
         n49483, n49484, n49485, n49486, n49487, n49488, n49489, n49490,
         n49491, n49492, n49493, n49494, n49495, n49496, n49497, n49498,
         n49499, n49500, n49501, n49502, n49503, n49504, n49505, n49506,
         n49507, n49508, n49509, n49510, n49511, n49512, n49513, n49514,
         n49515, n49516, n49517, n49518, n49519, n49520, n49521, n49522,
         n49523, n49524, n49525, n49526, n49527, n49528, n49529, n49530,
         n49531, n49532, n49533, n49534, n49535, n49536, n49537, n49538,
         n49539, n49540, n49541, n49542, n49543, n49544, n49545, n49546,
         n49547, n49548, n49549, n49550, n49551, n49552, n49553, n49554,
         n49555, n49556, n49557, n49558, n49559, n49560, n49561, n49562,
         n49563, n49564, n49565, n49566, n49567, n49568, n49569, n49570,
         n49571, n49572, n49573, n49574, n49575, n49576, n49577, n49578,
         n49579, n49580, n49581, n49582, n49583, n49584, n49585, n49586,
         n49587, n49588, n49589, n49590, n49591, n49592, n49593, n49594,
         n49595, n49596, n49597, n49598, n49599, n49600, n49601, n49602,
         n49603, n49604, n49605, n49606, n49607, n49608, n49609, n49610,
         n49611, n49612, n49613, n49614, n49615, n49616, n49617, n49618,
         n49619, n49620, n49621, n49622, n49623, n49624, n49625, n49626,
         n49627, n49628, n49629, n49630, n49631, n49632, n49633, n49634,
         n49635, n49636, n49637, n49638, n49639, n49640, n49641, n49642,
         n49643, n49644, n49645, n49646, n49647, n49648, n49649, n49650,
         n49651, n49652, n49653, n49654, n49655, n49656, n49657, n49658,
         n49659, n49660, n49661, n49662, n49663, n49664, n49665, n49666,
         n49667, n49668, n49669, n49670, n49671, n49672, n49673, n49674,
         n49675, n49676, n49677, n49678, n49679, n49680, n49681, n49682,
         n49683, n49684, n49685, n49686, n49687, n49688, n49689, n49690,
         n49691, n49692, n49693, n49694, n49695, n49696, n49697, n49698,
         n49699, n49700, n49701, n49702, n49703, n49704, n49705, n49706,
         n49707, n49708, n49709, n49710, n49711, n49712, n49713, n49714,
         n49715, n49716, n49717, n49718, n49719, n49720, n49721, n49722,
         n49723, n49724, n49725, n49726, n49727, n49728, n49729, n49730,
         n49731, n49732, n49733, n49734, n49735, n49736, n49737, n49738,
         n49739, n49740, n49741, n49742, n49743, n49744, n49745, n49746,
         n49747, n49748, n49749, n49750, n49751, n49752, n49753, n49754,
         n49755, n49756, n49757, n49758, n49759, n49760, n49761, n49762,
         n49763, n49764, n49765, n49766, n49767, n49768, n49769, n49770,
         n49771, n49772, n49773, n49774, n49775, n49776, n49777, n49778,
         n49779, n49780, n49781, n49782, n49783, n49784, n49785, n49786,
         n49787, n49788, n49789, n49790, n49791, n49792, n49793, n49794,
         n49795, n49796, n49797, n49798, n49799, n49800, n49801, n49802,
         n49803, n49804, n49805, n49806, n49807, n49808, n49809, n49810,
         n49811, n49812, n49813, n49814, n49815, n49816, n49817, n49818,
         n49819, n49820, n49821, n49822, n49823, n49824, n49825, n49826,
         n49827, n49828, n49829, n49830, n49831, n49832, n49833, n49834,
         n49835, n49836, n49837, n49838, n49839, n49840, n49841, n49842,
         n49843, n49844, n49845, n49846, n49847, n49848, n49849, n49850,
         n49851, n49852, n49853, n49854, n49855, n49856, n49857, n49858,
         n49859, n49860, n49861, n49862, n49863, n49864, n49865, n49866,
         n49867, n49868, n49869, n49870, n49871, n49872, n49873, n49874,
         n49875, n49876, n49877, n49878, n49879, n49880, n49881, n49882,
         n49883, n49884, n49885, n49886, n49887, n49888, n49889, n49890,
         n49891, n49892, n49893, n49894, n49895, n49896, n49897, n49898,
         n49899, n49900, n49901, n49902, n49903, n49904, n49905, n49906,
         n49907, n49908, n49909, n49910, n49911, n49912, n49913, n49914,
         n49915, n49916, n49917, n49918, n49919, n49920, n49921, n49922,
         n49923, n49924, n49925, n49926, n49927, n49928, n49929, n49930,
         n49931, n49932, n49933, n49934, n49935, n49936, n49937, n49938,
         n49939, n49940, n49941, n49942, n49943, n49944, n49945, n49946,
         n49947, n49948, n49949, n49950, n49951, n49952, n49953, n49954,
         n49955, n49956, n49957, n49958, n49959, n49960, n49961, n49962,
         n49963, n49964, n49965, n49966, n49967, n49968, n49969, n49970,
         n49971, n49972, n49973, n49974, n49975, n49976, n49977, n49978,
         n49979, n49980, n49981, n49982, n49983, n49984, n49985, n49986,
         n49987, n49988, n49989, n49990, n49991, n49992, n49993, n49994,
         n49995, n49996, n49997, n49998, n49999, n50000, n50001, n50002,
         n50003, n50004, n50005, n50006, n50007, n50008, n50009, n50010,
         n50011, n50012, n50013, n50014, n50015, n50016, n50017, n50018,
         n50019, n50020, n50021, n50022, n50023, n50024, n50025, n50026,
         n50027, n50028, n50029, n50030, n50031, n50032, n50033, n50034,
         n50035, n50036, n50037, n50038, n50039, n50040, n50041, n50042,
         n50043, n50044, n50045, n50046, n50047, n50048, n50049, n50050,
         n50051, n50052, n50053, n50054, n50055, n50056, n50057, n50058,
         n50059, n50060, n50061, n50062, n50063, n50064, n50065, n50066,
         n50067, n50068, n50069, n50070, n50071, n50072, n50073, n50074,
         n50075, n50076, n50077, n50078, n50079, n50080, n50081, n50082,
         n50083, n50084, n50085, n50086, n50087, n50088, n50089, n50090,
         n50091, n50092, n50093, n50094, n50095, n50096, n50097, n50098,
         n50099, n50100, n50101, n50102, n50103, n50104, n50105, n50106,
         n50107, n50108, n50109, n50110, n50111, n50112, n50113, n50114,
         n50115, n50116, n50117, n50118, n50119, n50120, n50121, n50122,
         n50123, n50124, n50125, n50126, n50127, n50128, n50129, n50130,
         n50131, n50132, n50133, n50134, n50135, n50136, n50137, n50138,
         n50139, n50140, n50141, n50142, n50143, n50144, n50145, n50146,
         n50147, n50148, n50149, n50150, n50151, n50152, n50153, n50154,
         n50155, n50156, n50157, n50158, n50159, n50160, n50161, n50162,
         n50163, n50164, n50165, n50166, n50167, n50168, n50169, n50170,
         n50171, n50172, n50173, n50174, n50175, n50176, n50177, n50178,
         n50179, n50180, n50181, n50182, n50183, n50184, n50185, n50186,
         n50187, n50188, n50189, n50190, n50191, n50192, n50193, n50194,
         n50195, n50196, n50197, n50198, n50199, n50200, n50201, n50202,
         n50203, n50204, n50205, n50206, n50207, n50208, n50209, n50210,
         n50211, n50212, n50213, n50214, n50215, n50216, n50217, n50218,
         n50219, n50220, n50221, n50222, n50223, n50224, n50225, n50226,
         n50227, n50228, n50229, n50230, n50231, n50232, n50233, n50234,
         n50235, n50236, n50237, n50238, n50239, n50240, n50241, n50242,
         n50243, n50244, n50245, n50246, n50247, n50248, n50249, n50250,
         n50251, n50252, n50253, n50254, n50255, n50256, n50257, n50258,
         n50259, n50260, n50261, n50262, n50263, n50264, n50265, n50266,
         n50267, n50268, n50269, n50270, n50271, n50272, n50273, n50274,
         n50275, n50276, n50277, n50278, n50279, n50280, n50281, n50282,
         n50283, n50284, n50285, n50286, n50287, n50288, n50289, n50290,
         n50291, n50292, n50293, n50294, n50295, n50296, n50297, n50298,
         n50299, n50300, n50301, n50302, n50303, n50304, n50305, n50306,
         n50307, n50308, n50309, n50310, n50311, n50312, n50313, n50314,
         n50315, n50316, n50317, n50318, n50319, n50320, n50321, n50322,
         n50323, n50324, n50325, n50326, n50327, n50328, n50329, n50330,
         n50331, n50332, n50333, n50334, n50335, n50336, n50337, n50338,
         n50339, n50340, n50341, n50342, n50343, n50344, n50345, n50346,
         n50347, n50348, n50349, n50350, n50351, n50352, n50353, n50354,
         n50355, n50356, n50357, n50358, n50359, n50360, n50361, n50362,
         n50363, n50364, n50365, n50366, n50367, n50368, n50369, n50370,
         n50371, n50372, n50373, n50374, n50375, n50376, n50377, n50378,
         n50379, n50380, n50381, n50382, n50383, n50384, n50385, n50386,
         n50387, n50388, n50389, n50390, n50391, n50392, n50393, n50394,
         n50395, n50396, n50397, n50398, n50399, n50400, n50401, n50402,
         n50403, n50404, n50405, n50406, n50407, n50408, n50409, n50410,
         n50411, n50412, n50413, n50414, n50415, n50416, n50417, n50418,
         n50419, n50420, n50421, n50422, n50423, n50424, n50425, n50426,
         n50427, n50428, n50429, n50430, n50431, n50432, n50433, n50434,
         n50435, n50436, n50437, n50438, n50439, n50440, n50441, n50442,
         n50443, n50444, n50445, n50446, n50447, n50448, n50449, n50450,
         n50451, n50452, n50453, n50454, n50455, n50456, n50457, n50458,
         n50459, n50460, n50461, n50462, n50463, n50464, n50465, n50466,
         n50467, n50468, n50469, n50470, n50471, n50472, n50473, n50474,
         n50475, n50476, n50477, n50478, n50479, n50480, n50481, n50482,
         n50483, n50484, n50485, n50486, n50487, n50488, n50489, n50490,
         n50491, n50492, n50493, n50494, n50495, n50496, n50497, n50498,
         n50499, n50500, n50501, n50502, n50503, n50504, n50505, n50506,
         n50507, n50508, n50509, n50510, n50511, n50512, n50513, n50514,
         n50515, n50516, n50517, n50518, n50519, n50520, n50521, n50522,
         n50523, n50524, n50525, n50526, n50527, n50528, n50529, n50530,
         n50531, n50532, n50533, n50534, n50535, n50536, n50537, n50538,
         n50539, n50540, n50541, n50542, n50543, n50544, n50545, n50546,
         n50547, n50548, n50549, n50550, n50551, n50552, n50553, n50554,
         n50555, n50556, n50557, n50558, n50559, n50560, n50561, n50562,
         n50563, n50564, n50565, n50566, n50567, n50568, n50569, n50570,
         n50571, n50572, n50573, n50574, n50575, n50576, n50577, n50578,
         n50579, n50580, n50581, n50582, n50583, n50584, n50585, n50586,
         n50587, n50588, n50589, n50590, n50591, n50592, n50593, n50594,
         n50595, n50596, n50597, n50598, n50599, n50600, n50601, n50602,
         n50603, n50604, n50605, n50606, n50607, n50608, n50609, n50610,
         n50611, n50612, n50613, n50614, n50615, n50616, n50617, n50618,
         n50619, n50620, n50621, n50622, n50623, n50624, n50625, n50626,
         n50627, n50628, n50629, n50630, n50631, n50632, n50633, n50634,
         n50635, n50636, n50637, n50638, n50639, n50640, n50641, n50642,
         n50643, n50644, n50645, n50646, n50647, n50648, n50649, n50650,
         n50651, n50652, n50653, n50654, n50655, n50656, n50657, n50658,
         n50659, n50660, n50661, n50662, n50663, n50664, n50665, n50666,
         n50667, n50668, n50669, n50670, n50671, n50672, n50673, n50674,
         n50675, n50676, n50677, n50678, n50679, n50680, n50681, n50682,
         n50683, n50684, n50685, n50686, n50687, n50688, n50689, n50690,
         n50691, n50692, n50693, n50694, n50695, n50696, n50697, n50698,
         n50699, n50700, n50701, n50702, n50703, n50704, n50705, n50706,
         n50707, n50708, n50709, n50710, n50711, n50712, n50713, n50714,
         n50715, n50716, n50717, n50718, n50719, n50720, n50721, n50722,
         n50723, n50724, n50725, n50726, n50727, n50728, n50729, n50730,
         n50731, n50732, n50733, n50734, n50735, n50736, n50737, n50738,
         n50739, n50740, n50741, n50742, n50743, n50744, n50745, n50746,
         n50747, n50748, n50749, n50750, n50751, n50752, n50753, n50754,
         n50755, n50756, n50757, n50758, n50759, n50760, n50761, n50762,
         n50763, n50764, n50765, n50766, n50767, n50768, n50769, n50770,
         n50771, n50772, n50773, n50774, n50775, n50776, n50777, n50778,
         n50779, n50780, n50781, n50782, n50783, n50784, n50785, n50786,
         n50787, n50788, n50789, n50790, n50791, n50792, n50793, n50794,
         n50795, n50796, n50797, n50798, n50799, n50800, n50801, n50802,
         n50803, n50804, n50805, n50806, n50807, n50808, n50809, n50810,
         n50811, n50812, n50813, n50814, n50815, n50816, n50817, n50818,
         n50819, n50820, n50821, n50822, n50823, n50824, n50825, n50826,
         n50827, n50828, n50829, n50830, n50831, n50832, n50833, n50834,
         n50835, n50836, n50837, n50838, n50839, n50840, n50841, n50842,
         n50843, n50844, n50845, n50846, n50847, n50848, n50849, n50850,
         n50851, n50852, n50853, n50854, n50855, n50856, n50857, n50858,
         n50859, n50860, n50861, n50862, n50863, n50864, n50865, n50866,
         n50867, n50868, n50869, n50870, n50871, n50872, n50873, n50874,
         n50875, n50876, n50877, n50878, n50879, n50880, n50881, n50882,
         n50883, n50884, n50885, n50886, n50887, n50888, n50889, n50890,
         n50891, n50892, n50893, n50894, n50895, n50896, n50897, n50898,
         n50899, n50900, n50901, n50902, n50903, n50904, n50905, n50906,
         n50907, n50908, n50909, n50910, n50911, n50912, n50913, n50914,
         n50915, n50916, n50917, n50918, n50919, n50920, n50921, n50922,
         n50923, n50924, n50925, n50926, n50927, n50928, n50929, n50930,
         n50931, n50932, n50933, n50934, n50935, n50936, n50937, n50938,
         n50939, n50940, n50941, n50942, n50943, n50944, n50945, n50946,
         n50947, n50948, n50949, n50950, n50951, n50952, n50953, n50954,
         n50955, n50956, n50957, n50958, n50959, n50960, n50961, n50962,
         n50963, n50964, n50965, n50966, n50967, n50968, n50969, n50970,
         n50971, n50972, n50973, n50974, n50975, n50976, n50977, n50978,
         n50979, n50980, n50981, n50982, n50983, n50984, n50985, n50986,
         n50987, n50988, n50989, n50990, n50991, n50992, n50993, n50994,
         n50995, n50996, n50997, n50998, n50999, n51000, n51001, n51002,
         n51003, n51004, n51005, n51006, n51007, n51008, n51009, n51010,
         n51011, n51012, n51013, n51014, n51015, n51016, n51017, n51018,
         n51019, n51020, n51021, n51022, n51023, n51024, n51025, n51026,
         n51027, n51028, n51029, n51030, n51031, n51032, n51033, n51034,
         n51035, n51036, n51037, n51038, n51039, n51040, n51041, n51042,
         n51043, n51044, n51045, n51046, n51047, n51048, n51049, n51050,
         n51051, n51052, n51053, n51054, n51055, n51056, n51057, n51058,
         n51059, n51060, n51061, n51062, n51063, n51064, n51065, n51066,
         n51067, n51068, n51069, n51070, n51071, n51072, n51073, n51074,
         n51075, n51076, n51077, n51078, n51079, n51080, n51081, n51082,
         n51083, n51084, n51085, n51086, n51087, n51088, n51089, n51090,
         n51091, n51092, n51093, n51094, n51095, n51096, n51097, n51098,
         n51099, n51100, n51101, n51102, n51103, n51104, n51105, n51106,
         n51107, n51108, n51109, n51110, n51111, n51112, n51113, n51114,
         n51115, n51116, n51117, n51118, n51119, n51120, n51121, n51122,
         n51123, n51124, n51125, n51126, n51127, n51128, n51129, n51130,
         n51131, n51132, n51133, n51134, n51135, n51136, n51137, n51138,
         n51139, n51140, n51141, n51142, n51143, n51144, n51145, n51146,
         n51147, n51148, n51149, n51150, n51151, n51152, n51153, n51154,
         n51155, n51156, n51157, n51158, n51159, n51160, n51161, n51162,
         n51163, n51164, n51165, n51166, n51167, n51168, n51169, n51170,
         n51171, n51172, n51173, n51174, n51175, n51176, n51177, n51178,
         n51179, n51180, n51181, n51182, n51183, n51184, n51185, n51186,
         n51187, n51188, n51189, n51190, n51191, n51192, n51193, n51194,
         n51195, n51196, n51197, n51198, n51199, n51200, n51201, n51202,
         n51203, n51204, n51205, n51206, n51207, n51208, n51209, n51210,
         n51211, n51212, n51213, n51214, n51215, n51216, n51217, n51218,
         n51219, n51220, n51221, n51222, n51223, n51224, n51225, n51226,
         n51227, n51228, n51229, n51230, n51231, n51232, n51233, n51234,
         n51235, n51236, n51237, n51238, n51239, n51240, n51241, n51242,
         n51243, n51244, n51245, n51246, n51247, n51248, n51249, n51250,
         n51251, n51252, n51253, n51254, n51255, n51256, n51257, n51258,
         n51259, n51260, n51261, n51262, n51263, n51264, n51265, n51266,
         n51267, n51268, n51269, n51270, n51271, n51272, n51273, n51274,
         n51275, n51276, n51277, n51278, n51279, n51280, n51281, n51282,
         n51283, n51284, n51285, n51286, n51287, n51288, n51289, n51290,
         n51291, n51292, n51293, n51294, n51295, n51296, n51297, n51298,
         n51299, n51300, n51301, n51302, n51303, n51304, n51305, n51306,
         n51307, n51308, n51309, n51310, n51311, n51312, n51313, n51314,
         n51315, n51316, n51317, n51318, n51319, n51320, n51321, n51322,
         n51323, n51324, n51325, n51326, n51327, n51328, n51329, n51330,
         n51331, n51332, n51333, n51334, n51335, n51336, n51337, n51338,
         n51339, n51340, n51341, n51342, n51343, n51344, n51345, n51346,
         n51347, n51348, n51349, n51350, n51351, n51352, n51353, n51354,
         n51355, n51356, n51357, n51358, n51359, n51360, n51361, n51362,
         n51363, n51364, n51365, n51366, n51367, n51368, n51369, n51370,
         n51371, n51372, n51373, n51374, n51375, n51376, n51377, n51378,
         n51379, n51380, n51381, n51382, n51383, n51384, n51385, n51386,
         n51387, n51388, n51389, n51390, n51391, n51392, n51393, n51394,
         n51395, n51396, n51397, n51398, n51399, n51400, n51401, n51402,
         n51403, n51404, n51405, n51406, n51407, n51408, n51409, n51410,
         n51411, n51412, n51413, n51414, n51415, n51416, n51417, n51418,
         n51419, n51420, n51421, n51422, n51423, n51424, n51425, n51426,
         n51427, n51428, n51429, n51430, n51431, n51432, n51433, n51434,
         n51435, n51436, n51437, n51438, n51439, n51440, n51441, n51442,
         n51443, n51444, n51445, n51446, n51447, n51448, n51449, n51450,
         n51451, n51452, n51453, n51454, n51455, n51456, n51457, n51458,
         n51459, n51460, n51461, n51462, n51463, n51464, n51465, n51466,
         n51467, n51468, n51469, n51470, n51471, n51472, n51473, n51474,
         n51475, n51476, n51477, n51478, n51479, n51480, n51481, n51482,
         n51483, n51484, n51485, n51486, n51487, n51488, n51489, n51490,
         n51491, n51492, n51493, n51494, n51495, n51496, n51497, n51498,
         n51499, n51500, n51501, n51502, n51503, n51504, n51505, n51506,
         n51507, n51508, n51509, n51510, n51511, n51512, n51513, n51514,
         n51515, n51516, n51517, n51518, n51519, n51520, n51522, n51523,
         n51524, n51525, n51526, n51527, n51528, n51529, n51530, n51531,
         n51532, n51533, n51534, n51535, n51536, n51537, n51538, n51539,
         n51540, n51541, n51542, n51543, n51544, n51545, n51546, n51547,
         n51548, n51549, n51550, n51551, n51552, n51553, n51554, n51555,
         n51556, n51557, n51558, n51560, n51561, n51562, n51563, n51564,
         n51565, n51566, n51567, n51568, n51569, n51570, n51571, n51572,
         n51573, n51574, n51575, n51576, n51577, n51578, n51579, n51580,
         n51581, n51582, n51583, n51584, n51585, n51586, n51587, n51588,
         n51589, n51590, n51591, n51592, n51593, n51594, n51595, n51596,
         n51597, n51598, n51599, n51600, n51601, n51602, n51603, n51604,
         n51605, n51606, n51607, n51608, n51609, n51610, n51611, n51612,
         n51613, n51614, n51615, n51616, n51617, n51618, n51619, n51620,
         n51621, n51622, n51623, n51624, n51625, n51626, n51627, n51628,
         n51629, n51630, n51631, n51632, n51633, n51634, n51635, n51636,
         n51637, n51638, n51639, n51640, n51641, n51642, n51643, n51644,
         n51645, n51646, n51647, n51648, n51649, n51650, n51651, n51652,
         n51653, n51654, n51655, n51656, n51657, n51658, n51659, n51660,
         n51661, n51662, n51663, n51664, n51665, n51666, n51667, n51668,
         n51669, n51670, n51671, n51672, n51673, n51674, n51675, n51676,
         n51677, n51678, n51679, n51680, n51681, n51682, n51683, n51684,
         n51685, n51686, n51687, n51688, n51689, n51690, n51691, n51692,
         n51693, n51694, n51695, n51696, n51697, n51698, n51699, n51700,
         n51701, n51702, n51703, n51704, n51705, n51706, n51707, n51708,
         n51709, n51710, n51711, n51712, n51713, n51714, n51715, n51716,
         n51717, n51718, n51719, n51720, n51721, n51722, n51723, n51724,
         n51725, n51726, n51727, n51728, n51729, n51730, n51731, n51732,
         n51733, n51734, n51735, n51736, n51737, n51738, n51739, n51740,
         n51741, n51742, n51743, n51744, n51745, n51746, n51747, n51748,
         n51749, n51750, n51751, n51752, n51753, n51754, n51755, n51756,
         n51757, n51758, n51759, n51760, n51761, n51762, n51763, n51764,
         n51765, n51766, n51767, n51768, n51769, n51770, n51771, n51772,
         n51773, n51774, n51775, n51776, n51777, n51778, n51779, n51780,
         n51781, n51782, n51783, n51784, n51785, n51786, n51787, n51788,
         n51789, n51790, n51791, n51792, n51793, n51794, n51795, n51796,
         n51797, n51798, n51799, n51800, n51801, n51802, n51803, n51804,
         n51805, n51806, n51807, n51808, n51809, n51810, n51811, n51812,
         n51813, n51814, n51815, n51816, n51817, n51818, n51819, n51820,
         n51821, n51822, n51823, n51824, n51825, n51826, n51827, n51828,
         n51829, n51830, n51831, n51832, n51833, n51834, n51835, n51836,
         n51837, n51838, n51839, n51840, n51841, n51842, n51843, n51844,
         n51845, n51846, n51847, n51848, n51849, n51850, n51851, n51852,
         n51853, n51854, n51855, n51856, n51857, n51858, n51859, n51860,
         n51861, n51862, n51863, n51864, n51865, n51866, n51867, n51868,
         n51869, n51870, n51871, n51872, n51873, n51874, n51875, n51876,
         n51877, n51878, n51879, n51880, n51881, n51882, n51883, n51884,
         n51885, n51886, n51887, n51888, n51889, n51890, n51891, n51892,
         n51893, n51894, n51895, n51896, n51897, n51898, n51899, n51900,
         n51901, n51902, n51903, n51904, n51905, n51906, n51907, n51908,
         n51909, n51910, n51911, n51912, n51913, n51914, n51915, n51916,
         n51917, n51918, n51919, n51920, n51921, n51922, n51923, n51924,
         n51925, n51926, n51927, n51928, n51929, n51930, n51931, n51932,
         n51933, n51934, n51935, n51936, n51937, n51938, n51939, n51940,
         n51941, n51942, n51943, n51944, n51945, n51946, n51947, n51948,
         n51949, n51950, n51951, n51952, n51953, n51954, n51955, n51956,
         n51957, n51958, n51959, n51960, n51961, n51962, n51963, n51964,
         n51965, n51966, n51967, n51968, n51969, n51970, n51971, n51972,
         n51973, n51974, n51975, n51976, n51977, n51978, n51979, n51980,
         n51981, n51982, n51983, n51984, n51985, n51986, n51987, n51988,
         n51989, n51990, n51991, n51992, n51993, n51994, n51995, n51996,
         n51997, n51998, n51999, n52000, n52001, n52002, n52003, n52004,
         n52005, n52006, n52007, n52008, n52009, n52010, n52011, n52012,
         n52013, n52014, n52015, n52016, n52017, n52018, n52019, n52020,
         n52021, n52022, n52023, n52024, n52025, n52026, n52027, n52028,
         n52029, n52030, n52031, n52032, n52033, n52034, n52035, n52036,
         n52037, n52038, n52039, n52040, n52041, n52042, n52043, n52044,
         n52045, n52046, n52047, n52048, n52049, n52050, n52051, n52052,
         n52053, n52054, n52055, n52056, n52057, n52058, n52059, n52060,
         n52061, n52062, n52063, n52064, n52065, n52066, n52067, n52068,
         n52069, n52070, n52071, n52072, n52073, n52074, n52075, n52076,
         n52077, n52078, n52079, n52080, n52081, n52082, n52083, n52084,
         n52085, n52086, n52087, n52088, n52089, n52090, n52091, n52092,
         n52093, n52094, n52095, n52096, n52097, n52098, n52099, n52100,
         n52101, n52102, n52103, n52104, n52105, n52106, n52107, n52108,
         n52109, n52110, n52111, n52112, n52113, n52114, n52115, n52116,
         n52117, n52118, n52119, n52120, n52121, n52122, n52123, n52124,
         n52125, n52126, n52127, n52128, n52129, n52130, n52131, n52132,
         n52133, n52134, n52135, n52136, n52137, n52138, n52139, n52140,
         n52141, n52142, n52143, n52144, n52145, n52146, n52147, n52148,
         n52149, n52150, n52151, n52152, n52153, n52154, n52155, n52156,
         n52157, n52158, n52159, n52160, n52161, n52162, n52163, n52164,
         n52165, n52166, n52167, n52168, n52169, n52170, n52171, n52172,
         n52173, n52174, n52175, n52176, n52177, n52178, n52179, n52180,
         n52181, n52182, n52183, n52184, n52185, n52186, n52187, n52188,
         n52189, n52190, n52191, n52192, n52193, n52194, n52195, n52196,
         n52197, n52198, n52199, n52200, n52201, n52202, n52203, n52204,
         n52205, n52206, n52207, n52208, n52209, n52210, n52211, n52212,
         n52213, n52214, n52215, n52216, n52217, n52218, n52219, n52220,
         n52221, n52222, n52223, n52224, n52225, n52226, n52227, n52228,
         n52229, n52230, n52231, n52232, n52233, n52234, n52235, n52236,
         n52237, n52238, n52239, n52240, n52241, n52242, n52243, n52244,
         n52245, n52246, n52247, n52248, n52249, n52250, n52251, n52252,
         n52253, n52254, n52255, n52256, n52257, n52258, n52259, n52260,
         n52261, n52262, n52263, n52264, n52265, n52266, n52267, n52268,
         n52269, n52270, n52271, n52272, n52273, n52274, n52275, n52276,
         n52277, n52278, n52279, n52280, n52281, n52282, n52283, n52284,
         n52285, n52286, n52287, n52288, n52289, n52290, n52291, n52292,
         n52293, n52294, n52295, n52296, n52297, n52298, n52299, n52300,
         n52301, n52302, n52303, n52304, n52305, n52306, n52307, n52308,
         n52309, n52310, n52311, n52312, n52313, n52314, n52315, n52316,
         n52317, n52318, n52319, n52320, n52321, n52322, n52323, n52324,
         n52325, n52326, n52327, n52328, n52329, n52330, n52331, n52332,
         n52333, n52334, n52335, n52336, n52337, n52338, n52339, n52340,
         n52341, n52342, n52343, n52344, n52345, n52346, n52347, n52348,
         n52349, n52350, n52351, n52352, n52353, n52354, n52355, n52356,
         n52357, n52358, n52359, n52360, n52361, n52362, n52363, n52364,
         n52365, n52366, n52367, n52368, n52369, n52370, n52371, n52372,
         n52373, n52374, n52375, n52376, n52377, n52378, n52379, n52380,
         n52381, n52382, n52383, n52384, n52385, n52386, n52387, n52388,
         n52389, n52390, n52391, n52392, n52393, n52394, n52395, n52396,
         n52397, n52398, n52399, n52400, n52401, n52402, n52403, n52404,
         n52405, n52406, n52407, n52408, n52409, n52410, n52411, n52412,
         n52413, n52414, n52415, n52416, n52417, n52418, n52419, n52420,
         n52421, n52422, n52423, n52424, n52425, n52426, n52427, n52428,
         n52429, n52430, n52431, n52432, n52433, n52434, n52435, n52436,
         n52437, n52438, n52439, n52440, n52441, n52442, n52443, n52444,
         n52445, n52446, n52447, n52448, n52449, n52450, n52451, n52452,
         n52453, n52454, n52455, n52456, n52457, n52458, n52459, n52460,
         n52461, n52462, n52463, n52464, n52465, n52466, n52467, n52468,
         n52469, n52470, n52471, n52472, n52473, n52474, n52475, n52476,
         n52477, n52478, n52479, n52480, n52481, n52482, n52483, n52484,
         n52485, n52486, n52487, n52488, n52489, n52490, n52491, n52492,
         n52493, n52494, n52495, n52496, n52497, n52498, n52499, n52500,
         n52501, n52502, n52503, n52504, n52505, n52506, n52507, n52508,
         n52509, n52510, n52511, n52512, n52513, n52514, n52515, n52516,
         n52517, n52518, n52519, n52520, n52521, n52522, n52523, n52524,
         n52525, n52526, n52527, n52528, n52529, n52530, n52531, n52532,
         n52533, n52534, n52535, n52536, n52537, n52538, n52539, n52540,
         n52541, n52542, n52543, n52544, n52545, n52546, n52547, n52548,
         n52549, n52550, n52551, n52552, n52553, n52554, n52555, n52556,
         n52557, n52558, n52559, n52560, n52561, n52562, n52563, n52564,
         n52565, n52566, n52567, n52568, n52569, n52570, n52571, n52572,
         n52573, n52574, n52575, n52576, n52577, n52578, n52579, n52580,
         n52581, n52582, n52583, n52584, n52585, n52586, n52587, n52588,
         n52589, n52590, n52591, n52592, n52593, n52594, n52595, n52596,
         n52597, n52598, n52599, n52600, n52601, n52602, n52603, n52604,
         n52605, n52606, n52607, n52608, n52609, n52610, n52611, n52612,
         n52613, n52614, n52615, n52616, n52617, n52618, n52619, n52620,
         n52621, n52622, n52623, n52624, n52625, n52626, n52627, n52628,
         n52629, n52630, n52631, n52632, n52633, n52634, n52635, n52636,
         n52637, n52638, n52639, n52640, n52641, n52642, n52643, n52644,
         n52645, n52646, n52647, n52648, n52649, n52650, n52651, n52652,
         n52653, n52654, n52655, n52656, n52657, n52658, n52659, n52660,
         n52661, n52662, n52663, n52664, n52665, n52666, n52667, n52668,
         n52669, n52670, n52671, n52672, n52673, n52674, n52675, n52676,
         n52677, n52678, n52679, n52680, n52681, n52682, n52683, n52684,
         n52685, n52686, n52687, n52688, n52689, n52690, n52691, n52692,
         n52693, n52694, n52695, n52696, n52697, n52698, n52699, n52700,
         n52701, n52702, n52703, n52704, n52705, n52706, n52707, n52708,
         n52709, n52710, n52711, n52712, n52713, n52714, n52715, n52716,
         n52717, n52718, n52719, n52720, n52721, n52722, n52723, n52724,
         n52725, n52726, n52727, n52728, n52729, n52730, n52731, n52732,
         n52733, n52734, n52735, n52736, n52737, n52738, n52739, n52740,
         n52741, n52742, n52743, n52744, n52745, n52746, n52747, n52748,
         n52749, n52750, n52751, n52752, n52753, n52754, n52755, n52756,
         n52757, n52758, n52759, n52760, n52761, n52762, n52763, n52764,
         n52765, n52766, n52767, n52768, n52769, n52770, n52771, n52772,
         n52773, n52774, n52775, n52776, n52777, n52778, n52779, n52780,
         n52781, n52782, n52783, n52784, n52785, n52786, n52787, n52788,
         n52789, n52790, n52791, n52792, n52793, n52794, n52795, n52796,
         n52797, n52798, n52799, n52800, n52801, n52802, n52803, n52804,
         n52805, n52806, n52807, n52808, n52809, n52810, n52811, n52812,
         n52813, n52814, n52815, n52816, n52817, n52818, n52819, n52820,
         n52821, n52822, n52823, n52824, n52825, n52826, n52827, n52828,
         n52829, n52830, n52831, n52832, n52833, n52834, n52835, n52836,
         n52837, n52838, n52839, n52840, n52841, n52842, n52843, n52844,
         n52845, n52846, n52847, n52848, n52849, n52850, n52851, n52852,
         n52853, n52854, n52855, n52856, n52857, n52858, n52859, n52860,
         n52861, n52862, n52863, n52864, n52865, n52866, n52867, n52868,
         n52869, n52870, n52871, n52872, n52873, n52874, n52875, n52876,
         n52877, n52878, n52879, n52880, n52881, n52882, n52883, n52884,
         n52885, n52886, n52887, n52888, n52889, n52890, n52891, n52892,
         n52893, n52894, n52895, n52896, n52897, n52898, n52899, n52900,
         n52901, n52902, n52903, n52904, n52905, n52906, n52907, n52908,
         n52909, n52910, n52911, n52912, n52913, n52914, n52915, n52916,
         n52917, n52918, n52919, n52920, n52921, n52922, n52923, n52924,
         n52925, n52926, n52927, n52928, n52929, n52930, n52931, n52932,
         n52933, n52934, n52935, n52936, n52937, n52938, n52939, n52940,
         n52941, n52942, n52943, n52944, n52945, n52946, n52947, n52948,
         n52949, n52950, n52951, n52952, n52953, n52954, n52955, n52956,
         n52957, n52958, n52959, n52960, n52961, n52962, n52963, n52964,
         n52965, n52966, n52967, n52968, n52969, n52970, n52971, n52972,
         n52973, n52974, n52975, n52976, n52977, n52978, n52979, n52980,
         n52981, n52982, n52983, n52984, n52985, n52986, n52987, n52988,
         n52989, n52990, n52991, n52992, n52993, n52994, n52995, n52996,
         n52997, n52998, n52999, n53000, n53001, n53002, n53003, n53004,
         n53005, n53006, n53007, n53008, n53009, n53010, n53011, n53012,
         n53013, n53014, n53015, n53016, n53017, n53018, n53019, n53020,
         n53021, n53022, n53023, n53024, n53025, n53026, n53027, n53028,
         n53029, n53030, n53031, n53032, n53033, n53034, n53035, n53036,
         n53037, n53038, n53039, n53040, n53041, n53042, n53043, n53044,
         n53045, n53046, n53047, n53048, n53049, n53050, n53051, n53052,
         n53053, n53054, n53055, n53056, n53057, n53058, n53059, n53060,
         n53061, n53062, n53063, n53064, n53065, n53066, n53067, n53068,
         n53069, n53070, n53071, n53072, n53073, n53074, n53075, n53076,
         n53077, n53078, n53079, n53080, n53081, n53082, n53083, n53084,
         n53085, n53086, n53087, n53088, n53089, n53090, n53091, n53092,
         n53093, n53094, n53095, n53096, n53097, n53098, n53099, n53100,
         n53101, n53102, n53103, n53104, n53105, n53106, n53107, n53108,
         n53109, n53110, n53111, n53112, n53113, n53114, n53115, n53116,
         n53117, n53118, n53119, n53120, n53121, n53122, n53123, n53124,
         n53125, n53126, n53127, n53128, n53129, n53130, n53131, n53132,
         n53133, n53134, n53135, n53136, n53137, n53138, n53139, n53140,
         n53141, n53142, n53143, n53144, n53145, n53146, n53147, n53148,
         n53149, n53150, n53151, n53152, n53153, n53154, n53155, n53156,
         n53157, n53158, n53159, n53160, n53161, n53162, n53163, n53164,
         n53165, n53166, n53167, n53168, n53169, n53170, n53171, n53172,
         n53173, n53174, n53175, n53176, n53177, n53178, n53179, n53180,
         n53181, n53182, n53183, n53184, n53185, n53186, n53187, n53188,
         n53189, n53190, n53191, n53192, n53193, n53194, n53195, n53196,
         n53197, n53198, n53199, n53200, n53201, n53202, n53203, n53204,
         n53205, n53206, n53207, n53208, n53209, n53210, n53211, n53212,
         n53213, n53214, n53215, n53216, n53217, n53218, n53219, n53220,
         n53221, n53222, n53223, n53224, n53225, n53226, n53227, n53228,
         n53229, n53230, n53231, n53232, n53233, n53234, n53235, n53236,
         n53237, n53238, n53239, n53240, n53241, n53242, n53243, n53244,
         n53245, n53246, n53247, n53248, n53249, n53250, n53251, n53252,
         n53253, n53254, n53255, n53256, n53257, n53258, n53259, n53260,
         n53261, n53262, n53263, n53264, n53265, n53266, n53267, n53268,
         n53269, n53270, n53271, n53272, n53273, n53274, n53275, n53276,
         n53277, n53278, n53279, n53280, n53281, n53282, n53283, n53284,
         n53285, n53286, n53287, n53288, n53289, n53290, n53291, n53292,
         n53293, n53294, n53295, n53296, n53297, n53298, n53299, n53300,
         n53301, n53302, n53303, n53304, n53305, n53306, n53307, n53308,
         n53309, n53310, n53311, n53312, n53313, n53314, n53315, n53316,
         n53317, n53318, n53319, n53320, n53321, n53322, n53323, n53324,
         n53325, n53326, n53327, n53328, n53329, n53330, n53331, n53332,
         n53333, n53334, n53335, n53336, n53337, n53338, n53339, n53340,
         n53341, n53342, n53343, n53344, n53345, n53346, n53347, n53348,
         n53349, n53350, n53351, n53352, n53353, n53354, n53355, n53356,
         n53357, n53358, n53359, n53360, n53361, n53362, n53363, n53364,
         n53365, n53366, n53367, n53368, n53369, n53370, n53371, n53372,
         n53373, n53374, n53375, n53376, n53377, n53378, n53379, n53380,
         n53381, n53382, n53383, n53384, n53385, n53386, n53387, n53388,
         n53389, n53390, n53391, n53392, n53393, n53394, n53395, n53396,
         n53397, n53398, n53399, n53400, n53401, n53402, n53403, n53404,
         n53405, n53406, n53407, n53408, n53409, n53410, n53411, n53412,
         n53413, n53414, n53415, n53416, n53417, n53418, n53419, n53420,
         n53421, n53422, n53423, n53424, n53425, n53426, n53427, n53428,
         n53429, n53430, n53431, n53432, n53433, n53434, n53435, n53436,
         n53437, n53438, n53439, n53440, n53441, n53442, n53443, n53444,
         n53445, n53446, n53447, n53448, n53449, n53450, n53451, n53452,
         n53453, n53454, n53455, n53456, n53457, n53458, n53459, n53460,
         n53461, n53462, n53463, n53464, n53465, n53466, n53467, n53468,
         n53469, n53470, n53471, n53472, n53473, n53474, n53475, n53476,
         n53477, n53478, n53479, n53480, n53481, n53482, n53483, n53484,
         n53485, n53486, n53487, n53488, n53489, n53490, n53491, n53492,
         n53493, n53494, n53495, n53496, n53497, n53498, n53499, n53500,
         n53501, n53502, n53503, n53504, n53505, n53506, n53507, n53508,
         n53509, n53510, n53511, n53512, n53513, n53514, n53515, n53516,
         n53517, n53518, n53519, n53520, n53521, n53522, n53523, n53524,
         n53525, n53526, n53527, n53528, n53529, n53530, n53531, n53532,
         n53533, n53534, n53535, n53536, n53537, n53538, n53539, n53540,
         n53541, n53542, n53543, n53544, n53545, n53546, n53547, n53548,
         n53549, n53550, n53551, n53552, n53553, n53554, n53555, n53556,
         n53557, n53558, n53559, n53560, n53561, n53562, n53563, n53564,
         n53565, n53566, n53567, n53568, n53569, n53570, n53571, n53572,
         n53573, n53574, n53575, n53576, n53577, n53578, n53579, n53580,
         n53581, n53582, n53583, n53584, n53585, n53586, n53587, n53588,
         n53589, n53590, n53591, n53592, n53593, n53594, n53595, n53596,
         n53597, n53598, n53599, n53600, n53601, n53602, n53603, n53604,
         n53605, n53606, n53607, n53608, n53609, n53610, n53611, n53612,
         n53613, n53614, n53615, n53616, n53617, n53618, n53619, n53620,
         n53621, n53622, n53623, n53624, n53625, n53626, n53627, n53628,
         n53629, n53630, n53631, n53632, n53633, n53634, n53635, n53636,
         n53637, n53638, n53639, n53640, n53641, n53642, n53643, n53644,
         n53645, n53646, n53647, n53648, n53649, n53650, n53651, n53652,
         n53653, n53654, n53655, n53656, n53657, n53658, n53659, n53660,
         n53661, n53662, n53663, n53664, n53665, n53666, n53667, n53668,
         n53669, n53670, n53671, n53672, n53673, n53674, n53675, n53676,
         n53677, n53678, n53679, n53680, n53681, n53682, n53683, n53684,
         n53685, n53686, n53687, n53688, n53689, n53690, n53691, n53692,
         n53693, n53694, n53695, n53696, n53697, n53698, n53699, n53700,
         n53701, n53702, n53703, n53704, n53705, n53706, n53707, n53708,
         n53709, n53710, n53711, n53712, n53713, n53714, n53715, n53716,
         n53717, n53718, n53720, n53722, n53724, n53726, n53728, n53730,
         n53732, n53734, n53736, n53738, n53740, n53742, n53744, n53746,
         n53748, n53750, n53752, n53754, n53756, n53758, n53760, n53762,
         n53764, n53766, n53768, n53770, n53772, n53774, n53776, n53778,
         n53780, n53782, n53784, n53786, n53788, n53790, n53792, n53794,
         n53796, n53798, n53800, n53802, n53804, n53806, n53808, n53810,
         n53812, n53814, n53816, n53818, n53820, n53822, n53824, n53826,
         n53828, n53830, n53832, n53834, n53836, n53838, n53840, n53842,
         n53844, n53846, n53848, n53850, n53852, n53854, n53856, n53858,
         n53860, n53862, n53864, n53866, n53868, n53870, n53872, n53874,
         n53876, n53878, n53880, n53882, n53884, n53886, n53888, n53890,
         n53892, n53894, n53896, n53898, n53900, n53902, n53904, n53906,
         n53908, n53910, n53912, n53914, n53916, n53918, n53920, n53922,
         n53924, n53926, n53928, n53930, n53932, n53934, n53936, n53938,
         n53940, n53942, n53944, n53946, n53948, n53950, n53952, n53954,
         n53956, n53958, n53960, n53962, n53964, n53966, n53968, n53970,
         n53972, n53974, n53976, n53978, n53980, n53982, n53984, n53986,
         n53988, n53990, n53992, n53994, n53996, n53998, n54000, n54002,
         n54004, n54006, n54008, n54010, n54012, n54014, n54016, n54018,
         n54020, n54022, n54024, n54026, n54028, n54030, n54032, n54034,
         n54036, n54038, n54040, n54042, n54044, n54046, n54048, n54050,
         n54052, n54054, n54056, n54058, n54060, n54062, n54064, n54066,
         n54068, n54070, n54072, n54074, n54076, n54078, n54080, n54082,
         n54084, n54086, n54088, n54090, n54092, n54094, n54096, n54098,
         n54100, n54102, n54104, n54106, n54108, n54110, n54112, n54114,
         n54116, n54118, n54120, n54122, n54124, n54126, n54128, n54130,
         n54132, n54134, n54136, n54138, n54140, n54142, n54144, n54146,
         n54148, n54150, n54152, n54154, n54156, n54158, n54160, n54162,
         n54164, n54166, n54168, n54170, n54172, n54174, n54176, n54178,
         n54180, n54182, n54184, n54186, n54188, n54190, n54192, n54194,
         n54196, n54198, n54200, n54202, n54204, n54206, n54208, n54210,
         n54212, n54214, n54216, n54218, n54220, n54222, n54224, n54226,
         n54228, n54230, n54232, n54234, n54236, n54238, n54240, n54242,
         n54244, n54246, n54248, n54250, n54252, n54254, n54256, n54258,
         n54260, n54262, n54264, n54266, n54268, n54270, n54272, n54274,
         n54276, n54278, n54280, n54282, n54284, n54286, n54288, n54290,
         n54292, n54294, n54296, n54298, n54300, n54302, n54304, n54306,
         n54308, n54310, n54312, n54314, n54316, n54318, n54320, n54322,
         n54324, n54326, n54328, n54330, n54332, n54334, n54336, n54338,
         n54340, n54342, n54344, n54346, n54348, n54350, n54352, n54354,
         n54356, n54358, n54360, n54362, n54364, n54366, n54368, n54370,
         n54372, n54374, n54376, n54378, n54380, n54382, n54384, n54386,
         n54388, n54390, n54392, n54394, n54396, n54398, n54400, n54402,
         n54404, n54406, n54408, n54410, n54412, n54414, n54416, n54418,
         n54420, n54422, n54424, n54426, n54428, n54430, n54432, n54434,
         n54436, n54438, n54440, n54442, n54444, n54446, n54448, n54450,
         n54452, n54454, n54456, n54458, n54460, n54462, n54464, n54466,
         n54468, n54470, n54472, n54474, n54476, n54478, n54480, n54482,
         n54484, n54486, n54488, n54490, n54492, n54494, n54496, n54498,
         n54500, n54502, n54504, n54506, n54508, n54510, n54512, n54514,
         n54516, n54518, n54520, n54522, n54524, n54526, n54528, n54530,
         n54532, n54534, n54536, n54538, n54540, n54542, n54544, n54546,
         n54548, n54550, n54552, n54554, n54556, n54558, n54560, n54562,
         n54564, n54566, n54568, n54570, n54572, n54574, n54576, n54578,
         n54580, n54582, n54584, n54586, n54588, n54590, n54592, n54594,
         n54596, n54598, n54600, n54602, n54604, n54606, n54608, n54610,
         n54612, n54614, n54616, n54618, n54620, n54622, n54624, n54626,
         n54628, n54630, n54632, n54634, n54636, n54638, n54640, n54642,
         n54644, n54646, n54648, n54650, n54652, n54654, n54656, n54658,
         n54660, n54662, n54664, n54666, n54668, n54670, n54672, n54674,
         n54676, n54678, n54680, n54682, n54684, n54686, n54688, n54690,
         n54692, n54694, n54696, n54698, n54700, n54702, n54704, n54706,
         n54708, n54710, n54712, n54714, n54716, n54718, n54720, n54722,
         n54724, n54726, n54728, n54730, n54732, n54734, n54736, n54738,
         n54740, n54742, n54744, n54746, n54748, n54750, n54752, n54754,
         n54756, n54758, n54760, n54762, n54764, n54766, n54768, n54770,
         n54772, n54774, n54776, n54778, n54780, n54782, n54784, n54786,
         n54788, n54790, n54792, n54794, n54796, n54798, n54800, n54802,
         n54804, n54806, n54808, n54810, n54812, n54814, n54816, n54818,
         n54820, n54822, n54824, n54826, n54828, n54830, n54832, n54834,
         n54836, n54838, n54840, n54842, n54844, n54846, n54848, n54850,
         n54852, n54854, n54856, n54858, n54860, n54862, n54864, n54866,
         n54868, n54870, n54872, n54874, n54876, n54878, n54880, n54882,
         n54884, n54886, n54888, n54890, n54892, n54894, n54896, n54898,
         n54900, n54902, n54904, n54906, n54908, n54910, n54912, n54914,
         n54916, n54918, n54920, n54922, n54924, n54926, n54928, n54930,
         n54932, n54934, n54936, n54938, n54940, n54942, n54944, n54946,
         n54948, n54950, n54952, n54954, n54956, n54958, n54960, n54962,
         n54964, n54966, n54968, n54970, n54972, n54974, n54976, n54978,
         n54980, n54982, n54984, n54986, n54988, n54990, n54992, n54994,
         n54996, n54998, n54999, n55000, n55001, n55002, n55003, n55004,
         n55005, n55006, n55007, n55008, n55009, n55010, n55011, n55012,
         n55013, n55014, n55015, n55016, n55017, n55018, n55019, n55020,
         n55021, n55022, n55023, n55024, n55025, n55026, n55027, n55028,
         n55029, n55030, n55031, n55032, n55033, n55034, n55035, n55036,
         n55037, n55038, n55039, n55040, n55041, n55042, n55043, n55044,
         n55045, n55046, n55047, n55048, n55049, n55050, n55051, n55052,
         n55053, n55054, n55055, n55056, n55057, n55058, n55059, n55060,
         n55061, n55062, n55063, n55064, n55065, n55066, n55067, n55068,
         n55069, n55070, n55071, n55072, n55073, n55074, n55075, n55076,
         n55077, n55078, n55079, n55080, n55081, n55082, n55083, n55084,
         n55085, n55086, n55087, n55088, n55089, n55090, n55091, n55092,
         n55093, n55094, n55095, n55096, n55097, n55098, n55099, n55100,
         n55101, n55102, n55103, n55104, n55105, n55106, n55107, n55108,
         n55109, n55110, n55111, n55112, n55113, n55114, n55115, n55116,
         n55117, n55118, n55119, n55120, n55121, n55122, n55123, n55124,
         n55125, n55126, n55127, n55128, n55129, n55130, n55131, n55132,
         n55133, n55134, n55135, n55136, n55137, n55138, n55139, n55140,
         n55141, n55142, n55143, n55144, n55145, n55146, n55147, n55148,
         n55149, n55150, n55151, n55152, n55153, n55154, n55155, n55156,
         n55157, n55158, n55159, n55160, n55161, n55162, n55163, n55164,
         n55165, n55166, n55167, n55168, n55169, n55170, n55171, n55172,
         n55173, n55174, n55175, n55176, n55177, n55178, n55179, n55180,
         n55181, n55182, n55183, n55184, n55185, n55186, n55187, n55188,
         n55189, n55190, n55191, n55192, n55193, n55194, n55195, n55196,
         n55197, n55198, n55199, n55200, n55201, n55202, n55203, n55204,
         n55205, n55206, n55207, n55208, n55209, n55210, n55211, n55212,
         n55213, n55214, n55215, n55216, n55217, n55218, n55219, n55220,
         n55221, n55222, n55223, n55224, n55225, n55226, n55227, n55228,
         n55229, n55230, n55231, n55232, n55233, n55234, n55235, n55236,
         n55237, n55238, n55239, n55240, n55241, n55242, n55243, n55244,
         n55245, n55246, n55247, n55248, n55249, n55250, n55251, n55252,
         n55253, n55254, n55255, n55256, n55257, n55258, n55259, n55260,
         n55261, n55262, n55263, n55264, n55265, n55266, n55267, n55268,
         n55269, n55270, n55271, n55272, n55273, n55274, n55275, n55276,
         n55277, n55278, n55279, n55280, n55281, n55282, n55283, n55284,
         n55285, n55286, n55287, n55288, n55289, n55290, n55291, n55292,
         n55293, n55294, n55295, n55296, n55297, n55298, n55299, n55300,
         n55301, n55302, n55303, n55304, n55305, n55306, n55307, n55308,
         n55309, n55310, n55311, n55312, n55313, n55314, n55315, n55316,
         n55317, n55318, n55319, n55320, n55321, n55322, n55323, n55324,
         n55325, n55326, n55327, n55328, n55329, n55330, n55331, n55332,
         n55333, n55334, n55335, n55336, n55337, n55338, n55339, n55340,
         n55341, n55342, n55343, n55344, n55345, n55346, n55347, n55348,
         n55349, n55350, n55351, n55352, n55353, n55354, n55355, n55356,
         n55357, n55358, n55359, n55360, n55361, n55362, n55363, n55364,
         n55365, n55366, n55367, n55368, n55369, n55370, n55371, n55372,
         n55373, n55374, n55375, n55376, n55377, n55378, n55379, n55380,
         n55381, n55382, n55383, n55384, n55385, n55386, n55387, n55388,
         n55389, n55390, n55391, n55392, n55393, n55394, n55395, n55396,
         n55397, n55398, n55399, n55400, n55401, n55402, n55403, n55404,
         n55405, n55406, n55407, n55408, n55409, n55410, n55411, n55412,
         n55413, n55414, n55415, n55416, n55417, n55418, n55419, n55420,
         n55421, n55422, n55423, n55424, n55425, n55426, n55427, n55428,
         n55429, n55430, n55431, n55432, n55433, n55434, n55435, n55436,
         n55437, n55438, n55439, n55440, n55441, n55442, n55443, n55444,
         n55445, n55446, n55447, n55448, n55449, n55450, n55451, n55452,
         n55453, n55454, n55455, n55456, n55457, n55458, n55459, n55460,
         n55461, n55462, n55463, n55464, n55465, n55466, n55467, n55468,
         n55469, n55470, n55471, n55472, n55473, n55474, n55475, n55476,
         n55477, n55478, n55479, n55480, n55481, n55482, n55483, n55484,
         n55485, n55486, n55487, n55488, n55489, n55490, n55491, n55492,
         n55493, n55494, n55495, n55496, n55497, n55498, n55499, n55500,
         n55501, n55502, n55503, n55504, n55505, n55506, n55507, n55508,
         n55509, n55510, n55511, n55512, n55513, n55514, n55515, n55516,
         n55517, n55518, n55519, n55520, n55521, n55522, n55523, n55524,
         n55525, n55526, n55527, n55528, n55529, n55530, n55531, n55532,
         n55533, n55534, n55535, n55536, n55537, n55538, n55539, n55540,
         n55541, n55542, n55543, n55544, n55545, n55546, n55547, n55548,
         n55549, n55550, n55551, n55552, n55553, n55554, n55555, n55556,
         n55557, n55558, n55559, n55560, n55561, n55562, n55563, n55564,
         n55565, n55566, n55567, n55568, n55569, n55570, n55571, n55572,
         n55573, n55574, n55575, n55576, n55577, n55578, n55579, n55580,
         n55581, n55582, n55583, n55584, n55585, n55586, n55587, n55588,
         n55589, n55590, n55591, n55592, n55593, n55594, n55595, n55596,
         n55597, n55598, n55599, n55600, n55601, n55602, n55603, n55604,
         n55605, n55606, n55607, n55608, n55609, n55610, n55611, n55612,
         n55613, n55614, n55615, n55616, n55617, n55618, n55619, n55620,
         n55621, n55622, n55623, n55624, n55625, n55626, n55627, n55628,
         n55629, n55630, n55631, n55632, n55633, n55634, n55635, n55636,
         n55637, n55638, n55639, n55640, n55641, n55642, n55643, n55644,
         n55645, n55646, n55647, n55648, n55649, n55650, n55651, n55652,
         n55653, n55654, n55655, n55656, n55657, n55658, n55659, n55660,
         n55661, n55662, n55663, n55664, n55665, n55666, n55667, n55668,
         n55669, n55670, n55671, n55672, n55673, n55674, n55675, n55676,
         n55677, n55678, n55679, n55680, n55681, n55682, n55683, n55684,
         n55685, n55686, n55687, n55688, n55689, n55690, n55691, n55692,
         n55693, n55694, n55695, n55696, n55697, n55698, n55699, n55700,
         n55701, n55702, n55703, n55704, n55705, n55706, n55707, n55708,
         n55709, n55710, n55711, n55712, n55713, n55714, n55715, n55716,
         n55717, n55718, n55719, n55720, n55721, n55722, n55723, n55724,
         n55725, n55726, n55727, n55728, n55729, n55730, n55731, n55732,
         n55733, n55734, n55735, n55736, n55737, n55738, n55739, n55740,
         n55741, n55742, n55743, n55744, n55745, n55746, n55747, n55748,
         n55749, n55750, n55751, n55752, n55753, n55754, n55755, n55756,
         n55757, n55758, n55759, n55760, n55761, n55762, n55763, n55764,
         n55765, n55766, n55767, n55768, n55769, n55770, n55771, n55772,
         n55773, n55774, n55775, n55776, n55777, n55778, n55779, n55780,
         n55781, n55782, n55783, n55784, n55785, n55786, n55787, n55788,
         n55789, n55790, n55791, n55792, n55793, n55794, n55795, n55796,
         n55797, n55798, n55799, n55800, n55801, n55802, n55803, n55804,
         n55805, n55806, n55807, n55808, n55809, n55810, n55811, n55812,
         n55813, n55814, n55815, n55816, n55817, n55818, n55819, n55820,
         n55821, n55822, n55823, n55824, n55825, n55826, n55827, n55828,
         n55829, n55830, n55831, n55832, n55833, n55834, n55835, n55836,
         n55837, n55838, n55839, n55840, n55841, n55842, n55843, n55844,
         n55845, n55846, n55847, n55848, n55849, n55850, n55851, n55852,
         n55853, n55854, n55855, n55856, n55857, n55858, n55859, n55860,
         n55861, n55862, n55863, n55864, n55865, n55866, n55867, n55868,
         n55869, n55870, n55871, n55872, n55873, n55874, n55875, n55876,
         n55877, n55878, n55879, n55880, n55881, n55882, n55883, n55884,
         n55885, n55886, n55887, n55888, n55889, n55890, n55891, n55892,
         n55893, n55894, n55895, n55896, n55897, n55898, n55899, n55900,
         n55901, n55902, n55903, n55904, n55905, n55906, n55907, n55908,
         n55909, n55910, n55911, n55912, n55913, n55914, n55915, n55916,
         n55917, n55918, n55919, n55920, n55921, n55922, n55923, n55924,
         n55925, n55926, n55927, n55928, n55929, n55930, n55931, n55932,
         n55933, n55934, n55935, n55936, n55937, n55938, n55939, n55940,
         n55941, n55942, n55943, n55944, n55945, n55946, n55947, n55948,
         n55949, n55950, n55951, n55952, n55953, n55954, n55955, n55956,
         n55957, n55958, n55959, n55960, n55961, n55962, n55963, n55964,
         n55965, n55966, n55967, n55968, n55969, n55970, n55971, n55972,
         n55973, n55974, n55975, n55976, n55977, n55978, n55979, n55980,
         n55981, n55982, n55983, n55984, n55985, n55986, n55987, n55988,
         n55989, n55990, n55991, n55992, n55993, n55994, n55995, n55996,
         n55997, n55998, n55999, n56000, n56001, n56002, n56003, n56004,
         n56005, n56006, n56007, n56008, n56009, n56010, n56011, n56012,
         n56013, n56014, n56015, n56016, n56017, n56018, n56019, n56020,
         n56021, n56022, n56023, n56024, n56025, n56026, n56027, n56028,
         n56029, n56030, n56031, n56032, n56033, n56034, n56035, n56036,
         n56037, n56038, n56039, n56040, n56041, n56042, n56043, n56044,
         n56045, n56046, n56047, n56048, n56049, n56050, n56051, n56052,
         n56053, n56054, n56055, n56056, n56057, n56058, n56059, n56060,
         n56061, n56062, n56063, n56064, n56065, n56066, n56067, n56068,
         n56069, n56070, n56071, n56072, n56073, n56074, n56075, n56076,
         n56077, n56078, n56079, n56080, n56081, n56082, n56083, n56084,
         n56085, n56086, n56087, n56088, n56089, n56090, n56091, n56092,
         n56093, n56094, n56095, n56096, n56097, n56098, n56099, n56100,
         n56101, n56102, n56103, n56104, n56105, n56106, n56107, n56108,
         n56109, n56110, n56111, n56112, n56113, n56114, n56115, n56116,
         n56117, n56118, n56119, n56120, n56121, n56122, n56123, n56124,
         n56125, n56126, n56127, n56128, n56129, n56130, n56131, n56132,
         n56133, n56134, n56135, n56136, n56137, n56138, n56139, n56140,
         n56141, n56142, n56143, n56144, n56145, n56146, n56147, n56148,
         n56149, n56150, n56151, n56152, n56153, n56154, n56155, n56156,
         n56157, n56158, n56159, n56160, n56161, n56162, n56163, n56164,
         n56165, n56166, n56167, n56168, n56169, n56170, n56171, n56172,
         n56173, n56174, n56175, n56176, n56177, n56178, n56179, n56180,
         n56181, n56182, n56183, n56184, n56185, n56186, n56187, n56188,
         n56189, n56190, n56191, n56192, n56193, n56194, n56195, n56196,
         n56197, n56198, n56199, n56200, n56201, n56202, n56203, n56204,
         n56205, n56206, n56207, n56208, n56209, n56210, n56211, n56212,
         n56213, n56214, n56215, n56216, n56217, n56218, n56219, n56220,
         n56221, n56222, n56223, n56224, n56225, n56226, n56227, n56228,
         n56229, n56230, n56231, n56232, n56233, n56234, n56235, n56236,
         n56237, n56238, n56239, n56240, n56241, n56242, n56243, n56244,
         n56245, n56246, n56247, n56248, n56249, n56250, n56251, n56252,
         n56253, n56254, n56255, n56256, n56257, n56258, n56259, n56260,
         n56261, n56262, n56263, n56264, n56265, n56266, n56267, n56268,
         n56269, n56270, n56271, n56272, n56273, n56274, n56275, n56276,
         n56277, n56278, n56279, n56280, n56281, n56282, n56283, n56284,
         n56285, n56286, n56287, n56288, n56289, n56290, n56291, n56292,
         n56293, n56294, n56295, n56296, n56297, n56298, n56299, n56300,
         n56301, n56302, n56303, n56304, n56305, n56306, n56307, n56308,
         n56309, n56310, n56311, n56312, n56313, n56314, n56315, n56316,
         n56317, n56318, n56319, n56320, n56321, n56322, n56323, n56324,
         n56325, n56326, n56327, n56328, n56329, n56330, n56331, n56332,
         n56333, n56334, n56335, n56336, n56337, n56338, n56339, n56340,
         n56341, n56342, n56343, n56344, n56345, n56346, n56347, n56348,
         n56349, n56350, n56351, n56352, n56353, n56354, n56355, n56356,
         n56357, n56358, n56359, n56360, n56361, n56362, n56363, n56364,
         n56365, n56366, n56367, n56368, n56369, n56370, n56371, n56372,
         n56373, n56374, n56375, n56376, n56377, n56378, n56379, n56380,
         n56381, n56382, n56383, n56384, n56385, n56386, n56387, n56388,
         n56389, n56390, n56391, n56392, n56393, n56394, n56395, n56396,
         n56397, n56398, n56399, n56400, n56401, n56402, n56403, n56404,
         n56405, n56406, n56407, n56408, n56409, n56410, n56411, n56412,
         n56413, n56414, n56415, n56416, n56417, n56418, n56419, n56420,
         n56421, n56422, n56423, n56424, n56425, n56426, n56427, n56428,
         n56429, n56430, n56431, n56432, n56433, n56434, n56435, n56436,
         n56437, n56438, n56439, n56440, n56441, n56442, n56443, n56444,
         n56445, n56446, n56447, n56448, n56449, n56450, n56451, n56452,
         n56453, n56454, n56455, n56456, n56457, n56458, n56459, n56460,
         n56461, n56462, n56463, n56464, n56465, n56466, n56467, n56468,
         n56469, n56470, n56471, n56472, n56473, n56474, n56475, n56476,
         n56477, n56478, n56479, n56480, n56481, n56482, n56483, n56484,
         n56485, n56486, n56487, n56488, n56489, n56490, n56491, n56492,
         n56493, n56494, n56495, n56496, n56497, n56498, n56499, n56500,
         n56501, n56502, n56503, n56504, n56505, n56506, n56507, n56508,
         n56509, n56510, n56511, n56512, n56513, n56514, n56515, n56516,
         n56517, n56518, n56519, n56520, n56521, n56522, n56523, n56524,
         n56525, n56526, n56527, n56528, n56529, n56530, n56531, n56532,
         n56533, n56534, n56535, n56536, n56537, n56538, n56539, n56540,
         n56541, n56542, n56543, n56544, n56545, n56546, n56547, n56548,
         n56549, n56550, n56551, n56552, n56553, n56554, n56555, n56556,
         n56557, n56558, n56559, n56560, n56561, n56562, n56563, n56564,
         n56565, n56566, n56567, n56568, n56569, n56570, n56571, n56572,
         n56573, n56574, n56575, n56576, n56577, n56578, n56579, n56580,
         n56581, n56582, n56583, n56584, n56585, n56586, n56587, n56588,
         n56589, n56590, n56591, n56592, n56593, n56594, n56595, n56596,
         n56598, n56600, n56602, n56604, n56606, n56608, n56610, n56612,
         n56614, n56616, n56618, n56620, n56622, n56624, n56626, n56628,
         n56630, n56632, n56634, n56636, n56638, n56640, n56642, n56644,
         n56646, n56648, n56650, n56652, n56654, n56656, n56658, n56660,
         n56661, n56662, n56663, n56664, n56665, n56666, n56667, n56668,
         n56669, n56670, n56671, n56672, n56673, n56674, n56675, n56676,
         n56677, n56678, n56679, n56680, n56681, n56682, n56683, n56684,
         n56685, n56686, n56687, n56688, n56689, n56690, n56691, n56692,
         n56693, n56694, n56695, n56696, n56697, n56698, n56699, n56700,
         n56701, n56702, n56703, n56704, n56705, n56706, n56707, n56708,
         n56709, n56710, n56711, n56712, n56713, n56714, n56715, n56716,
         n56717, n56718, n56719, n56720, n56721, n56722, n56723, n56724,
         n56725, n56726, n56727, n56728, n56729, n56730, n56731, n56732,
         n56733, n56734, n56735, n56736, n56737, n56738, n56739, n56740,
         n56741, n56742, n56743, n56744, n56745, n56746, n56747, n56748,
         n56749, n56750, n56751, n56752, n56753, n56754, n56755, n56756,
         n56757, n56758, n56759, n56760, n56761, n56762, n56763, n56764,
         n56765, n56766, n56767, n56768, n56769, n56770, n56771, n56772,
         n56773, n56774, n56775, n56776, n56777, n56778, n56779, n56780,
         n56781, n56782, n56783, n56784, n56785, n56786, n56787, n56788,
         n56789, n56790, n56791, n56792, n56793, n56794, n56795, n56796,
         n56797, n56798, n56799, n56800, n56801, n56802, n56803, n56804,
         n56805, n56806, n56807, n56808, n56809, n56810, n56811, n56812,
         n56813, n56814, n56815, n56816, n56817, n56818, n56819, n56820,
         n56821, n56822, n56823, n56824, n56825, n56826, n56827, n56828,
         n56829, n56830, n56831, n56832, n56833, n56834, n56835, n56836,
         n56837, n56838, n56839, n56840, n56841, n56842, n56843, n56844,
         n56845, n56846, n56847, n56848, n56849, n56850, n56851, n56852,
         n56853, n56854, n56855, n56856, n56857, n56858, n56859, n56860,
         n56861, n56862, n56863, n56864, n56865, n56866, n56867, n56868,
         n56869, n56870, n56871, n56872, n56873, n56874, n56875, n56876,
         n56877, n56878, n56879, n56880, n56881, n56882, n56883, n56884,
         n56885, n56886, n56887, n56888, n56889, n56890, n56891, n56892,
         n56893, n56894, n56895, n56896, n56897, n56898, n56899, n56900,
         n56901, n56902, n56903, n56904, n56905, n56906, n56907, n56908,
         n56909, n56910, n56911, n56912, n56913, n56914, n56915, n56916,
         n56917, n56918, n56919, n56920, n56921, n56922, n56923, n56924,
         n56925, n56926, n56927, n56928, n56929, n56930, n56931, n56932,
         n56933, n56934, n56935, n56936, n56937, n56938, n56939, n56940,
         n56941, n56942, n56943, n56944, n56945, n56946, n56947, n56948,
         n56949, n56950, n56951, n56952, n56953, n56954, n56955, n56956,
         n56957, n56958, n56959, n56960, n56961, n56962, n56963, n56964,
         n56965, n56966, n56967, n56968, n56969, n56970, n56971, n56972,
         n56973, n56974, n56975, n56976, n56977, n56978, n56979, n56980,
         n56981, n56982, n56983, n56984, n56985, n56986, n56987, n56988,
         n56989, n56990, n56991, n56992, n56993, n56994, n56995, n56996,
         n56997, n56998, n56999, n57000, n57001, n57002, n57003, n57004,
         n57005, n57006, n57007, n57008, n57009, n57010, n57011, n57012,
         n57013, n57014, n57015, n57016, n57017, n57018, n57019, n57020,
         n57021, n57022, n57023, n57024, n57025, n57026, n57027, n57028,
         n57029, n57030, n57031, n57032, n57033, n57034, n57035, n57036,
         n57037, n57038, n57039, n57040, n57041, n57042, n57043, n57044,
         n57045, n57046, n57047, n57048, n57049, n57050, n57051, n57052,
         n57053, n57054, n57055, n57056, n57057, n57058, n57059, n57060,
         n57061, n57062, n57063, n57064, n57065, n57066, n57067, n57068,
         n57069, n57070, n57071, n57072, n57073, n57074, n57075, n57076,
         n57077, n57078, n57079, n57080, n57081, n57082, n57083, n57084,
         n57085, n57086, n57087, n57088, n57089, n57090, n57091, n57092,
         n57093, n57094, n57095, n57096, n57097, n57098, n57099, n57100,
         n57101, n57102, n57103, n57104, n57105, n57106, n57107, n57108,
         n57109, n57110, n57111, n57112, n57113, n57114, n57115, n57116,
         n57117, n57118, n57119, n57120, n57121, n57122, n57123, n57124,
         n57125, n57126, n57127, n57128, n57129, n57130, n57131, n57132,
         n57133, n57134, n57135, n57136, n57137, n57138, n57139, n57140,
         n57141, n57142, n57143, n57144, n57145, n57146, n57147, n57148,
         n57149, n57150, n57151, n57152, n57153, n57154, n57155, n57156,
         n57157, n57158, n57159, n57160, n57161, n57162, n57163, n57164,
         n57165, n57166, n57167, n57168, n57169, n57170, n57171, n57172,
         n57173, n57174, n57175, n57176, n57177, n57178, n57179, n57180,
         n57181, n57182, n57183, n57184, n57185, n57186, n57187, n57188,
         n57189, n57190, n57191, n57192, n57193, n57194, n57195, n57196,
         n57197, n57198, n57199, n57200, n57201, n57202, n57203, n57204,
         n57205, n57206, n57207, n57208, n57209, n57210, n57211, n57212,
         n57213, n57214, n57215, n57216, n57217, n57218, n57219, n57220,
         n57221, n57222, n57223, n57224, n57225, n57226, n57227, n57228,
         n57229, n57230, n57231, n57232, n57233, n57234, n57235, n57236,
         n57237, n57238, n57239, n57240, n57241, n57242, n57243, n57244,
         n57245, n57246, n57247, n57248, n57249, n57250, n57251, n57252,
         n57253, n57254, n57255, n57256, n57257, n57258, n57259, n57260,
         n57261, n57262, n57263, n57264, n57265, n57266, n57267, n57268,
         n57269, n57270, n57271, n57272, n57273, n57274, n57275, n57276,
         n57277, n57278, n57279, n57280, n57281, n57282, n57283, n57284,
         n57285, n57286, n57287, n57288, n57289, n57290, n57291, n57292,
         n57293, n57294, n57295, n57296, n57297, n57298, n57299, n57300,
         n57301, n57302, n57303, n57304, n57305, n57306, n57307, n57308,
         n57309, n57310, n57311, n57312, n57313, n57314, n57315, n57316,
         n57317, n57318, n57319, n57320, n57321, n57322, n57323, n57324,
         n57325, n57326, n57327, n57328, n57329, n57330, n57331, n57332,
         n57333, n57334, n57335, n57336, n57337, n57338, n57339, n57340,
         n57341, n57342, n57343, n57344, n57345, n57346, n57347, n57348,
         n57349, n57350, n57351, n57352, n57353, n57354, n57355, n57356,
         n57357, n57358, n57359, n57360, n57361, n57362, n57363, n57364,
         n57365, n57366, n57367, n57368, n57369, n57370, n57371, n57372,
         n57373, n57374, n57375, n57376, n57377, n57378, n57379, n57380,
         n57381, n57382, n57383, n57384, n57385, n57386, n57387, n57388,
         n57389, n57390, n57391, n57392, n57393, n57394, n57395, n57396,
         n57397, n57398, n57399, n57400, n57401, n57402, n57403, n57404,
         n57405, n57406, n57407, n57408, n57409, n57410, n57411, n57412,
         n57413, n57414, n57415, n57416, n57417, n57418, n57419, n57420,
         n57421, n57422, n57423, n57424, n57425, n57426, n57427, n57428,
         n57429, n57430, n57431, n57432, n57433, n57434, n57435, n57436,
         n57437, n57438, n57439, n57440, n57441, n57442, n57443, n57444,
         n57445, n57446, n57447, n57448, n57449, n57450, n57451, n57452,
         n57453, n57454, n57455, n57456, n57457, n57458, n57459, n57460,
         n57461, n57462, n57463, n57464, n57465, n57466, n57467, n57468,
         n57469, n57470, n57471, n57472, n57473, n57474, n57475, n57476,
         n57477, n57478, n57479, n57480, n57481, n57482, n57483, n57484,
         n57485, n57486, n57487, n57488, n57489, n57490, n57491, n57492,
         n57493, n57494, n57495, n57496, n57497, n57498, n57499, n57500,
         n57501, n57502, n57503, n57504, n57505, n57506, n57507, n57508,
         n57509, n57510, n57511, n57512, n57513, n57514, n57515, n57516,
         n57517, n57518, n57519, n57520, n57521, n57522, n57523, n57524,
         n57525, n57526, n57527, n57528, n57529, n57530, n57531, n57532,
         n57533, n57534, n57535, n57536, n57537, n57538, n57539, n57540,
         n57541, n57542, n57543, n57544, n57545, n57546, n57547, n57548,
         n57549, n57550, n57551, n57552, n57553, n57554, n57555, n57556,
         n57557, n57558, n57559, n57560, n57561, n57562, n57563, n57564,
         n57565, n57566, n57567, n57568, n57569, n57570, n57571, n57572,
         n57573, n57574, n57575, n57576, n57577, n57578, n57579, n57580,
         n57581, n57582, n57583, n57584, n57585, n57586, n57587, n57588,
         n57589, n57590, n57591, n57592, n57593, n57594, n57595, n57596,
         n57597, n57598, n57599, n57600, n57601, n57602, n57603, n57604,
         n57605, n57606, n57607, n57608, n57609, n57610, n57611, n57612,
         n57613, n57614, n57615, n57616, n57617, n57618, n57619, n57620,
         n57621, n57622, n57623, n57624, n57625, n57626, n57627, n57628,
         n57629, n57630, n57631, n57632, n57633, n57634, n57635, n57636,
         n57637, n57638, n57639, n57640, n57641, n57642, n57643, n57644,
         n57645, n57646, n57647, n57648, n57649, n57650, n57651, n57652,
         n57653, n57654, n57655, n57656, n57657, n57658, n57659, n57660,
         n57661, n57662, n57663, n57664, n57665, n57666, n57667, n57668,
         n57669, n57670, n57671, n57672, n57673, n57674, n57675, n57676,
         n57677, n57678, n57679, n57680, n57681, n57682, n57683, n57684,
         n57685, n57686, n57687, n57688, n57689, n57690, n57691, n57692,
         n57693, n57694, n57695, n57696, n57697, n57698, n57699, n57700,
         n57701, n57702, n57703, n57704, n57705, n57706, n57707, n57708,
         n57709, n57710, n57711, n57712, n57713, n57714, n57715, n57716,
         n57717, n57718, n57719, n57720, n57721, n57722, n57723, n57724,
         n57725, n57726, n57727, n57728, n57729, n57730, n57731, n57732,
         n57733, n57734, n57735, n57736, n57737, n57738, n57739, n57740,
         n57741, n57742, n57743, n57744, n57745, n57746, n57747, n57748,
         n57749, n57750, n57751, n57752, n57753, n57754, n57755, n57756,
         n57757, n57758, n57759, n57760, n57761, n57762, n57763, n57764,
         n57765, n57766, n57767, n57768, n57769, n57770, n57771, n57772,
         n57773, n57774, n57775, n57776, n57777, n57778, n57779, n57780,
         n57781, n57782, n57783, n57784, n57785, n57786, n57787, n57788,
         n57789, n57790, n57791, n57792, n57793, n57794, n57795, n57796,
         n57797, n57798, n57799, n57800, n57801, n57802, n57803, n57804,
         n57805, n57806, n57807, n57808, n57809, n57810, n57811, n57812,
         n57813, n57814, n57815, n57816, n57817, n57818, n57819, n57820,
         n57821, n57822, n57823, n57824, n57825, n57826, n57827, n57828,
         n57829, n57830, n57831, n57832, n57833, n57834, n57835, n57836,
         n57837, n57838, n57839, n57840, n57841, n57842, n57843, n57844,
         n57845, n57846, n57847, n57848, n57849, n57850, n57851, n57852,
         n57853, n57854, n57855, n57856, n57857, n57858, n57859, n57860,
         n57861, n57862, n57863, n57864, n57865, n57866, n57867, n57868,
         n57869, n57870, n57871, n57872, n57873, n57874, n57875, n57876,
         n57877, n57878, n57879, n57880, n57881, n57882, n57883, n57884,
         n57885, n57886, n57887, n57888, n57889, n57890, n57891, n57892,
         n57893, n57894, n57895, n57896, n57897, n57898, n57899, n57900,
         n57901, n57902, n57903, n57904, n57905, n57906, n57907, n57908,
         n57909, n57910, n57911, n57912, n57913, n57914, n57915, n57916,
         n57917, n57918, n57919, n57920, n57921, n57922, n57923, n57924,
         n57925, n57926, n57927, n57928, n57929, n57930, n57931, n57932,
         n57933, n57934, n57935, n57936, n57937, n57938, n57939, n57940,
         n57941, n57942, n57943, n57944, n57945, n57946, n57947, n57948,
         n57949, n57950, n57951, n57952, n57953, n57954, n57955, n57956,
         n57957, n57958, n57959, n57960, n57961, n57962, n57963, n57964,
         n57965, n57966, n57967, n57968, n57969, n57970, n57971, n57972,
         n57973, n57974, n57975, n57976, n57977, n57978, n57979, n57980,
         n57981, n57982, n57983, n57984, n57985, n57986, n57987, n57988,
         n57989, n57990, n57991, n57992, n57993, n57994, n57995, n57996,
         n57997, n57998, n57999, n58000, n58001, n58002, n58003, n58004,
         n58005, n58006, n58007, n58008, n58009, n58010, n58011, n58012,
         n58013, n58014, n58015, n58016, n58017, n58018, n58019, n58020,
         n58021, n58022, n58023, n58024, n58025, n58026, n58027, n58028,
         n58029, n58030, n58031, n58032, n58033, n58034, n58035, n58036,
         n58037, n58038, n58039, n58040, n58041, n58042, n58043, n58044,
         n58045, n58046, n58047, n58048, n58049, n58050, n58051, n58052,
         n58053, n58054, n58055, n58056, n58057, n58058, n58059, n58060,
         n58061, n58062, n58063, n58064, n58065, n58066, n58067, n58068,
         n58069, n58070, n58071, n58072, n58073, n58074, n58075, n58076,
         n58077, n58078, n58079, n58080, n58081, n58082, n58083, n58084,
         n58085, n58086, n58087, n58088, n58089, n58090, n58091, n58092,
         n58093, n58094, n58095, n58096, n58097, n58098, n58099, n58100,
         n58101, n58102, n58103, n58104, n58105, n58106, n58107, n58108,
         n58109, n58110, n58111, n58112, n58113, n58114, n58115, n58116,
         n58117, n58118, n58119, n58120, n58121, n58122, n58123, n58124,
         n58125, n58126, n58127, n58128, n58129, n58130, n58131, n58132,
         n58133, n58134, n58135, n58136, n58137, n58138, n58139, n58140,
         n58141, n58142, n58143, n58144, n58145, n58146, n58147, n58148,
         n58149, n58150, n58151, n58152, n58153, n58154, n58155, n58156,
         n58157, n58158, n58159, n58160, n58161, n58162, n58163, n58164,
         n58165, n58166, n58167, n58168, n58169, n58170, n58171, n58172,
         n58173, n58174, n58175, n58176, n58177, n58178, n58179, n58180,
         n58181, n58182, n58183, n58184, n58185, n58186, n58187, n58188,
         n58189, n58190, n58191, n58192, n58193, n58194, n58195, n58196,
         n58197, n58198, n58199, n58200, n58201, n58202, n58203, n58204,
         n58205, n58206, n58207, n58208, n58209, n58210, n58211, n58212,
         n58213, n58214, n58215, n58216, n58217, n58218, n58219, n58220,
         n58221, n58222, n58223, n58224, n58225, n58226, n58227, n58228,
         n58229, n58230, n58231, n58232, n58233, n58234, n58235, n58236,
         n58237, n58238, n58239, n58240, n58241, n58242, n58243, n58244,
         n58245, n58246, n58247, n58248, n58249, n58250, n58251, n58252,
         n58253, n58254, n58255, n58256, n58257, n58258, n58259, n58260,
         n58261, n58262, n58263, n58264, n58265, n58266, n58267, n58268,
         n58269, n58270, n58271, n58272, n58273, n58274, n58275, n58276,
         n58277, n58278, n58279, n58280, n58281, n58282, n58283, n58284,
         n58285, n58286, n58287, n58288, n58289, n58290, n58291, n58292,
         n58293, n58294, n58295, n58296, n58297, n58298, n58299, n58300,
         n58301, n58302, n58303, n58304, n58305, n58306, n58307, n58308,
         n58309, n58310, n58311, n58312, n58313, n58314, n58315, n58316,
         n58317, n58318, n58319, n58320, n58321, n58322, n58323, n58324,
         n58325, n58326, n58327, n58328, n58329, n58330, n58331, n58332,
         n58333, n58334, n58335, n58336, n58337, n58338, n58339, n58340,
         n58341, n58342, n58343, n58344, n58345, n58346, n58347, n58348,
         n58349, n58350, n58351, n58352, n58353, n58354, n58355, n58356,
         n58357, n58358, n58359, n58360, n58361, n58362, n58363, n58364,
         n58365, n58366, n58367, n58368, n58369, n58370, n58371, n58372,
         n58373, n58374, n58375, n58376, n58377, n58378, n58379, n58380,
         n58381, n58382, n58383, n58384, n58385, n58386, n58387, n58388,
         n58389, n58390, n58391, n58392, n58393, n58394, n58395, n58396,
         n58397, n58398, n58399, n58400, n58401, n58402, n58403, n58404,
         n58405, n58406, n58407, n58408, n58409, n58410, n58411, n58412,
         n58413, n58414, n58415, n58416, n58417, n58418, n58419, n58420,
         n58421, n58422, n58423, n58424, n58425, n58426, n58427, n58428,
         n58429, n58430, n58431, n58432, n58433, n58434, n58435, n58436,
         n58437, n58438, n58439, n58440, n58441, n58442, n58443, n58444,
         n58445, n58446, n58447, n58448, n58449, n58450, n58451, n58452,
         n58453, n58454, n58455, n58456, n58457, n58458, n58459, n58460,
         n58461, n58462, n58463, n58464, n58465, n58466, n58467, n58468,
         n58469, n58470, n58471, n58472, n58473, n58474, n58475, n58476,
         n58477, n58478, n58479, n58480, n58481, n58482, n58483, n58484,
         n58485, n58486, n58487, n58488, n58489, n58490, n58491, n58492,
         n58493, n58494, n58495, n58496, n58497, n58498, n58499, n58500,
         n58501, n58502, n58503, n58504, n58505, n58506, n58507, n58508,
         n58509, n58510, n58511, n58512, n58513, n58514, n58515, n58516,
         n58517, n58518, n58519, n58520, n58521, n58522, n58523, n58524,
         n58525, n58526, n58527, n58528, n58529, n58530, n58531, n58532,
         n58533, n58534, n58535, n58536, n58537, n58538, n58539, n58540,
         n58541, n58542, n58543, n58544, n58545, n58546, n58547, n58548,
         n58549, n58550, n58551, n58552, n58553, n58554, n58555, n58556,
         n58557, n58558, n58559, n58560, n58561, n58562, n58563, n58564,
         n58565, n58566, n58567, n58568, n58569, n58570, n58571, n58572,
         n58573, n58574, n58575, n58576, n58577, n58578, n58579, n58580,
         n58581, n58582, n58583, n58584, n58585, n58586, n58587, n58588,
         n58589, n58590, n58591, n58592, n58593, n58594, n58595, n58596,
         n58597, n58598, n58599, n58600, n58601, n58602, n58603, n58604,
         n58605, n58606, n58607, n58608, n58609, n58610, n58611, n58612,
         n58613, n58614, n58615, n58616, n58617, n58618, n58619, n58620,
         n58621, n58622, n58623, n58624, n58625, n58626, n58627, n58628,
         n58629, n58630, n58631, n58632, n58633, n58634, n58635, n58636,
         n58637, n58638, n58639, n58640, n58641, n58642, n58643, n58644,
         n58645, n58646, n58647, n58648, n58649, n58650, n58651, n58652,
         n58653, n58654, n58655, n58656, n58657, n58658, n58659, n58660,
         n58661, n58662, n58663, n58664, n58665, n58666, n58667, n58668,
         n58669, n58670, n58671, n58672, n58673, n58674, n58675, n58676,
         n58677, n58678, n58679, n58680, n58681, n58682, n58683, n58684,
         n58685, n58686, n58687, n58688, n58689, n58690, n58691, n58692,
         n58693, n58694, n58695, n58696, n58697, n58698, n58699, n58700,
         n58701, n58702, n58703, n58704, n58705, n58706, n58707, n58708,
         n58709, n58710, n58711, n58712, n58713, n58714, n58715, n58716,
         n58717, n58718, n58719, n58720, n58721, n58722, n58723, n58724,
         n58725, n58726, n58727, n58728, n58729, n58730, n58731, n58732,
         n58733, n58734, n58735, n58736, n58737, n58738, n58739, n58740,
         n58741, n58742, n58743, n58744, n58745, n58746, n58747, n58748,
         n58749, n58750, n58751, n58752, n58753, n58754, n58755, n58756,
         n58757, n58758, n58759, n58760, n58761, n58762, n58763, n58764,
         n58765, n58766, n58767, n58768, n58769, n58770, n58771, n58772,
         n58773, n58774, n58775, n58776, n58777, n58778, n58779, n58780,
         n58781, n58782, n58783, n58784, n58785, n58786, n58787, n58788,
         n58789, n58790, n58791, n58792, n58793, n58794, n58795, n58796,
         n58797, n58798, n58799, n58800, n58801, n58802, n58803, n58804,
         n58805, n58806, n58807, n58808, n58809, n58810, n58811, n58812,
         n58813, n58814, n58815, n58816, n58817, n58818, n58819, n58820,
         n58821, n58822, n58823, n58824, n58825, n58826, n58827, n58828,
         n58829, n58830, n58831, n58832, n58833, n58834, n58835, n58836,
         n58837, n58838, n58839, n58840, n58841, n58842, n58843, n58844,
         n58845, n58846, n58847, n58848, n58849, n58850, n58851, n58852,
         n58853, n58854, n58855, n58856, n58857, n58858, n58859, n58860,
         n58861, n58862, n58863, n58864, n58865, n58866, n58867, n58868,
         n58869, n58870, n58871, n58872, n58873, n58874, n58875, n58876,
         n58877, n58878, n58879, n58880, n58881, n58882, n58883, n58884,
         n58885, n58886, n58887, n58888, n58889, n58890, n58891, n58892,
         n58893, n58894, n58895, n58896, n58897, n58898, n58899, n58900,
         n58901, n58902, n58903, n58904, n58905, n58906, n58907, n58908,
         n58909, n58910, n58911, n58912, n58913, n58914, n58915, n58916,
         n58917, n58918, n58919, n58920, n58921, n58922, n58923, n58924,
         n58925, n58926, n58927, n58928, n58929, n58930, n58931, n58932,
         n58933, n58934, n58935, n58936, n58937, n58938, n58939, n58940,
         n58941, n58942, n58943, n58944, n58945, n58946, n58947, n58948,
         n58949, n58950, n58951, n58952, n58953, n58954, n58955, n58956,
         n58957, n58958, n58959, n58960, n58961, n58962, n58963, n58964,
         n58965, n58966, n58967, n58968, n58969, n58970, n58971, n58972,
         n58973, n58974, n58975, n58976, n58977, n58978, n58979, n58980,
         n58981, n58982, n58983, n58984, n58985, n58986, n58987, n58988,
         n58989, n58990, n58991, n58992, n58993, n58994, n58995, n58996,
         n58997, n58998, n58999, n59000, n59001, n59002, n59003, n59004,
         n59005, n59006, n59007, n59008, n59009, n59010, n59011, n59012,
         n59013, n59014, n59015, n59016, n59017, n59018, n59019, n59020,
         n59021, n59022, n59023, n59024, n59025, n59026, n59027, n59028,
         n59029, n59030, n59031, n59032, n59033, n59034, n59035, n59036,
         n59037, n59038, n59039, n59040, n59041, n59042, n59043, n59044,
         n59045, n59046, n59047, n59048, n59049, n59050, n59051, n59052,
         n59053, n59054, n59055, n59056, n59057, n59058, n59059, n59060,
         n59061, n59062, n59063, n59064, n59065, n59066, n59067, n59068,
         n59069, n59070, n59071, n59072, n59073, n59074, n59075, n59076,
         n59077, n59078, n59079, n59080, n59081, n59082, n59083, n59084,
         n59085, n59086, n59087, n59088, n59089, n59090, n59091, n59092,
         n59093, n59094, n59095, n59096, n59097, n59098, n59099, n59100,
         n59101, n59102, n59103, n59104, n59105, n59106, n59107, n59108,
         n59109, n59110, n59111, n59112, n59113, n59114, n59115, n59116,
         n59117, n59118, n59119, n59120, n59121, n59122, n59123, n59124,
         n59125, n59126, n59127, n59128, n59129, n59130, n59131, n59132,
         n59133, n59134, n59135, n59136, n59137, n59138, n59139, n59140,
         n59141, n59142, n59143, n59144, n59145, n59146, n59147, n59148,
         n59149, n59150, n59151, n59152, n59153, n59154, n59155, n59156,
         n59157, n59158, n59159, n59160, n59161, n59162, n59163, n59164,
         n59165, n59166, n59167, n59168, n59169, n59170, n59171, n59172,
         n59173, n59174, n59175, n59176, n59177, n59178, n59179, n59180,
         n59181, n59182, n59183, n59184, n59185, n59186, n59187, n59188,
         n59189, n59190, n59191, n59192, n59193, n59194, n59195, n59196,
         n59197, n59198, n59199, n59200, n59201, n59202, n59203, n59204,
         n59205, n59206, n59207, n59208, n59209, n59210, n59211, n59212,
         n59213, n59214, n59215, n59216, n59217, n59218, n59219, n59220,
         n59221, n59222, n59223, n59224, n59225, n59226, n59227, n59228,
         n59229, n59230, n59231, n59232, n59233, n59234, n59235, n59236,
         n59237, n59238, n59239, n59240, n59241, n59242, n59243, n59244,
         n59245, n59246, n59247, n59248, n59249, n59250, n59251, n59252,
         n59253, n59254, n59255, n59256, n59257, n59258, n59259, n59260,
         n59261, n59262, n59263, n59264, n59265, n59266, n59267, n59268,
         n59269, n59270, n59271, n59272, n59273, n59274, n59275, n59276,
         n59277, n59278, n59279, n59280, n59281, n59282, n59283, n59284,
         n59285, n59286, n59287, n59288, n59289, n59290, n59291, n59292,
         n59293, n59294, n59295, n59296, n59297, n59298, n59299, n59300,
         n59301, n59302, n59303, n59304, n59305, n59306, n59307, n59308,
         n59309, n59310, n59311, n59312, n59313, n59314, n59315, n59316,
         n59317, n59318, n59319, n59320, n59321, n59322, n59323, n59324,
         n59325, n59326, n59327, n59328, n59329, n59330, n59331, n59332,
         n59333, n59334, n59335, n59336, n59337, n59338, n59339, n59340,
         n59341, n59342, n59343, n59344, n59345, n59346, n59347, n59348,
         n59349, n59350, n59351, n59352, n59353, n59354, n59355, n59356,
         n59357, n59358, n59359, n59360, n59361, n59362, n59363, n59364,
         n59365, n59366, n59367, n59368, n59369, n59370, n59371, n59372,
         n59373, n59374, n59375, n59376, n59377, n59378, n59379, n59380,
         n59381, n59382, n59383, n59384, n59385, n59386, n59387, n59388,
         n59389, n59390, n59391, n59392, n59393, n59394, n59395, n59396,
         n59397, n59398, n59399, n59400, n59401, n59402, n59403, n59404,
         n59405, n59406, n59407, n59408, n59409, n59410, n59411, n59412,
         n59413, n59414, n59415, n59416, n59417, n59418, n59419, n59420,
         n59421, n59422, n59423, n59424, n59425, n59426, n59427, n59428,
         n59429, n59430, n59431, n59432, n59433, n59434, n59435, n59436,
         n59437, n59438, n59439, n59440, n59441, n59442, n59443, n59444,
         n59445, n59446, n59447, n59448, n59449, n59450, n59451, n59452,
         n59453, n59454, n59455, n59456, n59457, n59458, n59459, n59460,
         n59461, n59462, n59463, n59464, n59465, n59466, n59467, n59468,
         n59469, n59470, n59471, n59472, n59473, n59474, n59475, n59476,
         n59477, n59478, n59479, n59480, n59481, n59482, n59483, n59484,
         n59485, n59486, n59487, n59488, n59489, n59490, n59491, n59492,
         n59493, n59494, n59495, n59496, n59497, n59498, n59499, n59500,
         n59501, n59502, n59503, n59504, n59505, n59506, n59507, n59508,
         n59509, n59510, n59511, n59512, n59513, n59514, n59515, n59516,
         n59517, n59518, n59519, n59520, n59521, n59522, n59523, n59524,
         n59525, n59526, n59527, n59528, n59529, n59530, n59531, n59532,
         n59533, n59534, n59535, n59536, n59537, n59538, n59539, n59540,
         n59541, n59542, n59543, n59544, n59545, n59546, n59547, n59548,
         n59549, n59550, n59551, n59552, n59553, n59554, n59555, n59556,
         n59557, n59558, n59559, n59560, n59561, n59562, n59563, n59564,
         n59565, n59566, n59567, n59568, n59569, n59570, n59571, n59572,
         n59573, n59574, n59575, n59576, n59577, n59578, n59579, n59580,
         n59581, n59582, n59583, n59584, n59585, n59586, n59587, n59588,
         n59589, n59590, n59591, n59592, n59593, n59594, n59595, n59596,
         n59597, n59598, n59599, n59600, n59601, n59602, n59603, n59604,
         n59605, n59606, n59607, n59608, n59609, n59610, n59611, n59612,
         n59613, n59614, n59615, n59616, n59617, n59618, n59619, n59620,
         n59621, n59622, n59623, n59624, n59625, n59626, n59627, n59628,
         n59629, n59630, n59631, n59632, n59633, n59634, n59635, n59636,
         n59637, n59638, n59639, n59640, n59641, n59642, n59643, n59644,
         n59645, n59646, n59647, n59648, n59649, n59650, n59651, n59652,
         n59653, n59654, n59655, n59656, n59657, n59658, n59659, n59660,
         n59661, n59662, n59663, n59664, n59665, n59666, n59667, n59668,
         n59669, n59670, n59671, n59672, n59673, n59674, n59675, n59676,
         n59677, n59678, n59679, n59680, n59681, n59682, n59683, n59684,
         n59685, n59686, n59687, n59688, n59689, n59690, n59691, n59692,
         n59693, n59694, n59695, n59696, n59697, n59698, n59699, n59700,
         n59701, n59702, n59703, n59704, n59705, n59706, n59707, n59708,
         n59709, n59710, n59711, n59712, n59713, n59714, n59715, n59716,
         n59717, n59718, n59719, n59720, n59721, n59722, n59723, n59724,
         n59725, n59726, n59727, n59728, n59729, n59730, n59731, n59732,
         n59733, n59734, n59735, n59736, n59737, n59738, n59739, n59740,
         n59741, n59742, n59743, n59744, n59745, n59746, n59747, n59748,
         n59749, n59750, n59751, n59752, n59753, n59754, n59755, n59756,
         n59757, n59758, n59759, n59760, n59761, n59762, n59763, n59764,
         n59765, n59766, n59767, n59768, n59769, n59770, n59771, n59772,
         n59773, n59774, n59775, n59776, n59777, n59778, n59779, n59780,
         n59781, n59782, n59783, n59784, n59785, n59786, n59787, n59788,
         n59789, n59790, n59791, n59792, n59793, n59794, n59795, n59796,
         n59797, n59798, n59799, n59800, n59801, n59802, n59803, n59804,
         n59805, n59806, n59807, n59808, n59809, n59810, n59811, n59812,
         n59813, n59814, n59815, n59816, n59817, n59818, n59819, n59820,
         n59821, n59822, n59823, n59824, n59825, n59826, n59827, n59828,
         n59829, n59830, n59831, n59832, n59833, n59834, n59835, n59836,
         n59837, n59838, n59839, n59840, n59841, n59842, n59843, n59844,
         n59845, n59846, n59847, n59848, n59849, n59850, n59851, n59852,
         n59853, n59854, n59855, n59856, n59857, n59858, n59859, n59860,
         n59861, n59862, n59863, n59864, n59865, n59866, n59867, n59868,
         n59869, n59870, n59871, n59872, n59873, n59874, n59875, n59876,
         n59877, n59878, n59879, n59880, n59881, n59882, n59883, n59884,
         n59885, n59886, n59887, n59888, n59889, n59890, n59891, n59892,
         n59893, n59894, n59895, n59896, n59897, n59898, n59899, n59900,
         n59901, n59902, n59903, n59904, n59905, n59906, n59907, n59908,
         n59909, n59910, n59911, n59912, n59913, n59914, n59915, n59916,
         n59917, n59918, n59919, n59920, n59921, n59922, n59923, n59924,
         n59925, n59926, n59927, n59928, n59929, n59930, n59931, n59932,
         n59933, n59934, n59935, n59936, n59937, n59938, n59939, n59940,
         n59941, n59942, n59943, n59944, n59945, n59946, n59947, n59948,
         n59949, n59950, n59951, n59952, n59953, n59954, n59955, n59956,
         n59957, n59958, n59959, n59960, n59961, n59962, n59963, n59964,
         n59965, n59966, n59967, n59968, n59969, n59970, n59971, n59972,
         n59973, n59974, n59975, n59976, n59977, n59978, n59979, n59980,
         n59981, n59982, n59983, n59984, n59985, n59986, n59987, n59988,
         n59989, n59990, n59991, n59992, n59993, n59994, n59995, n59996,
         n59997, n59998, n59999, n60000, n60001, n60002, n60003, n60004,
         n60005, n60006, n60007, n60008, n60009, n60010, n60011, n60012,
         n60013, n60014, n60015, n60016, n60017, n60018, n60019, n60020,
         n60021, n60022, n60023, n60024, n60025, n60026, n60027, n60028,
         n60029, n60030, n60031, n60032, n60033, n60034, n60035, n60036,
         n60037, n60038, n60039, n60040, n60041, n60042, n60043, n60044,
         n60045, n60046, n60047, n60048, n60049, n60050, n60051, n60052,
         n60053, n60054, n60055, n60056, n60057, n60058, n60059, n60060,
         n60061, n60062, n60063, n60064, n60065, n60066, n60067, n60068,
         n60069, n60070, n60071, n60072, n60073, n60074, n60075, n60076,
         n60077, n60078, n60079, n60080, n60081, n60082, n60083, n60084,
         n60085, n60086, n60087, n60088, n60089, n60090, n60091, n60092,
         n60093, n60094, n60095, n60096, n60097, n60098, n60099, n60100,
         n60101, n60102, n60103, n60104, n60105, n60106, n60107, n60108,
         n60109, n60110, n60111, n60112, n60113, n60114, n60115, n60116,
         n60117, n60118, n60119, n60120, n60121, n60122, n60123, n60124,
         n60125, n60126, n60127, n60128, n60129, n60130, n60131, n60132,
         n60133, n60134, n60135, n60136, n60137, n60138, n60139, n60140,
         n60141, n60142, n60143, n60144, n60145, n60146, n60147, n60148,
         n60149, n60150, n60151, n60152, n60153, n60154, n60155, n60156,
         n60157, n60158, n60159, n60160, n60161, n60162, n60163, n60164,
         n60165, n60166, n60167, n60168, n60169, n60170, n60171, n60172,
         n60173, n60174, n60175, n60176, n60177, n60178, n60179, n60180,
         n60181, n60182, n60183, n60184, n60185, n60186, n60187, n60188,
         n60189, n60190, n60191, n60192, n60193, n60194, n60195, n60196,
         n60197, n60198, n60199, n60200, n60201, n60202, n60203, n60204,
         n60205, n60206, n60207, n60208, n60209, n60210, n60211, n60212,
         n60213, n60214, n60215, n60216, n60217, n60218, n60219, n60220,
         n60221, n60222, n60223, n60224, n60225, n60226, n60227, n60228,
         n60229, n60230, n60231, n60232, n60233, n60234, n60235, n60236,
         n60237, n60238, n60239, n60240, n60241, n60242, n60243, n60244,
         n60245, n60246, n60247, n60248, n60249, n60250, n60251, n60252,
         n60253, n60254, n60255, n60256, n60257, n60258, n60259, n60260,
         n60261, n60262, n60263, n60264, n60265, n60266, n60267, n60268,
         n60269, n60270, n60271, n60272, n60273, n60274, n60275, n60276,
         n60277, n60278, n60279, n60280, n60281, n60282, n60283, n60284,
         n60285, n60286, n60287, n60288, n60289, n60290, n60291, n60292,
         n60293, n60294, n60295, n60296, n60297, n60298, n60299, n60300,
         n60301, n60302, n60303, n60304, n60305, n60306, n60307, n60308,
         n60309, n60310, n60311, n60312, n60313, n60314, n60315, n60316,
         n60317, n60318, n60319, n60320, n60321, n60322, n60323, n60324,
         n60325, n60326, n60327, n60328, n60329, n60330, n60331, n60332,
         n60333, n60334, n60335, n60336, n60337, n60338, n60339, n60340,
         n60341, n60342, n60343, n60344, n60345, n60346, n60347, n60348,
         n60349, n60350, n60351, n60352, n60353, n60354, n60355, n60356,
         n60357, n60358, n60359, n60360, n60361, n60362, n60363, n60364,
         n60365, n60366, n60367, n60368, n60369, n60370, n60371, n60372,
         n60373, n60374, n60375, n60376, n60377, n60378, n60379, n60380,
         n60381, n60382, n60383, n60384, n60385, n60386, n60387, n60388,
         n60389, n60390, n60391, n60392, n60393, n60394, n60395, n60396,
         n60397, n60398, n60399, n60400, n60401, n60402, n60403, n60404,
         n60405, n60406, n60407, n60408, n60409, n60410, n60411, n60412,
         n60413, n60414, n60415, n60416, n60417, n60418, n60419, n60420,
         n60421, n60422, n60423, n60424, n60425, n60426, n60427, n60428,
         n60429, n60430, n60431, n60432, n60433, n60434, n60435, n60436,
         n60437, n60438, n60439, n60440, n60441, n60442, n60443, n60444,
         n60445, n60446, n60447, n60448, n60449, n60450, n60451, n60452,
         n60453, n60454, n60455, n60456, n60457, n60458, n60459, n60460,
         n60461, n60462, n60463, n60464, n60465, n60466, n60467, n60468,
         n60469, n60470, n60471, n60472, n60473, n60474, n60475, n60476,
         n60477, n60478, n60479, n60480, n60481, n60482, n60483, n60484,
         n60485, n60486, n60487, n60488, n60489, n60490, n60491, n60492,
         n60493, n60494, n60495, n60496, n60497, n60498, n60499, n60500,
         n60501, n60502, n60503, n60504, n60505, n60506, n60507, n60508,
         n60509, n60510, n60511, n60512, n60513, n60514, n60515, n60516,
         n60517, n60518, n60519, n60520, n60521, n60522, n60523, n60524,
         n60525, n60526, n60527, n60528, n60529, n60530, n60531, n60532,
         n60533, n60534, n60535, n60536, n60537, n60538, n60539, n60540,
         n60541, n60542, n60543, n60544, n60545, n60546, n60547, n60548,
         n60549, n60550, n60551, n60552, n60553, n60554, n60555, n60556,
         n60557, n60558, n60559, n60560, n60561, n60562, n60563, n60564,
         n60565, n60566, n60567, n60568, n60569, n60570, n60571, n60572,
         n60573, n60574, n60575, n60576, n60577, n60578, n60579, n60580,
         n60581, n60582, n60583, n60584, n60585, n60586, n60587, n60588,
         n60589, n60590, n60591, n60592, n60593, n60594, n60595, n60596,
         n60597, n60598, n60599, n60600, n60601, n60602, n60603, n60604,
         n60605, n60606, n60607, n60608, n60609, n60610, n60611, n60612,
         n60613, n60614, n60615, n60616, n60617, n60618, n60619, n60620,
         n60621, n60622, n60623, n60624, n60625, n60626, n60627, n60628,
         n60629, n60630, n60631, n60632, n60633, n60634, n60635, n60636,
         n60637, n60638, n60639, n60640, n60641, n60642, n60643, n60644,
         n60645, n60646, n60647, n60648, n60649, n60650, n60651, n60652,
         n60653, n60654, n60655, n60656, n60657, n60658, n60659, n60660,
         n60661, n60662, n60663, n60664, n60665, n60666, n60667, n60668,
         n60669, n60670, n60671, n60672, n60673, n60674, n60675, n60676,
         n60677, n60678, n60679, n60680, n60681, n60682, n60683, n60684,
         n60685, n60686, n60687, n60688, n60689, n60690, n60691, n60692,
         n60693, n60694, n60695, n60696, n60697, n60698, n60699, n60700,
         n60701, n60702, n60703, n60704, n60705, n60706, n60707, n60708,
         n60709, n60710, n60711, n60712, n60713, n60714, n60715, n60716,
         n60717, n60718, n60719, n60720, n60721, n60722, n60723, n60724,
         n60725, n60726, n60727, n60728, n60729, n60730, n60731, n60732,
         n60733, n60734, n60735, n60736, n60737, n60738, n60739, n60740,
         n60741, n60742, n60743, n60744, n60745, n60746, n60747, n60748,
         n60749, n60750, n60751, n60752, n60753, n60754, n60755, n60756,
         n60757, n60758, n60759, n60760, n60761, n60762, n60763, n60764,
         n60765, n60766, n60767, n60768, n60769, n60770, n60771, n60772,
         n60773, n60774, n60775, n60776, n60777, n60778, n60779, n60780,
         n60781, n60782, n60783, n60784, n60785, n60786, n60787, n60788,
         n60789, n60790, n60791, n60792, n60793, n60794, n60795, n60796,
         n60797, n60798, n60799, n60800, n60801, n60802, n60803, n60804,
         n60805, n60806, n60807, n60808, n60809, n60810, n60811, n60812,
         n60813, n60814, n60815, n60816, n60817, n60818, n60819, n60820,
         n60821, n60822, n60823, n60824, n60825, n60826, n60827, n60828,
         n60829, n60830, n60831, n60832, n60833, n60834, n60835, n60836,
         n60837, n60838, n60839, n60840, n60841, n60842, n60843, n60844,
         n60845, n60846, n60847, n60848, n60849, n60850, n60851, n60852,
         n60853, n60854, n60855, n60856, n60857, n60858, n60859, n60860,
         n60861, n60862, n60863, n60864, n60865, n60866, n60867, n60868,
         n60869, n60870, n60871, n60872, n60873, n60874, n60875, n60876,
         n60877, n60878, n60879, n60880, n60881, n60882, n60883, n60884,
         n60885, n60886, n60887, n60888, n60889, n60890, n60891, n60892,
         n60893, n60894, n60895, n60896, n60897, n60898, n60899, n60900,
         n60901, n60902, n60903, n60904, n60905, n60906, n60907, n60908,
         n60909, n60910, n60911, n60912, n60913, n60914, n60915, n60916,
         n60917, n60918, n60919, n60920, n60921, n60922, n60923, n60924,
         n60925, n60926, n60927, n60928, n60929, n60930, n60931, n60932,
         n60933, n60934, n60935, n60936, n60937, n60938, n60939, n60940,
         n60941, n60942, n60943, n60944, n60945, n60946, n60947, n60948,
         n60949, n60950, n60951, n60952, n60953, n60954, n60955, n60956,
         n60957, n60958, n60959, n60960, n60961, n60962, n60963, n60964,
         n60965, n60966, n60967, n60968, n60969, n60970, n60971, n60972,
         n60973, n60974, n60975, n60976, n60977, n60978, n60979, n60980,
         n60981, n60982, n60983, n60984, n60985, n60986, n60987, n60988,
         n60989, n60990, n60991, n60992, n60993, n60994, n60995, n60996,
         n60997, n60998, n60999, n61000, n61001, n61002, n61003, n61004,
         n61005, n61006, n61007, n61008, n61009, n61010, n61011, n61012,
         n61013, n61014, n61015, n61016, n61017, n61018, n61019, n61020,
         n61021, n61022, n61023, n61024, n61025, n61026, n61027, n61028,
         n61029, n61030, n61031, n61032, n61033, n61034, n61035, n61036,
         n61037, n61038, n61039, n61040, n61041, n61042, n61043, n61044,
         n61045, n61046, n61047, n61048, n61049, n61050, n61051, n61052,
         n61053, n61054, n61055, n61056, n61057, n61058, n61059, n61060,
         n61061, n61062, n61063, n61064, n61065, n61066, n61067, n61068,
         n61069, n61070, n61071, n61072, n61073, n61074, n61075, n61076,
         n61077, n61078, n61079, n61080, n61081, n61082, n61083, n61084,
         n61085, n61086, n61087, n61088, n61089, n61090, n61091, n61092,
         n61093, n61094, n61095, n61096, n61097, n61098, n61099, n61100,
         n61101, n61102, n61103, n61104, n61105, n61106, n61107, n61108,
         n61109, n61110, n61111, n61112, n61113, n61114, n61115, n61116,
         n61117, n61118, n61119, n61120, n61121, n61122, n61123, n61124,
         n61125, n61126, n61127, n61128, n61129, n61130, n61131, n61132,
         n61133, n61134, n61135, n61136, n61137, n61138, n61139, n61140,
         n61141, n61142, n61143, n61144, n61145, n61146, n61147, n61148,
         n61149, n61150, n61151, n61152, n61153, n61154, n61155, n61156,
         n61157, n61158, n61159, n61160, n61161, n61162, n61163, n61164,
         n61165, n61166, n61167, n61168, n61169, n61170, n61171, n61172,
         n61173, n61174, n61175, n61176, n61177, n61178, n61179, n61180,
         n61181, n61182, n61183, n61184, n61185, n61186, n61187, n61188,
         n61189, n61190, n61191, n61192, n61193, n61194, n61195, n61196,
         n61197, n61198, n61199, n61200, n61201, n61202, n61203, n61204,
         n61205, n61206, n61207, n61208, n61209, n61210, n61211, n61212,
         n61213, n61214, n61215, n61216, n61217, n61218, n61219, n61220,
         n61221, n61222, n61223, n61224, n61225, n61226, n61227, n61228,
         n61229, n61230, n61231, n61232, n61233, n61234, n61235, n61236,
         n61237, n61238, n61239, n61240, n61241, n61242, n61243, n61244,
         n61245, n61246, n61247, n61248, n61249, n61250, n61251, n61252,
         n61253, n61254, n61255, n61256, n61257, n61258, n61259, n61260,
         n61261, n61262, n61263, n61264, n61265, n61266, n61267, n61268,
         n61269, n61270, n61271, n61272, n61273, n61274, n61275, n61276,
         n61277, n61278, n61279, n61280, n61281, n61282, n61283, n61284,
         n61285, n61286, n61287, n61288, n61289, n61290, n61291, n61292,
         n61293, n61294, n61295, n61296, n61297, n61298, n61299, n61300,
         n61301, n61302, n61303, n61304, n61305, n61306, n61307, n61308,
         n61309, n61310, n61311, n61312, n61313, n61314, n61315, n61316,
         n61317, n61318, n61319, n61320, n61321, n61322, n61323, n61324,
         n61325, n61326, n61327, n61328, n61329, n61330, n61331, n61332,
         n61333, n61334, n61335, n61336, n61337, n61338, n61339, n61340,
         n61341, n61342, n61343, n61344, n61345, n61346, n61347, n61348,
         n61349, n61350, n61351, n61352, n61353, n61354, n61355, n61356,
         n61357, n61358, n61359, n61360, n61361, n61362, n61363, n61364,
         n61365, n61366, n61367, n61368, n61369, n61370, n61371, n61372,
         n61373, n61374, n61375, n61376, n61377, n61378, n61379, n61380,
         n61381, n61382, n61383, n61384, n61385, n61386, n61387, n61388,
         n61389, n61390, n61391, n61392, n61393, n61394, n61395, n61396,
         n61397, n61398, n61399, n61400, n61401, n61402, n61403, n61404,
         n61405, n61406, n61407, n61408, n61409, n61410, n61411, n61412,
         n61413, n61414, n61415, n61416, n61417, n61418, n61419, n61420,
         n61421, n61422, n61423, n61424, n61425, n61426, n61427, n61428,
         n61429, n61430, n61431, n61432, n61433, n61434, n61435, n61436,
         n61437, n61438, n61439, n61440, n61441, n61442, n61443, n61444,
         n61445, n61446, n61447, n61448, n61449, n61450, n61451, n61452,
         n61453, n61454, n61455, n61456, n61457, n61458, n61459, n61460,
         n61461, n61462, n61463, n61464, n61465, n61466, n61467, n61468,
         n61469, n61470, n61471, n61472, n61473, n61474, n61475, n61476,
         n61477, n61478, n61479, n61480, n61481, n61482, n61483, n61484,
         n61485, n61486, n61487, n61488, n61489, n61490, n61491, n61492,
         n61493, n61494, n61495, n61496, n61497, n61498, n61499, n61500,
         n61501, n61502, n61503, n61504, n61505, n61506, n61507, n61508,
         n61509, n61510, n61511, n61512, n61513, n61514, n61515, n61516,
         n61517, n61518, n61519, n61520, n61521, n61522, n61523, n61524,
         n61525, n61526, n61527, n61528, n61529, n61530, n61531, n61532,
         n61533, n61534, n61535, n61536, n61537, n61538, n61539, n61540,
         n61541, n61542, n61543, n61544, n61545, n61546, n61547, n61548,
         n61549, n61550, n61551, n61552, n61553, n61554, n61555, n61556,
         n61557, n61558, n61559, n61560, n61561, n61562, n61563, n61564,
         n61565, n61566, n61567, n61568, n61569, n61570, n61571, n61572,
         n61573, n61574, n61575, n61576, n61577, n61578, n61579, n61580,
         n61581, n61582, n61583, n61584, n61585, n61586, n61587, n61588,
         n61589, n61590, n61591, n61592, n61593, n61594, n61595, n61596,
         n61597, n61598, n61599, n61600, n61601, n61602, n61603, n61604,
         n61605, n61606, n61607, n61608, n61609, n61610, n61611, n61612,
         n61613, n61614, n61615, n61616, n61617, n61618, n61619, n61620,
         n61621, n61622, n61623, n61624, n61625, n61626, n61627, n61628,
         n61629, n61630, n61631, n61632, n61633, n61634, n61635, n61636,
         n61637, n61638, n61639, n61640, n61641, n61642, n61643, n61644,
         n61645, n61646, n61647, n61648, n61649, n61650, n61651, n61652,
         n61653, n61654, n61655, n61656, n61657, n61658, n61659, n61660,
         n61661, n61662, n61663, n61664, n61665, n61666, n61667, n61668,
         n61669, n61670, n61671, n61672, n61673, n61674, n61675, n61676,
         n61677, n61678, n61679, n61680, n61681, n61682, n61683, n61684,
         n61685, n61686, n61687, n61688, n61689, n61690, n61691, n61692,
         n61693, n61694, n61695, n61696, n61697, n61698, n61699, n61700,
         n61701, n61702, n61703, n61704, n61705, n61706, n61707, n61708,
         n61709, n61710, n61711, n61712, n61713, n61714, n61715, n61716,
         n61717, n61718, n61719, n61720, n61721, n61722, n61723, n61724,
         n61725, n61726, n61727, n61728, n61729, n61730, n61731, n61732,
         n61733, n61734, n61735, n61736, n61737, n61738, n61739, n61740,
         n61741, n61742, n61743, n61744, n61745, n61746, n61747, n61748,
         n61749, n61750, n61751, n61752, n61753, n61754, n61755, n61756,
         n61757, n61758, n61759, n61760, n61761, n61762, n61763, n61764,
         n61765, n61766, n61767, n61768, n61769, n61770, n61771, n61772,
         n61773, n61774, n61775, n61776, n61777, n61778, n61779, n61780,
         n61781, n61782, n61783, n61784, n61785, n61786, n61787, n61788,
         n61789, n61790, n61791, n61792, n61793, n61794, n61795, n61796,
         n61797, n61798, n61799, n61800, n61801, n61802, n61803, n61804,
         n61805, n61806, n61807, n61808, n61809, n61810, n61811, n61812,
         n61813, n61814, n61815, n61816, n61817, n61818, n61819, n61820,
         n61821, n61822, n61823, n61824, n61825, n61826, n61827, n61828,
         n61829, n61830, n61831, n61832, n61833, n61834, n61835, n61836,
         n61837, n61838, n61839, n61840, n61841, n61842, n61843, n61844,
         n61845, n61846, n61847, n61848, n61849, n61850, n61851, n61852,
         n61853, n61854, n61855, n61856, n61857, n61858, n61859, n61860,
         n61861, n61862, n61863, n61864, n61865, n61866, n61867, n61868,
         n61869, n61870, n61871, n61872, n61873, n61874, n61875, n61876,
         n61877, n61878, n61879, n61880, n61881, n61882, n61883, n61884,
         n61885, n61886, n61887, n61888, n61889, n61890, n61891, n61892,
         n61893, n61894, n61895, n61896, n61897, n61898, n61899, n61900,
         n61901, n61902, n61903, n61904, n61905, n61906, n61907, n61908,
         n61909, n61910, n61911, n67084, n67085, n67086, n67087, n67088,
         n67089, n67090, n67091, n67092, n67093, n67094, n67095, n67096,
         n67097, n67098, n67099, n67100, n67101, n67102, n67103, n67104,
         n67105, n67106, n67107, n67108, n67109, n67110, n67111, n67112,
         n67113, n67114, n67115, n67116, n67117, n67118, n67119, n67120,
         n67121, n67122, n67123, n67124, n67125, n67126, n67127, n67128,
         n67129, n67130, n67131, n67132, n67133, n67134, n67135, n67136,
         n67137, n67138, n67139, n67140, n67141, n67142, n67143, n67144,
         n67145, n67146, n67147, n67148, n67149, n67150, n67151, n67152,
         n67153, n67154, n67155, n67156, n67157, n67158, n67159, n67160,
         n67161, n67162, n67163, n67164, n67165, n67166, n67167, n67168,
         n67169, n67170, n67171, n67172, n67173, n67174, n67175, n67176,
         n67177, n67178, n67179, n67180, n67181, n67182, n67183, n67184,
         n67185, n67186, n67187, n67188, n67189, n67190, n67191, n67192,
         n67193, n67194, n67195, n67196, n67197, n67198, n67199, n67200,
         n67201, n67202, n67203, n67204, n67205, n67206, n67207, n67208,
         n67209, n67210, n67211, n67212, n67213, n67214, n67215, n67216,
         n67217, n67218, n67219, n67220, n67221, n67222, n67223, n67224,
         n67225, n67226, n67227, n67228, n67229, n67230, n67231, n67232,
         n67233, n67234, n67235, n67236, n67237, n67238, n67239, n67240,
         n67241, n67242, n67243, n67244, n67245, n67246, n67247, n67248,
         n67249, n67250, n67251, n67252, n67253, n67254, n67255, n67256,
         n67257, n67258, n67259, n67260, n67261, n67262, n67263, n67264,
         n67265, n67266, n67267, n67268, n67269, n67270, n67271, n67272,
         n67273, n67274, n67275, n67276, n67277, n67278, n67279, n67280,
         n67281, n67282, n67283, n67284, n67285, n67286, n67287, n67288,
         n67289, n67290, n67291, n67292, n67293, n67294, n67295, n67296,
         n67297, n67298, n67299, n67300, n67301, n67302, n67303, n67304,
         n67305, n67306, n67307, n67308, n67309, n67310, n67311, n67312,
         n67313, n67314, n67315, n67316, n67317, n67318, n67319, n67320,
         n67321, n67322, n67323, n67324, n67325, n67326, n67327, n67328,
         n67329, n67330, n67331, n67332, n67333, n67334, n67335, n67336,
         n67337, n67338, n67339, n67340, n67341, n67342, n67343, n67344,
         n67345, n67346, n67347, n67348, n67349, n67350, n67351, n67352,
         n67353, n67354, n67355, n67356, n67357, n67358, n67359, n67360,
         n67361, n67362, n67363, n67364, n67365, n67366, n67367, n67368,
         n67369, n67370, n67371, n67372, n67373, n67374, n67375, n67376,
         n67377, n67378, n67379, n67380, n67381, n67382, n67383, n67384,
         n67385, n67386, n67387, n67388, n67389, n67390, n67391, n67392,
         n67393, n67394, n67395, n67396, n67397, n67398, n67399, n67400,
         n67401, n67402, n67403, n67404, n67405, n67406, n67407, n67408,
         n67409, n67410, n67411, n67412, n67413, n67414, n67415, n67416,
         n67417, n67418, n67419, n67420, n67421, n67422, n67423, n67424,
         n67425, n67426, n67427, n67428, n67429, n67430, n67431, n67432,
         n67433, n67434, n67435, n67436, n67437, n67438, n67439, n67440,
         n67441, n67442, n67443, n67444, n67445, n67446, n67447, n67448,
         n67449, n67450, n67451, n67452, n67453, n67454, n67455, n67456,
         n67457, n67458, n67459, n67460, n67461, n67462, n67463, n67464,
         n67465, n67466, n67467, n67468, n67469, n67470, n67471, n67472,
         n67473, n67474, n67475, n67476, n67477, n67478, n67479, n67480,
         n67481, n67482, n67483, n67484, n67485, n67486, n67487, n67488,
         n67489, n67490, n67491, n67492, n67493, n67494, n67495, n67496,
         n67497, n67498, n67499, n67500, n67501, n67502, n67503, n67504,
         n67505, n67506, n67507, n67508, n67509, n67510, n67511, n67512,
         n67513, n67514, n67515, n67516, n67517, n67518, n67519, n67520,
         n67521, n67522, n67523, n67524, n67525, n67526, n67527, n67528,
         n67529, n67530, n67531, n67532, n67533, n67534, n67535, n67536,
         n67537, n67538, n67539, n67540, n67541, n67542, n67543, n67544,
         n67545, n67546, n67547, n67548, n67549, n67550, n67551, n67552,
         n67553, n67554, n67555, n67556, n67557, n67558, n67559, n67560,
         n67561, n67562, n67563, n67564, n67565, n67566, n67567, n67568,
         n67569, n67570, n67571, n67572, n67573, n67574, n67575, n67576,
         n67577, n67578, n67579, n67580, n67581, n67582, n67583, n67584,
         n67585, n67586, n67587, n67588, n67589, n67590, n67591, n67592,
         n67593, n67594, n67595, n67596, n67597, n67598, n67599, n67600,
         n67601, n67602, n67603, n67604, n67605, n67606, n67607, n67608,
         n67609, n67610, n67611, n67612, n67613, n67614, n67615, n67616,
         n67617, n67618, n67619, n67620, n67621, n67622, n67623, n67624,
         n67625, n67626, n67627, n67628, n67629, n67630, n67631, n67632,
         n67633, n67634, n67635, n67636, n67637, n67638, n67639, n67640,
         n67641, n67642, n67643, n67644, n67645, n67646, n67647, n67648,
         n67649, n67650, n67651, n67652, n67653, n67654, n67655, n67656,
         n67657, n67658, n67659, n67660, n67661, n67662, n67663, n67664,
         n67665, n67666, n67667, n67668, n67669, n67670, n67671, n67672,
         n67673, n67674, n67675, n67676, n67677, n67678, n67679, n67680,
         n67681, n67682, n67683, n67684, n67685, n67686, n67687, n67688,
         n67689, n67690, n67691, n67692, n67693, n67694, n67695, n67696,
         n67697, n67698, n67699, n67700, n67701, n67702, n67703, n67704,
         n67705, n67706, n67707, n67708, n67709, n67710, n67711, n67712,
         n67713, n67714, n67715, n67716, n67717, n67718, n67719, n67720,
         n67721, n67722, n67723, n67724, n67725, n67726, n67727, n67728,
         n67729, n67730, n67731, n67732, n67733, n67734, n67735, n67736,
         n67737, n67738, n67739, n67740, n67741, n67742, n67743, n67744,
         n67745, n67746, n67747, n67748, n67749, n67750, n67751, n67752,
         n67753, n67754, n67755, n67756, n67757, n67758, n67759, n67760,
         n67761, n67762, n67763, n67764, n67765, n67766, n67767, n67768,
         n67769, n67770, n67771, n67772, n67773, n67774, n67775, n67776,
         n67777, n67778, n67779, n67780, n67781, n67782, n67783, n67784,
         n67785, n67786, n67787, n67788, n67789, n67790, n67791, n67792,
         n67793, n67794, n67795, n67796, n67797, n67798, n67799, n67800,
         n67801, n67802, n67803, n67804, n67805, n67806, n67807, n67808,
         n67809, n67810, n67811, n67812, n67813, n67814, n67815, n67816,
         n67817, n67818, n67819, n67820, n67821, n67822, n67823, n67824,
         n67825, n67826, n67827, n67828, n67829, n67830, n67831, n67832,
         n67833, n67834, n67835, n67836, n67837, n67838, n67839, n67840,
         n67841, n67842, n67843, n67844, n67845, n67846, n67847, n67848,
         n67849, n67850, n67851, n67852, n67853, n67854, n67855, n67856,
         n67857, n67858, n67859, n67860, n67861, n67862, n67863, n67864,
         n67865, n67866, n67867, n67868, n67869, n67870, n67871, n67872,
         n67873, n67874, n67875, n67876, n67877, n67878, n67879, n67880,
         n67881, n67882, n67883, n67884, n67885, n67886, n67887, n67888,
         n67889, n67890, n67891, n67892, n67893, n67894, n67895, n67896,
         n67897, n67898, n67899, n67900, n67901, n67902, n67903, n67904,
         n67905, n67906, n67907, n67908, n67909, n67910, n67911, n67912,
         n67913, n67914, n67915, n67916, n67917, n67918, n67919, n67920,
         n67921, n67922, n67923, n67924, n67925, n67926, n67927, n67928,
         n67929, n67930, n67931, n67932, n67933, n67934, n67935, n67936,
         n67937, n67938, n67939, n67940, n67941, n67942, n67943, n67944,
         n67945, n67946, n67947, n67948, n67949, n67950, n67951, n67952,
         n67953, n67954, n67955, n67956, n67957, n67958, n67959, n67960,
         n67961, n67962, n67963, n67964, n67965, n67966, n67967, n67968,
         n67969, n67970, n67971, n67972, n67973, n67974, n67975, n67976,
         n67977, n67978, n67979, n67980, n67981, n67982, n67983, n67984,
         n67985, n67986, n67987, n67988, n67989, n67990, n67991, n67992,
         n67993, n67994, n67995, n67996, n67997, n67998, n67999, n68000,
         n68001, n68002, n68003, n68004, n68005, n68006, n68007, n68008,
         n68009, n68010, n68011, n68012, n68013, n68014, n68015, n68016,
         n68017, n68018, n68019, n68020, n68021, n68022, n68023, n68024,
         n68025, n68026, n68027, n68028, n68029, n68030, n68031, n68032,
         n68033, n68034, n68035, n68036, n68037, n68038, n68039, n68040,
         n68041, n68042, n68043, n68044, n68045, n68046, n68047, n68048,
         n68049, n68050, n68051, n68052, n68053, n68054, n68055, n68056,
         n68057, n68058, n68059, n68060, n68061, n68062, n68063, n68064,
         n68065, n68066, n68067, n68068, n68069, n68070, n68071, n68072,
         n68073, n68074, n68075, n68076, n68077, n68078, n68079, n68080,
         n68081, n68082, n68083, n68084, n68085, n68086, n68087, n68088,
         n68089, n68090, n68091, n68092, n68093, n68094, n68095, n68096,
         n68097, n68098, n68099, n68100, n68101, n68102, n68103, n68104,
         n68105, n68106, n68107, n68108, n68109, n68110, n68111, n68112,
         n68113, n68114, n68115, n68116, n68117, n68118, n68119, n68120,
         n68121, n68122, n68123, n68124, n68125, n68126, n68127, n68128,
         n68129, n68130, n68131, n68132, n68133, n68134, n68135, n68136,
         n68137, n68138, n68139, n68140, n68141, n68142, n68143, n68144,
         n68145, n68146, n68147, n68148, n68149, n68150, n68151, n68152,
         n68153, n68154, n68155, n68156, n68157, n68158, n68159, n68160,
         n68161, n68162, n68163, n68164, n68165, n68166, n68167, n68168,
         n68169, n68170, n68171, n68172, n68173, n68174, n68175, n68176,
         n68177, n68178, n68179, n68180, n68181, n68182, n68183, n68184,
         n68185, n68186, n68187, n68188, n68189, n68190, n68191, n68192,
         n68193, n68194, n68195, n68196, n68197, n68198, n68199, n68200,
         n68201, n68202, n68203, n68204, n68205, n68206, n68207, n68208,
         n68209, n68210, n68211, n68212, n68213, n68214, n68215, n68216,
         n68217, n68218, n68219, n68220, n68221, n68222, n68223, n68224,
         n68225, n68226, n68227, n68228, n68229, n68230, n68231, n68232,
         n68233, n68234, n68235, n68236, n68237, n68238, n68239, n68240,
         n68241, n68242, n68243, n68244, n68245, n68246, n68247, n68248,
         n68249, n68250, n68251, n68252, n68253, n68254, n68255, n68256,
         n68257, n68258, n68259, n68260, n68261, n68262, n68263, n68264,
         n68265, n68266, n68267, n68268, n68269, n68270, n68271, n68272,
         n68273, n68274, n68275, n68276, n68277, n68278, n68279, n68280,
         n68281, n68282, n68283, n68284, n68285, n68286, n68287, n68288,
         n68289, n68290, n68291, n68292, n68293, n68294, n68295, n68296,
         n68297, n68298, n68299, n68300, n68301, n68302, n68303, n68304,
         n68305, n68306, n68307, n68308, n68309, n68310, n68311, n68312,
         n68313, n68314, n68315, n68316, n68317, n68318, n68319, n68320,
         n68321, n68322, n68323, n68324, n68325, n68326, n68327, n68328,
         n68329, n68330, n68331, n68332, n68333, n68334, n68335, n68336,
         n68337, n68338, n68339, n68340, n68341, n68342, n68343, n68344,
         n68345, n68346, n68347, n68348, n68349, n68350, n68351, n68352,
         n68353, n68354, n68355, n68356, n68357, n68358, n68359, n68360,
         n68361, n68362, n68363, n68364, n68365, n68366, n68367, n68368,
         n68369, n68370, n68371, n68372, n68373, n68374, n68375, n68376,
         n68377, n68378, n68379, n68380, n68381, n68382, n68383, n68384,
         n68385, n68386, n68387, n68388, n68389, n68390, n68391, n68392,
         n68393, n68394, n68395, n68396, n68397, n68398, n68399, n68400,
         n68401, n68402, n68403, n68404, n68405, n68406, n68407, n68408,
         n68409, n68410, n68411, n68412, n68413, n68414, n68415, n68416,
         n68417, n68418, n68419, n68420, n68421, n68422, n68423, n68424,
         n68425, n68426, n68427, n68428, n68429, n68430, n68431, n68432,
         n68433, n68434, n68435, n68436, n68437, n68438, n68439, n68440,
         n68441, n68442, n68443, n68444, n68445, n68446, n68447, n68448,
         n68449, n68450, n68451, n68452, n68453, n68454, n68455, n68456,
         n68457, n68458, n68459, n68460, n68461, n68462, n68463, n68464,
         n68465, n68466, n68467, n68468, n68469, n68470, n68471, n68472,
         n68473, n68474, n68475, n68476, n68477, n68478, n68479, n68480,
         n68481, n68482, n68483, n68484, n68485, n68486, n68487, n68488,
         n68489, n68490, n68491, n68492, n68493, n68494, n68495, n68496,
         n68497, n68498, n68499, n68500, n68501, n68502, n68503, n68504,
         n68505, n68506, n68507, n68508, n68509, n68510, n68511, n68512,
         n68513, n68514, n68515, n68516, n68517, n68518, n68519, n68520,
         n68521, n68522, n68523, n68524, n68525, n68526, n68527, n68528,
         n68529, n68530, n68531, n68532, n68533, n68534, n68535, n68536,
         n68537, n68538, n68539, n68540, n68541, n68542, n68543, n68544,
         n68545, n68546, n68547, n68548, n68549, n68550, n68551, n68552,
         n68553, n68554, n68555, n68556, n68557, n68558, n68559, n68560,
         n68561, n68562, n68563, n68564, n68565, n68566, n68567, n68568,
         n68569, n68570, n68571, n68572, n68573, n68574, n68575, n68576,
         n68577, n68578, n68579, n68580, n68581, n68582, n68583, n68584,
         n68585, n68586, n68587, n68588, n68589, n68590, n68591;
  wire   [19:0] reg_i_0;
  wire   [19:0] reg_i_1;
  wire   [19:0] reg_i_2;
  wire   [19:0] reg_i_3;
  wire   [19:0] reg_i_4;
  wire   [19:0] reg_i_5;
  wire   [19:0] reg_i_6;
  wire   [19:0] reg_i_7;
  wire   [19:0] reg_i_8;
  wire   [19:0] reg_i_9;
  wire   [19:0] reg_i_10;
  wire   [19:0] reg_i_11;
  wire   [19:0] reg_i_12;
  wire   [19:0] reg_i_13;
  wire   [19:0] reg_i_14;
  wire   [19:0] reg_i_15;
  wire   [19:0] reg_w_0;
  wire   [19:0] reg_w_1;
  wire   [19:0] reg_w_2;
  wire   [19:0] reg_w_3;
  wire   [19:0] reg_w_4;
  wire   [19:0] reg_w_5;
  wire   [19:0] reg_w_6;
  wire   [19:0] reg_w_7;
  wire   [19:0] reg_w_8;
  wire   [19:0] reg_w_9;
  wire   [19:0] reg_w_10;
  wire   [19:0] reg_w_11;
  wire   [19:0] reg_w_12;
  wire   [19:0] reg_w_13;
  wire   [19:0] reg_w_14;
  wire   [19:0] reg_w_15;
  wire   [19:0] reg_ii_0;
  wire   [19:0] reg_ii_1;
  wire   [19:0] reg_ii_2;
  wire   [19:0] reg_ii_3;
  wire   [19:0] reg_ii_4;
  wire   [19:0] reg_ii_5;
  wire   [19:0] reg_ii_6;
  wire   [19:0] reg_ii_7;
  wire   [19:0] reg_ii_8;
  wire   [19:0] reg_ii_9;
  wire   [19:0] reg_ii_10;
  wire   [19:0] reg_ii_11;
  wire   [19:0] reg_ii_12;
  wire   [19:0] reg_ii_13;
  wire   [19:0] reg_ii_14;
  wire   [19:0] reg_ii_15;
  wire   [19:0] reg_ww_0;
  wire   [19:0] reg_ww_1;
  wire   [19:0] reg_ww_2;
  wire   [19:0] reg_ww_3;
  wire   [19:0] reg_ww_4;
  wire   [19:0] reg_ww_5;
  wire   [19:0] reg_ww_6;
  wire   [19:0] reg_ww_7;
  wire   [19:0] reg_ww_8;
  wire   [19:0] reg_ww_9;
  wire   [19:0] reg_ww_10;
  wire   [19:0] reg_ww_11;
  wire   [19:0] reg_ww_12;
  wire   [19:0] reg_ww_13;
  wire   [19:0] reg_ww_14;
  wire   [19:0] reg_ww_15;
  wire   [19:0] reg_iii_0;
  wire   [19:0] reg_iii_1;
  wire   [19:0] reg_iii_2;
  wire   [19:0] reg_iii_3;
  wire   [19:0] reg_iii_4;
  wire   [19:0] reg_iii_5;
  wire   [19:0] reg_iii_6;
  wire   [19:0] reg_iii_7;
  wire   [19:0] reg_iii_8;
  wire   [19:0] reg_iii_9;
  wire   [19:0] reg_iii_10;
  wire   [19:0] reg_iii_11;
  wire   [19:0] reg_iii_12;
  wire   [19:0] reg_iii_13;
  wire   [19:0] reg_iii_14;
  wire   [19:0] reg_iii_15;
  wire   [19:0] reg_www_0;
  wire   [19:0] reg_www_1;
  wire   [19:0] reg_www_2;
  wire   [19:0] reg_www_3;
  wire   [19:0] reg_www_4;
  wire   [19:0] reg_www_5;
  wire   [19:0] reg_www_6;
  wire   [19:0] reg_www_7;
  wire   [19:0] reg_www_8;
  wire   [19:0] reg_www_9;
  wire   [19:0] reg_www_10;
  wire   [19:0] reg_www_11;
  wire   [19:0] reg_www_12;
  wire   [19:0] reg_www_13;
  wire   [19:0] reg_www_14;
  wire   [19:0] reg_www_15;
  wire   [31:0] reg_i_mask;
  wire   [31:0] reg_w_mask;
  wire   [31:0] \mask_0/reg_ww_mask ;
  wire   [31:0] \mask_0/reg_ii_mask ;
  wire   [1:0] \mask_0/counter ;
  wire   [31:0] \mask_0/reg_w_mask ;
  wire   [31:0] \mask_0/reg_i_mask ;
  wire   [3:0] \filter_0/w_pointer ;
  wire   [3:0] \filter_0/i_pointer ;
  wire   [31:0] \filter_0/reg_xor_w_mask ;
  wire   [31:0] \filter_0/reg_xor_i_mask ;
  wire   [31:0] \filter_0/reg_o_mask ;
  wire   [19:0] \filter_0/reg_w_15 ;
  wire   [19:0] \filter_0/reg_w_14 ;
  wire   [19:0] \filter_0/reg_w_13 ;
  wire   [19:0] \filter_0/reg_w_12 ;
  wire   [19:0] \filter_0/reg_w_11 ;
  wire   [19:0] \filter_0/reg_w_10 ;
  wire   [19:0] \filter_0/reg_w_9 ;
  wire   [19:0] \filter_0/reg_w_8 ;
  wire   [19:0] \filter_0/reg_w_7 ;
  wire   [19:0] \filter_0/reg_w_6 ;
  wire   [19:0] \filter_0/reg_w_5 ;
  wire   [19:0] \filter_0/reg_w_4 ;
  wire   [19:0] \filter_0/reg_w_3 ;
  wire   [19:0] \filter_0/reg_w_2 ;
  wire   [19:0] \filter_0/reg_w_1 ;
  wire   [19:0] \filter_0/reg_w_0 ;
  wire   [19:0] \filter_0/reg_i_15 ;
  wire   [19:0] \filter_0/reg_i_14 ;
  wire   [19:0] \filter_0/reg_i_13 ;
  wire   [19:0] \filter_0/reg_i_12 ;
  wire   [19:0] \filter_0/reg_i_11 ;
  wire   [19:0] \filter_0/reg_i_10 ;
  wire   [19:0] \filter_0/reg_i_9 ;
  wire   [19:0] \filter_0/reg_i_8 ;
  wire   [19:0] \filter_0/reg_i_7 ;
  wire   [19:0] \filter_0/reg_i_6 ;
  wire   [19:0] \filter_0/reg_i_5 ;
  wire   [19:0] \filter_0/reg_i_4 ;
  wire   [19:0] \filter_0/reg_i_3 ;
  wire   [19:0] \filter_0/reg_i_2 ;
  wire   [19:0] \filter_0/reg_i_1 ;
  wire   [19:0] \filter_0/reg_i_0 ;
  wire   [3:0] \shifter_0/w_pointer ;
  wire   [3:0] \shifter_0/i_pointer ;
  wire   [3:0] \shifter_0/pointer ;
  wire   [19:0] \shifter_0/reg_w_15 ;
  wire   [19:0] \shifter_0/reg_w_14 ;
  wire   [19:0] \shifter_0/reg_w_13 ;
  wire   [19:0] \shifter_0/reg_w_12 ;
  wire   [19:0] \shifter_0/reg_w_11 ;
  wire   [19:0] \shifter_0/reg_w_10 ;
  wire   [19:0] \shifter_0/reg_w_9 ;
  wire   [19:0] \shifter_0/reg_w_8 ;
  wire   [19:0] \shifter_0/reg_w_7 ;
  wire   [19:0] \shifter_0/reg_w_6 ;
  wire   [19:0] \shifter_0/reg_w_5 ;
  wire   [19:0] \shifter_0/reg_w_4 ;
  wire   [19:0] \shifter_0/reg_w_3 ;
  wire   [19:0] \shifter_0/reg_w_2 ;
  wire   [19:0] \shifter_0/reg_w_1 ;
  wire   [19:0] \shifter_0/reg_w_0 ;
  wire   [19:0] \shifter_0/reg_i_15 ;
  wire   [19:0] \shifter_0/reg_i_14 ;
  wire   [19:0] \shifter_0/reg_i_13 ;
  wire   [19:0] \shifter_0/reg_i_12 ;
  wire   [19:0] \shifter_0/reg_i_11 ;
  wire   [19:0] \shifter_0/reg_i_10 ;
  wire   [19:0] \shifter_0/reg_i_9 ;
  wire   [19:0] \shifter_0/reg_i_8 ;
  wire   [19:0] \shifter_0/reg_i_7 ;
  wire   [19:0] \shifter_0/reg_i_6 ;
  wire   [19:0] \shifter_0/reg_i_5 ;
  wire   [19:0] \shifter_0/reg_i_4 ;
  wire   [19:0] \shifter_0/reg_i_3 ;
  wire   [19:0] \shifter_0/reg_i_2 ;
  wire   [19:0] \shifter_0/reg_i_1 ;
  wire   [19:0] \shifter_0/reg_i_0 ;

  dff_sg mask_input_ready_reg ( .D(input_ready), .CP(clk), .Q(mask_input_ready) );
  dff_sg delayed_input_ready_reg ( .D(n55071), .CP(clk), .Q(
        delayed_input_ready) );
  dff_sg filter_input_ready_reg ( .D(delayed_input_ready), .CP(clk), .Q(
        filter_input_ready) );
  dff_sg \state_reg[1]  ( .D(n45552), .CP(clk), .Q(n69264) );
  dff_sg \state_reg[0]  ( .D(n45553), .CP(clk), .Q(n69265) );
  dff_sg \reg_w_mask_reg[31]  ( .D(n10399), .CP(clk), .Q(reg_w_mask[31]) );
  dff_sg \reg_w_mask_reg[30]  ( .D(n10400), .CP(clk), .Q(reg_w_mask[30]) );
  dff_sg \reg_w_mask_reg[29]  ( .D(n10401), .CP(clk), .Q(reg_w_mask[29]) );
  dff_sg \reg_w_mask_reg[28]  ( .D(n10402), .CP(clk), .Q(reg_w_mask[28]) );
  dff_sg \reg_w_mask_reg[27]  ( .D(n10403), .CP(clk), .Q(reg_w_mask[27]) );
  dff_sg \reg_w_mask_reg[26]  ( .D(n10404), .CP(clk), .Q(reg_w_mask[26]) );
  dff_sg \reg_w_mask_reg[25]  ( .D(n10405), .CP(clk), .Q(reg_w_mask[25]) );
  dff_sg \reg_w_mask_reg[24]  ( .D(n10406), .CP(clk), .Q(reg_w_mask[24]) );
  dff_sg \reg_w_mask_reg[23]  ( .D(n10407), .CP(clk), .Q(reg_w_mask[23]) );
  dff_sg \reg_w_mask_reg[22]  ( .D(n10408), .CP(clk), .Q(reg_w_mask[22]) );
  dff_sg \reg_w_mask_reg[21]  ( .D(n10409), .CP(clk), .Q(reg_w_mask[21]) );
  dff_sg \reg_w_mask_reg[20]  ( .D(n10410), .CP(clk), .Q(reg_w_mask[20]) );
  dff_sg \reg_w_mask_reg[19]  ( .D(n10411), .CP(clk), .Q(reg_w_mask[19]) );
  dff_sg \reg_w_mask_reg[18]  ( .D(n10412), .CP(clk), .Q(reg_w_mask[18]) );
  dff_sg \reg_w_mask_reg[17]  ( .D(n10413), .CP(clk), .Q(reg_w_mask[17]) );
  dff_sg \reg_w_mask_reg[16]  ( .D(n10414), .CP(clk), .Q(reg_w_mask[16]) );
  dff_sg \reg_w_mask_reg[15]  ( .D(n10415), .CP(clk), .Q(reg_w_mask[15]) );
  dff_sg \reg_w_mask_reg[14]  ( .D(n10416), .CP(clk), .Q(reg_w_mask[14]) );
  dff_sg \reg_w_mask_reg[13]  ( .D(n10417), .CP(clk), .Q(reg_w_mask[13]) );
  dff_sg \reg_w_mask_reg[12]  ( .D(n10418), .CP(clk), .Q(reg_w_mask[12]) );
  dff_sg \reg_w_mask_reg[11]  ( .D(n10419), .CP(clk), .Q(reg_w_mask[11]) );
  dff_sg \reg_w_mask_reg[10]  ( .D(n10420), .CP(clk), .Q(reg_w_mask[10]) );
  dff_sg \reg_w_mask_reg[9]  ( .D(n10421), .CP(clk), .Q(reg_w_mask[9]) );
  dff_sg \reg_w_mask_reg[8]  ( .D(n10422), .CP(clk), .Q(reg_w_mask[8]) );
  dff_sg \reg_w_mask_reg[7]  ( .D(n10423), .CP(clk), .Q(reg_w_mask[7]) );
  dff_sg \reg_w_mask_reg[6]  ( .D(n10424), .CP(clk), .Q(reg_w_mask[6]) );
  dff_sg \reg_w_mask_reg[5]  ( .D(n10425), .CP(clk), .Q(reg_w_mask[5]) );
  dff_sg \reg_w_mask_reg[4]  ( .D(n10426), .CP(clk), .Q(reg_w_mask[4]) );
  dff_sg \reg_w_mask_reg[3]  ( .D(n10427), .CP(clk), .Q(reg_w_mask[3]) );
  dff_sg \reg_w_mask_reg[2]  ( .D(n10428), .CP(clk), .Q(reg_w_mask[2]) );
  dff_sg \reg_w_mask_reg[1]  ( .D(n10429), .CP(clk), .Q(reg_w_mask[1]) );
  dff_sg \reg_w_mask_reg[0]  ( .D(n10430), .CP(clk), .Q(reg_w_mask[0]) );
  dff_sg \reg_i_mask_reg[31]  ( .D(n10431), .CP(clk), .Q(reg_i_mask[31]) );
  dff_sg \reg_i_mask_reg[30]  ( .D(n10432), .CP(clk), .Q(reg_i_mask[30]) );
  dff_sg \reg_i_mask_reg[29]  ( .D(n10433), .CP(clk), .Q(reg_i_mask[29]) );
  dff_sg \reg_i_mask_reg[28]  ( .D(n10434), .CP(clk), .Q(reg_i_mask[28]) );
  dff_sg \reg_i_mask_reg[27]  ( .D(n10435), .CP(clk), .Q(reg_i_mask[27]) );
  dff_sg \reg_i_mask_reg[26]  ( .D(n10436), .CP(clk), .Q(reg_i_mask[26]) );
  dff_sg \reg_i_mask_reg[25]  ( .D(n10437), .CP(clk), .Q(reg_i_mask[25]) );
  dff_sg \reg_i_mask_reg[24]  ( .D(n10438), .CP(clk), .Q(reg_i_mask[24]) );
  dff_sg \reg_i_mask_reg[23]  ( .D(n10439), .CP(clk), .Q(reg_i_mask[23]) );
  dff_sg \reg_i_mask_reg[22]  ( .D(n10440), .CP(clk), .Q(reg_i_mask[22]) );
  dff_sg \reg_i_mask_reg[21]  ( .D(n10441), .CP(clk), .Q(reg_i_mask[21]) );
  dff_sg \reg_i_mask_reg[20]  ( .D(n10442), .CP(clk), .Q(reg_i_mask[20]) );
  dff_sg \reg_i_mask_reg[19]  ( .D(n10443), .CP(clk), .Q(reg_i_mask[19]) );
  dff_sg \reg_i_mask_reg[18]  ( .D(n10444), .CP(clk), .Q(reg_i_mask[18]) );
  dff_sg \reg_i_mask_reg[17]  ( .D(n10445), .CP(clk), .Q(reg_i_mask[17]) );
  dff_sg \reg_i_mask_reg[16]  ( .D(n10446), .CP(clk), .Q(reg_i_mask[16]) );
  dff_sg \reg_i_mask_reg[15]  ( .D(n10447), .CP(clk), .Q(reg_i_mask[15]) );
  dff_sg \reg_i_mask_reg[14]  ( .D(n10448), .CP(clk), .Q(reg_i_mask[14]) );
  dff_sg \reg_i_mask_reg[13]  ( .D(n10449), .CP(clk), .Q(reg_i_mask[13]) );
  dff_sg \reg_i_mask_reg[12]  ( .D(n10450), .CP(clk), .Q(reg_i_mask[12]) );
  dff_sg \reg_i_mask_reg[11]  ( .D(n10451), .CP(clk), .Q(reg_i_mask[11]) );
  dff_sg \reg_i_mask_reg[10]  ( .D(n10452), .CP(clk), .Q(reg_i_mask[10]) );
  dff_sg \reg_i_mask_reg[9]  ( .D(n10453), .CP(clk), .Q(reg_i_mask[9]) );
  dff_sg \reg_i_mask_reg[8]  ( .D(n10454), .CP(clk), .Q(reg_i_mask[8]) );
  dff_sg \reg_i_mask_reg[7]  ( .D(n10455), .CP(clk), .Q(reg_i_mask[7]) );
  dff_sg \reg_i_mask_reg[6]  ( .D(n10456), .CP(clk), .Q(reg_i_mask[6]) );
  dff_sg \reg_i_mask_reg[5]  ( .D(n10457), .CP(clk), .Q(reg_i_mask[5]) );
  dff_sg \reg_i_mask_reg[4]  ( .D(n10458), .CP(clk), .Q(reg_i_mask[4]) );
  dff_sg \reg_i_mask_reg[3]  ( .D(n10459), .CP(clk), .Q(reg_i_mask[3]) );
  dff_sg \reg_i_mask_reg[2]  ( .D(n10460), .CP(clk), .Q(reg_i_mask[2]) );
  dff_sg \reg_i_mask_reg[1]  ( .D(n10461), .CP(clk), .Q(reg_i_mask[1]) );
  dff_sg \reg_i_mask_reg[0]  ( .D(n10462), .CP(clk), .Q(reg_i_mask[0]) );
  dff_sg \reg_i_0_reg[0]  ( .D(n45712), .CP(clk), .Q(reg_i_0[0]) );
  dff_sg \reg_i_0_reg[1]  ( .D(n45711), .CP(clk), .Q(reg_i_0[1]) );
  dff_sg \reg_i_0_reg[2]  ( .D(n45837), .CP(clk), .Q(reg_i_0[2]) );
  dff_sg \reg_i_0_reg[3]  ( .D(n45836), .CP(clk), .Q(reg_i_0[3]) );
  dff_sg \reg_i_0_reg[4]  ( .D(n45840), .CP(clk), .Q(reg_i_0[4]) );
  dff_sg \reg_i_0_reg[5]  ( .D(n45839), .CP(clk), .Q(reg_i_0[5]) );
  dff_sg \reg_i_0_reg[6]  ( .D(n45831), .CP(clk), .Q(reg_i_0[6]) );
  dff_sg \reg_i_0_reg[7]  ( .D(n45830), .CP(clk), .Q(reg_i_0[7]) );
  dff_sg \reg_i_0_reg[8]  ( .D(n45834), .CP(clk), .Q(reg_i_0[8]) );
  dff_sg \reg_i_0_reg[9]  ( .D(n45833), .CP(clk), .Q(reg_i_0[9]) );
  dff_sg \reg_i_0_reg[10]  ( .D(n45844), .CP(clk), .Q(reg_i_0[10]) );
  dff_sg \reg_i_0_reg[11]  ( .D(n45843), .CP(clk), .Q(reg_i_0[11]) );
  dff_sg \reg_i_0_reg[12]  ( .D(n45847), .CP(clk), .Q(reg_i_0[12]) );
  dff_sg \reg_i_0_reg[13]  ( .D(n45846), .CP(clk), .Q(reg_i_0[13]) );
  dff_sg \reg_i_0_reg[14]  ( .D(n45845), .CP(clk), .Q(reg_i_0[14]) );
  dff_sg \reg_i_0_reg[15]  ( .D(n45842), .CP(clk), .Q(reg_i_0[15]) );
  dff_sg \reg_i_0_reg[16]  ( .D(n45841), .CP(clk), .Q(reg_i_0[16]) );
  dff_sg \reg_i_0_reg[17]  ( .D(n45832), .CP(clk), .Q(reg_i_0[17]) );
  dff_sg \reg_i_0_reg[18]  ( .D(n45821), .CP(clk), .Q(reg_i_0[18]) );
  dff_sg \reg_i_0_reg[19]  ( .D(n45820), .CP(clk), .Q(reg_i_0[19]) );
  dff_sg \reg_i_1_reg[0]  ( .D(n45801), .CP(clk), .Q(reg_i_1[0]) );
  dff_sg \reg_i_1_reg[1]  ( .D(n45819), .CP(clk), .Q(reg_i_1[1]) );
  dff_sg \reg_i_1_reg[2]  ( .D(n45803), .CP(clk), .Q(reg_i_1[2]) );
  dff_sg \reg_i_1_reg[3]  ( .D(n45802), .CP(clk), .Q(reg_i_1[3]) );
  dff_sg \reg_i_1_reg[4]  ( .D(n45806), .CP(clk), .Q(reg_i_1[4]) );
  dff_sg \reg_i_1_reg[5]  ( .D(n45805), .CP(clk), .Q(reg_i_1[5]) );
  dff_sg \reg_i_1_reg[6]  ( .D(n45822), .CP(clk), .Q(reg_i_1[6]) );
  dff_sg \reg_i_1_reg[7]  ( .D(n45826), .CP(clk), .Q(reg_i_1[7]) );
  dff_sg \reg_i_1_reg[8]  ( .D(n45823), .CP(clk), .Q(reg_i_1[8]) );
  dff_sg \reg_i_1_reg[9]  ( .D(n45829), .CP(clk), .Q(reg_i_1[9]) );
  dff_sg \reg_i_1_reg[10]  ( .D(n45825), .CP(clk), .Q(reg_i_1[10]) );
  dff_sg \reg_i_1_reg[11]  ( .D(n45824), .CP(clk), .Q(reg_i_1[11]) );
  dff_sg \reg_i_1_reg[12]  ( .D(n45828), .CP(clk), .Q(reg_i_1[12]) );
  dff_sg \reg_i_1_reg[13]  ( .D(n45827), .CP(clk), .Q(reg_i_1[13]) );
  dff_sg \reg_i_1_reg[14]  ( .D(n45874), .CP(clk), .Q(reg_i_1[14]) );
  dff_sg \reg_i_1_reg[15]  ( .D(n45873), .CP(clk), .Q(reg_i_1[15]) );
  dff_sg \reg_i_1_reg[16]  ( .D(n45877), .CP(clk), .Q(reg_i_1[16]) );
  dff_sg \reg_i_1_reg[17]  ( .D(n45876), .CP(clk), .Q(reg_i_1[17]) );
  dff_sg \reg_i_1_reg[18]  ( .D(n45868), .CP(clk), .Q(reg_i_1[18]) );
  dff_sg \reg_i_1_reg[19]  ( .D(n45867), .CP(clk), .Q(reg_i_1[19]) );
  dff_sg \reg_i_2_reg[0]  ( .D(n45871), .CP(clk), .Q(reg_i_2[0]) );
  dff_sg \reg_i_2_reg[1]  ( .D(n45870), .CP(clk), .Q(reg_i_2[1]) );
  dff_sg \reg_i_2_reg[2]  ( .D(n45879), .CP(clk), .Q(reg_i_2[2]) );
  dff_sg \reg_i_2_reg[3]  ( .D(n45878), .CP(clk), .Q(reg_i_2[3]) );
  dff_sg \reg_i_2_reg[4]  ( .D(n45708), .CP(clk), .Q(reg_i_2[4]) );
  dff_sg \reg_i_2_reg[5]  ( .D(n45707), .CP(clk), .Q(reg_i_2[5]) );
  dff_sg \reg_i_2_reg[6]  ( .D(n45869), .CP(clk), .Q(reg_i_2[6]) );
  dff_sg \reg_i_2_reg[7]  ( .D(n45866), .CP(clk), .Q(reg_i_2[7]) );
  dff_sg \reg_i_2_reg[8]  ( .D(n45859), .CP(clk), .Q(reg_i_2[8]) );
  dff_sg \reg_i_2_reg[9]  ( .D(n45880), .CP(clk), .Q(reg_i_2[9]) );
  dff_sg \reg_i_2_reg[10]  ( .D(n45856), .CP(clk), .Q(reg_i_2[10]) );
  dff_sg \reg_i_2_reg[11]  ( .D(n45848), .CP(clk), .Q(reg_i_2[11]) );
  dff_sg \reg_i_2_reg[12]  ( .D(n45858), .CP(clk), .Q(reg_i_2[12]) );
  dff_sg \reg_i_2_reg[13]  ( .D(n45857), .CP(clk), .Q(reg_i_2[13]) );
  dff_sg \reg_i_2_reg[14]  ( .D(n45850), .CP(clk), .Q(reg_i_2[14]) );
  dff_sg \reg_i_2_reg[15]  ( .D(n45849), .CP(clk), .Q(reg_i_2[15]) );
  dff_sg \reg_i_2_reg[16]  ( .D(n45852), .CP(clk), .Q(reg_i_2[16]) );
  dff_sg \reg_i_2_reg[17]  ( .D(n45851), .CP(clk), .Q(reg_i_2[17]) );
  dff_sg \reg_i_2_reg[18]  ( .D(n45855), .CP(clk), .Q(reg_i_2[18]) );
  dff_sg \reg_i_2_reg[19]  ( .D(n45854), .CP(clk), .Q(reg_i_2[19]) );
  dff_sg \reg_i_3_reg[0]  ( .D(n45860), .CP(clk), .Q(reg_i_3[0]) );
  dff_sg \reg_i_3_reg[1]  ( .D(n45853), .CP(clk), .Q(reg_i_3[1]) );
  dff_sg \reg_i_3_reg[2]  ( .D(n45862), .CP(clk), .Q(reg_i_3[2]) );
  dff_sg \reg_i_3_reg[3]  ( .D(n45861), .CP(clk), .Q(reg_i_3[3]) );
  dff_sg \reg_i_3_reg[4]  ( .D(n45865), .CP(clk), .Q(reg_i_3[4]) );
  dff_sg \reg_i_3_reg[5]  ( .D(n45864), .CP(clk), .Q(reg_i_3[5]) );
  dff_sg \reg_i_3_reg[6]  ( .D(n45752), .CP(clk), .Q(reg_i_3[6]) );
  dff_sg \reg_i_3_reg[7]  ( .D(n45751), .CP(clk), .Q(reg_i_3[7]) );
  dff_sg \reg_i_3_reg[8]  ( .D(n45755), .CP(clk), .Q(reg_i_3[8]) );
  dff_sg \reg_i_3_reg[9]  ( .D(n45754), .CP(clk), .Q(reg_i_3[9]) );
  dff_sg \reg_i_3_reg[10]  ( .D(n45746), .CP(clk), .Q(reg_i_3[10]) );
  dff_sg \reg_i_3_reg[11]  ( .D(n45745), .CP(clk), .Q(reg_i_3[11]) );
  dff_sg \reg_i_3_reg[12]  ( .D(n45749), .CP(clk), .Q(reg_i_3[12]) );
  dff_sg \reg_i_3_reg[13]  ( .D(n45748), .CP(clk), .Q(reg_i_3[13]) );
  dff_sg \reg_i_3_reg[14]  ( .D(n45764), .CP(clk), .Q(reg_i_3[14]) );
  dff_sg \reg_i_3_reg[15]  ( .D(n45763), .CP(clk), .Q(reg_i_3[15]) );
  dff_sg \reg_i_3_reg[16]  ( .D(n45767), .CP(clk), .Q(reg_i_3[16]) );
  dff_sg \reg_i_3_reg[17]  ( .D(n45766), .CP(clk), .Q(reg_i_3[17]) );
  dff_sg \reg_i_3_reg[18]  ( .D(n45758), .CP(clk), .Q(reg_i_3[18]) );
  dff_sg \reg_i_3_reg[19]  ( .D(n45757), .CP(clk), .Q(reg_i_3[19]) );
  dff_sg \reg_i_4_reg[0]  ( .D(n45761), .CP(clk), .Q(reg_i_4[0]) );
  dff_sg \reg_i_4_reg[1]  ( .D(n45760), .CP(clk), .Q(reg_i_4[1]) );
  dff_sg \reg_i_4_reg[2]  ( .D(n45728), .CP(clk), .Q(reg_i_4[2]) );
  dff_sg \reg_i_4_reg[3]  ( .D(n45727), .CP(clk), .Q(reg_i_4[3]) );
  dff_sg \reg_i_4_reg[4]  ( .D(n45731), .CP(clk), .Q(reg_i_4[4]) );
  dff_sg \reg_i_4_reg[5]  ( .D(n45730), .CP(clk), .Q(reg_i_4[5]) );
  dff_sg \reg_i_4_reg[6]  ( .D(n45722), .CP(clk), .Q(reg_i_4[6]) );
  dff_sg \reg_i_4_reg[7]  ( .D(n45721), .CP(clk), .Q(reg_i_4[7]) );
  dff_sg \reg_i_4_reg[8]  ( .D(n45725), .CP(clk), .Q(reg_i_4[8]) );
  dff_sg \reg_i_4_reg[9]  ( .D(n45724), .CP(clk), .Q(reg_i_4[9]) );
  dff_sg \reg_i_4_reg[10]  ( .D(n45740), .CP(clk), .Q(reg_i_4[10]) );
  dff_sg \reg_i_4_reg[11]  ( .D(n45739), .CP(clk), .Q(reg_i_4[11]) );
  dff_sg \reg_i_4_reg[12]  ( .D(n45743), .CP(clk), .Q(reg_i_4[12]) );
  dff_sg \reg_i_4_reg[13]  ( .D(n45742), .CP(clk), .Q(reg_i_4[13]) );
  dff_sg \reg_i_4_reg[14]  ( .D(n45734), .CP(clk), .Q(reg_i_4[14]) );
  dff_sg \reg_i_4_reg[15]  ( .D(n45733), .CP(clk), .Q(reg_i_4[15]) );
  dff_sg \reg_i_4_reg[16]  ( .D(n45737), .CP(clk), .Q(reg_i_4[16]) );
  dff_sg \reg_i_4_reg[17]  ( .D(n45736), .CP(clk), .Q(reg_i_4[17]) );
  dff_sg \reg_i_4_reg[18]  ( .D(n45790), .CP(clk), .Q(reg_i_4[18]) );
  dff_sg \reg_i_4_reg[19]  ( .D(n45789), .CP(clk), .Q(reg_i_4[19]) );
  dff_sg \reg_i_5_reg[0]  ( .D(n45793), .CP(clk), .Q(reg_i_5[0]) );
  dff_sg \reg_i_5_reg[1]  ( .D(n45792), .CP(clk), .Q(reg_i_5[1]) );
  dff_sg \reg_i_5_reg[2]  ( .D(n45778), .CP(clk), .Q(reg_i_5[2]) );
  dff_sg \reg_i_5_reg[3]  ( .D(n45787), .CP(clk), .Q(reg_i_5[3]) );
  dff_sg \reg_i_5_reg[4]  ( .D(n45775), .CP(clk), .Q(reg_i_5[4]) );
  dff_sg \reg_i_5_reg[5]  ( .D(n45781), .CP(clk), .Q(reg_i_5[5]) );
  dff_sg \reg_i_5_reg[6]  ( .D(n45795), .CP(clk), .Q(reg_i_5[6]) );
  dff_sg \reg_i_5_reg[7]  ( .D(n45794), .CP(clk), .Q(reg_i_5[7]) );
  dff_sg \reg_i_5_reg[8]  ( .D(n45788), .CP(clk), .Q(reg_i_5[8]) );
  dff_sg \reg_i_5_reg[9]  ( .D(n45798), .CP(clk), .Q(reg_i_5[9]) );
  dff_sg \reg_i_5_reg[10]  ( .D(n45797), .CP(clk), .Q(reg_i_5[10]) );
  dff_sg \reg_i_5_reg[11]  ( .D(n45796), .CP(clk), .Q(reg_i_5[11]) );
  dff_sg \reg_i_5_reg[12]  ( .D(n45800), .CP(clk), .Q(reg_i_5[12]) );
  dff_sg \reg_i_5_reg[13]  ( .D(n45799), .CP(clk), .Q(reg_i_5[13]) );
  dff_sg \reg_i_5_reg[14]  ( .D(n45769), .CP(clk), .Q(reg_i_5[14]) );
  dff_sg \reg_i_5_reg[15]  ( .D(n45768), .CP(clk), .Q(reg_i_5[15]) );
  dff_sg \reg_i_5_reg[16]  ( .D(n45772), .CP(clk), .Q(reg_i_5[16]) );
  dff_sg \reg_i_5_reg[17]  ( .D(n45710), .CP(clk), .Q(reg_i_5[17]) );
  dff_sg \reg_i_5_reg[18]  ( .D(n45771), .CP(clk), .Q(reg_i_5[18]) );
  dff_sg \reg_i_5_reg[19]  ( .D(n45770), .CP(clk), .Q(reg_i_5[19]) );
  dff_sg \reg_i_6_reg[0]  ( .D(n45774), .CP(clk), .Q(reg_i_6[0]) );
  dff_sg \reg_i_6_reg[1]  ( .D(n45773), .CP(clk), .Q(reg_i_6[1]) );
  dff_sg \reg_i_6_reg[2]  ( .D(n45783), .CP(clk), .Q(reg_i_6[2]) );
  dff_sg \reg_i_6_reg[3]  ( .D(n45782), .CP(clk), .Q(reg_i_6[3]) );
  dff_sg \reg_i_6_reg[4]  ( .D(n45786), .CP(clk), .Q(reg_i_6[4]) );
  dff_sg \reg_i_6_reg[5]  ( .D(n45785), .CP(clk), .Q(reg_i_6[5]) );
  dff_sg \reg_i_6_reg[6]  ( .D(n45777), .CP(clk), .Q(reg_i_6[6]) );
  dff_sg \reg_i_6_reg[7]  ( .D(n45776), .CP(clk), .Q(reg_i_6[7]) );
  dff_sg \reg_i_6_reg[8]  ( .D(n45780), .CP(clk), .Q(reg_i_6[8]) );
  dff_sg \reg_i_6_reg[9]  ( .D(n45779), .CP(clk), .Q(reg_i_6[9]) );
  dff_sg \reg_i_6_reg[10]  ( .D(n45573), .CP(clk), .Q(reg_i_6[10]) );
  dff_sg \reg_i_6_reg[11]  ( .D(n45572), .CP(clk), .Q(reg_i_6[11]) );
  dff_sg \reg_i_6_reg[12]  ( .D(n45744), .CP(clk), .Q(reg_i_6[12]) );
  dff_sg \reg_i_6_reg[13]  ( .D(n45741), .CP(clk), .Q(reg_i_6[13]) );
  dff_sg \reg_i_6_reg[14]  ( .D(n45987), .CP(clk), .Q(reg_i_6[14]) );
  dff_sg \reg_i_6_reg[15]  ( .D(n45720), .CP(clk), .Q(reg_i_6[15]) );
  dff_sg \reg_i_6_reg[16]  ( .D(n46143), .CP(clk), .Q(reg_i_6[16]) );
  dff_sg \reg_i_6_reg[17]  ( .D(n46155), .CP(clk), .Q(reg_i_6[17]) );
  dff_sg \reg_i_6_reg[18]  ( .D(n45732), .CP(clk), .Q(reg_i_6[18]) );
  dff_sg \reg_i_6_reg[19]  ( .D(n45729), .CP(clk), .Q(reg_i_6[19]) );
  dff_sg \reg_i_7_reg[0]  ( .D(n45726), .CP(clk), .Q(reg_i_7[0]) );
  dff_sg \reg_i_7_reg[1]  ( .D(n45723), .CP(clk), .Q(reg_i_7[1]) );
  dff_sg \reg_i_7_reg[2]  ( .D(n45568), .CP(clk), .Q(reg_i_7[2]) );
  dff_sg \reg_i_7_reg[3]  ( .D(n45574), .CP(clk), .Q(reg_i_7[3]) );
  dff_sg \reg_i_7_reg[4]  ( .D(n45738), .CP(clk), .Q(reg_i_7[4]) );
  dff_sg \reg_i_7_reg[5]  ( .D(n45735), .CP(clk), .Q(reg_i_7[5]) );
  dff_sg \reg_i_7_reg[6]  ( .D(n46089), .CP(clk), .Q(reg_i_7[6]) );
  dff_sg \reg_i_7_reg[7]  ( .D(n46059), .CP(clk), .Q(reg_i_7[7]) );
  dff_sg \reg_i_7_reg[8]  ( .D(n45984), .CP(clk), .Q(reg_i_7[8]) );
  dff_sg \reg_i_7_reg[9]  ( .D(n45969), .CP(clk), .Q(reg_i_7[9]) );
  dff_sg \reg_i_7_reg[10]  ( .D(n46131), .CP(clk), .Q(reg_i_7[10]) );
  dff_sg \reg_i_7_reg[11]  ( .D(n46128), .CP(clk), .Q(reg_i_7[11]) );
  dff_sg \reg_i_7_reg[12]  ( .D(n46122), .CP(clk), .Q(reg_i_7[12]) );
  dff_sg \reg_i_7_reg[13]  ( .D(n46113), .CP(clk), .Q(reg_i_7[13]) );
  dff_sg \reg_i_7_reg[14]  ( .D(n46152), .CP(clk), .Q(reg_i_7[14]) );
  dff_sg \reg_i_7_reg[15]  ( .D(n46149), .CP(clk), .Q(reg_i_7[15]) );
  dff_sg \reg_i_7_reg[16]  ( .D(n46140), .CP(clk), .Q(reg_i_7[16]) );
  dff_sg \reg_i_7_reg[17]  ( .D(n46137), .CP(clk), .Q(reg_i_7[17]) );
  dff_sg \reg_i_7_reg[18]  ( .D(n46179), .CP(clk), .Q(reg_i_7[18]) );
  dff_sg \reg_i_7_reg[19]  ( .D(n46176), .CP(clk), .Q(reg_i_7[19]) );
  dff_sg \reg_i_8_reg[0]  ( .D(n46173), .CP(clk), .Q(reg_i_8[0]) );
  dff_sg \reg_i_8_reg[1]  ( .D(n46170), .CP(clk), .Q(reg_i_8[1]) );
  dff_sg \reg_i_8_reg[2]  ( .D(n46116), .CP(clk), .Q(reg_i_8[2]) );
  dff_sg \reg_i_8_reg[3]  ( .D(n46083), .CP(clk), .Q(reg_i_8[3]) );
  dff_sg \reg_i_8_reg[4]  ( .D(n46080), .CP(clk), .Q(reg_i_8[4]) );
  dff_sg \reg_i_8_reg[5]  ( .D(n46077), .CP(clk), .Q(reg_i_8[5]) );
  dff_sg \reg_i_8_reg[6]  ( .D(n45807), .CP(clk), .Q(reg_i_8[6]) );
  dff_sg \reg_i_8_reg[7]  ( .D(n45906), .CP(clk), .Q(reg_i_8[7]) );
  dff_sg \reg_i_8_reg[8]  ( .D(n46119), .CP(clk), .Q(reg_i_8[8]) );
  dff_sg \reg_i_8_reg[9]  ( .D(n45554), .CP(clk), .Q(reg_i_8[9]) );
  dff_sg \reg_i_8_reg[10]  ( .D(n46020), .CP(clk), .Q(reg_i_8[10]) );
  dff_sg \reg_i_8_reg[11]  ( .D(n45963), .CP(clk), .Q(reg_i_8[11]) );
  dff_sg \reg_i_8_reg[12]  ( .D(n45586), .CP(clk), .Q(reg_i_8[12]) );
  dff_sg \reg_i_8_reg[13]  ( .D(n45585), .CP(clk), .Q(reg_i_8[13]) );
  dff_sg \reg_i_8_reg[14]  ( .D(n46074), .CP(clk), .Q(reg_i_8[14]) );
  dff_sg \reg_i_8_reg[15]  ( .D(n46035), .CP(clk), .Q(reg_i_8[15]) );
  dff_sg \reg_i_8_reg[16]  ( .D(n46029), .CP(clk), .Q(reg_i_8[16]) );
  dff_sg \reg_i_8_reg[17]  ( .D(n46026), .CP(clk), .Q(reg_i_8[17]) );
  dff_sg \reg_i_8_reg[18]  ( .D(n45756), .CP(clk), .Q(reg_i_8[18]) );
  dff_sg \reg_i_8_reg[19]  ( .D(n45753), .CP(clk), .Q(reg_i_8[19]) );
  dff_sg \reg_i_9_reg[0]  ( .D(n45750), .CP(clk), .Q(reg_i_9[0]) );
  dff_sg \reg_i_9_reg[1]  ( .D(n45747), .CP(clk), .Q(reg_i_9[1]) );
  dff_sg \reg_i_9_reg[2]  ( .D(n45784), .CP(clk), .Q(reg_i_9[2]) );
  dff_sg \reg_i_9_reg[3]  ( .D(n45875), .CP(clk), .Q(reg_i_9[3]) );
  dff_sg \reg_i_9_reg[4]  ( .D(n45762), .CP(clk), .Q(reg_i_9[4]) );
  dff_sg \reg_i_9_reg[5]  ( .D(n45759), .CP(clk), .Q(reg_i_9[5]) );
  dff_sg \reg_i_9_reg[6]  ( .D(n45894), .CP(clk), .Q(reg_i_9[6]) );
  dff_sg \reg_i_9_reg[7]  ( .D(n45810), .CP(clk), .Q(reg_i_9[7]) );
  dff_sg \reg_i_9_reg[8]  ( .D(n45765), .CP(clk), .Q(reg_i_9[8]) );
  dff_sg \reg_i_9_reg[9]  ( .D(n45581), .CP(clk), .Q(reg_i_9[9]) );
  dff_sg \reg_i_9_reg[10]  ( .D(n45960), .CP(clk), .Q(reg_i_9[10]) );
  dff_sg \reg_i_9_reg[11]  ( .D(n45957), .CP(clk), .Q(reg_i_9[11]) );
  dff_sg \reg_i_9_reg[12]  ( .D(n45954), .CP(clk), .Q(reg_i_9[12]) );
  dff_sg \reg_i_9_reg[13]  ( .D(n45909), .CP(clk), .Q(reg_i_9[13]) );
  dff_sg \reg_i_9_reg[14]  ( .D(n45885), .CP(clk), .Q(reg_i_9[14]) );
  dff_sg \reg_i_9_reg[15]  ( .D(n45897), .CP(clk), .Q(reg_i_9[15]) );
  dff_sg \reg_i_9_reg[16]  ( .D(n45816), .CP(clk), .Q(reg_i_9[16]) );
  dff_sg \reg_i_9_reg[17]  ( .D(n45882), .CP(clk), .Q(reg_i_9[17]) );
  dff_sg \reg_i_9_reg[18]  ( .D(n45891), .CP(clk), .Q(reg_i_9[18]) );
  dff_sg \reg_i_9_reg[19]  ( .D(n45888), .CP(clk), .Q(reg_i_9[19]) );
  dff_sg \reg_i_10_reg[0]  ( .D(n45881), .CP(clk), .Q(reg_i_10[0]) );
  dff_sg \reg_i_10_reg[1]  ( .D(n45654), .CP(clk), .Q(reg_i_10[1]) );
  dff_sg \reg_i_10_reg[2]  ( .D(n45936), .CP(clk), .Q(reg_i_10[2]) );
  dff_sg \reg_i_10_reg[3]  ( .D(n45927), .CP(clk), .Q(reg_i_10[3]) );
  dff_sg \reg_i_10_reg[4]  ( .D(n45930), .CP(clk), .Q(reg_i_10[4]) );
  dff_sg \reg_i_10_reg[5]  ( .D(n45918), .CP(clk), .Q(reg_i_10[5]) );
  dff_sg \reg_i_10_reg[6]  ( .D(n45933), .CP(clk), .Q(reg_i_10[6]) );
  dff_sg \reg_i_10_reg[7]  ( .D(n45555), .CP(clk), .Q(reg_i_10[7]) );
  dff_sg \reg_i_10_reg[8]  ( .D(n45924), .CP(clk), .Q(reg_i_10[8]) );
  dff_sg \reg_i_10_reg[9]  ( .D(n45921), .CP(clk), .Q(reg_i_10[9]) );
  dff_sg \reg_i_10_reg[10]  ( .D(n46158), .CP(clk), .Q(reg_i_10[10]) );
  dff_sg \reg_i_10_reg[11]  ( .D(n45558), .CP(clk), .Q(reg_i_10[11]) );
  dff_sg \reg_i_10_reg[12]  ( .D(n45675), .CP(clk), .Q(reg_i_10[12]) );
  dff_sg \reg_i_10_reg[13]  ( .D(n46164), .CP(clk), .Q(reg_i_10[13]) );
  dff_sg \reg_i_10_reg[14]  ( .D(n45556), .CP(clk), .Q(reg_i_10[14]) );
  dff_sg \reg_i_10_reg[15]  ( .D(n45557), .CP(clk), .Q(reg_i_10[15]) );
  dff_sg \reg_i_10_reg[16]  ( .D(n45672), .CP(clk), .Q(reg_i_10[16]) );
  dff_sg \reg_i_10_reg[17]  ( .D(n46167), .CP(clk), .Q(reg_i_10[17]) );
  dff_sg \reg_i_10_reg[18]  ( .D(n45915), .CP(clk), .Q(reg_i_10[18]) );
  dff_sg \reg_i_10_reg[19]  ( .D(n45560), .CP(clk), .Q(reg_i_10[19]) );
  dff_sg \reg_i_11_reg[0]  ( .D(n45912), .CP(clk), .Q(reg_i_11[0]) );
  dff_sg \reg_i_11_reg[1]  ( .D(n45903), .CP(clk), .Q(reg_i_11[1]) );
  dff_sg \reg_i_11_reg[2]  ( .D(n45900), .CP(clk), .Q(reg_i_11[2]) );
  dff_sg \reg_i_11_reg[3]  ( .D(n45559), .CP(clk), .Q(reg_i_11[3]) );
  dff_sg \reg_i_11_reg[4]  ( .D(n45813), .CP(clk), .Q(reg_i_11[4]) );
  dff_sg \reg_i_11_reg[5]  ( .D(n45561), .CP(clk), .Q(reg_i_11[5]) );
  dff_sg \reg_i_11_reg[6]  ( .D(n46056), .CP(clk), .Q(reg_i_11[6]) );
  dff_sg \reg_i_11_reg[7]  ( .D(n46101), .CP(clk), .Q(reg_i_11[7]) );
  dff_sg \reg_i_11_reg[8]  ( .D(n46107), .CP(clk), .Q(reg_i_11[8]) );
  dff_sg \reg_i_11_reg[9]  ( .D(n46104), .CP(clk), .Q(reg_i_11[9]) );
  dff_sg \reg_i_11_reg[10]  ( .D(n46014), .CP(clk), .Q(reg_i_11[10]) );
  dff_sg \reg_i_11_reg[11]  ( .D(n45575), .CP(clk), .Q(reg_i_11[11]) );
  dff_sg \reg_i_11_reg[12]  ( .D(n46053), .CP(clk), .Q(reg_i_11[12]) );
  dff_sg \reg_i_11_reg[13]  ( .D(n46017), .CP(clk), .Q(reg_i_11[13]) );
  dff_sg \reg_i_11_reg[14]  ( .D(n46086), .CP(clk), .Q(reg_i_11[14]) );
  dff_sg \reg_i_11_reg[15]  ( .D(n46098), .CP(clk), .Q(reg_i_11[15]) );
  dff_sg \reg_i_11_reg[16]  ( .D(n46062), .CP(clk), .Q(reg_i_11[16]) );
  dff_sg \reg_i_11_reg[17]  ( .D(n46071), .CP(clk), .Q(reg_i_11[17]) );
  dff_sg \reg_i_11_reg[18]  ( .D(n46095), .CP(clk), .Q(reg_i_11[18]) );
  dff_sg \reg_i_11_reg[19]  ( .D(n46092), .CP(clk), .Q(reg_i_11[19]) );
  dff_sg \reg_i_12_reg[0]  ( .D(n46068), .CP(clk), .Q(reg_i_12[0]) );
  dff_sg \reg_i_12_reg[1]  ( .D(n46065), .CP(clk), .Q(reg_i_12[1]) );
  dff_sg \reg_i_12_reg[2]  ( .D(n45990), .CP(clk), .Q(reg_i_12[2]) );
  dff_sg \reg_i_12_reg[3]  ( .D(n45564), .CP(clk), .Q(reg_i_12[3]) );
  dff_sg \reg_i_12_reg[4]  ( .D(n45972), .CP(clk), .Q(reg_i_12[4]) );
  dff_sg \reg_i_12_reg[5]  ( .D(n45993), .CP(clk), .Q(reg_i_12[5]) );
  dff_sg \reg_i_12_reg[6]  ( .D(n45562), .CP(clk), .Q(reg_i_12[6]) );
  dff_sg \reg_i_12_reg[7]  ( .D(n45563), .CP(clk), .Q(reg_i_12[7]) );
  dff_sg \reg_i_12_reg[8]  ( .D(n45999), .CP(clk), .Q(reg_i_12[8]) );
  dff_sg \reg_i_12_reg[9]  ( .D(n45996), .CP(clk), .Q(reg_i_12[9]) );
  dff_sg \reg_i_12_reg[10]  ( .D(n45565), .CP(clk), .Q(reg_i_12[10]) );
  dff_sg \reg_i_12_reg[11]  ( .D(n45566), .CP(clk), .Q(reg_i_12[11]) );
  dff_sg \reg_i_12_reg[12]  ( .D(n46050), .CP(clk), .Q(reg_i_12[12]) );
  dff_sg \reg_i_12_reg[13]  ( .D(n46032), .CP(clk), .Q(reg_i_12[13]) );
  dff_sg \reg_i_12_reg[14]  ( .D(n46002), .CP(clk), .Q(reg_i_12[14]) );
  dff_sg \reg_i_12_reg[15]  ( .D(n45567), .CP(clk), .Q(reg_i_12[15]) );
  dff_sg \reg_i_12_reg[16]  ( .D(n46005), .CP(clk), .Q(reg_i_12[16]) );
  dff_sg \reg_i_12_reg[17]  ( .D(n45939), .CP(clk), .Q(reg_i_12[17]) );
  dff_sg \reg_i_12_reg[18]  ( .D(n45659), .CP(clk), .Q(reg_i_12[18]) );
  dff_sg \reg_i_12_reg[19]  ( .D(n45658), .CP(clk), .Q(reg_i_12[19]) );
  dff_sg \reg_i_13_reg[0]  ( .D(n45651), .CP(clk), .Q(reg_i_13[0]) );
  dff_sg \reg_i_13_reg[1]  ( .D(n45657), .CP(clk), .Q(reg_i_13[1]) );
  dff_sg \reg_i_13_reg[2]  ( .D(n45653), .CP(clk), .Q(reg_i_13[2]) );
  dff_sg \reg_i_13_reg[3]  ( .D(n45652), .CP(clk), .Q(reg_i_13[3]) );
  dff_sg \reg_i_13_reg[4]  ( .D(n45656), .CP(clk), .Q(reg_i_13[4]) );
  dff_sg \reg_i_13_reg[5]  ( .D(n45655), .CP(clk), .Q(reg_i_13[5]) );
  dff_sg \reg_i_13_reg[6]  ( .D(n45680), .CP(clk), .Q(reg_i_13[6]) );
  dff_sg \reg_i_13_reg[7]  ( .D(n45679), .CP(clk), .Q(reg_i_13[7]) );
  dff_sg \reg_i_13_reg[8]  ( .D(n45660), .CP(clk), .Q(reg_i_13[8]) );
  dff_sg \reg_i_13_reg[9]  ( .D(n45678), .CP(clk), .Q(reg_i_13[9]) );
  dff_sg \reg_i_13_reg[10]  ( .D(n45662), .CP(clk), .Q(reg_i_13[10]) );
  dff_sg \reg_i_13_reg[11]  ( .D(n45661), .CP(clk), .Q(reg_i_13[11]) );
  dff_sg \reg_i_13_reg[12]  ( .D(n45665), .CP(clk), .Q(reg_i_13[12]) );
  dff_sg \reg_i_13_reg[13]  ( .D(n45664), .CP(clk), .Q(reg_i_13[13]) );
  dff_sg \reg_i_13_reg[14]  ( .D(n45640), .CP(clk), .Q(reg_i_13[14]) );
  dff_sg \reg_i_13_reg[15]  ( .D(n45639), .CP(clk), .Q(reg_i_13[15]) );
  dff_sg \reg_i_13_reg[16]  ( .D(n45643), .CP(clk), .Q(reg_i_13[16]) );
  dff_sg \reg_i_13_reg[17]  ( .D(n45642), .CP(clk), .Q(reg_i_13[17]) );
  dff_sg \reg_i_13_reg[18]  ( .D(n45634), .CP(clk), .Q(reg_i_13[18]) );
  dff_sg \reg_i_13_reg[19]  ( .D(n45633), .CP(clk), .Q(reg_i_13[19]) );
  dff_sg \reg_i_14_reg[0]  ( .D(n45637), .CP(clk), .Q(reg_i_14[0]) );
  dff_sg \reg_i_14_reg[1]  ( .D(n45636), .CP(clk), .Q(reg_i_14[1]) );
  dff_sg \reg_i_14_reg[2]  ( .D(n45647), .CP(clk), .Q(reg_i_14[2]) );
  dff_sg \reg_i_14_reg[3]  ( .D(n45646), .CP(clk), .Q(reg_i_14[3]) );
  dff_sg \reg_i_14_reg[4]  ( .D(n45650), .CP(clk), .Q(reg_i_14[4]) );
  dff_sg \reg_i_14_reg[5]  ( .D(n45649), .CP(clk), .Q(reg_i_14[5]) );
  dff_sg \reg_i_14_reg[6]  ( .D(n45648), .CP(clk), .Q(reg_i_14[6]) );
  dff_sg \reg_i_14_reg[7]  ( .D(n45645), .CP(clk), .Q(reg_i_14[7]) );
  dff_sg \reg_i_14_reg[8]  ( .D(n45638), .CP(clk), .Q(reg_i_14[8]) );
  dff_sg \reg_i_14_reg[9]  ( .D(n45644), .CP(clk), .Q(reg_i_14[9]) );
  dff_sg \reg_i_14_reg[10]  ( .D(n45694), .CP(clk), .Q(reg_i_14[10]) );
  dff_sg \reg_i_14_reg[11]  ( .D(n45701), .CP(clk), .Q(reg_i_14[11]) );
  dff_sg \reg_i_14_reg[12]  ( .D(n45703), .CP(clk), .Q(reg_i_14[12]) );
  dff_sg \reg_i_14_reg[13]  ( .D(n45702), .CP(clk), .Q(reg_i_14[13]) );
  dff_sg \reg_i_14_reg[14]  ( .D(n45706), .CP(clk), .Q(reg_i_14[14]) );
  dff_sg \reg_i_14_reg[15]  ( .D(n45705), .CP(clk), .Q(reg_i_14[15]) );
  dff_sg \reg_i_14_reg[16]  ( .D(n45697), .CP(clk), .Q(reg_i_14[16]) );
  dff_sg \reg_i_14_reg[17]  ( .D(n45704), .CP(clk), .Q(reg_i_14[17]) );
  dff_sg \reg_i_14_reg[18]  ( .D(n45569), .CP(clk), .Q(reg_i_14[18]) );
  dff_sg \reg_i_14_reg[19]  ( .D(n45709), .CP(clk), .Q(reg_i_14[19]) );
  dff_sg \reg_i_15_reg[0]  ( .D(n45700), .CP(clk), .Q(reg_i_15[0]) );
  dff_sg \reg_i_15_reg[1]  ( .D(n45641), .CP(clk), .Q(reg_i_15[1]) );
  dff_sg \reg_i_15_reg[2]  ( .D(n45571), .CP(clk), .Q(reg_i_15[2]) );
  dff_sg \reg_i_15_reg[3]  ( .D(n45570), .CP(clk), .Q(reg_i_15[3]) );
  dff_sg \reg_i_15_reg[4]  ( .D(n45591), .CP(clk), .Q(reg_i_15[4]) );
  dff_sg \reg_i_15_reg[5]  ( .D(n45608), .CP(clk), .Q(reg_i_15[5]) );
  dff_sg \reg_i_15_reg[6]  ( .D(n45689), .CP(clk), .Q(reg_i_15[6]) );
  dff_sg \reg_i_15_reg[7]  ( .D(n45688), .CP(clk), .Q(reg_i_15[7]) );
  dff_sg \reg_i_15_reg[8]  ( .D(n45692), .CP(clk), .Q(reg_i_15[8]) );
  dff_sg \reg_i_15_reg[9]  ( .D(n45691), .CP(clk), .Q(reg_i_15[9]) );
  dff_sg \reg_i_15_reg[10]  ( .D(n45683), .CP(clk), .Q(reg_i_15[10]) );
  dff_sg \reg_i_15_reg[11]  ( .D(n45682), .CP(clk), .Q(reg_i_15[11]) );
  dff_sg \reg_i_15_reg[12]  ( .D(n45686), .CP(clk), .Q(reg_i_15[12]) );
  dff_sg \reg_i_15_reg[13]  ( .D(n45685), .CP(clk), .Q(reg_i_15[13]) );
  dff_sg \reg_i_15_reg[14]  ( .D(n45696), .CP(clk), .Q(reg_i_15[14]) );
  dff_sg \reg_i_15_reg[15]  ( .D(n45695), .CP(clk), .Q(reg_i_15[15]) );
  dff_sg \reg_i_15_reg[16]  ( .D(n45699), .CP(clk), .Q(reg_i_15[16]) );
  dff_sg \reg_i_15_reg[17]  ( .D(n45698), .CP(clk), .Q(reg_i_15[17]) );
  dff_sg \reg_i_15_reg[18]  ( .D(n45687), .CP(clk), .Q(reg_i_15[18]) );
  dff_sg \reg_i_15_reg[19]  ( .D(n45684), .CP(clk), .Q(reg_i_15[19]) );
  dff_sg \reg_w_0_reg[0]  ( .D(n45681), .CP(clk), .Q(reg_w_0[0]) );
  dff_sg \reg_w_0_reg[1]  ( .D(n45693), .CP(clk), .Q(reg_w_0[1]) );
  dff_sg \reg_w_0_reg[2]  ( .D(n45596), .CP(clk), .Q(reg_w_0[2]) );
  dff_sg \reg_w_0_reg[3]  ( .D(n45595), .CP(clk), .Q(reg_w_0[3]) );
  dff_sg \reg_w_0_reg[4]  ( .D(n46023), .CP(clk), .Q(reg_w_0[4]) );
  dff_sg \reg_w_0_reg[5]  ( .D(n45594), .CP(clk), .Q(reg_w_0[5]) );
  dff_sg \reg_w_0_reg[6]  ( .D(n45590), .CP(clk), .Q(reg_w_0[6]) );
  dff_sg \reg_w_0_reg[7]  ( .D(n45589), .CP(clk), .Q(reg_w_0[7]) );
  dff_sg \reg_w_0_reg[8]  ( .D(n45593), .CP(clk), .Q(reg_w_0[8]) );
  dff_sg \reg_w_0_reg[9]  ( .D(n45592), .CP(clk), .Q(reg_w_0[9]) );
  dff_sg \reg_w_0_reg[10]  ( .D(n45600), .CP(clk), .Q(reg_w_0[10]) );
  dff_sg \reg_w_0_reg[11]  ( .D(n45599), .CP(clk), .Q(reg_w_0[11]) );
  dff_sg \reg_w_0_reg[12]  ( .D(n45603), .CP(clk), .Q(reg_w_0[12]) );
  dff_sg \reg_w_0_reg[13]  ( .D(n45602), .CP(clk), .Q(reg_w_0[13]) );
  dff_sg \reg_w_0_reg[14]  ( .D(n45588), .CP(clk), .Q(reg_w_0[14]) );
  dff_sg \reg_w_0_reg[15]  ( .D(n45582), .CP(clk), .Q(reg_w_0[15]) );
  dff_sg \reg_w_0_reg[16]  ( .D(n45584), .CP(clk), .Q(reg_w_0[16]) );
  dff_sg \reg_w_0_reg[17]  ( .D(n45583), .CP(clk), .Q(reg_w_0[17]) );
  dff_sg \reg_w_0_reg[18]  ( .D(n45578), .CP(clk), .Q(reg_w_0[18]) );
  dff_sg \reg_w_0_reg[19]  ( .D(n45577), .CP(clk), .Q(reg_w_0[19]) );
  dff_sg \reg_w_1_reg[0]  ( .D(n46011), .CP(clk), .Q(reg_w_1[0]) );
  dff_sg \reg_w_1_reg[1]  ( .D(n45580), .CP(clk), .Q(reg_w_1[1]) );
  dff_sg \reg_w_1_reg[2]  ( .D(n45576), .CP(clk), .Q(reg_w_1[2]) );
  dff_sg \reg_w_1_reg[3]  ( .D(n46134), .CP(clk), .Q(reg_w_1[3]) );
  dff_sg \reg_w_1_reg[4]  ( .D(n45579), .CP(clk), .Q(reg_w_1[4]) );
  dff_sg \reg_w_1_reg[5]  ( .D(n45587), .CP(clk), .Q(reg_w_1[5]) );
  dff_sg \reg_w_1_reg[6]  ( .D(n46008), .CP(clk), .Q(reg_w_1[6]) );
  dff_sg \reg_w_1_reg[7]  ( .D(n46188), .CP(clk), .Q(reg_w_1[7]) );
  dff_sg \reg_w_1_reg[8]  ( .D(n46191), .CP(clk), .Q(reg_w_1[8]) );
  dff_sg \reg_w_1_reg[9]  ( .D(n46146), .CP(clk), .Q(reg_w_1[9]) );
  dff_sg \reg_w_1_reg[10]  ( .D(n45975), .CP(clk), .Q(reg_w_1[10]) );
  dff_sg \reg_w_1_reg[11]  ( .D(n45966), .CP(clk), .Q(reg_w_1[11]) );
  dff_sg \reg_w_1_reg[12]  ( .D(n46185), .CP(clk), .Q(reg_w_1[12]) );
  dff_sg \reg_w_1_reg[13]  ( .D(n46182), .CP(clk), .Q(reg_w_1[13]) );
  dff_sg \reg_w_1_reg[14]  ( .D(n45618), .CP(clk), .Q(reg_w_1[14]) );
  dff_sg \reg_w_1_reg[15]  ( .D(n45622), .CP(clk), .Q(reg_w_1[15]) );
  dff_sg \reg_w_1_reg[16]  ( .D(n45619), .CP(clk), .Q(reg_w_1[16]) );
  dff_sg \reg_w_1_reg[17]  ( .D(n45629), .CP(clk), .Q(reg_w_1[17]) );
  dff_sg \reg_w_1_reg[18]  ( .D(n45621), .CP(clk), .Q(reg_w_1[18]) );
  dff_sg \reg_w_1_reg[19]  ( .D(n45620), .CP(clk), .Q(reg_w_1[19]) );
  dff_sg \reg_w_2_reg[0]  ( .D(n45624), .CP(clk), .Q(reg_w_2[0]) );
  dff_sg \reg_w_2_reg[1]  ( .D(n45623), .CP(clk), .Q(reg_w_2[1]) );
  dff_sg \reg_w_2_reg[2]  ( .D(n45625), .CP(clk), .Q(reg_w_2[2]) );
  dff_sg \reg_w_2_reg[3]  ( .D(n45626), .CP(clk), .Q(reg_w_2[3]) );
  dff_sg \reg_w_2_reg[4]  ( .D(n45632), .CP(clk), .Q(reg_w_2[4]) );
  dff_sg \reg_w_2_reg[5]  ( .D(n45635), .CP(clk), .Q(reg_w_2[5]) );
  dff_sg \reg_w_2_reg[6]  ( .D(n45628), .CP(clk), .Q(reg_w_2[6]) );
  dff_sg \reg_w_2_reg[7]  ( .D(n45627), .CP(clk), .Q(reg_w_2[7]) );
  dff_sg \reg_w_2_reg[8]  ( .D(n45631), .CP(clk), .Q(reg_w_2[8]) );
  dff_sg \reg_w_2_reg[9]  ( .D(n45630), .CP(clk), .Q(reg_w_2[9]) );
  dff_sg \reg_w_2_reg[10]  ( .D(n45607), .CP(clk), .Q(reg_w_2[10]) );
  dff_sg \reg_w_2_reg[11]  ( .D(n45606), .CP(clk), .Q(reg_w_2[11]) );
  dff_sg \reg_w_2_reg[12]  ( .D(n45610), .CP(clk), .Q(reg_w_2[12]) );
  dff_sg \reg_w_2_reg[13]  ( .D(n45609), .CP(clk), .Q(reg_w_2[13]) );
  dff_sg \reg_w_2_reg[14]  ( .D(n45597), .CP(clk), .Q(reg_w_2[14]) );
  dff_sg \reg_w_2_reg[15]  ( .D(n45604), .CP(clk), .Q(reg_w_2[15]) );
  dff_sg \reg_w_2_reg[16]  ( .D(n45601), .CP(clk), .Q(reg_w_2[16]) );
  dff_sg \reg_w_2_reg[17]  ( .D(n45598), .CP(clk), .Q(reg_w_2[17]) );
  dff_sg \reg_w_2_reg[18]  ( .D(n45612), .CP(clk), .Q(reg_w_2[18]) );
  dff_sg \reg_w_2_reg[19]  ( .D(n45611), .CP(clk), .Q(reg_w_2[19]) );
  dff_sg \reg_w_3_reg[0]  ( .D(n45605), .CP(clk), .Q(reg_w_3[0]) );
  dff_sg \reg_w_3_reg[1]  ( .D(n45615), .CP(clk), .Q(reg_w_3[1]) );
  dff_sg \reg_w_3_reg[2]  ( .D(n45614), .CP(clk), .Q(reg_w_3[2]) );
  dff_sg \reg_w_3_reg[3]  ( .D(n45613), .CP(clk), .Q(reg_w_3[3]) );
  dff_sg \reg_w_3_reg[4]  ( .D(n45617), .CP(clk), .Q(reg_w_3[4]) );
  dff_sg \reg_w_3_reg[5]  ( .D(n45616), .CP(clk), .Q(reg_w_3[5]) );
  dff_sg \reg_w_3_reg[6]  ( .D(n45974), .CP(clk), .Q(reg_w_3[6]) );
  dff_sg \reg_w_3_reg[7]  ( .D(n45973), .CP(clk), .Q(reg_w_3[7]) );
  dff_sg \reg_w_3_reg[8]  ( .D(n45977), .CP(clk), .Q(reg_w_3[8]) );
  dff_sg \reg_w_3_reg[9]  ( .D(n45976), .CP(clk), .Q(reg_w_3[9]) );
  dff_sg \reg_w_3_reg[10]  ( .D(n45968), .CP(clk), .Q(reg_w_3[10]) );
  dff_sg \reg_w_3_reg[11]  ( .D(n45967), .CP(clk), .Q(reg_w_3[11]) );
  dff_sg \reg_w_3_reg[12]  ( .D(n45971), .CP(clk), .Q(reg_w_3[12]) );
  dff_sg \reg_w_3_reg[13]  ( .D(n45970), .CP(clk), .Q(reg_w_3[13]) );
  dff_sg \reg_w_3_reg[14]  ( .D(n45986), .CP(clk), .Q(reg_w_3[14]) );
  dff_sg \reg_w_3_reg[15]  ( .D(n45985), .CP(clk), .Q(reg_w_3[15]) );
  dff_sg \reg_w_3_reg[16]  ( .D(n45989), .CP(clk), .Q(reg_w_3[16]) );
  dff_sg \reg_w_3_reg[17]  ( .D(n45988), .CP(clk), .Q(reg_w_3[17]) );
  dff_sg \reg_w_3_reg[18]  ( .D(n45980), .CP(clk), .Q(reg_w_3[18]) );
  dff_sg \reg_w_3_reg[19]  ( .D(n45979), .CP(clk), .Q(reg_w_3[19]) );
  dff_sg \reg_w_4_reg[0]  ( .D(n45983), .CP(clk), .Q(reg_w_4[0]) );
  dff_sg \reg_w_4_reg[1]  ( .D(n45982), .CP(clk), .Q(reg_w_4[1]) );
  dff_sg \reg_w_4_reg[2]  ( .D(n45950), .CP(clk), .Q(reg_w_4[2]) );
  dff_sg \reg_w_4_reg[3]  ( .D(n45949), .CP(clk), .Q(reg_w_4[3]) );
  dff_sg \reg_w_4_reg[4]  ( .D(n45953), .CP(clk), .Q(reg_w_4[4]) );
  dff_sg \reg_w_4_reg[5]  ( .D(n45952), .CP(clk), .Q(reg_w_4[5]) );
  dff_sg \reg_w_4_reg[6]  ( .D(n45944), .CP(clk), .Q(reg_w_4[6]) );
  dff_sg \reg_w_4_reg[7]  ( .D(n45943), .CP(clk), .Q(reg_w_4[7]) );
  dff_sg \reg_w_4_reg[8]  ( .D(n45947), .CP(clk), .Q(reg_w_4[8]) );
  dff_sg \reg_w_4_reg[9]  ( .D(n45946), .CP(clk), .Q(reg_w_4[9]) );
  dff_sg \reg_w_4_reg[10]  ( .D(n45962), .CP(clk), .Q(reg_w_4[10]) );
  dff_sg \reg_w_4_reg[11]  ( .D(n45961), .CP(clk), .Q(reg_w_4[11]) );
  dff_sg \reg_w_4_reg[12]  ( .D(n45965), .CP(clk), .Q(reg_w_4[12]) );
  dff_sg \reg_w_4_reg[13]  ( .D(n45964), .CP(clk), .Q(reg_w_4[13]) );
  dff_sg \reg_w_4_reg[14]  ( .D(n45956), .CP(clk), .Q(reg_w_4[14]) );
  dff_sg \reg_w_4_reg[15]  ( .D(n45955), .CP(clk), .Q(reg_w_4[15]) );
  dff_sg \reg_w_4_reg[16]  ( .D(n45959), .CP(clk), .Q(reg_w_4[16]) );
  dff_sg \reg_w_4_reg[17]  ( .D(n45958), .CP(clk), .Q(reg_w_4[17]) );
  dff_sg \reg_w_4_reg[18]  ( .D(n46022), .CP(clk), .Q(reg_w_4[18]) );
  dff_sg \reg_w_4_reg[19]  ( .D(n46021), .CP(clk), .Q(reg_w_4[19]) );
  dff_sg \reg_w_5_reg[0]  ( .D(n46025), .CP(clk), .Q(reg_w_5[0]) );
  dff_sg \reg_w_5_reg[1]  ( .D(n46024), .CP(clk), .Q(reg_w_5[1]) );
  dff_sg \reg_w_5_reg[2]  ( .D(n46016), .CP(clk), .Q(reg_w_5[2]) );
  dff_sg \reg_w_5_reg[3]  ( .D(n46015), .CP(clk), .Q(reg_w_5[3]) );
  dff_sg \reg_w_5_reg[4]  ( .D(n46019), .CP(clk), .Q(reg_w_5[4]) );
  dff_sg \reg_w_5_reg[5]  ( .D(n46018), .CP(clk), .Q(reg_w_5[5]) );
  dff_sg \reg_w_5_reg[6]  ( .D(n46034), .CP(clk), .Q(reg_w_5[6]) );
  dff_sg \reg_w_5_reg[7]  ( .D(n46033), .CP(clk), .Q(reg_w_5[7]) );
  dff_sg \reg_w_5_reg[8]  ( .D(n46037), .CP(clk), .Q(reg_w_5[8]) );
  dff_sg \reg_w_5_reg[9]  ( .D(n46036), .CP(clk), .Q(reg_w_5[9]) );
  dff_sg \reg_w_5_reg[10]  ( .D(n46028), .CP(clk), .Q(reg_w_5[10]) );
  dff_sg \reg_w_5_reg[11]  ( .D(n46027), .CP(clk), .Q(reg_w_5[11]) );
  dff_sg \reg_w_5_reg[12]  ( .D(n46031), .CP(clk), .Q(reg_w_5[12]) );
  dff_sg \reg_w_5_reg[13]  ( .D(n46030), .CP(clk), .Q(reg_w_5[13]) );
  dff_sg \reg_w_5_reg[14]  ( .D(n45998), .CP(clk), .Q(reg_w_5[14]) );
  dff_sg \reg_w_5_reg[15]  ( .D(n45997), .CP(clk), .Q(reg_w_5[15]) );
  dff_sg \reg_w_5_reg[16]  ( .D(n46001), .CP(clk), .Q(reg_w_5[16]) );
  dff_sg \reg_w_5_reg[17]  ( .D(n46000), .CP(clk), .Q(reg_w_5[17]) );
  dff_sg \reg_w_5_reg[18]  ( .D(n45992), .CP(clk), .Q(reg_w_5[18]) );
  dff_sg \reg_w_5_reg[19]  ( .D(n45991), .CP(clk), .Q(reg_w_5[19]) );
  dff_sg \reg_w_6_reg[0]  ( .D(n45995), .CP(clk), .Q(reg_w_6[0]) );
  dff_sg \reg_w_6_reg[1]  ( .D(n45994), .CP(clk), .Q(reg_w_6[1]) );
  dff_sg \reg_w_6_reg[2]  ( .D(n46010), .CP(clk), .Q(reg_w_6[2]) );
  dff_sg \reg_w_6_reg[3]  ( .D(n46009), .CP(clk), .Q(reg_w_6[3]) );
  dff_sg \reg_w_6_reg[4]  ( .D(n46013), .CP(clk), .Q(reg_w_6[4]) );
  dff_sg \reg_w_6_reg[5]  ( .D(n46012), .CP(clk), .Q(reg_w_6[5]) );
  dff_sg \reg_w_6_reg[6]  ( .D(n46004), .CP(clk), .Q(reg_w_6[6]) );
  dff_sg \reg_w_6_reg[7]  ( .D(n46003), .CP(clk), .Q(reg_w_6[7]) );
  dff_sg \reg_w_6_reg[8]  ( .D(n46007), .CP(clk), .Q(reg_w_6[8]) );
  dff_sg \reg_w_6_reg[9]  ( .D(n46006), .CP(clk), .Q(reg_w_6[9]) );
  dff_sg \reg_w_6_reg[10]  ( .D(n45809), .CP(clk), .Q(reg_w_6[10]) );
  dff_sg \reg_w_6_reg[11]  ( .D(n45808), .CP(clk), .Q(reg_w_6[11]) );
  dff_sg \reg_w_6_reg[12]  ( .D(n45812), .CP(clk), .Q(reg_w_6[12]) );
  dff_sg \reg_w_6_reg[13]  ( .D(n45811), .CP(clk), .Q(reg_w_6[13]) );
  dff_sg \reg_w_6_reg[14]  ( .D(n45838), .CP(clk), .Q(reg_w_6[14]) );
  dff_sg \reg_w_6_reg[15]  ( .D(n45872), .CP(clk), .Q(reg_w_6[15]) );
  dff_sg \reg_w_6_reg[16]  ( .D(n45835), .CP(clk), .Q(reg_w_6[16]) );
  dff_sg \reg_w_6_reg[17]  ( .D(n45804), .CP(clk), .Q(reg_w_6[17]) );
  dff_sg \reg_w_6_reg[18]  ( .D(n45890), .CP(clk), .Q(reg_w_6[18]) );
  dff_sg \reg_w_6_reg[19]  ( .D(n45889), .CP(clk), .Q(reg_w_6[19]) );
  dff_sg \reg_w_7_reg[0]  ( .D(n45893), .CP(clk), .Q(reg_w_7[0]) );
  dff_sg \reg_w_7_reg[1]  ( .D(n45892), .CP(clk), .Q(reg_w_7[1]) );
  dff_sg \reg_w_7_reg[2]  ( .D(n45884), .CP(clk), .Q(reg_w_7[2]) );
  dff_sg \reg_w_7_reg[3]  ( .D(n45883), .CP(clk), .Q(reg_w_7[3]) );
  dff_sg \reg_w_7_reg[4]  ( .D(n45887), .CP(clk), .Q(reg_w_7[4]) );
  dff_sg \reg_w_7_reg[5]  ( .D(n45886), .CP(clk), .Q(reg_w_7[5]) );
  dff_sg \reg_w_7_reg[6]  ( .D(n45674), .CP(clk), .Q(reg_w_7[6]) );
  dff_sg \reg_w_7_reg[7]  ( .D(n45673), .CP(clk), .Q(reg_w_7[7]) );
  dff_sg \reg_w_7_reg[8]  ( .D(n45677), .CP(clk), .Q(reg_w_7[8]) );
  dff_sg \reg_w_7_reg[9]  ( .D(n45676), .CP(clk), .Q(reg_w_7[9]) );
  dff_sg \reg_w_7_reg[10]  ( .D(n45668), .CP(clk), .Q(reg_w_7[10]) );
  dff_sg \reg_w_7_reg[11]  ( .D(n45667), .CP(clk), .Q(reg_w_7[11]) );
  dff_sg \reg_w_7_reg[12]  ( .D(n45671), .CP(clk), .Q(reg_w_7[12]) );
  dff_sg \reg_w_7_reg[13]  ( .D(n45670), .CP(clk), .Q(reg_w_7[13]) );
  dff_sg \reg_w_7_reg[14]  ( .D(n45690), .CP(clk), .Q(reg_w_7[14]) );
  dff_sg \reg_w_7_reg[15]  ( .D(n45663), .CP(clk), .Q(reg_w_7[15]) );
  dff_sg \reg_w_7_reg[16]  ( .D(n45791), .CP(clk), .Q(reg_w_7[16]) );
  dff_sg \reg_w_7_reg[17]  ( .D(n45863), .CP(clk), .Q(reg_w_7[17]) );
  dff_sg \reg_w_7_reg[18]  ( .D(n45815), .CP(clk), .Q(reg_w_7[18]) );
  dff_sg \reg_w_7_reg[19]  ( .D(n45814), .CP(clk), .Q(reg_w_7[19]) );
  dff_sg \reg_w_8_reg[0]  ( .D(n45818), .CP(clk), .Q(reg_w_8[0]) );
  dff_sg \reg_w_8_reg[1]  ( .D(n45817), .CP(clk), .Q(reg_w_8[1]) );
  dff_sg \reg_w_8_reg[2]  ( .D(n45926), .CP(clk), .Q(reg_w_8[2]) );
  dff_sg \reg_w_8_reg[3]  ( .D(n45925), .CP(clk), .Q(reg_w_8[3]) );
  dff_sg \reg_w_8_reg[4]  ( .D(n45929), .CP(clk), .Q(reg_w_8[4]) );
  dff_sg \reg_w_8_reg[5]  ( .D(n45928), .CP(clk), .Q(reg_w_8[5]) );
  dff_sg \reg_w_8_reg[6]  ( .D(n45920), .CP(clk), .Q(reg_w_8[6]) );
  dff_sg \reg_w_8_reg[7]  ( .D(n45919), .CP(clk), .Q(reg_w_8[7]) );
  dff_sg \reg_w_8_reg[8]  ( .D(n45923), .CP(clk), .Q(reg_w_8[8]) );
  dff_sg \reg_w_8_reg[9]  ( .D(n45922), .CP(clk), .Q(reg_w_8[9]) );
  dff_sg \reg_w_8_reg[10]  ( .D(n45938), .CP(clk), .Q(reg_w_8[10]) );
  dff_sg \reg_w_8_reg[11]  ( .D(n45937), .CP(clk), .Q(reg_w_8[11]) );
  dff_sg \reg_w_8_reg[12]  ( .D(n45941), .CP(clk), .Q(reg_w_8[12]) );
  dff_sg \reg_w_8_reg[13]  ( .D(n45940), .CP(clk), .Q(reg_w_8[13]) );
  dff_sg \reg_w_8_reg[14]  ( .D(n45932), .CP(clk), .Q(reg_w_8[14]) );
  dff_sg \reg_w_8_reg[15]  ( .D(n45931), .CP(clk), .Q(reg_w_8[15]) );
  dff_sg \reg_w_8_reg[16]  ( .D(n45935), .CP(clk), .Q(reg_w_8[16]) );
  dff_sg \reg_w_8_reg[17]  ( .D(n45934), .CP(clk), .Q(reg_w_8[17]) );
  dff_sg \reg_w_8_reg[18]  ( .D(n45902), .CP(clk), .Q(reg_w_8[18]) );
  dff_sg \reg_w_8_reg[19]  ( .D(n45901), .CP(clk), .Q(reg_w_8[19]) );
  dff_sg \reg_w_9_reg[0]  ( .D(n45905), .CP(clk), .Q(reg_w_9[0]) );
  dff_sg \reg_w_9_reg[1]  ( .D(n45904), .CP(clk), .Q(reg_w_9[1]) );
  dff_sg \reg_w_9_reg[2]  ( .D(n45896), .CP(clk), .Q(reg_w_9[2]) );
  dff_sg \reg_w_9_reg[3]  ( .D(n45895), .CP(clk), .Q(reg_w_9[3]) );
  dff_sg \reg_w_9_reg[4]  ( .D(n45899), .CP(clk), .Q(reg_w_9[4]) );
  dff_sg \reg_w_9_reg[5]  ( .D(n45898), .CP(clk), .Q(reg_w_9[5]) );
  dff_sg \reg_w_9_reg[6]  ( .D(n45914), .CP(clk), .Q(reg_w_9[6]) );
  dff_sg \reg_w_9_reg[7]  ( .D(n45913), .CP(clk), .Q(reg_w_9[7]) );
  dff_sg \reg_w_9_reg[8]  ( .D(n45917), .CP(clk), .Q(reg_w_9[8]) );
  dff_sg \reg_w_9_reg[9]  ( .D(n45916), .CP(clk), .Q(reg_w_9[9]) );
  dff_sg \reg_w_9_reg[10]  ( .D(n45908), .CP(clk), .Q(reg_w_9[10]) );
  dff_sg \reg_w_9_reg[11]  ( .D(n45907), .CP(clk), .Q(reg_w_9[11]) );
  dff_sg \reg_w_9_reg[12]  ( .D(n45911), .CP(clk), .Q(reg_w_9[12]) );
  dff_sg \reg_w_9_reg[13]  ( .D(n45910), .CP(clk), .Q(reg_w_9[13]) );
  dff_sg \reg_w_9_reg[14]  ( .D(n46130), .CP(clk), .Q(reg_w_9[14]) );
  dff_sg \reg_w_9_reg[15]  ( .D(n46129), .CP(clk), .Q(reg_w_9[15]) );
  dff_sg \reg_w_9_reg[16]  ( .D(n46133), .CP(clk), .Q(reg_w_9[16]) );
  dff_sg \reg_w_9_reg[17]  ( .D(n46132), .CP(clk), .Q(reg_w_9[17]) );
  dff_sg \reg_w_9_reg[18]  ( .D(n46124), .CP(clk), .Q(reg_w_9[18]) );
  dff_sg \reg_w_9_reg[19]  ( .D(n46123), .CP(clk), .Q(reg_w_9[19]) );
  dff_sg \reg_w_10_reg[0]  ( .D(n46127), .CP(clk), .Q(reg_w_10[0]) );
  dff_sg \reg_w_10_reg[1]  ( .D(n46126), .CP(clk), .Q(reg_w_10[1]) );
  dff_sg \reg_w_10_reg[2]  ( .D(n46142), .CP(clk), .Q(reg_w_10[2]) );
  dff_sg \reg_w_10_reg[3]  ( .D(n46141), .CP(clk), .Q(reg_w_10[3]) );
  dff_sg \reg_w_10_reg[4]  ( .D(n46145), .CP(clk), .Q(reg_w_10[4]) );
  dff_sg \reg_w_10_reg[5]  ( .D(n46144), .CP(clk), .Q(reg_w_10[5]) );
  dff_sg \reg_w_10_reg[6]  ( .D(n46136), .CP(clk), .Q(reg_w_10[6]) );
  dff_sg \reg_w_10_reg[7]  ( .D(n46135), .CP(clk), .Q(reg_w_10[7]) );
  dff_sg \reg_w_10_reg[8]  ( .D(n46139), .CP(clk), .Q(reg_w_10[8]) );
  dff_sg \reg_w_10_reg[9]  ( .D(n46138), .CP(clk), .Q(reg_w_10[9]) );
  dff_sg \reg_w_10_reg[10]  ( .D(n46106), .CP(clk), .Q(reg_w_10[10]) );
  dff_sg \reg_w_10_reg[11]  ( .D(n46105), .CP(clk), .Q(reg_w_10[11]) );
  dff_sg \reg_w_10_reg[12]  ( .D(n46109), .CP(clk), .Q(reg_w_10[12]) );
  dff_sg \reg_w_10_reg[13]  ( .D(n46108), .CP(clk), .Q(reg_w_10[13]) );
  dff_sg \reg_w_10_reg[14]  ( .D(n46100), .CP(clk), .Q(reg_w_10[14]) );
  dff_sg \reg_w_10_reg[15]  ( .D(n46099), .CP(clk), .Q(reg_w_10[15]) );
  dff_sg \reg_w_10_reg[16]  ( .D(n46103), .CP(clk), .Q(reg_w_10[16]) );
  dff_sg \reg_w_10_reg[17]  ( .D(n46102), .CP(clk), .Q(reg_w_10[17]) );
  dff_sg \reg_w_10_reg[18]  ( .D(n46118), .CP(clk), .Q(reg_w_10[18]) );
  dff_sg \reg_w_10_reg[19]  ( .D(n46117), .CP(clk), .Q(reg_w_10[19]) );
  dff_sg \reg_w_11_reg[0]  ( .D(n46121), .CP(clk), .Q(reg_w_11[0]) );
  dff_sg \reg_w_11_reg[1]  ( .D(n46120), .CP(clk), .Q(reg_w_11[1]) );
  dff_sg \reg_w_11_reg[2]  ( .D(n46112), .CP(clk), .Q(reg_w_11[2]) );
  dff_sg \reg_w_11_reg[3]  ( .D(n46111), .CP(clk), .Q(reg_w_11[3]) );
  dff_sg \reg_w_11_reg[4]  ( .D(n46115), .CP(clk), .Q(reg_w_11[4]) );
  dff_sg \reg_w_11_reg[5]  ( .D(n46114), .CP(clk), .Q(reg_w_11[5]) );
  dff_sg \reg_w_11_reg[6]  ( .D(n46178), .CP(clk), .Q(reg_w_11[6]) );
  dff_sg \reg_w_11_reg[7]  ( .D(n46177), .CP(clk), .Q(reg_w_11[7]) );
  dff_sg \reg_w_11_reg[8]  ( .D(n46181), .CP(clk), .Q(reg_w_11[8]) );
  dff_sg \reg_w_11_reg[9]  ( .D(n46180), .CP(clk), .Q(reg_w_11[9]) );
  dff_sg \reg_w_11_reg[10]  ( .D(n46172), .CP(clk), .Q(reg_w_11[10]) );
  dff_sg \reg_w_11_reg[11]  ( .D(n46171), .CP(clk), .Q(reg_w_11[11]) );
  dff_sg \reg_w_11_reg[12]  ( .D(n46175), .CP(clk), .Q(reg_w_11[12]) );
  dff_sg \reg_w_11_reg[13]  ( .D(n46174), .CP(clk), .Q(reg_w_11[13]) );
  dff_sg \reg_w_11_reg[14]  ( .D(n46190), .CP(clk), .Q(reg_w_11[14]) );
  dff_sg \reg_w_11_reg[15]  ( .D(n46189), .CP(clk), .Q(reg_w_11[15]) );
  dff_sg \reg_w_11_reg[16]  ( .D(n46193), .CP(clk), .Q(reg_w_11[16]) );
  dff_sg \reg_w_11_reg[17]  ( .D(n46192), .CP(clk), .Q(reg_w_11[17]) );
  dff_sg \reg_w_11_reg[18]  ( .D(n46184), .CP(clk), .Q(reg_w_11[18]) );
  dff_sg \reg_w_11_reg[19]  ( .D(n46183), .CP(clk), .Q(reg_w_11[19]) );
  dff_sg \reg_w_12_reg[0]  ( .D(n46187), .CP(clk), .Q(reg_w_12[0]) );
  dff_sg \reg_w_12_reg[1]  ( .D(n46186), .CP(clk), .Q(reg_w_12[1]) );
  dff_sg \reg_w_12_reg[2]  ( .D(n46154), .CP(clk), .Q(reg_w_12[2]) );
  dff_sg \reg_w_12_reg[3]  ( .D(n46153), .CP(clk), .Q(reg_w_12[3]) );
  dff_sg \reg_w_12_reg[4]  ( .D(n46157), .CP(clk), .Q(reg_w_12[4]) );
  dff_sg \reg_w_12_reg[5]  ( .D(n46156), .CP(clk), .Q(reg_w_12[5]) );
  dff_sg \reg_w_12_reg[6]  ( .D(n46148), .CP(clk), .Q(reg_w_12[6]) );
  dff_sg \reg_w_12_reg[7]  ( .D(n46147), .CP(clk), .Q(reg_w_12[7]) );
  dff_sg \reg_w_12_reg[8]  ( .D(n46151), .CP(clk), .Q(reg_w_12[8]) );
  dff_sg \reg_w_12_reg[9]  ( .D(n46150), .CP(clk), .Q(reg_w_12[9]) );
  dff_sg \reg_w_12_reg[10]  ( .D(n46166), .CP(clk), .Q(reg_w_12[10]) );
  dff_sg \reg_w_12_reg[11]  ( .D(n46165), .CP(clk), .Q(reg_w_12[11]) );
  dff_sg \reg_w_12_reg[12]  ( .D(n46169), .CP(clk), .Q(reg_w_12[12]) );
  dff_sg \reg_w_12_reg[13]  ( .D(n46168), .CP(clk), .Q(reg_w_12[13]) );
  dff_sg \reg_w_12_reg[14]  ( .D(n46160), .CP(clk), .Q(reg_w_12[14]) );
  dff_sg \reg_w_12_reg[15]  ( .D(n46159), .CP(clk), .Q(reg_w_12[15]) );
  dff_sg \reg_w_12_reg[16]  ( .D(n46163), .CP(clk), .Q(reg_w_12[16]) );
  dff_sg \reg_w_12_reg[17]  ( .D(n46162), .CP(clk), .Q(reg_w_12[17]) );
  dff_sg \reg_w_12_reg[18]  ( .D(n46082), .CP(clk), .Q(reg_w_12[18]) );
  dff_sg \reg_w_12_reg[19]  ( .D(n46081), .CP(clk), .Q(reg_w_12[19]) );
  dff_sg \reg_w_13_reg[0]  ( .D(n46085), .CP(clk), .Q(reg_w_13[0]) );
  dff_sg \reg_w_13_reg[1]  ( .D(n46084), .CP(clk), .Q(reg_w_13[1]) );
  dff_sg \reg_w_13_reg[2]  ( .D(n46076), .CP(clk), .Q(reg_w_13[2]) );
  dff_sg \reg_w_13_reg[3]  ( .D(n46075), .CP(clk), .Q(reg_w_13[3]) );
  dff_sg \reg_w_13_reg[4]  ( .D(n46079), .CP(clk), .Q(reg_w_13[4]) );
  dff_sg \reg_w_13_reg[5]  ( .D(n46078), .CP(clk), .Q(reg_w_13[5]) );
  dff_sg \reg_w_13_reg[6]  ( .D(n46094), .CP(clk), .Q(reg_w_13[6]) );
  dff_sg \reg_w_13_reg[7]  ( .D(n46093), .CP(clk), .Q(reg_w_13[7]) );
  dff_sg \reg_w_13_reg[8]  ( .D(n46097), .CP(clk), .Q(reg_w_13[8]) );
  dff_sg \reg_w_13_reg[9]  ( .D(n46096), .CP(clk), .Q(reg_w_13[9]) );
  dff_sg \reg_w_13_reg[10]  ( .D(n46088), .CP(clk), .Q(reg_w_13[10]) );
  dff_sg \reg_w_13_reg[11]  ( .D(n46087), .CP(clk), .Q(reg_w_13[11]) );
  dff_sg \reg_w_13_reg[12]  ( .D(n46091), .CP(clk), .Q(reg_w_13[12]) );
  dff_sg \reg_w_13_reg[13]  ( .D(n46090), .CP(clk), .Q(reg_w_13[13]) );
  dff_sg \reg_w_13_reg[14]  ( .D(n46058), .CP(clk), .Q(reg_w_13[14]) );
  dff_sg \reg_w_13_reg[15]  ( .D(n46057), .CP(clk), .Q(reg_w_13[15]) );
  dff_sg \reg_w_13_reg[16]  ( .D(n46061), .CP(clk), .Q(reg_w_13[16]) );
  dff_sg \reg_w_13_reg[17]  ( .D(n46060), .CP(clk), .Q(reg_w_13[17]) );
  dff_sg \reg_w_13_reg[18]  ( .D(n46052), .CP(clk), .Q(reg_w_13[18]) );
  dff_sg \reg_w_13_reg[19]  ( .D(n46051), .CP(clk), .Q(reg_w_13[19]) );
  dff_sg \reg_w_14_reg[0]  ( .D(n46055), .CP(clk), .Q(reg_w_14[0]) );
  dff_sg \reg_w_14_reg[1]  ( .D(n46054), .CP(clk), .Q(reg_w_14[1]) );
  dff_sg \reg_w_14_reg[2]  ( .D(n46070), .CP(clk), .Q(reg_w_14[2]) );
  dff_sg \reg_w_14_reg[3]  ( .D(n46069), .CP(clk), .Q(reg_w_14[3]) );
  dff_sg \reg_w_14_reg[4]  ( .D(n46073), .CP(clk), .Q(reg_w_14[4]) );
  dff_sg \reg_w_14_reg[5]  ( .D(n46072), .CP(clk), .Q(reg_w_14[5]) );
  dff_sg \reg_w_14_reg[6]  ( .D(n46064), .CP(clk), .Q(reg_w_14[6]) );
  dff_sg \reg_w_14_reg[7]  ( .D(n46063), .CP(clk), .Q(reg_w_14[7]) );
  dff_sg \reg_w_14_reg[8]  ( .D(n46067), .CP(clk), .Q(reg_w_14[8]) );
  dff_sg \reg_w_14_reg[9]  ( .D(n46066), .CP(clk), .Q(reg_w_14[9]) );
  dff_sg \reg_w_14_reg[10]  ( .D(n46046), .CP(clk), .Q(reg_w_14[10]) );
  dff_sg \reg_w_14_reg[11]  ( .D(n46045), .CP(clk), .Q(reg_w_14[11]) );
  dff_sg \reg_w_14_reg[12]  ( .D(n46049), .CP(clk), .Q(reg_w_14[12]) );
  dff_sg \reg_w_14_reg[13]  ( .D(n46048), .CP(clk), .Q(reg_w_14[13]) );
  dff_sg \reg_w_14_reg[14]  ( .D(n46040), .CP(clk), .Q(reg_w_14[14]) );
  dff_sg \reg_w_14_reg[15]  ( .D(n46039), .CP(clk), .Q(reg_w_14[15]) );
  dff_sg \reg_w_14_reg[16]  ( .D(n46043), .CP(clk), .Q(reg_w_14[16]) );
  dff_sg \reg_w_14_reg[17]  ( .D(n46042), .CP(clk), .Q(reg_w_14[17]) );
  dff_sg \reg_w_14_reg[18]  ( .D(n45716), .CP(clk), .Q(reg_w_14[18]) );
  dff_sg \reg_w_14_reg[19]  ( .D(n45715), .CP(clk), .Q(reg_w_14[19]) );
  dff_sg \reg_w_15_reg[0]  ( .D(n45719), .CP(clk), .Q(reg_w_15[0]) );
  dff_sg \reg_w_15_reg[1]  ( .D(n45718), .CP(clk), .Q(reg_w_15[1]) );
  dff_sg \reg_w_15_reg[2]  ( .D(n45978), .CP(clk), .Q(reg_w_15[2]) );
  dff_sg \reg_w_15_reg[3]  ( .D(n45951), .CP(clk), .Q(reg_w_15[3]) );
  dff_sg \reg_w_15_reg[4]  ( .D(n45948), .CP(clk), .Q(reg_w_15[4]) );
  dff_sg \reg_w_15_reg[5]  ( .D(n45945), .CP(clk), .Q(reg_w_15[5]) );
  dff_sg \reg_w_15_reg[6]  ( .D(n45714), .CP(clk), .Q(reg_w_15[6]) );
  dff_sg \reg_w_15_reg[7]  ( .D(n45942), .CP(clk), .Q(reg_w_15[7]) );
  dff_sg \reg_w_15_reg[8]  ( .D(n45713), .CP(clk), .Q(reg_w_15[8]) );
  dff_sg \reg_w_15_reg[9]  ( .D(n46047), .CP(clk), .Q(reg_w_15[9]) );
  dff_sg \reg_w_15_reg[10]  ( .D(n46044), .CP(clk), .Q(reg_w_15[10]) );
  dff_sg \reg_w_15_reg[11]  ( .D(n45717), .CP(clk), .Q(reg_w_15[11]) );
  dff_sg \reg_w_15_reg[12]  ( .D(n46041), .CP(clk), .Q(reg_w_15[12]) );
  dff_sg \reg_w_15_reg[13]  ( .D(n46038), .CP(clk), .Q(reg_w_15[13]) );
  dff_sg \reg_w_15_reg[14]  ( .D(n45666), .CP(clk), .Q(reg_w_15[14]) );
  dff_sg \reg_w_15_reg[15]  ( .D(n45981), .CP(clk), .Q(reg_w_15[15]) );
  dff_sg \reg_w_15_reg[16]  ( .D(n46110), .CP(clk), .Q(reg_w_15[16]) );
  dff_sg \reg_w_15_reg[17]  ( .D(n46125), .CP(clk), .Q(reg_w_15[17]) );
  dff_sg \reg_w_15_reg[18]  ( .D(n46161), .CP(clk), .Q(reg_w_15[18]) );
  dff_sg \reg_w_15_reg[19]  ( .D(n45669), .CP(clk), .Q(reg_w_15[19]) );
  dff_sg input_taken_reg ( .D(n10398), .CP(clk), .Q(n69266) );
  dff_sg \reg_ii_4_reg[18]  ( .D(n44476), .CP(clk), .Q(reg_ii_4[18]) );
  dff_sg \reg_iii_4_reg[18]  ( .D(n45436), .CP(clk), .Q(reg_iii_4[18]) );
  dff_sg \reg_ii_4_reg[17]  ( .D(n45342), .CP(clk), .Q(reg_ii_4[17]) );
  dff_sg \reg_iii_4_reg[17]  ( .D(n44669), .CP(clk), .Q(reg_iii_4[17]) );
  dff_sg \reg_ii_4_reg[16]  ( .D(n45501), .CP(clk), .Q(reg_ii_4[16]) );
  dff_sg \reg_iii_4_reg[16]  ( .D(n45403), .CP(clk), .Q(reg_iii_4[16]) );
  dff_sg \reg_ii_4_reg[15]  ( .D(n45502), .CP(clk), .Q(reg_ii_4[15]) );
  dff_sg \reg_iii_4_reg[15]  ( .D(n44660), .CP(clk), .Q(reg_iii_4[15]) );
  dff_sg \reg_ii_4_reg[14]  ( .D(n45331), .CP(clk), .Q(reg_ii_4[14]) );
  dff_sg \reg_iii_4_reg[14]  ( .D(n44654), .CP(clk), .Q(reg_iii_4[14]) );
  dff_sg \reg_ii_4_reg[13]  ( .D(n45332), .CP(clk), .Q(reg_ii_4[13]) );
  dff_sg \reg_iii_4_reg[13]  ( .D(n44567), .CP(clk), .Q(reg_iii_4[13]) );
  dff_sg \reg_ii_4_reg[12]  ( .D(n45329), .CP(clk), .Q(reg_ii_4[12]) );
  dff_sg \reg_iii_4_reg[12]  ( .D(n45407), .CP(clk), .Q(reg_iii_4[12]) );
  dff_sg \reg_ii_4_reg[11]  ( .D(n45330), .CP(clk), .Q(reg_ii_4[11]) );
  dff_sg \reg_iii_4_reg[11]  ( .D(n44666), .CP(clk), .Q(reg_iii_4[11]) );
  dff_sg \reg_ii_4_reg[10]  ( .D(n45335), .CP(clk), .Q(reg_ii_4[10]) );
  dff_sg \reg_iii_4_reg[10]  ( .D(n44690), .CP(clk), .Q(reg_iii_4[10]) );
  dff_sg \reg_ii_4_reg[9]  ( .D(n45336), .CP(clk), .Q(reg_ii_4[9]) );
  dff_sg \reg_iii_4_reg[9]  ( .D(n44777), .CP(clk), .Q(reg_iii_4[9]) );
  dff_sg \reg_ii_4_reg[8]  ( .D(n45333), .CP(clk), .Q(reg_ii_4[8]) );
  dff_sg \reg_iii_4_reg[8]  ( .D(n45326), .CP(clk), .Q(reg_iii_4[8]) );
  dff_sg \reg_ii_4_reg[7]  ( .D(n45334), .CP(clk), .Q(reg_ii_4[7]) );
  dff_sg \reg_iii_4_reg[7]  ( .D(n44735), .CP(clk), .Q(reg_iii_4[7]) );
  dff_sg \reg_ii_4_reg[6]  ( .D(n45302), .CP(clk), .Q(reg_ii_4[6]) );
  dff_sg \reg_iii_4_reg[6]  ( .D(n45328), .CP(clk), .Q(reg_iii_4[6]) );
  dff_sg \reg_ii_4_reg[5]  ( .D(n45303), .CP(clk), .Q(reg_ii_4[5]) );
  dff_sg \reg_iii_4_reg[5]  ( .D(n44741), .CP(clk), .Q(reg_iii_4[5]) );
  dff_sg \reg_ii_4_reg[4]  ( .D(n45300), .CP(clk), .Q(reg_ii_4[4]) );
  dff_sg \reg_iii_4_reg[4]  ( .D(n44723), .CP(clk), .Q(reg_iii_4[4]) );
  dff_sg \reg_ii_4_reg[3]  ( .D(n45301), .CP(clk), .Q(reg_ii_4[3]) );
  dff_sg \reg_iii_4_reg[3]  ( .D(n45338), .CP(clk), .Q(reg_iii_4[3]) );
  dff_sg \reg_ii_4_reg[2]  ( .D(n45306), .CP(clk), .Q(reg_ii_4[2]) );
  dff_sg \reg_iii_4_reg[2]  ( .D(n45339), .CP(clk), .Q(reg_iii_4[2]) );
  dff_sg \reg_ii_4_reg[1]  ( .D(n45307), .CP(clk), .Q(reg_ii_4[1]) );
  dff_sg \reg_iii_4_reg[1]  ( .D(n45073), .CP(clk), .Q(reg_iii_4[1]) );
  dff_sg \reg_ii_4_reg[0]  ( .D(n45304), .CP(clk), .Q(reg_ii_4[0]) );
  dff_sg \reg_iii_4_reg[0]  ( .D(n45337), .CP(clk), .Q(reg_iii_4[0]) );
  dff_sg \reg_ii_3_reg[19]  ( .D(n45310), .CP(clk), .Q(reg_ii_3[19]) );
  dff_sg \reg_iii_3_reg[19]  ( .D(n45305), .CP(clk), .Q(reg_iii_3[19]) );
  dff_sg \reg_ii_3_reg[18]  ( .D(n45315), .CP(clk), .Q(reg_ii_3[18]) );
  dff_sg \reg_iii_3_reg[18]  ( .D(n45295), .CP(clk), .Q(reg_iii_3[18]) );
  dff_sg \reg_ii_3_reg[17]  ( .D(n45316), .CP(clk), .Q(reg_ii_3[17]) );
  dff_sg \reg_iii_3_reg[17]  ( .D(n45296), .CP(clk), .Q(reg_iii_3[17]) );
  dff_sg \reg_ii_3_reg[16]  ( .D(n45107), .CP(clk), .Q(reg_ii_3[16]) );
  dff_sg \reg_iii_3_reg[16]  ( .D(n44478), .CP(clk), .Q(reg_iii_3[16]) );
  dff_sg \reg_ii_3_reg[15]  ( .D(n45104), .CP(clk), .Q(reg_ii_3[15]) );
  dff_sg \reg_iii_3_reg[15]  ( .D(n44477), .CP(clk), .Q(reg_iii_3[15]) );
  dff_sg \reg_ii_3_reg[14]  ( .D(n45101), .CP(clk), .Q(reg_ii_3[14]) );
  dff_sg \reg_iii_3_reg[14]  ( .D(n45075), .CP(clk), .Q(reg_iii_3[14]) );
  dff_sg \reg_ii_3_reg[13]  ( .D(n45384), .CP(clk), .Q(reg_ii_3[13]) );
  dff_sg \reg_iii_3_reg[13]  ( .D(n45074), .CP(clk), .Q(reg_iii_3[13]) );
  dff_sg \reg_ii_3_reg[12]  ( .D(n45114), .CP(clk), .Q(reg_ii_3[12]) );
  dff_sg \reg_iii_3_reg[12]  ( .D(n45298), .CP(clk), .Q(reg_iii_3[12]) );
  dff_sg \reg_ii_3_reg[11]  ( .D(n45383), .CP(clk), .Q(reg_ii_3[11]) );
  dff_sg \reg_iii_3_reg[11]  ( .D(n45299), .CP(clk), .Q(reg_iii_3[11]) );
  dff_sg \reg_ii_3_reg[10]  ( .D(n45117), .CP(clk), .Q(reg_ii_3[10]) );
  dff_sg \reg_iii_3_reg[10]  ( .D(n45320), .CP(clk), .Q(reg_iii_3[10]) );
  dff_sg \reg_ii_3_reg[9]  ( .D(n45110), .CP(clk), .Q(reg_ii_3[9]) );
  dff_sg \reg_iii_3_reg[9]  ( .D(n45321), .CP(clk), .Q(reg_iii_3[9]) );
  dff_sg \reg_ii_3_reg[8]  ( .D(n45388), .CP(clk), .Q(reg_ii_3[8]) );
  dff_sg \reg_iii_3_reg[8]  ( .D(n45317), .CP(clk), .Q(reg_iii_3[8]) );
  dff_sg \reg_ii_3_reg[7]  ( .D(n45389), .CP(clk), .Q(reg_ii_3[7]) );
  dff_sg \reg_iii_3_reg[7]  ( .D(n45318), .CP(clk), .Q(reg_iii_3[7]) );
  dff_sg \reg_ii_3_reg[6]  ( .D(n45376), .CP(clk), .Q(reg_ii_3[6]) );
  dff_sg \reg_iii_3_reg[6]  ( .D(n45325), .CP(clk), .Q(reg_iii_3[6]) );
  dff_sg \reg_ii_3_reg[5]  ( .D(n45373), .CP(clk), .Q(reg_ii_3[5]) );
  dff_sg \reg_iii_3_reg[5]  ( .D(n44498), .CP(clk), .Q(reg_iii_3[5]) );
  dff_sg \reg_ii_3_reg[4]  ( .D(n45380), .CP(clk), .Q(reg_ii_3[4]) );
  dff_sg \reg_iii_3_reg[4]  ( .D(n45323), .CP(clk), .Q(reg_iii_3[4]) );
  dff_sg \reg_ii_3_reg[3]  ( .D(n45377), .CP(clk), .Q(reg_ii_3[3]) );
  dff_sg \reg_iii_3_reg[3]  ( .D(n45324), .CP(clk), .Q(reg_iii_3[3]) );
  dff_sg \reg_ii_3_reg[2]  ( .D(n45381), .CP(clk), .Q(reg_ii_3[2]) );
  dff_sg \reg_iii_3_reg[2]  ( .D(n45312), .CP(clk), .Q(reg_iii_3[2]) );
  dff_sg \reg_ii_3_reg[1]  ( .D(n45382), .CP(clk), .Q(reg_ii_3[1]) );
  dff_sg \reg_iii_3_reg[1]  ( .D(n45313), .CP(clk), .Q(reg_iii_3[1]) );
  dff_sg \reg_ii_3_reg[0]  ( .D(n45378), .CP(clk), .Q(reg_ii_3[0]) );
  dff_sg \reg_iii_3_reg[0]  ( .D(n45309), .CP(clk), .Q(reg_iii_3[0]) );
  dff_sg \reg_ii_2_reg[19]  ( .D(n44801), .CP(clk), .Q(reg_ii_2[19]) );
  dff_sg \reg_iii_2_reg[19]  ( .D(n45379), .CP(clk), .Q(reg_iii_2[19]) );
  dff_sg \reg_ii_2_reg[18]  ( .D(n45357), .CP(clk), .Q(reg_ii_2[18]) );
  dff_sg \reg_iii_2_reg[18]  ( .D(n45390), .CP(clk), .Q(reg_iii_2[18]) );
  dff_sg \reg_ii_2_reg[17]  ( .D(n45353), .CP(clk), .Q(reg_ii_2[17]) );
  dff_sg \reg_iii_2_reg[17]  ( .D(n45397), .CP(clk), .Q(reg_iii_2[17]) );
  dff_sg \reg_ii_2_reg[16]  ( .D(n45358), .CP(clk), .Q(reg_ii_2[16]) );
  dff_sg \reg_iii_2_reg[16]  ( .D(n45398), .CP(clk), .Q(reg_iii_2[16]) );
  dff_sg \reg_ii_2_reg[15]  ( .D(n45359), .CP(clk), .Q(reg_ii_2[15]) );
  dff_sg \reg_iii_2_reg[15]  ( .D(n45391), .CP(clk), .Q(reg_iii_2[15]) );
  dff_sg \reg_ii_2_reg[14]  ( .D(n45345), .CP(clk), .Q(reg_ii_2[14]) );
  dff_sg \reg_iii_2_reg[14]  ( .D(n45399), .CP(clk), .Q(reg_iii_2[14]) );
  dff_sg \reg_ii_2_reg[13]  ( .D(n45346), .CP(clk), .Q(reg_ii_2[13]) );
  dff_sg \reg_iii_2_reg[13]  ( .D(n45400), .CP(clk), .Q(reg_iii_2[13]) );
  dff_sg \reg_ii_2_reg[12]  ( .D(n45343), .CP(clk), .Q(reg_ii_2[12]) );
  dff_sg \reg_iii_2_reg[12]  ( .D(n44873), .CP(clk), .Q(reg_iii_2[12]) );
  dff_sg \reg_ii_2_reg[11]  ( .D(n45344), .CP(clk), .Q(reg_ii_2[11]) );
  dff_sg \reg_iii_2_reg[11]  ( .D(n44840), .CP(clk), .Q(reg_iii_2[11]) );
  dff_sg \reg_ii_2_reg[10]  ( .D(n45148), .CP(clk), .Q(reg_ii_2[10]) );
  dff_sg \reg_iii_2_reg[10]  ( .D(n45394), .CP(clk), .Q(reg_iii_2[10]) );
  dff_sg \reg_ii_2_reg[9]  ( .D(n45350), .CP(clk), .Q(reg_ii_2[9]) );
  dff_sg \reg_iii_2_reg[9]  ( .D(n44843), .CP(clk), .Q(reg_iii_2[9]) );
  dff_sg \reg_ii_2_reg[8]  ( .D(n45351), .CP(clk), .Q(reg_ii_2[8]) );
  dff_sg \reg_iii_2_reg[8]  ( .D(n44834), .CP(clk), .Q(reg_iii_2[8]) );
  dff_sg \reg_ii_2_reg[7]  ( .D(n45352), .CP(clk), .Q(reg_ii_2[7]) );
  dff_sg \reg_iii_2_reg[7]  ( .D(n45392), .CP(clk), .Q(reg_iii_2[7]) );
  dff_sg \reg_ii_2_reg[6]  ( .D(n45368), .CP(clk), .Q(reg_ii_2[6]) );
  dff_sg \reg_iii_2_reg[6]  ( .D(n45395), .CP(clk), .Q(reg_iii_2[6]) );
  dff_sg \reg_ii_2_reg[5]  ( .D(n45362), .CP(clk), .Q(reg_ii_2[5]) );
  dff_sg \reg_iii_2_reg[5]  ( .D(n45393), .CP(clk), .Q(reg_iii_2[5]) );
  dff_sg \reg_ii_2_reg[4]  ( .D(n45365), .CP(clk), .Q(reg_ii_2[4]) );
  dff_sg \reg_iii_2_reg[4]  ( .D(n44816), .CP(clk), .Q(reg_iii_2[4]) );
  dff_sg \reg_ii_2_reg[3]  ( .D(n45370), .CP(clk), .Q(reg_ii_2[3]) );
  dff_sg \reg_iii_2_reg[3]  ( .D(n45396), .CP(clk), .Q(reg_iii_2[3]) );
  dff_sg \reg_ii_2_reg[2]  ( .D(n45374), .CP(clk), .Q(reg_ii_2[2]) );
  dff_sg \reg_iii_2_reg[2]  ( .D(n45354), .CP(clk), .Q(reg_iii_2[2]) );
  dff_sg \reg_ii_2_reg[1]  ( .D(n45375), .CP(clk), .Q(reg_ii_2[1]) );
  dff_sg \reg_iii_2_reg[1]  ( .D(n45355), .CP(clk), .Q(reg_iii_2[1]) );
  dff_sg \reg_ii_2_reg[0]  ( .D(n45371), .CP(clk), .Q(reg_ii_2[0]) );
  dff_sg \reg_iii_2_reg[0]  ( .D(n44807), .CP(clk), .Q(reg_iii_2[0]) );
  dff_sg \reg_ii_1_reg[19]  ( .D(n45227), .CP(clk), .Q(reg_ii_1[19]) );
  dff_sg \reg_iii_1_reg[19]  ( .D(n45372), .CP(clk), .Q(reg_iii_1[19]) );
  dff_sg \reg_ii_1_reg[18]  ( .D(n45012), .CP(clk), .Q(reg_ii_1[18]) );
  dff_sg \reg_iii_1_reg[18]  ( .D(n45363), .CP(clk), .Q(reg_iii_1[18]) );
  dff_sg \reg_ii_1_reg[17]  ( .D(n44275), .CP(clk), .Q(reg_ii_1[17]) );
  dff_sg \reg_iii_1_reg[17]  ( .D(n45364), .CP(clk), .Q(reg_iii_1[17]) );
  dff_sg \reg_ii_1_reg[16]  ( .D(n45228), .CP(clk), .Q(reg_ii_1[16]) );
  dff_sg \reg_iii_1_reg[16]  ( .D(n45360), .CP(clk), .Q(reg_iii_1[16]) );
  dff_sg \reg_ii_1_reg[15]  ( .D(n44289), .CP(clk), .Q(reg_ii_1[15]) );
  dff_sg \reg_iii_1_reg[15]  ( .D(n45361), .CP(clk), .Q(reg_iii_1[15]) );
  dff_sg \reg_ii_1_reg[14]  ( .D(n44849), .CP(clk), .Q(reg_ii_1[14]) );
  dff_sg \reg_iii_1_reg[14]  ( .D(n45369), .CP(clk), .Q(reg_iii_1[14]) );
  dff_sg \reg_ii_1_reg[13]  ( .D(n44846), .CP(clk), .Q(reg_ii_1[13]) );
  dff_sg \reg_iii_1_reg[13]  ( .D(n44272), .CP(clk), .Q(reg_iii_1[13]) );
  dff_sg \reg_ii_1_reg[12]  ( .D(n45236), .CP(clk), .Q(reg_ii_1[12]) );
  dff_sg \reg_iii_1_reg[12]  ( .D(n45366), .CP(clk), .Q(reg_iii_1[12]) );
  dff_sg \reg_ii_1_reg[11]  ( .D(n44288), .CP(clk), .Q(reg_ii_1[11]) );
  dff_sg \reg_iii_1_reg[11]  ( .D(n45367), .CP(clk), .Q(reg_iii_1[11]) );
  dff_sg \reg_ii_1_reg[10]  ( .D(n45238), .CP(clk), .Q(reg_ii_1[10]) );
  dff_sg \reg_iii_1_reg[10]  ( .D(n45231), .CP(clk), .Q(reg_iii_1[10]) );
  dff_sg \reg_ii_1_reg[9]  ( .D(n45239), .CP(clk), .Q(reg_ii_1[9]) );
  dff_sg \reg_iii_1_reg[9]  ( .D(n45232), .CP(clk), .Q(reg_iii_1[9]) );
  dff_sg \reg_ii_1_reg[8]  ( .D(n44714), .CP(clk), .Q(reg_ii_1[8]) );
  dff_sg \reg_iii_1_reg[8]  ( .D(n45229), .CP(clk), .Q(reg_iii_1[8]) );
  dff_sg \reg_ii_1_reg[7]  ( .D(n44284), .CP(clk), .Q(reg_ii_1[7]) );
  dff_sg \reg_iii_1_reg[7]  ( .D(n45230), .CP(clk), .Q(reg_iii_1[7]) );
  dff_sg \reg_ii_1_reg[6]  ( .D(n44630), .CP(clk), .Q(reg_ii_1[6]) );
  dff_sg \reg_iii_1_reg[6]  ( .D(n45234), .CP(clk), .Q(reg_iii_1[6]) );
  dff_sg \reg_ii_1_reg[5]  ( .D(n44762), .CP(clk), .Q(reg_ii_1[5]) );
  dff_sg \reg_iii_1_reg[5]  ( .D(n45235), .CP(clk), .Q(reg_iii_1[5]) );
  dff_sg \reg_ii_1_reg[4]  ( .D(n44286), .CP(clk), .Q(reg_ii_1[4]) );
  dff_sg \reg_iii_1_reg[4]  ( .D(n45233), .CP(clk), .Q(reg_iii_1[4]) );
  dff_sg \reg_ii_1_reg[3]  ( .D(n44771), .CP(clk), .Q(reg_ii_1[3]) );
  dff_sg \reg_iii_1_reg[3]  ( .D(n44615), .CP(clk), .Q(reg_iii_1[3]) );
  dff_sg \reg_ii_1_reg[2]  ( .D(n44831), .CP(clk), .Q(reg_ii_1[2]) );
  dff_sg \reg_iii_1_reg[2]  ( .D(n44991), .CP(clk), .Q(reg_iii_1[2]) );
  dff_sg \reg_ii_1_reg[1]  ( .D(n44813), .CP(clk), .Q(reg_ii_1[1]) );
  dff_sg \reg_iii_1_reg[1]  ( .D(n44287), .CP(clk), .Q(reg_iii_1[1]) );
  dff_sg \reg_ii_1_reg[0]  ( .D(n44858), .CP(clk), .Q(reg_ii_1[0]) );
  dff_sg \reg_iii_1_reg[0]  ( .D(n45226), .CP(clk), .Q(reg_iii_1[0]) );
  dff_sg \reg_ii_0_reg[19]  ( .D(n44882), .CP(clk), .Q(reg_ii_0[19]) );
  dff_sg \reg_iii_0_reg[19]  ( .D(n44789), .CP(clk), .Q(reg_iii_0[19]) );
  dff_sg \reg_ii_0_reg[18]  ( .D(n44648), .CP(clk), .Q(reg_ii_0[18]) );
  dff_sg \reg_iii_0_reg[18]  ( .D(n44988), .CP(clk), .Q(reg_iii_0[18]) );
  dff_sg \reg_ii_0_reg[17]  ( .D(n45224), .CP(clk), .Q(reg_ii_0[17]) );
  dff_sg \reg_iii_0_reg[17]  ( .D(n45217), .CP(clk), .Q(reg_iii_0[17]) );
  dff_sg \reg_ii_0_reg[16]  ( .D(n44281), .CP(clk), .Q(reg_ii_0[16]) );
  dff_sg \reg_iii_0_reg[16]  ( .D(n44322), .CP(clk), .Q(reg_iii_0[16]) );
  dff_sg \reg_ii_0_reg[15]  ( .D(n44900), .CP(clk), .Q(reg_ii_0[15]) );
  dff_sg \reg_iii_0_reg[15]  ( .D(n44323), .CP(clk), .Q(reg_iii_0[15]) );
  dff_sg \reg_ii_0_reg[14]  ( .D(n45221), .CP(clk), .Q(reg_ii_0[14]) );
  dff_sg \reg_iii_0_reg[14]  ( .D(n44531), .CP(clk), .Q(reg_iii_0[14]) );
  dff_sg \reg_ii_0_reg[13]  ( .D(n44963), .CP(clk), .Q(reg_ii_0[13]) );
  dff_sg \reg_iii_0_reg[13]  ( .D(n44324), .CP(clk), .Q(reg_iii_0[13]) );
  dff_sg \reg_ii_0_reg[12]  ( .D(n45219), .CP(clk), .Q(reg_ii_0[12]) );
  dff_sg \reg_iii_0_reg[12]  ( .D(n45218), .CP(clk), .Q(reg_iii_0[12]) );
  dff_sg \reg_ii_0_reg[11]  ( .D(n45220), .CP(clk), .Q(reg_ii_0[11]) );
  dff_sg \reg_iii_0_reg[11]  ( .D(n44618), .CP(clk), .Q(reg_iii_0[11]) );
  dff_sg \reg_ii_0_reg[10]  ( .D(n44909), .CP(clk), .Q(reg_ii_0[10]) );
  dff_sg \reg_iii_0_reg[10]  ( .D(n45214), .CP(clk), .Q(reg_iii_0[10]) );
  dff_sg \reg_ii_0_reg[9]  ( .D(n44942), .CP(clk), .Q(reg_ii_0[9]) );
  dff_sg \reg_iii_0_reg[9]  ( .D(n45215), .CP(clk), .Q(reg_iii_0[9]) );
  dff_sg \reg_ii_0_reg[8]  ( .D(n45222), .CP(clk), .Q(reg_ii_0[8]) );
  dff_sg \reg_iii_0_reg[8]  ( .D(n44891), .CP(clk), .Q(reg_iii_0[8]) );
  dff_sg \reg_ii_0_reg[7]  ( .D(n45223), .CP(clk), .Q(reg_ii_0[7]) );
  dff_sg \reg_iii_0_reg[7]  ( .D(n44795), .CP(clk), .Q(reg_iii_0[7]) );
  dff_sg \reg_ii_0_reg[6]  ( .D(n45276), .CP(clk), .Q(reg_ii_0[6]) );
  dff_sg \reg_iii_0_reg[6]  ( .D(n44804), .CP(clk), .Q(reg_iii_0[6]) );
  dff_sg \reg_ii_0_reg[5]  ( .D(n45277), .CP(clk), .Q(reg_ii_0[5]) );
  dff_sg \reg_iii_0_reg[5]  ( .D(n44798), .CP(clk), .Q(reg_iii_0[5]) );
  dff_sg \reg_ii_0_reg[4]  ( .D(n45274), .CP(clk), .Q(reg_ii_0[4]) );
  dff_sg \reg_iii_0_reg[4]  ( .D(n45216), .CP(clk), .Q(reg_iii_0[4]) );
  dff_sg \reg_ii_0_reg[3]  ( .D(n45275), .CP(clk), .Q(reg_ii_0[3]) );
  dff_sg \reg_iii_0_reg[3]  ( .D(n44620), .CP(clk), .Q(reg_iii_0[3]) );
  dff_sg \reg_ii_0_reg[2]  ( .D(n45278), .CP(clk), .Q(reg_ii_0[2]) );
  dff_sg \reg_iii_0_reg[2]  ( .D(n44750), .CP(clk), .Q(reg_iii_0[2]) );
  dff_sg \reg_ii_0_reg[1]  ( .D(n45279), .CP(clk), .Q(reg_ii_0[1]) );
  dff_sg \reg_iii_0_reg[1]  ( .D(n44753), .CP(clk), .Q(reg_iii_0[1]) );
  dff_sg \reg_ii_0_reg[0]  ( .D(n44530), .CP(clk), .Q(reg_ii_0[0]) );
  dff_sg \reg_iii_0_reg[0]  ( .D(n44619), .CP(clk), .Q(reg_iii_0[0]) );
  dff_sg \reg_ii_9_reg[17]  ( .D(n45281), .CP(clk), .Q(reg_ii_9[17]) );
  dff_sg \reg_iii_9_reg[17]  ( .D(n44924), .CP(clk), .Q(reg_iii_9[17]) );
  dff_sg \reg_ii_9_reg[16]  ( .D(n45287), .CP(clk), .Q(reg_ii_9[16]) );
  dff_sg \reg_iii_9_reg[16]  ( .D(n44975), .CP(clk), .Q(reg_iii_9[16]) );
  dff_sg \reg_ii_9_reg[15]  ( .D(n45288), .CP(clk), .Q(reg_ii_9[15]) );
  dff_sg \reg_iii_9_reg[15]  ( .D(n44933), .CP(clk), .Q(reg_iii_9[15]) );
  dff_sg \reg_ii_9_reg[14]  ( .D(n45285), .CP(clk), .Q(reg_ii_9[14]) );
  dff_sg \reg_iii_9_reg[14]  ( .D(n45273), .CP(clk), .Q(reg_iii_9[14]) );
  dff_sg \reg_ii_9_reg[13]  ( .D(n45286), .CP(clk), .Q(reg_ii_9[13]) );
  dff_sg \reg_iii_9_reg[13]  ( .D(n44915), .CP(clk), .Q(reg_iii_9[13]) );
  dff_sg \reg_ii_9_reg[12]  ( .D(n45251), .CP(clk), .Q(reg_ii_9[12]) );
  dff_sg \reg_iii_9_reg[12]  ( .D(n45142), .CP(clk), .Q(reg_iii_9[12]) );
  dff_sg \reg_ii_9_reg[11]  ( .D(n45252), .CP(clk), .Q(reg_ii_9[11]) );
  dff_sg \reg_iii_9_reg[11]  ( .D(n44445), .CP(clk), .Q(reg_iii_9[11]) );
  dff_sg \reg_ii_9_reg[10]  ( .D(n45249), .CP(clk), .Q(reg_ii_9[10]) );
  dff_sg \reg_iii_9_reg[10]  ( .D(n45139), .CP(clk), .Q(reg_iii_9[10]) );
  dff_sg \reg_ii_9_reg[9]  ( .D(n45250), .CP(clk), .Q(reg_ii_9[9]) );
  dff_sg \reg_iii_9_reg[9]  ( .D(n44535), .CP(clk), .Q(reg_iii_9[9]) );
  dff_sg \reg_ii_9_reg[8]  ( .D(n45256), .CP(clk), .Q(reg_ii_9[8]) );
  dff_sg \reg_iii_9_reg[8]  ( .D(n45290), .CP(clk), .Q(reg_iii_9[8]) );
  dff_sg \reg_ii_9_reg[7]  ( .D(n45257), .CP(clk), .Q(reg_ii_9[7]) );
  dff_sg \reg_iii_9_reg[7]  ( .D(n44444), .CP(clk), .Q(reg_iii_9[7]) );
  dff_sg \reg_ii_9_reg[6]  ( .D(n45253), .CP(clk), .Q(reg_ii_9[6]) );
  dff_sg \reg_iii_9_reg[6]  ( .D(n44280), .CP(clk), .Q(reg_iii_9[6]) );
  dff_sg \reg_ii_9_reg[5]  ( .D(n45254), .CP(clk), .Q(reg_ii_9[5]) );
  dff_sg \reg_iii_9_reg[5]  ( .D(n44446), .CP(clk), .Q(reg_iii_9[5]) );
  dff_sg \reg_ii_9_reg[4]  ( .D(n45242), .CP(clk), .Q(reg_ii_9[4]) );
  dff_sg \reg_iii_9_reg[4]  ( .D(n45292), .CP(clk), .Q(reg_iii_9[4]) );
  dff_sg \reg_ii_9_reg[3]  ( .D(n45243), .CP(clk), .Q(reg_ii_9[3]) );
  dff_sg \reg_iii_9_reg[3]  ( .D(n45293), .CP(clk), .Q(reg_iii_9[3]) );
  dff_sg \reg_ii_9_reg[2]  ( .D(n45240), .CP(clk), .Q(reg_ii_9[2]) );
  dff_sg \reg_iii_9_reg[2]  ( .D(n45282), .CP(clk), .Q(reg_iii_9[2]) );
  dff_sg \reg_ii_9_reg[1]  ( .D(n45241), .CP(clk), .Q(reg_ii_9[1]) );
  dff_sg \reg_iii_9_reg[1]  ( .D(n45283), .CP(clk), .Q(reg_iii_9[1]) );
  dff_sg \reg_ii_9_reg[0]  ( .D(n45246), .CP(clk), .Q(reg_ii_9[0]) );
  dff_sg \reg_iii_9_reg[0]  ( .D(n45280), .CP(clk), .Q(reg_iii_9[0]) );
  dff_sg \reg_ii_8_reg[19]  ( .D(n45524), .CP(clk), .Q(reg_ii_8[19]) );
  dff_sg \reg_iii_8_reg[19]  ( .D(n45247), .CP(clk), .Q(reg_iii_8[19]) );
  dff_sg \reg_ii_8_reg[18]  ( .D(n45153), .CP(clk), .Q(reg_ii_8[18]) );
  dff_sg \reg_iii_8_reg[18]  ( .D(n45244), .CP(clk), .Q(reg_iii_8[18]) );
  dff_sg \reg_ii_8_reg[17]  ( .D(n45154), .CP(clk), .Q(reg_ii_8[17]) );
  dff_sg \reg_iii_8_reg[17]  ( .D(n45245), .CP(clk), .Q(reg_iii_8[17]) );
  dff_sg \reg_ii_8_reg[16]  ( .D(n45515), .CP(clk), .Q(reg_ii_8[16]) );
  dff_sg \reg_iii_8_reg[16]  ( .D(n45268), .CP(clk), .Q(reg_iii_8[16]) );
  dff_sg \reg_ii_8_reg[15]  ( .D(n45516), .CP(clk), .Q(reg_ii_8[15]) );
  dff_sg \reg_iii_8_reg[15]  ( .D(n45269), .CP(clk), .Q(reg_iii_8[15]) );
  dff_sg \reg_ii_8_reg[14]  ( .D(n45340), .CP(clk), .Q(reg_ii_8[14]) );
  dff_sg \reg_iii_8_reg[14]  ( .D(n45266), .CP(clk), .Q(reg_iii_8[14]) );
  dff_sg \reg_ii_8_reg[13]  ( .D(n45341), .CP(clk), .Q(reg_ii_8[13]) );
  dff_sg \reg_iii_8_reg[13]  ( .D(n45267), .CP(clk), .Q(reg_iii_8[13]) );
  dff_sg \reg_ii_8_reg[12]  ( .D(n45525), .CP(clk), .Q(reg_ii_8[12]) );
  dff_sg \reg_iii_8_reg[12]  ( .D(n45270), .CP(clk), .Q(reg_iii_8[12]) );
  dff_sg \reg_ii_8_reg[11]  ( .D(n45526), .CP(clk), .Q(reg_ii_8[11]) );
  dff_sg \reg_iii_8_reg[11]  ( .D(n45271), .CP(clk), .Q(reg_iii_8[11]) );
  dff_sg \reg_ii_8_reg[10]  ( .D(n45491), .CP(clk), .Q(reg_ii_8[10]) );
  dff_sg \reg_iii_8_reg[10]  ( .D(n44441), .CP(clk), .Q(reg_iii_8[10]) );
  dff_sg \reg_ii_8_reg[9]  ( .D(n45225), .CP(clk), .Q(reg_ii_8[9]) );
  dff_sg \reg_iii_8_reg[9]  ( .D(n44526), .CP(clk), .Q(reg_iii_8[9]) );
  dff_sg \reg_ii_8_reg[8]  ( .D(n45158), .CP(clk), .Q(reg_ii_8[8]) );
  dff_sg \reg_iii_8_reg[8]  ( .D(n45260), .CP(clk), .Q(reg_iii_8[8]) );
  dff_sg \reg_ii_8_reg[7]  ( .D(n45159), .CP(clk), .Q(reg_ii_8[7]) );
  dff_sg \reg_iii_8_reg[7]  ( .D(n44605), .CP(clk), .Q(reg_iii_8[7]) );
  dff_sg \reg_ii_8_reg[6]  ( .D(n45156), .CP(clk), .Q(reg_ii_8[6]) );
  dff_sg \reg_iii_8_reg[6]  ( .D(n45258), .CP(clk), .Q(reg_iii_8[6]) );
  dff_sg \reg_ii_8_reg[5]  ( .D(n45157), .CP(clk), .Q(reg_ii_8[5]) );
  dff_sg \reg_iii_8_reg[5]  ( .D(n45259), .CP(clk), .Q(reg_iii_8[5]) );
  dff_sg \reg_ii_8_reg[4]  ( .D(n45166), .CP(clk), .Q(reg_ii_8[4]) );
  dff_sg \reg_iii_8_reg[4]  ( .D(n45264), .CP(clk), .Q(reg_iii_8[4]) );
  dff_sg \reg_ii_8_reg[3]  ( .D(n45167), .CP(clk), .Q(reg_ii_8[3]) );
  dff_sg \reg_iii_8_reg[3]  ( .D(n45265), .CP(clk), .Q(reg_iii_8[3]) );
  dff_sg \reg_ii_8_reg[2]  ( .D(n45163), .CP(clk), .Q(reg_ii_8[2]) );
  dff_sg \reg_iii_8_reg[2]  ( .D(n45262), .CP(clk), .Q(reg_iii_8[2]) );
  dff_sg \reg_ii_8_reg[1]  ( .D(n45164), .CP(clk), .Q(reg_ii_8[1]) );
  dff_sg \reg_iii_8_reg[1]  ( .D(n45263), .CP(clk), .Q(reg_iii_8[1]) );
  dff_sg \reg_ii_8_reg[0]  ( .D(n45169), .CP(clk), .Q(reg_ii_8[0]) );
  dff_sg \reg_iii_8_reg[0]  ( .D(n45523), .CP(clk), .Q(reg_iii_8[0]) );
  dff_sg \reg_ii_7_reg[19]  ( .D(n44364), .CP(clk), .Q(reg_ii_7[19]) );
  dff_sg \reg_iii_7_reg[19]  ( .D(n45170), .CP(clk), .Q(reg_iii_7[19]) );
  dff_sg \reg_ii_7_reg[18]  ( .D(n45151), .CP(clk), .Q(reg_ii_7[18]) );
  dff_sg \reg_iii_7_reg[18]  ( .D(n45168), .CP(clk), .Q(reg_iii_7[18]) );
  dff_sg \reg_ii_7_reg[17]  ( .D(n44410), .CP(clk), .Q(reg_ii_7[17]) );
  dff_sg \reg_iii_7_reg[17]  ( .D(n44389), .CP(clk), .Q(reg_iii_7[17]) );
  dff_sg \reg_ii_7_reg[16]  ( .D(n45255), .CP(clk), .Q(reg_ii_7[16]) );
  dff_sg \reg_iii_7_reg[16]  ( .D(n45161), .CP(clk), .Q(reg_iii_7[16]) );
  dff_sg \reg_ii_7_reg[15]  ( .D(n45272), .CP(clk), .Q(reg_ii_7[15]) );
  dff_sg \reg_iii_7_reg[15]  ( .D(n45327), .CP(clk), .Q(reg_iii_7[15]) );
  dff_sg \reg_ii_7_reg[14]  ( .D(n45150), .CP(clk), .Q(reg_ii_7[14]) );
  dff_sg \reg_iii_7_reg[14]  ( .D(n45160), .CP(clk), .Q(reg_iii_7[14]) );
  dff_sg \reg_ii_7_reg[13]  ( .D(n45284), .CP(clk), .Q(reg_ii_7[13]) );
  dff_sg \reg_iii_7_reg[13]  ( .D(n44386), .CP(clk), .Q(reg_iii_7[13]) );
  dff_sg \reg_ii_7_reg[12]  ( .D(n45494), .CP(clk), .Q(reg_ii_7[12]) );
  dff_sg \reg_iii_7_reg[12]  ( .D(n45518), .CP(clk), .Q(reg_iii_7[12]) );
  dff_sg \reg_ii_7_reg[11]  ( .D(n45490), .CP(clk), .Q(reg_ii_7[11]) );
  dff_sg \reg_iii_7_reg[11]  ( .D(n45519), .CP(clk), .Q(reg_iii_7[11]) );
  dff_sg \reg_ii_7_reg[10]  ( .D(n45493), .CP(clk), .Q(reg_ii_7[10]) );
  dff_sg \reg_iii_7_reg[10]  ( .D(n44403), .CP(clk), .Q(reg_iii_7[10]) );
  dff_sg \reg_ii_7_reg[9]  ( .D(n45499), .CP(clk), .Q(reg_ii_7[9]) );
  dff_sg \reg_iii_7_reg[9]  ( .D(n44358), .CP(clk), .Q(reg_iii_7[9]) );
  dff_sg \reg_ii_7_reg[8]  ( .D(n45472), .CP(clk), .Q(reg_ii_7[8]) );
  dff_sg \reg_iii_7_reg[8]  ( .D(n44822), .CP(clk), .Q(reg_iii_7[8]) );
  dff_sg \reg_ii_7_reg[7]  ( .D(n45473), .CP(clk), .Q(reg_ii_7[7]) );
  dff_sg \reg_iii_7_reg[7]  ( .D(n44819), .CP(clk), .Q(reg_iii_7[7]) );
  dff_sg \reg_ii_7_reg[6]  ( .D(n45485), .CP(clk), .Q(reg_ii_7[6]) );
  dff_sg \reg_iii_7_reg[6]  ( .D(n45504), .CP(clk), .Q(reg_iii_7[6]) );
  dff_sg \reg_ii_7_reg[5]  ( .D(n45486), .CP(clk), .Q(reg_ii_7[5]) );
  dff_sg \reg_iii_7_reg[5]  ( .D(n44306), .CP(clk), .Q(reg_iii_7[5]) );
  dff_sg \reg_ii_7_reg[4]  ( .D(n45322), .CP(clk), .Q(reg_ii_7[4]) );
  dff_sg \reg_iii_7_reg[4]  ( .D(n44810), .CP(clk), .Q(reg_iii_7[4]) );
  dff_sg \reg_ii_7_reg[3]  ( .D(n45319), .CP(clk), .Q(reg_ii_7[3]) );
  dff_sg \reg_iii_7_reg[3]  ( .D(n45492), .CP(clk), .Q(reg_iii_7[3]) );
  dff_sg \reg_ii_7_reg[2]  ( .D(n45522), .CP(clk), .Q(reg_ii_7[2]) );
  dff_sg \reg_iii_7_reg[2]  ( .D(n45248), .CP(clk), .Q(reg_iii_7[2]) );
  dff_sg \reg_ii_7_reg[1]  ( .D(n45311), .CP(clk), .Q(reg_ii_7[1]) );
  dff_sg \reg_iii_7_reg[1]  ( .D(n44319), .CP(clk), .Q(reg_iii_7[1]) );
  dff_sg \reg_ii_7_reg[0]  ( .D(n45291), .CP(clk), .Q(reg_ii_7[0]) );
  dff_sg \reg_iii_7_reg[0]  ( .D(n45503), .CP(clk), .Q(reg_iii_7[0]) );
  dff_sg \reg_ii_6_reg[19]  ( .D(n45548), .CP(clk), .Q(reg_ii_6[19]) );
  dff_sg \reg_iii_6_reg[19]  ( .D(n45297), .CP(clk), .Q(reg_iii_6[19]) );
  dff_sg \reg_ii_6_reg[18]  ( .D(n45546), .CP(clk), .Q(reg_ii_6[18]) );
  dff_sg \reg_iii_6_reg[18]  ( .D(n45308), .CP(clk), .Q(reg_iii_6[18]) );
  dff_sg \reg_ii_6_reg[17]  ( .D(n45547), .CP(clk), .Q(reg_ii_6[17]) );
  dff_sg \reg_iii_6_reg[17]  ( .D(n45314), .CP(clk), .Q(reg_iii_6[17]) );
  dff_sg \reg_ii_6_reg[16]  ( .D(n45550), .CP(clk), .Q(reg_ii_6[16]) );
  dff_sg \reg_iii_6_reg[16]  ( .D(n45538), .CP(clk), .Q(reg_iii_6[16]) );
  dff_sg \reg_ii_6_reg[15]  ( .D(n45551), .CP(clk), .Q(reg_ii_6[15]) );
  dff_sg \reg_iii_6_reg[15]  ( .D(n45539), .CP(clk), .Q(reg_iii_6[15]) );
  dff_sg \reg_ii_6_reg[14]  ( .D(n44923), .CP(clk), .Q(reg_ii_6[14]) );
  dff_sg \reg_iii_6_reg[14]  ( .D(n44837), .CP(clk), .Q(reg_iii_6[14]) );
  dff_sg \reg_ii_6_reg[13]  ( .D(n44922), .CP(clk), .Q(reg_ii_6[13]) );
  dff_sg \reg_iii_6_reg[13]  ( .D(n45537), .CP(clk), .Q(reg_iii_6[13]) );
  dff_sg \reg_ii_6_reg[12]  ( .D(n44926), .CP(clk), .Q(reg_ii_6[12]) );
  dff_sg \reg_iii_6_reg[12]  ( .D(n45543), .CP(clk), .Q(reg_iii_6[12]) );
  dff_sg \reg_ii_6_reg[11]  ( .D(n44925), .CP(clk), .Q(reg_ii_6[11]) );
  dff_sg \reg_iii_6_reg[11]  ( .D(n45544), .CP(clk), .Q(reg_iii_6[11]) );
  dff_sg \reg_ii_6_reg[10]  ( .D(n44917), .CP(clk), .Q(reg_ii_6[10]) );
  dff_sg \reg_iii_6_reg[10]  ( .D(n45541), .CP(clk), .Q(reg_iii_6[10]) );
  dff_sg \reg_ii_6_reg[9]  ( .D(n44916), .CP(clk), .Q(reg_ii_6[9]) );
  dff_sg \reg_iii_6_reg[9]  ( .D(n45542), .CP(clk), .Q(reg_iii_6[9]) );
  dff_sg \reg_ii_6_reg[8]  ( .D(n44920), .CP(clk), .Q(reg_ii_6[8]) );
  dff_sg \reg_iii_6_reg[8]  ( .D(n45531), .CP(clk), .Q(reg_iii_6[8]) );
  dff_sg \reg_ii_6_reg[7]  ( .D(n44919), .CP(clk), .Q(reg_ii_6[7]) );
  dff_sg \reg_iii_6_reg[7]  ( .D(n45532), .CP(clk), .Q(reg_iii_6[7]) );
  dff_sg \reg_ii_6_reg[6]  ( .D(n44935), .CP(clk), .Q(reg_ii_6[6]) );
  dff_sg \reg_iii_6_reg[6]  ( .D(n45528), .CP(clk), .Q(reg_iii_6[6]) );
  dff_sg \reg_ii_6_reg[5]  ( .D(n44934), .CP(clk), .Q(reg_ii_6[5]) );
  dff_sg \reg_iii_6_reg[5]  ( .D(n45529), .CP(clk), .Q(reg_iii_6[5]) );
  dff_sg \reg_ii_6_reg[4]  ( .D(n44938), .CP(clk), .Q(reg_ii_6[4]) );
  dff_sg \reg_iii_6_reg[4]  ( .D(n44825), .CP(clk), .Q(reg_iii_6[4]) );
  dff_sg \reg_ii_6_reg[3]  ( .D(n44937), .CP(clk), .Q(reg_ii_6[3]) );
  dff_sg \reg_iii_6_reg[3]  ( .D(n45536), .CP(clk), .Q(reg_iii_6[3]) );
  dff_sg \reg_ii_6_reg[2]  ( .D(n44929), .CP(clk), .Q(reg_ii_6[2]) );
  dff_sg \reg_iii_6_reg[2]  ( .D(n45534), .CP(clk), .Q(reg_iii_6[2]) );
  dff_sg \reg_ii_6_reg[1]  ( .D(n44928), .CP(clk), .Q(reg_ii_6[1]) );
  dff_sg \reg_iii_6_reg[1]  ( .D(n45535), .CP(clk), .Q(reg_iii_6[1]) );
  dff_sg \reg_ii_6_reg[0]  ( .D(n44932), .CP(clk), .Q(reg_ii_6[0]) );
  dff_sg \reg_iii_6_reg[0]  ( .D(n44828), .CP(clk), .Q(reg_iii_6[0]) );
  dff_sg \reg_ii_5_reg[19]  ( .D(n44973), .CP(clk), .Q(reg_ii_5[19]) );
  dff_sg \reg_iii_5_reg[19]  ( .D(n44931), .CP(clk), .Q(reg_iii_5[19]) );
  dff_sg \reg_ii_5_reg[18]  ( .D(n44965), .CP(clk), .Q(reg_ii_5[18]) );
  dff_sg \reg_iii_5_reg[18]  ( .D(n44899), .CP(clk), .Q(reg_iii_5[18]) );
  dff_sg \reg_ii_5_reg[17]  ( .D(n44964), .CP(clk), .Q(reg_ii_5[17]) );
  dff_sg \reg_iii_5_reg[17]  ( .D(n44898), .CP(clk), .Q(reg_iii_5[17]) );
  dff_sg \reg_ii_5_reg[16]  ( .D(n44968), .CP(clk), .Q(reg_ii_5[16]) );
  dff_sg \reg_iii_5_reg[16]  ( .D(n44902), .CP(clk), .Q(reg_iii_5[16]) );
  dff_sg \reg_ii_5_reg[15]  ( .D(n44967), .CP(clk), .Q(reg_ii_5[15]) );
  dff_sg \reg_iii_5_reg[15]  ( .D(n44901), .CP(clk), .Q(reg_iii_5[15]) );
  dff_sg \reg_ii_5_reg[14]  ( .D(n44983), .CP(clk), .Q(reg_ii_5[14]) );
  dff_sg \reg_iii_5_reg[14]  ( .D(n44893), .CP(clk), .Q(reg_iii_5[14]) );
  dff_sg \reg_ii_5_reg[13]  ( .D(n44982), .CP(clk), .Q(reg_ii_5[13]) );
  dff_sg \reg_iii_5_reg[13]  ( .D(n44892), .CP(clk), .Q(reg_iii_5[13]) );
  dff_sg \reg_ii_5_reg[12]  ( .D(n44986), .CP(clk), .Q(reg_ii_5[12]) );
  dff_sg \reg_iii_5_reg[12]  ( .D(n44896), .CP(clk), .Q(reg_iii_5[12]) );
  dff_sg \reg_ii_5_reg[11]  ( .D(n44985), .CP(clk), .Q(reg_ii_5[11]) );
  dff_sg \reg_iii_5_reg[11]  ( .D(n44895), .CP(clk), .Q(reg_iii_5[11]) );
  dff_sg \reg_ii_5_reg[10]  ( .D(n44977), .CP(clk), .Q(reg_ii_5[10]) );
  dff_sg \reg_iii_5_reg[10]  ( .D(n44911), .CP(clk), .Q(reg_iii_5[10]) );
  dff_sg \reg_ii_5_reg[9]  ( .D(n44976), .CP(clk), .Q(reg_ii_5[9]) );
  dff_sg \reg_iii_5_reg[9]  ( .D(n44910), .CP(clk), .Q(reg_iii_5[9]) );
  dff_sg \reg_ii_5_reg[8]  ( .D(n44980), .CP(clk), .Q(reg_ii_5[8]) );
  dff_sg \reg_iii_5_reg[8]  ( .D(n44914), .CP(clk), .Q(reg_iii_5[8]) );
  dff_sg \reg_ii_5_reg[7]  ( .D(n44979), .CP(clk), .Q(reg_ii_5[7]) );
  dff_sg \reg_iii_5_reg[7]  ( .D(n44913), .CP(clk), .Q(reg_iii_5[7]) );
  dff_sg \reg_ii_5_reg[6]  ( .D(n44947), .CP(clk), .Q(reg_ii_5[6]) );
  dff_sg \reg_iii_5_reg[6]  ( .D(n44905), .CP(clk), .Q(reg_iii_5[6]) );
  dff_sg \reg_ii_5_reg[5]  ( .D(n44946), .CP(clk), .Q(reg_ii_5[5]) );
  dff_sg \reg_iii_5_reg[5]  ( .D(n44904), .CP(clk), .Q(reg_iii_5[5]) );
  dff_sg \reg_ii_5_reg[4]  ( .D(n44950), .CP(clk), .Q(reg_ii_5[4]) );
  dff_sg \reg_iii_5_reg[4]  ( .D(n44908), .CP(clk), .Q(reg_iii_5[4]) );
  dff_sg \reg_ii_5_reg[3]  ( .D(n44949), .CP(clk), .Q(reg_ii_5[3]) );
  dff_sg \reg_iii_5_reg[3]  ( .D(n44907), .CP(clk), .Q(reg_iii_5[3]) );
  dff_sg \reg_ii_5_reg[2]  ( .D(n44941), .CP(clk), .Q(reg_ii_5[2]) );
  dff_sg \reg_iii_5_reg[2]  ( .D(n44971), .CP(clk), .Q(reg_iii_5[2]) );
  dff_sg \reg_ii_5_reg[1]  ( .D(n44940), .CP(clk), .Q(reg_ii_5[1]) );
  dff_sg \reg_iii_5_reg[1]  ( .D(n44970), .CP(clk), .Q(reg_iii_5[1]) );
  dff_sg \reg_ii_5_reg[0]  ( .D(n44944), .CP(clk), .Q(reg_ii_5[0]) );
  dff_sg \reg_iii_5_reg[0]  ( .D(n44974), .CP(clk), .Q(reg_iii_5[0]) );
  dff_sg \reg_ii_4_reg[19]  ( .D(n44943), .CP(clk), .Q(reg_ii_4[19]) );
  dff_sg \reg_iii_4_reg[19]  ( .D(n45152), .CP(clk), .Q(reg_iii_4[19]) );
  dff_sg \reg_ii_14_reg[16]  ( .D(n44833), .CP(clk), .Q(reg_ii_14[16]) );
  dff_sg \reg_iii_14_reg[16]  ( .D(n44961), .CP(clk), .Q(reg_iii_14[16]) );
  dff_sg \reg_ii_14_reg[15]  ( .D(n44832), .CP(clk), .Q(reg_ii_14[15]) );
  dff_sg \reg_iii_14_reg[15]  ( .D(n44953), .CP(clk), .Q(reg_iii_14[15]) );
  dff_sg \reg_ii_14_reg[14]  ( .D(n44836), .CP(clk), .Q(reg_ii_14[14]) );
  dff_sg \reg_iii_14_reg[14]  ( .D(n44952), .CP(clk), .Q(reg_iii_14[14]) );
  dff_sg \reg_ii_14_reg[13]  ( .D(n44835), .CP(clk), .Q(reg_ii_14[13]) );
  dff_sg \reg_iii_14_reg[13]  ( .D(n44956), .CP(clk), .Q(reg_iii_14[13]) );
  dff_sg \reg_ii_14_reg[12]  ( .D(n44803), .CP(clk), .Q(reg_ii_14[12]) );
  dff_sg \reg_iii_14_reg[12]  ( .D(n44955), .CP(clk), .Q(reg_iii_14[12]) );
  dff_sg \reg_ii_14_reg[11]  ( .D(n44802), .CP(clk), .Q(reg_ii_14[11]) );
  dff_sg \reg_iii_14_reg[11]  ( .D(n44827), .CP(clk), .Q(reg_iii_14[11]) );
  dff_sg \reg_ii_14_reg[10]  ( .D(n44806), .CP(clk), .Q(reg_ii_14[10]) );
  dff_sg \reg_iii_14_reg[10]  ( .D(n44826), .CP(clk), .Q(reg_iii_14[10]) );
  dff_sg \reg_ii_14_reg[9]  ( .D(n44805), .CP(clk), .Q(reg_ii_14[9]) );
  dff_sg \reg_iii_14_reg[9]  ( .D(n44830), .CP(clk), .Q(reg_iii_14[9]) );
  dff_sg \reg_ii_14_reg[8]  ( .D(n44797), .CP(clk), .Q(reg_ii_14[8]) );
  dff_sg \reg_iii_14_reg[8]  ( .D(n44829), .CP(clk), .Q(reg_iii_14[8]) );
  dff_sg \reg_ii_14_reg[7]  ( .D(n44796), .CP(clk), .Q(reg_ii_14[7]) );
  dff_sg \reg_iii_14_reg[7]  ( .D(n44821), .CP(clk), .Q(reg_iii_14[7]) );
  dff_sg \reg_ii_14_reg[6]  ( .D(n44800), .CP(clk), .Q(reg_ii_14[6]) );
  dff_sg \reg_iii_14_reg[6]  ( .D(n44820), .CP(clk), .Q(reg_iii_14[6]) );
  dff_sg \reg_ii_14_reg[5]  ( .D(n44799), .CP(clk), .Q(reg_ii_14[5]) );
  dff_sg \reg_iii_14_reg[5]  ( .D(n44824), .CP(clk), .Q(reg_iii_14[5]) );
  dff_sg \reg_ii_14_reg[4]  ( .D(n44815), .CP(clk), .Q(reg_ii_14[4]) );
  dff_sg \reg_iii_14_reg[4]  ( .D(n44823), .CP(clk), .Q(reg_iii_14[4]) );
  dff_sg \reg_ii_14_reg[3]  ( .D(n44814), .CP(clk), .Q(reg_ii_14[3]) );
  dff_sg \reg_iii_14_reg[3]  ( .D(n44839), .CP(clk), .Q(reg_iii_14[3]) );
  dff_sg \reg_ii_14_reg[2]  ( .D(n44818), .CP(clk), .Q(reg_ii_14[2]) );
  dff_sg \reg_iii_14_reg[2]  ( .D(n44838), .CP(clk), .Q(reg_iii_14[2]) );
  dff_sg \reg_ii_14_reg[1]  ( .D(n44817), .CP(clk), .Q(reg_ii_14[1]) );
  dff_sg \reg_iii_14_reg[1]  ( .D(n44842), .CP(clk), .Q(reg_iii_14[1]) );
  dff_sg \reg_ii_14_reg[0]  ( .D(n44809), .CP(clk), .Q(reg_ii_14[0]) );
  dff_sg \reg_iii_14_reg[0]  ( .D(n44841), .CP(clk), .Q(reg_iii_14[0]) );
  dff_sg \reg_ii_13_reg[19]  ( .D(n44850), .CP(clk), .Q(reg_ii_13[19]) );
  dff_sg \reg_iii_13_reg[19]  ( .D(n44808), .CP(clk), .Q(reg_iii_13[19]) );
  dff_sg \reg_ii_13_reg[18]  ( .D(n44854), .CP(clk), .Q(reg_ii_13[18]) );
  dff_sg \reg_iii_13_reg[18]  ( .D(n44812), .CP(clk), .Q(reg_iii_13[18]) );
  dff_sg \reg_ii_13_reg[17]  ( .D(n44853), .CP(clk), .Q(reg_ii_13[17]) );
  dff_sg \reg_iii_13_reg[17]  ( .D(n44811), .CP(clk), .Q(reg_iii_13[17]) );
  dff_sg \reg_ii_13_reg[16]  ( .D(n44845), .CP(clk), .Q(reg_ii_13[16]) );
  dff_sg \reg_iii_13_reg[16]  ( .D(n44875), .CP(clk), .Q(reg_iii_13[16]) );
  dff_sg \reg_ii_13_reg[15]  ( .D(n44844), .CP(clk), .Q(reg_ii_13[15]) );
  dff_sg \reg_iii_13_reg[15]  ( .D(n44874), .CP(clk), .Q(reg_iii_13[15]) );
  dff_sg \reg_ii_13_reg[14]  ( .D(n44848), .CP(clk), .Q(reg_ii_13[14]) );
  dff_sg \reg_iii_13_reg[14]  ( .D(n44878), .CP(clk), .Q(reg_iii_13[14]) );
  dff_sg \reg_ii_13_reg[13]  ( .D(n44847), .CP(clk), .Q(reg_ii_13[13]) );
  dff_sg \reg_iii_13_reg[13]  ( .D(n44877), .CP(clk), .Q(reg_iii_13[13]) );
  dff_sg \reg_ii_13_reg[12]  ( .D(n44863), .CP(clk), .Q(reg_ii_13[12]) );
  dff_sg \reg_iii_13_reg[12]  ( .D(n44869), .CP(clk), .Q(reg_iii_13[12]) );
  dff_sg \reg_ii_13_reg[11]  ( .D(n44862), .CP(clk), .Q(reg_ii_13[11]) );
  dff_sg \reg_iii_13_reg[11]  ( .D(n44868), .CP(clk), .Q(reg_iii_13[11]) );
  dff_sg \reg_ii_13_reg[10]  ( .D(n44866), .CP(clk), .Q(reg_ii_13[10]) );
  dff_sg \reg_iii_13_reg[10]  ( .D(n44872), .CP(clk), .Q(reg_iii_13[10]) );
  dff_sg \reg_ii_13_reg[9]  ( .D(n44865), .CP(clk), .Q(reg_ii_13[9]) );
  dff_sg \reg_iii_13_reg[9]  ( .D(n44871), .CP(clk), .Q(reg_iii_13[9]) );
  dff_sg \reg_ii_13_reg[8]  ( .D(n44857), .CP(clk), .Q(reg_ii_13[8]) );
  dff_sg \reg_iii_13_reg[8]  ( .D(n44887), .CP(clk), .Q(reg_iii_13[8]) );
  dff_sg \reg_ii_13_reg[7]  ( .D(n44856), .CP(clk), .Q(reg_ii_13[7]) );
  dff_sg \reg_iii_13_reg[7]  ( .D(n44886), .CP(clk), .Q(reg_iii_13[7]) );
  dff_sg \reg_ii_13_reg[6]  ( .D(n44860), .CP(clk), .Q(reg_ii_13[6]) );
  dff_sg \reg_iii_13_reg[6]  ( .D(n44890), .CP(clk), .Q(reg_iii_13[6]) );
  dff_sg \reg_ii_13_reg[5]  ( .D(n44859), .CP(clk), .Q(reg_ii_13[5]) );
  dff_sg \reg_iii_13_reg[5]  ( .D(n44889), .CP(clk), .Q(reg_iii_13[5]) );
  dff_sg \reg_ii_13_reg[4]  ( .D(n44504), .CP(clk), .Q(reg_ii_13[4]) );
  dff_sg \reg_iii_13_reg[4]  ( .D(n44881), .CP(clk), .Q(reg_iii_13[4]) );
  dff_sg \reg_ii_13_reg[3]  ( .D(n44503), .CP(clk), .Q(reg_ii_13[3]) );
  dff_sg \reg_iii_13_reg[3]  ( .D(n44880), .CP(clk), .Q(reg_iii_13[3]) );
  dff_sg \reg_ii_13_reg[2]  ( .D(n44507), .CP(clk), .Q(reg_ii_13[2]) );
  dff_sg \reg_iii_13_reg[2]  ( .D(n44884), .CP(clk), .Q(reg_iii_13[2]) );
  dff_sg \reg_ii_13_reg[1]  ( .D(n44506), .CP(clk), .Q(reg_ii_13[1]) );
  dff_sg \reg_iii_13_reg[1]  ( .D(n44883), .CP(clk), .Q(reg_iii_13[1]) );
  dff_sg \reg_ii_13_reg[0]  ( .D(n44505), .CP(clk), .Q(reg_ii_13[0]) );
  dff_sg \reg_iii_13_reg[0]  ( .D(n44851), .CP(clk), .Q(reg_iii_13[0]) );
  dff_sg \reg_ii_12_reg[19]  ( .D(n44496), .CP(clk), .Q(reg_ii_12[19]) );
  dff_sg \reg_iii_12_reg[19]  ( .D(n44502), .CP(clk), .Q(reg_iii_12[19]) );
  dff_sg \reg_ii_12_reg[18]  ( .D(n44500), .CP(clk), .Q(reg_ii_12[18]) );
  dff_sg \reg_iii_12_reg[18]  ( .D(n44495), .CP(clk), .Q(reg_iii_12[18]) );
  dff_sg \reg_ii_12_reg[17]  ( .D(n44499), .CP(clk), .Q(reg_ii_12[17]) );
  dff_sg \reg_iii_12_reg[17]  ( .D(n44501), .CP(clk), .Q(reg_iii_12[17]) );
  dff_sg \reg_ii_12_reg[16]  ( .D(n44483), .CP(clk), .Q(reg_ii_12[16]) );
  dff_sg \reg_iii_12_reg[16]  ( .D(n44519), .CP(clk), .Q(reg_iii_12[16]) );
  dff_sg \reg_ii_12_reg[15]  ( .D(n44492), .CP(clk), .Q(reg_ii_12[15]) );
  dff_sg \reg_iii_12_reg[15]  ( .D(n44518), .CP(clk), .Q(reg_iii_12[15]) );
  dff_sg \reg_ii_12_reg[14]  ( .D(n44494), .CP(clk), .Q(reg_ii_12[14]) );
  dff_sg \reg_iii_12_reg[14]  ( .D(n44508), .CP(clk), .Q(reg_iii_12[14]) );
  dff_sg \reg_ii_12_reg[13]  ( .D(n44493), .CP(clk), .Q(reg_ii_12[13]) );
  dff_sg \reg_iii_12_reg[13]  ( .D(n44517), .CP(clk), .Q(reg_iii_12[13]) );
  dff_sg \reg_ii_12_reg[12]  ( .D(n45091), .CP(clk), .Q(reg_ii_12[12]) );
  dff_sg \reg_iii_12_reg[12]  ( .D(n44510), .CP(clk), .Q(reg_iii_12[12]) );
  dff_sg \reg_ii_12_reg[11]  ( .D(n45090), .CP(clk), .Q(reg_ii_12[11]) );
  dff_sg \reg_iii_12_reg[11]  ( .D(n44509), .CP(clk), .Q(reg_iii_12[11]) );
  dff_sg \reg_ii_12_reg[10]  ( .D(n45094), .CP(clk), .Q(reg_ii_12[10]) );
  dff_sg \reg_iii_12_reg[10]  ( .D(n44513), .CP(clk), .Q(reg_iii_12[10]) );
  dff_sg \reg_ii_12_reg[9]  ( .D(n45093), .CP(clk), .Q(reg_ii_12[9]) );
  dff_sg \reg_iii_12_reg[9]  ( .D(n44512), .CP(clk), .Q(reg_iii_12[9]) );
  dff_sg \reg_ii_12_reg[8]  ( .D(n45082), .CP(clk), .Q(reg_ii_12[8]) );
  dff_sg \reg_iii_12_reg[8]  ( .D(n44491), .CP(clk), .Q(reg_iii_12[8]) );
  dff_sg \reg_ii_12_reg[7]  ( .D(n45088), .CP(clk), .Q(reg_ii_12[7]) );
  dff_sg \reg_iii_12_reg[7]  ( .D(n44490), .CP(clk), .Q(reg_iii_12[7]) );
  dff_sg \reg_ii_12_reg[6]  ( .D(n45079), .CP(clk), .Q(reg_ii_12[6]) );
  dff_sg \reg_iii_12_reg[6]  ( .D(n44486), .CP(clk), .Q(reg_iii_12[6]) );
  dff_sg \reg_ii_12_reg[5]  ( .D(n45085), .CP(clk), .Q(reg_ii_12[5]) );
  dff_sg \reg_iii_12_reg[5]  ( .D(n44489), .CP(clk), .Q(reg_iii_12[5]) );
  dff_sg \reg_ii_12_reg[4]  ( .D(n45096), .CP(clk), .Q(reg_ii_12[4]) );
  dff_sg \reg_iii_12_reg[4]  ( .D(n44485), .CP(clk), .Q(reg_iii_12[4]) );
  dff_sg \reg_ii_12_reg[3]  ( .D(n45095), .CP(clk), .Q(reg_ii_12[3]) );
  dff_sg \reg_iii_12_reg[3]  ( .D(n44484), .CP(clk), .Q(reg_iii_12[3]) );
  dff_sg \reg_ii_12_reg[2]  ( .D(n45089), .CP(clk), .Q(reg_ii_12[2]) );
  dff_sg \reg_iii_12_reg[2]  ( .D(n44488), .CP(clk), .Q(reg_iii_12[2]) );
  dff_sg \reg_ii_12_reg[1]  ( .D(n45092), .CP(clk), .Q(reg_ii_12[1]) );
  dff_sg \reg_iii_12_reg[1]  ( .D(n44487), .CP(clk), .Q(reg_iii_12[1]) );
  dff_sg \reg_ii_12_reg[0]  ( .D(n45098), .CP(clk), .Q(reg_ii_12[0]) );
  dff_sg \reg_iii_12_reg[0]  ( .D(n44497), .CP(clk), .Q(reg_iii_12[0]) );
  dff_sg \reg_ii_11_reg[19]  ( .D(n45029), .CP(clk), .Q(reg_ii_11[19]) );
  dff_sg \reg_iii_11_reg[19]  ( .D(n45097), .CP(clk), .Q(reg_iii_11[19]) );
  dff_sg \reg_ii_11_reg[18]  ( .D(n45015), .CP(clk), .Q(reg_ii_11[18]) );
  dff_sg \reg_iii_11_reg[18]  ( .D(n45100), .CP(clk), .Q(reg_iii_11[18]) );
  dff_sg \reg_ii_11_reg[17]  ( .D(n45028), .CP(clk), .Q(reg_ii_11[17]) );
  dff_sg \reg_iii_11_reg[17]  ( .D(n45099), .CP(clk), .Q(reg_iii_11[17]) );
  dff_sg \reg_ii_11_reg[16]  ( .D(n45014), .CP(clk), .Q(reg_ii_11[16]) );
  dff_sg \reg_iii_11_reg[16]  ( .D(n44511), .CP(clk), .Q(reg_iii_11[16]) );
  dff_sg \reg_ii_11_reg[15]  ( .D(n45013), .CP(clk), .Q(reg_ii_11[15]) );
  dff_sg \reg_iii_11_reg[15]  ( .D(n45070), .CP(clk), .Q(reg_iii_11[15]) );
  dff_sg \reg_ii_11_reg[14]  ( .D(n45017), .CP(clk), .Q(reg_ii_11[14]) );
  dff_sg \reg_iii_11_reg[14]  ( .D(n44514), .CP(clk), .Q(reg_iii_11[14]) );
  dff_sg \reg_ii_11_reg[13]  ( .D(n45016), .CP(clk), .Q(reg_ii_11[13]) );
  dff_sg \reg_iii_11_reg[13]  ( .D(n45076), .CP(clk), .Q(reg_iii_11[13]) );
  dff_sg \reg_ii_11_reg[12]  ( .D(n45032), .CP(clk), .Q(reg_ii_11[12]) );
  dff_sg \reg_iii_11_reg[12]  ( .D(n44516), .CP(clk), .Q(reg_iii_11[12]) );
  dff_sg \reg_ii_11_reg[11]  ( .D(n45031), .CP(clk), .Q(reg_ii_11[11]) );
  dff_sg \reg_iii_11_reg[11]  ( .D(n44515), .CP(clk), .Q(reg_iii_11[11]) );
  dff_sg \reg_ii_11_reg[10]  ( .D(n45038), .CP(clk), .Q(reg_ii_11[10]) );
  dff_sg \reg_iii_11_reg[10]  ( .D(n45072), .CP(clk), .Q(reg_iii_11[10]) );
  dff_sg \reg_ii_11_reg[9]  ( .D(n45035), .CP(clk), .Q(reg_ii_11[9]) );
  dff_sg \reg_iii_11_reg[9]  ( .D(n45071), .CP(clk), .Q(reg_iii_11[9]) );
  dff_sg \reg_ii_11_reg[8]  ( .D(n45034), .CP(clk), .Q(reg_ii_11[8]) );
  dff_sg \reg_iii_11_reg[8]  ( .D(n45084), .CP(clk), .Q(reg_iii_11[8]) );
  dff_sg \reg_ii_11_reg[7]  ( .D(n45033), .CP(clk), .Q(reg_ii_11[7]) );
  dff_sg \reg_iii_11_reg[7]  ( .D(n45083), .CP(clk), .Q(reg_iii_11[7]) );
  dff_sg \reg_ii_11_reg[6]  ( .D(n45037), .CP(clk), .Q(reg_ii_11[6]) );
  dff_sg \reg_iii_11_reg[6]  ( .D(n45087), .CP(clk), .Q(reg_iii_11[6]) );
  dff_sg \reg_ii_11_reg[5]  ( .D(n45036), .CP(clk), .Q(reg_ii_11[5]) );
  dff_sg \reg_iii_11_reg[5]  ( .D(n45086), .CP(clk), .Q(reg_iii_11[5]) );
  dff_sg \reg_ii_11_reg[4]  ( .D(n44996), .CP(clk), .Q(reg_ii_11[4]) );
  dff_sg \reg_iii_11_reg[4]  ( .D(n45078), .CP(clk), .Q(reg_iii_11[4]) );
  dff_sg \reg_ii_11_reg[3]  ( .D(n44995), .CP(clk), .Q(reg_ii_11[3]) );
  dff_sg \reg_iii_11_reg[3]  ( .D(n45077), .CP(clk), .Q(reg_iii_11[3]) );
  dff_sg \reg_ii_11_reg[2]  ( .D(n44999), .CP(clk), .Q(reg_ii_11[2]) );
  dff_sg \reg_iii_11_reg[2]  ( .D(n45081), .CP(clk), .Q(reg_iii_11[2]) );
  dff_sg \reg_ii_11_reg[1]  ( .D(n44998), .CP(clk), .Q(reg_ii_11[1]) );
  dff_sg \reg_iii_11_reg[1]  ( .D(n45080), .CP(clk), .Q(reg_iii_11[1]) );
  dff_sg \reg_ii_11_reg[0]  ( .D(n44990), .CP(clk), .Q(reg_ii_11[0]) );
  dff_sg \reg_iii_11_reg[0]  ( .D(n45030), .CP(clk), .Q(reg_iii_11[0]) );
  dff_sg \reg_ii_10_reg[19]  ( .D(n45067), .CP(clk), .Q(reg_ii_10[19]) );
  dff_sg \reg_iii_10_reg[19]  ( .D(n44989), .CP(clk), .Q(reg_iii_10[19]) );
  dff_sg \reg_ii_10_reg[18]  ( .D(n45064), .CP(clk), .Q(reg_ii_10[18]) );
  dff_sg \reg_iii_10_reg[18]  ( .D(n44993), .CP(clk), .Q(reg_iii_10[18]) );
  dff_sg \reg_ii_10_reg[17]  ( .D(n45057), .CP(clk), .Q(reg_ii_10[17]) );
  dff_sg \reg_iii_10_reg[17]  ( .D(n44992), .CP(clk), .Q(reg_iii_10[17]) );
  dff_sg \reg_ii_10_reg[16]  ( .D(n45066), .CP(clk), .Q(reg_ii_10[16]) );
  dff_sg \reg_iii_10_reg[16]  ( .D(n45008), .CP(clk), .Q(reg_iii_10[16]) );
  dff_sg \reg_ii_10_reg[15]  ( .D(n45065), .CP(clk), .Q(reg_ii_10[15]) );
  dff_sg \reg_iii_10_reg[15]  ( .D(n45007), .CP(clk), .Q(reg_iii_10[15]) );
  dff_sg \reg_ii_10_reg[14]  ( .D(n45069), .CP(clk), .Q(reg_ii_10[14]) );
  dff_sg \reg_iii_10_reg[14]  ( .D(n45011), .CP(clk), .Q(reg_iii_10[14]) );
  dff_sg \reg_ii_10_reg[13]  ( .D(n45068), .CP(clk), .Q(reg_ii_10[13]) );
  dff_sg \reg_iii_10_reg[13]  ( .D(n45010), .CP(clk), .Q(reg_iii_10[13]) );
  dff_sg \reg_ii_10_reg[12]  ( .D(n45046), .CP(clk), .Q(reg_ii_10[12]) );
  dff_sg \reg_iii_10_reg[12]  ( .D(n45002), .CP(clk), .Q(reg_iii_10[12]) );
  dff_sg \reg_ii_10_reg[11]  ( .D(n45045), .CP(clk), .Q(reg_ii_10[11]) );
  dff_sg \reg_iii_10_reg[11]  ( .D(n45001), .CP(clk), .Q(reg_iii_10[11]) );
  dff_sg \reg_ii_10_reg[10]  ( .D(n45049), .CP(clk), .Q(reg_ii_10[10]) );
  dff_sg \reg_iii_10_reg[10]  ( .D(n45005), .CP(clk), .Q(reg_iii_10[10]) );
  dff_sg \reg_ii_10_reg[9]  ( .D(n45048), .CP(clk), .Q(reg_ii_10[9]) );
  dff_sg \reg_iii_10_reg[9]  ( .D(n45004), .CP(clk), .Q(reg_iii_10[9]) );
  dff_sg \reg_ii_10_reg[8]  ( .D(n45040), .CP(clk), .Q(reg_ii_10[8]) );
  dff_sg \reg_iii_10_reg[8]  ( .D(n45063), .CP(clk), .Q(reg_iii_10[8]) );
  dff_sg \reg_ii_10_reg[7]  ( .D(n45039), .CP(clk), .Q(reg_ii_10[7]) );
  dff_sg \reg_iii_10_reg[7]  ( .D(n45062), .CP(clk), .Q(reg_iii_10[7]) );
  dff_sg \reg_ii_10_reg[6]  ( .D(n45043), .CP(clk), .Q(reg_ii_10[6]) );
  dff_sg \reg_iii_10_reg[6]  ( .D(n45058), .CP(clk), .Q(reg_iii_10[6]) );
  dff_sg \reg_ii_10_reg[5]  ( .D(n45042), .CP(clk), .Q(reg_ii_10[5]) );
  dff_sg \reg_iii_10_reg[5]  ( .D(n45061), .CP(clk), .Q(reg_iii_10[5]) );
  dff_sg \reg_ii_10_reg[4]  ( .D(n45053), .CP(clk), .Q(reg_ii_10[4]) );
  dff_sg \reg_iii_10_reg[4]  ( .D(n45047), .CP(clk), .Q(reg_iii_10[4]) );
  dff_sg \reg_ii_10_reg[3]  ( .D(n45052), .CP(clk), .Q(reg_ii_10[3]) );
  dff_sg \reg_iii_10_reg[3]  ( .D(n45044), .CP(clk), .Q(reg_iii_10[3]) );
  dff_sg \reg_ii_10_reg[2]  ( .D(n45056), .CP(clk), .Q(reg_ii_10[2]) );
  dff_sg \reg_iii_10_reg[2]  ( .D(n45060), .CP(clk), .Q(reg_iii_10[2]) );
  dff_sg \reg_ii_10_reg[1]  ( .D(n45055), .CP(clk), .Q(reg_ii_10[1]) );
  dff_sg \reg_iii_10_reg[1]  ( .D(n45059), .CP(clk), .Q(reg_iii_10[1]) );
  dff_sg \reg_ii_10_reg[0]  ( .D(n45054), .CP(clk), .Q(reg_ii_10[0]) );
  dff_sg \reg_iii_10_reg[0]  ( .D(n44987), .CP(clk), .Q(reg_iii_10[0]) );
  dff_sg \reg_ii_9_reg[19]  ( .D(n45051), .CP(clk), .Q(reg_ii_9[19]) );
  dff_sg \reg_iii_9_reg[19]  ( .D(n44529), .CP(clk), .Q(reg_iii_9[19]) );
  dff_sg \reg_ii_9_reg[18]  ( .D(n45041), .CP(clk), .Q(reg_ii_9[18]) );
  dff_sg \reg_iii_9_reg[18]  ( .D(n44864), .CP(clk), .Q(reg_iii_9[18]) );
  dff_sg \reg_ww_3_reg[15]  ( .D(n44978), .CP(clk), .Q(reg_ww_3[15]) );
  dff_sg \reg_www_3_reg[15]  ( .D(n44867), .CP(clk), .Q(reg_www_3[15]) );
  dff_sg \reg_ww_3_reg[14]  ( .D(n44997), .CP(clk), .Q(reg_ww_3[14]) );
  dff_sg \reg_www_3_reg[14]  ( .D(n44897), .CP(clk), .Q(reg_www_3[14]) );
  dff_sg \reg_ww_3_reg[13]  ( .D(n44994), .CP(clk), .Q(reg_ww_3[13]) );
  dff_sg \reg_www_3_reg[13]  ( .D(n44894), .CP(clk), .Q(reg_www_3[13]) );
  dff_sg \reg_ww_3_reg[12]  ( .D(n44939), .CP(clk), .Q(reg_ww_3[12]) );
  dff_sg \reg_www_3_reg[12]  ( .D(n44888), .CP(clk), .Q(reg_www_3[12]) );
  dff_sg \reg_ww_3_reg[11]  ( .D(n44936), .CP(clk), .Q(reg_ww_3[11]) );
  dff_sg \reg_www_3_reg[11]  ( .D(n44885), .CP(clk), .Q(reg_www_3[11]) );
  dff_sg \reg_ww_3_reg[10]  ( .D(n44951), .CP(clk), .Q(reg_ww_3[10]) );
  dff_sg \reg_www_3_reg[10]  ( .D(n44969), .CP(clk), .Q(reg_www_3[10]) );
  dff_sg \reg_ww_3_reg[9]  ( .D(n44912), .CP(clk), .Q(reg_ww_3[9]) );
  dff_sg \reg_www_3_reg[9]  ( .D(n44960), .CP(clk), .Q(reg_www_3[9]) );
  dff_sg \reg_ww_3_reg[8]  ( .D(n44906), .CP(clk), .Q(reg_ww_3[8]) );
  dff_sg \reg_www_3_reg[8]  ( .D(n44957), .CP(clk), .Q(reg_www_3[8]) );
  dff_sg \reg_ww_3_reg[7]  ( .D(n44903), .CP(clk), .Q(reg_ww_3[7]) );
  dff_sg \reg_www_3_reg[7]  ( .D(n44954), .CP(clk), .Q(reg_www_3[7]) );
  dff_sg \reg_ww_3_reg[6]  ( .D(n44972), .CP(clk), .Q(reg_ww_3[6]) );
  dff_sg \reg_www_3_reg[6]  ( .D(n44617), .CP(clk), .Q(reg_www_3[6]) );
  dff_sg \reg_ww_3_reg[5]  ( .D(n44966), .CP(clk), .Q(reg_ww_3[5]) );
  dff_sg \reg_www_3_reg[5]  ( .D(n44616), .CP(clk), .Q(reg_www_3[5]) );
  dff_sg \reg_ww_3_reg[4]  ( .D(n44948), .CP(clk), .Q(reg_ww_3[4]) );
  dff_sg \reg_www_3_reg[4]  ( .D(n45003), .CP(clk), .Q(reg_www_3[4]) );
  dff_sg \reg_ww_3_reg[3]  ( .D(n44945), .CP(clk), .Q(reg_ww_3[3]) );
  dff_sg \reg_www_3_reg[3]  ( .D(n45000), .CP(clk), .Q(reg_www_3[3]) );
  dff_sg \reg_ww_3_reg[2]  ( .D(n45141), .CP(clk), .Q(reg_ww_3[2]) );
  dff_sg \reg_www_3_reg[2]  ( .D(n44984), .CP(clk), .Q(reg_www_3[2]) );
  dff_sg \reg_ww_3_reg[1]  ( .D(n45140), .CP(clk), .Q(reg_ww_3[1]) );
  dff_sg \reg_www_3_reg[1]  ( .D(n45495), .CP(clk), .Q(reg_www_3[1]) );
  dff_sg \reg_ww_3_reg[0]  ( .D(n45144), .CP(clk), .Q(reg_ww_3[0]) );
  dff_sg \reg_www_3_reg[0]  ( .D(n44981), .CP(clk), .Q(reg_www_3[0]) );
  dff_sg \reg_ww_2_reg[19]  ( .D(n45427), .CP(clk), .Q(reg_ww_2[19]) );
  dff_sg \reg_www_2_reg[19]  ( .D(n45143), .CP(clk), .Q(reg_www_2[19]) );
  dff_sg \reg_ww_2_reg[18]  ( .D(n44283), .CP(clk), .Q(reg_ww_2[18]) );
  dff_sg \reg_www_2_reg[18]  ( .D(n44274), .CP(clk), .Q(reg_www_2[18]) );
  dff_sg \reg_ww_2_reg[17]  ( .D(n44282), .CP(clk), .Q(reg_ww_2[17]) );
  dff_sg \reg_www_2_reg[17]  ( .D(n44273), .CP(clk), .Q(reg_www_2[17]) );
  dff_sg \reg_ww_2_reg[16]  ( .D(n44482), .CP(clk), .Q(reg_ww_2[16]) );
  dff_sg \reg_www_2_reg[16]  ( .D(n44277), .CP(clk), .Q(reg_www_2[16]) );
  dff_sg \reg_ww_2_reg[15]  ( .D(n45439), .CP(clk), .Q(reg_ww_2[15]) );
  dff_sg \reg_www_2_reg[15]  ( .D(n44276), .CP(clk), .Q(reg_www_2[15]) );
  dff_sg \reg_ww_2_reg[14]  ( .D(n45437), .CP(clk), .Q(reg_ww_2[14]) );
  dff_sg \reg_www_2_reg[14]  ( .D(n45496), .CP(clk), .Q(reg_www_2[14]) );
  dff_sg \reg_ww_2_reg[13]  ( .D(n45438), .CP(clk), .Q(reg_ww_2[13]) );
  dff_sg \reg_www_2_reg[13]  ( .D(n45497), .CP(clk), .Q(reg_www_2[13]) );
  dff_sg \reg_ww_2_reg[12]  ( .D(n44564), .CP(clk), .Q(reg_ww_2[12]) );
  dff_sg \reg_www_2_reg[12]  ( .D(n45430), .CP(clk), .Q(reg_www_2[12]) );
  dff_sg \reg_ww_2_reg[11]  ( .D(n44551), .CP(clk), .Q(reg_ww_2[11]) );
  dff_sg \reg_www_2_reg[11]  ( .D(n45431), .CP(clk), .Q(reg_www_2[11]) );
  dff_sg \reg_ww_2_reg[10]  ( .D(n44711), .CP(clk), .Q(reg_ww_2[10]) );
  dff_sg \reg_www_2_reg[10]  ( .D(n45428), .CP(clk), .Q(reg_www_2[10]) );
  dff_sg \reg_ww_2_reg[9]  ( .D(n44708), .CP(clk), .Q(reg_ww_2[9]) );
  dff_sg \reg_www_2_reg[9]  ( .D(n45429), .CP(clk), .Q(reg_www_2[9]) );
  dff_sg \reg_ww_2_reg[8]  ( .D(n44702), .CP(clk), .Q(reg_ww_2[8]) );
  dff_sg \reg_www_2_reg[8]  ( .D(n45434), .CP(clk), .Q(reg_www_2[8]) );
  dff_sg \reg_ww_2_reg[7]  ( .D(n44699), .CP(clk), .Q(reg_ww_2[7]) );
  dff_sg \reg_www_2_reg[7]  ( .D(n45435), .CP(clk), .Q(reg_www_2[7]) );
  dff_sg \reg_ww_2_reg[6]  ( .D(n44759), .CP(clk), .Q(reg_ww_2[6]) );
  dff_sg \reg_www_2_reg[6]  ( .D(n45432), .CP(clk), .Q(reg_www_2[6]) );
  dff_sg \reg_ww_2_reg[5]  ( .D(n44768), .CP(clk), .Q(reg_ww_2[5]) );
  dff_sg \reg_www_2_reg[5]  ( .D(n45433), .CP(clk), .Q(reg_www_2[5]) );
  dff_sg \reg_ww_2_reg[4]  ( .D(n44720), .CP(clk), .Q(reg_ww_2[4]) );
  dff_sg \reg_www_2_reg[4]  ( .D(n45009), .CP(clk), .Q(reg_www_2[4]) );
  dff_sg \reg_ww_2_reg[3]  ( .D(n44717), .CP(clk), .Q(reg_ww_2[3]) );
  dff_sg \reg_www_2_reg[3]  ( .D(n45006), .CP(clk), .Q(reg_www_2[3]) );
  dff_sg \reg_ww_2_reg[2]  ( .D(n44663), .CP(clk), .Q(reg_ww_2[2]) );
  dff_sg \reg_www_2_reg[2]  ( .D(n45424), .CP(clk), .Q(reg_www_2[2]) );
  dff_sg \reg_ww_2_reg[1]  ( .D(n44285), .CP(clk), .Q(reg_ww_2[1]) );
  dff_sg \reg_www_2_reg[1]  ( .D(n45425), .CP(clk), .Q(reg_www_2[1]) );
  dff_sg \reg_ww_2_reg[0]  ( .D(n44645), .CP(clk), .Q(reg_ww_2[0]) );
  dff_sg \reg_www_2_reg[0]  ( .D(n45426), .CP(clk), .Q(reg_www_2[0]) );
  dff_sg \reg_ww_1_reg[19]  ( .D(n44621), .CP(clk), .Q(reg_ww_1[19]) );
  dff_sg \reg_www_1_reg[19]  ( .D(n44642), .CP(clk), .Q(reg_www_1[19]) );
  dff_sg \reg_ww_1_reg[18]  ( .D(n44786), .CP(clk), .Q(reg_ww_1[18]) );
  dff_sg \reg_www_1_reg[18]  ( .D(n44696), .CP(clk), .Q(reg_www_1[18]) );
  dff_sg \reg_ww_1_reg[17]  ( .D(n44783), .CP(clk), .Q(reg_ww_1[17]) );
  dff_sg \reg_www_1_reg[17]  ( .D(n44693), .CP(clk), .Q(reg_www_1[17]) );
  dff_sg \reg_ww_1_reg[16]  ( .D(n44765), .CP(clk), .Q(reg_ww_1[16]) );
  dff_sg \reg_www_1_reg[16]  ( .D(n44678), .CP(clk), .Q(reg_www_1[16]) );
  dff_sg \reg_ww_1_reg[15]  ( .D(n44756), .CP(clk), .Q(reg_ww_1[15]) );
  dff_sg \reg_www_1_reg[15]  ( .D(n44675), .CP(clk), .Q(reg_www_1[15]) );
  dff_sg \reg_ww_1_reg[14]  ( .D(n44855), .CP(clk), .Q(reg_ww_1[14]) );
  dff_sg \reg_www_1_reg[14]  ( .D(n44687), .CP(clk), .Q(reg_www_1[14]) );
  dff_sg \reg_ww_1_reg[13]  ( .D(n44861), .CP(clk), .Q(reg_ww_1[13]) );
  dff_sg \reg_www_1_reg[13]  ( .D(n44672), .CP(clk), .Q(reg_www_1[13]) );
  dff_sg \reg_ww_1_reg[12]  ( .D(n44852), .CP(clk), .Q(reg_ww_1[12]) );
  dff_sg \reg_www_1_reg[12]  ( .D(n44367), .CP(clk), .Q(reg_www_1[12]) );
  dff_sg \reg_ww_1_reg[11]  ( .D(n44792), .CP(clk), .Q(reg_ww_1[11]) );
  dff_sg \reg_www_1_reg[11]  ( .D(n45405), .CP(clk), .Q(reg_www_1[11]) );
  dff_sg \reg_ww_1_reg[10]  ( .D(n45416), .CP(clk), .Q(reg_ww_1[10]) );
  dff_sg \reg_www_1_reg[10]  ( .D(n45404), .CP(clk), .Q(reg_www_1[10]) );
  dff_sg \reg_ww_1_reg[9]  ( .D(n45417), .CP(clk), .Q(reg_ww_1[9]) );
  dff_sg \reg_www_1_reg[9]  ( .D(n44633), .CP(clk), .Q(reg_www_1[9]) );
  dff_sg \reg_ww_1_reg[8]  ( .D(n44279), .CP(clk), .Q(reg_ww_1[8]) );
  dff_sg \reg_www_1_reg[8]  ( .D(n45408), .CP(clk), .Q(reg_www_1[8]) );
  dff_sg \reg_ww_1_reg[7]  ( .D(n44278), .CP(clk), .Q(reg_ww_1[7]) );
  dff_sg \reg_www_1_reg[7]  ( .D(n45409), .CP(clk), .Q(reg_www_1[7]) );
  dff_sg \reg_ww_1_reg[6]  ( .D(n44930), .CP(clk), .Q(reg_ww_1[6]) );
  dff_sg \reg_www_1_reg[6]  ( .D(n44627), .CP(clk), .Q(reg_www_1[6]) );
  dff_sg \reg_ww_1_reg[5]  ( .D(n44927), .CP(clk), .Q(reg_ww_1[5]) );
  dff_sg \reg_www_1_reg[5]  ( .D(n44576), .CP(clk), .Q(reg_www_1[5]) );
  dff_sg \reg_ww_1_reg[4]  ( .D(n44921), .CP(clk), .Q(reg_ww_1[4]) );
  dff_sg \reg_www_1_reg[4]  ( .D(n44573), .CP(clk), .Q(reg_www_1[4]) );
  dff_sg \reg_ww_1_reg[3]  ( .D(n44918), .CP(clk), .Q(reg_ww_1[3]) );
  dff_sg \reg_www_1_reg[3]  ( .D(n44570), .CP(clk), .Q(reg_www_1[3]) );
  dff_sg \reg_ww_1_reg[2]  ( .D(n45475), .CP(clk), .Q(reg_ww_1[2]) );
  dff_sg \reg_www_1_reg[2]  ( .D(n44651), .CP(clk), .Q(reg_www_1[2]) );
  dff_sg \reg_ww_1_reg[1]  ( .D(n45476), .CP(clk), .Q(reg_ww_1[1]) );
  dff_sg \reg_www_1_reg[1]  ( .D(n44657), .CP(clk), .Q(reg_www_1[1]) );
  dff_sg \reg_ww_1_reg[0]  ( .D(n44747), .CP(clk), .Q(reg_ww_1[0]) );
  dff_sg \reg_www_1_reg[0]  ( .D(n44624), .CP(clk), .Q(reg_www_1[0]) );
  dff_sg \reg_ww_0_reg[19]  ( .D(n45484), .CP(clk), .Q(reg_ww_0[19]) );
  dff_sg \reg_www_0_reg[19]  ( .D(n44744), .CP(clk), .Q(reg_www_0[19]) );
  dff_sg \reg_ww_0_reg[18]  ( .D(n45481), .CP(clk), .Q(reg_ww_0[18]) );
  dff_sg \reg_www_0_reg[18]  ( .D(n44636), .CP(clk), .Q(reg_www_0[18]) );
  dff_sg \reg_ww_0_reg[17]  ( .D(n45482), .CP(clk), .Q(reg_ww_0[17]) );
  dff_sg \reg_www_0_reg[17]  ( .D(n44780), .CP(clk), .Q(reg_www_0[17]) );
  dff_sg \reg_ww_0_reg[16]  ( .D(n45450), .CP(clk), .Q(reg_ww_0[16]) );
  dff_sg \reg_www_0_reg[16]  ( .D(n44774), .CP(clk), .Q(reg_www_0[16]) );
  dff_sg \reg_ww_0_reg[15]  ( .D(n45451), .CP(clk), .Q(reg_ww_0[15]) );
  dff_sg \reg_www_0_reg[15]  ( .D(n45474), .CP(clk), .Q(reg_www_0[15]) );
  dff_sg \reg_ww_0_reg[14]  ( .D(n45448), .CP(clk), .Q(reg_ww_0[14]) );
  dff_sg \reg_www_0_reg[14]  ( .D(n44705), .CP(clk), .Q(reg_www_0[14]) );
  dff_sg \reg_ww_0_reg[13]  ( .D(n45449), .CP(clk), .Q(reg_ww_0[13]) );
  dff_sg \reg_www_0_reg[13]  ( .D(n44684), .CP(clk), .Q(reg_www_0[13]) );
  dff_sg \reg_ww_0_reg[12]  ( .D(n45454), .CP(clk), .Q(reg_ww_0[12]) );
  dff_sg \reg_www_0_reg[12]  ( .D(n44681), .CP(clk), .Q(reg_www_0[12]) );
  dff_sg \reg_ww_0_reg[11]  ( .D(n45455), .CP(clk), .Q(reg_ww_0[11]) );
  dff_sg \reg_www_0_reg[11]  ( .D(n44639), .CP(clk), .Q(reg_www_0[11]) );
  dff_sg \reg_ww_0_reg[10]  ( .D(n45452), .CP(clk), .Q(reg_ww_0[10]) );
  dff_sg \reg_www_0_reg[10]  ( .D(n44732), .CP(clk), .Q(reg_www_0[10]) );
  dff_sg \reg_ww_0_reg[9]  ( .D(n45453), .CP(clk), .Q(reg_ww_0[9]) );
  dff_sg \reg_www_0_reg[9]  ( .D(n44738), .CP(clk), .Q(reg_www_0[9]) );
  dff_sg \reg_ww_0_reg[8]  ( .D(n45442), .CP(clk), .Q(reg_ww_0[8]) );
  dff_sg \reg_www_0_reg[8]  ( .D(n44729), .CP(clk), .Q(reg_www_0[8]) );
  dff_sg \reg_ww_0_reg[7]  ( .D(n45443), .CP(clk), .Q(reg_ww_0[7]) );
  dff_sg \reg_www_0_reg[7]  ( .D(n44726), .CP(clk), .Q(reg_www_0[7]) );
  dff_sg \reg_ww_0_reg[6]  ( .D(n45440), .CP(clk), .Q(reg_ww_0[6]) );
  dff_sg \reg_www_0_reg[6]  ( .D(n45487), .CP(clk), .Q(reg_www_0[6]) );
  dff_sg \reg_ww_0_reg[5]  ( .D(n45441), .CP(clk), .Q(reg_ww_0[5]) );
  dff_sg \reg_www_0_reg[5]  ( .D(n45488), .CP(clk), .Q(reg_www_0[5]) );
  dff_sg \reg_ww_0_reg[4]  ( .D(n45446), .CP(clk), .Q(reg_ww_0[4]) );
  dff_sg \reg_www_0_reg[4]  ( .D(n45479), .CP(clk), .Q(reg_www_0[4]) );
  dff_sg \reg_ww_0_reg[3]  ( .D(n45447), .CP(clk), .Q(reg_ww_0[3]) );
  dff_sg \reg_www_0_reg[3]  ( .D(n45480), .CP(clk), .Q(reg_www_0[3]) );
  dff_sg \reg_ww_0_reg[2]  ( .D(n45444), .CP(clk), .Q(reg_ww_0[2]) );
  dff_sg \reg_www_0_reg[2]  ( .D(n45477), .CP(clk), .Q(reg_www_0[2]) );
  dff_sg \reg_ww_0_reg[1]  ( .D(n45445), .CP(clk), .Q(reg_ww_0[1]) );
  dff_sg \reg_www_0_reg[1]  ( .D(n45478), .CP(clk), .Q(reg_www_0[1]) );
  dff_sg \reg_ww_0_reg[0]  ( .D(n45466), .CP(clk), .Q(reg_ww_0[0]) );
  dff_sg \reg_www_0_reg[0]  ( .D(n45483), .CP(clk), .Q(reg_www_0[0]) );
  dff_sg \reg_ii_15_reg[19]  ( .D(n45520), .CP(clk), .Q(reg_ii_15[19]) );
  dff_sg \reg_iii_15_reg[19]  ( .D(n45467), .CP(clk), .Q(reg_iii_15[19]) );
  dff_sg \reg_ii_15_reg[18]  ( .D(n45410), .CP(clk), .Q(reg_ii_15[18]) );
  dff_sg \reg_iii_15_reg[18]  ( .D(n45464), .CP(clk), .Q(reg_iii_15[18]) );
  dff_sg \reg_ii_15_reg[17]  ( .D(n45412), .CP(clk), .Q(reg_ii_15[17]) );
  dff_sg \reg_iii_15_reg[17]  ( .D(n45465), .CP(clk), .Q(reg_iii_15[17]) );
  dff_sg \reg_ii_15_reg[16]  ( .D(n45401), .CP(clk), .Q(reg_ii_15[16]) );
  dff_sg \reg_iii_15_reg[16]  ( .D(n45470), .CP(clk), .Q(reg_iii_15[16]) );
  dff_sg \reg_ii_15_reg[15]  ( .D(n45149), .CP(clk), .Q(reg_ii_15[15]) );
  dff_sg \reg_iii_15_reg[15]  ( .D(n45471), .CP(clk), .Q(reg_iii_15[15]) );
  dff_sg \reg_ii_15_reg[14]  ( .D(n45419), .CP(clk), .Q(reg_ii_15[14]) );
  dff_sg \reg_iii_15_reg[14]  ( .D(n45468), .CP(clk), .Q(reg_iii_15[14]) );
  dff_sg \reg_ii_15_reg[13]  ( .D(n45420), .CP(clk), .Q(reg_ii_15[13]) );
  dff_sg \reg_iii_15_reg[13]  ( .D(n45469), .CP(clk), .Q(reg_iii_15[13]) );
  dff_sg \reg_ii_15_reg[12]  ( .D(n45181), .CP(clk), .Q(reg_ii_15[12]) );
  dff_sg \reg_iii_15_reg[12]  ( .D(n45458), .CP(clk), .Q(reg_iii_15[12]) );
  dff_sg \reg_ii_15_reg[11]  ( .D(n45237), .CP(clk), .Q(reg_ii_15[11]) );
  dff_sg \reg_iii_15_reg[11]  ( .D(n45459), .CP(clk), .Q(reg_iii_15[11]) );
  dff_sg \reg_ii_15_reg[10]  ( .D(n45402), .CP(clk), .Q(reg_ii_15[10]) );
  dff_sg \reg_iii_15_reg[10]  ( .D(n45456), .CP(clk), .Q(reg_iii_15[10]) );
  dff_sg \reg_ii_15_reg[9]  ( .D(n45545), .CP(clk), .Q(reg_ii_15[9]) );
  dff_sg \reg_iii_15_reg[9]  ( .D(n45457), .CP(clk), .Q(reg_iii_15[9]) );
  dff_sg \reg_ii_15_reg[8]  ( .D(n45192), .CP(clk), .Q(reg_ii_15[8]) );
  dff_sg \reg_iii_15_reg[8]  ( .D(n45462), .CP(clk), .Q(reg_iii_15[8]) );
  dff_sg \reg_ii_15_reg[7]  ( .D(n45193), .CP(clk), .Q(reg_ii_15[7]) );
  dff_sg \reg_iii_15_reg[7]  ( .D(n45463), .CP(clk), .Q(reg_iii_15[7]) );
  dff_sg \reg_ii_15_reg[6]  ( .D(n45191), .CP(clk), .Q(reg_ii_15[6]) );
  dff_sg \reg_iii_15_reg[6]  ( .D(n45460), .CP(clk), .Q(reg_iii_15[6]) );
  dff_sg \reg_ii_15_reg[5]  ( .D(n45182), .CP(clk), .Q(reg_ii_15[5]) );
  dff_sg \reg_iii_15_reg[5]  ( .D(n45461), .CP(clk), .Q(reg_iii_15[5]) );
  dff_sg \reg_ii_15_reg[4]  ( .D(n45196), .CP(clk), .Q(reg_ii_15[4]) );
  dff_sg \reg_iii_15_reg[4]  ( .D(n45517), .CP(clk), .Q(reg_iii_15[4]) );
  dff_sg \reg_ii_15_reg[3]  ( .D(n45197), .CP(clk), .Q(reg_ii_15[3]) );
  dff_sg \reg_iii_15_reg[3]  ( .D(n45261), .CP(clk), .Q(reg_iii_15[3]) );
  dff_sg \reg_ii_15_reg[2]  ( .D(n45194), .CP(clk), .Q(reg_ii_15[2]) );
  dff_sg \reg_iii_15_reg[2]  ( .D(n45406), .CP(clk), .Q(reg_iii_15[2]) );
  dff_sg \reg_ii_15_reg[1]  ( .D(n45195), .CP(clk), .Q(reg_ii_15[1]) );
  dff_sg \reg_iii_15_reg[1]  ( .D(n45411), .CP(clk), .Q(reg_iii_15[1]) );
  dff_sg \reg_ii_15_reg[0]  ( .D(n45186), .CP(clk), .Q(reg_ii_15[0]) );
  dff_sg \reg_iii_15_reg[0]  ( .D(n45521), .CP(clk), .Q(reg_iii_15[0]) );
  dff_sg \reg_ii_14_reg[19]  ( .D(n45187), .CP(clk), .Q(reg_ii_14[19]) );
  dff_sg \reg_iii_14_reg[19]  ( .D(n44959), .CP(clk), .Q(reg_iii_14[19]) );
  dff_sg \reg_ii_14_reg[18]  ( .D(n45183), .CP(clk), .Q(reg_ii_14[18]) );
  dff_sg \reg_iii_14_reg[18]  ( .D(n44958), .CP(clk), .Q(reg_iii_14[18]) );
  dff_sg \reg_ii_14_reg[17]  ( .D(n45184), .CP(clk), .Q(reg_ii_14[17]) );
  dff_sg \reg_iii_14_reg[17]  ( .D(n44962), .CP(clk), .Q(reg_iii_14[17]) );
  dff_sg \reg_ww_8_reg[14]  ( .D(n45165), .CP(clk), .Q(reg_ww_8[14]) );
  dff_sg \reg_www_8_reg[14]  ( .D(n45423), .CP(clk), .Q(reg_www_8[14]) );
  dff_sg \reg_ww_8_reg[13]  ( .D(n45540), .CP(clk), .Q(reg_ww_8[13]) );
  dff_sg \reg_www_8_reg[13]  ( .D(n45507), .CP(clk), .Q(reg_www_8[13]) );
  dff_sg \reg_ww_8_reg[12]  ( .D(n45180), .CP(clk), .Q(reg_ww_8[12]) );
  dff_sg \reg_www_8_reg[12]  ( .D(n45500), .CP(clk), .Q(reg_www_8[12]) );
  dff_sg \reg_ww_8_reg[11]  ( .D(n45533), .CP(clk), .Q(reg_ww_8[11]) );
  dff_sg \reg_www_8_reg[11]  ( .D(n45421), .CP(clk), .Q(reg_www_8[11]) );
  dff_sg \reg_ww_8_reg[10]  ( .D(n45549), .CP(clk), .Q(reg_ww_8[10]) );
  dff_sg \reg_www_8_reg[10]  ( .D(n45356), .CP(clk), .Q(reg_www_8[10]) );
  dff_sg \reg_ww_8_reg[9]  ( .D(n45294), .CP(clk), .Q(reg_ww_8[9]) );
  dff_sg \reg_www_8_reg[9]  ( .D(n45489), .CP(clk), .Q(reg_www_8[9]) );
  dff_sg \reg_ww_8_reg[8]  ( .D(n45179), .CP(clk), .Q(reg_ww_8[8]) );
  dff_sg \reg_www_8_reg[8]  ( .D(n45498), .CP(clk), .Q(reg_www_8[8]) );
  dff_sg \reg_ww_8_reg[7]  ( .D(n45178), .CP(clk), .Q(reg_ww_8[7]) );
  dff_sg \reg_www_8_reg[7]  ( .D(n45418), .CP(clk), .Q(reg_www_8[7]) );
  dff_sg \reg_ww_8_reg[6]  ( .D(n45527), .CP(clk), .Q(reg_ww_8[6]) );
  dff_sg \reg_www_8_reg[6]  ( .D(n45414), .CP(clk), .Q(reg_www_8[6]) );
  dff_sg \reg_ww_8_reg[5]  ( .D(n45530), .CP(clk), .Q(reg_ww_8[5]) );
  dff_sg \reg_www_8_reg[5]  ( .D(n45174), .CP(clk), .Q(reg_www_8[5]) );
  dff_sg \reg_ww_8_reg[4]  ( .D(n45176), .CP(clk), .Q(reg_ww_8[4]) );
  dff_sg \reg_www_8_reg[4]  ( .D(n45415), .CP(clk), .Q(reg_www_8[4]) );
  dff_sg \reg_ww_8_reg[3]  ( .D(n45175), .CP(clk), .Q(reg_ww_8[3]) );
  dff_sg \reg_www_8_reg[3]  ( .D(n45173), .CP(clk), .Q(reg_www_8[3]) );
  dff_sg \reg_ww_8_reg[2]  ( .D(n45289), .CP(clk), .Q(reg_ww_8[2]) );
  dff_sg \reg_www_8_reg[2]  ( .D(n45171), .CP(clk), .Q(reg_www_8[2]) );
  dff_sg \reg_ww_8_reg[1]  ( .D(n45155), .CP(clk), .Q(reg_ww_8[1]) );
  dff_sg \reg_www_8_reg[1]  ( .D(n45172), .CP(clk), .Q(reg_www_8[1]) );
  dff_sg \reg_ww_8_reg[0]  ( .D(n45177), .CP(clk), .Q(reg_ww_8[0]) );
  dff_sg \reg_www_8_reg[0]  ( .D(n45413), .CP(clk), .Q(reg_www_8[0]) );
  dff_sg \reg_ww_7_reg[19]  ( .D(n45349), .CP(clk), .Q(reg_ww_7[19]) );
  dff_sg \reg_www_7_reg[19]  ( .D(n45162), .CP(clk), .Q(reg_www_7[19]) );
  dff_sg \reg_ww_7_reg[18]  ( .D(n45385), .CP(clk), .Q(reg_ww_7[18]) );
  dff_sg \reg_www_7_reg[18]  ( .D(n45207), .CP(clk), .Q(reg_www_7[18]) );
  dff_sg \reg_ww_7_reg[17]  ( .D(n45347), .CP(clk), .Q(reg_ww_7[17]) );
  dff_sg \reg_www_7_reg[17]  ( .D(n45200), .CP(clk), .Q(reg_www_7[17]) );
  dff_sg \reg_ww_7_reg[16]  ( .D(n44388), .CP(clk), .Q(reg_ww_7[16]) );
  dff_sg \reg_www_7_reg[16]  ( .D(n45208), .CP(clk), .Q(reg_www_7[16]) );
  dff_sg \reg_ww_7_reg[15]  ( .D(n44387), .CP(clk), .Q(reg_ww_7[15]) );
  dff_sg \reg_www_7_reg[15]  ( .D(n45211), .CP(clk), .Q(reg_www_7[15]) );
  dff_sg \reg_ww_7_reg[14]  ( .D(n44391), .CP(clk), .Q(reg_ww_7[14]) );
  dff_sg \reg_www_7_reg[14]  ( .D(n45212), .CP(clk), .Q(reg_www_7[14]) );
  dff_sg \reg_ww_7_reg[13]  ( .D(n44390), .CP(clk), .Q(reg_ww_7[13]) );
  dff_sg \reg_www_7_reg[13]  ( .D(n45213), .CP(clk), .Q(reg_www_7[13]) );
  dff_sg \reg_ww_7_reg[12]  ( .D(n44382), .CP(clk), .Q(reg_ww_7[12]) );
  dff_sg \reg_www_7_reg[12]  ( .D(n45209), .CP(clk), .Q(reg_www_7[12]) );
  dff_sg \reg_ww_7_reg[11]  ( .D(n44381), .CP(clk), .Q(reg_ww_7[11]) );
  dff_sg \reg_www_7_reg[11]  ( .D(n45210), .CP(clk), .Q(reg_www_7[11]) );
  dff_sg \reg_ww_7_reg[10]  ( .D(n44385), .CP(clk), .Q(reg_ww_7[10]) );
  dff_sg \reg_www_7_reg[10]  ( .D(n45201), .CP(clk), .Q(reg_www_7[10]) );
  dff_sg \reg_ww_7_reg[9]  ( .D(n44384), .CP(clk), .Q(reg_ww_7[9]) );
  dff_sg \reg_www_7_reg[9]  ( .D(n45202), .CP(clk), .Q(reg_www_7[9]) );
  dff_sg \reg_ww_7_reg[8]  ( .D(n44395), .CP(clk), .Q(reg_ww_7[8]) );
  dff_sg \reg_www_7_reg[8]  ( .D(n45198), .CP(clk), .Q(reg_www_7[8]) );
  dff_sg \reg_ww_7_reg[7]  ( .D(n44394), .CP(clk), .Q(reg_ww_7[7]) );
  dff_sg \reg_www_7_reg[7]  ( .D(n45199), .CP(clk), .Q(reg_www_7[7]) );
  dff_sg \reg_ww_7_reg[6]  ( .D(n44398), .CP(clk), .Q(reg_ww_7[6]) );
  dff_sg \reg_www_7_reg[6]  ( .D(n45205), .CP(clk), .Q(reg_www_7[6]) );
  dff_sg \reg_ww_7_reg[5]  ( .D(n44397), .CP(clk), .Q(reg_ww_7[5]) );
  dff_sg \reg_www_7_reg[5]  ( .D(n45206), .CP(clk), .Q(reg_www_7[5]) );
  dff_sg \reg_ww_7_reg[4]  ( .D(n44396), .CP(clk), .Q(reg_ww_7[4]) );
  dff_sg \reg_www_7_reg[4]  ( .D(n45203), .CP(clk), .Q(reg_www_7[4]) );
  dff_sg \reg_ww_7_reg[3]  ( .D(n44393), .CP(clk), .Q(reg_ww_7[3]) );
  dff_sg \reg_www_7_reg[3]  ( .D(n45204), .CP(clk), .Q(reg_www_7[3]) );
  dff_sg \reg_ww_7_reg[2]  ( .D(n44383), .CP(clk), .Q(reg_ww_7[2]) );
  dff_sg \reg_www_7_reg[2]  ( .D(n45386), .CP(clk), .Q(reg_www_7[2]) );
  dff_sg \reg_ww_7_reg[1]  ( .D(n44392), .CP(clk), .Q(reg_ww_7[1]) );
  dff_sg \reg_www_7_reg[1]  ( .D(n45387), .CP(clk), .Q(reg_www_7[1]) );
  dff_sg \reg_ww_7_reg[0]  ( .D(n44372), .CP(clk), .Q(reg_ww_7[0]) );
  dff_sg \reg_www_7_reg[0]  ( .D(n45348), .CP(clk), .Q(reg_www_7[0]) );
  dff_sg \reg_ww_6_reg[19]  ( .D(n45019), .CP(clk), .Q(reg_ww_6[19]) );
  dff_sg \reg_www_6_reg[19]  ( .D(n44371), .CP(clk), .Q(reg_www_6[19]) );
  dff_sg \reg_ww_6_reg[18]  ( .D(n45023), .CP(clk), .Q(reg_ww_6[18]) );
  dff_sg \reg_www_6_reg[18]  ( .D(n44361), .CP(clk), .Q(reg_www_6[18]) );
  dff_sg \reg_ww_6_reg[17]  ( .D(n45022), .CP(clk), .Q(reg_ww_6[17]) );
  dff_sg \reg_www_6_reg[17]  ( .D(n44370), .CP(clk), .Q(reg_www_6[17]) );
  dff_sg \reg_ww_6_reg[16]  ( .D(n44409), .CP(clk), .Q(reg_ww_6[16]) );
  dff_sg \reg_www_6_reg[16]  ( .D(n44363), .CP(clk), .Q(reg_www_6[16]) );
  dff_sg \reg_ww_6_reg[15]  ( .D(n44408), .CP(clk), .Q(reg_ww_6[15]) );
  dff_sg \reg_www_6_reg[15]  ( .D(n44362), .CP(clk), .Q(reg_www_6[15]) );
  dff_sg \reg_ww_6_reg[14]  ( .D(n44412), .CP(clk), .Q(reg_ww_6[14]) );
  dff_sg \reg_www_6_reg[14]  ( .D(n44366), .CP(clk), .Q(reg_www_6[14]) );
  dff_sg \reg_ww_6_reg[13]  ( .D(n44411), .CP(clk), .Q(reg_ww_6[13]) );
  dff_sg \reg_www_6_reg[13]  ( .D(n44365), .CP(clk), .Q(reg_www_6[13]) );
  dff_sg \reg_ww_6_reg[12]  ( .D(n45018), .CP(clk), .Q(reg_ww_6[12]) );
  dff_sg \reg_www_6_reg[12]  ( .D(n44373), .CP(clk), .Q(reg_www_6[12]) );
  dff_sg \reg_ww_6_reg[11]  ( .D(n44406), .CP(clk), .Q(reg_ww_6[11]) );
  dff_sg \reg_www_6_reg[11]  ( .D(n44377), .CP(clk), .Q(reg_www_6[11]) );
  dff_sg \reg_ww_6_reg[10]  ( .D(n45021), .CP(clk), .Q(reg_ww_6[10]) );
  dff_sg \reg_www_6_reg[10]  ( .D(n44374), .CP(clk), .Q(reg_www_6[10]) );
  dff_sg \reg_ww_6_reg[9]  ( .D(n44290), .CP(clk), .Q(reg_ww_6[9]) );
  dff_sg \reg_www_6_reg[9]  ( .D(n44380), .CP(clk), .Q(reg_www_6[9]) );
  dff_sg \reg_ww_6_reg[8]  ( .D(n44400), .CP(clk), .Q(reg_ww_6[8]) );
  dff_sg \reg_www_6_reg[8]  ( .D(n44376), .CP(clk), .Q(reg_www_6[8]) );
  dff_sg \reg_ww_6_reg[7]  ( .D(n44413), .CP(clk), .Q(reg_ww_6[7]) );
  dff_sg \reg_www_6_reg[7]  ( .D(n44375), .CP(clk), .Q(reg_www_6[7]) );
  dff_sg \reg_ww_6_reg[6]  ( .D(n44415), .CP(clk), .Q(reg_ww_6[6]) );
  dff_sg \reg_www_6_reg[6]  ( .D(n44379), .CP(clk), .Q(reg_www_6[6]) );
  dff_sg \reg_ww_6_reg[5]  ( .D(n44414), .CP(clk), .Q(reg_ww_6[5]) );
  dff_sg \reg_www_6_reg[5]  ( .D(n44378), .CP(clk), .Q(reg_www_6[5]) );
  dff_sg \reg_ww_6_reg[4]  ( .D(n44402), .CP(clk), .Q(reg_ww_6[4]) );
  dff_sg \reg_www_6_reg[4]  ( .D(n45025), .CP(clk), .Q(reg_www_6[4]) );
  dff_sg \reg_ww_6_reg[3]  ( .D(n44401), .CP(clk), .Q(reg_ww_6[3]) );
  dff_sg \reg_www_6_reg[3]  ( .D(n45024), .CP(clk), .Q(reg_www_6[3]) );
  dff_sg \reg_ww_6_reg[2]  ( .D(n44405), .CP(clk), .Q(reg_ww_6[2]) );
  dff_sg \reg_www_6_reg[2]  ( .D(n45027), .CP(clk), .Q(reg_www_6[2]) );
  dff_sg \reg_ww_6_reg[1]  ( .D(n44404), .CP(clk), .Q(reg_ww_6[1]) );
  dff_sg \reg_www_6_reg[1]  ( .D(n45026), .CP(clk), .Q(reg_www_6[1]) );
  dff_sg \reg_ww_6_reg[0]  ( .D(n44416), .CP(clk), .Q(reg_ww_6[0]) );
  dff_sg \reg_www_6_reg[0]  ( .D(n45020), .CP(clk), .Q(reg_www_6[0]) );
  dff_sg \reg_ww_5_reg[19]  ( .D(n44317), .CP(clk), .Q(reg_ww_5[19]) );
  dff_sg \reg_www_5_reg[19]  ( .D(n44420), .CP(clk), .Q(reg_www_5[19]) );
  dff_sg \reg_ww_5_reg[18]  ( .D(n44321), .CP(clk), .Q(reg_ww_5[18]) );
  dff_sg \reg_www_5_reg[18]  ( .D(n44417), .CP(clk), .Q(reg_www_5[18]) );
  dff_sg \reg_ww_5_reg[17]  ( .D(n44320), .CP(clk), .Q(reg_ww_5[17]) );
  dff_sg \reg_www_5_reg[17]  ( .D(n44399), .CP(clk), .Q(reg_www_5[17]) );
  dff_sg \reg_ww_5_reg[16]  ( .D(n44299), .CP(clk), .Q(reg_ww_5[16]) );
  dff_sg \reg_www_5_reg[16]  ( .D(n44419), .CP(clk), .Q(reg_www_5[16]) );
  dff_sg \reg_ww_5_reg[15]  ( .D(n44298), .CP(clk), .Q(reg_ww_5[15]) );
  dff_sg \reg_www_5_reg[15]  ( .D(n44418), .CP(clk), .Q(reg_www_5[15]) );
  dff_sg \reg_ww_5_reg[14]  ( .D(n44291), .CP(clk), .Q(reg_ww_5[14]) );
  dff_sg \reg_www_5_reg[14]  ( .D(n44422), .CP(clk), .Q(reg_www_5[14]) );
  dff_sg \reg_ww_5_reg[13]  ( .D(n44297), .CP(clk), .Q(reg_ww_5[13]) );
  dff_sg \reg_www_5_reg[13]  ( .D(n44421), .CP(clk), .Q(reg_www_5[13]) );
  dff_sg \reg_ww_5_reg[12]  ( .D(n44293), .CP(clk), .Q(reg_ww_5[12]) );
  dff_sg \reg_www_5_reg[12]  ( .D(n44312), .CP(clk), .Q(reg_www_5[12]) );
  dff_sg \reg_ww_5_reg[11]  ( .D(n44292), .CP(clk), .Q(reg_ww_5[11]) );
  dff_sg \reg_www_5_reg[11]  ( .D(n44311), .CP(clk), .Q(reg_www_5[11]) );
  dff_sg \reg_ww_5_reg[10]  ( .D(n44296), .CP(clk), .Q(reg_ww_5[10]) );
  dff_sg \reg_www_5_reg[10]  ( .D(n44315), .CP(clk), .Q(reg_www_5[10]) );
  dff_sg \reg_ww_5_reg[9]  ( .D(n44295), .CP(clk), .Q(reg_ww_5[9]) );
  dff_sg \reg_www_5_reg[9]  ( .D(n44314), .CP(clk), .Q(reg_www_5[9]) );
  dff_sg \reg_ww_5_reg[8]  ( .D(n44305), .CP(clk), .Q(reg_ww_5[8]) );
  dff_sg \reg_www_5_reg[8]  ( .D(n44309), .CP(clk), .Q(reg_www_5[8]) );
  dff_sg \reg_ww_5_reg[7]  ( .D(n44304), .CP(clk), .Q(reg_ww_5[7]) );
  dff_sg \reg_www_5_reg[7]  ( .D(n44313), .CP(clk), .Q(reg_www_5[7]) );
  dff_sg \reg_ww_5_reg[6]  ( .D(n44308), .CP(clk), .Q(reg_ww_5[6]) );
  dff_sg \reg_www_5_reg[6]  ( .D(n44310), .CP(clk), .Q(reg_www_5[6]) );
  dff_sg \reg_ww_5_reg[5]  ( .D(n44307), .CP(clk), .Q(reg_ww_5[5]) );
  dff_sg \reg_www_5_reg[5]  ( .D(n44303), .CP(clk), .Q(reg_www_5[5]) );
  dff_sg \reg_ww_5_reg[4]  ( .D(n44294), .CP(clk), .Q(reg_ww_5[4]) );
  dff_sg \reg_www_5_reg[4]  ( .D(n44327), .CP(clk), .Q(reg_www_5[4]) );
  dff_sg \reg_ww_5_reg[3]  ( .D(n44300), .CP(clk), .Q(reg_ww_5[3]) );
  dff_sg \reg_www_5_reg[3]  ( .D(n44326), .CP(clk), .Q(reg_www_5[3]) );
  dff_sg \reg_ww_5_reg[2]  ( .D(n44302), .CP(clk), .Q(reg_ww_5[2]) );
  dff_sg \reg_www_5_reg[2]  ( .D(n44316), .CP(clk), .Q(reg_www_5[2]) );
  dff_sg \reg_ww_5_reg[1]  ( .D(n44301), .CP(clk), .Q(reg_ww_5[1]) );
  dff_sg \reg_www_5_reg[1]  ( .D(n44325), .CP(clk), .Q(reg_www_5[1]) );
  dff_sg \reg_ww_5_reg[0]  ( .D(n44350), .CP(clk), .Q(reg_ww_5[0]) );
  dff_sg \reg_www_5_reg[0]  ( .D(n44318), .CP(clk), .Q(reg_www_5[0]) );
  dff_sg \reg_ww_4_reg[19]  ( .D(n44330), .CP(clk), .Q(reg_ww_4[19]) );
  dff_sg \reg_www_4_reg[19]  ( .D(n44349), .CP(clk), .Q(reg_www_4[19]) );
  dff_sg \reg_ww_4_reg[18]  ( .D(n44334), .CP(clk), .Q(reg_ww_4[18]) );
  dff_sg \reg_www_4_reg[18]  ( .D(n44353), .CP(clk), .Q(reg_www_4[18]) );
  dff_sg \reg_ww_4_reg[17]  ( .D(n44333), .CP(clk), .Q(reg_ww_4[17]) );
  dff_sg \reg_www_4_reg[17]  ( .D(n44352), .CP(clk), .Q(reg_www_4[17]) );
  dff_sg \reg_ww_4_reg[16]  ( .D(n44343), .CP(clk), .Q(reg_ww_4[16]) );
  dff_sg \reg_www_4_reg[16]  ( .D(n44341), .CP(clk), .Q(reg_www_4[16]) );
  dff_sg \reg_ww_4_reg[15]  ( .D(n44342), .CP(clk), .Q(reg_ww_4[15]) );
  dff_sg \reg_www_4_reg[15]  ( .D(n44347), .CP(clk), .Q(reg_www_4[15]) );
  dff_sg \reg_ww_4_reg[14]  ( .D(n44346), .CP(clk), .Q(reg_ww_4[14]) );
  dff_sg \reg_www_4_reg[14]  ( .D(n44338), .CP(clk), .Q(reg_www_4[14]) );
  dff_sg \reg_ww_4_reg[13]  ( .D(n44345), .CP(clk), .Q(reg_ww_4[13]) );
  dff_sg \reg_www_4_reg[13]  ( .D(n44344), .CP(clk), .Q(reg_www_4[13]) );
  dff_sg \reg_ww_4_reg[12]  ( .D(n44337), .CP(clk), .Q(reg_ww_4[12]) );
  dff_sg \reg_www_4_reg[12]  ( .D(n44348), .CP(clk), .Q(reg_www_4[12]) );
  dff_sg \reg_ww_4_reg[11]  ( .D(n44336), .CP(clk), .Q(reg_ww_4[11]) );
  dff_sg \reg_www_4_reg[11]  ( .D(n44354), .CP(clk), .Q(reg_www_4[11]) );
  dff_sg \reg_ww_4_reg[10]  ( .D(n44340), .CP(clk), .Q(reg_ww_4[10]) );
  dff_sg \reg_www_4_reg[10]  ( .D(n44351), .CP(clk), .Q(reg_www_4[10]) );
  dff_sg \reg_ww_4_reg[9]  ( .D(n44339), .CP(clk), .Q(reg_ww_4[9]) );
  dff_sg \reg_www_4_reg[9]  ( .D(n44355), .CP(clk), .Q(reg_www_4[9]) );
  dff_sg \reg_ww_4_reg[8]  ( .D(n44557), .CP(clk), .Q(reg_ww_4[8]) );
  dff_sg \reg_www_4_reg[8]  ( .D(n44357), .CP(clk), .Q(reg_www_4[8]) );
  dff_sg \reg_ww_4_reg[7]  ( .D(n44556), .CP(clk), .Q(reg_ww_4[7]) );
  dff_sg \reg_www_4_reg[7]  ( .D(n44356), .CP(clk), .Q(reg_www_4[7]) );
  dff_sg \reg_ww_4_reg[6]  ( .D(n44560), .CP(clk), .Q(reg_ww_4[6]) );
  dff_sg \reg_www_4_reg[6]  ( .D(n44360), .CP(clk), .Q(reg_www_4[6]) );
  dff_sg \reg_ww_4_reg[5]  ( .D(n44559), .CP(clk), .Q(reg_ww_4[5]) );
  dff_sg \reg_www_4_reg[5]  ( .D(n44359), .CP(clk), .Q(reg_www_4[5]) );
  dff_sg \reg_ww_4_reg[4]  ( .D(n44554), .CP(clk), .Q(reg_ww_4[4]) );
  dff_sg \reg_www_4_reg[4]  ( .D(n44328), .CP(clk), .Q(reg_www_4[4]) );
  dff_sg \reg_ww_4_reg[3]  ( .D(n44558), .CP(clk), .Q(reg_ww_4[3]) );
  dff_sg \reg_www_4_reg[3]  ( .D(n44332), .CP(clk), .Q(reg_www_4[3]) );
  dff_sg \reg_ww_4_reg[2]  ( .D(n44555), .CP(clk), .Q(reg_ww_4[2]) );
  dff_sg \reg_www_4_reg[2]  ( .D(n44329), .CP(clk), .Q(reg_www_4[2]) );
  dff_sg \reg_ww_4_reg[1]  ( .D(n44548), .CP(clk), .Q(reg_ww_4[1]) );
  dff_sg \reg_www_4_reg[1]  ( .D(n44335), .CP(clk), .Q(reg_www_4[1]) );
  dff_sg \reg_ww_4_reg[0]  ( .D(n44581), .CP(clk), .Q(reg_ww_4[0]) );
  dff_sg \reg_www_4_reg[0]  ( .D(n44331), .CP(clk), .Q(reg_www_4[0]) );
  dff_sg \reg_ww_3_reg[19]  ( .D(n44580), .CP(clk), .Q(reg_ww_3[19]) );
  dff_sg \reg_www_3_reg[19]  ( .D(n45050), .CP(clk), .Q(reg_www_3[19]) );
  dff_sg \reg_ww_3_reg[18]  ( .D(n44561), .CP(clk), .Q(reg_ww_3[18]) );
  dff_sg \reg_www_3_reg[18]  ( .D(n44879), .CP(clk), .Q(reg_www_3[18]) );
  dff_sg \reg_ww_3_reg[17]  ( .D(n44579), .CP(clk), .Q(reg_ww_3[17]) );
  dff_sg \reg_www_3_reg[17]  ( .D(n44876), .CP(clk), .Q(reg_www_3[17]) );
  dff_sg \reg_ww_3_reg[16]  ( .D(n44563), .CP(clk), .Q(reg_ww_3[16]) );
  dff_sg \reg_www_3_reg[16]  ( .D(n44870), .CP(clk), .Q(reg_www_3[16]) );
  dff_sg \reg_ww_13_reg[13]  ( .D(n44603), .CP(clk), .Q(reg_ww_13[13]) );
  dff_sg \reg_www_13_reg[13]  ( .D(n44542), .CP(clk), .Q(reg_www_13[13]) );
  dff_sg \reg_ww_13_reg[12]  ( .D(n44607), .CP(clk), .Q(reg_ww_13[12]) );
  dff_sg \reg_www_13_reg[12]  ( .D(n44538), .CP(clk), .Q(reg_www_13[12]) );
  dff_sg \reg_ww_13_reg[11]  ( .D(n44606), .CP(clk), .Q(reg_ww_13[11]) );
  dff_sg \reg_www_13_reg[11]  ( .D(n44537), .CP(clk), .Q(reg_www_13[11]) );
  dff_sg \reg_ww_13_reg[10]  ( .D(n44595), .CP(clk), .Q(reg_ww_13[10]) );
  dff_sg \reg_www_13_reg[10]  ( .D(n44541), .CP(clk), .Q(reg_www_13[10]) );
  dff_sg \reg_ww_13_reg[9]  ( .D(n44601), .CP(clk), .Q(reg_ww_13[9]) );
  dff_sg \reg_www_13_reg[9]  ( .D(n44540), .CP(clk), .Q(reg_www_13[9]) );
  dff_sg \reg_ww_13_reg[8]  ( .D(n44592), .CP(clk), .Q(reg_ww_13[8]) );
  dff_sg \reg_www_13_reg[8]  ( .D(n44550), .CP(clk), .Q(reg_www_13[8]) );
  dff_sg \reg_ww_13_reg[7]  ( .D(n44598), .CP(clk), .Q(reg_ww_13[7]) );
  dff_sg \reg_www_13_reg[7]  ( .D(n44549), .CP(clk), .Q(reg_www_13[7]) );
  dff_sg \reg_ww_13_reg[6]  ( .D(n44609), .CP(clk), .Q(reg_ww_13[6]) );
  dff_sg \reg_www_13_reg[6]  ( .D(n44553), .CP(clk), .Q(reg_www_13[6]) );
  dff_sg \reg_ww_13_reg[5]  ( .D(n44608), .CP(clk), .Q(reg_ww_13[5]) );
  dff_sg \reg_www_13_reg[5]  ( .D(n44552), .CP(clk), .Q(reg_www_13[5]) );
  dff_sg \reg_ww_13_reg[4]  ( .D(n44602), .CP(clk), .Q(reg_ww_13[4]) );
  dff_sg \reg_www_13_reg[4]  ( .D(n44536), .CP(clk), .Q(reg_www_13[4]) );
  dff_sg \reg_ww_13_reg[3]  ( .D(n44612), .CP(clk), .Q(reg_ww_13[3]) );
  dff_sg \reg_www_13_reg[3]  ( .D(n44545), .CP(clk), .Q(reg_www_13[3]) );
  dff_sg \reg_ww_13_reg[2]  ( .D(n44611), .CP(clk), .Q(reg_ww_13[2]) );
  dff_sg \reg_www_13_reg[2]  ( .D(n44547), .CP(clk), .Q(reg_www_13[2]) );
  dff_sg \reg_ww_13_reg[1]  ( .D(n44610), .CP(clk), .Q(reg_ww_13[1]) );
  dff_sg \reg_www_13_reg[1]  ( .D(n44546), .CP(clk), .Q(reg_www_13[1]) );
  dff_sg \reg_ww_13_reg[0]  ( .D(n44614), .CP(clk), .Q(reg_ww_13[0]) );
  dff_sg \reg_www_13_reg[0]  ( .D(n44604), .CP(clk), .Q(reg_www_13[0]) );
  dff_sg \reg_ww_12_reg[19]  ( .D(n44447), .CP(clk), .Q(reg_ww_12[19]) );
  dff_sg \reg_www_12_reg[19]  ( .D(n44613), .CP(clk), .Q(reg_www_12[19]) );
  dff_sg \reg_ww_12_reg[18]  ( .D(n44440), .CP(clk), .Q(reg_ww_12[18]) );
  dff_sg \reg_www_12_reg[18]  ( .D(n44582), .CP(clk), .Q(reg_www_12[18]) );
  dff_sg \reg_ww_12_reg[17]  ( .D(n44439), .CP(clk), .Q(reg_ww_12[17]) );
  dff_sg \reg_www_12_reg[17]  ( .D(n44586), .CP(clk), .Q(reg_www_12[17]) );
  dff_sg \reg_ww_12_reg[16]  ( .D(n44443), .CP(clk), .Q(reg_ww_12[16]) );
  dff_sg \reg_www_12_reg[16]  ( .D(n44583), .CP(clk), .Q(reg_www_12[16]) );
  dff_sg \reg_ww_12_reg[15]  ( .D(n44442), .CP(clk), .Q(reg_ww_12[15]) );
  dff_sg \reg_www_12_reg[15]  ( .D(n44589), .CP(clk), .Q(reg_www_12[15]) );
  dff_sg \reg_ww_12_reg[14]  ( .D(n44451), .CP(clk), .Q(reg_ww_12[14]) );
  dff_sg \reg_www_12_reg[14]  ( .D(n44585), .CP(clk), .Q(reg_www_12[14]) );
  dff_sg \reg_ww_12_reg[13]  ( .D(n44450), .CP(clk), .Q(reg_ww_12[13]) );
  dff_sg \reg_www_12_reg[13]  ( .D(n44584), .CP(clk), .Q(reg_www_12[13]) );
  dff_sg \reg_ww_12_reg[12]  ( .D(n44457), .CP(clk), .Q(reg_ww_12[12]) );
  dff_sg \reg_www_12_reg[12]  ( .D(n44588), .CP(clk), .Q(reg_www_12[12]) );
  dff_sg \reg_ww_12_reg[11]  ( .D(n44454), .CP(clk), .Q(reg_ww_12[11]) );
  dff_sg \reg_www_12_reg[11]  ( .D(n44587), .CP(clk), .Q(reg_www_12[11]) );
  dff_sg \reg_ww_12_reg[10]  ( .D(n44453), .CP(clk), .Q(reg_ww_12[10]) );
  dff_sg \reg_www_12_reg[10]  ( .D(n44597), .CP(clk), .Q(reg_www_12[10]) );
  dff_sg \reg_ww_12_reg[9]  ( .D(n44452), .CP(clk), .Q(reg_ww_12[9]) );
  dff_sg \reg_www_12_reg[9]  ( .D(n44596), .CP(clk), .Q(reg_www_12[9]) );
  dff_sg \reg_ww_12_reg[8]  ( .D(n44456), .CP(clk), .Q(reg_ww_12[8]) );
  dff_sg \reg_www_12_reg[8]  ( .D(n44600), .CP(clk), .Q(reg_www_12[8]) );
  dff_sg \reg_ww_12_reg[7]  ( .D(n44455), .CP(clk), .Q(reg_ww_12[7]) );
  dff_sg \reg_www_12_reg[7]  ( .D(n44599), .CP(clk), .Q(reg_www_12[7]) );
  dff_sg \reg_ww_12_reg[6]  ( .D(n44434), .CP(clk), .Q(reg_ww_12[6]) );
  dff_sg \reg_www_12_reg[6]  ( .D(n44591), .CP(clk), .Q(reg_www_12[6]) );
  dff_sg \reg_ww_12_reg[5]  ( .D(n44433), .CP(clk), .Q(reg_ww_12[5]) );
  dff_sg \reg_www_12_reg[5]  ( .D(n44590), .CP(clk), .Q(reg_www_12[5]) );
  dff_sg \reg_ww_12_reg[4]  ( .D(n44437), .CP(clk), .Q(reg_ww_12[4]) );
  dff_sg \reg_www_12_reg[4]  ( .D(n44594), .CP(clk), .Q(reg_www_12[4]) );
  dff_sg \reg_ww_12_reg[3]  ( .D(n44436), .CP(clk), .Q(reg_ww_12[3]) );
  dff_sg \reg_www_12_reg[3]  ( .D(n44593), .CP(clk), .Q(reg_www_12[3]) );
  dff_sg \reg_ww_12_reg[2]  ( .D(n44407), .CP(clk), .Q(reg_ww_12[2]) );
  dff_sg \reg_www_12_reg[2]  ( .D(n44449), .CP(clk), .Q(reg_www_12[2]) );
  dff_sg \reg_ww_12_reg[1]  ( .D(n44429), .CP(clk), .Q(reg_ww_12[1]) );
  dff_sg \reg_www_12_reg[1]  ( .D(n44448), .CP(clk), .Q(reg_www_12[1]) );
  dff_sg \reg_ww_12_reg[0]  ( .D(n44431), .CP(clk), .Q(reg_ww_12[0]) );
  dff_sg \reg_www_12_reg[0]  ( .D(n44438), .CP(clk), .Q(reg_www_12[0]) );
  dff_sg \reg_ww_11_reg[19]  ( .D(n44532), .CP(clk), .Q(reg_ww_11[19]) );
  dff_sg \reg_www_11_reg[19]  ( .D(n44430), .CP(clk), .Q(reg_www_11[19]) );
  dff_sg \reg_ww_11_reg[18]  ( .D(n44525), .CP(clk), .Q(reg_ww_11[18]) );
  dff_sg \reg_www_11_reg[18]  ( .D(n44426), .CP(clk), .Q(reg_www_11[18]) );
  dff_sg \reg_ww_11_reg[17]  ( .D(n44524), .CP(clk), .Q(reg_ww_11[17]) );
  dff_sg \reg_www_11_reg[17]  ( .D(n44423), .CP(clk), .Q(reg_www_11[17]) );
  dff_sg \reg_ww_11_reg[16]  ( .D(n44528), .CP(clk), .Q(reg_ww_11[16]) );
  dff_sg \reg_www_11_reg[16]  ( .D(n44425), .CP(clk), .Q(reg_www_11[16]) );
  dff_sg \reg_ww_11_reg[15]  ( .D(n44527), .CP(clk), .Q(reg_ww_11[15]) );
  dff_sg \reg_www_11_reg[15]  ( .D(n44424), .CP(clk), .Q(reg_www_11[15]) );
  dff_sg \reg_ww_11_reg[14]  ( .D(n44465), .CP(clk), .Q(reg_ww_11[14]) );
  dff_sg \reg_www_11_reg[14]  ( .D(n44428), .CP(clk), .Q(reg_www_11[14]) );
  dff_sg \reg_ww_11_reg[13]  ( .D(n44464), .CP(clk), .Q(reg_ww_11[13]) );
  dff_sg \reg_www_11_reg[13]  ( .D(n44427), .CP(clk), .Q(reg_www_11[13]) );
  dff_sg \reg_ww_11_reg[12]  ( .D(n44468), .CP(clk), .Q(reg_ww_11[12]) );
  dff_sg \reg_www_11_reg[12]  ( .D(n44435), .CP(clk), .Q(reg_www_11[12]) );
  dff_sg \reg_ww_11_reg[11]  ( .D(n44467), .CP(clk), .Q(reg_ww_11[11]) );
  dff_sg \reg_www_11_reg[11]  ( .D(n44432), .CP(clk), .Q(reg_www_11[11]) );
  dff_sg \reg_ww_11_reg[10]  ( .D(n44459), .CP(clk), .Q(reg_ww_11[10]) );
  dff_sg \reg_www_11_reg[10]  ( .D(n44522), .CP(clk), .Q(reg_www_11[10]) );
  dff_sg \reg_ww_11_reg[9]  ( .D(n44458), .CP(clk), .Q(reg_ww_11[9]) );
  dff_sg \reg_www_11_reg[9]  ( .D(n44521), .CP(clk), .Q(reg_www_11[9]) );
  dff_sg \reg_ww_11_reg[8]  ( .D(n44462), .CP(clk), .Q(reg_ww_11[8]) );
  dff_sg \reg_www_11_reg[8]  ( .D(n44479), .CP(clk), .Q(reg_www_11[8]) );
  dff_sg \reg_ww_11_reg[7]  ( .D(n44461), .CP(clk), .Q(reg_ww_11[7]) );
  dff_sg \reg_www_11_reg[7]  ( .D(n44520), .CP(clk), .Q(reg_www_11[7]) );
  dff_sg \reg_ww_11_reg[6]  ( .D(n44472), .CP(clk), .Q(reg_ww_11[6]) );
  dff_sg \reg_www_11_reg[6]  ( .D(n44466), .CP(clk), .Q(reg_www_11[6]) );
  dff_sg \reg_ww_11_reg[5]  ( .D(n44471), .CP(clk), .Q(reg_ww_11[5]) );
  dff_sg \reg_www_11_reg[5]  ( .D(n44463), .CP(clk), .Q(reg_www_11[5]) );
  dff_sg \reg_ww_11_reg[4]  ( .D(n44475), .CP(clk), .Q(reg_ww_11[4]) );
  dff_sg \reg_www_11_reg[4]  ( .D(n44481), .CP(clk), .Q(reg_www_11[4]) );
  dff_sg \reg_ww_11_reg[3]  ( .D(n44474), .CP(clk), .Q(reg_ww_11[3]) );
  dff_sg \reg_www_11_reg[3]  ( .D(n44480), .CP(clk), .Q(reg_www_11[3]) );
  dff_sg \reg_ww_11_reg[2]  ( .D(n44473), .CP(clk), .Q(reg_ww_11[2]) );
  dff_sg \reg_www_11_reg[2]  ( .D(n44534), .CP(clk), .Q(reg_www_11[2]) );
  dff_sg \reg_ww_11_reg[1]  ( .D(n44470), .CP(clk), .Q(reg_ww_11[1]) );
  dff_sg \reg_www_11_reg[1]  ( .D(n44533), .CP(clk), .Q(reg_www_11[1]) );
  dff_sg \reg_ww_11_reg[0]  ( .D(n44460), .CP(clk), .Q(reg_ww_11[0]) );
  dff_sg \reg_www_11_reg[0]  ( .D(n44523), .CP(clk), .Q(reg_www_11[0]) );
  dff_sg \reg_ww_10_reg[19]  ( .D(n44709), .CP(clk), .Q(reg_ww_10[19]) );
  dff_sg \reg_www_10_reg[19]  ( .D(n44469), .CP(clk), .Q(reg_www_10[19]) );
  dff_sg \reg_ww_10_reg[18]  ( .D(n44701), .CP(clk), .Q(reg_ww_10[18]) );
  dff_sg \reg_www_10_reg[18]  ( .D(n44731), .CP(clk), .Q(reg_www_10[18]) );
  dff_sg \reg_ww_10_reg[17]  ( .D(n44700), .CP(clk), .Q(reg_ww_10[17]) );
  dff_sg \reg_www_10_reg[17]  ( .D(n44730), .CP(clk), .Q(reg_www_10[17]) );
  dff_sg \reg_ww_10_reg[16]  ( .D(n44704), .CP(clk), .Q(reg_ww_10[16]) );
  dff_sg \reg_www_10_reg[16]  ( .D(n44734), .CP(clk), .Q(reg_www_10[16]) );
  dff_sg \reg_ww_10_reg[15]  ( .D(n44703), .CP(clk), .Q(reg_ww_10[15]) );
  dff_sg \reg_www_10_reg[15]  ( .D(n44733), .CP(clk), .Q(reg_www_10[15]) );
  dff_sg \reg_ww_10_reg[14]  ( .D(n44719), .CP(clk), .Q(reg_ww_10[14]) );
  dff_sg \reg_www_10_reg[14]  ( .D(n44725), .CP(clk), .Q(reg_www_10[14]) );
  dff_sg \reg_ww_10_reg[13]  ( .D(n44718), .CP(clk), .Q(reg_ww_10[13]) );
  dff_sg \reg_www_10_reg[13]  ( .D(n44724), .CP(clk), .Q(reg_www_10[13]) );
  dff_sg \reg_ww_10_reg[12]  ( .D(n44722), .CP(clk), .Q(reg_ww_10[12]) );
  dff_sg \reg_www_10_reg[12]  ( .D(n44728), .CP(clk), .Q(reg_www_10[12]) );
  dff_sg \reg_ww_10_reg[11]  ( .D(n44721), .CP(clk), .Q(reg_ww_10[11]) );
  dff_sg \reg_www_10_reg[11]  ( .D(n44727), .CP(clk), .Q(reg_www_10[11]) );
  dff_sg \reg_ww_10_reg[10]  ( .D(n44713), .CP(clk), .Q(reg_ww_10[10]) );
  dff_sg \reg_www_10_reg[10]  ( .D(n44743), .CP(clk), .Q(reg_www_10[10]) );
  dff_sg \reg_ww_10_reg[9]  ( .D(n44712), .CP(clk), .Q(reg_ww_10[9]) );
  dff_sg \reg_www_10_reg[9]  ( .D(n44742), .CP(clk), .Q(reg_www_10[9]) );
  dff_sg \reg_ww_10_reg[8]  ( .D(n44716), .CP(clk), .Q(reg_ww_10[8]) );
  dff_sg \reg_www_10_reg[8]  ( .D(n44746), .CP(clk), .Q(reg_www_10[8]) );
  dff_sg \reg_ww_10_reg[7]  ( .D(n44715), .CP(clk), .Q(reg_ww_10[7]) );
  dff_sg \reg_www_10_reg[7]  ( .D(n44745), .CP(clk), .Q(reg_www_10[7]) );
  dff_sg \reg_ww_10_reg[6]  ( .D(n44779), .CP(clk), .Q(reg_ww_10[6]) );
  dff_sg \reg_www_10_reg[6]  ( .D(n44737), .CP(clk), .Q(reg_www_10[6]) );
  dff_sg \reg_ww_10_reg[5]  ( .D(n44778), .CP(clk), .Q(reg_ww_10[5]) );
  dff_sg \reg_www_10_reg[5]  ( .D(n44736), .CP(clk), .Q(reg_www_10[5]) );
  dff_sg \reg_ww_10_reg[4]  ( .D(n44782), .CP(clk), .Q(reg_ww_10[4]) );
  dff_sg \reg_www_10_reg[4]  ( .D(n44740), .CP(clk), .Q(reg_www_10[4]) );
  dff_sg \reg_ww_10_reg[3]  ( .D(n44781), .CP(clk), .Q(reg_ww_10[3]) );
  dff_sg \reg_www_10_reg[3]  ( .D(n44739), .CP(clk), .Q(reg_www_10[3]) );
  dff_sg \reg_ww_10_reg[2]  ( .D(n44773), .CP(clk), .Q(reg_ww_10[2]) );
  dff_sg \reg_www_10_reg[2]  ( .D(n44707), .CP(clk), .Q(reg_www_10[2]) );
  dff_sg \reg_ww_10_reg[1]  ( .D(n44772), .CP(clk), .Q(reg_ww_10[1]) );
  dff_sg \reg_www_10_reg[1]  ( .D(n44706), .CP(clk), .Q(reg_www_10[1]) );
  dff_sg \reg_ww_10_reg[0]  ( .D(n44776), .CP(clk), .Q(reg_ww_10[0]) );
  dff_sg \reg_www_10_reg[0]  ( .D(n44710), .CP(clk), .Q(reg_www_10[0]) );
  dff_sg \reg_ww_9_reg[19]  ( .D(n44769), .CP(clk), .Q(reg_ww_9[19]) );
  dff_sg \reg_www_9_reg[19]  ( .D(n44775), .CP(clk), .Q(reg_www_9[19]) );
  dff_sg \reg_ww_9_reg[18]  ( .D(n44761), .CP(clk), .Q(reg_ww_9[18]) );
  dff_sg \reg_www_9_reg[18]  ( .D(n44791), .CP(clk), .Q(reg_www_9[18]) );
  dff_sg \reg_ww_9_reg[17]  ( .D(n44760), .CP(clk), .Q(reg_ww_9[17]) );
  dff_sg \reg_www_9_reg[17]  ( .D(n44790), .CP(clk), .Q(reg_www_9[17]) );
  dff_sg \reg_ww_9_reg[16]  ( .D(n44764), .CP(clk), .Q(reg_ww_9[16]) );
  dff_sg \reg_www_9_reg[16]  ( .D(n44794), .CP(clk), .Q(reg_www_9[16]) );
  dff_sg \reg_ww_9_reg[15]  ( .D(n44763), .CP(clk), .Q(reg_ww_9[15]) );
  dff_sg \reg_www_9_reg[15]  ( .D(n44793), .CP(clk), .Q(reg_www_9[15]) );
  dff_sg \reg_ww_9_reg[14]  ( .D(n44575), .CP(clk), .Q(reg_ww_9[14]) );
  dff_sg \reg_www_9_reg[14]  ( .D(n44785), .CP(clk), .Q(reg_www_9[14]) );
  dff_sg \reg_ww_9_reg[13]  ( .D(n44574), .CP(clk), .Q(reg_ww_9[13]) );
  dff_sg \reg_www_9_reg[13]  ( .D(n44784), .CP(clk), .Q(reg_www_9[13]) );
  dff_sg \reg_ww_9_reg[12]  ( .D(n44578), .CP(clk), .Q(reg_ww_9[12]) );
  dff_sg \reg_www_9_reg[12]  ( .D(n44788), .CP(clk), .Q(reg_www_9[12]) );
  dff_sg \reg_ww_9_reg[11]  ( .D(n44577), .CP(clk), .Q(reg_ww_9[11]) );
  dff_sg \reg_www_9_reg[11]  ( .D(n44787), .CP(clk), .Q(reg_www_9[11]) );
  dff_sg \reg_ww_9_reg[10]  ( .D(n44569), .CP(clk), .Q(reg_ww_9[10]) );
  dff_sg \reg_www_9_reg[10]  ( .D(n44755), .CP(clk), .Q(reg_www_9[10]) );
  dff_sg \reg_ww_9_reg[9]  ( .D(n44568), .CP(clk), .Q(reg_ww_9[9]) );
  dff_sg \reg_www_9_reg[9]  ( .D(n44754), .CP(clk), .Q(reg_www_9[9]) );
  dff_sg \reg_ww_9_reg[8]  ( .D(n44572), .CP(clk), .Q(reg_ww_9[8]) );
  dff_sg \reg_www_9_reg[8]  ( .D(n44758), .CP(clk), .Q(reg_www_9[8]) );
  dff_sg \reg_ww_9_reg[7]  ( .D(n44571), .CP(clk), .Q(reg_ww_9[7]) );
  dff_sg \reg_www_9_reg[7]  ( .D(n44757), .CP(clk), .Q(reg_www_9[7]) );
  dff_sg \reg_ww_9_reg[6]  ( .D(n44623), .CP(clk), .Q(reg_ww_9[6]) );
  dff_sg \reg_www_9_reg[6]  ( .D(n44749), .CP(clk), .Q(reg_www_9[6]) );
  dff_sg \reg_ww_9_reg[5]  ( .D(n44622), .CP(clk), .Q(reg_ww_9[5]) );
  dff_sg \reg_www_9_reg[5]  ( .D(n44748), .CP(clk), .Q(reg_www_9[5]) );
  dff_sg \reg_ww_9_reg[4]  ( .D(n44626), .CP(clk), .Q(reg_ww_9[4]) );
  dff_sg \reg_www_9_reg[4]  ( .D(n44752), .CP(clk), .Q(reg_www_9[4]) );
  dff_sg \reg_ww_9_reg[3]  ( .D(n44625), .CP(clk), .Q(reg_ww_9[3]) );
  dff_sg \reg_www_9_reg[3]  ( .D(n44751), .CP(clk), .Q(reg_www_9[3]) );
  dff_sg \reg_ww_9_reg[2]  ( .D(n44629), .CP(clk), .Q(reg_ww_9[2]) );
  dff_sg \reg_www_9_reg[2]  ( .D(n44767), .CP(clk), .Q(reg_www_9[2]) );
  dff_sg \reg_ww_9_reg[1]  ( .D(n44628), .CP(clk), .Q(reg_ww_9[1]) );
  dff_sg \reg_www_9_reg[1]  ( .D(n44766), .CP(clk), .Q(reg_www_9[1]) );
  dff_sg \reg_ww_9_reg[0]  ( .D(n44632), .CP(clk), .Q(reg_ww_9[0]) );
  dff_sg \reg_www_9_reg[0]  ( .D(n44770), .CP(clk), .Q(reg_www_9[0]) );
  dff_sg \reg_ww_8_reg[19]  ( .D(n44631), .CP(clk), .Q(reg_ww_8[19]) );
  dff_sg \reg_www_8_reg[19]  ( .D(n45188), .CP(clk), .Q(reg_www_8[19]) );
  dff_sg \reg_ww_8_reg[18]  ( .D(n45505), .CP(clk), .Q(reg_ww_8[18]) );
  dff_sg \reg_www_8_reg[18]  ( .D(n45185), .CP(clk), .Q(reg_www_8[18]) );
  dff_sg \reg_ww_8_reg[17]  ( .D(n45506), .CP(clk), .Q(reg_ww_8[17]) );
  dff_sg \reg_www_8_reg[17]  ( .D(n45189), .CP(clk), .Q(reg_www_8[17]) );
  dff_sg \reg_ww_8_reg[16]  ( .D(n44369), .CP(clk), .Q(reg_ww_8[16]) );
  dff_sg \reg_www_8_reg[16]  ( .D(n45190), .CP(clk), .Q(reg_www_8[16]) );
  dff_sg \reg_ww_8_reg[15]  ( .D(n44368), .CP(clk), .Q(reg_ww_8[15]) );
  dff_sg \reg_www_8_reg[15]  ( .D(n45422), .CP(clk), .Q(reg_www_8[15]) );
  dff_sg \reg_ww_15_reg[19]  ( .D(n44695), .CP(clk), .Q(reg_ww_15[19]) );
  dff_sg \reg_www_15_reg[19]  ( .D(n44635), .CP(clk), .Q(reg_www_15[19]) );
  dff_sg \reg_ww_15_reg[18]  ( .D(n44694), .CP(clk), .Q(reg_ww_15[18]) );
  dff_sg \reg_www_15_reg[18]  ( .D(n44634), .CP(clk), .Q(reg_www_15[18]) );
  dff_sg \reg_ww_15_reg[17]  ( .D(n44698), .CP(clk), .Q(reg_ww_15[17]) );
  dff_sg \reg_www_15_reg[17]  ( .D(n44638), .CP(clk), .Q(reg_www_15[17]) );
  dff_sg \reg_ww_15_reg[16]  ( .D(n44697), .CP(clk), .Q(reg_ww_15[16]) );
  dff_sg \reg_www_15_reg[16]  ( .D(n44637), .CP(clk), .Q(reg_www_15[16]) );
  dff_sg \reg_ww_15_reg[15]  ( .D(n44689), .CP(clk), .Q(reg_ww_15[15]) );
  dff_sg \reg_www_15_reg[15]  ( .D(n44647), .CP(clk), .Q(reg_www_15[15]) );
  dff_sg \reg_ww_15_reg[14]  ( .D(n44688), .CP(clk), .Q(reg_ww_15[14]) );
  dff_sg \reg_www_15_reg[14]  ( .D(n44646), .CP(clk), .Q(reg_www_15[14]) );
  dff_sg \reg_ww_15_reg[13]  ( .D(n44692), .CP(clk), .Q(reg_ww_15[13]) );
  dff_sg \reg_www_15_reg[13]  ( .D(n44650), .CP(clk), .Q(reg_www_15[13]) );
  dff_sg \reg_ww_15_reg[12]  ( .D(n44691), .CP(clk), .Q(reg_ww_15[12]) );
  dff_sg \reg_www_15_reg[12]  ( .D(n44649), .CP(clk), .Q(reg_www_15[12]) );
  dff_sg \reg_ww_15_reg[11]  ( .D(n44659), .CP(clk), .Q(reg_ww_15[11]) );
  dff_sg \reg_www_15_reg[11]  ( .D(n44641), .CP(clk), .Q(reg_www_15[11]) );
  dff_sg \reg_ww_15_reg[10]  ( .D(n44658), .CP(clk), .Q(reg_ww_15[10]) );
  dff_sg \reg_www_15_reg[10]  ( .D(n44640), .CP(clk), .Q(reg_www_15[10]) );
  dff_sg \reg_ww_15_reg[9]  ( .D(n44662), .CP(clk), .Q(reg_ww_15[9]) );
  dff_sg \reg_www_15_reg[9]  ( .D(n44644), .CP(clk), .Q(reg_www_15[9]) );
  dff_sg \reg_ww_15_reg[8]  ( .D(n44661), .CP(clk), .Q(reg_ww_15[8]) );
  dff_sg \reg_www_15_reg[8]  ( .D(n44643), .CP(clk), .Q(reg_www_15[8]) );
  dff_sg \reg_ww_15_reg[7]  ( .D(n44653), .CP(clk), .Q(reg_ww_15[7]) );
  dff_sg \reg_www_15_reg[7]  ( .D(n44683), .CP(clk), .Q(reg_www_15[7]) );
  dff_sg \reg_ww_15_reg[6]  ( .D(n44652), .CP(clk), .Q(reg_ww_15[6]) );
  dff_sg \reg_www_15_reg[6]  ( .D(n44682), .CP(clk), .Q(reg_www_15[6]) );
  dff_sg \reg_ww_15_reg[5]  ( .D(n44656), .CP(clk), .Q(reg_ww_15[5]) );
  dff_sg \reg_www_15_reg[5]  ( .D(n44686), .CP(clk), .Q(reg_www_15[5]) );
  dff_sg \reg_ww_15_reg[4]  ( .D(n44655), .CP(clk), .Q(reg_ww_15[4]) );
  dff_sg \reg_www_15_reg[4]  ( .D(n44685), .CP(clk), .Q(reg_www_15[4]) );
  dff_sg \reg_ww_15_reg[3]  ( .D(n44671), .CP(clk), .Q(reg_ww_15[3]) );
  dff_sg \reg_www_15_reg[3]  ( .D(n44677), .CP(clk), .Q(reg_www_15[3]) );
  dff_sg \reg_ww_15_reg[2]  ( .D(n44670), .CP(clk), .Q(reg_ww_15[2]) );
  dff_sg \reg_www_15_reg[2]  ( .D(n44676), .CP(clk), .Q(reg_www_15[2]) );
  dff_sg \reg_ww_15_reg[1]  ( .D(n44674), .CP(clk), .Q(reg_ww_15[1]) );
  dff_sg \reg_www_15_reg[1]  ( .D(n44680), .CP(clk), .Q(reg_www_15[1]) );
  dff_sg \reg_ww_15_reg[0]  ( .D(n44673), .CP(clk), .Q(reg_ww_15[0]) );
  dff_sg \reg_www_15_reg[0]  ( .D(n44679), .CP(clk), .Q(reg_www_15[0]) );
  dff_sg \reg_ww_14_reg[19]  ( .D(n45109), .CP(clk), .Q(reg_ww_14[19]) );
  dff_sg \reg_www_14_reg[19]  ( .D(n44665), .CP(clk), .Q(reg_www_14[19]) );
  dff_sg \reg_ww_14_reg[18]  ( .D(n45108), .CP(clk), .Q(reg_ww_14[18]) );
  dff_sg \reg_www_14_reg[18]  ( .D(n44664), .CP(clk), .Q(reg_www_14[18]) );
  dff_sg \reg_ww_14_reg[17]  ( .D(n45112), .CP(clk), .Q(reg_ww_14[17]) );
  dff_sg \reg_www_14_reg[17]  ( .D(n44668), .CP(clk), .Q(reg_www_14[17]) );
  dff_sg \reg_ww_14_reg[16]  ( .D(n45111), .CP(clk), .Q(reg_ww_14[16]) );
  dff_sg \reg_www_14_reg[16]  ( .D(n44667), .CP(clk), .Q(reg_www_14[16]) );
  dff_sg \reg_ww_14_reg[15]  ( .D(n45103), .CP(clk), .Q(reg_ww_14[15]) );
  dff_sg \reg_www_14_reg[15]  ( .D(n45128), .CP(clk), .Q(reg_www_14[15]) );
  dff_sg \reg_ww_14_reg[14]  ( .D(n45102), .CP(clk), .Q(reg_ww_14[14]) );
  dff_sg \reg_www_14_reg[14]  ( .D(n45127), .CP(clk), .Q(reg_www_14[14]) );
  dff_sg \reg_ww_14_reg[13]  ( .D(n45106), .CP(clk), .Q(reg_ww_14[13]) );
  dff_sg \reg_www_14_reg[13]  ( .D(n45131), .CP(clk), .Q(reg_www_14[13]) );
  dff_sg \reg_ww_14_reg[12]  ( .D(n45105), .CP(clk), .Q(reg_ww_14[12]) );
  dff_sg \reg_www_14_reg[12]  ( .D(n45130), .CP(clk), .Q(reg_www_14[12]) );
  dff_sg \reg_ww_14_reg[11]  ( .D(n45129), .CP(clk), .Q(reg_ww_14[11]) );
  dff_sg \reg_www_14_reg[11]  ( .D(n45122), .CP(clk), .Q(reg_www_14[11]) );
  dff_sg \reg_ww_14_reg[10]  ( .D(n45126), .CP(clk), .Q(reg_ww_14[10]) );
  dff_sg \reg_www_14_reg[10]  ( .D(n45121), .CP(clk), .Q(reg_www_14[10]) );
  dff_sg \reg_ww_14_reg[9]  ( .D(n45120), .CP(clk), .Q(reg_ww_14[9]) );
  dff_sg \reg_www_14_reg[9]  ( .D(n45125), .CP(clk), .Q(reg_www_14[9]) );
  dff_sg \reg_ww_14_reg[8]  ( .D(n45113), .CP(clk), .Q(reg_ww_14[8]) );
  dff_sg \reg_www_14_reg[8]  ( .D(n45124), .CP(clk), .Q(reg_www_14[8]) );
  dff_sg \reg_ww_14_reg[7]  ( .D(n45116), .CP(clk), .Q(reg_ww_14[7]) );
  dff_sg \reg_www_14_reg[7]  ( .D(n45135), .CP(clk), .Q(reg_www_14[7]) );
  dff_sg \reg_ww_14_reg[6]  ( .D(n45115), .CP(clk), .Q(reg_ww_14[6]) );
  dff_sg \reg_www_14_reg[6]  ( .D(n45134), .CP(clk), .Q(reg_www_14[6]) );
  dff_sg \reg_ww_14_reg[5]  ( .D(n45119), .CP(clk), .Q(reg_ww_14[5]) );
  dff_sg \reg_www_14_reg[5]  ( .D(n45138), .CP(clk), .Q(reg_www_14[5]) );
  dff_sg \reg_ww_14_reg[4]  ( .D(n45118), .CP(clk), .Q(reg_ww_14[4]) );
  dff_sg \reg_www_14_reg[4]  ( .D(n45137), .CP(clk), .Q(reg_www_14[4]) );
  dff_sg \reg_ww_14_reg[3]  ( .D(n45145), .CP(clk), .Q(reg_ww_14[3]) );
  dff_sg \reg_www_14_reg[3]  ( .D(n45136), .CP(clk), .Q(reg_www_14[3]) );
  dff_sg \reg_ww_14_reg[2]  ( .D(n45514), .CP(clk), .Q(reg_ww_14[2]) );
  dff_sg \reg_www_14_reg[2]  ( .D(n45133), .CP(clk), .Q(reg_www_14[2]) );
  dff_sg \reg_ww_14_reg[1]  ( .D(n45509), .CP(clk), .Q(reg_ww_14[1]) );
  dff_sg \reg_www_14_reg[1]  ( .D(n45123), .CP(clk), .Q(reg_www_14[1]) );
  dff_sg \reg_ww_14_reg[0]  ( .D(n45510), .CP(clk), .Q(reg_ww_14[0]) );
  dff_sg \reg_www_14_reg[0]  ( .D(n45132), .CP(clk), .Q(reg_www_14[0]) );
  dff_sg \reg_ww_13_reg[19]  ( .D(n45147), .CP(clk), .Q(reg_ww_13[19]) );
  dff_sg \reg_www_13_reg[19]  ( .D(n44562), .CP(clk), .Q(reg_www_13[19]) );
  dff_sg \reg_ww_13_reg[18]  ( .D(n45146), .CP(clk), .Q(reg_ww_13[18]) );
  dff_sg \reg_www_13_reg[18]  ( .D(n44566), .CP(clk), .Q(reg_www_13[18]) );
  dff_sg \reg_ww_13_reg[17]  ( .D(n45511), .CP(clk), .Q(reg_ww_13[17]) );
  dff_sg \reg_www_13_reg[17]  ( .D(n44565), .CP(clk), .Q(reg_www_13[17]) );
  dff_sg \reg_ww_13_reg[16]  ( .D(n45508), .CP(clk), .Q(reg_ww_13[16]) );
  dff_sg \reg_www_13_reg[16]  ( .D(n44544), .CP(clk), .Q(reg_www_13[16]) );
  dff_sg \reg_ww_13_reg[15]  ( .D(n45512), .CP(clk), .Q(reg_ww_13[15]) );
  dff_sg \reg_www_13_reg[15]  ( .D(n44543), .CP(clk), .Q(reg_www_13[15]) );
  dff_sg \reg_ww_13_reg[14]  ( .D(n45513), .CP(clk), .Q(reg_ww_13[14]) );
  dff_sg \reg_www_13_reg[14]  ( .D(n44539), .CP(clk), .Q(reg_www_13[14]) );
  dff_sg \mask_0/reg_ii_mask_reg[0]  ( .D(n44174), .CP(clk), .Q(
        \mask_0/reg_ii_mask [0]) );
  dff_sg \mask_0/reg_ii_mask_reg[1]  ( .D(n44175), .CP(clk), .Q(
        \mask_0/reg_ii_mask [1]) );
  dff_sg \mask_0/reg_ii_mask_reg[2]  ( .D(n44171), .CP(clk), .Q(
        \mask_0/reg_ii_mask [2]) );
  dff_sg \mask_0/reg_ii_mask_reg[3]  ( .D(n44172), .CP(clk), .Q(
        \mask_0/reg_ii_mask [3]) );
  dff_sg \mask_0/reg_ii_mask_reg[4]  ( .D(n44180), .CP(clk), .Q(
        \mask_0/reg_ii_mask [4]) );
  dff_sg \mask_0/reg_ii_mask_reg[5]  ( .D(n44181), .CP(clk), .Q(
        \mask_0/reg_ii_mask [5]) );
  dff_sg \mask_0/reg_ii_mask_reg[6]  ( .D(n44177), .CP(clk), .Q(
        \mask_0/reg_ii_mask [6]) );
  dff_sg \mask_0/reg_ii_mask_reg[7]  ( .D(n44178), .CP(clk), .Q(
        \mask_0/reg_ii_mask [7]) );
  dff_sg \mask_0/reg_ii_mask_reg[8]  ( .D(n44162), .CP(clk), .Q(
        \mask_0/reg_ii_mask [8]) );
  dff_sg \mask_0/reg_ii_mask_reg[9]  ( .D(n44163), .CP(clk), .Q(
        \mask_0/reg_ii_mask [9]) );
  dff_sg \mask_0/reg_ii_mask_reg[10]  ( .D(n44159), .CP(clk), .Q(
        \mask_0/reg_ii_mask [10]) );
  dff_sg \mask_0/reg_ii_mask_reg[11]  ( .D(n44160), .CP(clk), .Q(
        \mask_0/reg_ii_mask [11]) );
  dff_sg \mask_0/reg_ii_mask_reg[12]  ( .D(n44168), .CP(clk), .Q(
        \mask_0/reg_ii_mask [12]) );
  dff_sg \mask_0/reg_ii_mask_reg[13]  ( .D(n44169), .CP(clk), .Q(
        \mask_0/reg_ii_mask [13]) );
  dff_sg \mask_0/reg_ii_mask_reg[14]  ( .D(n44165), .CP(clk), .Q(
        \mask_0/reg_ii_mask [14]) );
  dff_sg \mask_0/reg_ii_mask_reg[15]  ( .D(n44166), .CP(clk), .Q(
        \mask_0/reg_ii_mask [15]) );
  dff_sg \mask_0/reg_ii_mask_reg[16]  ( .D(n44198), .CP(clk), .Q(
        \mask_0/reg_ii_mask [16]) );
  dff_sg \mask_0/reg_ii_mask_reg[17]  ( .D(n44199), .CP(clk), .Q(
        \mask_0/reg_ii_mask [17]) );
  dff_sg \mask_0/reg_ii_mask_reg[18]  ( .D(n44195), .CP(clk), .Q(
        \mask_0/reg_ii_mask [18]) );
  dff_sg \mask_0/reg_ii_mask_reg[19]  ( .D(n44196), .CP(clk), .Q(
        \mask_0/reg_ii_mask [19]) );
  dff_sg \mask_0/reg_ii_mask_reg[20]  ( .D(n44204), .CP(clk), .Q(
        \mask_0/reg_ii_mask [20]) );
  dff_sg \mask_0/reg_ii_mask_reg[21]  ( .D(n44205), .CP(clk), .Q(
        \mask_0/reg_ii_mask [21]) );
  dff_sg \mask_0/reg_ii_mask_reg[22]  ( .D(n44201), .CP(clk), .Q(
        \mask_0/reg_ii_mask [22]) );
  dff_sg \mask_0/reg_ii_mask_reg[23]  ( .D(n44202), .CP(clk), .Q(
        \mask_0/reg_ii_mask [23]) );
  dff_sg \mask_0/reg_ii_mask_reg[24]  ( .D(n44186), .CP(clk), .Q(
        \mask_0/reg_ii_mask [24]) );
  dff_sg \mask_0/reg_ii_mask_reg[25]  ( .D(n44187), .CP(clk), .Q(
        \mask_0/reg_ii_mask [25]) );
  dff_sg \mask_0/reg_ii_mask_reg[26]  ( .D(n44183), .CP(clk), .Q(
        \mask_0/reg_ii_mask [26]) );
  dff_sg \mask_0/reg_ii_mask_reg[27]  ( .D(n44184), .CP(clk), .Q(
        \mask_0/reg_ii_mask [27]) );
  dff_sg \mask_0/reg_ii_mask_reg[28]  ( .D(n44192), .CP(clk), .Q(
        \mask_0/reg_ii_mask [28]) );
  dff_sg \mask_0/reg_ii_mask_reg[29]  ( .D(n44193), .CP(clk), .Q(
        \mask_0/reg_ii_mask [29]) );
  dff_sg \mask_0/reg_ii_mask_reg[30]  ( .D(n44189), .CP(clk), .Q(
        \mask_0/reg_ii_mask [30]) );
  dff_sg \mask_0/reg_ii_mask_reg[31]  ( .D(n44190), .CP(clk), .Q(
        \mask_0/reg_ii_mask [31]) );
  dff_sg \mask_0/reg_ww_mask_reg[0]  ( .D(n44126), .CP(clk), .Q(
        \mask_0/reg_ww_mask [0]) );
  dff_sg \mask_0/reg_ww_mask_reg[1]  ( .D(n44127), .CP(clk), .Q(
        \mask_0/reg_ww_mask [1]) );
  dff_sg \mask_0/reg_ww_mask_reg[2]  ( .D(n44123), .CP(clk), .Q(
        \mask_0/reg_ww_mask [2]) );
  dff_sg \mask_0/reg_ww_mask_reg[3]  ( .D(n44124), .CP(clk), .Q(
        \mask_0/reg_ww_mask [3]) );
  dff_sg \mask_0/reg_ww_mask_reg[4]  ( .D(n44132), .CP(clk), .Q(
        \mask_0/reg_ww_mask [4]) );
  dff_sg \mask_0/reg_ww_mask_reg[5]  ( .D(n44133), .CP(clk), .Q(
        \mask_0/reg_ww_mask [5]) );
  dff_sg \mask_0/reg_ww_mask_reg[6]  ( .D(n44129), .CP(clk), .Q(
        \mask_0/reg_ww_mask [6]) );
  dff_sg \mask_0/reg_ww_mask_reg[7]  ( .D(n44130), .CP(clk), .Q(
        \mask_0/reg_ww_mask [7]) );
  dff_sg \mask_0/reg_ww_mask_reg[8]  ( .D(n44114), .CP(clk), .Q(
        \mask_0/reg_ww_mask [8]) );
  dff_sg \mask_0/reg_ww_mask_reg[9]  ( .D(n44115), .CP(clk), .Q(
        \mask_0/reg_ww_mask [9]) );
  dff_sg \mask_0/reg_ww_mask_reg[10]  ( .D(n44111), .CP(clk), .Q(
        \mask_0/reg_ww_mask [10]) );
  dff_sg \mask_0/reg_ww_mask_reg[11]  ( .D(n44112), .CP(clk), .Q(
        \mask_0/reg_ww_mask [11]) );
  dff_sg \mask_0/reg_ww_mask_reg[12]  ( .D(n44120), .CP(clk), .Q(
        \mask_0/reg_ww_mask [12]) );
  dff_sg \mask_0/reg_ww_mask_reg[13]  ( .D(n44121), .CP(clk), .Q(
        \mask_0/reg_ww_mask [13]) );
  dff_sg \mask_0/reg_ww_mask_reg[14]  ( .D(n44117), .CP(clk), .Q(
        \mask_0/reg_ww_mask [14]) );
  dff_sg \mask_0/reg_ww_mask_reg[15]  ( .D(n44118), .CP(clk), .Q(
        \mask_0/reg_ww_mask [15]) );
  dff_sg \mask_0/reg_ww_mask_reg[16]  ( .D(n44150), .CP(clk), .Q(
        \mask_0/reg_ww_mask [16]) );
  dff_sg \mask_0/reg_ww_mask_reg[17]  ( .D(n44151), .CP(clk), .Q(
        \mask_0/reg_ww_mask [17]) );
  dff_sg \mask_0/reg_ww_mask_reg[18]  ( .D(n44147), .CP(clk), .Q(
        \mask_0/reg_ww_mask [18]) );
  dff_sg \mask_0/reg_ww_mask_reg[19]  ( .D(n44148), .CP(clk), .Q(
        \mask_0/reg_ww_mask [19]) );
  dff_sg \mask_0/reg_ww_mask_reg[20]  ( .D(n44156), .CP(clk), .Q(
        \mask_0/reg_ww_mask [20]) );
  dff_sg \mask_0/reg_ww_mask_reg[21]  ( .D(n44157), .CP(clk), .Q(
        \mask_0/reg_ww_mask [21]) );
  dff_sg \mask_0/reg_ww_mask_reg[22]  ( .D(n44153), .CP(clk), .Q(
        \mask_0/reg_ww_mask [22]) );
  dff_sg \mask_0/reg_ww_mask_reg[23]  ( .D(n44154), .CP(clk), .Q(
        \mask_0/reg_ww_mask [23]) );
  dff_sg \mask_0/reg_ww_mask_reg[24]  ( .D(n44138), .CP(clk), .Q(
        \mask_0/reg_ww_mask [24]) );
  dff_sg \mask_0/reg_ww_mask_reg[25]  ( .D(n44139), .CP(clk), .Q(
        \mask_0/reg_ww_mask [25]) );
  dff_sg \mask_0/reg_ww_mask_reg[26]  ( .D(n44135), .CP(clk), .Q(
        \mask_0/reg_ww_mask [26]) );
  dff_sg \mask_0/reg_ww_mask_reg[27]  ( .D(n44136), .CP(clk), .Q(
        \mask_0/reg_ww_mask [27]) );
  dff_sg \mask_0/reg_ww_mask_reg[28]  ( .D(n44144), .CP(clk), .Q(
        \mask_0/reg_ww_mask [28]) );
  dff_sg \mask_0/reg_ww_mask_reg[29]  ( .D(n44145), .CP(clk), .Q(
        \mask_0/reg_ww_mask [29]) );
  dff_sg \mask_0/reg_ww_mask_reg[30]  ( .D(n44141), .CP(clk), .Q(
        \mask_0/reg_ww_mask [30]) );
  dff_sg \mask_0/reg_ww_mask_reg[31]  ( .D(n44142), .CP(clk), .Q(
        \mask_0/reg_ww_mask [31]) );
  dff_sg \mask_0/reg_o_mask_reg[0]  ( .D(n44122), .CP(clk), .Q(n69263) );
  dff_sg \mask_0/reg_o_mask_reg[1]  ( .D(n44197), .CP(clk), .Q(n69262) );
  dff_sg \mask_0/reg_o_mask_reg[2]  ( .D(n44134), .CP(clk), .Q(n69261) );
  dff_sg \mask_0/reg_o_mask_reg[3]  ( .D(n44131), .CP(clk), .Q(n69260) );
  dff_sg \mask_0/reg_o_mask_reg[4]  ( .D(n44125), .CP(clk), .Q(n69259) );
  dff_sg \mask_0/reg_o_mask_reg[5]  ( .D(n44128), .CP(clk), .Q(n69258) );
  dff_sg \mask_0/reg_o_mask_reg[6]  ( .D(n44137), .CP(clk), .Q(n69257) );
  dff_sg \mask_0/reg_o_mask_reg[7]  ( .D(n44140), .CP(clk), .Q(n69256) );
  dff_sg \mask_0/reg_o_mask_reg[8]  ( .D(n44158), .CP(clk), .Q(n69255) );
  dff_sg \mask_0/reg_o_mask_reg[9]  ( .D(n44164), .CP(clk), .Q(n69254) );
  dff_sg \mask_0/reg_o_mask_reg[10]  ( .D(n44155), .CP(clk), .Q(n69253) );
  dff_sg \mask_0/reg_o_mask_reg[11]  ( .D(n44152), .CP(clk), .Q(n69252) );
  dff_sg \mask_0/reg_o_mask_reg[12]  ( .D(n44146), .CP(clk), .Q(n69251) );
  dff_sg \mask_0/reg_o_mask_reg[13]  ( .D(n44149), .CP(clk), .Q(n69250) );
  dff_sg \mask_0/reg_o_mask_reg[14]  ( .D(n44161), .CP(clk), .Q(n69249) );
  dff_sg \mask_0/reg_o_mask_reg[15]  ( .D(n44173), .CP(clk), .Q(n69248) );
  dff_sg \mask_0/reg_o_mask_reg[16]  ( .D(n44194), .CP(clk), .Q(n69247) );
  dff_sg \mask_0/reg_o_mask_reg[17]  ( .D(n44143), .CP(clk), .Q(n69246) );
  dff_sg \mask_0/reg_o_mask_reg[18]  ( .D(n44185), .CP(clk), .Q(n69245) );
  dff_sg \mask_0/reg_o_mask_reg[19]  ( .D(n44182), .CP(clk), .Q(n69244) );
  dff_sg \mask_0/reg_o_mask_reg[20]  ( .D(n44176), .CP(clk), .Q(n69243) );
  dff_sg \mask_0/reg_o_mask_reg[21]  ( .D(n44179), .CP(clk), .Q(n69242) );
  dff_sg \mask_0/reg_o_mask_reg[22]  ( .D(n44188), .CP(clk), .Q(n69241) );
  dff_sg \mask_0/reg_o_mask_reg[23]  ( .D(n44191), .CP(clk), .Q(n69240) );
  dff_sg \mask_0/reg_o_mask_reg[24]  ( .D(n44167), .CP(clk), .Q(n69239) );
  dff_sg \mask_0/reg_o_mask_reg[25]  ( .D(n44170), .CP(clk), .Q(n69238) );
  dff_sg \mask_0/reg_o_mask_reg[26]  ( .D(n44200), .CP(clk), .Q(n69237) );
  dff_sg \mask_0/reg_o_mask_reg[27]  ( .D(n44203), .CP(clk), .Q(n69236) );
  dff_sg \mask_0/reg_o_mask_reg[28]  ( .D(n44110), .CP(clk), .Q(n69235) );
  dff_sg \mask_0/reg_o_mask_reg[29]  ( .D(n44113), .CP(clk), .Q(n69234) );
  dff_sg \mask_0/reg_o_mask_reg[30]  ( .D(n44116), .CP(clk), .Q(n69233) );
  dff_sg \mask_0/reg_o_mask_reg[31]  ( .D(n44119), .CP(clk), .Q(n69232) );
  dff_sg \mask_0/reg_i_mask_reg[0]  ( .D(n44234), .CP(clk), .Q(
        \mask_0/reg_i_mask [0]) );
  dff_sg \mask_0/reg_i_mask_reg[1]  ( .D(n44233), .CP(clk), .Q(
        \mask_0/reg_i_mask [1]) );
  dff_sg \mask_0/reg_i_mask_reg[2]  ( .D(n44232), .CP(clk), .Q(
        \mask_0/reg_i_mask [2]) );
  dff_sg \mask_0/reg_i_mask_reg[3]  ( .D(n44206), .CP(clk), .Q(
        \mask_0/reg_i_mask [3]) );
  dff_sg \mask_0/reg_i_mask_reg[4]  ( .D(n44228), .CP(clk), .Q(
        \mask_0/reg_i_mask [4]) );
  dff_sg \mask_0/reg_i_mask_reg[5]  ( .D(n44227), .CP(clk), .Q(
        \mask_0/reg_i_mask [5]) );
  dff_sg \mask_0/reg_i_mask_reg[6]  ( .D(n44231), .CP(clk), .Q(
        \mask_0/reg_i_mask [6]) );
  dff_sg \mask_0/reg_i_mask_reg[7]  ( .D(n44230), .CP(clk), .Q(
        \mask_0/reg_i_mask [7]) );
  dff_sg \mask_0/reg_i_mask_reg[8]  ( .D(n44238), .CP(clk), .Q(
        \mask_0/reg_i_mask [8]) );
  dff_sg \mask_0/reg_i_mask_reg[9]  ( .D(n44237), .CP(clk), .Q(
        \mask_0/reg_i_mask [9]) );
  dff_sg \mask_0/reg_i_mask_reg[10]  ( .D(n44241), .CP(clk), .Q(
        \mask_0/reg_i_mask [10]) );
  dff_sg \mask_0/reg_i_mask_reg[11]  ( .D(n44240), .CP(clk), .Q(
        \mask_0/reg_i_mask [11]) );
  dff_sg \mask_0/reg_i_mask_reg[12]  ( .D(n44235), .CP(clk), .Q(
        \mask_0/reg_i_mask [12]) );
  dff_sg \mask_0/reg_i_mask_reg[13]  ( .D(n44239), .CP(clk), .Q(
        \mask_0/reg_i_mask [13]) );
  dff_sg \mask_0/reg_i_mask_reg[14]  ( .D(n44229), .CP(clk), .Q(
        \mask_0/reg_i_mask [14]) );
  dff_sg \mask_0/reg_i_mask_reg[15]  ( .D(n44226), .CP(clk), .Q(
        \mask_0/reg_i_mask [15]) );
  dff_sg \mask_0/reg_i_mask_reg[16]  ( .D(n44215), .CP(clk), .Q(
        \mask_0/reg_i_mask [16]) );
  dff_sg \mask_0/reg_i_mask_reg[17]  ( .D(n44214), .CP(clk), .Q(
        \mask_0/reg_i_mask [17]) );
  dff_sg \mask_0/reg_i_mask_reg[18]  ( .D(n44218), .CP(clk), .Q(
        \mask_0/reg_i_mask [18]) );
  dff_sg \mask_0/reg_i_mask_reg[19]  ( .D(n44217), .CP(clk), .Q(
        \mask_0/reg_i_mask [19]) );
  dff_sg \mask_0/reg_i_mask_reg[20]  ( .D(n44209), .CP(clk), .Q(
        \mask_0/reg_i_mask [20]) );
  dff_sg \mask_0/reg_i_mask_reg[21]  ( .D(n44208), .CP(clk), .Q(
        \mask_0/reg_i_mask [21]) );
  dff_sg \mask_0/reg_i_mask_reg[22]  ( .D(n44212), .CP(clk), .Q(
        \mask_0/reg_i_mask [22]) );
  dff_sg \mask_0/reg_i_mask_reg[23]  ( .D(n44211), .CP(clk), .Q(
        \mask_0/reg_i_mask [23]) );
  dff_sg \mask_0/reg_i_mask_reg[24]  ( .D(n44222), .CP(clk), .Q(
        \mask_0/reg_i_mask [24]) );
  dff_sg \mask_0/reg_i_mask_reg[25]  ( .D(n44221), .CP(clk), .Q(
        \mask_0/reg_i_mask [25]) );
  dff_sg \mask_0/reg_i_mask_reg[26]  ( .D(n44225), .CP(clk), .Q(
        \mask_0/reg_i_mask [26]) );
  dff_sg \mask_0/reg_i_mask_reg[27]  ( .D(n44224), .CP(clk), .Q(
        \mask_0/reg_i_mask [27]) );
  dff_sg \mask_0/reg_i_mask_reg[28]  ( .D(n44219), .CP(clk), .Q(
        \mask_0/reg_i_mask [28]) );
  dff_sg \mask_0/reg_i_mask_reg[29]  ( .D(n44223), .CP(clk), .Q(
        \mask_0/reg_i_mask [29]) );
  dff_sg \mask_0/reg_i_mask_reg[30]  ( .D(n44236), .CP(clk), .Q(
        \mask_0/reg_i_mask [30]) );
  dff_sg \mask_0/reg_i_mask_reg[31]  ( .D(n44220), .CP(clk), .Q(
        \mask_0/reg_i_mask [31]) );
  dff_sg \mask_0/reg_w_mask_reg[0]  ( .D(n44216), .CP(clk), .Q(
        \mask_0/reg_w_mask [0]) );
  dff_sg \mask_0/reg_w_mask_reg[1]  ( .D(n44213), .CP(clk), .Q(
        \mask_0/reg_w_mask [1]) );
  dff_sg \mask_0/reg_w_mask_reg[2]  ( .D(n44210), .CP(clk), .Q(
        \mask_0/reg_w_mask [2]) );
  dff_sg \mask_0/reg_w_mask_reg[3]  ( .D(n44207), .CP(clk), .Q(
        \mask_0/reg_w_mask [3]) );
  dff_sg \mask_0/reg_w_mask_reg[4]  ( .D(n44259), .CP(clk), .Q(
        \mask_0/reg_w_mask [4]) );
  dff_sg \mask_0/reg_w_mask_reg[5]  ( .D(n44258), .CP(clk), .Q(
        \mask_0/reg_w_mask [5]) );
  dff_sg \mask_0/reg_w_mask_reg[6]  ( .D(n44262), .CP(clk), .Q(
        \mask_0/reg_w_mask [6]) );
  dff_sg \mask_0/reg_w_mask_reg[7]  ( .D(n44261), .CP(clk), .Q(
        \mask_0/reg_w_mask [7]) );
  dff_sg \mask_0/reg_w_mask_reg[8]  ( .D(n44266), .CP(clk), .Q(
        \mask_0/reg_w_mask [8]) );
  dff_sg \mask_0/reg_w_mask_reg[9]  ( .D(n44265), .CP(clk), .Q(
        \mask_0/reg_w_mask [9]) );
  dff_sg \mask_0/reg_w_mask_reg[10]  ( .D(n44269), .CP(clk), .Q(
        \mask_0/reg_w_mask [10]) );
  dff_sg \mask_0/reg_w_mask_reg[11]  ( .D(n44268), .CP(clk), .Q(
        \mask_0/reg_w_mask [11]) );
  dff_sg \mask_0/reg_w_mask_reg[12]  ( .D(n44263), .CP(clk), .Q(
        \mask_0/reg_w_mask [12]) );
  dff_sg \mask_0/reg_w_mask_reg[13]  ( .D(n44267), .CP(clk), .Q(
        \mask_0/reg_w_mask [13]) );
  dff_sg \mask_0/reg_w_mask_reg[14]  ( .D(n44256), .CP(clk), .Q(
        \mask_0/reg_w_mask [14]) );
  dff_sg \mask_0/reg_w_mask_reg[15]  ( .D(n44264), .CP(clk), .Q(
        \mask_0/reg_w_mask [15]) );
  dff_sg \mask_0/reg_w_mask_reg[16]  ( .D(n44245), .CP(clk), .Q(
        \mask_0/reg_w_mask [16]) );
  dff_sg \mask_0/reg_w_mask_reg[17]  ( .D(n44244), .CP(clk), .Q(
        \mask_0/reg_w_mask [17]) );
  dff_sg \mask_0/reg_w_mask_reg[18]  ( .D(n44248), .CP(clk), .Q(
        \mask_0/reg_w_mask [18]) );
  dff_sg \mask_0/reg_w_mask_reg[19]  ( .D(n44247), .CP(clk), .Q(
        \mask_0/reg_w_mask [19]) );
  dff_sg \mask_0/reg_w_mask_reg[20]  ( .D(n44242), .CP(clk), .Q(
        \mask_0/reg_w_mask [20]) );
  dff_sg \mask_0/reg_w_mask_reg[21]  ( .D(n44246), .CP(clk), .Q(
        \mask_0/reg_w_mask [21]) );
  dff_sg \mask_0/reg_w_mask_reg[22]  ( .D(n44260), .CP(clk), .Q(
        \mask_0/reg_w_mask [22]) );
  dff_sg \mask_0/reg_w_mask_reg[23]  ( .D(n44243), .CP(clk), .Q(
        \mask_0/reg_w_mask [23]) );
  dff_sg \mask_0/reg_w_mask_reg[24]  ( .D(n44252), .CP(clk), .Q(
        \mask_0/reg_w_mask [24]) );
  dff_sg \mask_0/reg_w_mask_reg[25]  ( .D(n44251), .CP(clk), .Q(
        \mask_0/reg_w_mask [25]) );
  dff_sg \mask_0/reg_w_mask_reg[26]  ( .D(n44255), .CP(clk), .Q(
        \mask_0/reg_w_mask [26]) );
  dff_sg \mask_0/reg_w_mask_reg[27]  ( .D(n44254), .CP(clk), .Q(
        \mask_0/reg_w_mask [27]) );
  dff_sg \mask_0/reg_w_mask_reg[28]  ( .D(n44249), .CP(clk), .Q(
        \mask_0/reg_w_mask [28]) );
  dff_sg \mask_0/reg_w_mask_reg[29]  ( .D(n44253), .CP(clk), .Q(
        \mask_0/reg_w_mask [29]) );
  dff_sg \mask_0/reg_w_mask_reg[30]  ( .D(n44257), .CP(clk), .Q(
        \mask_0/reg_w_mask [30]) );
  dff_sg \mask_0/reg_w_mask_reg[31]  ( .D(n44250), .CP(clk), .Q(
        \mask_0/reg_w_mask [31]) );
  dff_sg \mask_0/state_reg[0]  ( .D(n44271), .CP(clk), .Q(\mask_0/n1655 ) );
  dff_sg \mask_0/state_reg[1]  ( .D(n44270), .CP(clk), .Q(\mask_0/n1654 ) );
  dff_sg \mask_0/counter_reg[1]  ( .D(n46194), .CP(clk), .Q(
        \mask_0/counter [1]) );
  dff_sg \mask_0/counter_reg[0]  ( .D(n46195), .CP(clk), .Q(
        \mask_0/counter [0]) );
  dff_sg \filter_0/ow_0_reg[0]  ( .D(n43368), .CP(clk), .Q(\filter_0/n17648 )
         );
  dff_sg \filter_0/ow_0_reg[1]  ( .D(n43367), .CP(clk), .Q(\filter_0/n17647 )
         );
  dff_sg \filter_0/ow_0_reg[2]  ( .D(n43366), .CP(clk), .Q(\filter_0/n17646 )
         );
  dff_sg \filter_0/ow_0_reg[3]  ( .D(n43357), .CP(clk), .Q(\filter_0/n17645 )
         );
  dff_sg \filter_0/ow_0_reg[4]  ( .D(n43365), .CP(clk), .Q(\filter_0/n17644 )
         );
  dff_sg \filter_0/ow_0_reg[5]  ( .D(n43364), .CP(clk), .Q(\filter_0/n17643 )
         );
  dff_sg \filter_0/ow_0_reg[6]  ( .D(n43354), .CP(clk), .Q(\filter_0/n17642 )
         );
  dff_sg \filter_0/ow_0_reg[7]  ( .D(n43363), .CP(clk), .Q(\filter_0/n17641 )
         );
  dff_sg \filter_0/ow_0_reg[8]  ( .D(n43351), .CP(clk), .Q(\filter_0/n17640 )
         );
  dff_sg \filter_0/ow_0_reg[9]  ( .D(n43362), .CP(clk), .Q(\filter_0/n17639 )
         );
  dff_sg \filter_0/ow_0_reg[10]  ( .D(n43361), .CP(clk), .Q(\filter_0/n17638 )
         );
  dff_sg \filter_0/ow_0_reg[11]  ( .D(n43360), .CP(clk), .Q(\filter_0/n17637 )
         );
  dff_sg \filter_0/ow_0_reg[12]  ( .D(n43350), .CP(clk), .Q(\filter_0/n17636 )
         );
  dff_sg \filter_0/ow_0_reg[13]  ( .D(n43349), .CP(clk), .Q(\filter_0/n17635 )
         );
  dff_sg \filter_0/ow_0_reg[14]  ( .D(n43355), .CP(clk), .Q(\filter_0/n17634 )
         );
  dff_sg \filter_0/ow_0_reg[15]  ( .D(n43359), .CP(clk), .Q(\filter_0/n17633 )
         );
  dff_sg \filter_0/ow_0_reg[16]  ( .D(n43358), .CP(clk), .Q(\filter_0/n17632 )
         );
  dff_sg \filter_0/ow_0_reg[17]  ( .D(n43353), .CP(clk), .Q(\filter_0/n17631 )
         );
  dff_sg \filter_0/ow_0_reg[18]  ( .D(n43356), .CP(clk), .Q(\filter_0/n17630 )
         );
  dff_sg \filter_0/ow_0_reg[19]  ( .D(n43352), .CP(clk), .Q(\filter_0/n17629 )
         );
  dff_sg \filter_0/ow_8_reg[0]  ( .D(n43348), .CP(clk), .Q(\filter_0/n17808 )
         );
  dff_sg \filter_0/ow_8_reg[1]  ( .D(n43347), .CP(clk), .Q(\filter_0/n17807 )
         );
  dff_sg \filter_0/ow_8_reg[2]  ( .D(n43346), .CP(clk), .Q(\filter_0/n17806 )
         );
  dff_sg \filter_0/ow_8_reg[3]  ( .D(n43337), .CP(clk), .Q(\filter_0/n17805 )
         );
  dff_sg \filter_0/ow_8_reg[4]  ( .D(n43345), .CP(clk), .Q(\filter_0/n17804 )
         );
  dff_sg \filter_0/ow_8_reg[5]  ( .D(n43344), .CP(clk), .Q(\filter_0/n17803 )
         );
  dff_sg \filter_0/ow_8_reg[6]  ( .D(n43334), .CP(clk), .Q(\filter_0/n17802 )
         );
  dff_sg \filter_0/ow_8_reg[7]  ( .D(n43343), .CP(clk), .Q(\filter_0/n17801 )
         );
  dff_sg \filter_0/ow_8_reg[8]  ( .D(n43331), .CP(clk), .Q(\filter_0/n17800 )
         );
  dff_sg \filter_0/ow_8_reg[9]  ( .D(n43342), .CP(clk), .Q(\filter_0/n17799 )
         );
  dff_sg \filter_0/ow_8_reg[10]  ( .D(n43341), .CP(clk), .Q(\filter_0/n17798 )
         );
  dff_sg \filter_0/ow_8_reg[11]  ( .D(n43340), .CP(clk), .Q(\filter_0/n17797 )
         );
  dff_sg \filter_0/ow_8_reg[12]  ( .D(n43330), .CP(clk), .Q(\filter_0/n17796 )
         );
  dff_sg \filter_0/ow_8_reg[13]  ( .D(n43329), .CP(clk), .Q(\filter_0/n17795 )
         );
  dff_sg \filter_0/ow_8_reg[14]  ( .D(n43335), .CP(clk), .Q(\filter_0/n17794 )
         );
  dff_sg \filter_0/ow_8_reg[15]  ( .D(n43339), .CP(clk), .Q(\filter_0/n17793 )
         );
  dff_sg \filter_0/ow_8_reg[16]  ( .D(n43338), .CP(clk), .Q(\filter_0/n17792 )
         );
  dff_sg \filter_0/ow_8_reg[17]  ( .D(n43333), .CP(clk), .Q(\filter_0/n17791 )
         );
  dff_sg \filter_0/ow_8_reg[18]  ( .D(n43336), .CP(clk), .Q(\filter_0/n17790 )
         );
  dff_sg \filter_0/ow_8_reg[19]  ( .D(n43332), .CP(clk), .Q(\filter_0/n17789 )
         );
  dff_sg \filter_0/ow_9_reg[0]  ( .D(n43408), .CP(clk), .Q(\filter_0/n17828 )
         );
  dff_sg \filter_0/ow_9_reg[1]  ( .D(n43407), .CP(clk), .Q(\filter_0/n17827 )
         );
  dff_sg \filter_0/ow_9_reg[2]  ( .D(n43393), .CP(clk), .Q(\filter_0/n17826 )
         );
  dff_sg \filter_0/ow_9_reg[3]  ( .D(n43397), .CP(clk), .Q(\filter_0/n17825 )
         );
  dff_sg \filter_0/ow_9_reg[4]  ( .D(n43406), .CP(clk), .Q(\filter_0/n17824 )
         );
  dff_sg \filter_0/ow_9_reg[5]  ( .D(n43405), .CP(clk), .Q(\filter_0/n17823 )
         );
  dff_sg \filter_0/ow_9_reg[6]  ( .D(n43390), .CP(clk), .Q(\filter_0/n17822 )
         );
  dff_sg \filter_0/ow_9_reg[7]  ( .D(n43404), .CP(clk), .Q(\filter_0/n17821 )
         );
  dff_sg \filter_0/ow_9_reg[8]  ( .D(n43403), .CP(clk), .Q(\filter_0/n17820 )
         );
  dff_sg \filter_0/ow_9_reg[9]  ( .D(n43402), .CP(clk), .Q(\filter_0/n17819 )
         );
  dff_sg \filter_0/ow_9_reg[10]  ( .D(n43401), .CP(clk), .Q(\filter_0/n17818 )
         );
  dff_sg \filter_0/ow_9_reg[11]  ( .D(n43400), .CP(clk), .Q(\filter_0/n17817 )
         );
  dff_sg \filter_0/ow_9_reg[12]  ( .D(n43391), .CP(clk), .Q(\filter_0/n17816 )
         );
  dff_sg \filter_0/ow_9_reg[13]  ( .D(n43394), .CP(clk), .Q(\filter_0/n17815 )
         );
  dff_sg \filter_0/ow_9_reg[14]  ( .D(n43395), .CP(clk), .Q(\filter_0/n17814 )
         );
  dff_sg \filter_0/ow_9_reg[15]  ( .D(n43399), .CP(clk), .Q(\filter_0/n17813 )
         );
  dff_sg \filter_0/ow_9_reg[16]  ( .D(n43398), .CP(clk), .Q(\filter_0/n17812 )
         );
  dff_sg \filter_0/ow_9_reg[17]  ( .D(n43389), .CP(clk), .Q(\filter_0/n17811 )
         );
  dff_sg \filter_0/ow_9_reg[18]  ( .D(n43396), .CP(clk), .Q(\filter_0/n17810 )
         );
  dff_sg \filter_0/ow_9_reg[19]  ( .D(n43392), .CP(clk), .Q(\filter_0/n17809 )
         );
  dff_sg \filter_0/ow_10_reg[0]  ( .D(n43388), .CP(clk), .Q(\filter_0/n17848 )
         );
  dff_sg \filter_0/ow_10_reg[1]  ( .D(n43387), .CP(clk), .Q(\filter_0/n17847 )
         );
  dff_sg \filter_0/ow_10_reg[2]  ( .D(n43373), .CP(clk), .Q(\filter_0/n17846 )
         );
  dff_sg \filter_0/ow_10_reg[3]  ( .D(n43377), .CP(clk), .Q(\filter_0/n17845 )
         );
  dff_sg \filter_0/ow_10_reg[4]  ( .D(n43386), .CP(clk), .Q(\filter_0/n17844 )
         );
  dff_sg \filter_0/ow_10_reg[5]  ( .D(n43385), .CP(clk), .Q(\filter_0/n17843 )
         );
  dff_sg \filter_0/ow_10_reg[6]  ( .D(n43370), .CP(clk), .Q(\filter_0/n17842 )
         );
  dff_sg \filter_0/ow_10_reg[7]  ( .D(n43384), .CP(clk), .Q(\filter_0/n17841 )
         );
  dff_sg \filter_0/ow_10_reg[8]  ( .D(n43383), .CP(clk), .Q(\filter_0/n17840 )
         );
  dff_sg \filter_0/ow_10_reg[9]  ( .D(n43382), .CP(clk), .Q(\filter_0/n17839 )
         );
  dff_sg \filter_0/ow_10_reg[10]  ( .D(n43381), .CP(clk), .Q(\filter_0/n17838 ) );
  dff_sg \filter_0/ow_10_reg[11]  ( .D(n43380), .CP(clk), .Q(\filter_0/n17837 ) );
  dff_sg \filter_0/ow_10_reg[12]  ( .D(n43371), .CP(clk), .Q(\filter_0/n17836 ) );
  dff_sg \filter_0/ow_10_reg[13]  ( .D(n43374), .CP(clk), .Q(\filter_0/n17835 ) );
  dff_sg \filter_0/ow_10_reg[14]  ( .D(n43375), .CP(clk), .Q(\filter_0/n17834 ) );
  dff_sg \filter_0/ow_10_reg[15]  ( .D(n43379), .CP(clk), .Q(\filter_0/n17833 ) );
  dff_sg \filter_0/ow_10_reg[16]  ( .D(n43378), .CP(clk), .Q(\filter_0/n17832 ) );
  dff_sg \filter_0/ow_10_reg[17]  ( .D(n43369), .CP(clk), .Q(\filter_0/n17831 ) );
  dff_sg \filter_0/ow_10_reg[18]  ( .D(n43376), .CP(clk), .Q(\filter_0/n17830 ) );
  dff_sg \filter_0/ow_10_reg[19]  ( .D(n43372), .CP(clk), .Q(\filter_0/n17829 ) );
  dff_sg \filter_0/ow_11_reg[0]  ( .D(n42938), .CP(clk), .Q(\filter_0/n17868 )
         );
  dff_sg \filter_0/ow_11_reg[1]  ( .D(n42940), .CP(clk), .Q(\filter_0/n17867 )
         );
  dff_sg \filter_0/ow_11_reg[2]  ( .D(n42931), .CP(clk), .Q(\filter_0/n17866 )
         );
  dff_sg \filter_0/ow_11_reg[3]  ( .D(n42935), .CP(clk), .Q(\filter_0/n17865 )
         );
  dff_sg \filter_0/ow_11_reg[4]  ( .D(n42943), .CP(clk), .Q(\filter_0/n17864 )
         );
  dff_sg \filter_0/ow_11_reg[5]  ( .D(n42939), .CP(clk), .Q(\filter_0/n17863 )
         );
  dff_sg \filter_0/ow_11_reg[6]  ( .D(n42948), .CP(clk), .Q(\filter_0/n17862 )
         );
  dff_sg \filter_0/ow_11_reg[7]  ( .D(n42933), .CP(clk), .Q(\filter_0/n17861 )
         );
  dff_sg \filter_0/ow_11_reg[8]  ( .D(n42936), .CP(clk), .Q(\filter_0/n17860 )
         );
  dff_sg \filter_0/ow_11_reg[9]  ( .D(n42929), .CP(clk), .Q(\filter_0/n17859 )
         );
  dff_sg \filter_0/ow_11_reg[10]  ( .D(n42945), .CP(clk), .Q(\filter_0/n17858 ) );
  dff_sg \filter_0/ow_11_reg[11]  ( .D(n42934), .CP(clk), .Q(\filter_0/n17857 ) );
  dff_sg \filter_0/ow_11_reg[12]  ( .D(n42944), .CP(clk), .Q(\filter_0/n17856 ) );
  dff_sg \filter_0/ow_11_reg[13]  ( .D(n42930), .CP(clk), .Q(\filter_0/n17855 ) );
  dff_sg \filter_0/ow_11_reg[14]  ( .D(n42946), .CP(clk), .Q(\filter_0/n17854 ) );
  dff_sg \filter_0/ow_11_reg[15]  ( .D(n42947), .CP(clk), .Q(\filter_0/n17853 ) );
  dff_sg \filter_0/ow_11_reg[16]  ( .D(n42941), .CP(clk), .Q(\filter_0/n17852 ) );
  dff_sg \filter_0/ow_11_reg[17]  ( .D(n42932), .CP(clk), .Q(\filter_0/n17851 ) );
  dff_sg \filter_0/ow_11_reg[18]  ( .D(n42937), .CP(clk), .Q(\filter_0/n17850 ) );
  dff_sg \filter_0/ow_11_reg[19]  ( .D(n42942), .CP(clk), .Q(\filter_0/n17849 ) );
  dff_sg \filter_0/ow_12_reg[0]  ( .D(n43428), .CP(clk), .Q(\filter_0/n17888 )
         );
  dff_sg \filter_0/ow_12_reg[1]  ( .D(n43427), .CP(clk), .Q(\filter_0/n17887 )
         );
  dff_sg \filter_0/ow_12_reg[2]  ( .D(n43413), .CP(clk), .Q(\filter_0/n17886 )
         );
  dff_sg \filter_0/ow_12_reg[3]  ( .D(n43417), .CP(clk), .Q(\filter_0/n17885 )
         );
  dff_sg \filter_0/ow_12_reg[4]  ( .D(n43426), .CP(clk), .Q(\filter_0/n17884 )
         );
  dff_sg \filter_0/ow_12_reg[5]  ( .D(n43425), .CP(clk), .Q(\filter_0/n17883 )
         );
  dff_sg \filter_0/ow_12_reg[6]  ( .D(n43410), .CP(clk), .Q(\filter_0/n17882 )
         );
  dff_sg \filter_0/ow_12_reg[7]  ( .D(n43424), .CP(clk), .Q(\filter_0/n17881 )
         );
  dff_sg \filter_0/ow_12_reg[8]  ( .D(n43423), .CP(clk), .Q(\filter_0/n17880 )
         );
  dff_sg \filter_0/ow_12_reg[9]  ( .D(n43422), .CP(clk), .Q(\filter_0/n17879 )
         );
  dff_sg \filter_0/ow_12_reg[10]  ( .D(n43421), .CP(clk), .Q(\filter_0/n17878 ) );
  dff_sg \filter_0/ow_12_reg[11]  ( .D(n43420), .CP(clk), .Q(\filter_0/n17877 ) );
  dff_sg \filter_0/ow_12_reg[12]  ( .D(n43411), .CP(clk), .Q(\filter_0/n17876 ) );
  dff_sg \filter_0/ow_12_reg[13]  ( .D(n43414), .CP(clk), .Q(\filter_0/n17875 ) );
  dff_sg \filter_0/ow_12_reg[14]  ( .D(n43415), .CP(clk), .Q(\filter_0/n17874 ) );
  dff_sg \filter_0/ow_12_reg[15]  ( .D(n43419), .CP(clk), .Q(\filter_0/n17873 ) );
  dff_sg \filter_0/ow_12_reg[16]  ( .D(n43418), .CP(clk), .Q(\filter_0/n17872 ) );
  dff_sg \filter_0/ow_12_reg[17]  ( .D(n43409), .CP(clk), .Q(\filter_0/n17871 ) );
  dff_sg \filter_0/ow_12_reg[18]  ( .D(n43416), .CP(clk), .Q(\filter_0/n17870 ) );
  dff_sg \filter_0/ow_12_reg[19]  ( .D(n43412), .CP(clk), .Q(\filter_0/n17869 ) );
  dff_sg \filter_0/ow_13_reg[0]  ( .D(n43168), .CP(clk), .Q(\filter_0/n17908 )
         );
  dff_sg \filter_0/ow_13_reg[1]  ( .D(n43167), .CP(clk), .Q(\filter_0/n17907 )
         );
  dff_sg \filter_0/ow_13_reg[2]  ( .D(n43166), .CP(clk), .Q(\filter_0/n17906 )
         );
  dff_sg \filter_0/ow_13_reg[3]  ( .D(n43157), .CP(clk), .Q(\filter_0/n17905 )
         );
  dff_sg \filter_0/ow_13_reg[4]  ( .D(n43165), .CP(clk), .Q(\filter_0/n17904 )
         );
  dff_sg \filter_0/ow_13_reg[5]  ( .D(n43164), .CP(clk), .Q(\filter_0/n17903 )
         );
  dff_sg \filter_0/ow_13_reg[6]  ( .D(n43154), .CP(clk), .Q(\filter_0/n17902 )
         );
  dff_sg \filter_0/ow_13_reg[7]  ( .D(n43163), .CP(clk), .Q(\filter_0/n17901 )
         );
  dff_sg \filter_0/ow_13_reg[8]  ( .D(n43151), .CP(clk), .Q(\filter_0/n17900 )
         );
  dff_sg \filter_0/ow_13_reg[9]  ( .D(n43162), .CP(clk), .Q(\filter_0/n17899 )
         );
  dff_sg \filter_0/ow_13_reg[10]  ( .D(n43161), .CP(clk), .Q(\filter_0/n17898 ) );
  dff_sg \filter_0/ow_13_reg[11]  ( .D(n43160), .CP(clk), .Q(\filter_0/n17897 ) );
  dff_sg \filter_0/ow_13_reg[12]  ( .D(n43150), .CP(clk), .Q(\filter_0/n17896 ) );
  dff_sg \filter_0/ow_13_reg[13]  ( .D(n43149), .CP(clk), .Q(\filter_0/n17895 ) );
  dff_sg \filter_0/ow_13_reg[14]  ( .D(n43155), .CP(clk), .Q(\filter_0/n17894 ) );
  dff_sg \filter_0/ow_13_reg[15]  ( .D(n43159), .CP(clk), .Q(\filter_0/n17893 ) );
  dff_sg \filter_0/ow_13_reg[16]  ( .D(n43158), .CP(clk), .Q(\filter_0/n17892 ) );
  dff_sg \filter_0/ow_13_reg[17]  ( .D(n43153), .CP(clk), .Q(\filter_0/n17891 ) );
  dff_sg \filter_0/ow_13_reg[18]  ( .D(n43156), .CP(clk), .Q(\filter_0/n17890 ) );
  dff_sg \filter_0/ow_13_reg[19]  ( .D(n43152), .CP(clk), .Q(\filter_0/n17889 ) );
  dff_sg \filter_0/ow_14_reg[0]  ( .D(n43148), .CP(clk), .Q(\filter_0/n17928 )
         );
  dff_sg \filter_0/ow_14_reg[1]  ( .D(n43147), .CP(clk), .Q(\filter_0/n17927 )
         );
  dff_sg \filter_0/ow_14_reg[2]  ( .D(n43133), .CP(clk), .Q(\filter_0/n17926 )
         );
  dff_sg \filter_0/ow_14_reg[3]  ( .D(n43137), .CP(clk), .Q(\filter_0/n17925 )
         );
  dff_sg \filter_0/ow_14_reg[4]  ( .D(n43146), .CP(clk), .Q(\filter_0/n17924 )
         );
  dff_sg \filter_0/ow_14_reg[5]  ( .D(n43145), .CP(clk), .Q(\filter_0/n17923 )
         );
  dff_sg \filter_0/ow_14_reg[6]  ( .D(n43130), .CP(clk), .Q(\filter_0/n17922 )
         );
  dff_sg \filter_0/ow_14_reg[7]  ( .D(n43144), .CP(clk), .Q(\filter_0/n17921 )
         );
  dff_sg \filter_0/ow_14_reg[8]  ( .D(n43143), .CP(clk), .Q(\filter_0/n17920 )
         );
  dff_sg \filter_0/ow_14_reg[9]  ( .D(n43142), .CP(clk), .Q(\filter_0/n17919 )
         );
  dff_sg \filter_0/ow_14_reg[10]  ( .D(n43141), .CP(clk), .Q(\filter_0/n17918 ) );
  dff_sg \filter_0/ow_14_reg[11]  ( .D(n43140), .CP(clk), .Q(\filter_0/n17917 ) );
  dff_sg \filter_0/ow_14_reg[12]  ( .D(n43131), .CP(clk), .Q(\filter_0/n17916 ) );
  dff_sg \filter_0/ow_14_reg[13]  ( .D(n43134), .CP(clk), .Q(\filter_0/n17915 ) );
  dff_sg \filter_0/ow_14_reg[14]  ( .D(n43135), .CP(clk), .Q(\filter_0/n17914 ) );
  dff_sg \filter_0/ow_14_reg[15]  ( .D(n43139), .CP(clk), .Q(\filter_0/n17913 ) );
  dff_sg \filter_0/ow_14_reg[16]  ( .D(n43138), .CP(clk), .Q(\filter_0/n17912 ) );
  dff_sg \filter_0/ow_14_reg[17]  ( .D(n43129), .CP(clk), .Q(\filter_0/n17911 ) );
  dff_sg \filter_0/ow_14_reg[18]  ( .D(n43136), .CP(clk), .Q(\filter_0/n17910 ) );
  dff_sg \filter_0/ow_14_reg[19]  ( .D(n43132), .CP(clk), .Q(\filter_0/n17909 ) );
  dff_sg \filter_0/ow_15_reg[0]  ( .D(n42848), .CP(clk), .Q(\filter_0/n17948 )
         );
  dff_sg \filter_0/ow_15_reg[1]  ( .D(n42842), .CP(clk), .Q(\filter_0/n17947 )
         );
  dff_sg \filter_0/ow_15_reg[2]  ( .D(n42847), .CP(clk), .Q(\filter_0/n17946 )
         );
  dff_sg \filter_0/ow_15_reg[3]  ( .D(n42829), .CP(clk), .Q(\filter_0/n17945 )
         );
  dff_sg \filter_0/ow_15_reg[4]  ( .D(n42846), .CP(clk), .Q(\filter_0/n17944 )
         );
  dff_sg \filter_0/ow_15_reg[5]  ( .D(n42841), .CP(clk), .Q(\filter_0/n17943 )
         );
  dff_sg \filter_0/ow_15_reg[6]  ( .D(n42845), .CP(clk), .Q(\filter_0/n17942 )
         );
  dff_sg \filter_0/ow_15_reg[7]  ( .D(n42840), .CP(clk), .Q(\filter_0/n17941 )
         );
  dff_sg \filter_0/ow_15_reg[8]  ( .D(n42844), .CP(clk), .Q(\filter_0/n17940 )
         );
  dff_sg \filter_0/ow_15_reg[9]  ( .D(n42839), .CP(clk), .Q(\filter_0/n17939 )
         );
  dff_sg \filter_0/ow_15_reg[10]  ( .D(n42843), .CP(clk), .Q(\filter_0/n17938 ) );
  dff_sg \filter_0/ow_15_reg[11]  ( .D(n42838), .CP(clk), .Q(\filter_0/n17937 ) );
  dff_sg \filter_0/ow_15_reg[12]  ( .D(n42836), .CP(clk), .Q(\filter_0/n17936 ) );
  dff_sg \filter_0/ow_15_reg[13]  ( .D(n42837), .CP(clk), .Q(\filter_0/n17935 ) );
  dff_sg \filter_0/ow_15_reg[14]  ( .D(n42835), .CP(clk), .Q(\filter_0/n17934 ) );
  dff_sg \filter_0/ow_15_reg[15]  ( .D(n42834), .CP(clk), .Q(\filter_0/n17933 ) );
  dff_sg \filter_0/ow_15_reg[16]  ( .D(n42833), .CP(clk), .Q(\filter_0/n17932 ) );
  dff_sg \filter_0/ow_15_reg[17]  ( .D(n42832), .CP(clk), .Q(\filter_0/n17931 ) );
  dff_sg \filter_0/ow_15_reg[18]  ( .D(n42831), .CP(clk), .Q(\filter_0/n17930 ) );
  dff_sg \filter_0/ow_15_reg[19]  ( .D(n42830), .CP(clk), .Q(\filter_0/n17929 ) );
  dff_sg \filter_0/ow_7_reg[0]  ( .D(n43088), .CP(clk), .Q(\filter_0/n17788 )
         );
  dff_sg \filter_0/ow_7_reg[1]  ( .D(n43069), .CP(clk), .Q(\filter_0/n17787 )
         );
  dff_sg \filter_0/ow_7_reg[2]  ( .D(n43087), .CP(clk), .Q(\filter_0/n17786 )
         );
  dff_sg \filter_0/ow_7_reg[3]  ( .D(n43077), .CP(clk), .Q(\filter_0/n17785 )
         );
  dff_sg \filter_0/ow_7_reg[4]  ( .D(n43086), .CP(clk), .Q(\filter_0/n17784 )
         );
  dff_sg \filter_0/ow_7_reg[5]  ( .D(n43073), .CP(clk), .Q(\filter_0/n17783 )
         );
  dff_sg \filter_0/ow_7_reg[6]  ( .D(n43085), .CP(clk), .Q(\filter_0/n17782 )
         );
  dff_sg \filter_0/ow_7_reg[7]  ( .D(n43071), .CP(clk), .Q(\filter_0/n17781 )
         );
  dff_sg \filter_0/ow_7_reg[8]  ( .D(n43084), .CP(clk), .Q(\filter_0/n17780 )
         );
  dff_sg \filter_0/ow_7_reg[9]  ( .D(n43074), .CP(clk), .Q(\filter_0/n17779 )
         );
  dff_sg \filter_0/ow_7_reg[10]  ( .D(n43083), .CP(clk), .Q(\filter_0/n17778 )
         );
  dff_sg \filter_0/ow_7_reg[11]  ( .D(n43070), .CP(clk), .Q(\filter_0/n17777 )
         );
  dff_sg \filter_0/ow_7_reg[12]  ( .D(n43082), .CP(clk), .Q(\filter_0/n17776 )
         );
  dff_sg \filter_0/ow_7_reg[13]  ( .D(n43081), .CP(clk), .Q(\filter_0/n17775 )
         );
  dff_sg \filter_0/ow_7_reg[14]  ( .D(n43075), .CP(clk), .Q(\filter_0/n17774 )
         );
  dff_sg \filter_0/ow_7_reg[15]  ( .D(n43072), .CP(clk), .Q(\filter_0/n17773 )
         );
  dff_sg \filter_0/ow_7_reg[16]  ( .D(n43080), .CP(clk), .Q(\filter_0/n17772 )
         );
  dff_sg \filter_0/ow_7_reg[17]  ( .D(n43079), .CP(clk), .Q(\filter_0/n17771 )
         );
  dff_sg \filter_0/ow_7_reg[18]  ( .D(n43076), .CP(clk), .Q(\filter_0/n17770 )
         );
  dff_sg \filter_0/ow_7_reg[19]  ( .D(n43078), .CP(clk), .Q(\filter_0/n17769 )
         );
  dff_sg \filter_0/ow_6_reg[0]  ( .D(n43068), .CP(clk), .Q(\filter_0/n17768 )
         );
  dff_sg \filter_0/ow_6_reg[1]  ( .D(n43067), .CP(clk), .Q(\filter_0/n17767 )
         );
  dff_sg \filter_0/ow_6_reg[2]  ( .D(n43066), .CP(clk), .Q(\filter_0/n17766 )
         );
  dff_sg \filter_0/ow_6_reg[3]  ( .D(n43057), .CP(clk), .Q(\filter_0/n17765 )
         );
  dff_sg \filter_0/ow_6_reg[4]  ( .D(n43065), .CP(clk), .Q(\filter_0/n17764 )
         );
  dff_sg \filter_0/ow_6_reg[5]  ( .D(n43064), .CP(clk), .Q(\filter_0/n17763 )
         );
  dff_sg \filter_0/ow_6_reg[6]  ( .D(n43054), .CP(clk), .Q(\filter_0/n17762 )
         );
  dff_sg \filter_0/ow_6_reg[7]  ( .D(n43063), .CP(clk), .Q(\filter_0/n17761 )
         );
  dff_sg \filter_0/ow_6_reg[8]  ( .D(n43051), .CP(clk), .Q(\filter_0/n17760 )
         );
  dff_sg \filter_0/ow_6_reg[9]  ( .D(n43062), .CP(clk), .Q(\filter_0/n17759 )
         );
  dff_sg \filter_0/ow_6_reg[10]  ( .D(n43061), .CP(clk), .Q(\filter_0/n17758 )
         );
  dff_sg \filter_0/ow_6_reg[11]  ( .D(n43060), .CP(clk), .Q(\filter_0/n17757 )
         );
  dff_sg \filter_0/ow_6_reg[12]  ( .D(n43050), .CP(clk), .Q(\filter_0/n17756 )
         );
  dff_sg \filter_0/ow_6_reg[13]  ( .D(n43049), .CP(clk), .Q(\filter_0/n17755 )
         );
  dff_sg \filter_0/ow_6_reg[14]  ( .D(n43055), .CP(clk), .Q(\filter_0/n17754 )
         );
  dff_sg \filter_0/ow_6_reg[15]  ( .D(n43059), .CP(clk), .Q(\filter_0/n17753 )
         );
  dff_sg \filter_0/ow_6_reg[16]  ( .D(n43058), .CP(clk), .Q(\filter_0/n17752 )
         );
  dff_sg \filter_0/ow_6_reg[17]  ( .D(n43053), .CP(clk), .Q(\filter_0/n17751 )
         );
  dff_sg \filter_0/ow_6_reg[18]  ( .D(n43056), .CP(clk), .Q(\filter_0/n17750 )
         );
  dff_sg \filter_0/ow_6_reg[19]  ( .D(n43052), .CP(clk), .Q(\filter_0/n17749 )
         );
  dff_sg \filter_0/ow_5_reg[0]  ( .D(n43048), .CP(clk), .Q(\filter_0/n17748 )
         );
  dff_sg \filter_0/ow_5_reg[1]  ( .D(n43047), .CP(clk), .Q(\filter_0/n17747 )
         );
  dff_sg \filter_0/ow_5_reg[2]  ( .D(n43033), .CP(clk), .Q(\filter_0/n17746 )
         );
  dff_sg \filter_0/ow_5_reg[3]  ( .D(n43037), .CP(clk), .Q(\filter_0/n17745 )
         );
  dff_sg \filter_0/ow_5_reg[4]  ( .D(n43046), .CP(clk), .Q(\filter_0/n17744 )
         );
  dff_sg \filter_0/ow_5_reg[5]  ( .D(n43045), .CP(clk), .Q(\filter_0/n17743 )
         );
  dff_sg \filter_0/ow_5_reg[6]  ( .D(n43030), .CP(clk), .Q(\filter_0/n17742 )
         );
  dff_sg \filter_0/ow_5_reg[7]  ( .D(n43044), .CP(clk), .Q(\filter_0/n17741 )
         );
  dff_sg \filter_0/ow_5_reg[8]  ( .D(n43043), .CP(clk), .Q(\filter_0/n17740 )
         );
  dff_sg \filter_0/ow_5_reg[9]  ( .D(n43042), .CP(clk), .Q(\filter_0/n17739 )
         );
  dff_sg \filter_0/ow_5_reg[10]  ( .D(n43041), .CP(clk), .Q(\filter_0/n17738 )
         );
  dff_sg \filter_0/ow_5_reg[11]  ( .D(n43040), .CP(clk), .Q(\filter_0/n17737 )
         );
  dff_sg \filter_0/ow_5_reg[12]  ( .D(n43031), .CP(clk), .Q(\filter_0/n17736 )
         );
  dff_sg \filter_0/ow_5_reg[13]  ( .D(n43034), .CP(clk), .Q(\filter_0/n17735 )
         );
  dff_sg \filter_0/ow_5_reg[14]  ( .D(n43035), .CP(clk), .Q(\filter_0/n17734 )
         );
  dff_sg \filter_0/ow_5_reg[15]  ( .D(n43039), .CP(clk), .Q(\filter_0/n17733 )
         );
  dff_sg \filter_0/ow_5_reg[16]  ( .D(n43038), .CP(clk), .Q(\filter_0/n17732 )
         );
  dff_sg \filter_0/ow_5_reg[17]  ( .D(n43029), .CP(clk), .Q(\filter_0/n17731 )
         );
  dff_sg \filter_0/ow_5_reg[18]  ( .D(n43036), .CP(clk), .Q(\filter_0/n17730 )
         );
  dff_sg \filter_0/ow_5_reg[19]  ( .D(n43032), .CP(clk), .Q(\filter_0/n17729 )
         );
  dff_sg \filter_0/ow_4_reg[0]  ( .D(n43468), .CP(clk), .Q(\filter_0/n17728 )
         );
  dff_sg \filter_0/ow_4_reg[1]  ( .D(n43467), .CP(clk), .Q(\filter_0/n17727 )
         );
  dff_sg \filter_0/ow_4_reg[2]  ( .D(n43451), .CP(clk), .Q(\filter_0/n17726 )
         );
  dff_sg \filter_0/ow_4_reg[3]  ( .D(n43461), .CP(clk), .Q(\filter_0/n17725 )
         );
  dff_sg \filter_0/ow_4_reg[4]  ( .D(n43453), .CP(clk), .Q(\filter_0/n17724 )
         );
  dff_sg \filter_0/ow_4_reg[5]  ( .D(n43466), .CP(clk), .Q(\filter_0/n17723 )
         );
  dff_sg \filter_0/ow_4_reg[6]  ( .D(n43458), .CP(clk), .Q(\filter_0/n17722 )
         );
  dff_sg \filter_0/ow_4_reg[7]  ( .D(n43449), .CP(clk), .Q(\filter_0/n17721 )
         );
  dff_sg \filter_0/ow_4_reg[8]  ( .D(n43456), .CP(clk), .Q(\filter_0/n17720 )
         );
  dff_sg \filter_0/ow_4_reg[9]  ( .D(n43465), .CP(clk), .Q(\filter_0/n17719 )
         );
  dff_sg \filter_0/ow_4_reg[10]  ( .D(n43457), .CP(clk), .Q(\filter_0/n17718 )
         );
  dff_sg \filter_0/ow_4_reg[11]  ( .D(n43464), .CP(clk), .Q(\filter_0/n17717 )
         );
  dff_sg \filter_0/ow_4_reg[12]  ( .D(n43455), .CP(clk), .Q(\filter_0/n17716 )
         );
  dff_sg \filter_0/ow_4_reg[13]  ( .D(n43459), .CP(clk), .Q(\filter_0/n17715 )
         );
  dff_sg \filter_0/ow_4_reg[14]  ( .D(n43454), .CP(clk), .Q(\filter_0/n17714 )
         );
  dff_sg \filter_0/ow_4_reg[15]  ( .D(n43463), .CP(clk), .Q(\filter_0/n17713 )
         );
  dff_sg \filter_0/ow_4_reg[16]  ( .D(n43462), .CP(clk), .Q(\filter_0/n17712 )
         );
  dff_sg \filter_0/ow_4_reg[17]  ( .D(n43450), .CP(clk), .Q(\filter_0/n17711 )
         );
  dff_sg \filter_0/ow_4_reg[18]  ( .D(n43460), .CP(clk), .Q(\filter_0/n17710 )
         );
  dff_sg \filter_0/ow_4_reg[19]  ( .D(n43452), .CP(clk), .Q(\filter_0/n17709 )
         );
  dff_sg \filter_0/ow_3_reg[0]  ( .D(n42920), .CP(clk), .Q(\filter_0/n17708 )
         );
  dff_sg \filter_0/ow_3_reg[1]  ( .D(n42914), .CP(clk), .Q(\filter_0/n17707 )
         );
  dff_sg \filter_0/ow_3_reg[2]  ( .D(n42911), .CP(clk), .Q(\filter_0/n17706 )
         );
  dff_sg \filter_0/ow_3_reg[3]  ( .D(n42925), .CP(clk), .Q(\filter_0/n17705 )
         );
  dff_sg \filter_0/ow_3_reg[4]  ( .D(n42923), .CP(clk), .Q(\filter_0/n17704 )
         );
  dff_sg \filter_0/ow_3_reg[5]  ( .D(n42919), .CP(clk), .Q(\filter_0/n17703 )
         );
  dff_sg \filter_0/ow_3_reg[6]  ( .D(n42915), .CP(clk), .Q(\filter_0/n17702 )
         );
  dff_sg \filter_0/ow_3_reg[7]  ( .D(n42928), .CP(clk), .Q(\filter_0/n17701 )
         );
  dff_sg \filter_0/ow_3_reg[8]  ( .D(n42918), .CP(clk), .Q(\filter_0/n17700 )
         );
  dff_sg \filter_0/ow_3_reg[9]  ( .D(n42922), .CP(clk), .Q(\filter_0/n17699 )
         );
  dff_sg \filter_0/ow_3_reg[10]  ( .D(n42909), .CP(clk), .Q(\filter_0/n17698 )
         );
  dff_sg \filter_0/ow_3_reg[11]  ( .D(n42916), .CP(clk), .Q(\filter_0/n17697 )
         );
  dff_sg \filter_0/ow_3_reg[12]  ( .D(n42910), .CP(clk), .Q(\filter_0/n17696 )
         );
  dff_sg \filter_0/ow_3_reg[13]  ( .D(n42924), .CP(clk), .Q(\filter_0/n17695 )
         );
  dff_sg \filter_0/ow_3_reg[14]  ( .D(n42926), .CP(clk), .Q(\filter_0/n17694 )
         );
  dff_sg \filter_0/ow_3_reg[15]  ( .D(n42921), .CP(clk), .Q(\filter_0/n17693 )
         );
  dff_sg \filter_0/ow_3_reg[16]  ( .D(n42913), .CP(clk), .Q(\filter_0/n17692 )
         );
  dff_sg \filter_0/ow_3_reg[17]  ( .D(n42912), .CP(clk), .Q(\filter_0/n17691 )
         );
  dff_sg \filter_0/ow_3_reg[18]  ( .D(n42917), .CP(clk), .Q(\filter_0/n17690 )
         );
  dff_sg \filter_0/ow_3_reg[19]  ( .D(n42927), .CP(clk), .Q(\filter_0/n17689 )
         );
  dff_sg \filter_0/ow_2_reg[0]  ( .D(n43128), .CP(clk), .Q(\filter_0/n17688 )
         );
  dff_sg \filter_0/ow_2_reg[1]  ( .D(n43127), .CP(clk), .Q(\filter_0/n17687 )
         );
  dff_sg \filter_0/ow_2_reg[2]  ( .D(n43113), .CP(clk), .Q(\filter_0/n17686 )
         );
  dff_sg \filter_0/ow_2_reg[3]  ( .D(n43117), .CP(clk), .Q(\filter_0/n17685 )
         );
  dff_sg \filter_0/ow_2_reg[4]  ( .D(n43126), .CP(clk), .Q(\filter_0/n17684 )
         );
  dff_sg \filter_0/ow_2_reg[5]  ( .D(n43125), .CP(clk), .Q(\filter_0/n17683 )
         );
  dff_sg \filter_0/ow_2_reg[6]  ( .D(n43110), .CP(clk), .Q(\filter_0/n17682 )
         );
  dff_sg \filter_0/ow_2_reg[7]  ( .D(n43124), .CP(clk), .Q(\filter_0/n17681 )
         );
  dff_sg \filter_0/ow_2_reg[8]  ( .D(n43123), .CP(clk), .Q(\filter_0/n17680 )
         );
  dff_sg \filter_0/ow_2_reg[9]  ( .D(n43122), .CP(clk), .Q(\filter_0/n17679 )
         );
  dff_sg \filter_0/ow_2_reg[10]  ( .D(n43121), .CP(clk), .Q(\filter_0/n17678 )
         );
  dff_sg \filter_0/ow_2_reg[11]  ( .D(n43120), .CP(clk), .Q(\filter_0/n17677 )
         );
  dff_sg \filter_0/ow_2_reg[12]  ( .D(n43111), .CP(clk), .Q(\filter_0/n17676 )
         );
  dff_sg \filter_0/ow_2_reg[13]  ( .D(n43114), .CP(clk), .Q(\filter_0/n17675 )
         );
  dff_sg \filter_0/ow_2_reg[14]  ( .D(n43115), .CP(clk), .Q(\filter_0/n17674 )
         );
  dff_sg \filter_0/ow_2_reg[15]  ( .D(n43119), .CP(clk), .Q(\filter_0/n17673 )
         );
  dff_sg \filter_0/ow_2_reg[16]  ( .D(n43118), .CP(clk), .Q(\filter_0/n17672 )
         );
  dff_sg \filter_0/ow_2_reg[17]  ( .D(n43109), .CP(clk), .Q(\filter_0/n17671 )
         );
  dff_sg \filter_0/ow_2_reg[18]  ( .D(n43116), .CP(clk), .Q(\filter_0/n17670 )
         );
  dff_sg \filter_0/ow_2_reg[19]  ( .D(n43112), .CP(clk), .Q(\filter_0/n17669 )
         );
  dff_sg \filter_0/ow_1_reg[0]  ( .D(n43108), .CP(clk), .Q(\filter_0/n17668 )
         );
  dff_sg \filter_0/ow_1_reg[1]  ( .D(n43107), .CP(clk), .Q(\filter_0/n17667 )
         );
  dff_sg \filter_0/ow_1_reg[2]  ( .D(n43093), .CP(clk), .Q(\filter_0/n17666 )
         );
  dff_sg \filter_0/ow_1_reg[3]  ( .D(n43097), .CP(clk), .Q(\filter_0/n17665 )
         );
  dff_sg \filter_0/ow_1_reg[4]  ( .D(n43106), .CP(clk), .Q(\filter_0/n17664 )
         );
  dff_sg \filter_0/ow_1_reg[5]  ( .D(n43105), .CP(clk), .Q(\filter_0/n17663 )
         );
  dff_sg \filter_0/ow_1_reg[6]  ( .D(n43090), .CP(clk), .Q(\filter_0/n17662 )
         );
  dff_sg \filter_0/ow_1_reg[7]  ( .D(n43104), .CP(clk), .Q(\filter_0/n17661 )
         );
  dff_sg \filter_0/ow_1_reg[8]  ( .D(n43103), .CP(clk), .Q(\filter_0/n17660 )
         );
  dff_sg \filter_0/ow_1_reg[9]  ( .D(n43102), .CP(clk), .Q(\filter_0/n17659 )
         );
  dff_sg \filter_0/ow_1_reg[10]  ( .D(n43101), .CP(clk), .Q(\filter_0/n17658 )
         );
  dff_sg \filter_0/ow_1_reg[11]  ( .D(n43100), .CP(clk), .Q(\filter_0/n17657 )
         );
  dff_sg \filter_0/ow_1_reg[12]  ( .D(n43091), .CP(clk), .Q(\filter_0/n17656 )
         );
  dff_sg \filter_0/ow_1_reg[13]  ( .D(n43094), .CP(clk), .Q(\filter_0/n17655 )
         );
  dff_sg \filter_0/ow_1_reg[14]  ( .D(n43095), .CP(clk), .Q(\filter_0/n17654 )
         );
  dff_sg \filter_0/ow_1_reg[15]  ( .D(n43099), .CP(clk), .Q(\filter_0/n17653 )
         );
  dff_sg \filter_0/ow_1_reg[16]  ( .D(n43098), .CP(clk), .Q(\filter_0/n17652 )
         );
  dff_sg \filter_0/ow_1_reg[17]  ( .D(n43089), .CP(clk), .Q(\filter_0/n17651 )
         );
  dff_sg \filter_0/ow_1_reg[18]  ( .D(n43096), .CP(clk), .Q(\filter_0/n17650 )
         );
  dff_sg \filter_0/ow_1_reg[19]  ( .D(n43092), .CP(clk), .Q(\filter_0/n17649 )
         );
  dff_sg \filter_0/oi_0_reg[0]  ( .D(n43328), .CP(clk), .Q(\filter_0/n17328 )
         );
  dff_sg \filter_0/oi_0_reg[1]  ( .D(n43327), .CP(clk), .Q(\filter_0/n17327 )
         );
  dff_sg \filter_0/oi_0_reg[2]  ( .D(n43326), .CP(clk), .Q(\filter_0/n17326 )
         );
  dff_sg \filter_0/oi_0_reg[3]  ( .D(n43317), .CP(clk), .Q(\filter_0/n17325 )
         );
  dff_sg \filter_0/oi_0_reg[4]  ( .D(n43325), .CP(clk), .Q(\filter_0/n17324 )
         );
  dff_sg \filter_0/oi_0_reg[5]  ( .D(n43324), .CP(clk), .Q(\filter_0/n17323 )
         );
  dff_sg \filter_0/oi_0_reg[6]  ( .D(n43314), .CP(clk), .Q(\filter_0/n17322 )
         );
  dff_sg \filter_0/oi_0_reg[7]  ( .D(n43323), .CP(clk), .Q(\filter_0/n17321 )
         );
  dff_sg \filter_0/oi_0_reg[8]  ( .D(n43311), .CP(clk), .Q(\filter_0/n17320 )
         );
  dff_sg \filter_0/oi_0_reg[9]  ( .D(n43322), .CP(clk), .Q(\filter_0/n17319 )
         );
  dff_sg \filter_0/oi_0_reg[10]  ( .D(n43321), .CP(clk), .Q(\filter_0/n17318 )
         );
  dff_sg \filter_0/oi_0_reg[11]  ( .D(n43320), .CP(clk), .Q(\filter_0/n17317 )
         );
  dff_sg \filter_0/oi_0_reg[12]  ( .D(n43310), .CP(clk), .Q(\filter_0/n17316 )
         );
  dff_sg \filter_0/oi_0_reg[13]  ( .D(n43309), .CP(clk), .Q(\filter_0/n17315 )
         );
  dff_sg \filter_0/oi_0_reg[14]  ( .D(n43315), .CP(clk), .Q(\filter_0/n17314 )
         );
  dff_sg \filter_0/oi_0_reg[15]  ( .D(n43319), .CP(clk), .Q(\filter_0/n17313 )
         );
  dff_sg \filter_0/oi_0_reg[16]  ( .D(n43318), .CP(clk), .Q(\filter_0/n17312 )
         );
  dff_sg \filter_0/oi_0_reg[17]  ( .D(n43313), .CP(clk), .Q(\filter_0/n17311 )
         );
  dff_sg \filter_0/oi_0_reg[18]  ( .D(n43316), .CP(clk), .Q(\filter_0/n17310 )
         );
  dff_sg \filter_0/oi_0_reg[19]  ( .D(n43312), .CP(clk), .Q(\filter_0/n17309 )
         );
  dff_sg \filter_0/oi_8_reg[0]  ( .D(n43308), .CP(clk), .Q(\filter_0/n17488 )
         );
  dff_sg \filter_0/oi_8_reg[1]  ( .D(n43307), .CP(clk), .Q(\filter_0/n17487 )
         );
  dff_sg \filter_0/oi_8_reg[2]  ( .D(n43306), .CP(clk), .Q(\filter_0/n17486 )
         );
  dff_sg \filter_0/oi_8_reg[3]  ( .D(n43297), .CP(clk), .Q(\filter_0/n17485 )
         );
  dff_sg \filter_0/oi_8_reg[4]  ( .D(n43305), .CP(clk), .Q(\filter_0/n17484 )
         );
  dff_sg \filter_0/oi_8_reg[5]  ( .D(n43304), .CP(clk), .Q(\filter_0/n17483 )
         );
  dff_sg \filter_0/oi_8_reg[6]  ( .D(n43294), .CP(clk), .Q(\filter_0/n17482 )
         );
  dff_sg \filter_0/oi_8_reg[7]  ( .D(n43303), .CP(clk), .Q(\filter_0/n17481 )
         );
  dff_sg \filter_0/oi_8_reg[8]  ( .D(n43291), .CP(clk), .Q(\filter_0/n17480 )
         );
  dff_sg \filter_0/oi_8_reg[9]  ( .D(n43302), .CP(clk), .Q(\filter_0/n17479 )
         );
  dff_sg \filter_0/oi_8_reg[10]  ( .D(n43301), .CP(clk), .Q(\filter_0/n17478 )
         );
  dff_sg \filter_0/oi_8_reg[11]  ( .D(n43300), .CP(clk), .Q(\filter_0/n17477 )
         );
  dff_sg \filter_0/oi_8_reg[12]  ( .D(n43290), .CP(clk), .Q(\filter_0/n17476 )
         );
  dff_sg \filter_0/oi_8_reg[13]  ( .D(n43289), .CP(clk), .Q(\filter_0/n17475 )
         );
  dff_sg \filter_0/oi_8_reg[14]  ( .D(n43295), .CP(clk), .Q(\filter_0/n17474 )
         );
  dff_sg \filter_0/oi_8_reg[15]  ( .D(n43299), .CP(clk), .Q(\filter_0/n17473 )
         );
  dff_sg \filter_0/oi_8_reg[16]  ( .D(n43298), .CP(clk), .Q(\filter_0/n17472 )
         );
  dff_sg \filter_0/oi_8_reg[17]  ( .D(n43293), .CP(clk), .Q(\filter_0/n17471 )
         );
  dff_sg \filter_0/oi_8_reg[18]  ( .D(n43296), .CP(clk), .Q(\filter_0/n17470 )
         );
  dff_sg \filter_0/oi_8_reg[19]  ( .D(n43292), .CP(clk), .Q(\filter_0/n17469 )
         );
  dff_sg \filter_0/oi_9_reg[0]  ( .D(n43288), .CP(clk), .Q(\filter_0/n17508 )
         );
  dff_sg \filter_0/oi_9_reg[1]  ( .D(n43287), .CP(clk), .Q(\filter_0/n17507 )
         );
  dff_sg \filter_0/oi_9_reg[2]  ( .D(n43273), .CP(clk), .Q(\filter_0/n17506 )
         );
  dff_sg \filter_0/oi_9_reg[3]  ( .D(n43277), .CP(clk), .Q(\filter_0/n17505 )
         );
  dff_sg \filter_0/oi_9_reg[4]  ( .D(n43286), .CP(clk), .Q(\filter_0/n17504 )
         );
  dff_sg \filter_0/oi_9_reg[5]  ( .D(n43285), .CP(clk), .Q(\filter_0/n17503 )
         );
  dff_sg \filter_0/oi_9_reg[6]  ( .D(n43270), .CP(clk), .Q(\filter_0/n17502 )
         );
  dff_sg \filter_0/oi_9_reg[7]  ( .D(n43284), .CP(clk), .Q(\filter_0/n17501 )
         );
  dff_sg \filter_0/oi_9_reg[8]  ( .D(n43283), .CP(clk), .Q(\filter_0/n17500 )
         );
  dff_sg \filter_0/oi_9_reg[9]  ( .D(n43282), .CP(clk), .Q(\filter_0/n17499 )
         );
  dff_sg \filter_0/oi_9_reg[10]  ( .D(n43281), .CP(clk), .Q(\filter_0/n17498 )
         );
  dff_sg \filter_0/oi_9_reg[11]  ( .D(n43280), .CP(clk), .Q(\filter_0/n17497 )
         );
  dff_sg \filter_0/oi_9_reg[12]  ( .D(n43271), .CP(clk), .Q(\filter_0/n17496 )
         );
  dff_sg \filter_0/oi_9_reg[13]  ( .D(n43274), .CP(clk), .Q(\filter_0/n17495 )
         );
  dff_sg \filter_0/oi_9_reg[14]  ( .D(n43275), .CP(clk), .Q(\filter_0/n17494 )
         );
  dff_sg \filter_0/oi_9_reg[15]  ( .D(n43279), .CP(clk), .Q(\filter_0/n17493 )
         );
  dff_sg \filter_0/oi_9_reg[16]  ( .D(n43278), .CP(clk), .Q(\filter_0/n17492 )
         );
  dff_sg \filter_0/oi_9_reg[17]  ( .D(n43269), .CP(clk), .Q(\filter_0/n17491 )
         );
  dff_sg \filter_0/oi_9_reg[18]  ( .D(n43276), .CP(clk), .Q(\filter_0/n17490 )
         );
  dff_sg \filter_0/oi_9_reg[19]  ( .D(n43272), .CP(clk), .Q(\filter_0/n17489 )
         );
  dff_sg \filter_0/oi_10_reg[0]  ( .D(n43268), .CP(clk), .Q(\filter_0/n17528 )
         );
  dff_sg \filter_0/oi_10_reg[1]  ( .D(n43267), .CP(clk), .Q(\filter_0/n17527 )
         );
  dff_sg \filter_0/oi_10_reg[2]  ( .D(n43253), .CP(clk), .Q(\filter_0/n17526 )
         );
  dff_sg \filter_0/oi_10_reg[3]  ( .D(n43257), .CP(clk), .Q(\filter_0/n17525 )
         );
  dff_sg \filter_0/oi_10_reg[4]  ( .D(n43266), .CP(clk), .Q(\filter_0/n17524 )
         );
  dff_sg \filter_0/oi_10_reg[5]  ( .D(n43265), .CP(clk), .Q(\filter_0/n17523 )
         );
  dff_sg \filter_0/oi_10_reg[6]  ( .D(n43250), .CP(clk), .Q(\filter_0/n17522 )
         );
  dff_sg \filter_0/oi_10_reg[7]  ( .D(n43264), .CP(clk), .Q(\filter_0/n17521 )
         );
  dff_sg \filter_0/oi_10_reg[8]  ( .D(n43263), .CP(clk), .Q(\filter_0/n17520 )
         );
  dff_sg \filter_0/oi_10_reg[9]  ( .D(n43262), .CP(clk), .Q(\filter_0/n17519 )
         );
  dff_sg \filter_0/oi_10_reg[10]  ( .D(n43261), .CP(clk), .Q(\filter_0/n17518 ) );
  dff_sg \filter_0/oi_10_reg[11]  ( .D(n43260), .CP(clk), .Q(\filter_0/n17517 ) );
  dff_sg \filter_0/oi_10_reg[12]  ( .D(n43251), .CP(clk), .Q(\filter_0/n17516 ) );
  dff_sg \filter_0/oi_10_reg[13]  ( .D(n43254), .CP(clk), .Q(\filter_0/n17515 ) );
  dff_sg \filter_0/oi_10_reg[14]  ( .D(n43255), .CP(clk), .Q(\filter_0/n17514 ) );
  dff_sg \filter_0/oi_10_reg[15]  ( .D(n43259), .CP(clk), .Q(\filter_0/n17513 ) );
  dff_sg \filter_0/oi_10_reg[16]  ( .D(n43258), .CP(clk), .Q(\filter_0/n17512 ) );
  dff_sg \filter_0/oi_10_reg[17]  ( .D(n43249), .CP(clk), .Q(\filter_0/n17511 ) );
  dff_sg \filter_0/oi_10_reg[18]  ( .D(n43256), .CP(clk), .Q(\filter_0/n17510 ) );
  dff_sg \filter_0/oi_10_reg[19]  ( .D(n43252), .CP(clk), .Q(\filter_0/n17509 ) );
  dff_sg \filter_0/oi_11_reg[0]  ( .D(n42898), .CP(clk), .Q(\filter_0/n17548 )
         );
  dff_sg \filter_0/oi_11_reg[1]  ( .D(n42900), .CP(clk), .Q(\filter_0/n17547 )
         );
  dff_sg \filter_0/oi_11_reg[2]  ( .D(n42891), .CP(clk), .Q(\filter_0/n17546 )
         );
  dff_sg \filter_0/oi_11_reg[3]  ( .D(n42895), .CP(clk), .Q(\filter_0/n17545 )
         );
  dff_sg \filter_0/oi_11_reg[4]  ( .D(n42903), .CP(clk), .Q(\filter_0/n17544 )
         );
  dff_sg \filter_0/oi_11_reg[5]  ( .D(n42899), .CP(clk), .Q(\filter_0/n17543 )
         );
  dff_sg \filter_0/oi_11_reg[6]  ( .D(n42908), .CP(clk), .Q(\filter_0/n17542 )
         );
  dff_sg \filter_0/oi_11_reg[7]  ( .D(n42893), .CP(clk), .Q(\filter_0/n17541 )
         );
  dff_sg \filter_0/oi_11_reg[8]  ( .D(n42896), .CP(clk), .Q(\filter_0/n17540 )
         );
  dff_sg \filter_0/oi_11_reg[9]  ( .D(n42889), .CP(clk), .Q(\filter_0/n17539 )
         );
  dff_sg \filter_0/oi_11_reg[10]  ( .D(n42905), .CP(clk), .Q(\filter_0/n17538 ) );
  dff_sg \filter_0/oi_11_reg[11]  ( .D(n42894), .CP(clk), .Q(\filter_0/n17537 ) );
  dff_sg \filter_0/oi_11_reg[12]  ( .D(n42904), .CP(clk), .Q(\filter_0/n17536 ) );
  dff_sg \filter_0/oi_11_reg[13]  ( .D(n42890), .CP(clk), .Q(\filter_0/n17535 ) );
  dff_sg \filter_0/oi_11_reg[14]  ( .D(n42906), .CP(clk), .Q(\filter_0/n17534 ) );
  dff_sg \filter_0/oi_11_reg[15]  ( .D(n42907), .CP(clk), .Q(\filter_0/n17533 ) );
  dff_sg \filter_0/oi_11_reg[16]  ( .D(n42901), .CP(clk), .Q(\filter_0/n17532 ) );
  dff_sg \filter_0/oi_11_reg[17]  ( .D(n42892), .CP(clk), .Q(\filter_0/n17531 ) );
  dff_sg \filter_0/oi_11_reg[18]  ( .D(n42897), .CP(clk), .Q(\filter_0/n17530 ) );
  dff_sg \filter_0/oi_11_reg[19]  ( .D(n42902), .CP(clk), .Q(\filter_0/n17529 ) );
  dff_sg \filter_0/oi_12_reg[0]  ( .D(n43028), .CP(clk), .Q(\filter_0/n17568 )
         );
  dff_sg \filter_0/oi_12_reg[1]  ( .D(n43027), .CP(clk), .Q(\filter_0/n17567 )
         );
  dff_sg \filter_0/oi_12_reg[2]  ( .D(n43013), .CP(clk), .Q(\filter_0/n17566 )
         );
  dff_sg \filter_0/oi_12_reg[3]  ( .D(n43017), .CP(clk), .Q(\filter_0/n17565 )
         );
  dff_sg \filter_0/oi_12_reg[4]  ( .D(n43026), .CP(clk), .Q(\filter_0/n17564 )
         );
  dff_sg \filter_0/oi_12_reg[5]  ( .D(n43025), .CP(clk), .Q(\filter_0/n17563 )
         );
  dff_sg \filter_0/oi_12_reg[6]  ( .D(n43010), .CP(clk), .Q(\filter_0/n17562 )
         );
  dff_sg \filter_0/oi_12_reg[7]  ( .D(n43024), .CP(clk), .Q(\filter_0/n17561 )
         );
  dff_sg \filter_0/oi_12_reg[8]  ( .D(n43023), .CP(clk), .Q(\filter_0/n17560 )
         );
  dff_sg \filter_0/oi_12_reg[9]  ( .D(n43022), .CP(clk), .Q(\filter_0/n17559 )
         );
  dff_sg \filter_0/oi_12_reg[10]  ( .D(n43021), .CP(clk), .Q(\filter_0/n17558 ) );
  dff_sg \filter_0/oi_12_reg[11]  ( .D(n43020), .CP(clk), .Q(\filter_0/n17557 ) );
  dff_sg \filter_0/oi_12_reg[12]  ( .D(n43011), .CP(clk), .Q(\filter_0/n17556 ) );
  dff_sg \filter_0/oi_12_reg[13]  ( .D(n43014), .CP(clk), .Q(\filter_0/n17555 ) );
  dff_sg \filter_0/oi_12_reg[14]  ( .D(n43015), .CP(clk), .Q(\filter_0/n17554 ) );
  dff_sg \filter_0/oi_12_reg[15]  ( .D(n43019), .CP(clk), .Q(\filter_0/n17553 ) );
  dff_sg \filter_0/oi_12_reg[16]  ( .D(n43018), .CP(clk), .Q(\filter_0/n17552 ) );
  dff_sg \filter_0/oi_12_reg[17]  ( .D(n43009), .CP(clk), .Q(\filter_0/n17551 ) );
  dff_sg \filter_0/oi_12_reg[18]  ( .D(n43016), .CP(clk), .Q(\filter_0/n17550 ) );
  dff_sg \filter_0/oi_12_reg[19]  ( .D(n43012), .CP(clk), .Q(\filter_0/n17549 ) );
  dff_sg \filter_0/oi_13_reg[0]  ( .D(n43008), .CP(clk), .Q(\filter_0/n17588 )
         );
  dff_sg \filter_0/oi_13_reg[1]  ( .D(n43007), .CP(clk), .Q(\filter_0/n17587 )
         );
  dff_sg \filter_0/oi_13_reg[2]  ( .D(n43006), .CP(clk), .Q(\filter_0/n17586 )
         );
  dff_sg \filter_0/oi_13_reg[3]  ( .D(n42997), .CP(clk), .Q(\filter_0/n17585 )
         );
  dff_sg \filter_0/oi_13_reg[4]  ( .D(n43005), .CP(clk), .Q(\filter_0/n17584 )
         );
  dff_sg \filter_0/oi_13_reg[5]  ( .D(n43004), .CP(clk), .Q(\filter_0/n17583 )
         );
  dff_sg \filter_0/oi_13_reg[6]  ( .D(n42994), .CP(clk), .Q(\filter_0/n17582 )
         );
  dff_sg \filter_0/oi_13_reg[7]  ( .D(n43003), .CP(clk), .Q(\filter_0/n17581 )
         );
  dff_sg \filter_0/oi_13_reg[8]  ( .D(n42991), .CP(clk), .Q(\filter_0/n17580 )
         );
  dff_sg \filter_0/oi_13_reg[9]  ( .D(n43002), .CP(clk), .Q(\filter_0/n17579 )
         );
  dff_sg \filter_0/oi_13_reg[10]  ( .D(n43001), .CP(clk), .Q(\filter_0/n17578 ) );
  dff_sg \filter_0/oi_13_reg[11]  ( .D(n43000), .CP(clk), .Q(\filter_0/n17577 ) );
  dff_sg \filter_0/oi_13_reg[12]  ( .D(n42990), .CP(clk), .Q(\filter_0/n17576 ) );
  dff_sg \filter_0/oi_13_reg[13]  ( .D(n42989), .CP(clk), .Q(\filter_0/n17575 ) );
  dff_sg \filter_0/oi_13_reg[14]  ( .D(n42995), .CP(clk), .Q(\filter_0/n17574 ) );
  dff_sg \filter_0/oi_13_reg[15]  ( .D(n42999), .CP(clk), .Q(\filter_0/n17573 ) );
  dff_sg \filter_0/oi_13_reg[16]  ( .D(n42998), .CP(clk), .Q(\filter_0/n17572 ) );
  dff_sg \filter_0/oi_13_reg[17]  ( .D(n42993), .CP(clk), .Q(\filter_0/n17571 ) );
  dff_sg \filter_0/oi_13_reg[18]  ( .D(n42996), .CP(clk), .Q(\filter_0/n17570 ) );
  dff_sg \filter_0/oi_13_reg[19]  ( .D(n42992), .CP(clk), .Q(\filter_0/n17569 ) );
  dff_sg \filter_0/oi_14_reg[0]  ( .D(n42988), .CP(clk), .Q(\filter_0/n17608 )
         );
  dff_sg \filter_0/oi_14_reg[1]  ( .D(n42987), .CP(clk), .Q(\filter_0/n17607 )
         );
  dff_sg \filter_0/oi_14_reg[2]  ( .D(n42973), .CP(clk), .Q(\filter_0/n17606 )
         );
  dff_sg \filter_0/oi_14_reg[3]  ( .D(n42977), .CP(clk), .Q(\filter_0/n17605 )
         );
  dff_sg \filter_0/oi_14_reg[4]  ( .D(n42986), .CP(clk), .Q(\filter_0/n17604 )
         );
  dff_sg \filter_0/oi_14_reg[5]  ( .D(n42985), .CP(clk), .Q(\filter_0/n17603 )
         );
  dff_sg \filter_0/oi_14_reg[6]  ( .D(n42970), .CP(clk), .Q(\filter_0/n17602 )
         );
  dff_sg \filter_0/oi_14_reg[7]  ( .D(n42984), .CP(clk), .Q(\filter_0/n17601 )
         );
  dff_sg \filter_0/oi_14_reg[8]  ( .D(n42983), .CP(clk), .Q(\filter_0/n17600 )
         );
  dff_sg \filter_0/oi_14_reg[9]  ( .D(n42982), .CP(clk), .Q(\filter_0/n17599 )
         );
  dff_sg \filter_0/oi_14_reg[10]  ( .D(n42981), .CP(clk), .Q(\filter_0/n17598 ) );
  dff_sg \filter_0/oi_14_reg[11]  ( .D(n42980), .CP(clk), .Q(\filter_0/n17597 ) );
  dff_sg \filter_0/oi_14_reg[12]  ( .D(n42971), .CP(clk), .Q(\filter_0/n17596 ) );
  dff_sg \filter_0/oi_14_reg[13]  ( .D(n42974), .CP(clk), .Q(\filter_0/n17595 ) );
  dff_sg \filter_0/oi_14_reg[14]  ( .D(n42975), .CP(clk), .Q(\filter_0/n17594 ) );
  dff_sg \filter_0/oi_14_reg[15]  ( .D(n42979), .CP(clk), .Q(\filter_0/n17593 ) );
  dff_sg \filter_0/oi_14_reg[16]  ( .D(n42978), .CP(clk), .Q(\filter_0/n17592 ) );
  dff_sg \filter_0/oi_14_reg[17]  ( .D(n42969), .CP(clk), .Q(\filter_0/n17591 ) );
  dff_sg \filter_0/oi_14_reg[18]  ( .D(n42976), .CP(clk), .Q(\filter_0/n17590 ) );
  dff_sg \filter_0/oi_14_reg[19]  ( .D(n42972), .CP(clk), .Q(\filter_0/n17589 ) );
  dff_sg \filter_0/oi_15_reg[0]  ( .D(n42868), .CP(clk), .Q(\filter_0/n17628 )
         );
  dff_sg \filter_0/oi_15_reg[1]  ( .D(n42861), .CP(clk), .Q(\filter_0/n17627 )
         );
  dff_sg \filter_0/oi_15_reg[2]  ( .D(n42867), .CP(clk), .Q(\filter_0/n17626 )
         );
  dff_sg \filter_0/oi_15_reg[3]  ( .D(n42860), .CP(clk), .Q(\filter_0/n17625 )
         );
  dff_sg \filter_0/oi_15_reg[4]  ( .D(n42866), .CP(clk), .Q(\filter_0/n17624 )
         );
  dff_sg \filter_0/oi_15_reg[5]  ( .D(n42859), .CP(clk), .Q(\filter_0/n17623 )
         );
  dff_sg \filter_0/oi_15_reg[6]  ( .D(n42865), .CP(clk), .Q(\filter_0/n17622 )
         );
  dff_sg \filter_0/oi_15_reg[7]  ( .D(n42858), .CP(clk), .Q(\filter_0/n17621 )
         );
  dff_sg \filter_0/oi_15_reg[8]  ( .D(n42864), .CP(clk), .Q(\filter_0/n17620 )
         );
  dff_sg \filter_0/oi_15_reg[9]  ( .D(n42857), .CP(clk), .Q(\filter_0/n17619 )
         );
  dff_sg \filter_0/oi_15_reg[10]  ( .D(n42863), .CP(clk), .Q(\filter_0/n17618 ) );
  dff_sg \filter_0/oi_15_reg[11]  ( .D(n42856), .CP(clk), .Q(\filter_0/n17617 ) );
  dff_sg \filter_0/oi_15_reg[12]  ( .D(n42862), .CP(clk), .Q(\filter_0/n17616 ) );
  dff_sg \filter_0/oi_15_reg[13]  ( .D(n42855), .CP(clk), .Q(\filter_0/n17615 ) );
  dff_sg \filter_0/oi_15_reg[14]  ( .D(n42853), .CP(clk), .Q(\filter_0/n17614 ) );
  dff_sg \filter_0/oi_15_reg[15]  ( .D(n42854), .CP(clk), .Q(\filter_0/n17613 ) );
  dff_sg \filter_0/oi_15_reg[16]  ( .D(n42852), .CP(clk), .Q(\filter_0/n17612 ) );
  dff_sg \filter_0/oi_15_reg[17]  ( .D(n42851), .CP(clk), .Q(\filter_0/n17611 ) );
  dff_sg \filter_0/oi_15_reg[18]  ( .D(n42850), .CP(clk), .Q(\filter_0/n17610 ) );
  dff_sg \filter_0/oi_15_reg[19]  ( .D(n42849), .CP(clk), .Q(\filter_0/n17609 ) );
  dff_sg \filter_0/oi_7_reg[0]  ( .D(n43208), .CP(clk), .Q(\filter_0/n17468 )
         );
  dff_sg \filter_0/oi_7_reg[1]  ( .D(n43189), .CP(clk), .Q(\filter_0/n17467 )
         );
  dff_sg \filter_0/oi_7_reg[2]  ( .D(n43207), .CP(clk), .Q(\filter_0/n17466 )
         );
  dff_sg \filter_0/oi_7_reg[3]  ( .D(n43197), .CP(clk), .Q(\filter_0/n17465 )
         );
  dff_sg \filter_0/oi_7_reg[4]  ( .D(n43206), .CP(clk), .Q(\filter_0/n17464 )
         );
  dff_sg \filter_0/oi_7_reg[5]  ( .D(n43193), .CP(clk), .Q(\filter_0/n17463 )
         );
  dff_sg \filter_0/oi_7_reg[6]  ( .D(n43205), .CP(clk), .Q(\filter_0/n17462 )
         );
  dff_sg \filter_0/oi_7_reg[7]  ( .D(n43191), .CP(clk), .Q(\filter_0/n17461 )
         );
  dff_sg \filter_0/oi_7_reg[8]  ( .D(n43204), .CP(clk), .Q(\filter_0/n17460 )
         );
  dff_sg \filter_0/oi_7_reg[9]  ( .D(n43194), .CP(clk), .Q(\filter_0/n17459 )
         );
  dff_sg \filter_0/oi_7_reg[10]  ( .D(n43203), .CP(clk), .Q(\filter_0/n17458 )
         );
  dff_sg \filter_0/oi_7_reg[11]  ( .D(n43190), .CP(clk), .Q(\filter_0/n17457 )
         );
  dff_sg \filter_0/oi_7_reg[12]  ( .D(n43202), .CP(clk), .Q(\filter_0/n17456 )
         );
  dff_sg \filter_0/oi_7_reg[13]  ( .D(n43201), .CP(clk), .Q(\filter_0/n17455 )
         );
  dff_sg \filter_0/oi_7_reg[14]  ( .D(n43195), .CP(clk), .Q(\filter_0/n17454 )
         );
  dff_sg \filter_0/oi_7_reg[15]  ( .D(n43192), .CP(clk), .Q(\filter_0/n17453 )
         );
  dff_sg \filter_0/oi_7_reg[16]  ( .D(n43200), .CP(clk), .Q(\filter_0/n17452 )
         );
  dff_sg \filter_0/oi_7_reg[17]  ( .D(n43199), .CP(clk), .Q(\filter_0/n17451 )
         );
  dff_sg \filter_0/oi_7_reg[18]  ( .D(n43196), .CP(clk), .Q(\filter_0/n17450 )
         );
  dff_sg \filter_0/oi_7_reg[19]  ( .D(n43198), .CP(clk), .Q(\filter_0/n17449 )
         );
  dff_sg \filter_0/oi_6_reg[0]  ( .D(n43188), .CP(clk), .Q(\filter_0/n17448 )
         );
  dff_sg \filter_0/oi_6_reg[1]  ( .D(n43187), .CP(clk), .Q(\filter_0/n17447 )
         );
  dff_sg \filter_0/oi_6_reg[2]  ( .D(n43186), .CP(clk), .Q(\filter_0/n17446 )
         );
  dff_sg \filter_0/oi_6_reg[3]  ( .D(n43177), .CP(clk), .Q(\filter_0/n17445 )
         );
  dff_sg \filter_0/oi_6_reg[4]  ( .D(n43185), .CP(clk), .Q(\filter_0/n17444 )
         );
  dff_sg \filter_0/oi_6_reg[5]  ( .D(n43184), .CP(clk), .Q(\filter_0/n17443 )
         );
  dff_sg \filter_0/oi_6_reg[6]  ( .D(n43174), .CP(clk), .Q(\filter_0/n17442 )
         );
  dff_sg \filter_0/oi_6_reg[7]  ( .D(n43183), .CP(clk), .Q(\filter_0/n17441 )
         );
  dff_sg \filter_0/oi_6_reg[8]  ( .D(n43171), .CP(clk), .Q(\filter_0/n17440 )
         );
  dff_sg \filter_0/oi_6_reg[9]  ( .D(n43182), .CP(clk), .Q(\filter_0/n17439 )
         );
  dff_sg \filter_0/oi_6_reg[10]  ( .D(n43181), .CP(clk), .Q(\filter_0/n17438 )
         );
  dff_sg \filter_0/oi_6_reg[11]  ( .D(n43180), .CP(clk), .Q(\filter_0/n17437 )
         );
  dff_sg \filter_0/oi_6_reg[12]  ( .D(n43170), .CP(clk), .Q(\filter_0/n17436 )
         );
  dff_sg \filter_0/oi_6_reg[13]  ( .D(n43169), .CP(clk), .Q(\filter_0/n17435 )
         );
  dff_sg \filter_0/oi_6_reg[14]  ( .D(n43175), .CP(clk), .Q(\filter_0/n17434 )
         );
  dff_sg \filter_0/oi_6_reg[15]  ( .D(n43179), .CP(clk), .Q(\filter_0/n17433 )
         );
  dff_sg \filter_0/oi_6_reg[16]  ( .D(n43178), .CP(clk), .Q(\filter_0/n17432 )
         );
  dff_sg \filter_0/oi_6_reg[17]  ( .D(n43173), .CP(clk), .Q(\filter_0/n17431 )
         );
  dff_sg \filter_0/oi_6_reg[18]  ( .D(n43176), .CP(clk), .Q(\filter_0/n17430 )
         );
  dff_sg \filter_0/oi_6_reg[19]  ( .D(n43172), .CP(clk), .Q(\filter_0/n17429 )
         );
  dff_sg \filter_0/oi_5_reg[0]  ( .D(n43248), .CP(clk), .Q(\filter_0/n17428 )
         );
  dff_sg \filter_0/oi_5_reg[1]  ( .D(n43247), .CP(clk), .Q(\filter_0/n17427 )
         );
  dff_sg \filter_0/oi_5_reg[2]  ( .D(n43233), .CP(clk), .Q(\filter_0/n17426 )
         );
  dff_sg \filter_0/oi_5_reg[3]  ( .D(n43237), .CP(clk), .Q(\filter_0/n17425 )
         );
  dff_sg \filter_0/oi_5_reg[4]  ( .D(n43246), .CP(clk), .Q(\filter_0/n17424 )
         );
  dff_sg \filter_0/oi_5_reg[5]  ( .D(n43245), .CP(clk), .Q(\filter_0/n17423 )
         );
  dff_sg \filter_0/oi_5_reg[6]  ( .D(n43230), .CP(clk), .Q(\filter_0/n17422 )
         );
  dff_sg \filter_0/oi_5_reg[7]  ( .D(n43244), .CP(clk), .Q(\filter_0/n17421 )
         );
  dff_sg \filter_0/oi_5_reg[8]  ( .D(n43243), .CP(clk), .Q(\filter_0/n17420 )
         );
  dff_sg \filter_0/oi_5_reg[9]  ( .D(n43242), .CP(clk), .Q(\filter_0/n17419 )
         );
  dff_sg \filter_0/oi_5_reg[10]  ( .D(n43241), .CP(clk), .Q(\filter_0/n17418 )
         );
  dff_sg \filter_0/oi_5_reg[11]  ( .D(n43240), .CP(clk), .Q(\filter_0/n17417 )
         );
  dff_sg \filter_0/oi_5_reg[12]  ( .D(n43231), .CP(clk), .Q(\filter_0/n17416 )
         );
  dff_sg \filter_0/oi_5_reg[13]  ( .D(n43234), .CP(clk), .Q(\filter_0/n17415 )
         );
  dff_sg \filter_0/oi_5_reg[14]  ( .D(n43235), .CP(clk), .Q(\filter_0/n17414 )
         );
  dff_sg \filter_0/oi_5_reg[15]  ( .D(n43239), .CP(clk), .Q(\filter_0/n17413 )
         );
  dff_sg \filter_0/oi_5_reg[16]  ( .D(n43238), .CP(clk), .Q(\filter_0/n17412 )
         );
  dff_sg \filter_0/oi_5_reg[17]  ( .D(n43229), .CP(clk), .Q(\filter_0/n17411 )
         );
  dff_sg \filter_0/oi_5_reg[18]  ( .D(n43236), .CP(clk), .Q(\filter_0/n17410 )
         );
  dff_sg \filter_0/oi_5_reg[19]  ( .D(n43232), .CP(clk), .Q(\filter_0/n17409 )
         );
  dff_sg \filter_0/oi_4_reg[0]  ( .D(n43228), .CP(clk), .Q(\filter_0/n17408 )
         );
  dff_sg \filter_0/oi_4_reg[1]  ( .D(n43227), .CP(clk), .Q(\filter_0/n17407 )
         );
  dff_sg \filter_0/oi_4_reg[2]  ( .D(n43213), .CP(clk), .Q(\filter_0/n17406 )
         );
  dff_sg \filter_0/oi_4_reg[3]  ( .D(n43217), .CP(clk), .Q(\filter_0/n17405 )
         );
  dff_sg \filter_0/oi_4_reg[4]  ( .D(n43226), .CP(clk), .Q(\filter_0/n17404 )
         );
  dff_sg \filter_0/oi_4_reg[5]  ( .D(n43225), .CP(clk), .Q(\filter_0/n17403 )
         );
  dff_sg \filter_0/oi_4_reg[6]  ( .D(n43210), .CP(clk), .Q(\filter_0/n17402 )
         );
  dff_sg \filter_0/oi_4_reg[7]  ( .D(n43224), .CP(clk), .Q(\filter_0/n17401 )
         );
  dff_sg \filter_0/oi_4_reg[8]  ( .D(n43223), .CP(clk), .Q(\filter_0/n17400 )
         );
  dff_sg \filter_0/oi_4_reg[9]  ( .D(n43222), .CP(clk), .Q(\filter_0/n17399 )
         );
  dff_sg \filter_0/oi_4_reg[10]  ( .D(n43221), .CP(clk), .Q(\filter_0/n17398 )
         );
  dff_sg \filter_0/oi_4_reg[11]  ( .D(n43220), .CP(clk), .Q(\filter_0/n17397 )
         );
  dff_sg \filter_0/oi_4_reg[12]  ( .D(n43211), .CP(clk), .Q(\filter_0/n17396 )
         );
  dff_sg \filter_0/oi_4_reg[13]  ( .D(n43214), .CP(clk), .Q(\filter_0/n17395 )
         );
  dff_sg \filter_0/oi_4_reg[14]  ( .D(n43215), .CP(clk), .Q(\filter_0/n17394 )
         );
  dff_sg \filter_0/oi_4_reg[15]  ( .D(n43219), .CP(clk), .Q(\filter_0/n17393 )
         );
  dff_sg \filter_0/oi_4_reg[16]  ( .D(n43218), .CP(clk), .Q(\filter_0/n17392 )
         );
  dff_sg \filter_0/oi_4_reg[17]  ( .D(n43209), .CP(clk), .Q(\filter_0/n17391 )
         );
  dff_sg \filter_0/oi_4_reg[18]  ( .D(n43216), .CP(clk), .Q(\filter_0/n17390 )
         );
  dff_sg \filter_0/oi_4_reg[19]  ( .D(n43212), .CP(clk), .Q(\filter_0/n17389 )
         );
  dff_sg \filter_0/oi_3_reg[0]  ( .D(n42888), .CP(clk), .Q(\filter_0/n17388 )
         );
  dff_sg \filter_0/oi_3_reg[1]  ( .D(n42874), .CP(clk), .Q(\filter_0/n17387 )
         );
  dff_sg \filter_0/oi_3_reg[2]  ( .D(n42887), .CP(clk), .Q(\filter_0/n17386 )
         );
  dff_sg \filter_0/oi_3_reg[3]  ( .D(n42877), .CP(clk), .Q(\filter_0/n17385 )
         );
  dff_sg \filter_0/oi_3_reg[4]  ( .D(n42886), .CP(clk), .Q(\filter_0/n17384 )
         );
  dff_sg \filter_0/oi_3_reg[5]  ( .D(n42873), .CP(clk), .Q(\filter_0/n17383 )
         );
  dff_sg \filter_0/oi_3_reg[6]  ( .D(n42885), .CP(clk), .Q(\filter_0/n17382 )
         );
  dff_sg \filter_0/oi_3_reg[7]  ( .D(n42884), .CP(clk), .Q(\filter_0/n17381 )
         );
  dff_sg \filter_0/oi_3_reg[8]  ( .D(n42883), .CP(clk), .Q(\filter_0/n17380 )
         );
  dff_sg \filter_0/oi_3_reg[9]  ( .D(n42882), .CP(clk), .Q(\filter_0/n17379 )
         );
  dff_sg \filter_0/oi_3_reg[10]  ( .D(n42881), .CP(clk), .Q(\filter_0/n17378 )
         );
  dff_sg \filter_0/oi_3_reg[11]  ( .D(n42869), .CP(clk), .Q(\filter_0/n17377 )
         );
  dff_sg \filter_0/oi_3_reg[12]  ( .D(n42880), .CP(clk), .Q(\filter_0/n17376 )
         );
  dff_sg \filter_0/oi_3_reg[13]  ( .D(n42871), .CP(clk), .Q(\filter_0/n17375 )
         );
  dff_sg \filter_0/oi_3_reg[14]  ( .D(n42875), .CP(clk), .Q(\filter_0/n17374 )
         );
  dff_sg \filter_0/oi_3_reg[15]  ( .D(n42879), .CP(clk), .Q(\filter_0/n17373 )
         );
  dff_sg \filter_0/oi_3_reg[16]  ( .D(n42870), .CP(clk), .Q(\filter_0/n17372 )
         );
  dff_sg \filter_0/oi_3_reg[17]  ( .D(n42872), .CP(clk), .Q(\filter_0/n17371 )
         );
  dff_sg \filter_0/oi_3_reg[18]  ( .D(n42876), .CP(clk), .Q(\filter_0/n17370 )
         );
  dff_sg \filter_0/oi_3_reg[19]  ( .D(n42878), .CP(clk), .Q(\filter_0/n17369 )
         );
  dff_sg \filter_0/oi_2_reg[0]  ( .D(n42968), .CP(clk), .Q(\filter_0/n17368 )
         );
  dff_sg \filter_0/oi_2_reg[1]  ( .D(n42967), .CP(clk), .Q(\filter_0/n17367 )
         );
  dff_sg \filter_0/oi_2_reg[2]  ( .D(n42953), .CP(clk), .Q(\filter_0/n17366 )
         );
  dff_sg \filter_0/oi_2_reg[3]  ( .D(n42957), .CP(clk), .Q(\filter_0/n17365 )
         );
  dff_sg \filter_0/oi_2_reg[4]  ( .D(n42966), .CP(clk), .Q(\filter_0/n17364 )
         );
  dff_sg \filter_0/oi_2_reg[5]  ( .D(n42965), .CP(clk), .Q(\filter_0/n17363 )
         );
  dff_sg \filter_0/oi_2_reg[6]  ( .D(n42950), .CP(clk), .Q(\filter_0/n17362 )
         );
  dff_sg \filter_0/oi_2_reg[7]  ( .D(n42964), .CP(clk), .Q(\filter_0/n17361 )
         );
  dff_sg \filter_0/oi_2_reg[8]  ( .D(n42963), .CP(clk), .Q(\filter_0/n17360 )
         );
  dff_sg \filter_0/oi_2_reg[9]  ( .D(n42962), .CP(clk), .Q(\filter_0/n17359 )
         );
  dff_sg \filter_0/oi_2_reg[10]  ( .D(n42961), .CP(clk), .Q(\filter_0/n17358 )
         );
  dff_sg \filter_0/oi_2_reg[11]  ( .D(n42960), .CP(clk), .Q(\filter_0/n17357 )
         );
  dff_sg \filter_0/oi_2_reg[12]  ( .D(n42951), .CP(clk), .Q(\filter_0/n17356 )
         );
  dff_sg \filter_0/oi_2_reg[13]  ( .D(n42954), .CP(clk), .Q(\filter_0/n17355 )
         );
  dff_sg \filter_0/oi_2_reg[14]  ( .D(n42955), .CP(clk), .Q(\filter_0/n17354 )
         );
  dff_sg \filter_0/oi_2_reg[15]  ( .D(n42959), .CP(clk), .Q(\filter_0/n17353 )
         );
  dff_sg \filter_0/oi_2_reg[16]  ( .D(n42958), .CP(clk), .Q(\filter_0/n17352 )
         );
  dff_sg \filter_0/oi_2_reg[17]  ( .D(n42949), .CP(clk), .Q(\filter_0/n17351 )
         );
  dff_sg \filter_0/oi_2_reg[18]  ( .D(n42956), .CP(clk), .Q(\filter_0/n17350 )
         );
  dff_sg \filter_0/oi_2_reg[19]  ( .D(n42952), .CP(clk), .Q(\filter_0/n17349 )
         );
  dff_sg \filter_0/oi_1_reg[0]  ( .D(n43436), .CP(clk), .Q(\filter_0/n17348 )
         );
  dff_sg \filter_0/oi_1_reg[1]  ( .D(n43448), .CP(clk), .Q(\filter_0/n17347 )
         );
  dff_sg \filter_0/oi_1_reg[2]  ( .D(n43431), .CP(clk), .Q(\filter_0/n17346 )
         );
  dff_sg \filter_0/oi_1_reg[3]  ( .D(n43441), .CP(clk), .Q(\filter_0/n17345 )
         );
  dff_sg \filter_0/oi_1_reg[4]  ( .D(n43433), .CP(clk), .Q(\filter_0/n17344 )
         );
  dff_sg \filter_0/oi_1_reg[5]  ( .D(n43447), .CP(clk), .Q(\filter_0/n17343 )
         );
  dff_sg \filter_0/oi_1_reg[6]  ( .D(n43438), .CP(clk), .Q(\filter_0/n17342 )
         );
  dff_sg \filter_0/oi_1_reg[7]  ( .D(n43429), .CP(clk), .Q(\filter_0/n17341 )
         );
  dff_sg \filter_0/oi_1_reg[8]  ( .D(n43446), .CP(clk), .Q(\filter_0/n17340 )
         );
  dff_sg \filter_0/oi_1_reg[9]  ( .D(n43445), .CP(clk), .Q(\filter_0/n17339 )
         );
  dff_sg \filter_0/oi_1_reg[10]  ( .D(n43444), .CP(clk), .Q(\filter_0/n17338 )
         );
  dff_sg \filter_0/oi_1_reg[11]  ( .D(n43443), .CP(clk), .Q(\filter_0/n17337 )
         );
  dff_sg \filter_0/oi_1_reg[12]  ( .D(n43439), .CP(clk), .Q(\filter_0/n17336 )
         );
  dff_sg \filter_0/oi_1_reg[13]  ( .D(n43437), .CP(clk), .Q(\filter_0/n17335 )
         );
  dff_sg \filter_0/oi_1_reg[14]  ( .D(n43434), .CP(clk), .Q(\filter_0/n17334 )
         );
  dff_sg \filter_0/oi_1_reg[15]  ( .D(n43442), .CP(clk), .Q(\filter_0/n17333 )
         );
  dff_sg \filter_0/oi_1_reg[16]  ( .D(n43435), .CP(clk), .Q(\filter_0/n17332 )
         );
  dff_sg \filter_0/oi_1_reg[17]  ( .D(n43430), .CP(clk), .Q(\filter_0/n17331 )
         );
  dff_sg \filter_0/oi_1_reg[18]  ( .D(n43440), .CP(clk), .Q(\filter_0/n17330 )
         );
  dff_sg \filter_0/oi_1_reg[19]  ( .D(n43432), .CP(clk), .Q(\filter_0/n17329 )
         );
  dff_sg \filter_0/input_taken_reg  ( .D(\filter_0/n12237 ), .CP(clk), .Q(
        \filter_0/n17951 ) );
  dff_sg \filter_0/reg_i_0_reg[0]  ( .D(n43530), .CP(clk), .Q(
        \filter_0/reg_i_0 [0]) );
  dff_sg \filter_0/reg_i_0_reg[1]  ( .D(n43720), .CP(clk), .Q(
        \filter_0/reg_i_0 [1]) );
  dff_sg \filter_0/reg_i_0_reg[2]  ( .D(n43747), .CP(clk), .Q(
        \filter_0/reg_i_0 [2]) );
  dff_sg \filter_0/reg_i_0_reg[3]  ( .D(n43735), .CP(clk), .Q(
        \filter_0/reg_i_0 [3]) );
  dff_sg \filter_0/reg_i_0_reg[4]  ( .D(n43494), .CP(clk), .Q(
        \filter_0/reg_i_0 [4]) );
  dff_sg \filter_0/reg_i_0_reg[5]  ( .D(n43537), .CP(clk), .Q(
        \filter_0/reg_i_0 [5]) );
  dff_sg \filter_0/reg_i_0_reg[6]  ( .D(n43492), .CP(clk), .Q(
        \filter_0/reg_i_0 [6]) );
  dff_sg \filter_0/reg_i_0_reg[7]  ( .D(n43927), .CP(clk), .Q(
        \filter_0/reg_i_0 [7]) );
  dff_sg \filter_0/reg_i_0_reg[8]  ( .D(n43524), .CP(clk), .Q(
        \filter_0/reg_i_0 [8]) );
  dff_sg \filter_0/reg_i_0_reg[9]  ( .D(n43753), .CP(clk), .Q(
        \filter_0/reg_i_0 [9]) );
  dff_sg \filter_0/reg_i_0_reg[10]  ( .D(n43491), .CP(clk), .Q(
        \filter_0/reg_i_0 [10]) );
  dff_sg \filter_0/reg_i_0_reg[11]  ( .D(n43528), .CP(clk), .Q(
        \filter_0/reg_i_0 [11]) );
  dff_sg \filter_0/reg_i_0_reg[12]  ( .D(n43721), .CP(clk), .Q(
        \filter_0/reg_i_0 [12]) );
  dff_sg \filter_0/reg_i_0_reg[13]  ( .D(n43722), .CP(clk), .Q(
        \filter_0/reg_i_0 [13]) );
  dff_sg \filter_0/reg_i_0_reg[14]  ( .D(n43718), .CP(clk), .Q(
        \filter_0/reg_i_0 [14]) );
  dff_sg \filter_0/reg_i_0_reg[15]  ( .D(n43719), .CP(clk), .Q(
        \filter_0/reg_i_0 [15]) );
  dff_sg \filter_0/reg_i_0_reg[16]  ( .D(n43727), .CP(clk), .Q(
        \filter_0/reg_i_0 [16]) );
  dff_sg \filter_0/reg_i_0_reg[17]  ( .D(n43728), .CP(clk), .Q(
        \filter_0/reg_i_0 [17]) );
  dff_sg \filter_0/reg_i_0_reg[18]  ( .D(n43724), .CP(clk), .Q(
        \filter_0/reg_i_0 [18]) );
  dff_sg \filter_0/reg_i_0_reg[19]  ( .D(n43725), .CP(clk), .Q(
        \filter_0/reg_i_0 [19]) );
  dff_sg \filter_0/reg_i_1_reg[0]  ( .D(n43709), .CP(clk), .Q(
        \filter_0/reg_i_1 [0]) );
  dff_sg \filter_0/reg_i_1_reg[1]  ( .D(n43710), .CP(clk), .Q(
        \filter_0/reg_i_1 [1]) );
  dff_sg \filter_0/reg_i_1_reg[2]  ( .D(n43706), .CP(clk), .Q(
        \filter_0/reg_i_1 [2]) );
  dff_sg \filter_0/reg_i_1_reg[3]  ( .D(n43707), .CP(clk), .Q(
        \filter_0/reg_i_1 [3]) );
  dff_sg \filter_0/reg_i_1_reg[4]  ( .D(n43715), .CP(clk), .Q(
        \filter_0/reg_i_1 [4]) );
  dff_sg \filter_0/reg_i_1_reg[5]  ( .D(n43716), .CP(clk), .Q(
        \filter_0/reg_i_1 [5]) );
  dff_sg \filter_0/reg_i_1_reg[6]  ( .D(n43712), .CP(clk), .Q(
        \filter_0/reg_i_1 [6]) );
  dff_sg \filter_0/reg_i_1_reg[7]  ( .D(n43713), .CP(clk), .Q(
        \filter_0/reg_i_1 [7]) );
  dff_sg \filter_0/reg_i_1_reg[8]  ( .D(n43745), .CP(clk), .Q(
        \filter_0/reg_i_1 [8]) );
  dff_sg \filter_0/reg_i_1_reg[9]  ( .D(n43746), .CP(clk), .Q(
        \filter_0/reg_i_1 [9]) );
  dff_sg \filter_0/reg_i_1_reg[10]  ( .D(n43742), .CP(clk), .Q(
        \filter_0/reg_i_1 [10]) );
  dff_sg \filter_0/reg_i_1_reg[11]  ( .D(n43743), .CP(clk), .Q(
        \filter_0/reg_i_1 [11]) );
  dff_sg \filter_0/reg_i_1_reg[12]  ( .D(n43751), .CP(clk), .Q(
        \filter_0/reg_i_1 [12]) );
  dff_sg \filter_0/reg_i_1_reg[13]  ( .D(n43752), .CP(clk), .Q(
        \filter_0/reg_i_1 [13]) );
  dff_sg \filter_0/reg_i_1_reg[14]  ( .D(n43748), .CP(clk), .Q(
        \filter_0/reg_i_1 [14]) );
  dff_sg \filter_0/reg_i_1_reg[15]  ( .D(n43749), .CP(clk), .Q(
        \filter_0/reg_i_1 [15]) );
  dff_sg \filter_0/reg_i_1_reg[16]  ( .D(n43733), .CP(clk), .Q(
        \filter_0/reg_i_1 [16]) );
  dff_sg \filter_0/reg_i_1_reg[17]  ( .D(n43734), .CP(clk), .Q(
        \filter_0/reg_i_1 [17]) );
  dff_sg \filter_0/reg_i_1_reg[18]  ( .D(n43730), .CP(clk), .Q(
        \filter_0/reg_i_1 [18]) );
  dff_sg \filter_0/reg_i_1_reg[19]  ( .D(n43731), .CP(clk), .Q(
        \filter_0/reg_i_1 [19]) );
  dff_sg \filter_0/reg_i_2_reg[0]  ( .D(n43739), .CP(clk), .Q(
        \filter_0/reg_i_2 [0]) );
  dff_sg \filter_0/reg_i_2_reg[1]  ( .D(n43740), .CP(clk), .Q(
        \filter_0/reg_i_2 [1]) );
  dff_sg \filter_0/reg_i_2_reg[2]  ( .D(n43736), .CP(clk), .Q(
        \filter_0/reg_i_2 [2]) );
  dff_sg \filter_0/reg_i_2_reg[3]  ( .D(n43737), .CP(clk), .Q(
        \filter_0/reg_i_2 [3]) );
  dff_sg \filter_0/reg_i_2_reg[4]  ( .D(n43557), .CP(clk), .Q(
        \filter_0/reg_i_2 [4]) );
  dff_sg \filter_0/reg_i_2_reg[5]  ( .D(n43498), .CP(clk), .Q(
        \filter_0/reg_i_2 [5]) );
  dff_sg \filter_0/reg_i_2_reg[6]  ( .D(n43507), .CP(clk), .Q(
        \filter_0/reg_i_2 [6]) );
  dff_sg \filter_0/reg_i_2_reg[7]  ( .D(n43546), .CP(clk), .Q(
        \filter_0/reg_i_2 [7]) );
  dff_sg \filter_0/reg_i_2_reg[8]  ( .D(n43540), .CP(clk), .Q(
        \filter_0/reg_i_2 [8]) );
  dff_sg \filter_0/reg_i_2_reg[9]  ( .D(n43504), .CP(clk), .Q(
        \filter_0/reg_i_2 [9]) );
  dff_sg \filter_0/reg_i_2_reg[10]  ( .D(n43501), .CP(clk), .Q(
        \filter_0/reg_i_2 [10]) );
  dff_sg \filter_0/reg_i_2_reg[11]  ( .D(n44102), .CP(clk), .Q(
        \filter_0/reg_i_2 [11]) );
  dff_sg \filter_0/reg_i_2_reg[12]  ( .D(n43543), .CP(clk), .Q(
        \filter_0/reg_i_2 [12]) );
  dff_sg \filter_0/reg_i_2_reg[13]  ( .D(n43552), .CP(clk), .Q(
        \filter_0/reg_i_2 [13]) );
  dff_sg \filter_0/reg_i_2_reg[14]  ( .D(n43512), .CP(clk), .Q(
        \filter_0/reg_i_2 [14]) );
  dff_sg \filter_0/reg_i_2_reg[15]  ( .D(n43556), .CP(clk), .Q(
        \filter_0/reg_i_2 [15]) );
  dff_sg \filter_0/reg_i_2_reg[16]  ( .D(n43511), .CP(clk), .Q(
        \filter_0/reg_i_2 [16]) );
  dff_sg \filter_0/reg_i_2_reg[17]  ( .D(n43519), .CP(clk), .Q(
        \filter_0/reg_i_2 [17]) );
  dff_sg \filter_0/reg_i_2_reg[18]  ( .D(n43510), .CP(clk), .Q(
        \filter_0/reg_i_2 [18]) );
  dff_sg \filter_0/reg_i_2_reg[19]  ( .D(n44060), .CP(clk), .Q(
        \filter_0/reg_i_2 [19]) );
  dff_sg \filter_0/reg_i_3_reg[0]  ( .D(n43570), .CP(clk), .Q(
        \filter_0/reg_i_3 [0]) );
  dff_sg \filter_0/reg_i_3_reg[1]  ( .D(n43582), .CP(clk), .Q(
        \filter_0/reg_i_3 [1]) );
  dff_sg \filter_0/reg_i_3_reg[2]  ( .D(n43518), .CP(clk), .Q(
        \filter_0/reg_i_3 [2]) );
  dff_sg \filter_0/reg_i_3_reg[3]  ( .D(n43579), .CP(clk), .Q(
        \filter_0/reg_i_3 [3]) );
  dff_sg \filter_0/reg_i_3_reg[4]  ( .D(n43588), .CP(clk), .Q(
        \filter_0/reg_i_3 [4]) );
  dff_sg \filter_0/reg_i_3_reg[5]  ( .D(n43591), .CP(clk), .Q(
        \filter_0/reg_i_3 [5]) );
  dff_sg \filter_0/reg_i_3_reg[6]  ( .D(n43517), .CP(clk), .Q(
        \filter_0/reg_i_3 [6]) );
  dff_sg \filter_0/reg_i_3_reg[7]  ( .D(n43516), .CP(clk), .Q(
        \filter_0/reg_i_3 [7]) );
  dff_sg \filter_0/reg_i_3_reg[8]  ( .D(n43573), .CP(clk), .Q(
        \filter_0/reg_i_3 [8]) );
  dff_sg \filter_0/reg_i_3_reg[9]  ( .D(n43576), .CP(clk), .Q(
        \filter_0/reg_i_3 [9]) );
  dff_sg \filter_0/reg_i_3_reg[10]  ( .D(n43514), .CP(clk), .Q(
        \filter_0/reg_i_3 [10]) );
  dff_sg \filter_0/reg_i_3_reg[11]  ( .D(n43513), .CP(clk), .Q(
        \filter_0/reg_i_3 [11]) );
  dff_sg \filter_0/reg_i_3_reg[12]  ( .D(n44096), .CP(clk), .Q(
        \filter_0/reg_i_3 [12]) );
  dff_sg \filter_0/reg_i_3_reg[13]  ( .D(n43564), .CP(clk), .Q(
        \filter_0/reg_i_3 [13]) );
  dff_sg \filter_0/reg_i_3_reg[14]  ( .D(n43515), .CP(clk), .Q(
        \filter_0/reg_i_3 [14]) );
  dff_sg \filter_0/reg_i_3_reg[15]  ( .D(n43567), .CP(clk), .Q(
        \filter_0/reg_i_3 [15]) );
  dff_sg \filter_0/reg_i_3_reg[16]  ( .D(n43828), .CP(clk), .Q(
        \filter_0/reg_i_3 [16]) );
  dff_sg \filter_0/reg_i_3_reg[17]  ( .D(n43816), .CP(clk), .Q(
        \filter_0/reg_i_3 [17]) );
  dff_sg \filter_0/reg_i_3_reg[18]  ( .D(n43801), .CP(clk), .Q(
        \filter_0/reg_i_3 [18]) );
  dff_sg \filter_0/reg_i_3_reg[19]  ( .D(n43834), .CP(clk), .Q(
        \filter_0/reg_i_3 [19]) );
  dff_sg \filter_0/reg_i_4_reg[0]  ( .D(n43780), .CP(clk), .Q(
        \filter_0/reg_i_4 [0]) );
  dff_sg \filter_0/reg_i_4_reg[1]  ( .D(n43771), .CP(clk), .Q(
        \filter_0/reg_i_4 [1]) );
  dff_sg \filter_0/reg_i_4_reg[2]  ( .D(n43975), .CP(clk), .Q(
        \filter_0/reg_i_4 [2]) );
  dff_sg \filter_0/reg_i_4_reg[3]  ( .D(n43777), .CP(clk), .Q(
        \filter_0/reg_i_4 [3]) );
  dff_sg \filter_0/reg_i_4_reg[4]  ( .D(n43738), .CP(clk), .Q(
        \filter_0/reg_i_4 [4]) );
  dff_sg \filter_0/reg_i_4_reg[5]  ( .D(n43741), .CP(clk), .Q(
        \filter_0/reg_i_4 [5]) );
  dff_sg \filter_0/reg_i_4_reg[6]  ( .D(n43750), .CP(clk), .Q(
        \filter_0/reg_i_4 [6]) );
  dff_sg \filter_0/reg_i_4_reg[7]  ( .D(n43744), .CP(clk), .Q(
        \filter_0/reg_i_4 [7]) );
  dff_sg \filter_0/reg_i_4_reg[8]  ( .D(n43723), .CP(clk), .Q(
        \filter_0/reg_i_4 [8]) );
  dff_sg \filter_0/reg_i_4_reg[9]  ( .D(n43726), .CP(clk), .Q(
        \filter_0/reg_i_4 [9]) );
  dff_sg \filter_0/reg_i_4_reg[10]  ( .D(n43729), .CP(clk), .Q(
        \filter_0/reg_i_4 [10]) );
  dff_sg \filter_0/reg_i_4_reg[11]  ( .D(n43732), .CP(clk), .Q(
        \filter_0/reg_i_4 [11]) );
  dff_sg \filter_0/reg_i_4_reg[12]  ( .D(n43837), .CP(clk), .Q(
        \filter_0/reg_i_4 [12]) );
  dff_sg \filter_0/reg_i_4_reg[13]  ( .D(n43495), .CP(clk), .Q(
        \filter_0/reg_i_4 [13]) );
  dff_sg \filter_0/reg_i_4_reg[14]  ( .D(n44105), .CP(clk), .Q(
        \filter_0/reg_i_4 [14]) );
  dff_sg \filter_0/reg_i_4_reg[15]  ( .D(n43497), .CP(clk), .Q(
        \filter_0/reg_i_4 [15]) );
  dff_sg \filter_0/reg_i_4_reg[16]  ( .D(n43980), .CP(clk), .Q(
        \filter_0/reg_i_4 [16]) );
  dff_sg \filter_0/reg_i_4_reg[17]  ( .D(n43558), .CP(clk), .Q(
        \filter_0/reg_i_4 [17]) );
  dff_sg \filter_0/reg_i_4_reg[18]  ( .D(n43496), .CP(clk), .Q(
        \filter_0/reg_i_4 [18]) );
  dff_sg \filter_0/reg_i_4_reg[19]  ( .D(n43561), .CP(clk), .Q(
        \filter_0/reg_i_4 [19]) );
  dff_sg \filter_0/reg_i_5_reg[0]  ( .D(n43948), .CP(clk), .Q(
        \filter_0/reg_i_5 [0]) );
  dff_sg \filter_0/reg_i_5_reg[1]  ( .D(n43545), .CP(clk), .Q(
        \filter_0/reg_i_5 [1]) );
  dff_sg \filter_0/reg_i_5_reg[2]  ( .D(n43493), .CP(clk), .Q(
        \filter_0/reg_i_5 [2]) );
  dff_sg \filter_0/reg_i_5_reg[3]  ( .D(n43950), .CP(clk), .Q(
        \filter_0/reg_i_5 [3]) );
  dff_sg \filter_0/reg_i_5_reg[4]  ( .D(n43894), .CP(clk), .Q(
        \filter_0/reg_i_5 [4]) );
  dff_sg \filter_0/reg_i_5_reg[5]  ( .D(n43882), .CP(clk), .Q(
        \filter_0/reg_i_5 [5]) );
  dff_sg \filter_0/reg_i_5_reg[6]  ( .D(n43900), .CP(clk), .Q(
        \filter_0/reg_i_5 [6]) );
  dff_sg \filter_0/reg_i_5_reg[7]  ( .D(n43939), .CP(clk), .Q(
        \filter_0/reg_i_5 [7]) );
  dff_sg \filter_0/reg_i_5_reg[8]  ( .D(n43539), .CP(clk), .Q(
        \filter_0/reg_i_5 [8]) );
  dff_sg \filter_0/reg_i_5_reg[9]  ( .D(n43856), .CP(clk), .Q(
        \filter_0/reg_i_5 [9]) );
  dff_sg \filter_0/reg_i_5_reg[10]  ( .D(n43487), .CP(clk), .Q(
        \filter_0/reg_i_5 [10]) );
  dff_sg \filter_0/reg_i_5_reg[11]  ( .D(n43680), .CP(clk), .Q(
        \filter_0/reg_i_5 [11]) );
  dff_sg \filter_0/reg_i_5_reg[12]  ( .D(n43694), .CP(clk), .Q(
        \filter_0/reg_i_5 [12]) );
  dff_sg \filter_0/reg_i_5_reg[13]  ( .D(n43697), .CP(clk), .Q(
        \filter_0/reg_i_5 [13]) );
  dff_sg \filter_0/reg_i_5_reg[14]  ( .D(n43485), .CP(clk), .Q(
        \filter_0/reg_i_5 [14]) );
  dff_sg \filter_0/reg_i_5_reg[15]  ( .D(n43486), .CP(clk), .Q(
        \filter_0/reg_i_5 [15]) );
  dff_sg \filter_0/reg_i_5_reg[16]  ( .D(n43671), .CP(clk), .Q(
        \filter_0/reg_i_5 [16]) );
  dff_sg \filter_0/reg_i_5_reg[17]  ( .D(n43674), .CP(clk), .Q(
        \filter_0/reg_i_5 [17]) );
  dff_sg \filter_0/reg_i_5_reg[18]  ( .D(n43474), .CP(clk), .Q(
        \filter_0/reg_i_5 [18]) );
  dff_sg \filter_0/reg_i_5_reg[19]  ( .D(n43685), .CP(clk), .Q(
        \filter_0/reg_i_5 [19]) );
  dff_sg \filter_0/reg_i_6_reg[0]  ( .D(n43668), .CP(clk), .Q(
        \filter_0/reg_i_6 [0]) );
  dff_sg \filter_0/reg_i_6_reg[1]  ( .D(n43677), .CP(clk), .Q(
        \filter_0/reg_i_6 [1]) );
  dff_sg \filter_0/reg_i_6_reg[2]  ( .D(n43688), .CP(clk), .Q(
        \filter_0/reg_i_6 [2]) );
  dff_sg \filter_0/reg_i_6_reg[3]  ( .D(n43665), .CP(clk), .Q(
        \filter_0/reg_i_6 [3]) );
  dff_sg \filter_0/reg_i_6_reg[4]  ( .D(n44028), .CP(clk), .Q(
        \filter_0/reg_i_6 [4]) );
  dff_sg \filter_0/reg_i_6_reg[5]  ( .D(n44018), .CP(clk), .Q(
        \filter_0/reg_i_6 [5]) );
  dff_sg \filter_0/reg_i_6_reg[6]  ( .D(n43999), .CP(clk), .Q(
        \filter_0/reg_i_6 [6]) );
  dff_sg \filter_0/reg_i_6_reg[7]  ( .D(n44005), .CP(clk), .Q(
        \filter_0/reg_i_6 [7]) );
  dff_sg \filter_0/reg_i_6_reg[8]  ( .D(n43903), .CP(clk), .Q(
        \filter_0/reg_i_6 [8]) );
  dff_sg \filter_0/reg_i_6_reg[9]  ( .D(n44008), .CP(clk), .Q(
        \filter_0/reg_i_6 [9]) );
  dff_sg \filter_0/reg_i_6_reg[10]  ( .D(n43549), .CP(clk), .Q(
        \filter_0/reg_i_6 [10]) );
  dff_sg \filter_0/reg_i_6_reg[11]  ( .D(n43945), .CP(clk), .Q(
        \filter_0/reg_i_6 [11]) );
  dff_sg \filter_0/reg_i_6_reg[12]  ( .D(n43702), .CP(clk), .Q(
        \filter_0/reg_i_6 [12]) );
  dff_sg \filter_0/reg_i_6_reg[13]  ( .D(n43691), .CP(clk), .Q(
        \filter_0/reg_i_6 [13]) );
  dff_sg \filter_0/reg_i_6_reg[14]  ( .D(n44108), .CP(clk), .Q(
        \filter_0/reg_i_6 [14]) );
  dff_sg \filter_0/reg_i_6_reg[15]  ( .D(n44025), .CP(clk), .Q(
        \filter_0/reg_i_6 [15]) );
  dff_sg \filter_0/reg_i_6_reg[16]  ( .D(n44057), .CP(clk), .Q(
        \filter_0/reg_i_6 [16]) );
  dff_sg \filter_0/reg_i_6_reg[17]  ( .D(n43789), .CP(clk), .Q(
        \filter_0/reg_i_6 [17]) );
  dff_sg \filter_0/reg_i_6_reg[18]  ( .D(n43798), .CP(clk), .Q(
        \filter_0/reg_i_6 [18]) );
  dff_sg \filter_0/reg_i_6_reg[19]  ( .D(n44109), .CP(clk), .Q(
        \filter_0/reg_i_6 [19]) );
  dff_sg \filter_0/reg_i_7_reg[0]  ( .D(n43600), .CP(clk), .Q(
        \filter_0/reg_i_7 [0]) );
  dff_sg \filter_0/reg_i_7_reg[1]  ( .D(n43624), .CP(clk), .Q(
        \filter_0/reg_i_7 [1]) );
  dff_sg \filter_0/reg_i_7_reg[2]  ( .D(n43609), .CP(clk), .Q(
        \filter_0/reg_i_7 [2]) );
  dff_sg \filter_0/reg_i_7_reg[3]  ( .D(n43606), .CP(clk), .Q(
        \filter_0/reg_i_7 [3]) );
  dff_sg \filter_0/reg_i_7_reg[4]  ( .D(n43615), .CP(clk), .Q(
        \filter_0/reg_i_7 [4]) );
  dff_sg \filter_0/reg_i_7_reg[5]  ( .D(n43627), .CP(clk), .Q(
        \filter_0/reg_i_7 [5]) );
  dff_sg \filter_0/reg_i_7_reg[6]  ( .D(n43612), .CP(clk), .Q(
        \filter_0/reg_i_7 [6]) );
  dff_sg \filter_0/reg_i_7_reg[7]  ( .D(n43603), .CP(clk), .Q(
        \filter_0/reg_i_7 [7]) );
  dff_sg \filter_0/reg_i_7_reg[8]  ( .D(n43585), .CP(clk), .Q(
        \filter_0/reg_i_7 [8]) );
  dff_sg \filter_0/reg_i_7_reg[9]  ( .D(n43597), .CP(clk), .Q(
        \filter_0/reg_i_7 [9]) );
  dff_sg \filter_0/reg_i_7_reg[10]  ( .D(n43527), .CP(clk), .Q(
        \filter_0/reg_i_7 [10]) );
  dff_sg \filter_0/reg_i_7_reg[11]  ( .D(n43594), .CP(clk), .Q(
        \filter_0/reg_i_7 [11]) );
  dff_sg \filter_0/reg_i_7_reg[12]  ( .D(n43618), .CP(clk), .Q(
        \filter_0/reg_i_7 [12]) );
  dff_sg \filter_0/reg_i_7_reg[13]  ( .D(n43621), .CP(clk), .Q(
        \filter_0/reg_i_7 [13]) );
  dff_sg \filter_0/reg_i_7_reg[14]  ( .D(n43526), .CP(clk), .Q(
        \filter_0/reg_i_7 [14]) );
  dff_sg \filter_0/reg_i_7_reg[15]  ( .D(n43525), .CP(clk), .Q(
        \filter_0/reg_i_7 [15]) );
  dff_sg \filter_0/reg_i_7_reg[16]  ( .D(n43648), .CP(clk), .Q(
        \filter_0/reg_i_7 [16]) );
  dff_sg \filter_0/reg_i_7_reg[17]  ( .D(n43651), .CP(clk), .Q(
        \filter_0/reg_i_7 [17]) );
  dff_sg \filter_0/reg_i_7_reg[18]  ( .D(n43662), .CP(clk), .Q(
        \filter_0/reg_i_7 [18]) );
  dff_sg \filter_0/reg_i_7_reg[19]  ( .D(n43654), .CP(clk), .Q(
        \filter_0/reg_i_7 [19]) );
  dff_sg \filter_0/reg_i_8_reg[0]  ( .D(n43630), .CP(clk), .Q(
        \filter_0/reg_i_8 [0]) );
  dff_sg \filter_0/reg_i_8_reg[1]  ( .D(n43633), .CP(clk), .Q(
        \filter_0/reg_i_8 [1]) );
  dff_sg \filter_0/reg_i_8_reg[2]  ( .D(n43636), .CP(clk), .Q(
        \filter_0/reg_i_8 [2]) );
  dff_sg \filter_0/reg_i_8_reg[3]  ( .D(n43639), .CP(clk), .Q(
        \filter_0/reg_i_8 [3]) );
  dff_sg \filter_0/reg_i_8_reg[4]  ( .D(n43657), .CP(clk), .Q(
        \filter_0/reg_i_8 [4]) );
  dff_sg \filter_0/reg_i_8_reg[5]  ( .D(n43645), .CP(clk), .Q(
        \filter_0/reg_i_8 [5]) );
  dff_sg \filter_0/reg_i_8_reg[6]  ( .D(n43714), .CP(clk), .Q(
        \filter_0/reg_i_8 [6]) );
  dff_sg \filter_0/reg_i_8_reg[7]  ( .D(n43717), .CP(clk), .Q(
        \filter_0/reg_i_8 [7]) );
  dff_sg \filter_0/reg_i_8_reg[8]  ( .D(n43711), .CP(clk), .Q(
        \filter_0/reg_i_8 [8]) );
  dff_sg \filter_0/reg_i_8_reg[9]  ( .D(n43490), .CP(clk), .Q(
        \filter_0/reg_i_8 [9]) );
  dff_sg \filter_0/reg_i_8_reg[10]  ( .D(n43705), .CP(clk), .Q(
        \filter_0/reg_i_8 [10]) );
  dff_sg \filter_0/reg_i_8_reg[11]  ( .D(n43708), .CP(clk), .Q(
        \filter_0/reg_i_8 [11]) );
  dff_sg \filter_0/reg_i_8_reg[12]  ( .D(n43997), .CP(clk), .Q(
        \filter_0/reg_i_8 [12]) );
  dff_sg \filter_0/reg_i_8_reg[13]  ( .D(n43998), .CP(clk), .Q(
        \filter_0/reg_i_8 [13]) );
  dff_sg \filter_0/reg_i_8_reg[14]  ( .D(n43488), .CP(clk), .Q(
        \filter_0/reg_i_8 [14]) );
  dff_sg \filter_0/reg_i_8_reg[15]  ( .D(n43489), .CP(clk), .Q(
        \filter_0/reg_i_8 [15]) );
  dff_sg \filter_0/reg_i_8_reg[16]  ( .D(n44003), .CP(clk), .Q(
        \filter_0/reg_i_8 [16]) );
  dff_sg \filter_0/reg_i_8_reg[17]  ( .D(n44004), .CP(clk), .Q(
        \filter_0/reg_i_8 [17]) );
  dff_sg \filter_0/reg_i_8_reg[18]  ( .D(n44000), .CP(clk), .Q(
        \filter_0/reg_i_8 [18]) );
  dff_sg \filter_0/reg_i_8_reg[19]  ( .D(n44001), .CP(clk), .Q(
        \filter_0/reg_i_8 [19]) );
  dff_sg \filter_0/reg_i_9_reg[0]  ( .D(n43987), .CP(clk), .Q(
        \filter_0/reg_i_9 [0]) );
  dff_sg \filter_0/reg_i_9_reg[1]  ( .D(n43988), .CP(clk), .Q(
        \filter_0/reg_i_9 [1]) );
  dff_sg \filter_0/reg_i_9_reg[2]  ( .D(n43984), .CP(clk), .Q(
        \filter_0/reg_i_9 [2]) );
  dff_sg \filter_0/reg_i_9_reg[3]  ( .D(n43985), .CP(clk), .Q(
        \filter_0/reg_i_9 [3]) );
  dff_sg \filter_0/reg_i_9_reg[4]  ( .D(n43993), .CP(clk), .Q(
        \filter_0/reg_i_9 [4]) );
  dff_sg \filter_0/reg_i_9_reg[5]  ( .D(n43994), .CP(clk), .Q(
        \filter_0/reg_i_9 [5]) );
  dff_sg \filter_0/reg_i_9_reg[6]  ( .D(n43990), .CP(clk), .Q(
        \filter_0/reg_i_9 [6]) );
  dff_sg \filter_0/reg_i_9_reg[7]  ( .D(n43991), .CP(clk), .Q(
        \filter_0/reg_i_9 [7]) );
  dff_sg \filter_0/reg_i_9_reg[8]  ( .D(n44019), .CP(clk), .Q(
        \filter_0/reg_i_9 [8]) );
  dff_sg \filter_0/reg_i_9_reg[9]  ( .D(n44020), .CP(clk), .Q(
        \filter_0/reg_i_9 [9]) );
  dff_sg \filter_0/reg_i_9_reg[10]  ( .D(n43478), .CP(clk), .Q(
        \filter_0/reg_i_9 [10]) );
  dff_sg \filter_0/reg_i_9_reg[11]  ( .D(n44017), .CP(clk), .Q(
        \filter_0/reg_i_9 [11]) );
  dff_sg \filter_0/reg_i_9_reg[12]  ( .D(n43476), .CP(clk), .Q(
        \filter_0/reg_i_9 [12]) );
  dff_sg \filter_0/reg_i_9_reg[13]  ( .D(n44024), .CP(clk), .Q(
        \filter_0/reg_i_9 [13]) );
  dff_sg \filter_0/reg_i_9_reg[14]  ( .D(n43481), .CP(clk), .Q(
        \filter_0/reg_i_9 [14]) );
  dff_sg \filter_0/reg_i_9_reg[15]  ( .D(n44022), .CP(clk), .Q(
        \filter_0/reg_i_9 [15]) );
  dff_sg \filter_0/reg_i_9_reg[16]  ( .D(n43479), .CP(clk), .Q(
        \filter_0/reg_i_9 [16]) );
  dff_sg \filter_0/reg_i_9_reg[17]  ( .D(n44009), .CP(clk), .Q(
        \filter_0/reg_i_9 [17]) );
  dff_sg \filter_0/reg_i_9_reg[18]  ( .D(n44006), .CP(clk), .Q(
        \filter_0/reg_i_9 [18]) );
  dff_sg \filter_0/reg_i_9_reg[19]  ( .D(n44007), .CP(clk), .Q(
        \filter_0/reg_i_9 [19]) );
  dff_sg \filter_0/reg_i_10_reg[0]  ( .D(n44014), .CP(clk), .Q(
        \filter_0/reg_i_10 [0]) );
  dff_sg \filter_0/reg_i_10_reg[1]  ( .D(n44015), .CP(clk), .Q(
        \filter_0/reg_i_10 [1]) );
  dff_sg \filter_0/reg_i_10_reg[2]  ( .D(n44011), .CP(clk), .Q(
        \filter_0/reg_i_10 [2]) );
  dff_sg \filter_0/reg_i_10_reg[3]  ( .D(n44012), .CP(clk), .Q(
        \filter_0/reg_i_10 [3]) );
  dff_sg \filter_0/reg_i_10_reg[4]  ( .D(n43957), .CP(clk), .Q(
        \filter_0/reg_i_10 [4]) );
  dff_sg \filter_0/reg_i_10_reg[5]  ( .D(n43958), .CP(clk), .Q(
        \filter_0/reg_i_10 [5]) );
  dff_sg \filter_0/reg_i_10_reg[6]  ( .D(n43954), .CP(clk), .Q(
        \filter_0/reg_i_10 [6]) );
  dff_sg \filter_0/reg_i_10_reg[7]  ( .D(n43955), .CP(clk), .Q(
        \filter_0/reg_i_10 [7]) );
  dff_sg \filter_0/reg_i_10_reg[8]  ( .D(n43962), .CP(clk), .Q(
        \filter_0/reg_i_10 [8]) );
  dff_sg \filter_0/reg_i_10_reg[9]  ( .D(n43963), .CP(clk), .Q(
        \filter_0/reg_i_10 [9]) );
  dff_sg \filter_0/reg_i_10_reg[10]  ( .D(n43960), .CP(clk), .Q(
        \filter_0/reg_i_10 [10]) );
  dff_sg \filter_0/reg_i_10_reg[11]  ( .D(n43472), .CP(clk), .Q(
        \filter_0/reg_i_10 [11]) );
  dff_sg \filter_0/reg_i_10_reg[12]  ( .D(n43946), .CP(clk), .Q(
        \filter_0/reg_i_10 [12]) );
  dff_sg \filter_0/reg_i_10_reg[13]  ( .D(n43947), .CP(clk), .Q(
        \filter_0/reg_i_10 [13]) );
  dff_sg \filter_0/reg_i_10_reg[14]  ( .D(n43943), .CP(clk), .Q(
        \filter_0/reg_i_10 [14]) );
  dff_sg \filter_0/reg_i_10_reg[15]  ( .D(n43944), .CP(clk), .Q(
        \filter_0/reg_i_10 [15]) );
  dff_sg \filter_0/reg_i_10_reg[16]  ( .D(n43951), .CP(clk), .Q(
        \filter_0/reg_i_10 [16]) );
  dff_sg \filter_0/reg_i_10_reg[17]  ( .D(n43952), .CP(clk), .Q(
        \filter_0/reg_i_10 [17]) );
  dff_sg \filter_0/reg_i_10_reg[18]  ( .D(n43480), .CP(clk), .Q(
        \filter_0/reg_i_10 [18]) );
  dff_sg \filter_0/reg_i_10_reg[19]  ( .D(n43949), .CP(clk), .Q(
        \filter_0/reg_i_10 [19]) );
  dff_sg \filter_0/reg_i_11_reg[0]  ( .D(n43976), .CP(clk), .Q(
        \filter_0/reg_i_11 [0]) );
  dff_sg \filter_0/reg_i_11_reg[1]  ( .D(n43977), .CP(clk), .Q(
        \filter_0/reg_i_11 [1]) );
  dff_sg \filter_0/reg_i_11_reg[2]  ( .D(n43483), .CP(clk), .Q(
        \filter_0/reg_i_11 [2]) );
  dff_sg \filter_0/reg_i_11_reg[3]  ( .D(n43974), .CP(clk), .Q(
        \filter_0/reg_i_11 [3]) );
  dff_sg \filter_0/reg_i_11_reg[4]  ( .D(n43981), .CP(clk), .Q(
        \filter_0/reg_i_11 [4]) );
  dff_sg \filter_0/reg_i_11_reg[5]  ( .D(n43982), .CP(clk), .Q(
        \filter_0/reg_i_11 [5]) );
  dff_sg \filter_0/reg_i_11_reg[6]  ( .D(n43482), .CP(clk), .Q(
        \filter_0/reg_i_11 [6]) );
  dff_sg \filter_0/reg_i_11_reg[7]  ( .D(n43979), .CP(clk), .Q(
        \filter_0/reg_i_11 [7]) );
  dff_sg \filter_0/reg_i_11_reg[8]  ( .D(n43484), .CP(clk), .Q(
        \filter_0/reg_i_11 [8]) );
  dff_sg \filter_0/reg_i_11_reg[9]  ( .D(n43968), .CP(clk), .Q(
        \filter_0/reg_i_11 [9]) );
  dff_sg \filter_0/reg_i_11_reg[10]  ( .D(n43965), .CP(clk), .Q(
        \filter_0/reg_i_11 [10]) );
  dff_sg \filter_0/reg_i_11_reg[11]  ( .D(n43966), .CP(clk), .Q(
        \filter_0/reg_i_11 [11]) );
  dff_sg \filter_0/reg_i_11_reg[12]  ( .D(n43972), .CP(clk), .Q(
        \filter_0/reg_i_11 [12]) );
  dff_sg \filter_0/reg_i_11_reg[13]  ( .D(n43470), .CP(clk), .Q(
        \filter_0/reg_i_11 [13]) );
  dff_sg \filter_0/reg_i_11_reg[14]  ( .D(n43477), .CP(clk), .Q(
        \filter_0/reg_i_11 [14]) );
  dff_sg \filter_0/reg_i_11_reg[15]  ( .D(n43970), .CP(clk), .Q(
        \filter_0/reg_i_11 [15]) );
  dff_sg \filter_0/reg_i_11_reg[16]  ( .D(n44078), .CP(clk), .Q(
        \filter_0/reg_i_11 [16]) );
  dff_sg \filter_0/reg_i_11_reg[17]  ( .D(n44075), .CP(clk), .Q(
        \filter_0/reg_i_11 [17]) );
  dff_sg \filter_0/reg_i_11_reg[18]  ( .D(n44079), .CP(clk), .Q(
        \filter_0/reg_i_11 [18]) );
  dff_sg \filter_0/reg_i_11_reg[19]  ( .D(n44080), .CP(clk), .Q(
        \filter_0/reg_i_11 [19]) );
  dff_sg \filter_0/reg_i_12_reg[0]  ( .D(n44082), .CP(clk), .Q(
        \filter_0/reg_i_12 [0]) );
  dff_sg \filter_0/reg_i_12_reg[1]  ( .D(n44083), .CP(clk), .Q(
        \filter_0/reg_i_12 [1]) );
  dff_sg \filter_0/reg_i_12_reg[2]  ( .D(n44081), .CP(clk), .Q(
        \filter_0/reg_i_12 [2]) );
  dff_sg \filter_0/reg_i_12_reg[3]  ( .D(n44072), .CP(clk), .Q(
        \filter_0/reg_i_12 [3]) );
  dff_sg \filter_0/reg_i_12_reg[4]  ( .D(n43534), .CP(clk), .Q(
        \filter_0/reg_i_12 [4]) );
  dff_sg \filter_0/reg_i_12_reg[5]  ( .D(n43535), .CP(clk), .Q(
        \filter_0/reg_i_12 [5]) );
  dff_sg \filter_0/reg_i_12_reg[6]  ( .D(n43536), .CP(clk), .Q(
        \filter_0/reg_i_12 [6]) );
  dff_sg \filter_0/reg_i_12_reg[7]  ( .D(n44066), .CP(clk), .Q(
        \filter_0/reg_i_12 [7]) );
  dff_sg \filter_0/reg_i_12_reg[8]  ( .D(n44076), .CP(clk), .Q(
        \filter_0/reg_i_12 [8]) );
  dff_sg \filter_0/reg_i_12_reg[9]  ( .D(n44077), .CP(clk), .Q(
        \filter_0/reg_i_12 [9]) );
  dff_sg \filter_0/reg_i_12_reg[10]  ( .D(n44073), .CP(clk), .Q(
        \filter_0/reg_i_12 [10]) );
  dff_sg \filter_0/reg_i_12_reg[11]  ( .D(n44069), .CP(clk), .Q(
        \filter_0/reg_i_12 [11]) );
  dff_sg \filter_0/reg_i_12_reg[12]  ( .D(n44094), .CP(clk), .Q(
        \filter_0/reg_i_12 [12]) );
  dff_sg \filter_0/reg_i_12_reg[13]  ( .D(n44095), .CP(clk), .Q(
        \filter_0/reg_i_12 [13]) );
  dff_sg \filter_0/reg_i_12_reg[14]  ( .D(n44092), .CP(clk), .Q(
        \filter_0/reg_i_12 [14]) );
  dff_sg \filter_0/reg_i_12_reg[15]  ( .D(n44093), .CP(clk), .Q(
        \filter_0/reg_i_12 [15]) );
  dff_sg \filter_0/reg_i_12_reg[16]  ( .D(n44099), .CP(clk), .Q(
        \filter_0/reg_i_12 [16]) );
  dff_sg \filter_0/reg_i_12_reg[17]  ( .D(n44091), .CP(clk), .Q(
        \filter_0/reg_i_12 [17]) );
  dff_sg \filter_0/reg_i_12_reg[18]  ( .D(n44100), .CP(clk), .Q(
        \filter_0/reg_i_12 [18]) );
  dff_sg \filter_0/reg_i_12_reg[19]  ( .D(n44101), .CP(clk), .Q(
        \filter_0/reg_i_12 [19]) );
  dff_sg \filter_0/reg_i_13_reg[0]  ( .D(n44089), .CP(clk), .Q(
        \filter_0/reg_i_13 [0]) );
  dff_sg \filter_0/reg_i_13_reg[1]  ( .D(n44090), .CP(clk), .Q(
        \filter_0/reg_i_13 [1]) );
  dff_sg \filter_0/reg_i_13_reg[2]  ( .D(n44086), .CP(clk), .Q(
        \filter_0/reg_i_13 [2]) );
  dff_sg \filter_0/reg_i_13_reg[3]  ( .D(n44087), .CP(clk), .Q(
        \filter_0/reg_i_13 [3]) );
  dff_sg \filter_0/reg_i_13_reg[4]  ( .D(n44088), .CP(clk), .Q(
        \filter_0/reg_i_13 [4]) );
  dff_sg \filter_0/reg_i_13_reg[5]  ( .D(n44074), .CP(clk), .Q(
        \filter_0/reg_i_13 [5]) );
  dff_sg \filter_0/reg_i_13_reg[6]  ( .D(n44084), .CP(clk), .Q(
        \filter_0/reg_i_13 [6]) );
  dff_sg \filter_0/reg_i_13_reg[7]  ( .D(n44085), .CP(clk), .Q(
        \filter_0/reg_i_13 [7]) );
  dff_sg \filter_0/reg_i_13_reg[8]  ( .D(n44041), .CP(clk), .Q(
        \filter_0/reg_i_13 [8]) );
  dff_sg \filter_0/reg_i_13_reg[9]  ( .D(n44042), .CP(clk), .Q(
        \filter_0/reg_i_13 [9]) );
  dff_sg \filter_0/reg_i_13_reg[10]  ( .D(n44038), .CP(clk), .Q(
        \filter_0/reg_i_13 [10]) );
  dff_sg \filter_0/reg_i_13_reg[11]  ( .D(n44039), .CP(clk), .Q(
        \filter_0/reg_i_13 [11]) );
  dff_sg \filter_0/reg_i_13_reg[12]  ( .D(n44046), .CP(clk), .Q(
        \filter_0/reg_i_13 [12]) );
  dff_sg \filter_0/reg_i_13_reg[13]  ( .D(n44047), .CP(clk), .Q(
        \filter_0/reg_i_13 [13]) );
  dff_sg \filter_0/reg_i_13_reg[14]  ( .D(n44043), .CP(clk), .Q(
        \filter_0/reg_i_13 [14]) );
  dff_sg \filter_0/reg_i_13_reg[15]  ( .D(n44044), .CP(clk), .Q(
        \filter_0/reg_i_13 [15]) );
  dff_sg \filter_0/reg_i_13_reg[16]  ( .D(n44029), .CP(clk), .Q(
        \filter_0/reg_i_13 [16]) );
  dff_sg \filter_0/reg_i_13_reg[17]  ( .D(n44030), .CP(clk), .Q(
        \filter_0/reg_i_13 [17]) );
  dff_sg \filter_0/reg_i_13_reg[18]  ( .D(n44026), .CP(clk), .Q(
        \filter_0/reg_i_13 [18]) );
  dff_sg \filter_0/reg_i_13_reg[19]  ( .D(n44027), .CP(clk), .Q(
        \filter_0/reg_i_13 [19]) );
  dff_sg \filter_0/reg_i_14_reg[0]  ( .D(n44035), .CP(clk), .Q(
        \filter_0/reg_i_14 [0]) );
  dff_sg \filter_0/reg_i_14_reg[1]  ( .D(n44036), .CP(clk), .Q(
        \filter_0/reg_i_14 [1]) );
  dff_sg \filter_0/reg_i_14_reg[2]  ( .D(n44032), .CP(clk), .Q(
        \filter_0/reg_i_14 [2]) );
  dff_sg \filter_0/reg_i_14_reg[3]  ( .D(n44033), .CP(clk), .Q(
        \filter_0/reg_i_14 [3]) );
  dff_sg \filter_0/reg_i_14_reg[4]  ( .D(n44064), .CP(clk), .Q(
        \filter_0/reg_i_14 [4]) );
  dff_sg \filter_0/reg_i_14_reg[5]  ( .D(n44065), .CP(clk), .Q(
        \filter_0/reg_i_14 [5]) );
  dff_sg \filter_0/reg_i_14_reg[6]  ( .D(n44061), .CP(clk), .Q(
        \filter_0/reg_i_14 [6]) );
  dff_sg \filter_0/reg_i_14_reg[7]  ( .D(n44062), .CP(clk), .Q(
        \filter_0/reg_i_14 [7]) );
  dff_sg \filter_0/reg_i_14_reg[8]  ( .D(n44070), .CP(clk), .Q(
        \filter_0/reg_i_14 [8]) );
  dff_sg \filter_0/reg_i_14_reg[9]  ( .D(n44071), .CP(clk), .Q(
        \filter_0/reg_i_14 [9]) );
  dff_sg \filter_0/reg_i_14_reg[10]  ( .D(n44067), .CP(clk), .Q(
        \filter_0/reg_i_14 [10]) );
  dff_sg \filter_0/reg_i_14_reg[11]  ( .D(n44068), .CP(clk), .Q(
        \filter_0/reg_i_14 [11]) );
  dff_sg \filter_0/reg_i_14_reg[12]  ( .D(n44052), .CP(clk), .Q(
        \filter_0/reg_i_14 [12]) );
  dff_sg \filter_0/reg_i_14_reg[13]  ( .D(n44053), .CP(clk), .Q(
        \filter_0/reg_i_14 [13]) );
  dff_sg \filter_0/reg_i_14_reg[14]  ( .D(n44049), .CP(clk), .Q(
        \filter_0/reg_i_14 [14]) );
  dff_sg \filter_0/reg_i_14_reg[15]  ( .D(n44050), .CP(clk), .Q(
        \filter_0/reg_i_14 [15]) );
  dff_sg \filter_0/reg_i_14_reg[16]  ( .D(n44058), .CP(clk), .Q(
        \filter_0/reg_i_14 [16]) );
  dff_sg \filter_0/reg_i_14_reg[17]  ( .D(n44059), .CP(clk), .Q(
        \filter_0/reg_i_14 [17]) );
  dff_sg \filter_0/reg_i_14_reg[18]  ( .D(n44055), .CP(clk), .Q(
        \filter_0/reg_i_14 [18]) );
  dff_sg \filter_0/reg_i_14_reg[19]  ( .D(n44056), .CP(clk), .Q(
        \filter_0/reg_i_14 [19]) );
  dff_sg \filter_0/reg_i_15_reg[0]  ( .D(n43817), .CP(clk), .Q(
        \filter_0/reg_i_15 [0]) );
  dff_sg \filter_0/reg_i_15_reg[1]  ( .D(n43818), .CP(clk), .Q(
        \filter_0/reg_i_15 [1]) );
  dff_sg \filter_0/reg_i_15_reg[2]  ( .D(n43814), .CP(clk), .Q(
        \filter_0/reg_i_15 [2]) );
  dff_sg \filter_0/reg_i_15_reg[3]  ( .D(n43815), .CP(clk), .Q(
        \filter_0/reg_i_15 [3]) );
  dff_sg \filter_0/reg_i_15_reg[4]  ( .D(n43823), .CP(clk), .Q(
        \filter_0/reg_i_15 [4]) );
  dff_sg \filter_0/reg_i_15_reg[5]  ( .D(n43824), .CP(clk), .Q(
        \filter_0/reg_i_15 [5]) );
  dff_sg \filter_0/reg_i_15_reg[6]  ( .D(n43820), .CP(clk), .Q(
        \filter_0/reg_i_15 [6]) );
  dff_sg \filter_0/reg_i_15_reg[7]  ( .D(n43821), .CP(clk), .Q(
        \filter_0/reg_i_15 [7]) );
  dff_sg \filter_0/reg_i_15_reg[8]  ( .D(n43805), .CP(clk), .Q(
        \filter_0/reg_i_15 [8]) );
  dff_sg \filter_0/reg_i_15_reg[9]  ( .D(n43806), .CP(clk), .Q(
        \filter_0/reg_i_15 [9]) );
  dff_sg \filter_0/reg_i_15_reg[10]  ( .D(n43802), .CP(clk), .Q(
        \filter_0/reg_i_15 [10]) );
  dff_sg \filter_0/reg_i_15_reg[11]  ( .D(n43803), .CP(clk), .Q(
        \filter_0/reg_i_15 [11]) );
  dff_sg \filter_0/reg_i_15_reg[12]  ( .D(n43811), .CP(clk), .Q(
        \filter_0/reg_i_15 [12]) );
  dff_sg \filter_0/reg_i_15_reg[13]  ( .D(n43812), .CP(clk), .Q(
        \filter_0/reg_i_15 [13]) );
  dff_sg \filter_0/reg_i_15_reg[14]  ( .D(n43808), .CP(clk), .Q(
        \filter_0/reg_i_15 [14]) );
  dff_sg \filter_0/reg_i_15_reg[15]  ( .D(n43809), .CP(clk), .Q(
        \filter_0/reg_i_15 [15]) );
  dff_sg \filter_0/reg_i_15_reg[16]  ( .D(n43475), .CP(clk), .Q(
        \filter_0/reg_i_15 [16]) );
  dff_sg \filter_0/reg_i_15_reg[17]  ( .D(n43840), .CP(clk), .Q(
        \filter_0/reg_i_15 [17]) );
  dff_sg \filter_0/reg_i_15_reg[18]  ( .D(n43473), .CP(clk), .Q(
        \filter_0/reg_i_15 [18]) );
  dff_sg \filter_0/reg_i_15_reg[19]  ( .D(n43838), .CP(clk), .Q(
        \filter_0/reg_i_15 [19]) );
  dff_sg \filter_0/reg_w_0_reg[0]  ( .D(n43845), .CP(clk), .Q(
        \filter_0/reg_w_0 [0]) );
  dff_sg \filter_0/reg_w_0_reg[1]  ( .D(n43846), .CP(clk), .Q(
        \filter_0/reg_w_0 [1]) );
  dff_sg \filter_0/reg_w_0_reg[2]  ( .D(n43842), .CP(clk), .Q(
        \filter_0/reg_w_0 [2]) );
  dff_sg \filter_0/reg_w_0_reg[3]  ( .D(n43843), .CP(clk), .Q(
        \filter_0/reg_w_0 [3]) );
  dff_sg \filter_0/reg_w_0_reg[4]  ( .D(n43829), .CP(clk), .Q(
        \filter_0/reg_w_0 [4]) );
  dff_sg \filter_0/reg_w_0_reg[5]  ( .D(n43830), .CP(clk), .Q(
        \filter_0/reg_w_0 [5]) );
  dff_sg \filter_0/reg_w_0_reg[6]  ( .D(n43826), .CP(clk), .Q(
        \filter_0/reg_w_0 [6]) );
  dff_sg \filter_0/reg_w_0_reg[7]  ( .D(n43827), .CP(clk), .Q(
        \filter_0/reg_w_0 [7]) );
  dff_sg \filter_0/reg_w_0_reg[8]  ( .D(n43835), .CP(clk), .Q(
        \filter_0/reg_w_0 [8]) );
  dff_sg \filter_0/reg_w_0_reg[9]  ( .D(n43836), .CP(clk), .Q(
        \filter_0/reg_w_0 [9]) );
  dff_sg \filter_0/reg_w_0_reg[10]  ( .D(n43832), .CP(clk), .Q(
        \filter_0/reg_w_0 [10]) );
  dff_sg \filter_0/reg_w_0_reg[11]  ( .D(n43833), .CP(clk), .Q(
        \filter_0/reg_w_0 [11]) );
  dff_sg \filter_0/reg_w_0_reg[12]  ( .D(n43769), .CP(clk), .Q(
        \filter_0/reg_w_0 [12]) );
  dff_sg \filter_0/reg_w_0_reg[13]  ( .D(n43770), .CP(clk), .Q(
        \filter_0/reg_w_0 [13]) );
  dff_sg \filter_0/reg_w_0_reg[14]  ( .D(n43766), .CP(clk), .Q(
        \filter_0/reg_w_0 [14]) );
  dff_sg \filter_0/reg_w_0_reg[15]  ( .D(n43767), .CP(clk), .Q(
        \filter_0/reg_w_0 [15]) );
  dff_sg \filter_0/reg_w_0_reg[16]  ( .D(n43775), .CP(clk), .Q(
        \filter_0/reg_w_0 [16]) );
  dff_sg \filter_0/reg_w_0_reg[17]  ( .D(n43776), .CP(clk), .Q(
        \filter_0/reg_w_0 [17]) );
  dff_sg \filter_0/reg_w_0_reg[18]  ( .D(n43772), .CP(clk), .Q(
        \filter_0/reg_w_0 [18]) );
  dff_sg \filter_0/reg_w_0_reg[19]  ( .D(n43773), .CP(clk), .Q(
        \filter_0/reg_w_0 [19]) );
  dff_sg \filter_0/reg_w_1_reg[0]  ( .D(n43757), .CP(clk), .Q(
        \filter_0/reg_w_1 [0]) );
  dff_sg \filter_0/reg_w_1_reg[1]  ( .D(n43758), .CP(clk), .Q(
        \filter_0/reg_w_1 [1]) );
  dff_sg \filter_0/reg_w_1_reg[2]  ( .D(n43754), .CP(clk), .Q(
        \filter_0/reg_w_1 [2]) );
  dff_sg \filter_0/reg_w_1_reg[3]  ( .D(n43755), .CP(clk), .Q(
        \filter_0/reg_w_1 [3]) );
  dff_sg \filter_0/reg_w_1_reg[4]  ( .D(n43763), .CP(clk), .Q(
        \filter_0/reg_w_1 [4]) );
  dff_sg \filter_0/reg_w_1_reg[5]  ( .D(n43764), .CP(clk), .Q(
        \filter_0/reg_w_1 [5]) );
  dff_sg \filter_0/reg_w_1_reg[6]  ( .D(n43760), .CP(clk), .Q(
        \filter_0/reg_w_1 [6]) );
  dff_sg \filter_0/reg_w_1_reg[7]  ( .D(n43761), .CP(clk), .Q(
        \filter_0/reg_w_1 [7]) );
  dff_sg \filter_0/reg_w_1_reg[8]  ( .D(n43793), .CP(clk), .Q(
        \filter_0/reg_w_1 [8]) );
  dff_sg \filter_0/reg_w_1_reg[9]  ( .D(n43794), .CP(clk), .Q(
        \filter_0/reg_w_1 [9]) );
  dff_sg \filter_0/reg_w_1_reg[10]  ( .D(n43790), .CP(clk), .Q(
        \filter_0/reg_w_1 [10]) );
  dff_sg \filter_0/reg_w_1_reg[11]  ( .D(n43791), .CP(clk), .Q(
        \filter_0/reg_w_1 [11]) );
  dff_sg \filter_0/reg_w_1_reg[12]  ( .D(n43799), .CP(clk), .Q(
        \filter_0/reg_w_1 [12]) );
  dff_sg \filter_0/reg_w_1_reg[13]  ( .D(n43800), .CP(clk), .Q(
        \filter_0/reg_w_1 [13]) );
  dff_sg \filter_0/reg_w_1_reg[14]  ( .D(n43796), .CP(clk), .Q(
        \filter_0/reg_w_1 [14]) );
  dff_sg \filter_0/reg_w_1_reg[15]  ( .D(n43797), .CP(clk), .Q(
        \filter_0/reg_w_1 [15]) );
  dff_sg \filter_0/reg_w_1_reg[16]  ( .D(n43781), .CP(clk), .Q(
        \filter_0/reg_w_1 [16]) );
  dff_sg \filter_0/reg_w_1_reg[17]  ( .D(n43782), .CP(clk), .Q(
        \filter_0/reg_w_1 [17]) );
  dff_sg \filter_0/reg_w_1_reg[18]  ( .D(n43778), .CP(clk), .Q(
        \filter_0/reg_w_1 [18]) );
  dff_sg \filter_0/reg_w_1_reg[19]  ( .D(n43779), .CP(clk), .Q(
        \filter_0/reg_w_1 [19]) );
  dff_sg \filter_0/reg_w_2_reg[0]  ( .D(n43787), .CP(clk), .Q(
        \filter_0/reg_w_2 [0]) );
  dff_sg \filter_0/reg_w_2_reg[1]  ( .D(n43788), .CP(clk), .Q(
        \filter_0/reg_w_2 [1]) );
  dff_sg \filter_0/reg_w_2_reg[2]  ( .D(n43784), .CP(clk), .Q(
        \filter_0/reg_w_2 [2]) );
  dff_sg \filter_0/reg_w_2_reg[3]  ( .D(n43785), .CP(clk), .Q(
        \filter_0/reg_w_2 [3]) );
  dff_sg \filter_0/reg_w_2_reg[4]  ( .D(n43910), .CP(clk), .Q(
        \filter_0/reg_w_2 [4]) );
  dff_sg \filter_0/reg_w_2_reg[5]  ( .D(n43911), .CP(clk), .Q(
        \filter_0/reg_w_2 [5]) );
  dff_sg \filter_0/reg_w_2_reg[6]  ( .D(n43907), .CP(clk), .Q(
        \filter_0/reg_w_2 [6]) );
  dff_sg \filter_0/reg_w_2_reg[7]  ( .D(n43908), .CP(clk), .Q(
        \filter_0/reg_w_2 [7]) );
  dff_sg \filter_0/reg_w_2_reg[8]  ( .D(n43916), .CP(clk), .Q(
        \filter_0/reg_w_2 [8]) );
  dff_sg \filter_0/reg_w_2_reg[9]  ( .D(n43917), .CP(clk), .Q(
        \filter_0/reg_w_2 [9]) );
  dff_sg \filter_0/reg_w_2_reg[10]  ( .D(n43913), .CP(clk), .Q(
        \filter_0/reg_w_2 [10]) );
  dff_sg \filter_0/reg_w_2_reg[11]  ( .D(n43914), .CP(clk), .Q(
        \filter_0/reg_w_2 [11]) );
  dff_sg \filter_0/reg_w_2_reg[12]  ( .D(n43898), .CP(clk), .Q(
        \filter_0/reg_w_2 [12]) );
  dff_sg \filter_0/reg_w_2_reg[13]  ( .D(n43899), .CP(clk), .Q(
        \filter_0/reg_w_2 [13]) );
  dff_sg \filter_0/reg_w_2_reg[14]  ( .D(n43895), .CP(clk), .Q(
        \filter_0/reg_w_2 [14]) );
  dff_sg \filter_0/reg_w_2_reg[15]  ( .D(n43896), .CP(clk), .Q(
        \filter_0/reg_w_2 [15]) );
  dff_sg \filter_0/reg_w_2_reg[16]  ( .D(n43904), .CP(clk), .Q(
        \filter_0/reg_w_2 [16]) );
  dff_sg \filter_0/reg_w_2_reg[17]  ( .D(n43905), .CP(clk), .Q(
        \filter_0/reg_w_2 [17]) );
  dff_sg \filter_0/reg_w_2_reg[18]  ( .D(n43901), .CP(clk), .Q(
        \filter_0/reg_w_2 [18]) );
  dff_sg \filter_0/reg_w_2_reg[19]  ( .D(n43902), .CP(clk), .Q(
        \filter_0/reg_w_2 [19]) );
  dff_sg \filter_0/reg_w_3_reg[0]  ( .D(n43934), .CP(clk), .Q(
        \filter_0/reg_w_3 [0]) );
  dff_sg \filter_0/reg_w_3_reg[1]  ( .D(n43935), .CP(clk), .Q(
        \filter_0/reg_w_3 [1]) );
  dff_sg \filter_0/reg_w_3_reg[2]  ( .D(n43931), .CP(clk), .Q(
        \filter_0/reg_w_3 [2]) );
  dff_sg \filter_0/reg_w_3_reg[3]  ( .D(n43932), .CP(clk), .Q(
        \filter_0/reg_w_3 [3]) );
  dff_sg \filter_0/reg_w_3_reg[4]  ( .D(n43940), .CP(clk), .Q(
        \filter_0/reg_w_3 [4]) );
  dff_sg \filter_0/reg_w_3_reg[5]  ( .D(n43941), .CP(clk), .Q(
        \filter_0/reg_w_3 [5]) );
  dff_sg \filter_0/reg_w_3_reg[6]  ( .D(n43937), .CP(clk), .Q(
        \filter_0/reg_w_3 [6]) );
  dff_sg \filter_0/reg_w_3_reg[7]  ( .D(n43938), .CP(clk), .Q(
        \filter_0/reg_w_3 [7]) );
  dff_sg \filter_0/reg_w_3_reg[8]  ( .D(n43922), .CP(clk), .Q(
        \filter_0/reg_w_3 [8]) );
  dff_sg \filter_0/reg_w_3_reg[9]  ( .D(n43923), .CP(clk), .Q(
        \filter_0/reg_w_3 [9]) );
  dff_sg \filter_0/reg_w_3_reg[10]  ( .D(n43919), .CP(clk), .Q(
        \filter_0/reg_w_3 [10]) );
  dff_sg \filter_0/reg_w_3_reg[11]  ( .D(n43920), .CP(clk), .Q(
        \filter_0/reg_w_3 [11]) );
  dff_sg \filter_0/reg_w_3_reg[12]  ( .D(n43928), .CP(clk), .Q(
        \filter_0/reg_w_3 [12]) );
  dff_sg \filter_0/reg_w_3_reg[13]  ( .D(n43929), .CP(clk), .Q(
        \filter_0/reg_w_3 [13]) );
  dff_sg \filter_0/reg_w_3_reg[14]  ( .D(n43925), .CP(clk), .Q(
        \filter_0/reg_w_3 [14]) );
  dff_sg \filter_0/reg_w_3_reg[15]  ( .D(n43926), .CP(clk), .Q(
        \filter_0/reg_w_3 [15]) );
  dff_sg \filter_0/reg_w_3_reg[16]  ( .D(n43863), .CP(clk), .Q(
        \filter_0/reg_w_3 [16]) );
  dff_sg \filter_0/reg_w_3_reg[17]  ( .D(n43864), .CP(clk), .Q(
        \filter_0/reg_w_3 [17]) );
  dff_sg \filter_0/reg_w_3_reg[18]  ( .D(n43860), .CP(clk), .Q(
        \filter_0/reg_w_3 [18]) );
  dff_sg \filter_0/reg_w_3_reg[19]  ( .D(n43861), .CP(clk), .Q(
        \filter_0/reg_w_3 [19]) );
  dff_sg \filter_0/reg_w_4_reg[0]  ( .D(n43869), .CP(clk), .Q(
        \filter_0/reg_w_4 [0]) );
  dff_sg \filter_0/reg_w_4_reg[1]  ( .D(n43870), .CP(clk), .Q(
        \filter_0/reg_w_4 [1]) );
  dff_sg \filter_0/reg_w_4_reg[2]  ( .D(n43866), .CP(clk), .Q(
        \filter_0/reg_w_4 [2]) );
  dff_sg \filter_0/reg_w_4_reg[3]  ( .D(n43867), .CP(clk), .Q(
        \filter_0/reg_w_4 [3]) );
  dff_sg \filter_0/reg_w_4_reg[4]  ( .D(n43851), .CP(clk), .Q(
        \filter_0/reg_w_4 [4]) );
  dff_sg \filter_0/reg_w_4_reg[5]  ( .D(n43852), .CP(clk), .Q(
        \filter_0/reg_w_4 [5]) );
  dff_sg \filter_0/reg_w_4_reg[6]  ( .D(n43848), .CP(clk), .Q(
        \filter_0/reg_w_4 [6]) );
  dff_sg \filter_0/reg_w_4_reg[7]  ( .D(n43849), .CP(clk), .Q(
        \filter_0/reg_w_4 [7]) );
  dff_sg \filter_0/reg_w_4_reg[8]  ( .D(n43857), .CP(clk), .Q(
        \filter_0/reg_w_4 [8]) );
  dff_sg \filter_0/reg_w_4_reg[9]  ( .D(n43858), .CP(clk), .Q(
        \filter_0/reg_w_4 [9]) );
  dff_sg \filter_0/reg_w_4_reg[10]  ( .D(n43854), .CP(clk), .Q(
        \filter_0/reg_w_4 [10]) );
  dff_sg \filter_0/reg_w_4_reg[11]  ( .D(n43855), .CP(clk), .Q(
        \filter_0/reg_w_4 [11]) );
  dff_sg \filter_0/reg_w_4_reg[12]  ( .D(n43886), .CP(clk), .Q(
        \filter_0/reg_w_4 [12]) );
  dff_sg \filter_0/reg_w_4_reg[13]  ( .D(n43887), .CP(clk), .Q(
        \filter_0/reg_w_4 [13]) );
  dff_sg \filter_0/reg_w_4_reg[14]  ( .D(n43883), .CP(clk), .Q(
        \filter_0/reg_w_4 [14]) );
  dff_sg \filter_0/reg_w_4_reg[15]  ( .D(n43884), .CP(clk), .Q(
        \filter_0/reg_w_4 [15]) );
  dff_sg \filter_0/reg_w_4_reg[16]  ( .D(n43892), .CP(clk), .Q(
        \filter_0/reg_w_4 [16]) );
  dff_sg \filter_0/reg_w_4_reg[17]  ( .D(n43893), .CP(clk), .Q(
        \filter_0/reg_w_4 [17]) );
  dff_sg \filter_0/reg_w_4_reg[18]  ( .D(n43889), .CP(clk), .Q(
        \filter_0/reg_w_4 [18]) );
  dff_sg \filter_0/reg_w_4_reg[19]  ( .D(n43890), .CP(clk), .Q(
        \filter_0/reg_w_4 [19]) );
  dff_sg \filter_0/reg_w_5_reg[0]  ( .D(n43875), .CP(clk), .Q(
        \filter_0/reg_w_5 [0]) );
  dff_sg \filter_0/reg_w_5_reg[1]  ( .D(n43876), .CP(clk), .Q(
        \filter_0/reg_w_5 [1]) );
  dff_sg \filter_0/reg_w_5_reg[2]  ( .D(n43872), .CP(clk), .Q(
        \filter_0/reg_w_5 [2]) );
  dff_sg \filter_0/reg_w_5_reg[3]  ( .D(n43873), .CP(clk), .Q(
        \filter_0/reg_w_5 [3]) );
  dff_sg \filter_0/reg_w_5_reg[4]  ( .D(n43880), .CP(clk), .Q(
        \filter_0/reg_w_5 [4]) );
  dff_sg \filter_0/reg_w_5_reg[5]  ( .D(n43881), .CP(clk), .Q(
        \filter_0/reg_w_5 [5]) );
  dff_sg \filter_0/reg_w_5_reg[6]  ( .D(n43471), .CP(clk), .Q(
        \filter_0/reg_w_5 [6]) );
  dff_sg \filter_0/reg_w_5_reg[7]  ( .D(n43878), .CP(clk), .Q(
        \filter_0/reg_w_5 [7]) );
  dff_sg \filter_0/reg_w_5_reg[8]  ( .D(n43580), .CP(clk), .Q(
        \filter_0/reg_w_5 [8]) );
  dff_sg \filter_0/reg_w_5_reg[9]  ( .D(n43581), .CP(clk), .Q(
        \filter_0/reg_w_5 [9]) );
  dff_sg \filter_0/reg_w_5_reg[10]  ( .D(n43577), .CP(clk), .Q(
        \filter_0/reg_w_5 [10]) );
  dff_sg \filter_0/reg_w_5_reg[11]  ( .D(n43578), .CP(clk), .Q(
        \filter_0/reg_w_5 [11]) );
  dff_sg \filter_0/reg_w_5_reg[12]  ( .D(n43586), .CP(clk), .Q(
        \filter_0/reg_w_5 [12]) );
  dff_sg \filter_0/reg_w_5_reg[13]  ( .D(n43587), .CP(clk), .Q(
        \filter_0/reg_w_5 [13]) );
  dff_sg \filter_0/reg_w_5_reg[14]  ( .D(n43583), .CP(clk), .Q(
        \filter_0/reg_w_5 [14]) );
  dff_sg \filter_0/reg_w_5_reg[15]  ( .D(n43584), .CP(clk), .Q(
        \filter_0/reg_w_5 [15]) );
  dff_sg \filter_0/reg_w_5_reg[16]  ( .D(n43568), .CP(clk), .Q(
        \filter_0/reg_w_5 [16]) );
  dff_sg \filter_0/reg_w_5_reg[17]  ( .D(n43569), .CP(clk), .Q(
        \filter_0/reg_w_5 [17]) );
  dff_sg \filter_0/reg_w_5_reg[18]  ( .D(n43565), .CP(clk), .Q(
        \filter_0/reg_w_5 [18]) );
  dff_sg \filter_0/reg_w_5_reg[19]  ( .D(n43566), .CP(clk), .Q(
        \filter_0/reg_w_5 [19]) );
  dff_sg \filter_0/reg_w_6_reg[0]  ( .D(n43574), .CP(clk), .Q(
        \filter_0/reg_w_6 [0]) );
  dff_sg \filter_0/reg_w_6_reg[1]  ( .D(n43575), .CP(clk), .Q(
        \filter_0/reg_w_6 [1]) );
  dff_sg \filter_0/reg_w_6_reg[2]  ( .D(n43571), .CP(clk), .Q(
        \filter_0/reg_w_6 [2]) );
  dff_sg \filter_0/reg_w_6_reg[3]  ( .D(n43572), .CP(clk), .Q(
        \filter_0/reg_w_6 [3]) );
  dff_sg \filter_0/reg_w_6_reg[4]  ( .D(n43604), .CP(clk), .Q(
        \filter_0/reg_w_6 [4]) );
  dff_sg \filter_0/reg_w_6_reg[5]  ( .D(n43605), .CP(clk), .Q(
        \filter_0/reg_w_6 [5]) );
  dff_sg \filter_0/reg_w_6_reg[6]  ( .D(n43601), .CP(clk), .Q(
        \filter_0/reg_w_6 [6]) );
  dff_sg \filter_0/reg_w_6_reg[7]  ( .D(n43602), .CP(clk), .Q(
        \filter_0/reg_w_6 [7]) );
  dff_sg \filter_0/reg_w_6_reg[8]  ( .D(n43610), .CP(clk), .Q(
        \filter_0/reg_w_6 [8]) );
  dff_sg \filter_0/reg_w_6_reg[9]  ( .D(n43611), .CP(clk), .Q(
        \filter_0/reg_w_6 [9]) );
  dff_sg \filter_0/reg_w_6_reg[10]  ( .D(n43607), .CP(clk), .Q(
        \filter_0/reg_w_6 [10]) );
  dff_sg \filter_0/reg_w_6_reg[11]  ( .D(n43608), .CP(clk), .Q(
        \filter_0/reg_w_6 [11]) );
  dff_sg \filter_0/reg_w_6_reg[12]  ( .D(n43592), .CP(clk), .Q(
        \filter_0/reg_w_6 [12]) );
  dff_sg \filter_0/reg_w_6_reg[13]  ( .D(n43593), .CP(clk), .Q(
        \filter_0/reg_w_6 [13]) );
  dff_sg \filter_0/reg_w_6_reg[14]  ( .D(n43589), .CP(clk), .Q(
        \filter_0/reg_w_6 [14]) );
  dff_sg \filter_0/reg_w_6_reg[15]  ( .D(n43590), .CP(clk), .Q(
        \filter_0/reg_w_6 [15]) );
  dff_sg \filter_0/reg_w_6_reg[16]  ( .D(n43598), .CP(clk), .Q(
        \filter_0/reg_w_6 [16]) );
  dff_sg \filter_0/reg_w_6_reg[17]  ( .D(n43599), .CP(clk), .Q(
        \filter_0/reg_w_6 [17]) );
  dff_sg \filter_0/reg_w_6_reg[18]  ( .D(n43595), .CP(clk), .Q(
        \filter_0/reg_w_6 [18]) );
  dff_sg \filter_0/reg_w_6_reg[19]  ( .D(n43596), .CP(clk), .Q(
        \filter_0/reg_w_6 [19]) );
  dff_sg \filter_0/reg_w_7_reg[0]  ( .D(n43562), .CP(clk), .Q(
        \filter_0/reg_w_7 [0]) );
  dff_sg \filter_0/reg_w_7_reg[1]  ( .D(n43563), .CP(clk), .Q(
        \filter_0/reg_w_7 [1]) );
  dff_sg \filter_0/reg_w_7_reg[2]  ( .D(n43559), .CP(clk), .Q(
        \filter_0/reg_w_7 [2]) );
  dff_sg \filter_0/reg_w_7_reg[3]  ( .D(n43560), .CP(clk), .Q(
        \filter_0/reg_w_7 [3]) );
  dff_sg \filter_0/reg_w_7_reg[4]  ( .D(n43553), .CP(clk), .Q(
        \filter_0/reg_w_7 [4]) );
  dff_sg \filter_0/reg_w_7_reg[5]  ( .D(n43986), .CP(clk), .Q(
        \filter_0/reg_w_7 [5]) );
  dff_sg \filter_0/reg_w_7_reg[6]  ( .D(n43541), .CP(clk), .Q(
        \filter_0/reg_w_7 [6]) );
  dff_sg \filter_0/reg_w_7_reg[7]  ( .D(n43542), .CP(clk), .Q(
        \filter_0/reg_w_7 [7]) );
  dff_sg \filter_0/reg_w_7_reg[8]  ( .D(n44063), .CP(clk), .Q(
        \filter_0/reg_w_7 [8]) );
  dff_sg \filter_0/reg_w_7_reg[9]  ( .D(n43961), .CP(clk), .Q(
        \filter_0/reg_w_7 [9]) );
  dff_sg \filter_0/reg_w_7_reg[10]  ( .D(n43973), .CP(clk), .Q(
        \filter_0/reg_w_7 [10]) );
  dff_sg \filter_0/reg_w_7_reg[11]  ( .D(n43978), .CP(clk), .Q(
        \filter_0/reg_w_7 [11]) );
  dff_sg \filter_0/reg_w_7_reg[12]  ( .D(n43554), .CP(clk), .Q(
        \filter_0/reg_w_7 [12]) );
  dff_sg \filter_0/reg_w_7_reg[13]  ( .D(n43555), .CP(clk), .Q(
        \filter_0/reg_w_7 [13]) );
  dff_sg \filter_0/reg_w_7_reg[14]  ( .D(n44106), .CP(clk), .Q(
        \filter_0/reg_w_7 [14]) );
  dff_sg \filter_0/reg_w_7_reg[15]  ( .D(n44107), .CP(clk), .Q(
        \filter_0/reg_w_7 [15]) );
  dff_sg \filter_0/reg_w_7_reg[16]  ( .D(n44103), .CP(clk), .Q(
        \filter_0/reg_w_7 [16]) );
  dff_sg \filter_0/reg_w_7_reg[17]  ( .D(n44104), .CP(clk), .Q(
        \filter_0/reg_w_7 [17]) );
  dff_sg \filter_0/reg_w_7_reg[18]  ( .D(n43547), .CP(clk), .Q(
        \filter_0/reg_w_7 [18]) );
  dff_sg \filter_0/reg_w_7_reg[19]  ( .D(n43548), .CP(clk), .Q(
        \filter_0/reg_w_7 [19]) );
  dff_sg \filter_0/reg_w_8_reg[0]  ( .D(n44097), .CP(clk), .Q(
        \filter_0/reg_w_8 [0]) );
  dff_sg \filter_0/reg_w_8_reg[1]  ( .D(n44098), .CP(clk), .Q(
        \filter_0/reg_w_8 [1]) );
  dff_sg \filter_0/reg_w_8_reg[2]  ( .D(n43520), .CP(clk), .Q(
        \filter_0/reg_w_8 [2]) );
  dff_sg \filter_0/reg_w_8_reg[3]  ( .D(n43521), .CP(clk), .Q(
        \filter_0/reg_w_8 [3]) );
  dff_sg \filter_0/reg_w_8_reg[4]  ( .D(n43502), .CP(clk), .Q(
        \filter_0/reg_w_8 [4]) );
  dff_sg \filter_0/reg_w_8_reg[5]  ( .D(n43503), .CP(clk), .Q(
        \filter_0/reg_w_8 [5]) );
  dff_sg \filter_0/reg_w_8_reg[6]  ( .D(n43499), .CP(clk), .Q(
        \filter_0/reg_w_8 [6]) );
  dff_sg \filter_0/reg_w_8_reg[7]  ( .D(n43500), .CP(clk), .Q(
        \filter_0/reg_w_8 [7]) );
  dff_sg \filter_0/reg_w_8_reg[8]  ( .D(n43508), .CP(clk), .Q(
        \filter_0/reg_w_8 [8]) );
  dff_sg \filter_0/reg_w_8_reg[9]  ( .D(n43509), .CP(clk), .Q(
        \filter_0/reg_w_8 [9]) );
  dff_sg \filter_0/reg_w_8_reg[10]  ( .D(n43505), .CP(clk), .Q(
        \filter_0/reg_w_8 [10]) );
  dff_sg \filter_0/reg_w_8_reg[11]  ( .D(n43506), .CP(clk), .Q(
        \filter_0/reg_w_8 [11]) );
  dff_sg \filter_0/reg_w_8_reg[12]  ( .D(n43675), .CP(clk), .Q(
        \filter_0/reg_w_8 [12]) );
  dff_sg \filter_0/reg_w_8_reg[13]  ( .D(n43676), .CP(clk), .Q(
        \filter_0/reg_w_8 [13]) );
  dff_sg \filter_0/reg_w_8_reg[14]  ( .D(n43672), .CP(clk), .Q(
        \filter_0/reg_w_8 [14]) );
  dff_sg \filter_0/reg_w_8_reg[15]  ( .D(n43673), .CP(clk), .Q(
        \filter_0/reg_w_8 [15]) );
  dff_sg \filter_0/reg_w_8_reg[16]  ( .D(n43681), .CP(clk), .Q(
        \filter_0/reg_w_8 [16]) );
  dff_sg \filter_0/reg_w_8_reg[17]  ( .D(n43682), .CP(clk), .Q(
        \filter_0/reg_w_8 [17]) );
  dff_sg \filter_0/reg_w_8_reg[18]  ( .D(n43678), .CP(clk), .Q(
        \filter_0/reg_w_8 [18]) );
  dff_sg \filter_0/reg_w_8_reg[19]  ( .D(n43679), .CP(clk), .Q(
        \filter_0/reg_w_8 [19]) );
  dff_sg \filter_0/reg_w_9_reg[0]  ( .D(n43663), .CP(clk), .Q(
        \filter_0/reg_w_9 [0]) );
  dff_sg \filter_0/reg_w_9_reg[1]  ( .D(n43664), .CP(clk), .Q(
        \filter_0/reg_w_9 [1]) );
  dff_sg \filter_0/reg_w_9_reg[2]  ( .D(n43660), .CP(clk), .Q(
        \filter_0/reg_w_9 [2]) );
  dff_sg \filter_0/reg_w_9_reg[3]  ( .D(n43661), .CP(clk), .Q(
        \filter_0/reg_w_9 [3]) );
  dff_sg \filter_0/reg_w_9_reg[4]  ( .D(n43669), .CP(clk), .Q(
        \filter_0/reg_w_9 [4]) );
  dff_sg \filter_0/reg_w_9_reg[5]  ( .D(n43670), .CP(clk), .Q(
        \filter_0/reg_w_9 [5]) );
  dff_sg \filter_0/reg_w_9_reg[6]  ( .D(n43666), .CP(clk), .Q(
        \filter_0/reg_w_9 [6]) );
  dff_sg \filter_0/reg_w_9_reg[7]  ( .D(n43667), .CP(clk), .Q(
        \filter_0/reg_w_9 [7]) );
  dff_sg \filter_0/reg_w_9_reg[8]  ( .D(n43698), .CP(clk), .Q(
        \filter_0/reg_w_9 [8]) );
  dff_sg \filter_0/reg_w_9_reg[9]  ( .D(n43699), .CP(clk), .Q(
        \filter_0/reg_w_9 [9]) );
  dff_sg \filter_0/reg_w_9_reg[10]  ( .D(n43695), .CP(clk), .Q(
        \filter_0/reg_w_9 [10]) );
  dff_sg \filter_0/reg_w_9_reg[11]  ( .D(n43696), .CP(clk), .Q(
        \filter_0/reg_w_9 [11]) );
  dff_sg \filter_0/reg_w_9_reg[12]  ( .D(n43703), .CP(clk), .Q(
        \filter_0/reg_w_9 [12]) );
  dff_sg \filter_0/reg_w_9_reg[13]  ( .D(n43704), .CP(clk), .Q(
        \filter_0/reg_w_9 [13]) );
  dff_sg \filter_0/reg_w_9_reg[14]  ( .D(n43700), .CP(clk), .Q(
        \filter_0/reg_w_9 [14]) );
  dff_sg \filter_0/reg_w_9_reg[15]  ( .D(n43701), .CP(clk), .Q(
        \filter_0/reg_w_9 [15]) );
  dff_sg \filter_0/reg_w_9_reg[16]  ( .D(n43686), .CP(clk), .Q(
        \filter_0/reg_w_9 [16]) );
  dff_sg \filter_0/reg_w_9_reg[17]  ( .D(n43687), .CP(clk), .Q(
        \filter_0/reg_w_9 [17]) );
  dff_sg \filter_0/reg_w_9_reg[18]  ( .D(n43683), .CP(clk), .Q(
        \filter_0/reg_w_9 [18]) );
  dff_sg \filter_0/reg_w_9_reg[19]  ( .D(n43684), .CP(clk), .Q(
        \filter_0/reg_w_9 [19]) );
  dff_sg \filter_0/reg_w_10_reg[0]  ( .D(n43692), .CP(clk), .Q(
        \filter_0/reg_w_10 [0]) );
  dff_sg \filter_0/reg_w_10_reg[1]  ( .D(n43693), .CP(clk), .Q(
        \filter_0/reg_w_10 [1]) );
  dff_sg \filter_0/reg_w_10_reg[2]  ( .D(n43689), .CP(clk), .Q(
        \filter_0/reg_w_10 [2]) );
  dff_sg \filter_0/reg_w_10_reg[3]  ( .D(n43690), .CP(clk), .Q(
        \filter_0/reg_w_10 [3]) );
  dff_sg \filter_0/reg_w_10_reg[4]  ( .D(n43628), .CP(clk), .Q(
        \filter_0/reg_w_10 [4]) );
  dff_sg \filter_0/reg_w_10_reg[5]  ( .D(n43629), .CP(clk), .Q(
        \filter_0/reg_w_10 [5]) );
  dff_sg \filter_0/reg_w_10_reg[6]  ( .D(n43625), .CP(clk), .Q(
        \filter_0/reg_w_10 [6]) );
  dff_sg \filter_0/reg_w_10_reg[7]  ( .D(n43626), .CP(clk), .Q(
        \filter_0/reg_w_10 [7]) );
  dff_sg \filter_0/reg_w_10_reg[8]  ( .D(n43634), .CP(clk), .Q(
        \filter_0/reg_w_10 [8]) );
  dff_sg \filter_0/reg_w_10_reg[9]  ( .D(n43635), .CP(clk), .Q(
        \filter_0/reg_w_10 [9]) );
  dff_sg \filter_0/reg_w_10_reg[10]  ( .D(n43631), .CP(clk), .Q(
        \filter_0/reg_w_10 [10]) );
  dff_sg \filter_0/reg_w_10_reg[11]  ( .D(n43632), .CP(clk), .Q(
        \filter_0/reg_w_10 [11]) );
  dff_sg \filter_0/reg_w_10_reg[12]  ( .D(n43616), .CP(clk), .Q(
        \filter_0/reg_w_10 [12]) );
  dff_sg \filter_0/reg_w_10_reg[13]  ( .D(n43617), .CP(clk), .Q(
        \filter_0/reg_w_10 [13]) );
  dff_sg \filter_0/reg_w_10_reg[14]  ( .D(n43613), .CP(clk), .Q(
        \filter_0/reg_w_10 [14]) );
  dff_sg \filter_0/reg_w_10_reg[15]  ( .D(n43614), .CP(clk), .Q(
        \filter_0/reg_w_10 [15]) );
  dff_sg \filter_0/reg_w_10_reg[16]  ( .D(n43622), .CP(clk), .Q(
        \filter_0/reg_w_10 [16]) );
  dff_sg \filter_0/reg_w_10_reg[17]  ( .D(n43623), .CP(clk), .Q(
        \filter_0/reg_w_10 [17]) );
  dff_sg \filter_0/reg_w_10_reg[18]  ( .D(n43619), .CP(clk), .Q(
        \filter_0/reg_w_10 [18]) );
  dff_sg \filter_0/reg_w_10_reg[19]  ( .D(n43620), .CP(clk), .Q(
        \filter_0/reg_w_10 [19]) );
  dff_sg \filter_0/reg_w_11_reg[0]  ( .D(n43652), .CP(clk), .Q(
        \filter_0/reg_w_11 [0]) );
  dff_sg \filter_0/reg_w_11_reg[1]  ( .D(n43653), .CP(clk), .Q(
        \filter_0/reg_w_11 [1]) );
  dff_sg \filter_0/reg_w_11_reg[2]  ( .D(n43649), .CP(clk), .Q(
        \filter_0/reg_w_11 [2]) );
  dff_sg \filter_0/reg_w_11_reg[3]  ( .D(n43650), .CP(clk), .Q(
        \filter_0/reg_w_11 [3]) );
  dff_sg \filter_0/reg_w_11_reg[4]  ( .D(n43658), .CP(clk), .Q(
        \filter_0/reg_w_11 [4]) );
  dff_sg \filter_0/reg_w_11_reg[5]  ( .D(n43659), .CP(clk), .Q(
        \filter_0/reg_w_11 [5]) );
  dff_sg \filter_0/reg_w_11_reg[6]  ( .D(n43655), .CP(clk), .Q(
        \filter_0/reg_w_11 [6]) );
  dff_sg \filter_0/reg_w_11_reg[7]  ( .D(n43656), .CP(clk), .Q(
        \filter_0/reg_w_11 [7]) );
  dff_sg \filter_0/reg_w_11_reg[8]  ( .D(n43640), .CP(clk), .Q(
        \filter_0/reg_w_11 [8]) );
  dff_sg \filter_0/reg_w_11_reg[9]  ( .D(n43641), .CP(clk), .Q(
        \filter_0/reg_w_11 [9]) );
  dff_sg \filter_0/reg_w_11_reg[10]  ( .D(n43637), .CP(clk), .Q(
        \filter_0/reg_w_11 [10]) );
  dff_sg \filter_0/reg_w_11_reg[11]  ( .D(n43638), .CP(clk), .Q(
        \filter_0/reg_w_11 [11]) );
  dff_sg \filter_0/reg_w_11_reg[12]  ( .D(n43646), .CP(clk), .Q(
        \filter_0/reg_w_11 [12]) );
  dff_sg \filter_0/reg_w_11_reg[13]  ( .D(n43647), .CP(clk), .Q(
        \filter_0/reg_w_11 [13]) );
  dff_sg \filter_0/reg_w_11_reg[14]  ( .D(n43643), .CP(clk), .Q(
        \filter_0/reg_w_11 [14]) );
  dff_sg \filter_0/reg_w_11_reg[15]  ( .D(n43644), .CP(clk), .Q(
        \filter_0/reg_w_11 [15]) );
  dff_sg \filter_0/reg_w_11_reg[16]  ( .D(n43885), .CP(clk), .Q(
        \filter_0/reg_w_11 [16]) );
  dff_sg \filter_0/reg_w_11_reg[17]  ( .D(n43888), .CP(clk), .Q(
        \filter_0/reg_w_11 [17]) );
  dff_sg \filter_0/reg_w_11_reg[18]  ( .D(n43897), .CP(clk), .Q(
        \filter_0/reg_w_11 [18]) );
  dff_sg \filter_0/reg_w_11_reg[19]  ( .D(n43891), .CP(clk), .Q(
        \filter_0/reg_w_11 [19]) );
  dff_sg \filter_0/reg_w_12_reg[0]  ( .D(n43871), .CP(clk), .Q(
        \filter_0/reg_w_12 [0]) );
  dff_sg \filter_0/reg_w_12_reg[1]  ( .D(n43874), .CP(clk), .Q(
        \filter_0/reg_w_12 [1]) );
  dff_sg \filter_0/reg_w_12_reg[2]  ( .D(n43877), .CP(clk), .Q(
        \filter_0/reg_w_12 [2]) );
  dff_sg \filter_0/reg_w_12_reg[3]  ( .D(n43879), .CP(clk), .Q(
        \filter_0/reg_w_12 [3]) );
  dff_sg \filter_0/reg_w_12_reg[4]  ( .D(n43850), .CP(clk), .Q(
        \filter_0/reg_w_12 [4]) );
  dff_sg \filter_0/reg_w_12_reg[5]  ( .D(n43853), .CP(clk), .Q(
        \filter_0/reg_w_12 [5]) );
  dff_sg \filter_0/reg_w_12_reg[6]  ( .D(n43859), .CP(clk), .Q(
        \filter_0/reg_w_12 [6]) );
  dff_sg \filter_0/reg_w_12_reg[7]  ( .D(n43862), .CP(clk), .Q(
        \filter_0/reg_w_12 [7]) );
  dff_sg \filter_0/reg_w_12_reg[8]  ( .D(n43906), .CP(clk), .Q(
        \filter_0/reg_w_12 [8]) );
  dff_sg \filter_0/reg_w_12_reg[9]  ( .D(n43909), .CP(clk), .Q(
        \filter_0/reg_w_12 [9]) );
  dff_sg \filter_0/reg_w_12_reg[10]  ( .D(n43538), .CP(clk), .Q(
        \filter_0/reg_w_12 [10]) );
  dff_sg \filter_0/reg_w_12_reg[11]  ( .D(n43912), .CP(clk), .Q(
        \filter_0/reg_w_12 [11]) );
  dff_sg \filter_0/reg_w_12_reg[12]  ( .D(n43956), .CP(clk), .Q(
        \filter_0/reg_w_12 [12]) );
  dff_sg \filter_0/reg_w_12_reg[13]  ( .D(n43964), .CP(clk), .Q(
        \filter_0/reg_w_12 [13]) );
  dff_sg \filter_0/reg_w_12_reg[14]  ( .D(n43983), .CP(clk), .Q(
        \filter_0/reg_w_12 [14]) );
  dff_sg \filter_0/reg_w_12_reg[15]  ( .D(n43989), .CP(clk), .Q(
        \filter_0/reg_w_12 [15]) );
  dff_sg \filter_0/reg_w_12_reg[16]  ( .D(n43967), .CP(clk), .Q(
        \filter_0/reg_w_12 [16]) );
  dff_sg \filter_0/reg_w_12_reg[17]  ( .D(n43969), .CP(clk), .Q(
        \filter_0/reg_w_12 [17]) );
  dff_sg \filter_0/reg_w_12_reg[18]  ( .D(n43544), .CP(clk), .Q(
        \filter_0/reg_w_12 [18]) );
  dff_sg \filter_0/reg_w_12_reg[19]  ( .D(n43971), .CP(clk), .Q(
        \filter_0/reg_w_12 [19]) );
  dff_sg \filter_0/reg_w_13_reg[0]  ( .D(n43930), .CP(clk), .Q(
        \filter_0/reg_w_13 [0]) );
  dff_sg \filter_0/reg_w_13_reg[1]  ( .D(n43933), .CP(clk), .Q(
        \filter_0/reg_w_13 [1]) );
  dff_sg \filter_0/reg_w_13_reg[2]  ( .D(n43942), .CP(clk), .Q(
        \filter_0/reg_w_13 [2]) );
  dff_sg \filter_0/reg_w_13_reg[3]  ( .D(n43936), .CP(clk), .Q(
        \filter_0/reg_w_13 [3]) );
  dff_sg \filter_0/reg_w_13_reg[4]  ( .D(n43915), .CP(clk), .Q(
        \filter_0/reg_w_13 [4]) );
  dff_sg \filter_0/reg_w_13_reg[5]  ( .D(n43918), .CP(clk), .Q(
        \filter_0/reg_w_13 [5]) );
  dff_sg \filter_0/reg_w_13_reg[6]  ( .D(n43921), .CP(clk), .Q(
        \filter_0/reg_w_13 [6]) );
  dff_sg \filter_0/reg_w_13_reg[7]  ( .D(n43924), .CP(clk), .Q(
        \filter_0/reg_w_13 [7]) );
  dff_sg \filter_0/reg_w_13_reg[8]  ( .D(n43551), .CP(clk), .Q(
        \filter_0/reg_w_13 [8]) );
  dff_sg \filter_0/reg_w_13_reg[9]  ( .D(n43642), .CP(clk), .Q(
        \filter_0/reg_w_13 [9]) );
  dff_sg \filter_0/reg_w_13_reg[10]  ( .D(n43774), .CP(clk), .Q(
        \filter_0/reg_w_13 [10]) );
  dff_sg \filter_0/reg_w_13_reg[11]  ( .D(n43768), .CP(clk), .Q(
        \filter_0/reg_w_13 [11]) );
  dff_sg \filter_0/reg_w_13_reg[12]  ( .D(n43529), .CP(clk), .Q(
        \filter_0/reg_w_13 [12]) );
  dff_sg \filter_0/reg_w_13_reg[13]  ( .D(n43522), .CP(clk), .Q(
        \filter_0/reg_w_13 [13]) );
  dff_sg \filter_0/reg_w_13_reg[14]  ( .D(n43533), .CP(clk), .Q(
        \filter_0/reg_w_13 [14]) );
  dff_sg \filter_0/reg_w_13_reg[15]  ( .D(n43868), .CP(clk), .Q(
        \filter_0/reg_w_13 [15]) );
  dff_sg \filter_0/reg_w_13_reg[16]  ( .D(n43756), .CP(clk), .Q(
        \filter_0/reg_w_13 [16]) );
  dff_sg \filter_0/reg_w_13_reg[17]  ( .D(n43759), .CP(clk), .Q(
        \filter_0/reg_w_13 [17]) );
  dff_sg \filter_0/reg_w_13_reg[18]  ( .D(n43762), .CP(clk), .Q(
        \filter_0/reg_w_13 [18]) );
  dff_sg \filter_0/reg_w_13_reg[19]  ( .D(n43765), .CP(clk), .Q(
        \filter_0/reg_w_13 [19]) );
  dff_sg \filter_0/reg_w_14_reg[0]  ( .D(n43783), .CP(clk), .Q(
        \filter_0/reg_w_14 [0]) );
  dff_sg \filter_0/reg_w_14_reg[1]  ( .D(n43786), .CP(clk), .Q(
        \filter_0/reg_w_14 [1]) );
  dff_sg \filter_0/reg_w_14_reg[2]  ( .D(n43531), .CP(clk), .Q(
        \filter_0/reg_w_14 [2]) );
  dff_sg \filter_0/reg_w_14_reg[3]  ( .D(n43532), .CP(clk), .Q(
        \filter_0/reg_w_14 [3]) );
  dff_sg \filter_0/reg_w_14_reg[4]  ( .D(n43523), .CP(clk), .Q(
        \filter_0/reg_w_14 [4]) );
  dff_sg \filter_0/reg_w_14_reg[5]  ( .D(n43865), .CP(clk), .Q(
        \filter_0/reg_w_14 [5]) );
  dff_sg \filter_0/reg_w_14_reg[6]  ( .D(n43792), .CP(clk), .Q(
        \filter_0/reg_w_14 [6]) );
  dff_sg \filter_0/reg_w_14_reg[7]  ( .D(n43795), .CP(clk), .Q(
        \filter_0/reg_w_14 [7]) );
  dff_sg \filter_0/reg_w_14_reg[8]  ( .D(n43839), .CP(clk), .Q(
        \filter_0/reg_w_14 [8]) );
  dff_sg \filter_0/reg_w_14_reg[9]  ( .D(n43841), .CP(clk), .Q(
        \filter_0/reg_w_14 [9]) );
  dff_sg \filter_0/reg_w_14_reg[10]  ( .D(n43844), .CP(clk), .Q(
        \filter_0/reg_w_14 [10]) );
  dff_sg \filter_0/reg_w_14_reg[11]  ( .D(n43847), .CP(clk), .Q(
        \filter_0/reg_w_14 [11]) );
  dff_sg \filter_0/reg_w_14_reg[12]  ( .D(n43819), .CP(clk), .Q(
        \filter_0/reg_w_14 [12]) );
  dff_sg \filter_0/reg_w_14_reg[13]  ( .D(n43822), .CP(clk), .Q(
        \filter_0/reg_w_14 [13]) );
  dff_sg \filter_0/reg_w_14_reg[14]  ( .D(n43831), .CP(clk), .Q(
        \filter_0/reg_w_14 [14]) );
  dff_sg \filter_0/reg_w_14_reg[15]  ( .D(n43825), .CP(clk), .Q(
        \filter_0/reg_w_14 [15]) );
  dff_sg \filter_0/reg_w_14_reg[16]  ( .D(n43804), .CP(clk), .Q(
        \filter_0/reg_w_14 [16]) );
  dff_sg \filter_0/reg_w_14_reg[17]  ( .D(n43807), .CP(clk), .Q(
        \filter_0/reg_w_14 [17]) );
  dff_sg \filter_0/reg_w_14_reg[18]  ( .D(n43810), .CP(clk), .Q(
        \filter_0/reg_w_14 [18]) );
  dff_sg \filter_0/reg_w_14_reg[19]  ( .D(n43813), .CP(clk), .Q(
        \filter_0/reg_w_14 [19]) );
  dff_sg \filter_0/reg_w_15_reg[0]  ( .D(n43992), .CP(clk), .Q(
        \filter_0/reg_w_15 [0]) );
  dff_sg \filter_0/reg_w_15_reg[1]  ( .D(n43995), .CP(clk), .Q(
        \filter_0/reg_w_15 [1]) );
  dff_sg \filter_0/reg_w_15_reg[2]  ( .D(n44002), .CP(clk), .Q(
        \filter_0/reg_w_15 [2]) );
  dff_sg \filter_0/reg_w_15_reg[3]  ( .D(n43996), .CP(clk), .Q(
        \filter_0/reg_w_15 [3]) );
  dff_sg \filter_0/reg_w_15_reg[4]  ( .D(n44051), .CP(clk), .Q(
        \filter_0/reg_w_15 [4]) );
  dff_sg \filter_0/reg_w_15_reg[5]  ( .D(n44054), .CP(clk), .Q(
        \filter_0/reg_w_15 [5]) );
  dff_sg \filter_0/reg_w_15_reg[6]  ( .D(n43953), .CP(clk), .Q(
        \filter_0/reg_w_15 [6]) );
  dff_sg \filter_0/reg_w_15_reg[7]  ( .D(n43959), .CP(clk), .Q(
        \filter_0/reg_w_15 [7]) );
  dff_sg \filter_0/reg_w_15_reg[8]  ( .D(n44021), .CP(clk), .Q(
        \filter_0/reg_w_15 [8]) );
  dff_sg \filter_0/reg_w_15_reg[9]  ( .D(n44023), .CP(clk), .Q(
        \filter_0/reg_w_15 [9]) );
  dff_sg \filter_0/reg_w_15_reg[10]  ( .D(n44031), .CP(clk), .Q(
        \filter_0/reg_w_15 [10]) );
  dff_sg \filter_0/reg_w_15_reg[11]  ( .D(n44034), .CP(clk), .Q(
        \filter_0/reg_w_15 [11]) );
  dff_sg \filter_0/reg_w_15_reg[12]  ( .D(n44010), .CP(clk), .Q(
        \filter_0/reg_w_15 [12]) );
  dff_sg \filter_0/reg_w_15_reg[13]  ( .D(n44013), .CP(clk), .Q(
        \filter_0/reg_w_15 [13]) );
  dff_sg \filter_0/reg_w_15_reg[14]  ( .D(n43550), .CP(clk), .Q(
        \filter_0/reg_w_15 [14]) );
  dff_sg \filter_0/reg_w_15_reg[15]  ( .D(n44016), .CP(clk), .Q(
        \filter_0/reg_w_15 [15]) );
  dff_sg \filter_0/reg_w_15_reg[16]  ( .D(n44037), .CP(clk), .Q(
        \filter_0/reg_w_15 [16]) );
  dff_sg \filter_0/reg_w_15_reg[17]  ( .D(n44040), .CP(clk), .Q(
        \filter_0/reg_w_15 [17]) );
  dff_sg \filter_0/reg_w_15_reg[18]  ( .D(n44045), .CP(clk), .Q(
        \filter_0/reg_w_15 [18]) );
  dff_sg \filter_0/reg_w_15_reg[19]  ( .D(n44048), .CP(clk), .Q(
        \filter_0/reg_w_15 [19]) );
  dff_sg \filter_0/reg_o_mask_reg[0]  ( .D(\filter_0/n11596 ), .CP(clk), .Q(
        \filter_0/reg_o_mask [0]) );
  dff_sg \filter_0/reg_o_mask_reg[1]  ( .D(\filter_0/n11595 ), .CP(clk), .Q(
        \filter_0/reg_o_mask [1]) );
  dff_sg \filter_0/reg_o_mask_reg[2]  ( .D(\filter_0/n11594 ), .CP(clk), .Q(
        \filter_0/reg_o_mask [2]) );
  dff_sg \filter_0/reg_o_mask_reg[3]  ( .D(\filter_0/n11593 ), .CP(clk), .Q(
        \filter_0/reg_o_mask [3]) );
  dff_sg \filter_0/reg_o_mask_reg[4]  ( .D(\filter_0/n11592 ), .CP(clk), .Q(
        \filter_0/reg_o_mask [4]) );
  dff_sg \filter_0/reg_o_mask_reg[5]  ( .D(\filter_0/n11591 ), .CP(clk), .Q(
        \filter_0/reg_o_mask [5]) );
  dff_sg \filter_0/reg_o_mask_reg[6]  ( .D(\filter_0/n11590 ), .CP(clk), .Q(
        \filter_0/reg_o_mask [6]) );
  dff_sg \filter_0/reg_o_mask_reg[7]  ( .D(\filter_0/n11589 ), .CP(clk), .Q(
        \filter_0/reg_o_mask [7]) );
  dff_sg \filter_0/reg_o_mask_reg[8]  ( .D(\filter_0/n11588 ), .CP(clk), .Q(
        \filter_0/reg_o_mask [8]) );
  dff_sg \filter_0/reg_o_mask_reg[9]  ( .D(\filter_0/n11587 ), .CP(clk), .Q(
        \filter_0/reg_o_mask [9]) );
  dff_sg \filter_0/reg_o_mask_reg[10]  ( .D(\filter_0/n11586 ), .CP(clk), .Q(
        \filter_0/reg_o_mask [10]) );
  dff_sg \filter_0/reg_o_mask_reg[11]  ( .D(\filter_0/n11585 ), .CP(clk), .Q(
        \filter_0/reg_o_mask [11]) );
  dff_sg \filter_0/reg_o_mask_reg[12]  ( .D(\filter_0/n11584 ), .CP(clk), .Q(
        \filter_0/reg_o_mask [12]) );
  dff_sg \filter_0/reg_o_mask_reg[13]  ( .D(\filter_0/n11583 ), .CP(clk), .Q(
        \filter_0/reg_o_mask [13]) );
  dff_sg \filter_0/reg_o_mask_reg[14]  ( .D(\filter_0/n11582 ), .CP(clk), .Q(
        \filter_0/reg_o_mask [14]) );
  dff_sg \filter_0/reg_o_mask_reg[15]  ( .D(\filter_0/n11581 ), .CP(clk), .Q(
        \filter_0/reg_o_mask [15]) );
  dff_sg \filter_0/reg_o_mask_reg[16]  ( .D(\filter_0/n11580 ), .CP(clk), .Q(
        \filter_0/reg_o_mask [16]) );
  dff_sg \filter_0/reg_o_mask_reg[17]  ( .D(\filter_0/n11579 ), .CP(clk), .Q(
        \filter_0/reg_o_mask [17]) );
  dff_sg \filter_0/reg_o_mask_reg[18]  ( .D(\filter_0/n11578 ), .CP(clk), .Q(
        \filter_0/reg_o_mask [18]) );
  dff_sg \filter_0/reg_o_mask_reg[19]  ( .D(\filter_0/n11577 ), .CP(clk), .Q(
        \filter_0/reg_o_mask [19]) );
  dff_sg \filter_0/reg_o_mask_reg[20]  ( .D(\filter_0/n11576 ), .CP(clk), .Q(
        \filter_0/reg_o_mask [20]) );
  dff_sg \filter_0/reg_o_mask_reg[21]  ( .D(\filter_0/n11575 ), .CP(clk), .Q(
        \filter_0/reg_o_mask [21]) );
  dff_sg \filter_0/reg_o_mask_reg[22]  ( .D(\filter_0/n11574 ), .CP(clk), .Q(
        \filter_0/reg_o_mask [22]) );
  dff_sg \filter_0/reg_o_mask_reg[23]  ( .D(\filter_0/n11573 ), .CP(clk), .Q(
        \filter_0/reg_o_mask [23]) );
  dff_sg \filter_0/reg_o_mask_reg[24]  ( .D(\filter_0/n11572 ), .CP(clk), .Q(
        \filter_0/reg_o_mask [24]) );
  dff_sg \filter_0/reg_o_mask_reg[25]  ( .D(\filter_0/n11571 ), .CP(clk), .Q(
        \filter_0/reg_o_mask [25]) );
  dff_sg \filter_0/reg_o_mask_reg[26]  ( .D(\filter_0/n11570 ), .CP(clk), .Q(
        \filter_0/reg_o_mask [26]) );
  dff_sg \filter_0/reg_o_mask_reg[27]  ( .D(\filter_0/n11569 ), .CP(clk), .Q(
        \filter_0/reg_o_mask [27]) );
  dff_sg \filter_0/reg_o_mask_reg[28]  ( .D(\filter_0/n11568 ), .CP(clk), .Q(
        \filter_0/reg_o_mask [28]) );
  dff_sg \filter_0/reg_o_mask_reg[29]  ( .D(\filter_0/n11567 ), .CP(clk), .Q(
        \filter_0/reg_o_mask [29]) );
  dff_sg \filter_0/reg_o_mask_reg[30]  ( .D(\filter_0/n11566 ), .CP(clk), .Q(
        \filter_0/reg_o_mask [30]) );
  dff_sg \filter_0/reg_o_mask_reg[31]  ( .D(\filter_0/n11565 ), .CP(clk), .Q(
        \filter_0/reg_o_mask [31]) );
  dff_sg \filter_0/reg_xor_i_mask_reg[0]  ( .D(\filter_0/n11564 ), .CP(clk), 
        .Q(\filter_0/reg_xor_i_mask [0]) );
  dff_sg \filter_0/reg_xor_i_mask_reg[1]  ( .D(\filter_0/n11563 ), .CP(clk), 
        .Q(\filter_0/reg_xor_i_mask [1]) );
  dff_sg \filter_0/reg_xor_i_mask_reg[2]  ( .D(\filter_0/n11562 ), .CP(clk), 
        .Q(\filter_0/reg_xor_i_mask [2]) );
  dff_sg \filter_0/reg_xor_i_mask_reg[3]  ( .D(\filter_0/n11561 ), .CP(clk), 
        .Q(\filter_0/reg_xor_i_mask [3]) );
  dff_sg \filter_0/reg_xor_i_mask_reg[4]  ( .D(\filter_0/n11560 ), .CP(clk), 
        .Q(\filter_0/reg_xor_i_mask [4]) );
  dff_sg \filter_0/reg_xor_i_mask_reg[5]  ( .D(\filter_0/n11559 ), .CP(clk), 
        .Q(\filter_0/reg_xor_i_mask [5]) );
  dff_sg \filter_0/reg_xor_i_mask_reg[6]  ( .D(\filter_0/n11558 ), .CP(clk), 
        .Q(\filter_0/reg_xor_i_mask [6]) );
  dff_sg \filter_0/reg_xor_i_mask_reg[7]  ( .D(\filter_0/n11557 ), .CP(clk), 
        .Q(\filter_0/reg_xor_i_mask [7]) );
  dff_sg \filter_0/reg_xor_i_mask_reg[8]  ( .D(\filter_0/n11556 ), .CP(clk), 
        .Q(\filter_0/reg_xor_i_mask [8]) );
  dff_sg \filter_0/reg_xor_i_mask_reg[9]  ( .D(\filter_0/n11555 ), .CP(clk), 
        .Q(\filter_0/reg_xor_i_mask [9]) );
  dff_sg \filter_0/reg_xor_i_mask_reg[10]  ( .D(\filter_0/n11554 ), .CP(clk), 
        .Q(\filter_0/reg_xor_i_mask [10]) );
  dff_sg \filter_0/reg_xor_i_mask_reg[11]  ( .D(\filter_0/n11553 ), .CP(clk), 
        .Q(\filter_0/reg_xor_i_mask [11]) );
  dff_sg \filter_0/reg_xor_i_mask_reg[12]  ( .D(\filter_0/n11552 ), .CP(clk), 
        .Q(\filter_0/reg_xor_i_mask [12]) );
  dff_sg \filter_0/reg_xor_i_mask_reg[13]  ( .D(\filter_0/n11551 ), .CP(clk), 
        .Q(\filter_0/reg_xor_i_mask [13]) );
  dff_sg \filter_0/reg_xor_i_mask_reg[14]  ( .D(\filter_0/n11550 ), .CP(clk), 
        .Q(\filter_0/reg_xor_i_mask [14]) );
  dff_sg \filter_0/reg_xor_i_mask_reg[15]  ( .D(\filter_0/n11549 ), .CP(clk), 
        .Q(\filter_0/reg_xor_i_mask [15]) );
  dff_sg \filter_0/reg_xor_i_mask_reg[16]  ( .D(\filter_0/n11548 ), .CP(clk), 
        .Q(\filter_0/reg_xor_i_mask [16]) );
  dff_sg \filter_0/reg_xor_i_mask_reg[17]  ( .D(\filter_0/n11547 ), .CP(clk), 
        .Q(\filter_0/reg_xor_i_mask [17]) );
  dff_sg \filter_0/reg_xor_i_mask_reg[18]  ( .D(\filter_0/n11546 ), .CP(clk), 
        .Q(\filter_0/reg_xor_i_mask [18]) );
  dff_sg \filter_0/reg_xor_i_mask_reg[19]  ( .D(\filter_0/n11545 ), .CP(clk), 
        .Q(\filter_0/reg_xor_i_mask [19]) );
  dff_sg \filter_0/reg_xor_i_mask_reg[20]  ( .D(\filter_0/n11544 ), .CP(clk), 
        .Q(\filter_0/reg_xor_i_mask [20]) );
  dff_sg \filter_0/reg_xor_i_mask_reg[21]  ( .D(\filter_0/n11543 ), .CP(clk), 
        .Q(\filter_0/reg_xor_i_mask [21]) );
  dff_sg \filter_0/reg_xor_i_mask_reg[22]  ( .D(\filter_0/n11542 ), .CP(clk), 
        .Q(\filter_0/reg_xor_i_mask [22]) );
  dff_sg \filter_0/reg_xor_i_mask_reg[23]  ( .D(\filter_0/n11541 ), .CP(clk), 
        .Q(\filter_0/reg_xor_i_mask [23]) );
  dff_sg \filter_0/reg_xor_i_mask_reg[24]  ( .D(\filter_0/n11540 ), .CP(clk), 
        .Q(\filter_0/reg_xor_i_mask [24]) );
  dff_sg \filter_0/reg_xor_i_mask_reg[25]  ( .D(\filter_0/n11539 ), .CP(clk), 
        .Q(\filter_0/reg_xor_i_mask [25]) );
  dff_sg \filter_0/reg_xor_i_mask_reg[26]  ( .D(\filter_0/n11538 ), .CP(clk), 
        .Q(\filter_0/reg_xor_i_mask [26]) );
  dff_sg \filter_0/reg_xor_i_mask_reg[27]  ( .D(\filter_0/n11537 ), .CP(clk), 
        .Q(\filter_0/reg_xor_i_mask [27]) );
  dff_sg \filter_0/reg_xor_i_mask_reg[28]  ( .D(\filter_0/n11536 ), .CP(clk), 
        .Q(\filter_0/reg_xor_i_mask [28]) );
  dff_sg \filter_0/reg_xor_i_mask_reg[29]  ( .D(\filter_0/n11535 ), .CP(clk), 
        .Q(\filter_0/reg_xor_i_mask [29]) );
  dff_sg \filter_0/reg_xor_i_mask_reg[30]  ( .D(\filter_0/n11534 ), .CP(clk), 
        .Q(\filter_0/reg_xor_i_mask [30]) );
  dff_sg \filter_0/reg_xor_i_mask_reg[31]  ( .D(\filter_0/n11533 ), .CP(clk), 
        .Q(\filter_0/reg_xor_i_mask [31]) );
  dff_sg \filter_0/reg_xor_w_mask_reg[0]  ( .D(\filter_0/n11532 ), .CP(clk), 
        .Q(\filter_0/reg_xor_w_mask [0]) );
  dff_sg \filter_0/reg_xor_w_mask_reg[1]  ( .D(\filter_0/n11531 ), .CP(clk), 
        .Q(\filter_0/reg_xor_w_mask [1]) );
  dff_sg \filter_0/reg_xor_w_mask_reg[2]  ( .D(\filter_0/n11530 ), .CP(clk), 
        .Q(\filter_0/reg_xor_w_mask [2]) );
  dff_sg \filter_0/reg_xor_w_mask_reg[3]  ( .D(\filter_0/n11529 ), .CP(clk), 
        .Q(\filter_0/reg_xor_w_mask [3]) );
  dff_sg \filter_0/reg_xor_w_mask_reg[4]  ( .D(\filter_0/n11528 ), .CP(clk), 
        .Q(\filter_0/reg_xor_w_mask [4]) );
  dff_sg \filter_0/reg_xor_w_mask_reg[5]  ( .D(\filter_0/n11527 ), .CP(clk), 
        .Q(\filter_0/reg_xor_w_mask [5]) );
  dff_sg \filter_0/reg_xor_w_mask_reg[6]  ( .D(\filter_0/n11526 ), .CP(clk), 
        .Q(\filter_0/reg_xor_w_mask [6]) );
  dff_sg \filter_0/reg_xor_w_mask_reg[7]  ( .D(\filter_0/n11525 ), .CP(clk), 
        .Q(\filter_0/reg_xor_w_mask [7]) );
  dff_sg \filter_0/reg_xor_w_mask_reg[8]  ( .D(\filter_0/n11524 ), .CP(clk), 
        .Q(\filter_0/reg_xor_w_mask [8]) );
  dff_sg \filter_0/reg_xor_w_mask_reg[9]  ( .D(\filter_0/n11523 ), .CP(clk), 
        .Q(\filter_0/reg_xor_w_mask [9]) );
  dff_sg \filter_0/reg_xor_w_mask_reg[10]  ( .D(\filter_0/n11522 ), .CP(clk), 
        .Q(\filter_0/reg_xor_w_mask [10]) );
  dff_sg \filter_0/reg_xor_w_mask_reg[11]  ( .D(\filter_0/n11521 ), .CP(clk), 
        .Q(\filter_0/reg_xor_w_mask [11]) );
  dff_sg \filter_0/reg_xor_w_mask_reg[12]  ( .D(\filter_0/n11520 ), .CP(clk), 
        .Q(\filter_0/reg_xor_w_mask [12]) );
  dff_sg \filter_0/reg_xor_w_mask_reg[13]  ( .D(\filter_0/n11519 ), .CP(clk), 
        .Q(\filter_0/reg_xor_w_mask [13]) );
  dff_sg \filter_0/reg_xor_w_mask_reg[14]  ( .D(\filter_0/n11518 ), .CP(clk), 
        .Q(\filter_0/reg_xor_w_mask [14]) );
  dff_sg \filter_0/reg_xor_w_mask_reg[15]  ( .D(\filter_0/n11517 ), .CP(clk), 
        .Q(\filter_0/reg_xor_w_mask [15]) );
  dff_sg \filter_0/reg_xor_w_mask_reg[16]  ( .D(\filter_0/n11516 ), .CP(clk), 
        .Q(\filter_0/reg_xor_w_mask [16]) );
  dff_sg \filter_0/reg_xor_w_mask_reg[17]  ( .D(\filter_0/n11515 ), .CP(clk), 
        .Q(\filter_0/reg_xor_w_mask [17]) );
  dff_sg \filter_0/reg_xor_w_mask_reg[18]  ( .D(\filter_0/n11514 ), .CP(clk), 
        .Q(\filter_0/reg_xor_w_mask [18]) );
  dff_sg \filter_0/reg_xor_w_mask_reg[19]  ( .D(\filter_0/n11513 ), .CP(clk), 
        .Q(\filter_0/reg_xor_w_mask [19]) );
  dff_sg \filter_0/reg_xor_w_mask_reg[20]  ( .D(\filter_0/n11512 ), .CP(clk), 
        .Q(\filter_0/reg_xor_w_mask [20]) );
  dff_sg \filter_0/reg_xor_w_mask_reg[21]  ( .D(\filter_0/n11511 ), .CP(clk), 
        .Q(\filter_0/reg_xor_w_mask [21]) );
  dff_sg \filter_0/reg_xor_w_mask_reg[22]  ( .D(\filter_0/n11510 ), .CP(clk), 
        .Q(\filter_0/reg_xor_w_mask [22]) );
  dff_sg \filter_0/reg_xor_w_mask_reg[23]  ( .D(\filter_0/n11509 ), .CP(clk), 
        .Q(\filter_0/reg_xor_w_mask [23]) );
  dff_sg \filter_0/reg_xor_w_mask_reg[24]  ( .D(\filter_0/n11508 ), .CP(clk), 
        .Q(\filter_0/reg_xor_w_mask [24]) );
  dff_sg \filter_0/reg_xor_w_mask_reg[25]  ( .D(\filter_0/n11507 ), .CP(clk), 
        .Q(\filter_0/reg_xor_w_mask [25]) );
  dff_sg \filter_0/reg_xor_w_mask_reg[26]  ( .D(\filter_0/n11506 ), .CP(clk), 
        .Q(\filter_0/reg_xor_w_mask [26]) );
  dff_sg \filter_0/reg_xor_w_mask_reg[27]  ( .D(\filter_0/n11505 ), .CP(clk), 
        .Q(\filter_0/reg_xor_w_mask [27]) );
  dff_sg \filter_0/reg_xor_w_mask_reg[28]  ( .D(\filter_0/n11504 ), .CP(clk), 
        .Q(\filter_0/reg_xor_w_mask [28]) );
  dff_sg \filter_0/reg_xor_w_mask_reg[29]  ( .D(\filter_0/n11503 ), .CP(clk), 
        .Q(\filter_0/reg_xor_w_mask [29]) );
  dff_sg \filter_0/reg_xor_w_mask_reg[30]  ( .D(\filter_0/n11502 ), .CP(clk), 
        .Q(\filter_0/reg_xor_w_mask [30]) );
  dff_sg \filter_0/reg_xor_w_mask_reg[31]  ( .D(\filter_0/n11501 ), .CP(clk), 
        .Q(\filter_0/reg_xor_w_mask [31]) );
  dff_sg \filter_0/m_pointer_reg[4]  ( .D(n42815), .CP(clk), .Q(\filter_0/N16 ) );
  dff_sg \filter_0/m_pointer_reg[3]  ( .D(n42817), .CP(clk), .Q(\filter_0/N15 ) );
  dff_sg \filter_0/m_pointer_reg[2]  ( .D(n42819), .CP(clk), .Q(\filter_0/N14 ) );
  dff_sg \filter_0/m_pointer_reg[1]  ( .D(n42818), .CP(clk), .Q(\filter_0/N13 ) );
  dff_sg \filter_0/m_pointer_reg[0]  ( .D(n42827), .CP(clk), .Q(\filter_0/N12 ) );
  dff_sg \filter_0/i_pointer_reg[3]  ( .D(n42828), .CP(clk), .Q(
        \filter_0/i_pointer [3]) );
  dff_sg \filter_0/i_pointer_reg[2]  ( .D(n42824), .CP(clk), .Q(
        \filter_0/i_pointer [2]) );
  dff_sg \filter_0/i_pointer_reg[1]  ( .D(n42822), .CP(clk), .Q(
        \filter_0/i_pointer [1]) );
  dff_sg \filter_0/i_pointer_reg[0]  ( .D(n42826), .CP(clk), .Q(
        \filter_0/i_pointer [0]) );
  dff_sg \filter_0/w_pointer_reg[3]  ( .D(n42816), .CP(clk), .Q(
        \filter_0/w_pointer [3]) );
  dff_sg \filter_0/w_pointer_reg[2]  ( .D(n42825), .CP(clk), .Q(
        \filter_0/w_pointer [2]) );
  dff_sg \filter_0/w_pointer_reg[1]  ( .D(n42821), .CP(clk), .Q(
        \filter_0/w_pointer [1]) );
  dff_sg \filter_0/w_pointer_reg[0]  ( .D(n42820), .CP(clk), .Q(
        \filter_0/w_pointer [0]) );
  dff_sg \filter_0/state_reg[0]  ( .D(n43469), .CP(clk), .Q(\filter_0/n17950 )
         );
  dff_sg \filter_0/state_reg[1]  ( .D(n42823), .CP(clk), .Q(\filter_0/n17949 )
         );
  dff_sg \filter_0/done_reg  ( .D(\filter_0/N1845 ), .CP(clk), .Q(
        \filter_0/done ) );
  dff_sg \shifter_0/ow_14_reg[0]  ( .D(n42680), .CP(clk), .Q(n69211) );
  dff_sg \shifter_0/ow_14_reg[1]  ( .D(n42681), .CP(clk), .Q(n69210) );
  dff_sg \shifter_0/ow_14_reg[2]  ( .D(n42677), .CP(clk), .Q(n69209) );
  dff_sg \shifter_0/ow_14_reg[3]  ( .D(n42678), .CP(clk), .Q(n69208) );
  dff_sg \shifter_0/ow_14_reg[4]  ( .D(n42686), .CP(clk), .Q(n69207) );
  dff_sg \shifter_0/ow_14_reg[5]  ( .D(n42687), .CP(clk), .Q(n69206) );
  dff_sg \shifter_0/ow_14_reg[6]  ( .D(n42683), .CP(clk), .Q(n69205) );
  dff_sg \shifter_0/ow_14_reg[7]  ( .D(n42684), .CP(clk), .Q(n69204) );
  dff_sg \shifter_0/ow_14_reg[8]  ( .D(n42668), .CP(clk), .Q(n69203) );
  dff_sg \shifter_0/ow_14_reg[9]  ( .D(n42669), .CP(clk), .Q(n69202) );
  dff_sg \shifter_0/ow_14_reg[10]  ( .D(n42665), .CP(clk), .Q(n69201) );
  dff_sg \shifter_0/ow_14_reg[11]  ( .D(n42666), .CP(clk), .Q(n69200) );
  dff_sg \shifter_0/ow_14_reg[12]  ( .D(n42674), .CP(clk), .Q(n69199) );
  dff_sg \shifter_0/ow_14_reg[13]  ( .D(n42675), .CP(clk), .Q(n69198) );
  dff_sg \shifter_0/ow_14_reg[14]  ( .D(n42671), .CP(clk), .Q(n69197) );
  dff_sg \shifter_0/ow_14_reg[15]  ( .D(n42672), .CP(clk), .Q(n69196) );
  dff_sg \shifter_0/ow_14_reg[16]  ( .D(n42704), .CP(clk), .Q(n69195) );
  dff_sg \shifter_0/ow_14_reg[17]  ( .D(n42705), .CP(clk), .Q(n69194) );
  dff_sg \shifter_0/ow_14_reg[18]  ( .D(n42701), .CP(clk), .Q(n69193) );
  dff_sg \shifter_0/ow_14_reg[19]  ( .D(n42702), .CP(clk), .Q(n69192) );
  dff_sg \shifter_0/ow_13_reg[0]  ( .D(n42710), .CP(clk), .Q(n69191) );
  dff_sg \shifter_0/ow_13_reg[1]  ( .D(n42711), .CP(clk), .Q(n69190) );
  dff_sg \shifter_0/ow_13_reg[2]  ( .D(n42707), .CP(clk), .Q(n69189) );
  dff_sg \shifter_0/ow_13_reg[3]  ( .D(n42708), .CP(clk), .Q(n69188) );
  dff_sg \shifter_0/ow_13_reg[4]  ( .D(n42692), .CP(clk), .Q(n69187) );
  dff_sg \shifter_0/ow_13_reg[5]  ( .D(n42693), .CP(clk), .Q(n69186) );
  dff_sg \shifter_0/ow_13_reg[6]  ( .D(n42689), .CP(clk), .Q(n69185) );
  dff_sg \shifter_0/ow_13_reg[7]  ( .D(n42690), .CP(clk), .Q(n69184) );
  dff_sg \shifter_0/ow_13_reg[8]  ( .D(n42698), .CP(clk), .Q(n69183) );
  dff_sg \shifter_0/ow_13_reg[9]  ( .D(n42699), .CP(clk), .Q(n69182) );
  dff_sg \shifter_0/ow_13_reg[10]  ( .D(n42695), .CP(clk), .Q(n69181) );
  dff_sg \shifter_0/ow_13_reg[11]  ( .D(n42696), .CP(clk), .Q(n69180) );
  dff_sg \shifter_0/ow_13_reg[12]  ( .D(n42632), .CP(clk), .Q(n69179) );
  dff_sg \shifter_0/ow_13_reg[13]  ( .D(n42633), .CP(clk), .Q(n69178) );
  dff_sg \shifter_0/ow_13_reg[14]  ( .D(n42629), .CP(clk), .Q(n69177) );
  dff_sg \shifter_0/ow_13_reg[15]  ( .D(n42630), .CP(clk), .Q(n69176) );
  dff_sg \shifter_0/ow_13_reg[16]  ( .D(n42638), .CP(clk), .Q(n69175) );
  dff_sg \shifter_0/ow_13_reg[17]  ( .D(n42639), .CP(clk), .Q(n69174) );
  dff_sg \shifter_0/ow_13_reg[18]  ( .D(n42635), .CP(clk), .Q(n69173) );
  dff_sg \shifter_0/ow_13_reg[19]  ( .D(n42636), .CP(clk), .Q(n69172) );
  dff_sg \shifter_0/ow_12_reg[0]  ( .D(n42620), .CP(clk), .Q(n69171) );
  dff_sg \shifter_0/ow_12_reg[1]  ( .D(n42621), .CP(clk), .Q(n69170) );
  dff_sg \shifter_0/ow_12_reg[2]  ( .D(n42617), .CP(clk), .Q(n69169) );
  dff_sg \shifter_0/ow_12_reg[3]  ( .D(n42618), .CP(clk), .Q(n69168) );
  dff_sg \shifter_0/ow_12_reg[4]  ( .D(n42626), .CP(clk), .Q(n69167) );
  dff_sg \shifter_0/ow_12_reg[5]  ( .D(n42627), .CP(clk), .Q(n69166) );
  dff_sg \shifter_0/ow_12_reg[6]  ( .D(n42623), .CP(clk), .Q(n69165) );
  dff_sg \shifter_0/ow_12_reg[7]  ( .D(n42624), .CP(clk), .Q(n69164) );
  dff_sg \shifter_0/ow_12_reg[8]  ( .D(n42656), .CP(clk), .Q(n69163) );
  dff_sg \shifter_0/ow_12_reg[9]  ( .D(n42657), .CP(clk), .Q(n69162) );
  dff_sg \shifter_0/ow_12_reg[10]  ( .D(n42653), .CP(clk), .Q(n69161) );
  dff_sg \shifter_0/ow_12_reg[11]  ( .D(n42654), .CP(clk), .Q(n69160) );
  dff_sg \shifter_0/ow_12_reg[12]  ( .D(n42662), .CP(clk), .Q(n69159) );
  dff_sg \shifter_0/ow_12_reg[13]  ( .D(n42663), .CP(clk), .Q(n69158) );
  dff_sg \shifter_0/ow_12_reg[14]  ( .D(n42659), .CP(clk), .Q(n69157) );
  dff_sg \shifter_0/ow_12_reg[15]  ( .D(n42660), .CP(clk), .Q(n69156) );
  dff_sg \shifter_0/ow_12_reg[16]  ( .D(n42644), .CP(clk), .Q(n69155) );
  dff_sg \shifter_0/ow_12_reg[17]  ( .D(n42645), .CP(clk), .Q(n69154) );
  dff_sg \shifter_0/ow_12_reg[18]  ( .D(n42641), .CP(clk), .Q(n69153) );
  dff_sg \shifter_0/ow_12_reg[19]  ( .D(n42642), .CP(clk), .Q(n69152) );
  dff_sg \shifter_0/ow_11_reg[0]  ( .D(n42650), .CP(clk), .Q(n69151) );
  dff_sg \shifter_0/ow_11_reg[1]  ( .D(n42651), .CP(clk), .Q(n69150) );
  dff_sg \shifter_0/ow_11_reg[2]  ( .D(n42647), .CP(clk), .Q(n69149) );
  dff_sg \shifter_0/ow_11_reg[3]  ( .D(n42648), .CP(clk), .Q(n69148) );
  dff_sg \shifter_0/ow_11_reg[4]  ( .D(n42776), .CP(clk), .Q(n69147) );
  dff_sg \shifter_0/ow_11_reg[5]  ( .D(n42777), .CP(clk), .Q(n69146) );
  dff_sg \shifter_0/ow_11_reg[6]  ( .D(n42773), .CP(clk), .Q(n69145) );
  dff_sg \shifter_0/ow_11_reg[7]  ( .D(n42774), .CP(clk), .Q(n69144) );
  dff_sg \shifter_0/ow_11_reg[8]  ( .D(n42782), .CP(clk), .Q(n69143) );
  dff_sg \shifter_0/ow_11_reg[9]  ( .D(n42783), .CP(clk), .Q(n69142) );
  dff_sg \shifter_0/ow_11_reg[10]  ( .D(n42779), .CP(clk), .Q(n69141) );
  dff_sg \shifter_0/ow_11_reg[11]  ( .D(n42780), .CP(clk), .Q(n69140) );
  dff_sg \shifter_0/ow_11_reg[12]  ( .D(n42764), .CP(clk), .Q(n69139) );
  dff_sg \shifter_0/ow_11_reg[13]  ( .D(n42765), .CP(clk), .Q(n69138) );
  dff_sg \shifter_0/ow_11_reg[14]  ( .D(n42761), .CP(clk), .Q(n69137) );
  dff_sg \shifter_0/ow_11_reg[15]  ( .D(n42762), .CP(clk), .Q(n69136) );
  dff_sg \shifter_0/ow_11_reg[16]  ( .D(n42770), .CP(clk), .Q(n69135) );
  dff_sg \shifter_0/ow_11_reg[17]  ( .D(n42771), .CP(clk), .Q(n69134) );
  dff_sg \shifter_0/ow_11_reg[18]  ( .D(n42767), .CP(clk), .Q(n69133) );
  dff_sg \shifter_0/ow_11_reg[19]  ( .D(n42768), .CP(clk), .Q(n69132) );
  dff_sg \shifter_0/ow_10_reg[0]  ( .D(n42793), .CP(clk), .Q(n69131) );
  dff_sg \shifter_0/ow_10_reg[1]  ( .D(n42794), .CP(clk), .Q(n69130) );
  dff_sg \shifter_0/ow_10_reg[2]  ( .D(n42791), .CP(clk), .Q(n69129) );
  dff_sg \shifter_0/ow_10_reg[3]  ( .D(n42792), .CP(clk), .Q(n69128) );
  dff_sg \shifter_0/ow_10_reg[4]  ( .D(n42799), .CP(clk), .Q(n69127) );
  dff_sg \shifter_0/ow_10_reg[5]  ( .D(n42800), .CP(clk), .Q(n69126) );
  dff_sg \shifter_0/ow_10_reg[6]  ( .D(n42798), .CP(clk), .Q(n69125) );
  dff_sg \shifter_0/ow_10_reg[7]  ( .D(n42790), .CP(clk), .Q(n69124) );
  dff_sg \shifter_0/ow_10_reg[8]  ( .D(n42788), .CP(clk), .Q(n69123) );
  dff_sg \shifter_0/ow_10_reg[9]  ( .D(n42789), .CP(clk), .Q(n69122) );
  dff_sg \shifter_0/ow_10_reg[10]  ( .D(n42785), .CP(clk), .Q(n69121) );
  dff_sg \shifter_0/ow_10_reg[11]  ( .D(n42786), .CP(clk), .Q(n69120) );
  dff_sg \shifter_0/ow_10_reg[12]  ( .D(n42796), .CP(clk), .Q(n69119) );
  dff_sg \shifter_0/ow_10_reg[13]  ( .D(n42797), .CP(clk), .Q(n69118) );
  dff_sg \shifter_0/ow_10_reg[14]  ( .D(n42431), .CP(clk), .Q(n69117) );
  dff_sg \shifter_0/ow_10_reg[15]  ( .D(n42432), .CP(clk), .Q(n69116) );
  dff_sg \shifter_0/ow_10_reg[16]  ( .D(n42728), .CP(clk), .Q(n69115) );
  dff_sg \shifter_0/ow_10_reg[17]  ( .D(n42729), .CP(clk), .Q(n69114) );
  dff_sg \shifter_0/ow_10_reg[18]  ( .D(n42725), .CP(clk), .Q(n69113) );
  dff_sg \shifter_0/ow_10_reg[19]  ( .D(n42726), .CP(clk), .Q(n69112) );
  dff_sg \shifter_0/ow_9_reg[0]  ( .D(n42734), .CP(clk), .Q(n69111) );
  dff_sg \shifter_0/ow_9_reg[1]  ( .D(n42735), .CP(clk), .Q(n69110) );
  dff_sg \shifter_0/ow_9_reg[2]  ( .D(n42731), .CP(clk), .Q(n69109) );
  dff_sg \shifter_0/ow_9_reg[3]  ( .D(n42732), .CP(clk), .Q(n69108) );
  dff_sg \shifter_0/ow_9_reg[4]  ( .D(n42716), .CP(clk), .Q(n69107) );
  dff_sg \shifter_0/ow_9_reg[5]  ( .D(n42717), .CP(clk), .Q(n69106) );
  dff_sg \shifter_0/ow_9_reg[6]  ( .D(n42713), .CP(clk), .Q(n69105) );
  dff_sg \shifter_0/ow_9_reg[7]  ( .D(n42714), .CP(clk), .Q(n69104) );
  dff_sg \shifter_0/ow_9_reg[8]  ( .D(n42722), .CP(clk), .Q(n69103) );
  dff_sg \shifter_0/ow_9_reg[9]  ( .D(n42723), .CP(clk), .Q(n69102) );
  dff_sg \shifter_0/ow_9_reg[10]  ( .D(n42719), .CP(clk), .Q(n69101) );
  dff_sg \shifter_0/ow_9_reg[11]  ( .D(n42720), .CP(clk), .Q(n69100) );
  dff_sg \shifter_0/ow_9_reg[12]  ( .D(n42752), .CP(clk), .Q(n69099) );
  dff_sg \shifter_0/ow_9_reg[13]  ( .D(n42753), .CP(clk), .Q(n69098) );
  dff_sg \shifter_0/ow_9_reg[14]  ( .D(n42749), .CP(clk), .Q(n69097) );
  dff_sg \shifter_0/ow_9_reg[15]  ( .D(n42750), .CP(clk), .Q(n69096) );
  dff_sg \shifter_0/ow_9_reg[16]  ( .D(n42758), .CP(clk), .Q(n69095) );
  dff_sg \shifter_0/ow_9_reg[17]  ( .D(n42759), .CP(clk), .Q(n69094) );
  dff_sg \shifter_0/ow_9_reg[18]  ( .D(n42755), .CP(clk), .Q(n69093) );
  dff_sg \shifter_0/ow_9_reg[19]  ( .D(n42756), .CP(clk), .Q(n69092) );
  dff_sg \shifter_0/ow_8_reg[0]  ( .D(n42740), .CP(clk), .Q(n69091) );
  dff_sg \shifter_0/ow_8_reg[1]  ( .D(n42741), .CP(clk), .Q(n69090) );
  dff_sg \shifter_0/ow_8_reg[2]  ( .D(n42737), .CP(clk), .Q(n69089) );
  dff_sg \shifter_0/ow_8_reg[3]  ( .D(n42738), .CP(clk), .Q(n69088) );
  dff_sg \shifter_0/ow_8_reg[4]  ( .D(n42746), .CP(clk), .Q(n69087) );
  dff_sg \shifter_0/ow_8_reg[5]  ( .D(n42747), .CP(clk), .Q(n69086) );
  dff_sg \shifter_0/ow_8_reg[6]  ( .D(n42743), .CP(clk), .Q(n69085) );
  dff_sg \shifter_0/ow_8_reg[7]  ( .D(n42744), .CP(clk), .Q(n69084) );
  dff_sg \shifter_0/ow_8_reg[8]  ( .D(n42488), .CP(clk), .Q(n69083) );
  dff_sg \shifter_0/ow_8_reg[9]  ( .D(n42489), .CP(clk), .Q(n69082) );
  dff_sg \shifter_0/ow_8_reg[10]  ( .D(n42485), .CP(clk), .Q(n69081) );
  dff_sg \shifter_0/ow_8_reg[11]  ( .D(n42486), .CP(clk), .Q(n69080) );
  dff_sg \shifter_0/ow_8_reg[12]  ( .D(n42494), .CP(clk), .Q(n69079) );
  dff_sg \shifter_0/ow_8_reg[13]  ( .D(n42495), .CP(clk), .Q(n69078) );
  dff_sg \shifter_0/ow_8_reg[14]  ( .D(n42491), .CP(clk), .Q(n69077) );
  dff_sg \shifter_0/ow_8_reg[15]  ( .D(n42492), .CP(clk), .Q(n69076) );
  dff_sg \shifter_0/ow_8_reg[16]  ( .D(n42476), .CP(clk), .Q(n69075) );
  dff_sg \shifter_0/ow_8_reg[17]  ( .D(n42477), .CP(clk), .Q(n69074) );
  dff_sg \shifter_0/ow_8_reg[18]  ( .D(n42473), .CP(clk), .Q(n69073) );
  dff_sg \shifter_0/ow_8_reg[19]  ( .D(n42474), .CP(clk), .Q(n69072) );
  dff_sg \shifter_0/ow_7_reg[0]  ( .D(n42482), .CP(clk), .Q(n69071) );
  dff_sg \shifter_0/ow_7_reg[1]  ( .D(n42483), .CP(clk), .Q(n69070) );
  dff_sg \shifter_0/ow_7_reg[2]  ( .D(n42479), .CP(clk), .Q(n69069) );
  dff_sg \shifter_0/ow_7_reg[3]  ( .D(n42480), .CP(clk), .Q(n69068) );
  dff_sg \shifter_0/ow_7_reg[4]  ( .D(n42512), .CP(clk), .Q(n69067) );
  dff_sg \shifter_0/ow_7_reg[5]  ( .D(n42513), .CP(clk), .Q(n69066) );
  dff_sg \shifter_0/ow_7_reg[6]  ( .D(n42509), .CP(clk), .Q(n69065) );
  dff_sg \shifter_0/ow_7_reg[7]  ( .D(n42510), .CP(clk), .Q(n69064) );
  dff_sg \shifter_0/ow_7_reg[8]  ( .D(n42518), .CP(clk), .Q(n69063) );
  dff_sg \shifter_0/ow_7_reg[9]  ( .D(n42519), .CP(clk), .Q(n69062) );
  dff_sg \shifter_0/ow_7_reg[10]  ( .D(n42515), .CP(clk), .Q(n69061) );
  dff_sg \shifter_0/ow_7_reg[11]  ( .D(n42516), .CP(clk), .Q(n69060) );
  dff_sg \shifter_0/ow_7_reg[12]  ( .D(n42500), .CP(clk), .Q(n69059) );
  dff_sg \shifter_0/ow_7_reg[13]  ( .D(n42501), .CP(clk), .Q(n69058) );
  dff_sg \shifter_0/ow_7_reg[14]  ( .D(n42497), .CP(clk), .Q(n69057) );
  dff_sg \shifter_0/ow_7_reg[15]  ( .D(n42498), .CP(clk), .Q(n69056) );
  dff_sg \shifter_0/ow_7_reg[16]  ( .D(n42506), .CP(clk), .Q(n69055) );
  dff_sg \shifter_0/ow_7_reg[17]  ( .D(n42507), .CP(clk), .Q(n69054) );
  dff_sg \shifter_0/ow_7_reg[18]  ( .D(n42503), .CP(clk), .Q(n69053) );
  dff_sg \shifter_0/ow_7_reg[19]  ( .D(n42504), .CP(clk), .Q(n69052) );
  dff_sg \shifter_0/ow_6_reg[0]  ( .D(n42440), .CP(clk), .Q(n69051) );
  dff_sg \shifter_0/ow_6_reg[1]  ( .D(n42441), .CP(clk), .Q(n69050) );
  dff_sg \shifter_0/ow_6_reg[2]  ( .D(n42437), .CP(clk), .Q(n69049) );
  dff_sg \shifter_0/ow_6_reg[3]  ( .D(n42438), .CP(clk), .Q(n69048) );
  dff_sg \shifter_0/ow_6_reg[4]  ( .D(n42446), .CP(clk), .Q(n69047) );
  dff_sg \shifter_0/ow_6_reg[5]  ( .D(n42447), .CP(clk), .Q(n69046) );
  dff_sg \shifter_0/ow_6_reg[6]  ( .D(n42443), .CP(clk), .Q(n69045) );
  dff_sg \shifter_0/ow_6_reg[7]  ( .D(n42444), .CP(clk), .Q(n69044) );
  dff_sg \shifter_0/ow_6_reg[8]  ( .D(n42428), .CP(clk), .Q(n69043) );
  dff_sg \shifter_0/ow_6_reg[9]  ( .D(n42429), .CP(clk), .Q(n69042) );
  dff_sg \shifter_0/ow_6_reg[10]  ( .D(n42425), .CP(clk), .Q(n69041) );
  dff_sg \shifter_0/ow_6_reg[11]  ( .D(n42426), .CP(clk), .Q(n69040) );
  dff_sg \shifter_0/ow_6_reg[12]  ( .D(n42430), .CP(clk), .Q(n69039) );
  dff_sg \shifter_0/ow_6_reg[13]  ( .D(n42795), .CP(clk), .Q(n69038) );
  dff_sg \shifter_0/ow_6_reg[14]  ( .D(n42434), .CP(clk), .Q(n69037) );
  dff_sg \shifter_0/ow_6_reg[15]  ( .D(n42435), .CP(clk), .Q(n69036) );
  dff_sg \shifter_0/ow_6_reg[16]  ( .D(n42464), .CP(clk), .Q(n69035) );
  dff_sg \shifter_0/ow_6_reg[17]  ( .D(n42465), .CP(clk), .Q(n69034) );
  dff_sg \shifter_0/ow_6_reg[18]  ( .D(n42461), .CP(clk), .Q(n69033) );
  dff_sg \shifter_0/ow_6_reg[19]  ( .D(n42462), .CP(clk), .Q(n69032) );
  dff_sg \shifter_0/ow_5_reg[0]  ( .D(n42470), .CP(clk), .Q(n69031) );
  dff_sg \shifter_0/ow_5_reg[1]  ( .D(n42471), .CP(clk), .Q(n69030) );
  dff_sg \shifter_0/ow_5_reg[2]  ( .D(n42467), .CP(clk), .Q(n69029) );
  dff_sg \shifter_0/ow_5_reg[3]  ( .D(n42468), .CP(clk), .Q(n69028) );
  dff_sg \shifter_0/ow_5_reg[4]  ( .D(n42452), .CP(clk), .Q(n69027) );
  dff_sg \shifter_0/ow_5_reg[5]  ( .D(n42453), .CP(clk), .Q(n69026) );
  dff_sg \shifter_0/ow_5_reg[6]  ( .D(n42449), .CP(clk), .Q(n69025) );
  dff_sg \shifter_0/ow_5_reg[7]  ( .D(n42450), .CP(clk), .Q(n69024) );
  dff_sg \shifter_0/ow_5_reg[8]  ( .D(n42458), .CP(clk), .Q(n69023) );
  dff_sg \shifter_0/ow_5_reg[9]  ( .D(n42459), .CP(clk), .Q(n69022) );
  dff_sg \shifter_0/ow_5_reg[10]  ( .D(n42455), .CP(clk), .Q(n69021) );
  dff_sg \shifter_0/ow_5_reg[11]  ( .D(n42456), .CP(clk), .Q(n69020) );
  dff_sg \shifter_0/ow_5_reg[12]  ( .D(n42584), .CP(clk), .Q(n69019) );
  dff_sg \shifter_0/ow_5_reg[13]  ( .D(n42585), .CP(clk), .Q(n69018) );
  dff_sg \shifter_0/ow_5_reg[14]  ( .D(n42581), .CP(clk), .Q(n69017) );
  dff_sg \shifter_0/ow_5_reg[15]  ( .D(n42582), .CP(clk), .Q(n69016) );
  dff_sg \shifter_0/ow_5_reg[16]  ( .D(n42590), .CP(clk), .Q(n69015) );
  dff_sg \shifter_0/ow_5_reg[17]  ( .D(n42591), .CP(clk), .Q(n69014) );
  dff_sg \shifter_0/ow_5_reg[18]  ( .D(n42587), .CP(clk), .Q(n69013) );
  dff_sg \shifter_0/ow_5_reg[19]  ( .D(n42588), .CP(clk), .Q(n69012) );
  dff_sg \shifter_0/ow_4_reg[0]  ( .D(n42572), .CP(clk), .Q(n69011) );
  dff_sg \shifter_0/ow_4_reg[1]  ( .D(n42573), .CP(clk), .Q(n69010) );
  dff_sg \shifter_0/ow_4_reg[2]  ( .D(n42569), .CP(clk), .Q(n69009) );
  dff_sg \shifter_0/ow_4_reg[3]  ( .D(n42570), .CP(clk), .Q(n69008) );
  dff_sg \shifter_0/ow_4_reg[4]  ( .D(n42578), .CP(clk), .Q(n69007) );
  dff_sg \shifter_0/ow_4_reg[5]  ( .D(n42579), .CP(clk), .Q(n69006) );
  dff_sg \shifter_0/ow_4_reg[6]  ( .D(n42575), .CP(clk), .Q(n69005) );
  dff_sg \shifter_0/ow_4_reg[7]  ( .D(n42576), .CP(clk), .Q(n69004) );
  dff_sg \shifter_0/ow_4_reg[8]  ( .D(n42608), .CP(clk), .Q(n69003) );
  dff_sg \shifter_0/ow_4_reg[9]  ( .D(n42609), .CP(clk), .Q(n69002) );
  dff_sg \shifter_0/ow_4_reg[10]  ( .D(n42605), .CP(clk), .Q(n69001) );
  dff_sg \shifter_0/ow_4_reg[11]  ( .D(n42606), .CP(clk), .Q(n69000) );
  dff_sg \shifter_0/ow_4_reg[12]  ( .D(n42614), .CP(clk), .Q(n68999) );
  dff_sg \shifter_0/ow_4_reg[13]  ( .D(n42615), .CP(clk), .Q(n68998) );
  dff_sg \shifter_0/ow_4_reg[14]  ( .D(n42611), .CP(clk), .Q(n68997) );
  dff_sg \shifter_0/ow_4_reg[15]  ( .D(n42612), .CP(clk), .Q(n68996) );
  dff_sg \shifter_0/ow_4_reg[16]  ( .D(n42596), .CP(clk), .Q(n68995) );
  dff_sg \shifter_0/ow_4_reg[17]  ( .D(n42597), .CP(clk), .Q(n68994) );
  dff_sg \shifter_0/ow_4_reg[18]  ( .D(n42593), .CP(clk), .Q(n68993) );
  dff_sg \shifter_0/ow_4_reg[19]  ( .D(n42594), .CP(clk), .Q(n68992) );
  dff_sg \shifter_0/ow_3_reg[0]  ( .D(n42602), .CP(clk), .Q(n68991) );
  dff_sg \shifter_0/ow_3_reg[1]  ( .D(n42603), .CP(clk), .Q(n68990) );
  dff_sg \shifter_0/ow_3_reg[2]  ( .D(n42599), .CP(clk), .Q(n68989) );
  dff_sg \shifter_0/ow_3_reg[3]  ( .D(n42600), .CP(clk), .Q(n68988) );
  dff_sg \shifter_0/ow_3_reg[4]  ( .D(n42536), .CP(clk), .Q(n68987) );
  dff_sg \shifter_0/ow_3_reg[5]  ( .D(n42537), .CP(clk), .Q(n68986) );
  dff_sg \shifter_0/ow_3_reg[6]  ( .D(n42533), .CP(clk), .Q(n68985) );
  dff_sg \shifter_0/ow_3_reg[7]  ( .D(n42534), .CP(clk), .Q(n68984) );
  dff_sg \shifter_0/ow_3_reg[8]  ( .D(n42542), .CP(clk), .Q(n68983) );
  dff_sg \shifter_0/ow_3_reg[9]  ( .D(n42543), .CP(clk), .Q(n68982) );
  dff_sg \shifter_0/ow_3_reg[10]  ( .D(n42539), .CP(clk), .Q(n68981) );
  dff_sg \shifter_0/ow_3_reg[11]  ( .D(n42540), .CP(clk), .Q(n68980) );
  dff_sg \shifter_0/ow_3_reg[12]  ( .D(n42524), .CP(clk), .Q(n68979) );
  dff_sg \shifter_0/ow_3_reg[13]  ( .D(n42525), .CP(clk), .Q(n68978) );
  dff_sg \shifter_0/ow_3_reg[14]  ( .D(n42521), .CP(clk), .Q(n68977) );
  dff_sg \shifter_0/ow_3_reg[15]  ( .D(n42522), .CP(clk), .Q(n68976) );
  dff_sg \shifter_0/ow_3_reg[16]  ( .D(n42530), .CP(clk), .Q(n68975) );
  dff_sg \shifter_0/ow_3_reg[17]  ( .D(n42531), .CP(clk), .Q(n68974) );
  dff_sg \shifter_0/ow_3_reg[18]  ( .D(n42527), .CP(clk), .Q(n68973) );
  dff_sg \shifter_0/ow_3_reg[19]  ( .D(n42528), .CP(clk), .Q(n68972) );
  dff_sg \shifter_0/ow_2_reg[0]  ( .D(n42560), .CP(clk), .Q(n68971) );
  dff_sg \shifter_0/ow_2_reg[1]  ( .D(n42561), .CP(clk), .Q(n68970) );
  dff_sg \shifter_0/ow_2_reg[2]  ( .D(n42557), .CP(clk), .Q(n68969) );
  dff_sg \shifter_0/ow_2_reg[3]  ( .D(n42558), .CP(clk), .Q(n68968) );
  dff_sg \shifter_0/ow_2_reg[4]  ( .D(n42566), .CP(clk), .Q(n68967) );
  dff_sg \shifter_0/ow_2_reg[5]  ( .D(n42567), .CP(clk), .Q(n68966) );
  dff_sg \shifter_0/ow_2_reg[6]  ( .D(n42563), .CP(clk), .Q(n68965) );
  dff_sg \shifter_0/ow_2_reg[7]  ( .D(n42564), .CP(clk), .Q(n68964) );
  dff_sg \shifter_0/ow_2_reg[8]  ( .D(n42548), .CP(clk), .Q(n68963) );
  dff_sg \shifter_0/ow_2_reg[9]  ( .D(n42549), .CP(clk), .Q(n68962) );
  dff_sg \shifter_0/ow_2_reg[10]  ( .D(n42545), .CP(clk), .Q(n68961) );
  dff_sg \shifter_0/ow_2_reg[11]  ( .D(n42546), .CP(clk), .Q(n68960) );
  dff_sg \shifter_0/ow_2_reg[12]  ( .D(n42554), .CP(clk), .Q(n68959) );
  dff_sg \shifter_0/ow_2_reg[13]  ( .D(n42555), .CP(clk), .Q(n68958) );
  dff_sg \shifter_0/ow_2_reg[14]  ( .D(n42551), .CP(clk), .Q(n68957) );
  dff_sg \shifter_0/ow_2_reg[15]  ( .D(n42552), .CP(clk), .Q(n68956) );
  dff_sg \shifter_0/ow_2_reg[16]  ( .D(n42389), .CP(clk), .Q(n68955) );
  dff_sg \shifter_0/ow_2_reg[17]  ( .D(n42392), .CP(clk), .Q(n68954) );
  dff_sg \shifter_0/ow_2_reg[18]  ( .D(n42532), .CP(clk), .Q(n68953) );
  dff_sg \shifter_0/ow_2_reg[19]  ( .D(n42408), .CP(clk), .Q(n68952) );
  dff_sg \shifter_0/ow_1_reg[0]  ( .D(n42374), .CP(clk), .Q(n68951) );
  dff_sg \shifter_0/ow_1_reg[1]  ( .D(n42377), .CP(clk), .Q(n68950) );
  dff_sg \shifter_0/ow_1_reg[2]  ( .D(n42380), .CP(clk), .Q(n68949) );
  dff_sg \shifter_0/ow_1_reg[3]  ( .D(n42383), .CP(clk), .Q(n68948) );
  dff_sg \shifter_0/ow_1_reg[4]  ( .D(n42168), .CP(clk), .Q(n68947) );
  dff_sg \shifter_0/ow_1_reg[5]  ( .D(n42171), .CP(clk), .Q(n68946) );
  dff_sg \shifter_0/ow_1_reg[6]  ( .D(n42201), .CP(clk), .Q(n68945) );
  dff_sg \shifter_0/ow_1_reg[7]  ( .D(n42237), .CP(clk), .Q(n68944) );
  dff_sg \shifter_0/ow_1_reg[8]  ( .D(n42538), .CP(clk), .Q(n68943) );
  dff_sg \shifter_0/ow_1_reg[9]  ( .D(n42365), .CP(clk), .Q(n68942) );
  dff_sg \shifter_0/ow_1_reg[10]  ( .D(n42395), .CP(clk), .Q(n68941) );
  dff_sg \shifter_0/ow_1_reg[11]  ( .D(n42398), .CP(clk), .Q(n68940) );
  dff_sg \shifter_0/ow_1_reg[12]  ( .D(n42727), .CP(clk), .Q(n68939) );
  dff_sg \shifter_0/ow_1_reg[13]  ( .D(n42730), .CP(clk), .Q(n68938) );
  dff_sg \shifter_0/ow_1_reg[14]  ( .D(n42407), .CP(clk), .Q(n68937) );
  dff_sg \shifter_0/ow_1_reg[15]  ( .D(n42422), .CP(clk), .Q(n68936) );
  dff_sg \shifter_0/ow_1_reg[16]  ( .D(n42706), .CP(clk), .Q(n68935) );
  dff_sg \shifter_0/ow_1_reg[17]  ( .D(n42709), .CP(clk), .Q(n68934) );
  dff_sg \shifter_0/ow_1_reg[18]  ( .D(n42418), .CP(clk), .Q(n68933) );
  dff_sg \shifter_0/ow_1_reg[19]  ( .D(n42712), .CP(clk), .Q(n68932) );
  dff_sg \shifter_0/ow_0_reg[0]  ( .D(n42404), .CP(clk), .Q(n68931) );
  dff_sg \shifter_0/ow_0_reg[1]  ( .D(n42350), .CP(clk), .Q(n68930) );
  dff_sg \shifter_0/ow_0_reg[2]  ( .D(n42420), .CP(clk), .Q(n68929) );
  dff_sg \shifter_0/ow_0_reg[3]  ( .D(n42356), .CP(clk), .Q(n68928) );
  dff_sg \shifter_0/ow_0_reg[4]  ( .D(n42401), .CP(clk), .Q(n68927) );
  dff_sg \shifter_0/ow_0_reg[5]  ( .D(n42338), .CP(clk), .Q(n68926) );
  dff_sg \shifter_0/ow_0_reg[6]  ( .D(n42347), .CP(clk), .Q(n68925) );
  dff_sg \shifter_0/ow_0_reg[7]  ( .D(n42353), .CP(clk), .Q(n68924) );
  dff_sg \shifter_0/ow_0_reg[8]  ( .D(n42222), .CP(clk), .Q(n68923) );
  dff_sg \shifter_0/ow_0_reg[9]  ( .D(n42754), .CP(clk), .Q(n68922) );
  dff_sg \shifter_0/ow_0_reg[10]  ( .D(n42745), .CP(clk), .Q(n68921) );
  dff_sg \shifter_0/ow_0_reg[11]  ( .D(n42161), .CP(clk), .Q(n68920) );
  dff_sg \shifter_0/ow_0_reg[12]  ( .D(n42204), .CP(clk), .Q(n68919) );
  dff_sg \shifter_0/ow_0_reg[13]  ( .D(n42207), .CP(clk), .Q(n68918) );
  dff_sg \shifter_0/ow_0_reg[14]  ( .D(n42210), .CP(clk), .Q(n68917) );
  dff_sg \shifter_0/ow_0_reg[15]  ( .D(n42213), .CP(clk), .Q(n68916) );
  dff_sg \shifter_0/ow_0_reg[16]  ( .D(n42697), .CP(clk), .Q(n68915) );
  dff_sg \shifter_0/ow_0_reg[17]  ( .D(n42700), .CP(clk), .Q(n68914) );
  dff_sg \shifter_0/ow_0_reg[18]  ( .D(n42180), .CP(clk), .Q(n68913) );
  dff_sg \shifter_0/ow_0_reg[19]  ( .D(n42703), .CP(clk), .Q(n68912) );
  dff_sg \shifter_0/oi_15_reg[0]  ( .D(n42183), .CP(clk), .Q(n68911) );
  dff_sg \shifter_0/oi_15_reg[1]  ( .D(n42186), .CP(clk), .Q(n68910) );
  dff_sg \shifter_0/oi_15_reg[2]  ( .D(n42691), .CP(clk), .Q(n68909) );
  dff_sg \shifter_0/oi_15_reg[3]  ( .D(n42694), .CP(clk), .Q(n68908) );
  dff_sg \shifter_0/oi_15_reg[4]  ( .D(n42225), .CP(clk), .Q(n68907) );
  dff_sg \shifter_0/oi_15_reg[5]  ( .D(n42231), .CP(clk), .Q(n68906) );
  dff_sg \shifter_0/oi_15_reg[6]  ( .D(n42234), .CP(clk), .Q(n68905) );
  dff_sg \shifter_0/oi_15_reg[7]  ( .D(n42240), .CP(clk), .Q(n68904) );
  dff_sg \shifter_0/oi_15_reg[8]  ( .D(n42362), .CP(clk), .Q(n68903) );
  dff_sg \shifter_0/oi_15_reg[9]  ( .D(n42368), .CP(clk), .Q(n68902) );
  dff_sg \shifter_0/oi_15_reg[10]  ( .D(n42415), .CP(clk), .Q(n68901) );
  dff_sg \shifter_0/oi_15_reg[11]  ( .D(n42371), .CP(clk), .Q(n68900) );
  dff_sg \shifter_0/oi_15_reg[12]  ( .D(n42359), .CP(clk), .Q(n68899) );
  dff_sg \shifter_0/oi_15_reg[13]  ( .D(n42416), .CP(clk), .Q(n68898) );
  dff_sg \shifter_0/oi_15_reg[14]  ( .D(n42244), .CP(clk), .Q(n68897) );
  dff_sg \shifter_0/oi_15_reg[15]  ( .D(n42162), .CP(clk), .Q(n68896) );
  dff_sg \shifter_0/oi_15_reg[16]  ( .D(n42195), .CP(clk), .Q(n68895) );
  dff_sg \shifter_0/oi_15_reg[17]  ( .D(n42198), .CP(clk), .Q(n68894) );
  dff_sg \shifter_0/oi_15_reg[18]  ( .D(n42245), .CP(clk), .Q(n68893) );
  dff_sg \shifter_0/oi_15_reg[19]  ( .D(n42216), .CP(clk), .Q(n68892) );
  dff_sg \shifter_0/oi_14_reg[0]  ( .D(n42220), .CP(clk), .Q(n68891) );
  dff_sg \shifter_0/oi_14_reg[1]  ( .D(n42221), .CP(clk), .Q(n68890) );
  dff_sg \shifter_0/oi_14_reg[2]  ( .D(n42217), .CP(clk), .Q(n68889) );
  dff_sg \shifter_0/oi_14_reg[3]  ( .D(n42218), .CP(clk), .Q(n68888) );
  dff_sg \shifter_0/oi_14_reg[4]  ( .D(n42226), .CP(clk), .Q(n68887) );
  dff_sg \shifter_0/oi_14_reg[5]  ( .D(n42227), .CP(clk), .Q(n68886) );
  dff_sg \shifter_0/oi_14_reg[6]  ( .D(n42223), .CP(clk), .Q(n68885) );
  dff_sg \shifter_0/oi_14_reg[7]  ( .D(n42224), .CP(clk), .Q(n68884) );
  dff_sg \shifter_0/oi_14_reg[8]  ( .D(n42208), .CP(clk), .Q(n68883) );
  dff_sg \shifter_0/oi_14_reg[9]  ( .D(n42209), .CP(clk), .Q(n68882) );
  dff_sg \shifter_0/oi_14_reg[10]  ( .D(n42205), .CP(clk), .Q(n68881) );
  dff_sg \shifter_0/oi_14_reg[11]  ( .D(n42206), .CP(clk), .Q(n68880) );
  dff_sg \shifter_0/oi_14_reg[12]  ( .D(n42214), .CP(clk), .Q(n68879) );
  dff_sg \shifter_0/oi_14_reg[13]  ( .D(n42215), .CP(clk), .Q(n68878) );
  dff_sg \shifter_0/oi_14_reg[14]  ( .D(n42211), .CP(clk), .Q(n68877) );
  dff_sg \shifter_0/oi_14_reg[15]  ( .D(n42212), .CP(clk), .Q(n68876) );
  dff_sg \shifter_0/oi_14_reg[16]  ( .D(n42748), .CP(clk), .Q(n68875) );
  dff_sg \shifter_0/oi_14_reg[17]  ( .D(n42751), .CP(clk), .Q(n68874) );
  dff_sg \shifter_0/oi_14_reg[18]  ( .D(n42760), .CP(clk), .Q(n68873) );
  dff_sg \shifter_0/oi_14_reg[19]  ( .D(n42763), .CP(clk), .Q(n68872) );
  dff_sg \shifter_0/oi_13_reg[0]  ( .D(n42733), .CP(clk), .Q(n68871) );
  dff_sg \shifter_0/oi_13_reg[1]  ( .D(n42736), .CP(clk), .Q(n68870) );
  dff_sg \shifter_0/oi_13_reg[2]  ( .D(n42757), .CP(clk), .Q(n68869) );
  dff_sg \shifter_0/oi_13_reg[3]  ( .D(n42739), .CP(clk), .Q(n68868) );
  dff_sg \shifter_0/oi_13_reg[4]  ( .D(n42235), .CP(clk), .Q(n68867) );
  dff_sg \shifter_0/oi_13_reg[5]  ( .D(n42236), .CP(clk), .Q(n68866) );
  dff_sg \shifter_0/oi_13_reg[6]  ( .D(n42232), .CP(clk), .Q(n68865) );
  dff_sg \shifter_0/oi_13_reg[7]  ( .D(n42233), .CP(clk), .Q(n68864) );
  dff_sg \shifter_0/oi_13_reg[8]  ( .D(n42241), .CP(clk), .Q(n68863) );
  dff_sg \shifter_0/oi_13_reg[9]  ( .D(n42242), .CP(clk), .Q(n68862) );
  dff_sg \shifter_0/oi_13_reg[10]  ( .D(n42238), .CP(clk), .Q(n68861) );
  dff_sg \shifter_0/oi_13_reg[11]  ( .D(n42239), .CP(clk), .Q(n68860) );
  dff_sg \shifter_0/oi_13_reg[12]  ( .D(n42172), .CP(clk), .Q(n68859) );
  dff_sg \shifter_0/oi_13_reg[13]  ( .D(n42173), .CP(clk), .Q(n68858) );
  dff_sg \shifter_0/oi_13_reg[14]  ( .D(n42169), .CP(clk), .Q(n68857) );
  dff_sg \shifter_0/oi_13_reg[15]  ( .D(n42170), .CP(clk), .Q(n68856) );
  dff_sg \shifter_0/oi_13_reg[16]  ( .D(n42178), .CP(clk), .Q(n68855) );
  dff_sg \shifter_0/oi_13_reg[17]  ( .D(n42179), .CP(clk), .Q(n68854) );
  dff_sg \shifter_0/oi_13_reg[18]  ( .D(n42175), .CP(clk), .Q(n68853) );
  dff_sg \shifter_0/oi_13_reg[19]  ( .D(n42176), .CP(clk), .Q(n68852) );
  dff_sg \shifter_0/oi_12_reg[0]  ( .D(n42166), .CP(clk), .Q(n68851) );
  dff_sg \shifter_0/oi_12_reg[1]  ( .D(n42167), .CP(clk), .Q(n68850) );
  dff_sg \shifter_0/oi_12_reg[2]  ( .D(n42718), .CP(clk), .Q(n68849) );
  dff_sg \shifter_0/oi_12_reg[3]  ( .D(n42721), .CP(clk), .Q(n68848) );
  dff_sg \shifter_0/oi_12_reg[4]  ( .D(n42252), .CP(clk), .Q(n68847) );
  dff_sg \shifter_0/oi_12_reg[5]  ( .D(n42253), .CP(clk), .Q(n68846) );
  dff_sg \shifter_0/oi_12_reg[6]  ( .D(n42163), .CP(clk), .Q(n68845) );
  dff_sg \shifter_0/oi_12_reg[7]  ( .D(n42164), .CP(clk), .Q(n68844) );
  dff_sg \shifter_0/oi_12_reg[8]  ( .D(n42196), .CP(clk), .Q(n68843) );
  dff_sg \shifter_0/oi_12_reg[9]  ( .D(n42197), .CP(clk), .Q(n68842) );
  dff_sg \shifter_0/oi_12_reg[10]  ( .D(n42193), .CP(clk), .Q(n68841) );
  dff_sg \shifter_0/oi_12_reg[11]  ( .D(n42194), .CP(clk), .Q(n68840) );
  dff_sg \shifter_0/oi_12_reg[12]  ( .D(n42202), .CP(clk), .Q(n68839) );
  dff_sg \shifter_0/oi_12_reg[13]  ( .D(n42203), .CP(clk), .Q(n68838) );
  dff_sg \shifter_0/oi_12_reg[14]  ( .D(n42199), .CP(clk), .Q(n68837) );
  dff_sg \shifter_0/oi_12_reg[15]  ( .D(n42200), .CP(clk), .Q(n68836) );
  dff_sg \shifter_0/oi_12_reg[16]  ( .D(n42184), .CP(clk), .Q(n68835) );
  dff_sg \shifter_0/oi_12_reg[17]  ( .D(n42185), .CP(clk), .Q(n68834) );
  dff_sg \shifter_0/oi_12_reg[18]  ( .D(n42181), .CP(clk), .Q(n68833) );
  dff_sg \shifter_0/oi_12_reg[19]  ( .D(n42182), .CP(clk), .Q(n68832) );
  dff_sg \shifter_0/oi_11_reg[0]  ( .D(n42190), .CP(clk), .Q(n68831) );
  dff_sg \shifter_0/oi_11_reg[1]  ( .D(n42191), .CP(clk), .Q(n68830) );
  dff_sg \shifter_0/oi_11_reg[2]  ( .D(n42187), .CP(clk), .Q(n68829) );
  dff_sg \shifter_0/oi_11_reg[3]  ( .D(n42188), .CP(clk), .Q(n68828) );
  dff_sg \shifter_0/oi_11_reg[4]  ( .D(n42481), .CP(clk), .Q(n68827) );
  dff_sg \shifter_0/oi_11_reg[5]  ( .D(n42478), .CP(clk), .Q(n68826) );
  dff_sg \shifter_0/oi_11_reg[6]  ( .D(n42484), .CP(clk), .Q(n68825) );
  dff_sg \shifter_0/oi_11_reg[7]  ( .D(n42487), .CP(clk), .Q(n68824) );
  dff_sg \shifter_0/oi_11_reg[8]  ( .D(n42529), .CP(clk), .Q(n68823) );
  dff_sg \shifter_0/oi_11_reg[9]  ( .D(n42526), .CP(clk), .Q(n68822) );
  dff_sg \shifter_0/oi_11_reg[10]  ( .D(n42544), .CP(clk), .Q(n68821) );
  dff_sg \shifter_0/oi_11_reg[11]  ( .D(n42547), .CP(clk), .Q(n68820) );
  dff_sg \shifter_0/oi_11_reg[12]  ( .D(n42256), .CP(clk), .Q(n68819) );
  dff_sg \shifter_0/oi_11_reg[13]  ( .D(n42490), .CP(clk), .Q(n68818) );
  dff_sg \shifter_0/oi_11_reg[14]  ( .D(n42255), .CP(clk), .Q(n68817) );
  dff_sg \shifter_0/oi_11_reg[15]  ( .D(n42254), .CP(clk), .Q(n68816) );
  dff_sg \shifter_0/oi_11_reg[16]  ( .D(n42535), .CP(clk), .Q(n68815) );
  dff_sg \shifter_0/oi_11_reg[17]  ( .D(n42523), .CP(clk), .Q(n68814) );
  dff_sg \shifter_0/oi_11_reg[18]  ( .D(n42496), .CP(clk), .Q(n68813) );
  dff_sg \shifter_0/oi_11_reg[19]  ( .D(n42493), .CP(clk), .Q(n68812) );
  dff_sg \shifter_0/oi_10_reg[0]  ( .D(n42559), .CP(clk), .Q(n68811) );
  dff_sg \shifter_0/oi_10_reg[1]  ( .D(n42553), .CP(clk), .Q(n68810) );
  dff_sg \shifter_0/oi_10_reg[2]  ( .D(n42568), .CP(clk), .Q(n68809) );
  dff_sg \shifter_0/oi_10_reg[3]  ( .D(n42562), .CP(clk), .Q(n68808) );
  dff_sg \shifter_0/oi_10_reg[4]  ( .D(n42550), .CP(clk), .Q(n68807) );
  dff_sg \shifter_0/oi_10_reg[5]  ( .D(n42556), .CP(clk), .Q(n68806) );
  dff_sg \shifter_0/oi_10_reg[6]  ( .D(n42246), .CP(clk), .Q(n68805) );
  dff_sg \shifter_0/oi_10_reg[7]  ( .D(n42565), .CP(clk), .Q(n68804) );
  dff_sg \shifter_0/oi_10_reg[8]  ( .D(n42511), .CP(clk), .Q(n68803) );
  dff_sg \shifter_0/oi_10_reg[9]  ( .D(n42520), .CP(clk), .Q(n68802) );
  dff_sg \shifter_0/oi_10_reg[10]  ( .D(n42514), .CP(clk), .Q(n68801) );
  dff_sg \shifter_0/oi_10_reg[11]  ( .D(n42517), .CP(clk), .Q(n68800) );
  dff_sg \shifter_0/oi_10_reg[12]  ( .D(n42499), .CP(clk), .Q(n68799) );
  dff_sg \shifter_0/oi_10_reg[13]  ( .D(n42502), .CP(clk), .Q(n68798) );
  dff_sg \shifter_0/oi_10_reg[14]  ( .D(n42505), .CP(clk), .Q(n68797) );
  dff_sg \shifter_0/oi_10_reg[15]  ( .D(n42508), .CP(clk), .Q(n68796) );
  dff_sg \shifter_0/oi_10_reg[16]  ( .D(n42272), .CP(clk), .Q(n68795) );
  dff_sg \shifter_0/oi_10_reg[17]  ( .D(n42322), .CP(clk), .Q(n68794) );
  dff_sg \shifter_0/oi_10_reg[18]  ( .D(n42247), .CP(clk), .Q(n68793) );
  dff_sg \shifter_0/oi_10_reg[19]  ( .D(n42325), .CP(clk), .Q(n68792) );
  dff_sg \shifter_0/oi_9_reg[0]  ( .D(n42248), .CP(clk), .Q(n68791) );
  dff_sg \shifter_0/oi_9_reg[1]  ( .D(n42302), .CP(clk), .Q(n68790) );
  dff_sg \shifter_0/oi_9_reg[2]  ( .D(n42269), .CP(clk), .Q(n68789) );
  dff_sg \shifter_0/oi_9_reg[3]  ( .D(n42260), .CP(clk), .Q(n68788) );
  dff_sg \shifter_0/oi_9_reg[4]  ( .D(n42278), .CP(clk), .Q(n68787) );
  dff_sg \shifter_0/oi_9_reg[5]  ( .D(n42275), .CP(clk), .Q(n68786) );
  dff_sg \shifter_0/oi_9_reg[6]  ( .D(n42309), .CP(clk), .Q(n68785) );
  dff_sg \shifter_0/oi_9_reg[7]  ( .D(n42312), .CP(clk), .Q(n68784) );
  dff_sg \shifter_0/oi_9_reg[8]  ( .D(n42315), .CP(clk), .Q(n68783) );
  dff_sg \shifter_0/oi_9_reg[9]  ( .D(n42318), .CP(clk), .Q(n68782) );
  dff_sg \shifter_0/oi_9_reg[10]  ( .D(n42263), .CP(clk), .Q(n68781) );
  dff_sg \shifter_0/oi_9_reg[11]  ( .D(n42266), .CP(clk), .Q(n68780) );
  dff_sg \shifter_0/oi_9_reg[12]  ( .D(n42329), .CP(clk), .Q(n68779) );
  dff_sg \shifter_0/oi_9_reg[13]  ( .D(n42332), .CP(clk), .Q(n68778) );
  dff_sg \shifter_0/oi_9_reg[14]  ( .D(n42335), .CP(clk), .Q(n68777) );
  dff_sg \shifter_0/oi_9_reg[15]  ( .D(n42344), .CP(clk), .Q(n68776) );
  dff_sg \shifter_0/oi_9_reg[16]  ( .D(n42228), .CP(clk), .Q(n68775) );
  dff_sg \shifter_0/oi_9_reg[17]  ( .D(n42341), .CP(clk), .Q(n68774) );
  dff_sg \shifter_0/oi_9_reg[18]  ( .D(n42305), .CP(clk), .Q(n68773) );
  dff_sg \shifter_0/oi_9_reg[19]  ( .D(n42772), .CP(clk), .Q(n68772) );
  dff_sg \shifter_0/oi_8_reg[0]  ( .D(n42296), .CP(clk), .Q(n68771) );
  dff_sg \shifter_0/oi_8_reg[1]  ( .D(n42299), .CP(clk), .Q(n68770) );
  dff_sg \shifter_0/oi_8_reg[2]  ( .D(n42249), .CP(clk), .Q(n68769) );
  dff_sg \shifter_0/oi_8_reg[3]  ( .D(n42293), .CP(clk), .Q(n68768) );
  dff_sg \shifter_0/oi_8_reg[4]  ( .D(n42281), .CP(clk), .Q(n68767) );
  dff_sg \shifter_0/oi_8_reg[5]  ( .D(n42284), .CP(clk), .Q(n68766) );
  dff_sg \shifter_0/oi_8_reg[6]  ( .D(n42287), .CP(clk), .Q(n68765) );
  dff_sg \shifter_0/oi_8_reg[7]  ( .D(n42290), .CP(clk), .Q(n68764) );
  dff_sg \shifter_0/oi_8_reg[8]  ( .D(n42742), .CP(clk), .Q(n68763) );
  dff_sg \shifter_0/oi_8_reg[9]  ( .D(n42219), .CP(clk), .Q(n68762) );
  dff_sg \shifter_0/oi_8_reg[10]  ( .D(n42423), .CP(clk), .Q(n68761) );
  dff_sg \shifter_0/oi_8_reg[11]  ( .D(n42192), .CP(clk), .Q(n68760) );
  dff_sg \shifter_0/oi_8_reg[12]  ( .D(n42652), .CP(clk), .Q(n68759) );
  dff_sg \shifter_0/oi_8_reg[13]  ( .D(n42655), .CP(clk), .Q(n68758) );
  dff_sg \shifter_0/oi_8_reg[14]  ( .D(n42661), .CP(clk), .Q(n68757) );
  dff_sg \shifter_0/oi_8_reg[15]  ( .D(n42664), .CP(clk), .Q(n68756) );
  dff_sg \shifter_0/oi_8_reg[16]  ( .D(n42637), .CP(clk), .Q(n68755) );
  dff_sg \shifter_0/oi_8_reg[17]  ( .D(n42634), .CP(clk), .Q(n68754) );
  dff_sg \shifter_0/oi_8_reg[18]  ( .D(n42646), .CP(clk), .Q(n68753) );
  dff_sg \shifter_0/oi_8_reg[19]  ( .D(n42640), .CP(clk), .Q(n68752) );
  dff_sg \shifter_0/oi_7_reg[0]  ( .D(n42619), .CP(clk), .Q(n68751) );
  dff_sg \shifter_0/oi_7_reg[1]  ( .D(n42622), .CP(clk), .Q(n68750) );
  dff_sg \shifter_0/oi_7_reg[2]  ( .D(n42625), .CP(clk), .Q(n68749) );
  dff_sg \shifter_0/oi_7_reg[3]  ( .D(n42628), .CP(clk), .Q(n68748) );
  dff_sg \shifter_0/oi_7_reg[4]  ( .D(n42724), .CP(clk), .Q(n68747) );
  dff_sg \shifter_0/oi_7_reg[5]  ( .D(n42419), .CP(clk), .Q(n68746) );
  dff_sg \shifter_0/oi_7_reg[6]  ( .D(n42165), .CP(clk), .Q(n68745) );
  dff_sg \shifter_0/oi_7_reg[7]  ( .D(n42715), .CP(clk), .Q(n68744) );
  dff_sg \shifter_0/oi_7_reg[8]  ( .D(n42541), .CP(clk), .Q(n68743) );
  dff_sg \shifter_0/oi_7_reg[9]  ( .D(n42386), .CP(clk), .Q(n68742) );
  dff_sg \shifter_0/oi_7_reg[10]  ( .D(n42411), .CP(clk), .Q(n68741) );
  dff_sg \shifter_0/oi_7_reg[11]  ( .D(n42328), .CP(clk), .Q(n68740) );
  dff_sg \shifter_0/oi_7_reg[12]  ( .D(n42670), .CP(clk), .Q(n68739) );
  dff_sg \shifter_0/oi_7_reg[13]  ( .D(n42673), .CP(clk), .Q(n68738) );
  dff_sg \shifter_0/oi_7_reg[14]  ( .D(n42676), .CP(clk), .Q(n68737) );
  dff_sg \shifter_0/oi_7_reg[15]  ( .D(n42679), .CP(clk), .Q(n68736) );
  dff_sg \shifter_0/oi_7_reg[16]  ( .D(n42174), .CP(clk), .Q(n68735) );
  dff_sg \shifter_0/oi_7_reg[17]  ( .D(n42177), .CP(clk), .Q(n68734) );
  dff_sg \shifter_0/oi_7_reg[18]  ( .D(n42685), .CP(clk), .Q(n68733) );
  dff_sg \shifter_0/oi_7_reg[19]  ( .D(n42688), .CP(clk), .Q(n68732) );
  dff_sg \shifter_0/oi_6_reg[0]  ( .D(n42414), .CP(clk), .Q(n68731) );
  dff_sg \shifter_0/oi_6_reg[1]  ( .D(n42243), .CP(clk), .Q(n68730) );
  dff_sg \shifter_0/oi_6_reg[2]  ( .D(n42616), .CP(clk), .Q(n68729) );
  dff_sg \shifter_0/oi_6_reg[3]  ( .D(n42257), .CP(clk), .Q(n68728) );
  dff_sg \shifter_0/oi_6_reg[4]  ( .D(n42189), .CP(clk), .Q(n68727) );
  dff_sg \shifter_0/oi_6_reg[5]  ( .D(n42667), .CP(clk), .Q(n68726) );
  dff_sg \shifter_0/oi_6_reg[6]  ( .D(n42682), .CP(clk), .Q(n68725) );
  dff_sg \shifter_0/oi_6_reg[7]  ( .D(n42251), .CP(clk), .Q(n68724) );
  dff_sg \shifter_0/oi_6_reg[8]  ( .D(n42583), .CP(clk), .Q(n68723) );
  dff_sg \shifter_0/oi_6_reg[9]  ( .D(n42574), .CP(clk), .Q(n68722) );
  dff_sg \shifter_0/oi_6_reg[10]  ( .D(n42631), .CP(clk), .Q(n68721) );
  dff_sg \shifter_0/oi_6_reg[11]  ( .D(n42643), .CP(clk), .Q(n68720) );
  dff_sg \shifter_0/oi_6_reg[12]  ( .D(n42250), .CP(clk), .Q(n68719) );
  dff_sg \shifter_0/oi_6_reg[13]  ( .D(n42658), .CP(clk), .Q(n68718) );
  dff_sg \shifter_0/oi_6_reg[14]  ( .D(n42601), .CP(clk), .Q(n68717) );
  dff_sg \shifter_0/oi_6_reg[15]  ( .D(n42592), .CP(clk), .Q(n68716) );
  dff_sg \shifter_0/oi_6_reg[16]  ( .D(n42595), .CP(clk), .Q(n68715) );
  dff_sg \shifter_0/oi_6_reg[17]  ( .D(n42598), .CP(clk), .Q(n68714) );
  dff_sg \shifter_0/oi_6_reg[18]  ( .D(n42604), .CP(clk), .Q(n68713) );
  dff_sg \shifter_0/oi_6_reg[19]  ( .D(n42607), .CP(clk), .Q(n68712) );
  dff_sg \shifter_0/oi_5_reg[0]  ( .D(n42577), .CP(clk), .Q(n68711) );
  dff_sg \shifter_0/oi_5_reg[1]  ( .D(n42580), .CP(clk), .Q(n68710) );
  dff_sg \shifter_0/oi_5_reg[2]  ( .D(n42586), .CP(clk), .Q(n68709) );
  dff_sg \shifter_0/oi_5_reg[3]  ( .D(n42589), .CP(clk), .Q(n68708) );
  dff_sg \shifter_0/oi_5_reg[4]  ( .D(n42421), .CP(clk), .Q(n68707) );
  dff_sg \shifter_0/oi_5_reg[5]  ( .D(n42258), .CP(clk), .Q(n68706) );
  dff_sg \shifter_0/oi_5_reg[6]  ( .D(n42417), .CP(clk), .Q(n68705) );
  dff_sg \shifter_0/oi_5_reg[7]  ( .D(n42259), .CP(clk), .Q(n68704) );
  dff_sg \shifter_0/oi_5_reg[8]  ( .D(n42649), .CP(clk), .Q(n68703) );
  dff_sg \shifter_0/oi_5_reg[9]  ( .D(n42571), .CP(clk), .Q(n68702) );
  dff_sg \shifter_0/oi_5_reg[10]  ( .D(n42610), .CP(clk), .Q(n68701) );
  dff_sg \shifter_0/oi_5_reg[11]  ( .D(n42613), .CP(clk), .Q(n68700) );
  dff_sg \shifter_0/oi_5_reg[12]  ( .D(n42424), .CP(clk), .Q(n68699) );
  dff_sg \shifter_0/oi_5_reg[13]  ( .D(n42427), .CP(clk), .Q(n68698) );
  dff_sg \shifter_0/oi_5_reg[14]  ( .D(n42445), .CP(clk), .Q(n68697) );
  dff_sg \shifter_0/oi_5_reg[15]  ( .D(n42433), .CP(clk), .Q(n68696) );
  dff_sg \shifter_0/oi_5_reg[16]  ( .D(n42787), .CP(clk), .Q(n68695) );
  dff_sg \shifter_0/oi_5_reg[17]  ( .D(n42436), .CP(clk), .Q(n68694) );
  dff_sg \shifter_0/oi_5_reg[18]  ( .D(n42439), .CP(clk), .Q(n68693) );
  dff_sg \shifter_0/oi_5_reg[19]  ( .D(n42442), .CP(clk), .Q(n68692) );
  dff_sg \shifter_0/oi_4_reg[0]  ( .D(n42448), .CP(clk), .Q(n68691) );
  dff_sg \shifter_0/oi_4_reg[1]  ( .D(n42451), .CP(clk), .Q(n68690) );
  dff_sg \shifter_0/oi_4_reg[2]  ( .D(n42466), .CP(clk), .Q(n68689) );
  dff_sg \shifter_0/oi_4_reg[3]  ( .D(n42454), .CP(clk), .Q(n68688) );
  dff_sg \shifter_0/oi_4_reg[4]  ( .D(n42457), .CP(clk), .Q(n68687) );
  dff_sg \shifter_0/oi_4_reg[5]  ( .D(n42460), .CP(clk), .Q(n68686) );
  dff_sg \shifter_0/oi_4_reg[6]  ( .D(n42308), .CP(clk), .Q(n68685) );
  dff_sg \shifter_0/oi_4_reg[7]  ( .D(n42463), .CP(clk), .Q(n68684) );
  dff_sg \shifter_0/oi_4_reg[8]  ( .D(n42469), .CP(clk), .Q(n68683) );
  dff_sg \shifter_0/oi_4_reg[9]  ( .D(n42472), .CP(clk), .Q(n68682) );
  dff_sg \shifter_0/oi_4_reg[10]  ( .D(n42321), .CP(clk), .Q(n68681) );
  dff_sg \shifter_0/oi_4_reg[11]  ( .D(n42475), .CP(clk), .Q(n68680) );
  dff_sg \shifter_0/oi_4_reg[12]  ( .D(n42326), .CP(clk), .Q(n68679) );
  dff_sg \shifter_0/oi_4_reg[13]  ( .D(n42327), .CP(clk), .Q(n68678) );
  dff_sg \shifter_0/oi_4_reg[14]  ( .D(n42323), .CP(clk), .Q(n68677) );
  dff_sg \shifter_0/oi_4_reg[15]  ( .D(n42324), .CP(clk), .Q(n68676) );
  dff_sg \shifter_0/oi_4_reg[16]  ( .D(n42313), .CP(clk), .Q(n68675) );
  dff_sg \shifter_0/oi_4_reg[17]  ( .D(n42314), .CP(clk), .Q(n68674) );
  dff_sg \shifter_0/oi_4_reg[18]  ( .D(n42310), .CP(clk), .Q(n68673) );
  dff_sg \shifter_0/oi_4_reg[19]  ( .D(n42311), .CP(clk), .Q(n68672) );
  dff_sg \shifter_0/oi_3_reg[0]  ( .D(n42319), .CP(clk), .Q(n68671) );
  dff_sg \shifter_0/oi_3_reg[1]  ( .D(n42320), .CP(clk), .Q(n68670) );
  dff_sg \shifter_0/oi_3_reg[2]  ( .D(n42316), .CP(clk), .Q(n68669) );
  dff_sg \shifter_0/oi_3_reg[3]  ( .D(n42317), .CP(clk), .Q(n68668) );
  dff_sg \shifter_0/oi_3_reg[4]  ( .D(n42276), .CP(clk), .Q(n68667) );
  dff_sg \shifter_0/oi_3_reg[5]  ( .D(n42277), .CP(clk), .Q(n68666) );
  dff_sg \shifter_0/oi_3_reg[6]  ( .D(n42273), .CP(clk), .Q(n68665) );
  dff_sg \shifter_0/oi_3_reg[7]  ( .D(n42274), .CP(clk), .Q(n68664) );
  dff_sg \shifter_0/oi_3_reg[8]  ( .D(n42282), .CP(clk), .Q(n68663) );
  dff_sg \shifter_0/oi_3_reg[9]  ( .D(n42283), .CP(clk), .Q(n68662) );
  dff_sg \shifter_0/oi_3_reg[10]  ( .D(n42279), .CP(clk), .Q(n68661) );
  dff_sg \shifter_0/oi_3_reg[11]  ( .D(n42280), .CP(clk), .Q(n68660) );
  dff_sg \shifter_0/oi_3_reg[12]  ( .D(n42264), .CP(clk), .Q(n68659) );
  dff_sg \shifter_0/oi_3_reg[13]  ( .D(n42265), .CP(clk), .Q(n68658) );
  dff_sg \shifter_0/oi_3_reg[14]  ( .D(n42261), .CP(clk), .Q(n68657) );
  dff_sg \shifter_0/oi_3_reg[15]  ( .D(n42262), .CP(clk), .Q(n68656) );
  dff_sg \shifter_0/oi_3_reg[16]  ( .D(n42270), .CP(clk), .Q(n68655) );
  dff_sg \shifter_0/oi_3_reg[17]  ( .D(n42271), .CP(clk), .Q(n68654) );
  dff_sg \shifter_0/oi_3_reg[18]  ( .D(n42267), .CP(clk), .Q(n68653) );
  dff_sg \shifter_0/oi_3_reg[19]  ( .D(n42268), .CP(clk), .Q(n68652) );
  dff_sg \shifter_0/oi_2_reg[0]  ( .D(n42300), .CP(clk), .Q(n68651) );
  dff_sg \shifter_0/oi_2_reg[1]  ( .D(n42301), .CP(clk), .Q(n68650) );
  dff_sg \shifter_0/oi_2_reg[2]  ( .D(n42297), .CP(clk), .Q(n68649) );
  dff_sg \shifter_0/oi_2_reg[3]  ( .D(n42298), .CP(clk), .Q(n68648) );
  dff_sg \shifter_0/oi_2_reg[4]  ( .D(n42306), .CP(clk), .Q(n68647) );
  dff_sg \shifter_0/oi_2_reg[5]  ( .D(n42307), .CP(clk), .Q(n68646) );
  dff_sg \shifter_0/oi_2_reg[6]  ( .D(n42303), .CP(clk), .Q(n68645) );
  dff_sg \shifter_0/oi_2_reg[7]  ( .D(n42304), .CP(clk), .Q(n68644) );
  dff_sg \shifter_0/oi_2_reg[8]  ( .D(n42288), .CP(clk), .Q(n68643) );
  dff_sg \shifter_0/oi_2_reg[9]  ( .D(n42289), .CP(clk), .Q(n68642) );
  dff_sg \shifter_0/oi_2_reg[10]  ( .D(n42285), .CP(clk), .Q(n68641) );
  dff_sg \shifter_0/oi_2_reg[11]  ( .D(n42286), .CP(clk), .Q(n68640) );
  dff_sg \shifter_0/oi_2_reg[12]  ( .D(n42294), .CP(clk), .Q(n68639) );
  dff_sg \shifter_0/oi_2_reg[13]  ( .D(n42295), .CP(clk), .Q(n68638) );
  dff_sg \shifter_0/oi_2_reg[14]  ( .D(n42291), .CP(clk), .Q(n68637) );
  dff_sg \shifter_0/oi_2_reg[15]  ( .D(n42292), .CP(clk), .Q(n68636) );
  dff_sg \shifter_0/oi_2_reg[16]  ( .D(n42387), .CP(clk), .Q(n68635) );
  dff_sg \shifter_0/oi_2_reg[17]  ( .D(n42388), .CP(clk), .Q(n68634) );
  dff_sg \shifter_0/oi_2_reg[18]  ( .D(n42384), .CP(clk), .Q(n68633) );
  dff_sg \shifter_0/oi_2_reg[19]  ( .D(n42385), .CP(clk), .Q(n68632) );
  dff_sg \shifter_0/oi_1_reg[0]  ( .D(n42393), .CP(clk), .Q(n68631) );
  dff_sg \shifter_0/oi_1_reg[1]  ( .D(n42394), .CP(clk), .Q(n68630) );
  dff_sg \shifter_0/oi_1_reg[2]  ( .D(n42390), .CP(clk), .Q(n68629) );
  dff_sg \shifter_0/oi_1_reg[3]  ( .D(n42391), .CP(clk), .Q(n68628) );
  dff_sg \shifter_0/oi_1_reg[4]  ( .D(n42375), .CP(clk), .Q(n68627) );
  dff_sg \shifter_0/oi_1_reg[5]  ( .D(n42376), .CP(clk), .Q(n68626) );
  dff_sg \shifter_0/oi_1_reg[6]  ( .D(n42372), .CP(clk), .Q(n68625) );
  dff_sg \shifter_0/oi_1_reg[7]  ( .D(n42373), .CP(clk), .Q(n68624) );
  dff_sg \shifter_0/oi_1_reg[8]  ( .D(n42381), .CP(clk), .Q(n68623) );
  dff_sg \shifter_0/oi_1_reg[9]  ( .D(n42382), .CP(clk), .Q(n68622) );
  dff_sg \shifter_0/oi_1_reg[10]  ( .D(n42378), .CP(clk), .Q(n68621) );
  dff_sg \shifter_0/oi_1_reg[11]  ( .D(n42379), .CP(clk), .Q(n68620) );
  dff_sg \shifter_0/oi_1_reg[12]  ( .D(n42412), .CP(clk), .Q(n68619) );
  dff_sg \shifter_0/oi_1_reg[13]  ( .D(n42413), .CP(clk), .Q(n68618) );
  dff_sg \shifter_0/oi_1_reg[14]  ( .D(n42409), .CP(clk), .Q(n68617) );
  dff_sg \shifter_0/oi_1_reg[15]  ( .D(n42410), .CP(clk), .Q(n68616) );
  dff_sg \shifter_0/oi_1_reg[16]  ( .D(n42775), .CP(clk), .Q(n68615) );
  dff_sg \shifter_0/oi_1_reg[17]  ( .D(n42778), .CP(clk), .Q(n68614) );
  dff_sg \shifter_0/oi_1_reg[18]  ( .D(n42781), .CP(clk), .Q(n68613) );
  dff_sg \shifter_0/oi_1_reg[19]  ( .D(n42784), .CP(clk), .Q(n68612) );
  dff_sg \shifter_0/oi_0_reg[0]  ( .D(n42399), .CP(clk), .Q(n68611) );
  dff_sg \shifter_0/oi_0_reg[1]  ( .D(n42400), .CP(clk), .Q(n68610) );
  dff_sg \shifter_0/oi_0_reg[2]  ( .D(n42396), .CP(clk), .Q(n68609) );
  dff_sg \shifter_0/oi_0_reg[3]  ( .D(n42397), .CP(clk), .Q(n68608) );
  dff_sg \shifter_0/oi_0_reg[4]  ( .D(n42405), .CP(clk), .Q(n68607) );
  dff_sg \shifter_0/oi_0_reg[5]  ( .D(n42406), .CP(clk), .Q(n68606) );
  dff_sg \shifter_0/oi_0_reg[6]  ( .D(n42402), .CP(clk), .Q(n68605) );
  dff_sg \shifter_0/oi_0_reg[7]  ( .D(n42403), .CP(clk), .Q(n68604) );
  dff_sg \shifter_0/oi_0_reg[8]  ( .D(n42339), .CP(clk), .Q(n68603) );
  dff_sg \shifter_0/oi_0_reg[9]  ( .D(n42340), .CP(clk), .Q(n68602) );
  dff_sg \shifter_0/oi_0_reg[10]  ( .D(n42336), .CP(clk), .Q(n68601) );
  dff_sg \shifter_0/oi_0_reg[11]  ( .D(n42337), .CP(clk), .Q(n68600) );
  dff_sg \shifter_0/oi_0_reg[12]  ( .D(n42345), .CP(clk), .Q(n68599) );
  dff_sg \shifter_0/oi_0_reg[13]  ( .D(n42346), .CP(clk), .Q(n68598) );
  dff_sg \shifter_0/oi_0_reg[14]  ( .D(n42342), .CP(clk), .Q(n68597) );
  dff_sg \shifter_0/oi_0_reg[15]  ( .D(n42343), .CP(clk), .Q(n68596) );
  dff_sg \shifter_0/oi_0_reg[16]  ( .D(n42229), .CP(clk), .Q(n68595) );
  dff_sg \shifter_0/oi_0_reg[17]  ( .D(n42230), .CP(clk), .Q(n68594) );
  dff_sg \shifter_0/oi_0_reg[18]  ( .D(n42766), .CP(clk), .Q(n68593) );
  dff_sg \shifter_0/oi_0_reg[19]  ( .D(n42769), .CP(clk), .Q(n68592) );
  dff_sg \shifter_0/ow_15_reg[0]  ( .D(n42333), .CP(clk), .Q(n69231) );
  dff_sg \shifter_0/ow_15_reg[1]  ( .D(n42334), .CP(clk), .Q(n69230) );
  dff_sg \shifter_0/ow_15_reg[2]  ( .D(n42330), .CP(clk), .Q(n69229) );
  dff_sg \shifter_0/ow_15_reg[3]  ( .D(n42331), .CP(clk), .Q(n69228) );
  dff_sg \shifter_0/ow_15_reg[4]  ( .D(n42363), .CP(clk), .Q(n69227) );
  dff_sg \shifter_0/ow_15_reg[5]  ( .D(n42364), .CP(clk), .Q(n69226) );
  dff_sg \shifter_0/ow_15_reg[6]  ( .D(n42360), .CP(clk), .Q(n69225) );
  dff_sg \shifter_0/ow_15_reg[7]  ( .D(n42361), .CP(clk), .Q(n69224) );
  dff_sg \shifter_0/ow_15_reg[8]  ( .D(n42369), .CP(clk), .Q(n69223) );
  dff_sg \shifter_0/ow_15_reg[9]  ( .D(n42370), .CP(clk), .Q(n69222) );
  dff_sg \shifter_0/ow_15_reg[10]  ( .D(n42366), .CP(clk), .Q(n69221) );
  dff_sg \shifter_0/ow_15_reg[11]  ( .D(n42367), .CP(clk), .Q(n69220) );
  dff_sg \shifter_0/ow_15_reg[12]  ( .D(n42351), .CP(clk), .Q(n69219) );
  dff_sg \shifter_0/ow_15_reg[13]  ( .D(n42352), .CP(clk), .Q(n69218) );
  dff_sg \shifter_0/ow_15_reg[14]  ( .D(n42348), .CP(clk), .Q(n69217) );
  dff_sg \shifter_0/ow_15_reg[15]  ( .D(n42349), .CP(clk), .Q(n69216) );
  dff_sg \shifter_0/ow_15_reg[16]  ( .D(n42357), .CP(clk), .Q(n69215) );
  dff_sg \shifter_0/ow_15_reg[17]  ( .D(n42358), .CP(clk), .Q(n69214) );
  dff_sg \shifter_0/ow_15_reg[18]  ( .D(n42354), .CP(clk), .Q(n69213) );
  dff_sg \shifter_0/ow_15_reg[19]  ( .D(n42355), .CP(clk), .Q(n69212) );
  dff_sg \shifter_0/i_pointer_reg[0]  ( .D(n42813), .CP(clk), .Q(
        \shifter_0/i_pointer [0]) );
  dff_sg \shifter_0/i_pointer_reg[1]  ( .D(n42811), .CP(clk), .Q(
        \shifter_0/i_pointer [1]) );
  dff_sg \shifter_0/i_pointer_reg[2]  ( .D(n42812), .CP(clk), .Q(
        \shifter_0/i_pointer [2]) );
  dff_sg \shifter_0/i_pointer_reg[3]  ( .D(n42814), .CP(clk), .Q(
        \shifter_0/i_pointer [3]) );
  dff_sg \shifter_0/input_taken_reg  ( .D(\shifter_0/n14056 ), .CP(clk), .Q(
        \shifter_0/n27116 ) );
  dff_sg \shifter_0/reg_i_0_reg[0]  ( .D(n42049), .CP(clk), .Q(
        \shifter_0/reg_i_0 [0]) );
  dff_sg \shifter_0/reg_i_0_reg[1]  ( .D(n42134), .CP(clk), .Q(
        \shifter_0/reg_i_0 [1]) );
  dff_sg \shifter_0/reg_i_0_reg[2]  ( .D(n42113), .CP(clk), .Q(
        \shifter_0/reg_i_0 [2]) );
  dff_sg \shifter_0/reg_i_0_reg[3]  ( .D(n42109), .CP(clk), .Q(
        \shifter_0/reg_i_0 [3]) );
  dff_sg \shifter_0/reg_i_0_reg[4]  ( .D(n41916), .CP(clk), .Q(
        \shifter_0/reg_i_0 [4]) );
  dff_sg \shifter_0/reg_i_0_reg[5]  ( .D(n42149), .CP(clk), .Q(
        \shifter_0/reg_i_0 [5]) );
  dff_sg \shifter_0/reg_i_0_reg[6]  ( .D(n41723), .CP(clk), .Q(
        \shifter_0/reg_i_0 [6]) );
  dff_sg \shifter_0/reg_i_0_reg[7]  ( .D(n41962), .CP(clk), .Q(
        \shifter_0/reg_i_0 [7]) );
  dff_sg \shifter_0/reg_i_0_reg[8]  ( .D(n42128), .CP(clk), .Q(
        \shifter_0/reg_i_0 [8]) );
  dff_sg \shifter_0/reg_i_0_reg[9]  ( .D(n42131), .CP(clk), .Q(
        \shifter_0/reg_i_0 [9]) );
  dff_sg \shifter_0/reg_i_0_reg[10]  ( .D(n41917), .CP(clk), .Q(
        \shifter_0/reg_i_0 [10]) );
  dff_sg \shifter_0/reg_i_0_reg[11]  ( .D(n41980), .CP(clk), .Q(
        \shifter_0/reg_i_0 [11]) );
  dff_sg \shifter_0/reg_i_0_reg[12]  ( .D(n42129), .CP(clk), .Q(
        \shifter_0/reg_i_0 [12]) );
  dff_sg \shifter_0/reg_i_0_reg[13]  ( .D(n42130), .CP(clk), .Q(
        \shifter_0/reg_i_0 [13]) );
  dff_sg \shifter_0/reg_i_0_reg[14]  ( .D(n42126), .CP(clk), .Q(
        \shifter_0/reg_i_0 [14]) );
  dff_sg \shifter_0/reg_i_0_reg[15]  ( .D(n42127), .CP(clk), .Q(
        \shifter_0/reg_i_0 [15]) );
  dff_sg \shifter_0/reg_i_0_reg[16]  ( .D(n42135), .CP(clk), .Q(
        \shifter_0/reg_i_0 [16]) );
  dff_sg \shifter_0/reg_i_0_reg[17]  ( .D(n42136), .CP(clk), .Q(
        \shifter_0/reg_i_0 [17]) );
  dff_sg \shifter_0/reg_i_0_reg[18]  ( .D(n42132), .CP(clk), .Q(
        \shifter_0/reg_i_0 [18]) );
  dff_sg \shifter_0/reg_i_0_reg[19]  ( .D(n42133), .CP(clk), .Q(
        \shifter_0/reg_i_0 [19]) );
  dff_sg \shifter_0/reg_i_1_reg[0]  ( .D(n42117), .CP(clk), .Q(
        \shifter_0/reg_i_1 [0]) );
  dff_sg \shifter_0/reg_i_1_reg[1]  ( .D(n42118), .CP(clk), .Q(
        \shifter_0/reg_i_1 [1]) );
  dff_sg \shifter_0/reg_i_1_reg[2]  ( .D(n42114), .CP(clk), .Q(
        \shifter_0/reg_i_1 [2]) );
  dff_sg \shifter_0/reg_i_1_reg[3]  ( .D(n42115), .CP(clk), .Q(
        \shifter_0/reg_i_1 [3]) );
  dff_sg \shifter_0/reg_i_1_reg[4]  ( .D(n42123), .CP(clk), .Q(
        \shifter_0/reg_i_1 [4]) );
  dff_sg \shifter_0/reg_i_1_reg[5]  ( .D(n42124), .CP(clk), .Q(
        \shifter_0/reg_i_1 [5]) );
  dff_sg \shifter_0/reg_i_1_reg[6]  ( .D(n42120), .CP(clk), .Q(
        \shifter_0/reg_i_1 [6]) );
  dff_sg \shifter_0/reg_i_1_reg[7]  ( .D(n42121), .CP(clk), .Q(
        \shifter_0/reg_i_1 [7]) );
  dff_sg \shifter_0/reg_i_1_reg[8]  ( .D(n42153), .CP(clk), .Q(
        \shifter_0/reg_i_1 [8]) );
  dff_sg \shifter_0/reg_i_1_reg[9]  ( .D(n42154), .CP(clk), .Q(
        \shifter_0/reg_i_1 [9]) );
  dff_sg \shifter_0/reg_i_1_reg[10]  ( .D(n42150), .CP(clk), .Q(
        \shifter_0/reg_i_1 [10]) );
  dff_sg \shifter_0/reg_i_1_reg[11]  ( .D(n42151), .CP(clk), .Q(
        \shifter_0/reg_i_1 [11]) );
  dff_sg \shifter_0/reg_i_1_reg[12]  ( .D(n42159), .CP(clk), .Q(
        \shifter_0/reg_i_1 [12]) );
  dff_sg \shifter_0/reg_i_1_reg[13]  ( .D(n42160), .CP(clk), .Q(
        \shifter_0/reg_i_1 [13]) );
  dff_sg \shifter_0/reg_i_1_reg[14]  ( .D(n42156), .CP(clk), .Q(
        \shifter_0/reg_i_1 [14]) );
  dff_sg \shifter_0/reg_i_1_reg[15]  ( .D(n42157), .CP(clk), .Q(
        \shifter_0/reg_i_1 [15]) );
  dff_sg \shifter_0/reg_i_1_reg[16]  ( .D(n42141), .CP(clk), .Q(
        \shifter_0/reg_i_1 [16]) );
  dff_sg \shifter_0/reg_i_1_reg[17]  ( .D(n42142), .CP(clk), .Q(
        \shifter_0/reg_i_1 [17]) );
  dff_sg \shifter_0/reg_i_1_reg[18]  ( .D(n42138), .CP(clk), .Q(
        \shifter_0/reg_i_1 [18]) );
  dff_sg \shifter_0/reg_i_1_reg[19]  ( .D(n42139), .CP(clk), .Q(
        \shifter_0/reg_i_1 [19]) );
  dff_sg \shifter_0/reg_i_2_reg[0]  ( .D(n42147), .CP(clk), .Q(
        \shifter_0/reg_i_2 [0]) );
  dff_sg \shifter_0/reg_i_2_reg[1]  ( .D(n42148), .CP(clk), .Q(
        \shifter_0/reg_i_2 [1]) );
  dff_sg \shifter_0/reg_i_2_reg[2]  ( .D(n42144), .CP(clk), .Q(
        \shifter_0/reg_i_2 [2]) );
  dff_sg \shifter_0/reg_i_2_reg[3]  ( .D(n42145), .CP(clk), .Q(
        \shifter_0/reg_i_2 [3]) );
  dff_sg \shifter_0/reg_i_2_reg[4]  ( .D(n41981), .CP(clk), .Q(
        \shifter_0/reg_i_2 [4]) );
  dff_sg \shifter_0/reg_i_2_reg[5]  ( .D(n41982), .CP(clk), .Q(
        \shifter_0/reg_i_2 [5]) );
  dff_sg \shifter_0/reg_i_2_reg[6]  ( .D(n41978), .CP(clk), .Q(
        \shifter_0/reg_i_2 [6]) );
  dff_sg \shifter_0/reg_i_2_reg[7]  ( .D(n41979), .CP(clk), .Q(
        \shifter_0/reg_i_2 [7]) );
  dff_sg \shifter_0/reg_i_2_reg[8]  ( .D(n41987), .CP(clk), .Q(
        \shifter_0/reg_i_2 [8]) );
  dff_sg \shifter_0/reg_i_2_reg[9]  ( .D(n41988), .CP(clk), .Q(
        \shifter_0/reg_i_2 [9]) );
  dff_sg \shifter_0/reg_i_2_reg[10]  ( .D(n41984), .CP(clk), .Q(
        \shifter_0/reg_i_2 [10]) );
  dff_sg \shifter_0/reg_i_2_reg[11]  ( .D(n41985), .CP(clk), .Q(
        \shifter_0/reg_i_2 [11]) );
  dff_sg \shifter_0/reg_i_2_reg[12]  ( .D(n41969), .CP(clk), .Q(
        \shifter_0/reg_i_2 [12]) );
  dff_sg \shifter_0/reg_i_2_reg[13]  ( .D(n41970), .CP(clk), .Q(
        \shifter_0/reg_i_2 [13]) );
  dff_sg \shifter_0/reg_i_2_reg[14]  ( .D(n41966), .CP(clk), .Q(
        \shifter_0/reg_i_2 [14]) );
  dff_sg \shifter_0/reg_i_2_reg[15]  ( .D(n41967), .CP(clk), .Q(
        \shifter_0/reg_i_2 [15]) );
  dff_sg \shifter_0/reg_i_2_reg[16]  ( .D(n41975), .CP(clk), .Q(
        \shifter_0/reg_i_2 [16]) );
  dff_sg \shifter_0/reg_i_2_reg[17]  ( .D(n41976), .CP(clk), .Q(
        \shifter_0/reg_i_2 [17]) );
  dff_sg \shifter_0/reg_i_2_reg[18]  ( .D(n41972), .CP(clk), .Q(
        \shifter_0/reg_i_2 [18]) );
  dff_sg \shifter_0/reg_i_2_reg[19]  ( .D(n41973), .CP(clk), .Q(
        \shifter_0/reg_i_2 [19]) );
  dff_sg \shifter_0/reg_i_3_reg[0]  ( .D(n42005), .CP(clk), .Q(
        \shifter_0/reg_i_3 [0]) );
  dff_sg \shifter_0/reg_i_3_reg[1]  ( .D(n42006), .CP(clk), .Q(
        \shifter_0/reg_i_3 [1]) );
  dff_sg \shifter_0/reg_i_3_reg[2]  ( .D(n42002), .CP(clk), .Q(
        \shifter_0/reg_i_3 [2]) );
  dff_sg \shifter_0/reg_i_3_reg[3]  ( .D(n42003), .CP(clk), .Q(
        \shifter_0/reg_i_3 [3]) );
  dff_sg \shifter_0/reg_i_3_reg[4]  ( .D(n42011), .CP(clk), .Q(
        \shifter_0/reg_i_3 [4]) );
  dff_sg \shifter_0/reg_i_3_reg[5]  ( .D(n42012), .CP(clk), .Q(
        \shifter_0/reg_i_3 [5]) );
  dff_sg \shifter_0/reg_i_3_reg[6]  ( .D(n42008), .CP(clk), .Q(
        \shifter_0/reg_i_3 [6]) );
  dff_sg \shifter_0/reg_i_3_reg[7]  ( .D(n42009), .CP(clk), .Q(
        \shifter_0/reg_i_3 [7]) );
  dff_sg \shifter_0/reg_i_3_reg[8]  ( .D(n41993), .CP(clk), .Q(
        \shifter_0/reg_i_3 [8]) );
  dff_sg \shifter_0/reg_i_3_reg[9]  ( .D(n41994), .CP(clk), .Q(
        \shifter_0/reg_i_3 [9]) );
  dff_sg \shifter_0/reg_i_3_reg[10]  ( .D(n41990), .CP(clk), .Q(
        \shifter_0/reg_i_3 [10]) );
  dff_sg \shifter_0/reg_i_3_reg[11]  ( .D(n41991), .CP(clk), .Q(
        \shifter_0/reg_i_3 [11]) );
  dff_sg \shifter_0/reg_i_3_reg[12]  ( .D(n41999), .CP(clk), .Q(
        \shifter_0/reg_i_3 [12]) );
  dff_sg \shifter_0/reg_i_3_reg[13]  ( .D(n42000), .CP(clk), .Q(
        \shifter_0/reg_i_3 [13]) );
  dff_sg \shifter_0/reg_i_3_reg[14]  ( .D(n41996), .CP(clk), .Q(
        \shifter_0/reg_i_3 [14]) );
  dff_sg \shifter_0/reg_i_3_reg[15]  ( .D(n41997), .CP(clk), .Q(
        \shifter_0/reg_i_3 [15]) );
  dff_sg \shifter_0/reg_i_3_reg[16]  ( .D(n41933), .CP(clk), .Q(
        \shifter_0/reg_i_3 [16]) );
  dff_sg \shifter_0/reg_i_3_reg[17]  ( .D(n41934), .CP(clk), .Q(
        \shifter_0/reg_i_3 [17]) );
  dff_sg \shifter_0/reg_i_3_reg[18]  ( .D(n41930), .CP(clk), .Q(
        \shifter_0/reg_i_3 [18]) );
  dff_sg \shifter_0/reg_i_3_reg[19]  ( .D(n41931), .CP(clk), .Q(
        \shifter_0/reg_i_3 [19]) );
  dff_sg \shifter_0/reg_i_4_reg[0]  ( .D(n41939), .CP(clk), .Q(
        \shifter_0/reg_i_4 [0]) );
  dff_sg \shifter_0/reg_i_4_reg[1]  ( .D(n41940), .CP(clk), .Q(
        \shifter_0/reg_i_4 [1]) );
  dff_sg \shifter_0/reg_i_4_reg[2]  ( .D(n41936), .CP(clk), .Q(
        \shifter_0/reg_i_4 [2]) );
  dff_sg \shifter_0/reg_i_4_reg[3]  ( .D(n41937), .CP(clk), .Q(
        \shifter_0/reg_i_4 [3]) );
  dff_sg \shifter_0/reg_i_4_reg[4]  ( .D(n41921), .CP(clk), .Q(
        \shifter_0/reg_i_4 [4]) );
  dff_sg \shifter_0/reg_i_4_reg[5]  ( .D(n41922), .CP(clk), .Q(
        \shifter_0/reg_i_4 [5]) );
  dff_sg \shifter_0/reg_i_4_reg[6]  ( .D(n41918), .CP(clk), .Q(
        \shifter_0/reg_i_4 [6]) );
  dff_sg \shifter_0/reg_i_4_reg[7]  ( .D(n41919), .CP(clk), .Q(
        \shifter_0/reg_i_4 [7]) );
  dff_sg \shifter_0/reg_i_4_reg[8]  ( .D(n41927), .CP(clk), .Q(
        \shifter_0/reg_i_4 [8]) );
  dff_sg \shifter_0/reg_i_4_reg[9]  ( .D(n41928), .CP(clk), .Q(
        \shifter_0/reg_i_4 [9]) );
  dff_sg \shifter_0/reg_i_4_reg[10]  ( .D(n41924), .CP(clk), .Q(
        \shifter_0/reg_i_4 [10]) );
  dff_sg \shifter_0/reg_i_4_reg[11]  ( .D(n41925), .CP(clk), .Q(
        \shifter_0/reg_i_4 [11]) );
  dff_sg \shifter_0/reg_i_4_reg[12]  ( .D(n41957), .CP(clk), .Q(
        \shifter_0/reg_i_4 [12]) );
  dff_sg \shifter_0/reg_i_4_reg[13]  ( .D(n41958), .CP(clk), .Q(
        \shifter_0/reg_i_4 [13]) );
  dff_sg \shifter_0/reg_i_4_reg[14]  ( .D(n41954), .CP(clk), .Q(
        \shifter_0/reg_i_4 [14]) );
  dff_sg \shifter_0/reg_i_4_reg[15]  ( .D(n41955), .CP(clk), .Q(
        \shifter_0/reg_i_4 [15]) );
  dff_sg \shifter_0/reg_i_4_reg[16]  ( .D(n41963), .CP(clk), .Q(
        \shifter_0/reg_i_4 [16]) );
  dff_sg \shifter_0/reg_i_4_reg[17]  ( .D(n41964), .CP(clk), .Q(
        \shifter_0/reg_i_4 [17]) );
  dff_sg \shifter_0/reg_i_4_reg[18]  ( .D(n41960), .CP(clk), .Q(
        \shifter_0/reg_i_4 [18]) );
  dff_sg \shifter_0/reg_i_4_reg[19]  ( .D(n41961), .CP(clk), .Q(
        \shifter_0/reg_i_4 [19]) );
  dff_sg \shifter_0/reg_i_5_reg[0]  ( .D(n41945), .CP(clk), .Q(
        \shifter_0/reg_i_5 [0]) );
  dff_sg \shifter_0/reg_i_5_reg[1]  ( .D(n41946), .CP(clk), .Q(
        \shifter_0/reg_i_5 [1]) );
  dff_sg \shifter_0/reg_i_5_reg[2]  ( .D(n41942), .CP(clk), .Q(
        \shifter_0/reg_i_5 [2]) );
  dff_sg \shifter_0/reg_i_5_reg[3]  ( .D(n41943), .CP(clk), .Q(
        \shifter_0/reg_i_5 [3]) );
  dff_sg \shifter_0/reg_i_5_reg[4]  ( .D(n41951), .CP(clk), .Q(
        \shifter_0/reg_i_5 [4]) );
  dff_sg \shifter_0/reg_i_5_reg[5]  ( .D(n41952), .CP(clk), .Q(
        \shifter_0/reg_i_5 [5]) );
  dff_sg \shifter_0/reg_i_5_reg[6]  ( .D(n41948), .CP(clk), .Q(
        \shifter_0/reg_i_5 [6]) );
  dff_sg \shifter_0/reg_i_5_reg[7]  ( .D(n41949), .CP(clk), .Q(
        \shifter_0/reg_i_5 [7]) );
  dff_sg \shifter_0/reg_i_5_reg[8]  ( .D(n42077), .CP(clk), .Q(
        \shifter_0/reg_i_5 [8]) );
  dff_sg \shifter_0/reg_i_5_reg[9]  ( .D(n42078), .CP(clk), .Q(
        \shifter_0/reg_i_5 [9]) );
  dff_sg \shifter_0/reg_i_5_reg[10]  ( .D(n42074), .CP(clk), .Q(
        \shifter_0/reg_i_5 [10]) );
  dff_sg \shifter_0/reg_i_5_reg[11]  ( .D(n42075), .CP(clk), .Q(
        \shifter_0/reg_i_5 [11]) );
  dff_sg \shifter_0/reg_i_5_reg[12]  ( .D(n42083), .CP(clk), .Q(
        \shifter_0/reg_i_5 [12]) );
  dff_sg \shifter_0/reg_i_5_reg[13]  ( .D(n42084), .CP(clk), .Q(
        \shifter_0/reg_i_5 [13]) );
  dff_sg \shifter_0/reg_i_5_reg[14]  ( .D(n42080), .CP(clk), .Q(
        \shifter_0/reg_i_5 [14]) );
  dff_sg \shifter_0/reg_i_5_reg[15]  ( .D(n42081), .CP(clk), .Q(
        \shifter_0/reg_i_5 [15]) );
  dff_sg \shifter_0/reg_i_5_reg[16]  ( .D(n42065), .CP(clk), .Q(
        \shifter_0/reg_i_5 [16]) );
  dff_sg \shifter_0/reg_i_5_reg[17]  ( .D(n42066), .CP(clk), .Q(
        \shifter_0/reg_i_5 [17]) );
  dff_sg \shifter_0/reg_i_5_reg[18]  ( .D(n42062), .CP(clk), .Q(
        \shifter_0/reg_i_5 [18]) );
  dff_sg \shifter_0/reg_i_5_reg[19]  ( .D(n42063), .CP(clk), .Q(
        \shifter_0/reg_i_5 [19]) );
  dff_sg \shifter_0/reg_i_6_reg[0]  ( .D(n42071), .CP(clk), .Q(
        \shifter_0/reg_i_6 [0]) );
  dff_sg \shifter_0/reg_i_6_reg[1]  ( .D(n42072), .CP(clk), .Q(
        \shifter_0/reg_i_6 [1]) );
  dff_sg \shifter_0/reg_i_6_reg[2]  ( .D(n42068), .CP(clk), .Q(
        \shifter_0/reg_i_6 [2]) );
  dff_sg \shifter_0/reg_i_6_reg[3]  ( .D(n42069), .CP(clk), .Q(
        \shifter_0/reg_i_6 [3]) );
  dff_sg \shifter_0/reg_i_6_reg[4]  ( .D(n42101), .CP(clk), .Q(
        \shifter_0/reg_i_6 [4]) );
  dff_sg \shifter_0/reg_i_6_reg[5]  ( .D(n42102), .CP(clk), .Q(
        \shifter_0/reg_i_6 [5]) );
  dff_sg \shifter_0/reg_i_6_reg[6]  ( .D(n42098), .CP(clk), .Q(
        \shifter_0/reg_i_6 [6]) );
  dff_sg \shifter_0/reg_i_6_reg[7]  ( .D(n42099), .CP(clk), .Q(
        \shifter_0/reg_i_6 [7]) );
  dff_sg \shifter_0/reg_i_6_reg[8]  ( .D(n42107), .CP(clk), .Q(
        \shifter_0/reg_i_6 [8]) );
  dff_sg \shifter_0/reg_i_6_reg[9]  ( .D(n42108), .CP(clk), .Q(
        \shifter_0/reg_i_6 [9]) );
  dff_sg \shifter_0/reg_i_6_reg[10]  ( .D(n42104), .CP(clk), .Q(
        \shifter_0/reg_i_6 [10]) );
  dff_sg \shifter_0/reg_i_6_reg[11]  ( .D(n42105), .CP(clk), .Q(
        \shifter_0/reg_i_6 [11]) );
  dff_sg \shifter_0/reg_i_6_reg[12]  ( .D(n42089), .CP(clk), .Q(
        \shifter_0/reg_i_6 [12]) );
  dff_sg \shifter_0/reg_i_6_reg[13]  ( .D(n42090), .CP(clk), .Q(
        \shifter_0/reg_i_6 [13]) );
  dff_sg \shifter_0/reg_i_6_reg[14]  ( .D(n42086), .CP(clk), .Q(
        \shifter_0/reg_i_6 [14]) );
  dff_sg \shifter_0/reg_i_6_reg[15]  ( .D(n42087), .CP(clk), .Q(
        \shifter_0/reg_i_6 [15]) );
  dff_sg \shifter_0/reg_i_6_reg[16]  ( .D(n42095), .CP(clk), .Q(
        \shifter_0/reg_i_6 [16]) );
  dff_sg \shifter_0/reg_i_6_reg[17]  ( .D(n42096), .CP(clk), .Q(
        \shifter_0/reg_i_6 [17]) );
  dff_sg \shifter_0/reg_i_6_reg[18]  ( .D(n42092), .CP(clk), .Q(
        \shifter_0/reg_i_6 [18]) );
  dff_sg \shifter_0/reg_i_6_reg[19]  ( .D(n42093), .CP(clk), .Q(
        \shifter_0/reg_i_6 [19]) );
  dff_sg \shifter_0/reg_i_7_reg[0]  ( .D(n42029), .CP(clk), .Q(
        \shifter_0/reg_i_7 [0]) );
  dff_sg \shifter_0/reg_i_7_reg[1]  ( .D(n42030), .CP(clk), .Q(
        \shifter_0/reg_i_7 [1]) );
  dff_sg \shifter_0/reg_i_7_reg[2]  ( .D(n42026), .CP(clk), .Q(
        \shifter_0/reg_i_7 [2]) );
  dff_sg \shifter_0/reg_i_7_reg[3]  ( .D(n42027), .CP(clk), .Q(
        \shifter_0/reg_i_7 [3]) );
  dff_sg \shifter_0/reg_i_7_reg[4]  ( .D(n42035), .CP(clk), .Q(
        \shifter_0/reg_i_7 [4]) );
  dff_sg \shifter_0/reg_i_7_reg[5]  ( .D(n42036), .CP(clk), .Q(
        \shifter_0/reg_i_7 [5]) );
  dff_sg \shifter_0/reg_i_7_reg[6]  ( .D(n42032), .CP(clk), .Q(
        \shifter_0/reg_i_7 [6]) );
  dff_sg \shifter_0/reg_i_7_reg[7]  ( .D(n42033), .CP(clk), .Q(
        \shifter_0/reg_i_7 [7]) );
  dff_sg \shifter_0/reg_i_7_reg[8]  ( .D(n42017), .CP(clk), .Q(
        \shifter_0/reg_i_7 [8]) );
  dff_sg \shifter_0/reg_i_7_reg[9]  ( .D(n42018), .CP(clk), .Q(
        \shifter_0/reg_i_7 [9]) );
  dff_sg \shifter_0/reg_i_7_reg[10]  ( .D(n42014), .CP(clk), .Q(
        \shifter_0/reg_i_7 [10]) );
  dff_sg \shifter_0/reg_i_7_reg[11]  ( .D(n42015), .CP(clk), .Q(
        \shifter_0/reg_i_7 [11]) );
  dff_sg \shifter_0/reg_i_7_reg[12]  ( .D(n42023), .CP(clk), .Q(
        \shifter_0/reg_i_7 [12]) );
  dff_sg \shifter_0/reg_i_7_reg[13]  ( .D(n42024), .CP(clk), .Q(
        \shifter_0/reg_i_7 [13]) );
  dff_sg \shifter_0/reg_i_7_reg[14]  ( .D(n42020), .CP(clk), .Q(
        \shifter_0/reg_i_7 [14]) );
  dff_sg \shifter_0/reg_i_7_reg[15]  ( .D(n42021), .CP(clk), .Q(
        \shifter_0/reg_i_7 [15]) );
  dff_sg \shifter_0/reg_i_7_reg[16]  ( .D(n42053), .CP(clk), .Q(
        \shifter_0/reg_i_7 [16]) );
  dff_sg \shifter_0/reg_i_7_reg[17]  ( .D(n42054), .CP(clk), .Q(
        \shifter_0/reg_i_7 [17]) );
  dff_sg \shifter_0/reg_i_7_reg[18]  ( .D(n42050), .CP(clk), .Q(
        \shifter_0/reg_i_7 [18]) );
  dff_sg \shifter_0/reg_i_7_reg[19]  ( .D(n42051), .CP(clk), .Q(
        \shifter_0/reg_i_7 [19]) );
  dff_sg \shifter_0/reg_i_8_reg[0]  ( .D(n42059), .CP(clk), .Q(
        \shifter_0/reg_i_8 [0]) );
  dff_sg \shifter_0/reg_i_8_reg[1]  ( .D(n42060), .CP(clk), .Q(
        \shifter_0/reg_i_8 [1]) );
  dff_sg \shifter_0/reg_i_8_reg[2]  ( .D(n42056), .CP(clk), .Q(
        \shifter_0/reg_i_8 [2]) );
  dff_sg \shifter_0/reg_i_8_reg[3]  ( .D(n42057), .CP(clk), .Q(
        \shifter_0/reg_i_8 [3]) );
  dff_sg \shifter_0/reg_i_8_reg[4]  ( .D(n42041), .CP(clk), .Q(
        \shifter_0/reg_i_8 [4]) );
  dff_sg \shifter_0/reg_i_8_reg[5]  ( .D(n42042), .CP(clk), .Q(
        \shifter_0/reg_i_8 [5]) );
  dff_sg \shifter_0/reg_i_8_reg[6]  ( .D(n42038), .CP(clk), .Q(
        \shifter_0/reg_i_8 [6]) );
  dff_sg \shifter_0/reg_i_8_reg[7]  ( .D(n42039), .CP(clk), .Q(
        \shifter_0/reg_i_8 [7]) );
  dff_sg \shifter_0/reg_i_8_reg[8]  ( .D(n42047), .CP(clk), .Q(
        \shifter_0/reg_i_8 [8]) );
  dff_sg \shifter_0/reg_i_8_reg[9]  ( .D(n42048), .CP(clk), .Q(
        \shifter_0/reg_i_8 [9]) );
  dff_sg \shifter_0/reg_i_8_reg[10]  ( .D(n42044), .CP(clk), .Q(
        \shifter_0/reg_i_8 [10]) );
  dff_sg \shifter_0/reg_i_8_reg[11]  ( .D(n42045), .CP(clk), .Q(
        \shifter_0/reg_i_8 [11]) );
  dff_sg \shifter_0/reg_i_8_reg[12]  ( .D(n41563), .CP(clk), .Q(
        \shifter_0/reg_i_8 [12]) );
  dff_sg \shifter_0/reg_i_8_reg[13]  ( .D(n41569), .CP(clk), .Q(
        \shifter_0/reg_i_8 [13]) );
  dff_sg \shifter_0/reg_i_8_reg[14]  ( .D(n41575), .CP(clk), .Q(
        \shifter_0/reg_i_8 [14]) );
  dff_sg \shifter_0/reg_i_8_reg[15]  ( .D(n41581), .CP(clk), .Q(
        \shifter_0/reg_i_8 [15]) );
  dff_sg \shifter_0/reg_i_8_reg[16]  ( .D(n41551), .CP(clk), .Q(
        \shifter_0/reg_i_8 [16]) );
  dff_sg \shifter_0/reg_i_8_reg[17]  ( .D(n41771), .CP(clk), .Q(
        \shifter_0/reg_i_8 [17]) );
  dff_sg \shifter_0/reg_i_8_reg[18]  ( .D(n41557), .CP(clk), .Q(
        \shifter_0/reg_i_8 [18]) );
  dff_sg \shifter_0/reg_i_8_reg[19]  ( .D(n41584), .CP(clk), .Q(
        \shifter_0/reg_i_8 [19]) );
  dff_sg \shifter_0/reg_i_9_reg[0]  ( .D(n41828), .CP(clk), .Q(
        \shifter_0/reg_i_9 [0]) );
  dff_sg \shifter_0/reg_i_9_reg[1]  ( .D(n41907), .CP(clk), .Q(
        \shifter_0/reg_i_9 [1]) );
  dff_sg \shifter_0/reg_i_9_reg[2]  ( .D(n41539), .CP(clk), .Q(
        \shifter_0/reg_i_9 [2]) );
  dff_sg \shifter_0/reg_i_9_reg[3]  ( .D(n41523), .CP(clk), .Q(
        \shifter_0/reg_i_9 [3]) );
  dff_sg \shifter_0/reg_i_9_reg[4]  ( .D(n42110), .CP(clk), .Q(
        \shifter_0/reg_i_9 [4]) );
  dff_sg \shifter_0/reg_i_9_reg[5]  ( .D(n41904), .CP(clk), .Q(
        \shifter_0/reg_i_9 [5]) );
  dff_sg \shifter_0/reg_i_9_reg[6]  ( .D(n41587), .CP(clk), .Q(
        \shifter_0/reg_i_9 [6]) );
  dff_sg \shifter_0/reg_i_9_reg[7]  ( .D(n41590), .CP(clk), .Q(
        \shifter_0/reg_i_9 [7]) );
  dff_sg \shifter_0/reg_i_9_reg[8]  ( .D(n41859), .CP(clk), .Q(
        \shifter_0/reg_i_9 [8]) );
  dff_sg \shifter_0/reg_i_9_reg[9]  ( .D(n41862), .CP(clk), .Q(
        \shifter_0/reg_i_9 [9]) );
  dff_sg \shifter_0/reg_i_9_reg[10]  ( .D(n41566), .CP(clk), .Q(
        \shifter_0/reg_i_9 [10]) );
  dff_sg \shifter_0/reg_i_9_reg[11]  ( .D(n41544), .CP(clk), .Q(
        \shifter_0/reg_i_9 [11]) );
  dff_sg \shifter_0/reg_i_9_reg[12]  ( .D(n41553), .CP(clk), .Q(
        \shifter_0/reg_i_9 [12]) );
  dff_sg \shifter_0/reg_i_9_reg[13]  ( .D(n41841), .CP(clk), .Q(
        \shifter_0/reg_i_9 [13]) );
  dff_sg \shifter_0/reg_i_9_reg[14]  ( .D(n41840), .CP(clk), .Q(
        \shifter_0/reg_i_9 [14]) );
  dff_sg \shifter_0/reg_i_9_reg[15]  ( .D(n41847), .CP(clk), .Q(
        \shifter_0/reg_i_9 [15]) );
  dff_sg \shifter_0/reg_i_9_reg[16]  ( .D(n41554), .CP(clk), .Q(
        \shifter_0/reg_i_9 [16]) );
  dff_sg \shifter_0/reg_i_9_reg[17]  ( .D(n41578), .CP(clk), .Q(
        \shifter_0/reg_i_9 [17]) );
  dff_sg \shifter_0/reg_i_9_reg[18]  ( .D(n41883), .CP(clk), .Q(
        \shifter_0/reg_i_9 [18]) );
  dff_sg \shifter_0/reg_i_9_reg[19]  ( .D(n41732), .CP(clk), .Q(
        \shifter_0/reg_i_9 [19]) );
  dff_sg \shifter_0/reg_i_10_reg[0]  ( .D(n41596), .CP(clk), .Q(
        \shifter_0/reg_i_10 [0]) );
  dff_sg \shifter_0/reg_i_10_reg[1]  ( .D(n41599), .CP(clk), .Q(
        \shifter_0/reg_i_10 [1]) );
  dff_sg \shifter_0/reg_i_10_reg[2]  ( .D(n41605), .CP(clk), .Q(
        \shifter_0/reg_i_10 [2]) );
  dff_sg \shifter_0/reg_i_10_reg[3]  ( .D(n41819), .CP(clk), .Q(
        \shifter_0/reg_i_10 [3]) );
  dff_sg \shifter_0/reg_i_10_reg[4]  ( .D(n41747), .CP(clk), .Q(
        \shifter_0/reg_i_10 [4]) );
  dff_sg \shifter_0/reg_i_10_reg[5]  ( .D(n41898), .CP(clk), .Q(
        \shifter_0/reg_i_10 [5]) );
  dff_sg \shifter_0/reg_i_10_reg[6]  ( .D(n41550), .CP(clk), .Q(
        \shifter_0/reg_i_10 [6]) );
  dff_sg \shifter_0/reg_i_10_reg[7]  ( .D(n41789), .CP(clk), .Q(
        \shifter_0/reg_i_10 [7]) );
  dff_sg \shifter_0/reg_i_10_reg[8]  ( .D(n41765), .CP(clk), .Q(
        \shifter_0/reg_i_10 [8]) );
  dff_sg \shifter_0/reg_i_10_reg[9]  ( .D(n41768), .CP(clk), .Q(
        \shifter_0/reg_i_10 [9]) );
  dff_sg \shifter_0/reg_i_10_reg[10]  ( .D(n41543), .CP(clk), .Q(
        \shifter_0/reg_i_10 [10]) );
  dff_sg \shifter_0/reg_i_10_reg[11]  ( .D(n41844), .CP(clk), .Q(
        \shifter_0/reg_i_10 [11]) );
  dff_sg \shifter_0/reg_i_10_reg[12]  ( .D(n41623), .CP(clk), .Q(
        \shifter_0/reg_i_10 [12]) );
  dff_sg \shifter_0/reg_i_10_reg[13]  ( .D(n41629), .CP(clk), .Q(
        \shifter_0/reg_i_10 [13]) );
  dff_sg \shifter_0/reg_i_10_reg[14]  ( .D(n41780), .CP(clk), .Q(
        \shifter_0/reg_i_10 [14]) );
  dff_sg \shifter_0/reg_i_10_reg[15]  ( .D(n41774), .CP(clk), .Q(
        \shifter_0/reg_i_10 [15]) );
  dff_sg \shifter_0/reg_i_10_reg[16]  ( .D(n41738), .CP(clk), .Q(
        \shifter_0/reg_i_10 [16]) );
  dff_sg \shifter_0/reg_i_10_reg[17]  ( .D(n41602), .CP(clk), .Q(
        \shifter_0/reg_i_10 [17]) );
  dff_sg \shifter_0/reg_i_10_reg[18]  ( .D(n41762), .CP(clk), .Q(
        \shifter_0/reg_i_10 [18]) );
  dff_sg \shifter_0/reg_i_10_reg[19]  ( .D(n41756), .CP(clk), .Q(
        \shifter_0/reg_i_10 [19]) );
  dff_sg \shifter_0/reg_i_11_reg[0]  ( .D(n41783), .CP(clk), .Q(
        \shifter_0/reg_i_11 [0]) );
  dff_sg \shifter_0/reg_i_11_reg[1]  ( .D(n41792), .CP(clk), .Q(
        \shifter_0/reg_i_11 [1]) );
  dff_sg \shifter_0/reg_i_11_reg[2]  ( .D(n41786), .CP(clk), .Q(
        \shifter_0/reg_i_11 [2]) );
  dff_sg \shifter_0/reg_i_11_reg[3]  ( .D(n41735), .CP(clk), .Q(
        \shifter_0/reg_i_11 [3]) );
  dff_sg \shifter_0/reg_i_11_reg[4]  ( .D(n41560), .CP(clk), .Q(
        \shifter_0/reg_i_11 [4]) );
  dff_sg \shifter_0/reg_i_11_reg[5]  ( .D(n41538), .CP(clk), .Q(
        \shifter_0/reg_i_11 [5]) );
  dff_sg \shifter_0/reg_i_11_reg[6]  ( .D(n41853), .CP(clk), .Q(
        \shifter_0/reg_i_11 [6]) );
  dff_sg \shifter_0/reg_i_11_reg[7]  ( .D(n41525), .CP(clk), .Q(
        \shifter_0/reg_i_11 [7]) );
  dff_sg \shifter_0/reg_i_11_reg[8]  ( .D(n41795), .CP(clk), .Q(
        \shifter_0/reg_i_11 [8]) );
  dff_sg \shifter_0/reg_i_11_reg[9]  ( .D(n41695), .CP(clk), .Q(
        \shifter_0/reg_i_11 [9]) );
  dff_sg \shifter_0/reg_i_11_reg[10]  ( .D(n41547), .CP(clk), .Q(
        \shifter_0/reg_i_11 [10]) );
  dff_sg \shifter_0/reg_i_11_reg[11]  ( .D(n41548), .CP(clk), .Q(
        \shifter_0/reg_i_11 [11]) );
  dff_sg \shifter_0/reg_i_11_reg[12]  ( .D(n41753), .CP(clk), .Q(
        \shifter_0/reg_i_11 [12]) );
  dff_sg \shifter_0/reg_i_11_reg[13]  ( .D(n41635), .CP(clk), .Q(
        \shifter_0/reg_i_11 [13]) );
  dff_sg \shifter_0/reg_i_11_reg[14]  ( .D(n41653), .CP(clk), .Q(
        \shifter_0/reg_i_11 [14]) );
  dff_sg \shifter_0/reg_i_11_reg[15]  ( .D(n41665), .CP(clk), .Q(
        \shifter_0/reg_i_11 [15]) );
  dff_sg \shifter_0/reg_i_11_reg[16]  ( .D(n41585), .CP(clk), .Q(
        \shifter_0/reg_i_11 [16]) );
  dff_sg \shifter_0/reg_i_11_reg[17]  ( .D(n41586), .CP(clk), .Q(
        \shifter_0/reg_i_11 [17]) );
  dff_sg \shifter_0/reg_i_11_reg[18]  ( .D(n41582), .CP(clk), .Q(
        \shifter_0/reg_i_11 [18]) );
  dff_sg \shifter_0/reg_i_11_reg[19]  ( .D(n41583), .CP(clk), .Q(
        \shifter_0/reg_i_11 [19]) );
  dff_sg \shifter_0/reg_i_12_reg[0]  ( .D(n41591), .CP(clk), .Q(
        \shifter_0/reg_i_12 [0]) );
  dff_sg \shifter_0/reg_i_12_reg[1]  ( .D(n41592), .CP(clk), .Q(
        \shifter_0/reg_i_12 [1]) );
  dff_sg \shifter_0/reg_i_12_reg[2]  ( .D(n41588), .CP(clk), .Q(
        \shifter_0/reg_i_12 [2]) );
  dff_sg \shifter_0/reg_i_12_reg[3]  ( .D(n41589), .CP(clk), .Q(
        \shifter_0/reg_i_12 [3]) );
  dff_sg \shifter_0/reg_i_12_reg[4]  ( .D(n41573), .CP(clk), .Q(
        \shifter_0/reg_i_12 [4]) );
  dff_sg \shifter_0/reg_i_12_reg[5]  ( .D(n41574), .CP(clk), .Q(
        \shifter_0/reg_i_12 [5]) );
  dff_sg \shifter_0/reg_i_12_reg[6]  ( .D(n41570), .CP(clk), .Q(
        \shifter_0/reg_i_12 [6]) );
  dff_sg \shifter_0/reg_i_12_reg[7]  ( .D(n41571), .CP(clk), .Q(
        \shifter_0/reg_i_12 [7]) );
  dff_sg \shifter_0/reg_i_12_reg[8]  ( .D(n41579), .CP(clk), .Q(
        \shifter_0/reg_i_12 [8]) );
  dff_sg \shifter_0/reg_i_12_reg[9]  ( .D(n41580), .CP(clk), .Q(
        \shifter_0/reg_i_12 [9]) );
  dff_sg \shifter_0/reg_i_12_reg[10]  ( .D(n41576), .CP(clk), .Q(
        \shifter_0/reg_i_12 [10]) );
  dff_sg \shifter_0/reg_i_12_reg[11]  ( .D(n41577), .CP(clk), .Q(
        \shifter_0/reg_i_12 [11]) );
  dff_sg \shifter_0/reg_i_12_reg[12]  ( .D(n41825), .CP(clk), .Q(
        \shifter_0/reg_i_12 [12]) );
  dff_sg \shifter_0/reg_i_12_reg[13]  ( .D(n41822), .CP(clk), .Q(
        \shifter_0/reg_i_12 [13]) );
  dff_sg \shifter_0/reg_i_12_reg[14]  ( .D(n41606), .CP(clk), .Q(
        \shifter_0/reg_i_12 [14]) );
  dff_sg \shifter_0/reg_i_12_reg[15]  ( .D(n41816), .CP(clk), .Q(
        \shifter_0/reg_i_12 [15]) );
  dff_sg \shifter_0/reg_i_12_reg[16]  ( .D(n41555), .CP(clk), .Q(
        \shifter_0/reg_i_12 [16]) );
  dff_sg \shifter_0/reg_i_12_reg[17]  ( .D(n41810), .CP(clk), .Q(
        \shifter_0/reg_i_12 [17]) );
  dff_sg \shifter_0/reg_i_12_reg[18]  ( .D(n41813), .CP(clk), .Q(
        \shifter_0/reg_i_12 [18]) );
  dff_sg \shifter_0/reg_i_12_reg[19]  ( .D(n41607), .CP(clk), .Q(
        \shifter_0/reg_i_12 [19]) );
  dff_sg \shifter_0/reg_i_13_reg[0]  ( .D(n41597), .CP(clk), .Q(
        \shifter_0/reg_i_13 [0]) );
  dff_sg \shifter_0/reg_i_13_reg[1]  ( .D(n41598), .CP(clk), .Q(
        \shifter_0/reg_i_13 [1]) );
  dff_sg \shifter_0/reg_i_13_reg[2]  ( .D(n41594), .CP(clk), .Q(
        \shifter_0/reg_i_13 [2]) );
  dff_sg \shifter_0/reg_i_13_reg[3]  ( .D(n41595), .CP(clk), .Q(
        \shifter_0/reg_i_13 [3]) );
  dff_sg \shifter_0/reg_i_13_reg[4]  ( .D(n41603), .CP(clk), .Q(
        \shifter_0/reg_i_13 [4]) );
  dff_sg \shifter_0/reg_i_13_reg[5]  ( .D(n41604), .CP(clk), .Q(
        \shifter_0/reg_i_13 [5]) );
  dff_sg \shifter_0/reg_i_13_reg[6]  ( .D(n41600), .CP(clk), .Q(
        \shifter_0/reg_i_13 [6]) );
  dff_sg \shifter_0/reg_i_13_reg[7]  ( .D(n41601), .CP(clk), .Q(
        \shifter_0/reg_i_13 [7]) );
  dff_sg \shifter_0/reg_i_13_reg[8]  ( .D(n41889), .CP(clk), .Q(
        \shifter_0/reg_i_13 [8]) );
  dff_sg \shifter_0/reg_i_13_reg[9]  ( .D(n41892), .CP(clk), .Q(
        \shifter_0/reg_i_13 [9]) );
  dff_sg \shifter_0/reg_i_13_reg[10]  ( .D(n41901), .CP(clk), .Q(
        \shifter_0/reg_i_13 [10]) );
  dff_sg \shifter_0/reg_i_13_reg[11]  ( .D(n41895), .CP(clk), .Q(
        \shifter_0/reg_i_13 [11]) );
  dff_sg \shifter_0/reg_i_13_reg[12]  ( .D(n41545), .CP(clk), .Q(
        \shifter_0/reg_i_13 [12]) );
  dff_sg \shifter_0/reg_i_13_reg[13]  ( .D(n41546), .CP(clk), .Q(
        \shifter_0/reg_i_13 [13]) );
  dff_sg \shifter_0/reg_i_13_reg[14]  ( .D(n41877), .CP(clk), .Q(
        \shifter_0/reg_i_13 [14]) );
  dff_sg \shifter_0/reg_i_13_reg[15]  ( .D(n41880), .CP(clk), .Q(
        \shifter_0/reg_i_13 [15]) );
  dff_sg \shifter_0/reg_i_13_reg[16]  ( .D(n41913), .CP(clk), .Q(
        \shifter_0/reg_i_13 [16]) );
  dff_sg \shifter_0/reg_i_13_reg[17]  ( .D(n41807), .CP(clk), .Q(
        \shifter_0/reg_i_13 [17]) );
  dff_sg \shifter_0/reg_i_13_reg[18]  ( .D(n41837), .CP(clk), .Q(
        \shifter_0/reg_i_13 [18]) );
  dff_sg \shifter_0/reg_i_13_reg[19]  ( .D(n41834), .CP(clk), .Q(
        \shifter_0/reg_i_13 [19]) );
  dff_sg \shifter_0/reg_i_14_reg[0]  ( .D(n41865), .CP(clk), .Q(
        \shifter_0/reg_i_14 [0]) );
  dff_sg \shifter_0/reg_i_14_reg[1]  ( .D(n41868), .CP(clk), .Q(
        \shifter_0/reg_i_14 [1]) );
  dff_sg \shifter_0/reg_i_14_reg[2]  ( .D(n41524), .CP(clk), .Q(
        \shifter_0/reg_i_14 [2]) );
  dff_sg \shifter_0/reg_i_14_reg[3]  ( .D(n41874), .CP(clk), .Q(
        \shifter_0/reg_i_14 [3]) );
  dff_sg \shifter_0/reg_i_14_reg[4]  ( .D(n41561), .CP(clk), .Q(
        \shifter_0/reg_i_14 [4]) );
  dff_sg \shifter_0/reg_i_14_reg[5]  ( .D(n41562), .CP(clk), .Q(
        \shifter_0/reg_i_14 [5]) );
  dff_sg \shifter_0/reg_i_14_reg[6]  ( .D(n41558), .CP(clk), .Q(
        \shifter_0/reg_i_14 [6]) );
  dff_sg \shifter_0/reg_i_14_reg[7]  ( .D(n41559), .CP(clk), .Q(
        \shifter_0/reg_i_14 [7]) );
  dff_sg \shifter_0/reg_i_14_reg[8]  ( .D(n41567), .CP(clk), .Q(
        \shifter_0/reg_i_14 [8]) );
  dff_sg \shifter_0/reg_i_14_reg[9]  ( .D(n41568), .CP(clk), .Q(
        \shifter_0/reg_i_14 [9]) );
  dff_sg \shifter_0/reg_i_14_reg[10]  ( .D(n41564), .CP(clk), .Q(
        \shifter_0/reg_i_14 [10]) );
  dff_sg \shifter_0/reg_i_14_reg[11]  ( .D(n41565), .CP(clk), .Q(
        \shifter_0/reg_i_14 [11]) );
  dff_sg \shifter_0/reg_i_14_reg[12]  ( .D(n41705), .CP(clk), .Q(
        \shifter_0/reg_i_14 [12]) );
  dff_sg \shifter_0/reg_i_14_reg[13]  ( .D(n41706), .CP(clk), .Q(
        \shifter_0/reg_i_14 [13]) );
  dff_sg \shifter_0/reg_i_14_reg[14]  ( .D(n42111), .CP(clk), .Q(
        \shifter_0/reg_i_14 [14]) );
  dff_sg \shifter_0/reg_i_14_reg[15]  ( .D(n42112), .CP(clk), .Q(
        \shifter_0/reg_i_14 [15]) );
  dff_sg \shifter_0/reg_i_14_reg[16]  ( .D(n41744), .CP(clk), .Q(
        \shifter_0/reg_i_14 [16]) );
  dff_sg \shifter_0/reg_i_14_reg[17]  ( .D(n41750), .CP(clk), .Q(
        \shifter_0/reg_i_14 [17]) );
  dff_sg \shifter_0/reg_i_14_reg[18]  ( .D(n41521), .CP(clk), .Q(
        \shifter_0/reg_i_14 [18]) );
  dff_sg \shifter_0/reg_i_14_reg[19]  ( .D(n41556), .CP(clk), .Q(
        \shifter_0/reg_i_14 [19]) );
  dff_sg \shifter_0/reg_i_15_reg[0]  ( .D(n41929), .CP(clk), .Q(
        \shifter_0/reg_i_15 [0]) );
  dff_sg \shifter_0/reg_i_15_reg[1]  ( .D(n42100), .CP(clk), .Q(
        \shifter_0/reg_i_15 [1]) );
  dff_sg \shifter_0/reg_i_15_reg[2]  ( .D(n42043), .CP(clk), .Q(
        \shifter_0/reg_i_15 [2]) );
  dff_sg \shifter_0/reg_i_15_reg[3]  ( .D(n42088), .CP(clk), .Q(
        \shifter_0/reg_i_15 [3]) );
  dff_sg \shifter_0/reg_i_15_reg[4]  ( .D(n41529), .CP(clk), .Q(
        \shifter_0/reg_i_15 [4]) );
  dff_sg \shifter_0/reg_i_15_reg[5]  ( .D(n42067), .CP(clk), .Q(
        \shifter_0/reg_i_15 [5]) );
  dff_sg \shifter_0/reg_i_15_reg[6]  ( .D(n42106), .CP(clk), .Q(
        \shifter_0/reg_i_15 [6]) );
  dff_sg \shifter_0/reg_i_15_reg[7]  ( .D(n42016), .CP(clk), .Q(
        \shifter_0/reg_i_15 [7]) );
  dff_sg \shifter_0/reg_i_15_reg[8]  ( .D(n42055), .CP(clk), .Q(
        \shifter_0/reg_i_15 [8]) );
  dff_sg \shifter_0/reg_i_15_reg[9]  ( .D(n42058), .CP(clk), .Q(
        \shifter_0/reg_i_15 [9]) );
  dff_sg \shifter_0/reg_i_15_reg[10]  ( .D(n42064), .CP(clk), .Q(
        \shifter_0/reg_i_15 [10]) );
  dff_sg \shifter_0/reg_i_15_reg[11]  ( .D(n42073), .CP(clk), .Q(
        \shifter_0/reg_i_15 [11]) );
  dff_sg \shifter_0/reg_i_15_reg[12]  ( .D(n41932), .CP(clk), .Q(
        \shifter_0/reg_i_15 [12]) );
  dff_sg \shifter_0/reg_i_15_reg[13]  ( .D(n41938), .CP(clk), .Q(
        \shifter_0/reg_i_15 [13]) );
  dff_sg \shifter_0/reg_i_15_reg[14]  ( .D(n41534), .CP(clk), .Q(
        \shifter_0/reg_i_15 [14]) );
  dff_sg \shifter_0/reg_i_15_reg[15]  ( .D(n41533), .CP(clk), .Q(
        \shifter_0/reg_i_15 [15]) );
  dff_sg \shifter_0/reg_i_15_reg[16]  ( .D(n42097), .CP(clk), .Q(
        \shifter_0/reg_i_15 [16]) );
  dff_sg \shifter_0/reg_i_15_reg[17]  ( .D(n41965), .CP(clk), .Q(
        \shifter_0/reg_i_15 [17]) );
  dff_sg \shifter_0/reg_i_15_reg[18]  ( .D(n42025), .CP(clk), .Q(
        \shifter_0/reg_i_15 [18]) );
  dff_sg \shifter_0/reg_i_15_reg[19]  ( .D(n41977), .CP(clk), .Q(
        \shifter_0/reg_i_15 [19]) );
  dff_sg \shifter_0/reg_w_0_reg[0]  ( .D(n42022), .CP(clk), .Q(
        \shifter_0/reg_w_0 [0]) );
  dff_sg \shifter_0/reg_w_0_reg[1]  ( .D(n42034), .CP(clk), .Q(
        \shifter_0/reg_w_0 [1]) );
  dff_sg \shifter_0/reg_w_0_reg[2]  ( .D(n42046), .CP(clk), .Q(
        \shifter_0/reg_w_0 [2]) );
  dff_sg \shifter_0/reg_w_0_reg[3]  ( .D(n42076), .CP(clk), .Q(
        \shifter_0/reg_w_0 [3]) );
  dff_sg \shifter_0/reg_w_0_reg[4]  ( .D(n41986), .CP(clk), .Q(
        \shifter_0/reg_w_0 [4]) );
  dff_sg \shifter_0/reg_w_0_reg[5]  ( .D(n42091), .CP(clk), .Q(
        \shifter_0/reg_w_0 [5]) );
  dff_sg \shifter_0/reg_w_0_reg[6]  ( .D(n41536), .CP(clk), .Q(
        \shifter_0/reg_w_0 [6]) );
  dff_sg \shifter_0/reg_w_0_reg[7]  ( .D(n42094), .CP(clk), .Q(
        \shifter_0/reg_w_0 [7]) );
  dff_sg \shifter_0/reg_w_0_reg[8]  ( .D(n41968), .CP(clk), .Q(
        \shifter_0/reg_w_0 [8]) );
  dff_sg \shifter_0/reg_w_0_reg[9]  ( .D(n41971), .CP(clk), .Q(
        \shifter_0/reg_w_0 [9]) );
  dff_sg \shifter_0/reg_w_0_reg[10]  ( .D(n42082), .CP(clk), .Q(
        \shifter_0/reg_w_0 [10]) );
  dff_sg \shifter_0/reg_w_0_reg[11]  ( .D(n41974), .CP(clk), .Q(
        \shifter_0/reg_w_0 [11]) );
  dff_sg \shifter_0/reg_w_0_reg[12]  ( .D(n42119), .CP(clk), .Q(
        \shifter_0/reg_w_0 [12]) );
  dff_sg \shifter_0/reg_w_0_reg[13]  ( .D(n42122), .CP(clk), .Q(
        \shifter_0/reg_w_0 [13]) );
  dff_sg \shifter_0/reg_w_0_reg[14]  ( .D(n42137), .CP(clk), .Q(
        \shifter_0/reg_w_0 [14]) );
  dff_sg \shifter_0/reg_w_0_reg[15]  ( .D(n42140), .CP(clk), .Q(
        \shifter_0/reg_w_0 [15]) );
  dff_sg \shifter_0/reg_w_0_reg[16]  ( .D(n41959), .CP(clk), .Q(
        \shifter_0/reg_w_0 [16]) );
  dff_sg \shifter_0/reg_w_0_reg[17]  ( .D(n41956), .CP(clk), .Q(
        \shifter_0/reg_w_0 [17]) );
  dff_sg \shifter_0/reg_w_0_reg[18]  ( .D(n41522), .CP(clk), .Q(
        \shifter_0/reg_w_0 [18]) );
  dff_sg \shifter_0/reg_w_0_reg[19]  ( .D(n41711), .CP(clk), .Q(
        \shifter_0/reg_w_0 [19]) );
  dff_sg \shifter_0/reg_w_1_reg[0]  ( .D(n41717), .CP(clk), .Q(
        \shifter_0/reg_w_1 [0]) );
  dff_sg \shifter_0/reg_w_1_reg[1]  ( .D(n41720), .CP(clk), .Q(
        \shifter_0/reg_w_1 [1]) );
  dff_sg \shifter_0/reg_w_1_reg[2]  ( .D(n42116), .CP(clk), .Q(
        \shifter_0/reg_w_1 [2]) );
  dff_sg \shifter_0/reg_w_1_reg[3]  ( .D(n42143), .CP(clk), .Q(
        \shifter_0/reg_w_1 [3]) );
  dff_sg \shifter_0/reg_w_1_reg[4]  ( .D(n42155), .CP(clk), .Q(
        \shifter_0/reg_w_1 [4]) );
  dff_sg \shifter_0/reg_w_1_reg[5]  ( .D(n41920), .CP(clk), .Q(
        \shifter_0/reg_w_1 [5]) );
  dff_sg \shifter_0/reg_w_1_reg[6]  ( .D(n41708), .CP(clk), .Q(
        \shifter_0/reg_w_1 [6]) );
  dff_sg \shifter_0/reg_w_1_reg[7]  ( .D(n41729), .CP(clk), .Q(
        \shifter_0/reg_w_1 [7]) );
  dff_sg \shifter_0/reg_w_1_reg[8]  ( .D(n42079), .CP(clk), .Q(
        \shifter_0/reg_w_1 [8]) );
  dff_sg \shifter_0/reg_w_1_reg[9]  ( .D(n41535), .CP(clk), .Q(
        \shifter_0/reg_w_1 [9]) );
  dff_sg \shifter_0/reg_w_1_reg[10]  ( .D(n41526), .CP(clk), .Q(
        \shifter_0/reg_w_1 [10]) );
  dff_sg \shifter_0/reg_w_1_reg[11]  ( .D(n41527), .CP(clk), .Q(
        \shifter_0/reg_w_1 [11]) );
  dff_sg \shifter_0/reg_w_1_reg[12]  ( .D(n41941), .CP(clk), .Q(
        \shifter_0/reg_w_1 [12]) );
  dff_sg \shifter_0/reg_w_1_reg[13]  ( .D(n41944), .CP(clk), .Q(
        \shifter_0/reg_w_1 [13]) );
  dff_sg \shifter_0/reg_w_1_reg[14]  ( .D(n41950), .CP(clk), .Q(
        \shifter_0/reg_w_1 [14]) );
  dff_sg \shifter_0/reg_w_1_reg[15]  ( .D(n42037), .CP(clk), .Q(
        \shifter_0/reg_w_1 [15]) );
  dff_sg \shifter_0/reg_w_1_reg[16]  ( .D(n41528), .CP(clk), .Q(
        \shifter_0/reg_w_1 [16]) );
  dff_sg \shifter_0/reg_w_1_reg[17]  ( .D(n42061), .CP(clk), .Q(
        \shifter_0/reg_w_1 [17]) );
  dff_sg \shifter_0/reg_w_1_reg[18]  ( .D(n41935), .CP(clk), .Q(
        \shifter_0/reg_w_1 [18]) );
  dff_sg \shifter_0/reg_w_1_reg[19]  ( .D(n41926), .CP(clk), .Q(
        \shifter_0/reg_w_1 [19]) );
  dff_sg \shifter_0/reg_w_2_reg[0]  ( .D(n42040), .CP(clk), .Q(
        \shifter_0/reg_w_2 [0]) );
  dff_sg \shifter_0/reg_w_2_reg[1]  ( .D(n41947), .CP(clk), .Q(
        \shifter_0/reg_w_2 [1]) );
  dff_sg \shifter_0/reg_w_2_reg[2]  ( .D(n41714), .CP(clk), .Q(
        \shifter_0/reg_w_2 [2]) );
  dff_sg \shifter_0/reg_w_2_reg[3]  ( .D(n41726), .CP(clk), .Q(
        \shifter_0/reg_w_2 [3]) );
  dff_sg \shifter_0/reg_w_2_reg[4]  ( .D(n41704), .CP(clk), .Q(
        \shifter_0/reg_w_2 [4]) );
  dff_sg \shifter_0/reg_w_2_reg[5]  ( .D(n41804), .CP(clk), .Q(
        \shifter_0/reg_w_2 [5]) );
  dff_sg \shifter_0/reg_w_2_reg[6]  ( .D(n41537), .CP(clk), .Q(
        \shifter_0/reg_w_2 [6]) );
  dff_sg \shifter_0/reg_w_2_reg[7]  ( .D(n41871), .CP(clk), .Q(
        \shifter_0/reg_w_2 [7]) );
  dff_sg \shifter_0/reg_w_2_reg[8]  ( .D(n41593), .CP(clk), .Q(
        \shifter_0/reg_w_2 [8]) );
  dff_sg \shifter_0/reg_w_2_reg[9]  ( .D(n41801), .CP(clk), .Q(
        \shifter_0/reg_w_2 [9]) );
  dff_sg \shifter_0/reg_w_2_reg[10]  ( .D(n41549), .CP(clk), .Q(
        \shifter_0/reg_w_2 [10]) );
  dff_sg \shifter_0/reg_w_2_reg[11]  ( .D(n41741), .CP(clk), .Q(
        \shifter_0/reg_w_2 [11]) );
  dff_sg \shifter_0/reg_w_2_reg[12]  ( .D(n41644), .CP(clk), .Q(
        \shifter_0/reg_w_2 [12]) );
  dff_sg \shifter_0/reg_w_2_reg[13]  ( .D(n41611), .CP(clk), .Q(
        \shifter_0/reg_w_2 [13]) );
  dff_sg \shifter_0/reg_w_2_reg[14]  ( .D(n41620), .CP(clk), .Q(
        \shifter_0/reg_w_2 [14]) );
  dff_sg \shifter_0/reg_w_2_reg[15]  ( .D(n41626), .CP(clk), .Q(
        \shifter_0/reg_w_2 [15]) );
  dff_sg \shifter_0/reg_w_2_reg[16]  ( .D(n41608), .CP(clk), .Q(
        \shifter_0/reg_w_2 [16]) );
  dff_sg \shifter_0/reg_w_2_reg[17]  ( .D(n42028), .CP(clk), .Q(
        \shifter_0/reg_w_2 [17]) );
  dff_sg \shifter_0/reg_w_2_reg[18]  ( .D(n41632), .CP(clk), .Q(
        \shifter_0/reg_w_2 [18]) );
  dff_sg \shifter_0/reg_w_2_reg[19]  ( .D(n41638), .CP(clk), .Q(
        \shifter_0/reg_w_2 [19]) );
  dff_sg \shifter_0/reg_w_3_reg[0]  ( .D(n41671), .CP(clk), .Q(
        \shifter_0/reg_w_3 [0]) );
  dff_sg \shifter_0/reg_w_3_reg[1]  ( .D(n41674), .CP(clk), .Q(
        \shifter_0/reg_w_3 [1]) );
  dff_sg \shifter_0/reg_w_3_reg[2]  ( .D(n41677), .CP(clk), .Q(
        \shifter_0/reg_w_3 [2]) );
  dff_sg \shifter_0/reg_w_3_reg[3]  ( .D(n41686), .CP(clk), .Q(
        \shifter_0/reg_w_3 [3]) );
  dff_sg \shifter_0/reg_w_3_reg[4]  ( .D(n41650), .CP(clk), .Q(
        \shifter_0/reg_w_3 [4]) );
  dff_sg \shifter_0/reg_w_3_reg[5]  ( .D(n41656), .CP(clk), .Q(
        \shifter_0/reg_w_3 [5]) );
  dff_sg \shifter_0/reg_w_3_reg[6]  ( .D(n41659), .CP(clk), .Q(
        \shifter_0/reg_w_3 [6]) );
  dff_sg \shifter_0/reg_w_3_reg[7]  ( .D(n41662), .CP(clk), .Q(
        \shifter_0/reg_w_3 [7]) );
  dff_sg \shifter_0/reg_w_3_reg[8]  ( .D(n41680), .CP(clk), .Q(
        \shifter_0/reg_w_3 [8]) );
  dff_sg \shifter_0/reg_w_3_reg[9]  ( .D(n41683), .CP(clk), .Q(
        \shifter_0/reg_w_3 [9]) );
  dff_sg \shifter_0/reg_w_3_reg[10]  ( .D(n41668), .CP(clk), .Q(
        \shifter_0/reg_w_3 [10]) );
  dff_sg \shifter_0/reg_w_3_reg[11]  ( .D(n41777), .CP(clk), .Q(
        \shifter_0/reg_w_3 [11]) );
  dff_sg \shifter_0/reg_w_3_reg[12]  ( .D(n41689), .CP(clk), .Q(
        \shifter_0/reg_w_3 [12]) );
  dff_sg \shifter_0/reg_w_3_reg[13]  ( .D(n41692), .CP(clk), .Q(
        \shifter_0/reg_w_3 [13]) );
  dff_sg \shifter_0/reg_w_3_reg[14]  ( .D(n41541), .CP(clk), .Q(
        \shifter_0/reg_w_3 [14]) );
  dff_sg \shifter_0/reg_w_3_reg[15]  ( .D(n41701), .CP(clk), .Q(
        \shifter_0/reg_w_3 [15]) );
  dff_sg \shifter_0/reg_w_3_reg[16]  ( .D(n41759), .CP(clk), .Q(
        \shifter_0/reg_w_3 [16]) );
  dff_sg \shifter_0/reg_w_3_reg[17]  ( .D(n41572), .CP(clk), .Q(
        \shifter_0/reg_w_3 [17]) );
  dff_sg \shifter_0/reg_w_3_reg[18]  ( .D(n41552), .CP(clk), .Q(
        \shifter_0/reg_w_3 [18]) );
  dff_sg \shifter_0/reg_w_3_reg[19]  ( .D(n42001), .CP(clk), .Q(
        \shifter_0/reg_w_3 [19]) );
  dff_sg \shifter_0/reg_w_4_reg[0]  ( .D(n42103), .CP(clk), .Q(
        \shifter_0/reg_w_4 [0]) );
  dff_sg \shifter_0/reg_w_4_reg[1]  ( .D(n41953), .CP(clk), .Q(
        \shifter_0/reg_w_4 [1]) );
  dff_sg \shifter_0/reg_w_4_reg[2]  ( .D(n41531), .CP(clk), .Q(
        \shifter_0/reg_w_4 [2]) );
  dff_sg \shifter_0/reg_w_4_reg[3]  ( .D(n41530), .CP(clk), .Q(
        \shifter_0/reg_w_4 [3]) );
  dff_sg \shifter_0/reg_w_4_reg[4]  ( .D(n41532), .CP(clk), .Q(
        \shifter_0/reg_w_4 [4]) );
  dff_sg \shifter_0/reg_w_4_reg[5]  ( .D(n41641), .CP(clk), .Q(
        \shifter_0/reg_w_4 [5]) );
  dff_sg \shifter_0/reg_w_4_reg[6]  ( .D(n42070), .CP(clk), .Q(
        \shifter_0/reg_w_4 [6]) );
  dff_sg \shifter_0/reg_w_4_reg[7]  ( .D(n42085), .CP(clk), .Q(
        \shifter_0/reg_w_4 [7]) );
  dff_sg \shifter_0/reg_w_4_reg[8]  ( .D(n41995), .CP(clk), .Q(
        \shifter_0/reg_w_4 [8]) );
  dff_sg \shifter_0/reg_w_4_reg[9]  ( .D(n41698), .CP(clk), .Q(
        \shifter_0/reg_w_4 [9]) );
  dff_sg \shifter_0/reg_w_4_reg[10]  ( .D(n42010), .CP(clk), .Q(
        \shifter_0/reg_w_4 [10]) );
  dff_sg \shifter_0/reg_w_4_reg[11]  ( .D(n41983), .CP(clk), .Q(
        \shifter_0/reg_w_4 [11]) );
  dff_sg \shifter_0/reg_w_4_reg[12]  ( .D(n41614), .CP(clk), .Q(
        \shifter_0/reg_w_4 [12]) );
  dff_sg \shifter_0/reg_w_4_reg[13]  ( .D(n41617), .CP(clk), .Q(
        \shifter_0/reg_w_4 [13]) );
  dff_sg \shifter_0/reg_w_4_reg[14]  ( .D(n41798), .CP(clk), .Q(
        \shifter_0/reg_w_4 [14]) );
  dff_sg \shifter_0/reg_w_4_reg[15]  ( .D(n41647), .CP(clk), .Q(
        \shifter_0/reg_w_4 [15]) );
  dff_sg \shifter_0/reg_w_4_reg[16]  ( .D(n42019), .CP(clk), .Q(
        \shifter_0/reg_w_4 [16]) );
  dff_sg \shifter_0/reg_w_4_reg[17]  ( .D(n42031), .CP(clk), .Q(
        \shifter_0/reg_w_4 [17]) );
  dff_sg \shifter_0/reg_w_4_reg[18]  ( .D(n41923), .CP(clk), .Q(
        \shifter_0/reg_w_4 [18]) );
  dff_sg \shifter_0/reg_w_4_reg[19]  ( .D(n42052), .CP(clk), .Q(
        \shifter_0/reg_w_4 [19]) );
  dff_sg \shifter_0/reg_w_5_reg[0]  ( .D(n41989), .CP(clk), .Q(
        \shifter_0/reg_w_5 [0]) );
  dff_sg \shifter_0/reg_w_5_reg[1]  ( .D(n41992), .CP(clk), .Q(
        \shifter_0/reg_w_5 [1]) );
  dff_sg \shifter_0/reg_w_5_reg[2]  ( .D(n41998), .CP(clk), .Q(
        \shifter_0/reg_w_5 [2]) );
  dff_sg \shifter_0/reg_w_5_reg[3]  ( .D(n42004), .CP(clk), .Q(
        \shifter_0/reg_w_5 [3]) );
  dff_sg \shifter_0/reg_w_5_reg[4]  ( .D(n42013), .CP(clk), .Q(
        \shifter_0/reg_w_5 [4]) );
  dff_sg \shifter_0/reg_w_5_reg[5]  ( .D(n42007), .CP(clk), .Q(
        \shifter_0/reg_w_5 [5]) );
  dff_sg \shifter_0/reg_w_5_reg[6]  ( .D(n41542), .CP(clk), .Q(
        \shifter_0/reg_w_5 [6]) );
  dff_sg \shifter_0/reg_w_5_reg[7]  ( .D(n41540), .CP(clk), .Q(
        \shifter_0/reg_w_5 [7]) );
  dff_sg \shifter_0/reg_w_5_reg[8]  ( .D(n41796), .CP(clk), .Q(
        \shifter_0/reg_w_5 [8]) );
  dff_sg \shifter_0/reg_w_5_reg[9]  ( .D(n41797), .CP(clk), .Q(
        \shifter_0/reg_w_5 [9]) );
  dff_sg \shifter_0/reg_w_5_reg[10]  ( .D(n41793), .CP(clk), .Q(
        \shifter_0/reg_w_5 [10]) );
  dff_sg \shifter_0/reg_w_5_reg[11]  ( .D(n41794), .CP(clk), .Q(
        \shifter_0/reg_w_5 [11]) );
  dff_sg \shifter_0/reg_w_5_reg[12]  ( .D(n41802), .CP(clk), .Q(
        \shifter_0/reg_w_5 [12]) );
  dff_sg \shifter_0/reg_w_5_reg[13]  ( .D(n41803), .CP(clk), .Q(
        \shifter_0/reg_w_5 [13]) );
  dff_sg \shifter_0/reg_w_5_reg[14]  ( .D(n41799), .CP(clk), .Q(
        \shifter_0/reg_w_5 [14]) );
  dff_sg \shifter_0/reg_w_5_reg[15]  ( .D(n41800), .CP(clk), .Q(
        \shifter_0/reg_w_5 [15]) );
  dff_sg \shifter_0/reg_w_5_reg[16]  ( .D(n41784), .CP(clk), .Q(
        \shifter_0/reg_w_5 [16]) );
  dff_sg \shifter_0/reg_w_5_reg[17]  ( .D(n41785), .CP(clk), .Q(
        \shifter_0/reg_w_5 [17]) );
  dff_sg \shifter_0/reg_w_5_reg[18]  ( .D(n41781), .CP(clk), .Q(
        \shifter_0/reg_w_5 [18]) );
  dff_sg \shifter_0/reg_w_5_reg[19]  ( .D(n41782), .CP(clk), .Q(
        \shifter_0/reg_w_5 [19]) );
  dff_sg \shifter_0/reg_w_6_reg[0]  ( .D(n41790), .CP(clk), .Q(
        \shifter_0/reg_w_6 [0]) );
  dff_sg \shifter_0/reg_w_6_reg[1]  ( .D(n41791), .CP(clk), .Q(
        \shifter_0/reg_w_6 [1]) );
  dff_sg \shifter_0/reg_w_6_reg[2]  ( .D(n41787), .CP(clk), .Q(
        \shifter_0/reg_w_6 [2]) );
  dff_sg \shifter_0/reg_w_6_reg[3]  ( .D(n41788), .CP(clk), .Q(
        \shifter_0/reg_w_6 [3]) );
  dff_sg \shifter_0/reg_w_6_reg[4]  ( .D(n41820), .CP(clk), .Q(
        \shifter_0/reg_w_6 [4]) );
  dff_sg \shifter_0/reg_w_6_reg[5]  ( .D(n41821), .CP(clk), .Q(
        \shifter_0/reg_w_6 [5]) );
  dff_sg \shifter_0/reg_w_6_reg[6]  ( .D(n41817), .CP(clk), .Q(
        \shifter_0/reg_w_6 [6]) );
  dff_sg \shifter_0/reg_w_6_reg[7]  ( .D(n41818), .CP(clk), .Q(
        \shifter_0/reg_w_6 [7]) );
  dff_sg \shifter_0/reg_w_6_reg[8]  ( .D(n41826), .CP(clk), .Q(
        \shifter_0/reg_w_6 [8]) );
  dff_sg \shifter_0/reg_w_6_reg[9]  ( .D(n41827), .CP(clk), .Q(
        \shifter_0/reg_w_6 [9]) );
  dff_sg \shifter_0/reg_w_6_reg[10]  ( .D(n41823), .CP(clk), .Q(
        \shifter_0/reg_w_6 [10]) );
  dff_sg \shifter_0/reg_w_6_reg[11]  ( .D(n41824), .CP(clk), .Q(
        \shifter_0/reg_w_6 [11]) );
  dff_sg \shifter_0/reg_w_6_reg[12]  ( .D(n41808), .CP(clk), .Q(
        \shifter_0/reg_w_6 [12]) );
  dff_sg \shifter_0/reg_w_6_reg[13]  ( .D(n41809), .CP(clk), .Q(
        \shifter_0/reg_w_6 [13]) );
  dff_sg \shifter_0/reg_w_6_reg[14]  ( .D(n41805), .CP(clk), .Q(
        \shifter_0/reg_w_6 [14]) );
  dff_sg \shifter_0/reg_w_6_reg[15]  ( .D(n41806), .CP(clk), .Q(
        \shifter_0/reg_w_6 [15]) );
  dff_sg \shifter_0/reg_w_6_reg[16]  ( .D(n41814), .CP(clk), .Q(
        \shifter_0/reg_w_6 [16]) );
  dff_sg \shifter_0/reg_w_6_reg[17]  ( .D(n41815), .CP(clk), .Q(
        \shifter_0/reg_w_6 [17]) );
  dff_sg \shifter_0/reg_w_6_reg[18]  ( .D(n41811), .CP(clk), .Q(
        \shifter_0/reg_w_6 [18]) );
  dff_sg \shifter_0/reg_w_6_reg[19]  ( .D(n41812), .CP(clk), .Q(
        \shifter_0/reg_w_6 [19]) );
  dff_sg \shifter_0/reg_w_7_reg[0]  ( .D(n41748), .CP(clk), .Q(
        \shifter_0/reg_w_7 [0]) );
  dff_sg \shifter_0/reg_w_7_reg[1]  ( .D(n41749), .CP(clk), .Q(
        \shifter_0/reg_w_7 [1]) );
  dff_sg \shifter_0/reg_w_7_reg[2]  ( .D(n41745), .CP(clk), .Q(
        \shifter_0/reg_w_7 [2]) );
  dff_sg \shifter_0/reg_w_7_reg[3]  ( .D(n41746), .CP(clk), .Q(
        \shifter_0/reg_w_7 [3]) );
  dff_sg \shifter_0/reg_w_7_reg[4]  ( .D(n41754), .CP(clk), .Q(
        \shifter_0/reg_w_7 [4]) );
  dff_sg \shifter_0/reg_w_7_reg[5]  ( .D(n41755), .CP(clk), .Q(
        \shifter_0/reg_w_7 [5]) );
  dff_sg \shifter_0/reg_w_7_reg[6]  ( .D(n41751), .CP(clk), .Q(
        \shifter_0/reg_w_7 [6]) );
  dff_sg \shifter_0/reg_w_7_reg[7]  ( .D(n41752), .CP(clk), .Q(
        \shifter_0/reg_w_7 [7]) );
  dff_sg \shifter_0/reg_w_7_reg[8]  ( .D(n41736), .CP(clk), .Q(
        \shifter_0/reg_w_7 [8]) );
  dff_sg \shifter_0/reg_w_7_reg[9]  ( .D(n41737), .CP(clk), .Q(
        \shifter_0/reg_w_7 [9]) );
  dff_sg \shifter_0/reg_w_7_reg[10]  ( .D(n41733), .CP(clk), .Q(
        \shifter_0/reg_w_7 [10]) );
  dff_sg \shifter_0/reg_w_7_reg[11]  ( .D(n41734), .CP(clk), .Q(
        \shifter_0/reg_w_7 [11]) );
  dff_sg \shifter_0/reg_w_7_reg[12]  ( .D(n41742), .CP(clk), .Q(
        \shifter_0/reg_w_7 [12]) );
  dff_sg \shifter_0/reg_w_7_reg[13]  ( .D(n41743), .CP(clk), .Q(
        \shifter_0/reg_w_7 [13]) );
  dff_sg \shifter_0/reg_w_7_reg[14]  ( .D(n41739), .CP(clk), .Q(
        \shifter_0/reg_w_7 [14]) );
  dff_sg \shifter_0/reg_w_7_reg[15]  ( .D(n41740), .CP(clk), .Q(
        \shifter_0/reg_w_7 [15]) );
  dff_sg \shifter_0/reg_w_7_reg[16]  ( .D(n41772), .CP(clk), .Q(
        \shifter_0/reg_w_7 [16]) );
  dff_sg \shifter_0/reg_w_7_reg[17]  ( .D(n41773), .CP(clk), .Q(
        \shifter_0/reg_w_7 [17]) );
  dff_sg \shifter_0/reg_w_7_reg[18]  ( .D(n41769), .CP(clk), .Q(
        \shifter_0/reg_w_7 [18]) );
  dff_sg \shifter_0/reg_w_7_reg[19]  ( .D(n41770), .CP(clk), .Q(
        \shifter_0/reg_w_7 [19]) );
  dff_sg \shifter_0/reg_w_8_reg[0]  ( .D(n41778), .CP(clk), .Q(
        \shifter_0/reg_w_8 [0]) );
  dff_sg \shifter_0/reg_w_8_reg[1]  ( .D(n41779), .CP(clk), .Q(
        \shifter_0/reg_w_8 [1]) );
  dff_sg \shifter_0/reg_w_8_reg[2]  ( .D(n41775), .CP(clk), .Q(
        \shifter_0/reg_w_8 [2]) );
  dff_sg \shifter_0/reg_w_8_reg[3]  ( .D(n41776), .CP(clk), .Q(
        \shifter_0/reg_w_8 [3]) );
  dff_sg \shifter_0/reg_w_8_reg[4]  ( .D(n41760), .CP(clk), .Q(
        \shifter_0/reg_w_8 [4]) );
  dff_sg \shifter_0/reg_w_8_reg[5]  ( .D(n41761), .CP(clk), .Q(
        \shifter_0/reg_w_8 [5]) );
  dff_sg \shifter_0/reg_w_8_reg[6]  ( .D(n41757), .CP(clk), .Q(
        \shifter_0/reg_w_8 [6]) );
  dff_sg \shifter_0/reg_w_8_reg[7]  ( .D(n41758), .CP(clk), .Q(
        \shifter_0/reg_w_8 [7]) );
  dff_sg \shifter_0/reg_w_8_reg[8]  ( .D(n41766), .CP(clk), .Q(
        \shifter_0/reg_w_8 [8]) );
  dff_sg \shifter_0/reg_w_8_reg[9]  ( .D(n41767), .CP(clk), .Q(
        \shifter_0/reg_w_8 [9]) );
  dff_sg \shifter_0/reg_w_8_reg[10]  ( .D(n41763), .CP(clk), .Q(
        \shifter_0/reg_w_8 [10]) );
  dff_sg \shifter_0/reg_w_8_reg[11]  ( .D(n41764), .CP(clk), .Q(
        \shifter_0/reg_w_8 [11]) );
  dff_sg \shifter_0/reg_w_8_reg[12]  ( .D(n41887), .CP(clk), .Q(
        \shifter_0/reg_w_8 [12]) );
  dff_sg \shifter_0/reg_w_8_reg[13]  ( .D(n41888), .CP(clk), .Q(
        \shifter_0/reg_w_8 [13]) );
  dff_sg \shifter_0/reg_w_8_reg[14]  ( .D(n41884), .CP(clk), .Q(
        \shifter_0/reg_w_8 [14]) );
  dff_sg \shifter_0/reg_w_8_reg[15]  ( .D(n41885), .CP(clk), .Q(
        \shifter_0/reg_w_8 [15]) );
  dff_sg \shifter_0/reg_w_8_reg[16]  ( .D(n41893), .CP(clk), .Q(
        \shifter_0/reg_w_8 [16]) );
  dff_sg \shifter_0/reg_w_8_reg[17]  ( .D(n41894), .CP(clk), .Q(
        \shifter_0/reg_w_8 [17]) );
  dff_sg \shifter_0/reg_w_8_reg[18]  ( .D(n41890), .CP(clk), .Q(
        \shifter_0/reg_w_8 [18]) );
  dff_sg \shifter_0/reg_w_8_reg[19]  ( .D(n41891), .CP(clk), .Q(
        \shifter_0/reg_w_8 [19]) );
  dff_sg \shifter_0/reg_w_9_reg[0]  ( .D(n41875), .CP(clk), .Q(
        \shifter_0/reg_w_9 [0]) );
  dff_sg \shifter_0/reg_w_9_reg[1]  ( .D(n41876), .CP(clk), .Q(
        \shifter_0/reg_w_9 [1]) );
  dff_sg \shifter_0/reg_w_9_reg[2]  ( .D(n41872), .CP(clk), .Q(
        \shifter_0/reg_w_9 [2]) );
  dff_sg \shifter_0/reg_w_9_reg[3]  ( .D(n41873), .CP(clk), .Q(
        \shifter_0/reg_w_9 [3]) );
  dff_sg \shifter_0/reg_w_9_reg[4]  ( .D(n41881), .CP(clk), .Q(
        \shifter_0/reg_w_9 [4]) );
  dff_sg \shifter_0/reg_w_9_reg[5]  ( .D(n41882), .CP(clk), .Q(
        \shifter_0/reg_w_9 [5]) );
  dff_sg \shifter_0/reg_w_9_reg[6]  ( .D(n41878), .CP(clk), .Q(
        \shifter_0/reg_w_9 [6]) );
  dff_sg \shifter_0/reg_w_9_reg[7]  ( .D(n41879), .CP(clk), .Q(
        \shifter_0/reg_w_9 [7]) );
  dff_sg \shifter_0/reg_w_9_reg[8]  ( .D(n41911), .CP(clk), .Q(
        \shifter_0/reg_w_9 [8]) );
  dff_sg \shifter_0/reg_w_9_reg[9]  ( .D(n41912), .CP(clk), .Q(
        \shifter_0/reg_w_9 [9]) );
  dff_sg \shifter_0/reg_w_9_reg[10]  ( .D(n41908), .CP(clk), .Q(
        \shifter_0/reg_w_9 [10]) );
  dff_sg \shifter_0/reg_w_9_reg[11]  ( .D(n41909), .CP(clk), .Q(
        \shifter_0/reg_w_9 [11]) );
  dff_sg \shifter_0/reg_w_9_reg[12]  ( .D(n41910), .CP(clk), .Q(
        \shifter_0/reg_w_9 [12]) );
  dff_sg \shifter_0/reg_w_9_reg[13]  ( .D(n41886), .CP(clk), .Q(
        \shifter_0/reg_w_9 [13]) );
  dff_sg \shifter_0/reg_w_9_reg[14]  ( .D(n41914), .CP(clk), .Q(
        \shifter_0/reg_w_9 [14]) );
  dff_sg \shifter_0/reg_w_9_reg[15]  ( .D(n41915), .CP(clk), .Q(
        \shifter_0/reg_w_9 [15]) );
  dff_sg \shifter_0/reg_w_9_reg[16]  ( .D(n41899), .CP(clk), .Q(
        \shifter_0/reg_w_9 [16]) );
  dff_sg \shifter_0/reg_w_9_reg[17]  ( .D(n41900), .CP(clk), .Q(
        \shifter_0/reg_w_9 [17]) );
  dff_sg \shifter_0/reg_w_9_reg[18]  ( .D(n41896), .CP(clk), .Q(
        \shifter_0/reg_w_9 [18]) );
  dff_sg \shifter_0/reg_w_9_reg[19]  ( .D(n41897), .CP(clk), .Q(
        \shifter_0/reg_w_9 [19]) );
  dff_sg \shifter_0/reg_w_10_reg[0]  ( .D(n41905), .CP(clk), .Q(
        \shifter_0/reg_w_10 [0]) );
  dff_sg \shifter_0/reg_w_10_reg[1]  ( .D(n41906), .CP(clk), .Q(
        \shifter_0/reg_w_10 [1]) );
  dff_sg \shifter_0/reg_w_10_reg[2]  ( .D(n41902), .CP(clk), .Q(
        \shifter_0/reg_w_10 [2]) );
  dff_sg \shifter_0/reg_w_10_reg[3]  ( .D(n41903), .CP(clk), .Q(
        \shifter_0/reg_w_10 [3]) );
  dff_sg \shifter_0/reg_w_10_reg[4]  ( .D(n41845), .CP(clk), .Q(
        \shifter_0/reg_w_10 [4]) );
  dff_sg \shifter_0/reg_w_10_reg[5]  ( .D(n41846), .CP(clk), .Q(
        \shifter_0/reg_w_10 [5]) );
  dff_sg \shifter_0/reg_w_10_reg[6]  ( .D(n41842), .CP(clk), .Q(
        \shifter_0/reg_w_10 [6]) );
  dff_sg \shifter_0/reg_w_10_reg[7]  ( .D(n41843), .CP(clk), .Q(
        \shifter_0/reg_w_10 [7]) );
  dff_sg \shifter_0/reg_w_10_reg[8]  ( .D(n41850), .CP(clk), .Q(
        \shifter_0/reg_w_10 [8]) );
  dff_sg \shifter_0/reg_w_10_reg[9]  ( .D(n41856), .CP(clk), .Q(
        \shifter_0/reg_w_10 [9]) );
  dff_sg \shifter_0/reg_w_10_reg[10]  ( .D(n41707), .CP(clk), .Q(
        \shifter_0/reg_w_10 [10]) );
  dff_sg \shifter_0/reg_w_10_reg[11]  ( .D(n41831), .CP(clk), .Q(
        \shifter_0/reg_w_10 [11]) );
  dff_sg \shifter_0/reg_w_10_reg[12]  ( .D(n41832), .CP(clk), .Q(
        \shifter_0/reg_w_10 [12]) );
  dff_sg \shifter_0/reg_w_10_reg[13]  ( .D(n41833), .CP(clk), .Q(
        \shifter_0/reg_w_10 [13]) );
  dff_sg \shifter_0/reg_w_10_reg[14]  ( .D(n41829), .CP(clk), .Q(
        \shifter_0/reg_w_10 [14]) );
  dff_sg \shifter_0/reg_w_10_reg[15]  ( .D(n41830), .CP(clk), .Q(
        \shifter_0/reg_w_10 [15]) );
  dff_sg \shifter_0/reg_w_10_reg[16]  ( .D(n41838), .CP(clk), .Q(
        \shifter_0/reg_w_10 [16]) );
  dff_sg \shifter_0/reg_w_10_reg[17]  ( .D(n41839), .CP(clk), .Q(
        \shifter_0/reg_w_10 [17]) );
  dff_sg \shifter_0/reg_w_10_reg[18]  ( .D(n41835), .CP(clk), .Q(
        \shifter_0/reg_w_10 [18]) );
  dff_sg \shifter_0/reg_w_10_reg[19]  ( .D(n41836), .CP(clk), .Q(
        \shifter_0/reg_w_10 [19]) );
  dff_sg \shifter_0/reg_w_11_reg[0]  ( .D(n41863), .CP(clk), .Q(
        \shifter_0/reg_w_11 [0]) );
  dff_sg \shifter_0/reg_w_11_reg[1]  ( .D(n41864), .CP(clk), .Q(
        \shifter_0/reg_w_11 [1]) );
  dff_sg \shifter_0/reg_w_11_reg[2]  ( .D(n41860), .CP(clk), .Q(
        \shifter_0/reg_w_11 [2]) );
  dff_sg \shifter_0/reg_w_11_reg[3]  ( .D(n41861), .CP(clk), .Q(
        \shifter_0/reg_w_11 [3]) );
  dff_sg \shifter_0/reg_w_11_reg[4]  ( .D(n41869), .CP(clk), .Q(
        \shifter_0/reg_w_11 [4]) );
  dff_sg \shifter_0/reg_w_11_reg[5]  ( .D(n41870), .CP(clk), .Q(
        \shifter_0/reg_w_11 [5]) );
  dff_sg \shifter_0/reg_w_11_reg[6]  ( .D(n41866), .CP(clk), .Q(
        \shifter_0/reg_w_11 [6]) );
  dff_sg \shifter_0/reg_w_11_reg[7]  ( .D(n41867), .CP(clk), .Q(
        \shifter_0/reg_w_11 [7]) );
  dff_sg \shifter_0/reg_w_11_reg[8]  ( .D(n41851), .CP(clk), .Q(
        \shifter_0/reg_w_11 [8]) );
  dff_sg \shifter_0/reg_w_11_reg[9]  ( .D(n41852), .CP(clk), .Q(
        \shifter_0/reg_w_11 [9]) );
  dff_sg \shifter_0/reg_w_11_reg[10]  ( .D(n41848), .CP(clk), .Q(
        \shifter_0/reg_w_11 [10]) );
  dff_sg \shifter_0/reg_w_11_reg[11]  ( .D(n41849), .CP(clk), .Q(
        \shifter_0/reg_w_11 [11]) );
  dff_sg \shifter_0/reg_w_11_reg[12]  ( .D(n41857), .CP(clk), .Q(
        \shifter_0/reg_w_11 [12]) );
  dff_sg \shifter_0/reg_w_11_reg[13]  ( .D(n41858), .CP(clk), .Q(
        \shifter_0/reg_w_11 [13]) );
  dff_sg \shifter_0/reg_w_11_reg[14]  ( .D(n41854), .CP(clk), .Q(
        \shifter_0/reg_w_11 [14]) );
  dff_sg \shifter_0/reg_w_11_reg[15]  ( .D(n41855), .CP(clk), .Q(
        \shifter_0/reg_w_11 [15]) );
  dff_sg \shifter_0/reg_w_11_reg[16]  ( .D(n41672), .CP(clk), .Q(
        \shifter_0/reg_w_11 [16]) );
  dff_sg \shifter_0/reg_w_11_reg[17]  ( .D(n41673), .CP(clk), .Q(
        \shifter_0/reg_w_11 [17]) );
  dff_sg \shifter_0/reg_w_11_reg[18]  ( .D(n41669), .CP(clk), .Q(
        \shifter_0/reg_w_11 [18]) );
  dff_sg \shifter_0/reg_w_11_reg[19]  ( .D(n41670), .CP(clk), .Q(
        \shifter_0/reg_w_11 [19]) );
  dff_sg \shifter_0/reg_w_12_reg[0]  ( .D(n41678), .CP(clk), .Q(
        \shifter_0/reg_w_12 [0]) );
  dff_sg \shifter_0/reg_w_12_reg[1]  ( .D(n41679), .CP(clk), .Q(
        \shifter_0/reg_w_12 [1]) );
  dff_sg \shifter_0/reg_w_12_reg[2]  ( .D(n41675), .CP(clk), .Q(
        \shifter_0/reg_w_12 [2]) );
  dff_sg \shifter_0/reg_w_12_reg[3]  ( .D(n41676), .CP(clk), .Q(
        \shifter_0/reg_w_12 [3]) );
  dff_sg \shifter_0/reg_w_12_reg[4]  ( .D(n41660), .CP(clk), .Q(
        \shifter_0/reg_w_12 [4]) );
  dff_sg \shifter_0/reg_w_12_reg[5]  ( .D(n41661), .CP(clk), .Q(
        \shifter_0/reg_w_12 [5]) );
  dff_sg \shifter_0/reg_w_12_reg[6]  ( .D(n41657), .CP(clk), .Q(
        \shifter_0/reg_w_12 [6]) );
  dff_sg \shifter_0/reg_w_12_reg[7]  ( .D(n41658), .CP(clk), .Q(
        \shifter_0/reg_w_12 [7]) );
  dff_sg \shifter_0/reg_w_12_reg[8]  ( .D(n41666), .CP(clk), .Q(
        \shifter_0/reg_w_12 [8]) );
  dff_sg \shifter_0/reg_w_12_reg[9]  ( .D(n41667), .CP(clk), .Q(
        \shifter_0/reg_w_12 [9]) );
  dff_sg \shifter_0/reg_w_12_reg[10]  ( .D(n41663), .CP(clk), .Q(
        \shifter_0/reg_w_12 [10]) );
  dff_sg \shifter_0/reg_w_12_reg[11]  ( .D(n41664), .CP(clk), .Q(
        \shifter_0/reg_w_12 [11]) );
  dff_sg \shifter_0/reg_w_12_reg[12]  ( .D(n41696), .CP(clk), .Q(
        \shifter_0/reg_w_12 [12]) );
  dff_sg \shifter_0/reg_w_12_reg[13]  ( .D(n41697), .CP(clk), .Q(
        \shifter_0/reg_w_12 [13]) );
  dff_sg \shifter_0/reg_w_12_reg[14]  ( .D(n41693), .CP(clk), .Q(
        \shifter_0/reg_w_12 [14]) );
  dff_sg \shifter_0/reg_w_12_reg[15]  ( .D(n41694), .CP(clk), .Q(
        \shifter_0/reg_w_12 [15]) );
  dff_sg \shifter_0/reg_w_12_reg[16]  ( .D(n41702), .CP(clk), .Q(
        \shifter_0/reg_w_12 [16]) );
  dff_sg \shifter_0/reg_w_12_reg[17]  ( .D(n41703), .CP(clk), .Q(
        \shifter_0/reg_w_12 [17]) );
  dff_sg \shifter_0/reg_w_12_reg[18]  ( .D(n41699), .CP(clk), .Q(
        \shifter_0/reg_w_12 [18]) );
  dff_sg \shifter_0/reg_w_12_reg[19]  ( .D(n41700), .CP(clk), .Q(
        \shifter_0/reg_w_12 [19]) );
  dff_sg \shifter_0/reg_w_13_reg[0]  ( .D(n41684), .CP(clk), .Q(
        \shifter_0/reg_w_13 [0]) );
  dff_sg \shifter_0/reg_w_13_reg[1]  ( .D(n41685), .CP(clk), .Q(
        \shifter_0/reg_w_13 [1]) );
  dff_sg \shifter_0/reg_w_13_reg[2]  ( .D(n41681), .CP(clk), .Q(
        \shifter_0/reg_w_13 [2]) );
  dff_sg \shifter_0/reg_w_13_reg[3]  ( .D(n41682), .CP(clk), .Q(
        \shifter_0/reg_w_13 [3]) );
  dff_sg \shifter_0/reg_w_13_reg[4]  ( .D(n41690), .CP(clk), .Q(
        \shifter_0/reg_w_13 [4]) );
  dff_sg \shifter_0/reg_w_13_reg[5]  ( .D(n41691), .CP(clk), .Q(
        \shifter_0/reg_w_13 [5]) );
  dff_sg \shifter_0/reg_w_13_reg[6]  ( .D(n41687), .CP(clk), .Q(
        \shifter_0/reg_w_13 [6]) );
  dff_sg \shifter_0/reg_w_13_reg[7]  ( .D(n41688), .CP(clk), .Q(
        \shifter_0/reg_w_13 [7]) );
  dff_sg \shifter_0/reg_w_13_reg[8]  ( .D(n41624), .CP(clk), .Q(
        \shifter_0/reg_w_13 [8]) );
  dff_sg \shifter_0/reg_w_13_reg[9]  ( .D(n41625), .CP(clk), .Q(
        \shifter_0/reg_w_13 [9]) );
  dff_sg \shifter_0/reg_w_13_reg[10]  ( .D(n41621), .CP(clk), .Q(
        \shifter_0/reg_w_13 [10]) );
  dff_sg \shifter_0/reg_w_13_reg[11]  ( .D(n41622), .CP(clk), .Q(
        \shifter_0/reg_w_13 [11]) );
  dff_sg \shifter_0/reg_w_13_reg[12]  ( .D(n41630), .CP(clk), .Q(
        \shifter_0/reg_w_13 [12]) );
  dff_sg \shifter_0/reg_w_13_reg[13]  ( .D(n41631), .CP(clk), .Q(
        \shifter_0/reg_w_13 [13]) );
  dff_sg \shifter_0/reg_w_13_reg[14]  ( .D(n41627), .CP(clk), .Q(
        \shifter_0/reg_w_13 [14]) );
  dff_sg \shifter_0/reg_w_13_reg[15]  ( .D(n41628), .CP(clk), .Q(
        \shifter_0/reg_w_13 [15]) );
  dff_sg \shifter_0/reg_w_13_reg[16]  ( .D(n41612), .CP(clk), .Q(
        \shifter_0/reg_w_13 [16]) );
  dff_sg \shifter_0/reg_w_13_reg[17]  ( .D(n41613), .CP(clk), .Q(
        \shifter_0/reg_w_13 [17]) );
  dff_sg \shifter_0/reg_w_13_reg[18]  ( .D(n41609), .CP(clk), .Q(
        \shifter_0/reg_w_13 [18]) );
  dff_sg \shifter_0/reg_w_13_reg[19]  ( .D(n41610), .CP(clk), .Q(
        \shifter_0/reg_w_13 [19]) );
  dff_sg \shifter_0/reg_w_14_reg[0]  ( .D(n41618), .CP(clk), .Q(
        \shifter_0/reg_w_14 [0]) );
  dff_sg \shifter_0/reg_w_14_reg[1]  ( .D(n41619), .CP(clk), .Q(
        \shifter_0/reg_w_14 [1]) );
  dff_sg \shifter_0/reg_w_14_reg[2]  ( .D(n41615), .CP(clk), .Q(
        \shifter_0/reg_w_14 [2]) );
  dff_sg \shifter_0/reg_w_14_reg[3]  ( .D(n41616), .CP(clk), .Q(
        \shifter_0/reg_w_14 [3]) );
  dff_sg \shifter_0/reg_w_14_reg[4]  ( .D(n41648), .CP(clk), .Q(
        \shifter_0/reg_w_14 [4]) );
  dff_sg \shifter_0/reg_w_14_reg[5]  ( .D(n41649), .CP(clk), .Q(
        \shifter_0/reg_w_14 [5]) );
  dff_sg \shifter_0/reg_w_14_reg[6]  ( .D(n41645), .CP(clk), .Q(
        \shifter_0/reg_w_14 [6]) );
  dff_sg \shifter_0/reg_w_14_reg[7]  ( .D(n41646), .CP(clk), .Q(
        \shifter_0/reg_w_14 [7]) );
  dff_sg \shifter_0/reg_w_14_reg[8]  ( .D(n41654), .CP(clk), .Q(
        \shifter_0/reg_w_14 [8]) );
  dff_sg \shifter_0/reg_w_14_reg[9]  ( .D(n41655), .CP(clk), .Q(
        \shifter_0/reg_w_14 [9]) );
  dff_sg \shifter_0/reg_w_14_reg[10]  ( .D(n41651), .CP(clk), .Q(
        \shifter_0/reg_w_14 [10]) );
  dff_sg \shifter_0/reg_w_14_reg[11]  ( .D(n41652), .CP(clk), .Q(
        \shifter_0/reg_w_14 [11]) );
  dff_sg \shifter_0/reg_w_14_reg[12]  ( .D(n41636), .CP(clk), .Q(
        \shifter_0/reg_w_14 [12]) );
  dff_sg \shifter_0/reg_w_14_reg[13]  ( .D(n41637), .CP(clk), .Q(
        \shifter_0/reg_w_14 [13]) );
  dff_sg \shifter_0/reg_w_14_reg[14]  ( .D(n41633), .CP(clk), .Q(
        \shifter_0/reg_w_14 [14]) );
  dff_sg \shifter_0/reg_w_14_reg[15]  ( .D(n41634), .CP(clk), .Q(
        \shifter_0/reg_w_14 [15]) );
  dff_sg \shifter_0/reg_w_14_reg[16]  ( .D(n41642), .CP(clk), .Q(
        \shifter_0/reg_w_14 [16]) );
  dff_sg \shifter_0/reg_w_14_reg[17]  ( .D(n41643), .CP(clk), .Q(
        \shifter_0/reg_w_14 [17]) );
  dff_sg \shifter_0/reg_w_14_reg[18]  ( .D(n41639), .CP(clk), .Q(
        \shifter_0/reg_w_14 [18]) );
  dff_sg \shifter_0/reg_w_14_reg[19]  ( .D(n41640), .CP(clk), .Q(
        \shifter_0/reg_w_14 [19]) );
  dff_sg \shifter_0/w_pointer_reg[0]  ( .D(n42804), .CP(clk), .Q(
        \shifter_0/w_pointer [0]) );
  dff_sg \shifter_0/w_pointer_reg[1]  ( .D(n42805), .CP(clk), .Q(
        \shifter_0/w_pointer [1]) );
  dff_sg \shifter_0/w_pointer_reg[2]  ( .D(n42806), .CP(clk), .Q(
        \shifter_0/w_pointer [2]) );
  dff_sg \shifter_0/w_pointer_reg[3]  ( .D(n42807), .CP(clk), .Q(
        \shifter_0/w_pointer [3]) );
  dff_sg \shifter_0/reg_w_15_reg[0]  ( .D(n41724), .CP(clk), .Q(
        \shifter_0/reg_w_15 [0]) );
  dff_sg \shifter_0/reg_w_15_reg[1]  ( .D(n41725), .CP(clk), .Q(
        \shifter_0/reg_w_15 [1]) );
  dff_sg \shifter_0/reg_w_15_reg[2]  ( .D(n41721), .CP(clk), .Q(
        \shifter_0/reg_w_15 [2]) );
  dff_sg \shifter_0/reg_w_15_reg[3]  ( .D(n41722), .CP(clk), .Q(
        \shifter_0/reg_w_15 [3]) );
  dff_sg \shifter_0/reg_w_15_reg[4]  ( .D(n41730), .CP(clk), .Q(
        \shifter_0/reg_w_15 [4]) );
  dff_sg \shifter_0/reg_w_15_reg[5]  ( .D(n41731), .CP(clk), .Q(
        \shifter_0/reg_w_15 [5]) );
  dff_sg \shifter_0/reg_w_15_reg[6]  ( .D(n41727), .CP(clk), .Q(
        \shifter_0/reg_w_15 [6]) );
  dff_sg \shifter_0/reg_w_15_reg[7]  ( .D(n41728), .CP(clk), .Q(
        \shifter_0/reg_w_15 [7]) );
  dff_sg \shifter_0/reg_w_15_reg[8]  ( .D(n41712), .CP(clk), .Q(
        \shifter_0/reg_w_15 [8]) );
  dff_sg \shifter_0/reg_w_15_reg[9]  ( .D(n41713), .CP(clk), .Q(
        \shifter_0/reg_w_15 [9]) );
  dff_sg \shifter_0/reg_w_15_reg[10]  ( .D(n41709), .CP(clk), .Q(
        \shifter_0/reg_w_15 [10]) );
  dff_sg \shifter_0/reg_w_15_reg[11]  ( .D(n41710), .CP(clk), .Q(
        \shifter_0/reg_w_15 [11]) );
  dff_sg \shifter_0/reg_w_15_reg[12]  ( .D(n41718), .CP(clk), .Q(
        \shifter_0/reg_w_15 [12]) );
  dff_sg \shifter_0/reg_w_15_reg[13]  ( .D(n41719), .CP(clk), .Q(
        \shifter_0/reg_w_15 [13]) );
  dff_sg \shifter_0/reg_w_15_reg[14]  ( .D(n41715), .CP(clk), .Q(
        \shifter_0/reg_w_15 [14]) );
  dff_sg \shifter_0/reg_w_15_reg[15]  ( .D(n41716), .CP(clk), .Q(
        \shifter_0/reg_w_15 [15]) );
  dff_sg \shifter_0/reg_w_15_reg[16]  ( .D(n42146), .CP(clk), .Q(
        \shifter_0/reg_w_15 [16]) );
  dff_sg \shifter_0/reg_w_15_reg[17]  ( .D(n42125), .CP(clk), .Q(
        \shifter_0/reg_w_15 [17]) );
  dff_sg \shifter_0/reg_w_15_reg[18]  ( .D(n42152), .CP(clk), .Q(
        \shifter_0/reg_w_15 [18]) );
  dff_sg \shifter_0/reg_w_15_reg[19]  ( .D(n42158), .CP(clk), .Q(
        \shifter_0/reg_w_15 [19]) );
  dff_sg \shifter_0/pointer_reg[3]  ( .D(n42808), .CP(clk), .Q(
        \shifter_0/pointer [3]) );
  dff_sg \shifter_0/pointer_reg[1]  ( .D(n42810), .CP(clk), .Q(
        \shifter_0/pointer [1]) );
  dff_sg \shifter_0/state_reg[0]  ( .D(n42801), .CP(clk), .Q(
        \shifter_0/n27115 ) );
  dff_sg \shifter_0/state_reg[1]  ( .D(n42802), .CP(clk), .Q(
        \shifter_0/n27114 ) );
  dff_sg \shifter_0/pointer_reg[2]  ( .D(n42809), .CP(clk), .Q(
        \shifter_0/pointer [2]) );
  dff_sg \shifter_0/pointer_reg[0]  ( .D(n42803), .CP(clk), .Q(
        \shifter_0/pointer [0]) );
  nor_x2_sg U27436 ( .A(n68590), .B(n31941), .X(n31940) );
  nor_x2_sg U27440 ( .A(n68591), .B(n31945), .X(n31939) );
  nor_x2_sg U27446 ( .A(n31952), .B(n31953), .X(n31951) );
  nor_x2_sg U27450 ( .A(n57300), .B(n31957), .X(n31949) );
  nor_x2_sg U27451 ( .A(n31958), .B(n31959), .X(n31957) );
  nor_x2_sg U27463 ( .A(n47329), .B(n31967), .X(n31971) );
  nor_x2_sg U27472 ( .A(n47393), .B(n31967), .X(n31982) );
  nor_x2_sg U27527 ( .A(n47310), .B(n31967), .X(n31996) );
  nand_x8_sg U27528 ( .A(n47491), .B(n61910), .X(n31967) );
  nor_x2_sg U27563 ( .A(n32078), .B(n57859), .X(n32077) );
  nor_x2_sg U27564 ( .A(n32079), .B(n68587), .X(n32076) );
  nor_x2_sg U27572 ( .A(n68589), .B(n32089), .X(n32083) );
  nor_x2_sg U27872 ( .A(n47289), .B(n32374), .X(n32369) );
  nor_x2_sg U27881 ( .A(n47293), .B(n32374), .X(n32381) );
  nor_x2_sg U27903 ( .A(n68590), .B(n32409), .X(n32408) );
  nor_x2_sg U27907 ( .A(n68591), .B(n32413), .X(n32407) );
  nor_x2_sg U27913 ( .A(n32420), .B(n32421), .X(n32419) );
  nor_x2_sg U27917 ( .A(n57306), .B(n32424), .X(n32417) );
  nor_x2_sg U27918 ( .A(n32425), .B(n32426), .X(n32424) );
  nand_x8_sg U27933 ( .A(n31994), .B(n32437), .X(n32372) );
  nor_x2_sg U27977 ( .A(n47391), .B(n32374), .X(n32438) );
  nand_x8_sg U27978 ( .A(n68265), .B(n61910), .X(n32374) );
  nor_x2_sg U28021 ( .A(n32523), .B(n57859), .X(n32522) );
  nor_x2_sg U28022 ( .A(n32524), .B(n68587), .X(n32521) );
  nor_x2_sg U28030 ( .A(n68589), .B(n32534), .X(n32528) );
  nand_x8_sg U28545 ( .A(n68230), .B(n32965), .X(n32926) );
  nand_x8_sg U28607 ( .A(n68230), .B(n33008), .X(n32969) );
  nand_x8_sg U28669 ( .A(n68231), .B(n33051), .X(n33012) );
  nand_x8_sg U28731 ( .A(n68231), .B(n33094), .X(n33055) );
  nand_x8_sg U28793 ( .A(n68229), .B(n32965), .X(n33098) );
  nand_x8_sg U28855 ( .A(n68229), .B(n33179), .X(n33140) );
  nand_x8_sg U28917 ( .A(n33222), .B(n33179), .X(n33183) );
  nand_x8_sg U28979 ( .A(n33265), .B(n33179), .X(n33226) );
  nand_x8_sg U28980 ( .A(n57166), .B(n68376), .X(n33179) );
  nand_x8_sg U29042 ( .A(n33309), .B(n33310), .X(n33270) );
  nand_x8_sg U29104 ( .A(n68228), .B(n33310), .X(n33314) );
  nand_x8_sg U29166 ( .A(n68231), .B(n33310), .X(n33356) );
  nand_x8_sg U29230 ( .A(n33309), .B(n33051), .X(n33401) );
  nand_x8_sg U29292 ( .A(n68228), .B(n33051), .X(n33443) );
  nand_x8_sg U29354 ( .A(n68228), .B(n33524), .X(n33485) );
  nand_x8_sg U29416 ( .A(n33309), .B(n33524), .X(n33528) );
  nand_x8_sg U29478 ( .A(n68229), .B(n33609), .X(n33570) );
  nand_x8_sg U29540 ( .A(n68230), .B(n33609), .X(n33613) );
  nand_x8_sg U29604 ( .A(n33265), .B(n33609), .X(n33657) );
  nand_x8_sg U29666 ( .A(n33222), .B(n33609), .X(n33699) );
  nand_x8_sg U29667 ( .A(n57166), .B(n68378), .X(n33609) );
  nand_x8_sg U29793 ( .A(n33222), .B(n33008), .X(n33787) );
  nand_x8_sg U29855 ( .A(n33265), .B(n33008), .X(n33829) );
  nand_x8_sg U29856 ( .A(n57166), .B(n68375), .X(n33008) );
  nand_x8_sg U29982 ( .A(n33955), .B(n33094), .X(n33916) );
  nand_x8_sg U30044 ( .A(n33955), .B(n33051), .X(n33959) );
  nand_x8_sg U30045 ( .A(n57166), .B(n68383), .X(n33051) );
  nand_x8_sg U30172 ( .A(n57166), .B(n68382), .X(n33094) );
  nand_x8_sg U30236 ( .A(n33955), .B(n33524), .X(n34092) );
  nand_x8_sg U30237 ( .A(n57166), .B(n68381), .X(n33524) );
  nand_x8_sg U30300 ( .A(n57166), .B(n68377), .X(n32965) );
  nand_x8_sg U30367 ( .A(n57166), .B(n68384), .X(n33310) );
  nand_x8_sg U30372 ( .A(n57166), .B(n57855), .X(n33396) );
  nand_x8_sg U32792 ( .A(n35840), .B(n61908), .X(n35705) );
  \**FFGEN**  \filter_0/next_w_pointer_reg[0]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(n67586), .force_10(
        \filter_0/n8240 ), .force_11(1'b0), .Q(n40871) );
  \**FFGEN**  \filter_0/next_w_pointer_reg[1]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n8243 ), 
        .force_10(n67585), .force_11(1'b0), .Q(n40870) );
  \**FFGEN**  \filter_0/next_w_pointer_reg[2]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n8247 ), 
        .force_10(n67584), .force_11(1'b0), .Q(n40869) );
  \**FFGEN**  \filter_0/next_w_pointer_reg[3]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(n67583), .force_10(
        \filter_0/n8252 ), .force_11(1'b0), .Q(n40868) );
  \**FFGEN**  \filter_0/next_i_pointer_reg[1]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n8255 ), 
        .force_10(n67579), .force_11(1'b0), .Q(n40874) );
  \**FFGEN**  \filter_0/next_i_pointer_reg[2]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n8259 ), 
        .force_10(n67578), .force_11(1'b0), .Q(n40873) );
  \**FFGEN**  \filter_0/next_i_pointer_reg[3]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(n67577), .force_10(
        \filter_0/n8264 ), .force_11(1'b0), .Q(n40872) );
  \**FFGEN**  \filter_0/next_i_pointer_reg[0]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(n67580), .force_10(
        \filter_0/n8268 ), .force_11(1'b0), .Q(n40875) );
  \**FFGEN**  \filter_0/next_m_pointer_reg[0]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n8271 ), 
        .force_10(\filter_0/n8272 ), .force_11(1'b0), .Q(n40880) );
  \**FFGEN**  \filter_0/next_m_pointer_reg[1]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(n67531), .force_10(
        \filter_0/n8276 ), .force_11(1'b0), .Q(n40879) );
  \**FFGEN**  \filter_0/next_m_pointer_reg[2]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n8279 ), 
        .force_10(n67533), .force_11(1'b0), .Q(n40878) );
  \**FFGEN**  \filter_0/next_m_pointer_reg[3]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(n67538), .force_10(
        \filter_0/n8284 ), .force_11(1'b0), .Q(n40877) );
  \**FFGEN**  \filter_0/next_m_pointer_reg[4]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n8287 ), 
        .force_10(n67539), .force_11(1'b0), .Q(n40876) );
  \**FFGEN**  \filter_0/pre_ow_15_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8291 ), .force_10(
        \filter_0/n8292 ), .force_11(1'b0), .Q(n40774) );
  \**FFGEN**  \filter_0/pre_ow_15_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8295 ), .force_10(
        \filter_0/n8296 ), .force_11(1'b0), .Q(n40773) );
  \**FFGEN**  \filter_0/pre_ow_15_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8299 ), .force_10(
        \filter_0/n8300 ), .force_11(1'b0), .Q(n40772) );
  \**FFGEN**  \filter_0/pre_ow_15_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8303 ), .force_10(
        \filter_0/n8304 ), .force_11(1'b0), .Q(n40771) );
  \**FFGEN**  \filter_0/pre_ow_15_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8307 ), .force_10(
        \filter_0/n8308 ), .force_11(1'b0), .Q(n40483) );
  \**FFGEN**  \filter_0/pre_ow_15_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8311 ), .force_10(
        \filter_0/n8312 ), .force_11(1'b0), .Q(n40451) );
  \**FFGEN**  \filter_0/pre_ow_15_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8315 ), .force_10(
        \filter_0/n8316 ), .force_11(1'b0), .Q(n40355) );
  \**FFGEN**  \filter_0/pre_ow_15_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8319 ), .force_10(
        \filter_0/n8320 ), .force_11(1'b0), .Q(n40420) );
  \**FFGEN**  \filter_0/pre_ow_15_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8323 ), .force_10(
        \filter_0/n8324 ), .force_11(1'b0), .Q(n40321) );
  \**FFGEN**  \filter_0/pre_ow_15_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8327 ), .force_10(
        \filter_0/n8328 ), .force_11(1'b0), .Q(n40354) );
  \**FFGEN**  \filter_0/pre_ow_15_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8331 ), .force_10(
        \filter_0/n8332 ), .force_11(1'b0), .Q(n40287) );
  \**FFGEN**  \filter_0/pre_ow_15_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8335 ), .force_10(
        \filter_0/n8336 ), .force_11(1'b0), .Q(n40320) );
  \**FFGEN**  \filter_0/pre_ow_15_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8339 ), .force_10(
        \filter_0/n8340 ), .force_11(1'b0), .Q(n40257) );
  \**FFGEN**  \filter_0/pre_ow_15_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8343 ), .force_10(
        \filter_0/n8344 ), .force_11(1'b0), .Q(n40286) );
  \**FFGEN**  \filter_0/pre_ow_15_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8347 ), .force_10(
        \filter_0/n8348 ), .force_11(1'b0), .Q(n40239) );
  \**FFGEN**  \filter_0/pre_ow_15_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8351 ), .force_10(
        \filter_0/n8352 ), .force_11(1'b0), .Q(n40256) );
  \**FFGEN**  \filter_0/pre_ow_15_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8355 ), .force_10(
        \filter_0/n8356 ), .force_11(1'b0), .Q(n40232) );
  \**FFGEN**  \filter_0/pre_ow_15_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8359 ), .force_10(
        \filter_0/n8360 ), .force_11(1'b0), .Q(n40238) );
  \**FFGEN**  \filter_0/pre_ow_15_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8363 ), .force_10(
        \filter_0/n8364 ), .force_11(1'b0), .Q(n40229) );
  \**FFGEN**  \filter_0/pre_ow_15_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8367 ), .force_10(
        \filter_0/n8368 ), .force_11(1'b0), .Q(n40228) );
  \**FFGEN**  \filter_0/pre_ow_14_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8371 ), .force_10(
        \filter_0/n8372 ), .force_11(1'b0), .Q(n40785) );
  \**FFGEN**  \filter_0/pre_ow_14_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8375 ), .force_10(
        \filter_0/n8376 ), .force_11(1'b0), .Q(n40784) );
  \**FFGEN**  \filter_0/pre_ow_14_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8379 ), .force_10(
        \filter_0/n8380 ), .force_11(1'b0), .Q(n40783) );
  \**FFGEN**  \filter_0/pre_ow_14_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8383 ), .force_10(
        \filter_0/n8384 ), .force_11(1'b0), .Q(n40782) );
  \**FFGEN**  \filter_0/pre_ow_14_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8387 ), .force_10(
        \filter_0/n8388 ), .force_11(1'b0), .Q(n40781) );
  \**FFGEN**  \filter_0/pre_ow_14_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8391 ), .force_10(
        \filter_0/n8392 ), .force_11(1'b0), .Q(n40780) );
  \**FFGEN**  \filter_0/pre_ow_14_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8395 ), .force_10(
        \filter_0/n8396 ), .force_11(1'b0), .Q(n40779) );
  \**FFGEN**  \filter_0/pre_ow_14_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8399 ), .force_10(
        \filter_0/n8400 ), .force_11(1'b0), .Q(n40778) );
  \**FFGEN**  \filter_0/pre_ow_14_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8403 ), .force_10(
        \filter_0/n8404 ), .force_11(1'b0), .Q(n40482) );
  \**FFGEN**  \filter_0/pre_ow_14_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8407 ), .force_10(
        \filter_0/n8408 ), .force_11(1'b0), .Q(n40450) );
  \**FFGEN**  \filter_0/pre_ow_14_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8411 ), .force_10(
        \filter_0/n8412 ), .force_11(1'b0), .Q(n40419) );
  \**FFGEN**  \filter_0/pre_ow_14_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8415 ), .force_10(
        \filter_0/n8416 ), .force_11(1'b0), .Q(n40387) );
  \**FFGEN**  \filter_0/pre_ow_14_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8419 ), .force_10(
        \filter_0/n8420 ), .force_11(1'b0), .Q(n40353) );
  \**FFGEN**  \filter_0/pre_ow_14_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8423 ), .force_10(
        \filter_0/n8424 ), .force_11(1'b0), .Q(n40777) );
  \**FFGEN**  \filter_0/pre_ow_14_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8427 ), .force_10(
        \filter_0/n8428 ), .force_11(1'b0), .Q(n40319) );
  \**FFGEN**  \filter_0/pre_ow_14_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8431 ), .force_10(
        \filter_0/n8432 ), .force_11(1'b0), .Q(n40285) );
  \**FFGEN**  \filter_0/pre_ow_14_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8435 ), .force_10(
        \filter_0/n8436 ), .force_11(1'b0), .Q(n40776) );
  \**FFGEN**  \filter_0/pre_ow_14_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8439 ), .force_10(
        \filter_0/n8440 ), .force_11(1'b0), .Q(n40775) );
  \**FFGEN**  \filter_0/pre_ow_14_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8443 ), .force_10(
        \filter_0/n8444 ), .force_11(1'b0), .Q(n40255) );
  \**FFGEN**  \filter_0/pre_ow_14_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8447 ), .force_10(
        \filter_0/n8448 ), .force_11(1'b0), .Q(n40237) );
  \**FFGEN**  \filter_0/pre_ow_13_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8451 ), .force_10(
        \filter_0/n8452 ), .force_11(1'b0), .Q(n40796) );
  \**FFGEN**  \filter_0/pre_ow_13_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8455 ), .force_10(
        \filter_0/n8456 ), .force_11(1'b0), .Q(n40795) );
  \**FFGEN**  \filter_0/pre_ow_13_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8459 ), .force_10(
        \filter_0/n8460 ), .force_11(1'b0), .Q(n40794) );
  \**FFGEN**  \filter_0/pre_ow_13_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8463 ), .force_10(
        \filter_0/n8464 ), .force_11(1'b0), .Q(n40793) );
  \**FFGEN**  \filter_0/pre_ow_13_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8467 ), .force_10(
        \filter_0/n8468 ), .force_11(1'b0), .Q(n40792) );
  \**FFGEN**  \filter_0/pre_ow_13_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8471 ), .force_10(
        \filter_0/n8472 ), .force_11(1'b0), .Q(n40791) );
  \**FFGEN**  \filter_0/pre_ow_13_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8475 ), .force_10(
        \filter_0/n8476 ), .force_11(1'b0), .Q(n40790) );
  \**FFGEN**  \filter_0/pre_ow_13_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8479 ), .force_10(
        \filter_0/n8480 ), .force_11(1'b0), .Q(n40789) );
  \**FFGEN**  \filter_0/pre_ow_13_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8483 ), .force_10(
        \filter_0/n8484 ), .force_11(1'b0), .Q(n40481) );
  \**FFGEN**  \filter_0/pre_ow_13_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8487 ), .force_10(
        \filter_0/n8488 ), .force_11(1'b0), .Q(n40449) );
  \**FFGEN**  \filter_0/pre_ow_13_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8491 ), .force_10(
        \filter_0/n8492 ), .force_11(1'b0), .Q(n40418) );
  \**FFGEN**  \filter_0/pre_ow_13_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8495 ), .force_10(
        \filter_0/n8496 ), .force_11(1'b0), .Q(n40788) );
  \**FFGEN**  \filter_0/pre_ow_13_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8499 ), .force_10(
        \filter_0/n8500 ), .force_11(1'b0), .Q(n40386) );
  \**FFGEN**  \filter_0/pre_ow_13_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8503 ), .force_10(
        \filter_0/n8504 ), .force_11(1'b0), .Q(n40787) );
  \**FFGEN**  \filter_0/pre_ow_13_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8507 ), .force_10(
        \filter_0/n8508 ), .force_11(1'b0), .Q(n40352) );
  \**FFGEN**  \filter_0/pre_ow_13_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8511 ), .force_10(
        \filter_0/n8512 ), .force_11(1'b0), .Q(n40318) );
  \**FFGEN**  \filter_0/pre_ow_13_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8515 ), .force_10(
        \filter_0/n8516 ), .force_11(1'b0), .Q(n40786) );
  \**FFGEN**  \filter_0/pre_ow_13_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8519 ), .force_10(
        \filter_0/n8520 ), .force_11(1'b0), .Q(n40284) );
  \**FFGEN**  \filter_0/pre_ow_13_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8523 ), .force_10(
        \filter_0/n8524 ), .force_11(1'b0), .Q(n40254) );
  \**FFGEN**  \filter_0/pre_ow_13_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8527 ), .force_10(
        \filter_0/n8528 ), .force_11(1'b0), .Q(n40236) );
  \**FFGEN**  \filter_0/pre_ow_12_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8531 ), .force_10(
        \filter_0/n8532 ), .force_11(1'b0), .Q(n40808) );
  \**FFGEN**  \filter_0/pre_ow_12_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8535 ), .force_10(
        \filter_0/n8536 ), .force_11(1'b0), .Q(n40807) );
  \**FFGEN**  \filter_0/pre_ow_12_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8539 ), .force_10(
        \filter_0/n8540 ), .force_11(1'b0), .Q(n40806) );
  \**FFGEN**  \filter_0/pre_ow_12_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8543 ), .force_10(
        \filter_0/n8544 ), .force_11(1'b0), .Q(n40805) );
  \**FFGEN**  \filter_0/pre_ow_12_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8547 ), .force_10(
        \filter_0/n8548 ), .force_11(1'b0), .Q(n40804) );
  \**FFGEN**  \filter_0/pre_ow_12_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8551 ), .force_10(
        \filter_0/n8552 ), .force_11(1'b0), .Q(n40803) );
  \**FFGEN**  \filter_0/pre_ow_12_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8555 ), .force_10(
        \filter_0/n8556 ), .force_11(1'b0), .Q(n40802) );
  \**FFGEN**  \filter_0/pre_ow_12_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8559 ), .force_10(
        \filter_0/n8560 ), .force_11(1'b0), .Q(n40801) );
  \**FFGEN**  \filter_0/pre_ow_12_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8563 ), .force_10(
        \filter_0/n8564 ), .force_11(1'b0), .Q(n40800) );
  \**FFGEN**  \filter_0/pre_ow_12_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8567 ), .force_10(
        \filter_0/n8568 ), .force_11(1'b0), .Q(n40480) );
  \**FFGEN**  \filter_0/pre_ow_12_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8571 ), .force_10(
        \filter_0/n8572 ), .force_11(1'b0), .Q(n40448) );
  \**FFGEN**  \filter_0/pre_ow_12_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8575 ), .force_10(
        \filter_0/n8576 ), .force_11(1'b0), .Q(n40417) );
  \**FFGEN**  \filter_0/pre_ow_12_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8579 ), .force_10(
        \filter_0/n8580 ), .force_11(1'b0), .Q(n40385) );
  \**FFGEN**  \filter_0/pre_ow_12_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8583 ), .force_10(
        \filter_0/n8584 ), .force_11(1'b0), .Q(n40799) );
  \**FFGEN**  \filter_0/pre_ow_12_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8587 ), .force_10(
        \filter_0/n8588 ), .force_11(1'b0), .Q(n40351) );
  \**FFGEN**  \filter_0/pre_ow_12_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8591 ), .force_10(
        \filter_0/n8592 ), .force_11(1'b0), .Q(n40317) );
  \**FFGEN**  \filter_0/pre_ow_12_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8595 ), .force_10(
        \filter_0/n8596 ), .force_11(1'b0), .Q(n40798) );
  \**FFGEN**  \filter_0/pre_ow_12_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8599 ), .force_10(
        \filter_0/n8600 ), .force_11(1'b0), .Q(n40797) );
  \**FFGEN**  \filter_0/pre_ow_12_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8603 ), .force_10(
        \filter_0/n8604 ), .force_11(1'b0), .Q(n40283) );
  \**FFGEN**  \filter_0/pre_ow_12_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8607 ), .force_10(
        \filter_0/n8608 ), .force_11(1'b0), .Q(n40253) );
  \**FFGEN**  \filter_0/pre_ow_11_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8611 ), .force_10(
        \filter_0/n8612 ), .force_11(1'b0), .Q(n40820) );
  \**FFGEN**  \filter_0/pre_ow_11_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8615 ), .force_10(
        \filter_0/n8616 ), .force_11(1'b0), .Q(n40819) );
  \**FFGEN**  \filter_0/pre_ow_11_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8619 ), .force_10(
        \filter_0/n8620 ), .force_11(1'b0), .Q(n40818) );
  \**FFGEN**  \filter_0/pre_ow_11_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8623 ), .force_10(
        \filter_0/n8624 ), .force_11(1'b0), .Q(n40817) );
  \**FFGEN**  \filter_0/pre_ow_11_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8627 ), .force_10(
        \filter_0/n8628 ), .force_11(1'b0), .Q(n40816) );
  \**FFGEN**  \filter_0/pre_ow_11_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8631 ), .force_10(
        \filter_0/n8632 ), .force_11(1'b0), .Q(n40815) );
  \**FFGEN**  \filter_0/pre_ow_11_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8635 ), .force_10(
        \filter_0/n8636 ), .force_11(1'b0), .Q(n40479) );
  \**FFGEN**  \filter_0/pre_ow_11_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8639 ), .force_10(
        \filter_0/n8640 ), .force_11(1'b0), .Q(n40447) );
  \**FFGEN**  \filter_0/pre_ow_11_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8643 ), .force_10(
        \filter_0/n8644 ), .force_11(1'b0), .Q(n40814) );
  \**FFGEN**  \filter_0/pre_ow_11_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8647 ), .force_10(
        \filter_0/n8648 ), .force_11(1'b0), .Q(n40416) );
  \**FFGEN**  \filter_0/pre_ow_11_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8651 ), .force_10(
        \filter_0/n8652 ), .force_11(1'b0), .Q(n40813) );
  \**FFGEN**  \filter_0/pre_ow_11_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8655 ), .force_10(
        \filter_0/n8656 ), .force_11(1'b0), .Q(n40384) );
  \**FFGEN**  \filter_0/pre_ow_11_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8659 ), .force_10(
        \filter_0/n8660 ), .force_11(1'b0), .Q(n40812) );
  \**FFGEN**  \filter_0/pre_ow_11_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8663 ), .force_10(
        \filter_0/n8664 ), .force_11(1'b0), .Q(n40350) );
  \**FFGEN**  \filter_0/pre_ow_11_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8667 ), .force_10(
        \filter_0/n8668 ), .force_11(1'b0), .Q(n40811) );
  \**FFGEN**  \filter_0/pre_ow_11_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8671 ), .force_10(
        \filter_0/n8672 ), .force_11(1'b0), .Q(n40316) );
  \**FFGEN**  \filter_0/pre_ow_11_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8675 ), .force_10(
        \filter_0/n8676 ), .force_11(1'b0), .Q(n40810) );
  \**FFGEN**  \filter_0/pre_ow_11_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8679 ), .force_10(
        \filter_0/n8680 ), .force_11(1'b0), .Q(n40282) );
  \**FFGEN**  \filter_0/pre_ow_11_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8683 ), .force_10(
        \filter_0/n8684 ), .force_11(1'b0), .Q(n40809) );
  \**FFGEN**  \filter_0/pre_ow_11_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8687 ), .force_10(
        \filter_0/n8688 ), .force_11(1'b0), .Q(n40252) );
  \**FFGEN**  \filter_0/pre_ow_10_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8691 ), .force_10(
        \filter_0/n8692 ), .force_11(1'b0), .Q(n40831) );
  \**FFGEN**  \filter_0/pre_ow_10_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8695 ), .force_10(
        \filter_0/n8696 ), .force_11(1'b0), .Q(n40830) );
  \**FFGEN**  \filter_0/pre_ow_10_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8699 ), .force_10(
        \filter_0/n8700 ), .force_11(1'b0), .Q(n40829) );
  \**FFGEN**  \filter_0/pre_ow_10_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8703 ), .force_10(
        \filter_0/n8704 ), .force_11(1'b0), .Q(n40828) );
  \**FFGEN**  \filter_0/pre_ow_10_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8707 ), .force_10(
        \filter_0/n8708 ), .force_11(1'b0), .Q(n40827) );
  \**FFGEN**  \filter_0/pre_ow_10_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8711 ), .force_10(
        \filter_0/n8712 ), .force_11(1'b0), .Q(n40826) );
  \**FFGEN**  \filter_0/pre_ow_10_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8715 ), .force_10(
        \filter_0/n8716 ), .force_11(1'b0), .Q(n40825) );
  \**FFGEN**  \filter_0/pre_ow_10_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8719 ), .force_10(
        \filter_0/n8720 ), .force_11(1'b0), .Q(n40824) );
  \**FFGEN**  \filter_0/pre_ow_10_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8723 ), .force_10(
        \filter_0/n8724 ), .force_11(1'b0), .Q(n40478) );
  \**FFGEN**  \filter_0/pre_ow_10_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8727 ), .force_10(
        \filter_0/n8728 ), .force_11(1'b0), .Q(n40446) );
  \**FFGEN**  \filter_0/pre_ow_10_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8731 ), .force_10(
        \filter_0/n8732 ), .force_11(1'b0), .Q(n40415) );
  \**FFGEN**  \filter_0/pre_ow_10_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8735 ), .force_10(
        \filter_0/n8736 ), .force_11(1'b0), .Q(n40383) );
  \**FFGEN**  \filter_0/pre_ow_10_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8739 ), .force_10(
        \filter_0/n8740 ), .force_11(1'b0), .Q(n40349) );
  \**FFGEN**  \filter_0/pre_ow_10_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8743 ), .force_10(
        \filter_0/n8744 ), .force_11(1'b0), .Q(n40823) );
  \**FFGEN**  \filter_0/pre_ow_10_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8747 ), .force_10(
        \filter_0/n8748 ), .force_11(1'b0), .Q(n40315) );
  \**FFGEN**  \filter_0/pre_ow_10_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8751 ), .force_10(
        \filter_0/n8752 ), .force_11(1'b0), .Q(n40281) );
  \**FFGEN**  \filter_0/pre_ow_10_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8755 ), .force_10(
        \filter_0/n8756 ), .force_11(1'b0), .Q(n40822) );
  \**FFGEN**  \filter_0/pre_ow_10_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8759 ), .force_10(
        \filter_0/n8760 ), .force_11(1'b0), .Q(n40821) );
  \**FFGEN**  \filter_0/pre_ow_10_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8763 ), .force_10(
        \filter_0/n8764 ), .force_11(1'b0), .Q(n40251) );
  \**FFGEN**  \filter_0/pre_ow_10_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8767 ), .force_10(
        \filter_0/n8768 ), .force_11(1'b0), .Q(n40235) );
  \**FFGEN**  \filter_0/pre_ow_9_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8771 ), .force_10(
        \filter_0/n8772 ), .force_11(1'b0), .Q(n40842) );
  \**FFGEN**  \filter_0/pre_ow_9_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8775 ), .force_10(
        \filter_0/n8776 ), .force_11(1'b0), .Q(n40841) );
  \**FFGEN**  \filter_0/pre_ow_9_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8779 ), .force_10(
        \filter_0/n8780 ), .force_11(1'b0), .Q(n40840) );
  \**FFGEN**  \filter_0/pre_ow_9_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8783 ), .force_10(
        \filter_0/n8784 ), .force_11(1'b0), .Q(n40839) );
  \**FFGEN**  \filter_0/pre_ow_9_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8787 ), .force_10(
        \filter_0/n8788 ), .force_11(1'b0), .Q(n40838) );
  \**FFGEN**  \filter_0/pre_ow_9_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8791 ), .force_10(
        \filter_0/n8792 ), .force_11(1'b0), .Q(n40837) );
  \**FFGEN**  \filter_0/pre_ow_9_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8795 ), .force_10(
        \filter_0/n8796 ), .force_11(1'b0), .Q(n40836) );
  \**FFGEN**  \filter_0/pre_ow_9_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8799 ), .force_10(
        \filter_0/n8800 ), .force_11(1'b0), .Q(n40835) );
  \**FFGEN**  \filter_0/pre_ow_9_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8803 ), .force_10(
        \filter_0/n8804 ), .force_11(1'b0), .Q(n40477) );
  \**FFGEN**  \filter_0/pre_ow_9_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8807 ), .force_10(
        \filter_0/n8808 ), .force_11(1'b0), .Q(n40445) );
  \**FFGEN**  \filter_0/pre_ow_9_reg[9]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n8811 ), .force_10(\filter_0/n8812 ), 
        .force_11(1'b0), .Q(n40414) );
  \**FFGEN**  \filter_0/pre_ow_9_reg[8]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n8815 ), .force_10(\filter_0/n8816 ), 
        .force_11(1'b0), .Q(n40382) );
  \**FFGEN**  \filter_0/pre_ow_9_reg[7]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n8819 ), .force_10(\filter_0/n8820 ), 
        .force_11(1'b0), .Q(n40348) );
  \**FFGEN**  \filter_0/pre_ow_9_reg[6]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n8823 ), .force_10(\filter_0/n8824 ), 
        .force_11(1'b0), .Q(n40834) );
  \**FFGEN**  \filter_0/pre_ow_9_reg[5]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n8827 ), .force_10(\filter_0/n8828 ), 
        .force_11(1'b0), .Q(n40314) );
  \**FFGEN**  \filter_0/pre_ow_9_reg[4]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n8831 ), .force_10(\filter_0/n8832 ), 
        .force_11(1'b0), .Q(n40280) );
  \**FFGEN**  \filter_0/pre_ow_9_reg[3]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n8835 ), .force_10(\filter_0/n8836 ), 
        .force_11(1'b0), .Q(n40833) );
  \**FFGEN**  \filter_0/pre_ow_9_reg[2]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n8839 ), .force_10(\filter_0/n8840 ), 
        .force_11(1'b0), .Q(n40832) );
  \**FFGEN**  \filter_0/pre_ow_9_reg[1]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n8843 ), .force_10(\filter_0/n8844 ), 
        .force_11(1'b0), .Q(n40250) );
  \**FFGEN**  \filter_0/pre_ow_9_reg[0]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n8847 ), .force_10(\filter_0/n8848 ), 
        .force_11(1'b0), .Q(n40234) );
  \**FFGEN**  \filter_0/pre_ow_8_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8851 ), .force_10(
        \filter_0/n8852 ), .force_11(1'b0), .Q(n40854) );
  \**FFGEN**  \filter_0/pre_ow_8_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8855 ), .force_10(
        \filter_0/n8856 ), .force_11(1'b0), .Q(n40853) );
  \**FFGEN**  \filter_0/pre_ow_8_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8859 ), .force_10(
        \filter_0/n8860 ), .force_11(1'b0), .Q(n40852) );
  \**FFGEN**  \filter_0/pre_ow_8_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8863 ), .force_10(
        \filter_0/n8864 ), .force_11(1'b0), .Q(n40851) );
  \**FFGEN**  \filter_0/pre_ow_8_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8867 ), .force_10(
        \filter_0/n8868 ), .force_11(1'b0), .Q(n40850) );
  \**FFGEN**  \filter_0/pre_ow_8_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8871 ), .force_10(
        \filter_0/n8872 ), .force_11(1'b0), .Q(n40849) );
  \**FFGEN**  \filter_0/pre_ow_8_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8875 ), .force_10(
        \filter_0/n8876 ), .force_11(1'b0), .Q(n40848) );
  \**FFGEN**  \filter_0/pre_ow_8_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8879 ), .force_10(
        \filter_0/n8880 ), .force_11(1'b0), .Q(n40847) );
  \**FFGEN**  \filter_0/pre_ow_8_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8883 ), .force_10(
        \filter_0/n8884 ), .force_11(1'b0), .Q(n40846) );
  \**FFGEN**  \filter_0/pre_ow_8_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8887 ), .force_10(
        \filter_0/n8888 ), .force_11(1'b0), .Q(n40476) );
  \**FFGEN**  \filter_0/pre_ow_8_reg[9]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n8891 ), .force_10(\filter_0/n8892 ), 
        .force_11(1'b0), .Q(n40444) );
  \**FFGEN**  \filter_0/pre_ow_8_reg[8]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n8895 ), .force_10(\filter_0/n8896 ), 
        .force_11(1'b0), .Q(n40845) );
  \**FFGEN**  \filter_0/pre_ow_8_reg[7]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n8899 ), .force_10(\filter_0/n8900 ), 
        .force_11(1'b0), .Q(n40413) );
  \**FFGEN**  \filter_0/pre_ow_8_reg[6]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n8903 ), .force_10(\filter_0/n8904 ), 
        .force_11(1'b0), .Q(n40844) );
  \**FFGEN**  \filter_0/pre_ow_8_reg[5]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n8907 ), .force_10(\filter_0/n8908 ), 
        .force_11(1'b0), .Q(n40381) );
  \**FFGEN**  \filter_0/pre_ow_8_reg[4]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n8911 ), .force_10(\filter_0/n8912 ), 
        .force_11(1'b0), .Q(n40347) );
  \**FFGEN**  \filter_0/pre_ow_8_reg[3]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n8915 ), .force_10(\filter_0/n8916 ), 
        .force_11(1'b0), .Q(n40843) );
  \**FFGEN**  \filter_0/pre_ow_8_reg[2]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n8919 ), .force_10(\filter_0/n8920 ), 
        .force_11(1'b0), .Q(n40313) );
  \**FFGEN**  \filter_0/pre_ow_8_reg[1]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n8923 ), .force_10(\filter_0/n8924 ), 
        .force_11(1'b0), .Q(n40279) );
  \**FFGEN**  \filter_0/pre_ow_8_reg[0]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n8927 ), .force_10(\filter_0/n8928 ), 
        .force_11(1'b0), .Q(n40249) );
  \**FFGEN**  \filter_0/pre_ow_7_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8931 ), .force_10(
        \filter_0/n8932 ), .force_11(1'b0), .Q(n40770) );
  \**FFGEN**  \filter_0/pre_ow_7_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8935 ), .force_10(
        \filter_0/n8936 ), .force_11(1'b0), .Q(n40769) );
  \**FFGEN**  \filter_0/pre_ow_7_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8939 ), .force_10(
        \filter_0/n8940 ), .force_11(1'b0), .Q(n40768) );
  \**FFGEN**  \filter_0/pre_ow_7_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8943 ), .force_10(
        \filter_0/n8944 ), .force_11(1'b0), .Q(n40484) );
  \**FFGEN**  \filter_0/pre_ow_7_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8947 ), .force_10(
        \filter_0/n8948 ), .force_11(1'b0), .Q(n40767) );
  \**FFGEN**  \filter_0/pre_ow_7_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8951 ), .force_10(
        \filter_0/n8952 ), .force_11(1'b0), .Q(n40766) );
  \**FFGEN**  \filter_0/pre_ow_7_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8955 ), .force_10(
        \filter_0/n8956 ), .force_11(1'b0), .Q(n40452) );
  \**FFGEN**  \filter_0/pre_ow_7_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8959 ), .force_10(
        \filter_0/n8960 ), .force_11(1'b0), .Q(n40421) );
  \**FFGEN**  \filter_0/pre_ow_7_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8963 ), .force_10(
        \filter_0/n8964 ), .force_11(1'b0), .Q(n40765) );
  \**FFGEN**  \filter_0/pre_ow_7_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n8967 ), .force_10(
        \filter_0/n8968 ), .force_11(1'b0), .Q(n40388) );
  \**FFGEN**  \filter_0/pre_ow_7_reg[9]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n8971 ), .force_10(\filter_0/n8972 ), 
        .force_11(1'b0), .Q(n40764) );
  \**FFGEN**  \filter_0/pre_ow_7_reg[8]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n8975 ), .force_10(\filter_0/n8976 ), 
        .force_11(1'b0), .Q(n40356) );
  \**FFGEN**  \filter_0/pre_ow_7_reg[7]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n8979 ), .force_10(\filter_0/n8980 ), 
        .force_11(1'b0), .Q(n40763) );
  \**FFGEN**  \filter_0/pre_ow_7_reg[6]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n8983 ), .force_10(\filter_0/n8984 ), 
        .force_11(1'b0), .Q(n40322) );
  \**FFGEN**  \filter_0/pre_ow_7_reg[5]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n8987 ), .force_10(\filter_0/n8988 ), 
        .force_11(1'b0), .Q(n40762) );
  \**FFGEN**  \filter_0/pre_ow_7_reg[4]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n8991 ), .force_10(\filter_0/n8992 ), 
        .force_11(1'b0), .Q(n40288) );
  \**FFGEN**  \filter_0/pre_ow_7_reg[3]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n8995 ), .force_10(\filter_0/n8996 ), 
        .force_11(1'b0), .Q(n40761) );
  \**FFGEN**  \filter_0/pre_ow_7_reg[2]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n8999 ), .force_10(\filter_0/n9000 ), 
        .force_11(1'b0), .Q(n40258) );
  \**FFGEN**  \filter_0/pre_ow_7_reg[1]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n9003 ), .force_10(\filter_0/n9004 ), 
        .force_11(1'b0), .Q(n40760) );
  \**FFGEN**  \filter_0/pre_ow_7_reg[0]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n9007 ), .force_10(\filter_0/n9008 ), 
        .force_11(1'b0), .Q(n40240) );
  \**FFGEN**  \filter_0/pre_ow_6_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9011 ), .force_10(
        \filter_0/n9012 ), .force_11(1'b0), .Q(n40759) );
  \**FFGEN**  \filter_0/pre_ow_6_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9015 ), .force_10(
        \filter_0/n9016 ), .force_11(1'b0), .Q(n40758) );
  \**FFGEN**  \filter_0/pre_ow_6_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9019 ), .force_10(
        \filter_0/n9020 ), .force_11(1'b0), .Q(n40757) );
  \**FFGEN**  \filter_0/pre_ow_6_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9023 ), .force_10(
        \filter_0/n9024 ), .force_11(1'b0), .Q(n40756) );
  \**FFGEN**  \filter_0/pre_ow_6_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9027 ), .force_10(
        \filter_0/n9028 ), .force_11(1'b0), .Q(n40755) );
  \**FFGEN**  \filter_0/pre_ow_6_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9031 ), .force_10(
        \filter_0/n9032 ), .force_11(1'b0), .Q(n40754) );
  \**FFGEN**  \filter_0/pre_ow_6_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9035 ), .force_10(
        \filter_0/n9036 ), .force_11(1'b0), .Q(n40753) );
  \**FFGEN**  \filter_0/pre_ow_6_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9039 ), .force_10(
        \filter_0/n9040 ), .force_11(1'b0), .Q(n40752) );
  \**FFGEN**  \filter_0/pre_ow_6_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9043 ), .force_10(
        \filter_0/n9044 ), .force_11(1'b0), .Q(n40751) );
  \**FFGEN**  \filter_0/pre_ow_6_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9047 ), .force_10(
        \filter_0/n9048 ), .force_11(1'b0), .Q(n40485) );
  \**FFGEN**  \filter_0/pre_ow_6_reg[9]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n9051 ), .force_10(\filter_0/n9052 ), 
        .force_11(1'b0), .Q(n40453) );
  \**FFGEN**  \filter_0/pre_ow_6_reg[8]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n9055 ), .force_10(\filter_0/n9056 ), 
        .force_11(1'b0), .Q(n40750) );
  \**FFGEN**  \filter_0/pre_ow_6_reg[7]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n9059 ), .force_10(\filter_0/n9060 ), 
        .force_11(1'b0), .Q(n40422) );
  \**FFGEN**  \filter_0/pre_ow_6_reg[6]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n9063 ), .force_10(\filter_0/n9064 ), 
        .force_11(1'b0), .Q(n40749) );
  \**FFGEN**  \filter_0/pre_ow_6_reg[5]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n9067 ), .force_10(\filter_0/n9068 ), 
        .force_11(1'b0), .Q(n40389) );
  \**FFGEN**  \filter_0/pre_ow_6_reg[4]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n9071 ), .force_10(\filter_0/n9072 ), 
        .force_11(1'b0), .Q(n40357) );
  \**FFGEN**  \filter_0/pre_ow_6_reg[3]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n9075 ), .force_10(\filter_0/n9076 ), 
        .force_11(1'b0), .Q(n40748) );
  \**FFGEN**  \filter_0/pre_ow_6_reg[2]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n9079 ), .force_10(\filter_0/n9080 ), 
        .force_11(1'b0), .Q(n40323) );
  \**FFGEN**  \filter_0/pre_ow_6_reg[1]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n9083 ), .force_10(\filter_0/n9084 ), 
        .force_11(1'b0), .Q(n40289) );
  \**FFGEN**  \filter_0/pre_ow_6_reg[0]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n9087 ), .force_10(\filter_0/n9088 ), 
        .force_11(1'b0), .Q(n40259) );
  \**FFGEN**  \filter_0/pre_ow_5_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9091 ), .force_10(
        \filter_0/n9092 ), .force_11(1'b0), .Q(n40747) );
  \**FFGEN**  \filter_0/pre_ow_5_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9095 ), .force_10(
        \filter_0/n9096 ), .force_11(1'b0), .Q(n40746) );
  \**FFGEN**  \filter_0/pre_ow_5_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9099 ), .force_10(
        \filter_0/n9100 ), .force_11(1'b0), .Q(n40745) );
  \**FFGEN**  \filter_0/pre_ow_5_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9103 ), .force_10(
        \filter_0/n9104 ), .force_11(1'b0), .Q(n40744) );
  \**FFGEN**  \filter_0/pre_ow_5_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9107 ), .force_10(
        \filter_0/n9108 ), .force_11(1'b0), .Q(n40743) );
  \**FFGEN**  \filter_0/pre_ow_5_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9111 ), .force_10(
        \filter_0/n9112 ), .force_11(1'b0), .Q(n40742) );
  \**FFGEN**  \filter_0/pre_ow_5_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9115 ), .force_10(
        \filter_0/n9116 ), .force_11(1'b0), .Q(n40741) );
  \**FFGEN**  \filter_0/pre_ow_5_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9119 ), .force_10(
        \filter_0/n9120 ), .force_11(1'b0), .Q(n40740) );
  \**FFGEN**  \filter_0/pre_ow_5_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9123 ), .force_10(
        \filter_0/n9124 ), .force_11(1'b0), .Q(n40739) );
  \**FFGEN**  \filter_0/pre_ow_5_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9127 ), .force_10(
        \filter_0/n9128 ), .force_11(1'b0), .Q(n40486) );
  \**FFGEN**  \filter_0/pre_ow_5_reg[9]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n9131 ), .force_10(\filter_0/n9132 ), 
        .force_11(1'b0), .Q(n40454) );
  \**FFGEN**  \filter_0/pre_ow_5_reg[8]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n9135 ), .force_10(\filter_0/n9136 ), 
        .force_11(1'b0), .Q(n40423) );
  \**FFGEN**  \filter_0/pre_ow_5_reg[7]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n9139 ), .force_10(\filter_0/n9140 ), 
        .force_11(1'b0), .Q(n40390) );
  \**FFGEN**  \filter_0/pre_ow_5_reg[6]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n9143 ), .force_10(\filter_0/n9144 ), 
        .force_11(1'b0), .Q(n40738) );
  \**FFGEN**  \filter_0/pre_ow_5_reg[5]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n9147 ), .force_10(\filter_0/n9148 ), 
        .force_11(1'b0), .Q(n40358) );
  \**FFGEN**  \filter_0/pre_ow_5_reg[4]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n9151 ), .force_10(\filter_0/n9152 ), 
        .force_11(1'b0), .Q(n40324) );
  \**FFGEN**  \filter_0/pre_ow_5_reg[3]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n9155 ), .force_10(\filter_0/n9156 ), 
        .force_11(1'b0), .Q(n40737) );
  \**FFGEN**  \filter_0/pre_ow_5_reg[2]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n9159 ), .force_10(\filter_0/n9160 ), 
        .force_11(1'b0), .Q(n40736) );
  \**FFGEN**  \filter_0/pre_ow_5_reg[1]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n9163 ), .force_10(\filter_0/n9164 ), 
        .force_11(1'b0), .Q(n40290) );
  \**FFGEN**  \filter_0/pre_ow_5_reg[0]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n9167 ), .force_10(\filter_0/n9168 ), 
        .force_11(1'b0), .Q(n40260) );
  \**FFGEN**  \filter_0/pre_ow_4_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9171 ), .force_10(
        \filter_0/n9172 ), .force_11(1'b0), .Q(n40735) );
  \**FFGEN**  \filter_0/pre_ow_4_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9175 ), .force_10(
        \filter_0/n9176 ), .force_11(1'b0), .Q(n40734) );
  \**FFGEN**  \filter_0/pre_ow_4_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9179 ), .force_10(
        \filter_0/n9180 ), .force_11(1'b0), .Q(n40733) );
  \**FFGEN**  \filter_0/pre_ow_4_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9183 ), .force_10(
        \filter_0/n9184 ), .force_11(1'b0), .Q(n40732) );
  \**FFGEN**  \filter_0/pre_ow_4_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9187 ), .force_10(
        \filter_0/n9188 ), .force_11(1'b0), .Q(n40731) );
  \**FFGEN**  \filter_0/pre_ow_4_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9191 ), .force_10(
        \filter_0/n9192 ), .force_11(1'b0), .Q(n40730) );
  \**FFGEN**  \filter_0/pre_ow_4_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9195 ), .force_10(
        \filter_0/n9196 ), .force_11(1'b0), .Q(n40729) );
  \**FFGEN**  \filter_0/pre_ow_4_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9199 ), .force_10(
        \filter_0/n9200 ), .force_11(1'b0), .Q(n40728) );
  \**FFGEN**  \filter_0/pre_ow_4_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9203 ), .force_10(
        \filter_0/n9204 ), .force_11(1'b0), .Q(n40727) );
  \**FFGEN**  \filter_0/pre_ow_4_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9207 ), .force_10(
        \filter_0/n9208 ), .force_11(1'b0), .Q(n40726) );
  \**FFGEN**  \filter_0/pre_ow_4_reg[9]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n9211 ), .force_10(\filter_0/n9212 ), 
        .force_11(1'b0), .Q(n40487) );
  \**FFGEN**  \filter_0/pre_ow_4_reg[8]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n9215 ), .force_10(\filter_0/n9216 ), 
        .force_11(1'b0), .Q(n40455) );
  \**FFGEN**  \filter_0/pre_ow_4_reg[7]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n9219 ), .force_10(\filter_0/n9220 ), 
        .force_11(1'b0), .Q(n40424) );
  \**FFGEN**  \filter_0/pre_ow_4_reg[6]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n9223 ), .force_10(\filter_0/n9224 ), 
        .force_11(1'b0), .Q(n40725) );
  \**FFGEN**  \filter_0/pre_ow_4_reg[5]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n9227 ), .force_10(\filter_0/n9228 ), 
        .force_11(1'b0), .Q(n40391) );
  \**FFGEN**  \filter_0/pre_ow_4_reg[4]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n9231 ), .force_10(\filter_0/n9232 ), 
        .force_11(1'b0), .Q(n40359) );
  \**FFGEN**  \filter_0/pre_ow_4_reg[3]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n9235 ), .force_10(\filter_0/n9236 ), 
        .force_11(1'b0), .Q(n40724) );
  \**FFGEN**  \filter_0/pre_ow_4_reg[2]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n9239 ), .force_10(\filter_0/n9240 ), 
        .force_11(1'b0), .Q(n40723) );
  \**FFGEN**  \filter_0/pre_ow_4_reg[1]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n9243 ), .force_10(\filter_0/n9244 ), 
        .force_11(1'b0), .Q(n40325) );
  \**FFGEN**  \filter_0/pre_ow_4_reg[0]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n9247 ), .force_10(\filter_0/n9248 ), 
        .force_11(1'b0), .Q(n40291) );
  \**FFGEN**  \filter_0/pre_ow_3_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9251 ), .force_10(
        \filter_0/n9252 ), .force_11(1'b0), .Q(n40722) );
  \**FFGEN**  \filter_0/pre_ow_3_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9255 ), .force_10(
        \filter_0/n9256 ), .force_11(1'b0), .Q(n40721) );
  \**FFGEN**  \filter_0/pre_ow_3_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9259 ), .force_10(
        \filter_0/n9260 ), .force_11(1'b0), .Q(n40720) );
  \**FFGEN**  \filter_0/pre_ow_3_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9263 ), .force_10(
        \filter_0/n9264 ), .force_11(1'b0), .Q(n40719) );
  \**FFGEN**  \filter_0/pre_ow_3_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9267 ), .force_10(
        \filter_0/n9268 ), .force_11(1'b0), .Q(n40718) );
  \**FFGEN**  \filter_0/pre_ow_3_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9271 ), .force_10(
        \filter_0/n9272 ), .force_11(1'b0), .Q(n40717) );
  \**FFGEN**  \filter_0/pre_ow_3_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9275 ), .force_10(
        \filter_0/n9276 ), .force_11(1'b0), .Q(n40716) );
  \**FFGEN**  \filter_0/pre_ow_3_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9279 ), .force_10(
        \filter_0/n9280 ), .force_11(1'b0), .Q(n40715) );
  \**FFGEN**  \filter_0/pre_ow_3_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9283 ), .force_10(
        \filter_0/n9284 ), .force_11(1'b0), .Q(n40714) );
  \**FFGEN**  \filter_0/pre_ow_3_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9287 ), .force_10(
        \filter_0/n9288 ), .force_11(1'b0), .Q(n40488) );
  \**FFGEN**  \filter_0/pre_ow_3_reg[9]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n9291 ), .force_10(\filter_0/n9292 ), 
        .force_11(1'b0), .Q(n40456) );
  \**FFGEN**  \filter_0/pre_ow_3_reg[8]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n9295 ), .force_10(\filter_0/n9296 ), 
        .force_11(1'b0), .Q(n40425) );
  \**FFGEN**  \filter_0/pre_ow_3_reg[7]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n9299 ), .force_10(\filter_0/n9300 ), 
        .force_11(1'b0), .Q(n40392) );
  \**FFGEN**  \filter_0/pre_ow_3_reg[6]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n9303 ), .force_10(\filter_0/n9304 ), 
        .force_11(1'b0), .Q(n40360) );
  \**FFGEN**  \filter_0/pre_ow_3_reg[5]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n9307 ), .force_10(\filter_0/n9308 ), 
        .force_11(1'b0), .Q(n40713) );
  \**FFGEN**  \filter_0/pre_ow_3_reg[4]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n9311 ), .force_10(\filter_0/n9312 ), 
        .force_11(1'b0), .Q(n40326) );
  \**FFGEN**  \filter_0/pre_ow_3_reg[3]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n9315 ), .force_10(\filter_0/n9316 ), 
        .force_11(1'b0), .Q(n40712) );
  \**FFGEN**  \filter_0/pre_ow_3_reg[2]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n9319 ), .force_10(\filter_0/n9320 ), 
        .force_11(1'b0), .Q(n40292) );
  \**FFGEN**  \filter_0/pre_ow_3_reg[1]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n9323 ), .force_10(\filter_0/n9324 ), 
        .force_11(1'b0), .Q(n40711) );
  \**FFGEN**  \filter_0/pre_ow_3_reg[0]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n9327 ), .force_10(\filter_0/n9328 ), 
        .force_11(1'b0), .Q(n40261) );
  \**FFGEN**  \filter_0/pre_ow_2_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9331 ), .force_10(
        \filter_0/n9332 ), .force_11(1'b0), .Q(n40710) );
  \**FFGEN**  \filter_0/pre_ow_2_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9335 ), .force_10(
        \filter_0/n9336 ), .force_11(1'b0), .Q(n40709) );
  \**FFGEN**  \filter_0/pre_ow_2_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9339 ), .force_10(
        \filter_0/n9340 ), .force_11(1'b0), .Q(n40708) );
  \**FFGEN**  \filter_0/pre_ow_2_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9343 ), .force_10(
        \filter_0/n9344 ), .force_11(1'b0), .Q(n40707) );
  \**FFGEN**  \filter_0/pre_ow_2_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9347 ), .force_10(
        \filter_0/n9348 ), .force_11(1'b0), .Q(n40706) );
  \**FFGEN**  \filter_0/pre_ow_2_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9351 ), .force_10(
        \filter_0/n9352 ), .force_11(1'b0), .Q(n40705) );
  \**FFGEN**  \filter_0/pre_ow_2_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9355 ), .force_10(
        \filter_0/n9356 ), .force_11(1'b0), .Q(n40704) );
  \**FFGEN**  \filter_0/pre_ow_2_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9359 ), .force_10(
        \filter_0/n9360 ), .force_11(1'b0), .Q(n40703) );
  \**FFGEN**  \filter_0/pre_ow_2_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9363 ), .force_10(
        \filter_0/n9364 ), .force_11(1'b0), .Q(n40702) );
  \**FFGEN**  \filter_0/pre_ow_2_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9367 ), .force_10(
        \filter_0/n9368 ), .force_11(1'b0), .Q(n40489) );
  \**FFGEN**  \filter_0/pre_ow_2_reg[9]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n9371 ), .force_10(\filter_0/n9372 ), 
        .force_11(1'b0), .Q(n40457) );
  \**FFGEN**  \filter_0/pre_ow_2_reg[8]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n9375 ), .force_10(\filter_0/n9376 ), 
        .force_11(1'b0), .Q(n40426) );
  \**FFGEN**  \filter_0/pre_ow_2_reg[7]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n9379 ), .force_10(\filter_0/n9380 ), 
        .force_11(1'b0), .Q(n40393) );
  \**FFGEN**  \filter_0/pre_ow_2_reg[6]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n9383 ), .force_10(\filter_0/n9384 ), 
        .force_11(1'b0), .Q(n40701) );
  \**FFGEN**  \filter_0/pre_ow_2_reg[5]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n9387 ), .force_10(\filter_0/n9388 ), 
        .force_11(1'b0), .Q(n40361) );
  \**FFGEN**  \filter_0/pre_ow_2_reg[4]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n9391 ), .force_10(\filter_0/n9392 ), 
        .force_11(1'b0), .Q(n40327) );
  \**FFGEN**  \filter_0/pre_ow_2_reg[3]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n9395 ), .force_10(\filter_0/n9396 ), 
        .force_11(1'b0), .Q(n40700) );
  \**FFGEN**  \filter_0/pre_ow_2_reg[2]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n9399 ), .force_10(\filter_0/n9400 ), 
        .force_11(1'b0), .Q(n40699) );
  \**FFGEN**  \filter_0/pre_ow_2_reg[1]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n9403 ), .force_10(\filter_0/n9404 ), 
        .force_11(1'b0), .Q(n40293) );
  \**FFGEN**  \filter_0/pre_ow_2_reg[0]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n9407 ), .force_10(\filter_0/n9408 ), 
        .force_11(1'b0), .Q(n40262) );
  \**FFGEN**  \filter_0/pre_ow_1_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9411 ), .force_10(
        \filter_0/n9412 ), .force_11(1'b0), .Q(n40698) );
  \**FFGEN**  \filter_0/pre_ow_1_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9415 ), .force_10(
        \filter_0/n9416 ), .force_11(1'b0), .Q(n40697) );
  \**FFGEN**  \filter_0/pre_ow_1_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9419 ), .force_10(
        \filter_0/n9420 ), .force_11(1'b0), .Q(n40696) );
  \**FFGEN**  \filter_0/pre_ow_1_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9423 ), .force_10(
        \filter_0/n9424 ), .force_11(1'b0), .Q(n40695) );
  \**FFGEN**  \filter_0/pre_ow_1_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9427 ), .force_10(
        \filter_0/n9428 ), .force_11(1'b0), .Q(n40694) );
  \**FFGEN**  \filter_0/pre_ow_1_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9431 ), .force_10(
        \filter_0/n9432 ), .force_11(1'b0), .Q(n40693) );
  \**FFGEN**  \filter_0/pre_ow_1_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9435 ), .force_10(
        \filter_0/n9436 ), .force_11(1'b0), .Q(n40692) );
  \**FFGEN**  \filter_0/pre_ow_1_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9439 ), .force_10(
        \filter_0/n9440 ), .force_11(1'b0), .Q(n40691) );
  \**FFGEN**  \filter_0/pre_ow_1_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9443 ), .force_10(
        \filter_0/n9444 ), .force_11(1'b0), .Q(n40690) );
  \**FFGEN**  \filter_0/pre_ow_1_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9447 ), .force_10(
        \filter_0/n9448 ), .force_11(1'b0), .Q(n40490) );
  \**FFGEN**  \filter_0/pre_ow_1_reg[9]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n9451 ), .force_10(\filter_0/n9452 ), 
        .force_11(1'b0), .Q(n40458) );
  \**FFGEN**  \filter_0/pre_ow_1_reg[8]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n9455 ), .force_10(\filter_0/n9456 ), 
        .force_11(1'b0), .Q(n40427) );
  \**FFGEN**  \filter_0/pre_ow_1_reg[7]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n9459 ), .force_10(\filter_0/n9460 ), 
        .force_11(1'b0), .Q(n40394) );
  \**FFGEN**  \filter_0/pre_ow_1_reg[6]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n9463 ), .force_10(\filter_0/n9464 ), 
        .force_11(1'b0), .Q(n40689) );
  \**FFGEN**  \filter_0/pre_ow_1_reg[5]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n9467 ), .force_10(\filter_0/n9468 ), 
        .force_11(1'b0), .Q(n40362) );
  \**FFGEN**  \filter_0/pre_ow_1_reg[4]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n9471 ), .force_10(\filter_0/n9472 ), 
        .force_11(1'b0), .Q(n40328) );
  \**FFGEN**  \filter_0/pre_ow_1_reg[3]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n9475 ), .force_10(\filter_0/n9476 ), 
        .force_11(1'b0), .Q(n40688) );
  \**FFGEN**  \filter_0/pre_ow_1_reg[2]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n9479 ), .force_10(\filter_0/n9480 ), 
        .force_11(1'b0), .Q(n40687) );
  \**FFGEN**  \filter_0/pre_ow_1_reg[1]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n9483 ), .force_10(\filter_0/n9484 ), 
        .force_11(1'b0), .Q(n40294) );
  \**FFGEN**  \filter_0/pre_ow_1_reg[0]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n9487 ), .force_10(\filter_0/n9488 ), 
        .force_11(1'b0), .Q(n40263) );
  \**FFGEN**  \filter_0/pre_ow_0_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9491 ), .force_10(
        \filter_0/n9492 ), .force_11(1'b0), .Q(n40867) );
  \**FFGEN**  \filter_0/pre_ow_0_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9495 ), .force_10(
        \filter_0/n9496 ), .force_11(1'b0), .Q(n40866) );
  \**FFGEN**  \filter_0/pre_ow_0_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9499 ), .force_10(
        \filter_0/n9500 ), .force_11(1'b0), .Q(n40865) );
  \**FFGEN**  \filter_0/pre_ow_0_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9503 ), .force_10(
        \filter_0/n9504 ), .force_11(1'b0), .Q(n40864) );
  \**FFGEN**  \filter_0/pre_ow_0_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9507 ), .force_10(
        \filter_0/n9508 ), .force_11(1'b0), .Q(n40863) );
  \**FFGEN**  \filter_0/pre_ow_0_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9511 ), .force_10(
        \filter_0/n9512 ), .force_11(1'b0), .Q(n40862) );
  \**FFGEN**  \filter_0/pre_ow_0_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9515 ), .force_10(
        \filter_0/n9516 ), .force_11(1'b0), .Q(n40861) );
  \**FFGEN**  \filter_0/pre_ow_0_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9519 ), .force_10(
        \filter_0/n9520 ), .force_11(1'b0), .Q(n40860) );
  \**FFGEN**  \filter_0/pre_ow_0_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9523 ), .force_10(
        \filter_0/n9524 ), .force_11(1'b0), .Q(n40859) );
  \**FFGEN**  \filter_0/pre_ow_0_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9527 ), .force_10(
        \filter_0/n9528 ), .force_11(1'b0), .Q(n40858) );
  \**FFGEN**  \filter_0/pre_ow_0_reg[9]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n9531 ), .force_10(\filter_0/n9532 ), 
        .force_11(1'b0), .Q(n40475) );
  \**FFGEN**  \filter_0/pre_ow_0_reg[8]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n9535 ), .force_10(\filter_0/n9536 ), 
        .force_11(1'b0), .Q(n40857) );
  \**FFGEN**  \filter_0/pre_ow_0_reg[7]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n9539 ), .force_10(\filter_0/n9540 ), 
        .force_11(1'b0), .Q(n40443) );
  \**FFGEN**  \filter_0/pre_ow_0_reg[6]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n9543 ), .force_10(\filter_0/n9544 ), 
        .force_11(1'b0), .Q(n40856) );
  \**FFGEN**  \filter_0/pre_ow_0_reg[5]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n9547 ), .force_10(\filter_0/n9548 ), 
        .force_11(1'b0), .Q(n40412) );
  \**FFGEN**  \filter_0/pre_ow_0_reg[4]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n9551 ), .force_10(\filter_0/n9552 ), 
        .force_11(1'b0), .Q(n40380) );
  \**FFGEN**  \filter_0/pre_ow_0_reg[3]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n9555 ), .force_10(\filter_0/n9556 ), 
        .force_11(1'b0), .Q(n40855) );
  \**FFGEN**  \filter_0/pre_ow_0_reg[2]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n9559 ), .force_10(\filter_0/n9560 ), 
        .force_11(1'b0), .Q(n40346) );
  \**FFGEN**  \filter_0/pre_ow_0_reg[1]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n9563 ), .force_10(\filter_0/n9564 ), 
        .force_11(1'b0), .Q(n40312) );
  \**FFGEN**  \filter_0/pre_ow_0_reg[0]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n9567 ), .force_10(\filter_0/n9568 ), 
        .force_11(1'b0), .Q(n40278) );
  \**FFGEN**  \filter_0/pre_oi_15_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9571 ), .force_10(
        \filter_0/n9572 ), .force_11(1'b0), .Q(n40592) );
  \**FFGEN**  \filter_0/pre_oi_15_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9575 ), .force_10(
        \filter_0/n9576 ), .force_11(1'b0), .Q(n40591) );
  \**FFGEN**  \filter_0/pre_oi_15_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9579 ), .force_10(
        \filter_0/n9580 ), .force_11(1'b0), .Q(n40590) );
  \**FFGEN**  \filter_0/pre_oi_15_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9583 ), .force_10(
        \filter_0/n9584 ), .force_11(1'b0), .Q(n40499) );
  \**FFGEN**  \filter_0/pre_oi_15_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9587 ), .force_10(
        \filter_0/n9588 ), .force_11(1'b0), .Q(n40404) );
  \**FFGEN**  \filter_0/pre_oi_15_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9591 ), .force_10(
        \filter_0/n9592 ), .force_11(1'b0), .Q(n40467) );
  \**FFGEN**  \filter_0/pre_oi_15_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9595 ), .force_10(
        \filter_0/n9596 ), .force_11(1'b0), .Q(n40372) );
  \**FFGEN**  \filter_0/pre_oi_15_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9599 ), .force_10(
        \filter_0/n9600 ), .force_11(1'b0), .Q(n40403) );
  \**FFGEN**  \filter_0/pre_oi_15_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9603 ), .force_10(
        \filter_0/n9604 ), .force_11(1'b0), .Q(n40338) );
  \**FFGEN**  \filter_0/pre_oi_15_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9607 ), .force_10(
        \filter_0/n9608 ), .force_11(1'b0), .Q(n40371) );
  \**FFGEN**  \filter_0/pre_oi_15_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9611 ), .force_10(
        \filter_0/n9612 ), .force_11(1'b0), .Q(n40304) );
  \**FFGEN**  \filter_0/pre_oi_15_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9615 ), .force_10(
        \filter_0/n9616 ), .force_11(1'b0), .Q(n40337) );
  \**FFGEN**  \filter_0/pre_oi_15_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9619 ), .force_10(
        \filter_0/n9620 ), .force_11(1'b0), .Q(n40271) );
  \**FFGEN**  \filter_0/pre_oi_15_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9623 ), .force_10(
        \filter_0/n9624 ), .force_11(1'b0), .Q(n40303) );
  \**FFGEN**  \filter_0/pre_oi_15_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9627 ), .force_10(
        \filter_0/n9628 ), .force_11(1'b0), .Q(n40246) );
  \**FFGEN**  \filter_0/pre_oi_15_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9631 ), .force_10(
        \filter_0/n9632 ), .force_11(1'b0), .Q(n40270) );
  \**FFGEN**  \filter_0/pre_oi_15_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9635 ), .force_10(
        \filter_0/n9636 ), .force_11(1'b0), .Q(n40233) );
  \**FFGEN**  \filter_0/pre_oi_15_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9639 ), .force_10(
        \filter_0/n9640 ), .force_11(1'b0), .Q(n40245) );
  \**FFGEN**  \filter_0/pre_oi_15_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9643 ), .force_10(
        \filter_0/n9644 ), .force_11(1'b0), .Q(n40231) );
  \**FFGEN**  \filter_0/pre_oi_15_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9647 ), .force_10(
        \filter_0/n9648 ), .force_11(1'b0), .Q(n40230) );
  \**FFGEN**  \filter_0/pre_oi_14_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9651 ), .force_10(
        \filter_0/n9652 ), .force_11(1'b0), .Q(n40603) );
  \**FFGEN**  \filter_0/pre_oi_14_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9655 ), .force_10(
        \filter_0/n9656 ), .force_11(1'b0), .Q(n40602) );
  \**FFGEN**  \filter_0/pre_oi_14_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9659 ), .force_10(
        \filter_0/n9660 ), .force_11(1'b0), .Q(n40601) );
  \**FFGEN**  \filter_0/pre_oi_14_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9663 ), .force_10(
        \filter_0/n9664 ), .force_11(1'b0), .Q(n40600) );
  \**FFGEN**  \filter_0/pre_oi_14_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9667 ), .force_10(
        \filter_0/n9668 ), .force_11(1'b0), .Q(n40599) );
  \**FFGEN**  \filter_0/pre_oi_14_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9671 ), .force_10(
        \filter_0/n9672 ), .force_11(1'b0), .Q(n40598) );
  \**FFGEN**  \filter_0/pre_oi_14_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9675 ), .force_10(
        \filter_0/n9676 ), .force_11(1'b0), .Q(n40597) );
  \**FFGEN**  \filter_0/pre_oi_14_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9679 ), .force_10(
        \filter_0/n9680 ), .force_11(1'b0), .Q(n40596) );
  \**FFGEN**  \filter_0/pre_oi_14_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9683 ), .force_10(
        \filter_0/n9684 ), .force_11(1'b0), .Q(n40498) );
  \**FFGEN**  \filter_0/pre_oi_14_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9687 ), .force_10(
        \filter_0/n9688 ), .force_11(1'b0), .Q(n40466) );
  \**FFGEN**  \filter_0/pre_oi_14_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9691 ), .force_10(
        \filter_0/n9692 ), .force_11(1'b0), .Q(n40435) );
  \**FFGEN**  \filter_0/pre_oi_14_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9695 ), .force_10(
        \filter_0/n9696 ), .force_11(1'b0), .Q(n40402) );
  \**FFGEN**  \filter_0/pre_oi_14_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9699 ), .force_10(
        \filter_0/n9700 ), .force_11(1'b0), .Q(n40370) );
  \**FFGEN**  \filter_0/pre_oi_14_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9703 ), .force_10(
        \filter_0/n9704 ), .force_11(1'b0), .Q(n40595) );
  \**FFGEN**  \filter_0/pre_oi_14_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9707 ), .force_10(
        \filter_0/n9708 ), .force_11(1'b0), .Q(n40336) );
  \**FFGEN**  \filter_0/pre_oi_14_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9711 ), .force_10(
        \filter_0/n9712 ), .force_11(1'b0), .Q(n40302) );
  \**FFGEN**  \filter_0/pre_oi_14_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9715 ), .force_10(
        \filter_0/n9716 ), .force_11(1'b0), .Q(n40594) );
  \**FFGEN**  \filter_0/pre_oi_14_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9719 ), .force_10(
        \filter_0/n9720 ), .force_11(1'b0), .Q(n40593) );
  \**FFGEN**  \filter_0/pre_oi_14_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9723 ), .force_10(
        \filter_0/n9724 ), .force_11(1'b0), .Q(n40269) );
  \**FFGEN**  \filter_0/pre_oi_14_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9727 ), .force_10(
        \filter_0/n9728 ), .force_11(1'b0), .Q(n40244) );
  \**FFGEN**  \filter_0/pre_oi_13_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9731 ), .force_10(
        \filter_0/n9732 ), .force_11(1'b0), .Q(n40614) );
  \**FFGEN**  \filter_0/pre_oi_13_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9735 ), .force_10(
        \filter_0/n9736 ), .force_11(1'b0), .Q(n40613) );
  \**FFGEN**  \filter_0/pre_oi_13_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9739 ), .force_10(
        \filter_0/n9740 ), .force_11(1'b0), .Q(n40612) );
  \**FFGEN**  \filter_0/pre_oi_13_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9743 ), .force_10(
        \filter_0/n9744 ), .force_11(1'b0), .Q(n40611) );
  \**FFGEN**  \filter_0/pre_oi_13_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9747 ), .force_10(
        \filter_0/n9748 ), .force_11(1'b0), .Q(n40610) );
  \**FFGEN**  \filter_0/pre_oi_13_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9751 ), .force_10(
        \filter_0/n9752 ), .force_11(1'b0), .Q(n40609) );
  \**FFGEN**  \filter_0/pre_oi_13_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9755 ), .force_10(
        \filter_0/n9756 ), .force_11(1'b0), .Q(n40608) );
  \**FFGEN**  \filter_0/pre_oi_13_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9759 ), .force_10(
        \filter_0/n9760 ), .force_11(1'b0), .Q(n40607) );
  \**FFGEN**  \filter_0/pre_oi_13_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9763 ), .force_10(
        \filter_0/n9764 ), .force_11(1'b0), .Q(n40497) );
  \**FFGEN**  \filter_0/pre_oi_13_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9767 ), .force_10(
        \filter_0/n9768 ), .force_11(1'b0), .Q(n40465) );
  \**FFGEN**  \filter_0/pre_oi_13_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9771 ), .force_10(
        \filter_0/n9772 ), .force_11(1'b0), .Q(n40434) );
  \**FFGEN**  \filter_0/pre_oi_13_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9775 ), .force_10(
        \filter_0/n9776 ), .force_11(1'b0), .Q(n40606) );
  \**FFGEN**  \filter_0/pre_oi_13_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9779 ), .force_10(
        \filter_0/n9780 ), .force_11(1'b0), .Q(n40401) );
  \**FFGEN**  \filter_0/pre_oi_13_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9783 ), .force_10(
        \filter_0/n9784 ), .force_11(1'b0), .Q(n40605) );
  \**FFGEN**  \filter_0/pre_oi_13_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9787 ), .force_10(
        \filter_0/n9788 ), .force_11(1'b0), .Q(n40369) );
  \**FFGEN**  \filter_0/pre_oi_13_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9791 ), .force_10(
        \filter_0/n9792 ), .force_11(1'b0), .Q(n40335) );
  \**FFGEN**  \filter_0/pre_oi_13_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9795 ), .force_10(
        \filter_0/n9796 ), .force_11(1'b0), .Q(n40604) );
  \**FFGEN**  \filter_0/pre_oi_13_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9799 ), .force_10(
        \filter_0/n9800 ), .force_11(1'b0), .Q(n40301) );
  \**FFGEN**  \filter_0/pre_oi_13_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9803 ), .force_10(
        \filter_0/n9804 ), .force_11(1'b0), .Q(n40268) );
  \**FFGEN**  \filter_0/pre_oi_13_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9807 ), .force_10(
        \filter_0/n9808 ), .force_11(1'b0), .Q(n40243) );
  \**FFGEN**  \filter_0/pre_oi_12_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9811 ), .force_10(
        \filter_0/n9812 ), .force_11(1'b0), .Q(n40625) );
  \**FFGEN**  \filter_0/pre_oi_12_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9815 ), .force_10(
        \filter_0/n9816 ), .force_11(1'b0), .Q(n40624) );
  \**FFGEN**  \filter_0/pre_oi_12_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9819 ), .force_10(
        \filter_0/n9820 ), .force_11(1'b0), .Q(n40623) );
  \**FFGEN**  \filter_0/pre_oi_12_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9823 ), .force_10(
        \filter_0/n9824 ), .force_11(1'b0), .Q(n40622) );
  \**FFGEN**  \filter_0/pre_oi_12_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9827 ), .force_10(
        \filter_0/n9828 ), .force_11(1'b0), .Q(n40621) );
  \**FFGEN**  \filter_0/pre_oi_12_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9831 ), .force_10(
        \filter_0/n9832 ), .force_11(1'b0), .Q(n40620) );
  \**FFGEN**  \filter_0/pre_oi_12_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9835 ), .force_10(
        \filter_0/n9836 ), .force_11(1'b0), .Q(n40619) );
  \**FFGEN**  \filter_0/pre_oi_12_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9839 ), .force_10(
        \filter_0/n9840 ), .force_11(1'b0), .Q(n40618) );
  \**FFGEN**  \filter_0/pre_oi_12_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9843 ), .force_10(
        \filter_0/n9844 ), .force_11(1'b0), .Q(n40496) );
  \**FFGEN**  \filter_0/pre_oi_12_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9847 ), .force_10(
        \filter_0/n9848 ), .force_11(1'b0), .Q(n40464) );
  \**FFGEN**  \filter_0/pre_oi_12_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9851 ), .force_10(
        \filter_0/n9852 ), .force_11(1'b0), .Q(n40433) );
  \**FFGEN**  \filter_0/pre_oi_12_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9855 ), .force_10(
        \filter_0/n9856 ), .force_11(1'b0), .Q(n40400) );
  \**FFGEN**  \filter_0/pre_oi_12_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9859 ), .force_10(
        \filter_0/n9860 ), .force_11(1'b0), .Q(n40368) );
  \**FFGEN**  \filter_0/pre_oi_12_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9863 ), .force_10(
        \filter_0/n9864 ), .force_11(1'b0), .Q(n40617) );
  \**FFGEN**  \filter_0/pre_oi_12_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9867 ), .force_10(
        \filter_0/n9868 ), .force_11(1'b0), .Q(n40334) );
  \**FFGEN**  \filter_0/pre_oi_12_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9871 ), .force_10(
        \filter_0/n9872 ), .force_11(1'b0), .Q(n40300) );
  \**FFGEN**  \filter_0/pre_oi_12_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9875 ), .force_10(
        \filter_0/n9876 ), .force_11(1'b0), .Q(n40616) );
  \**FFGEN**  \filter_0/pre_oi_12_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9879 ), .force_10(
        \filter_0/n9880 ), .force_11(1'b0), .Q(n40615) );
  \**FFGEN**  \filter_0/pre_oi_12_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9883 ), .force_10(
        \filter_0/n9884 ), .force_11(1'b0), .Q(n40267) );
  \**FFGEN**  \filter_0/pre_oi_12_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9887 ), .force_10(
        \filter_0/n9888 ), .force_11(1'b0), .Q(n40242) );
  \**FFGEN**  \filter_0/pre_oi_11_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9891 ), .force_10(
        \filter_0/n9892 ), .force_11(1'b0), .Q(n40637) );
  \**FFGEN**  \filter_0/pre_oi_11_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9895 ), .force_10(
        \filter_0/n9896 ), .force_11(1'b0), .Q(n40636) );
  \**FFGEN**  \filter_0/pre_oi_11_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9899 ), .force_10(
        \filter_0/n9900 ), .force_11(1'b0), .Q(n40635) );
  \**FFGEN**  \filter_0/pre_oi_11_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9903 ), .force_10(
        \filter_0/n9904 ), .force_11(1'b0), .Q(n40634) );
  \**FFGEN**  \filter_0/pre_oi_11_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9907 ), .force_10(
        \filter_0/n9908 ), .force_11(1'b0), .Q(n40633) );
  \**FFGEN**  \filter_0/pre_oi_11_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9911 ), .force_10(
        \filter_0/n9912 ), .force_11(1'b0), .Q(n40632) );
  \**FFGEN**  \filter_0/pre_oi_11_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9915 ), .force_10(
        \filter_0/n9916 ), .force_11(1'b0), .Q(n40495) );
  \**FFGEN**  \filter_0/pre_oi_11_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9919 ), .force_10(
        \filter_0/n9920 ), .force_11(1'b0), .Q(n40463) );
  \**FFGEN**  \filter_0/pre_oi_11_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9923 ), .force_10(
        \filter_0/n9924 ), .force_11(1'b0), .Q(n40631) );
  \**FFGEN**  \filter_0/pre_oi_11_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9927 ), .force_10(
        \filter_0/n9928 ), .force_11(1'b0), .Q(n40432) );
  \**FFGEN**  \filter_0/pre_oi_11_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9931 ), .force_10(
        \filter_0/n9932 ), .force_11(1'b0), .Q(n40630) );
  \**FFGEN**  \filter_0/pre_oi_11_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9935 ), .force_10(
        \filter_0/n9936 ), .force_11(1'b0), .Q(n40399) );
  \**FFGEN**  \filter_0/pre_oi_11_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9939 ), .force_10(
        \filter_0/n9940 ), .force_11(1'b0), .Q(n40629) );
  \**FFGEN**  \filter_0/pre_oi_11_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9943 ), .force_10(
        \filter_0/n9944 ), .force_11(1'b0), .Q(n40367) );
  \**FFGEN**  \filter_0/pre_oi_11_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9947 ), .force_10(
        \filter_0/n9948 ), .force_11(1'b0), .Q(n40628) );
  \**FFGEN**  \filter_0/pre_oi_11_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9951 ), .force_10(
        \filter_0/n9952 ), .force_11(1'b0), .Q(n40333) );
  \**FFGEN**  \filter_0/pre_oi_11_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9955 ), .force_10(
        \filter_0/n9956 ), .force_11(1'b0), .Q(n40627) );
  \**FFGEN**  \filter_0/pre_oi_11_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9959 ), .force_10(
        \filter_0/n9960 ), .force_11(1'b0), .Q(n40299) );
  \**FFGEN**  \filter_0/pre_oi_11_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9963 ), .force_10(
        \filter_0/n9964 ), .force_11(1'b0), .Q(n40626) );
  \**FFGEN**  \filter_0/pre_oi_11_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9967 ), .force_10(
        \filter_0/n9968 ), .force_11(1'b0), .Q(n40266) );
  \**FFGEN**  \filter_0/pre_oi_10_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9971 ), .force_10(
        \filter_0/n9972 ), .force_11(1'b0), .Q(n40649) );
  \**FFGEN**  \filter_0/pre_oi_10_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9975 ), .force_10(
        \filter_0/n9976 ), .force_11(1'b0), .Q(n40648) );
  \**FFGEN**  \filter_0/pre_oi_10_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9979 ), .force_10(
        \filter_0/n9980 ), .force_11(1'b0), .Q(n40647) );
  \**FFGEN**  \filter_0/pre_oi_10_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9983 ), .force_10(
        \filter_0/n9984 ), .force_11(1'b0), .Q(n40646) );
  \**FFGEN**  \filter_0/pre_oi_10_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9987 ), .force_10(
        \filter_0/n9988 ), .force_11(1'b0), .Q(n40645) );
  \**FFGEN**  \filter_0/pre_oi_10_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9991 ), .force_10(
        \filter_0/n9992 ), .force_11(1'b0), .Q(n40644) );
  \**FFGEN**  \filter_0/pre_oi_10_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9995 ), .force_10(
        \filter_0/n9996 ), .force_11(1'b0), .Q(n40643) );
  \**FFGEN**  \filter_0/pre_oi_10_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n9999 ), .force_10(
        \filter_0/n10000 ), .force_11(1'b0), .Q(n40642) );
  \**FFGEN**  \filter_0/pre_oi_10_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10003 ), .force_10(
        \filter_0/n10004 ), .force_11(1'b0), .Q(n40641) );
  \**FFGEN**  \filter_0/pre_oi_10_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10007 ), .force_10(
        \filter_0/n10008 ), .force_11(1'b0), .Q(n40494) );
  \**FFGEN**  \filter_0/pre_oi_10_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10011 ), .force_10(
        \filter_0/n10012 ), .force_11(1'b0), .Q(n40462) );
  \**FFGEN**  \filter_0/pre_oi_10_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10015 ), .force_10(
        \filter_0/n10016 ), .force_11(1'b0), .Q(n40431) );
  \**FFGEN**  \filter_0/pre_oi_10_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10019 ), .force_10(
        \filter_0/n10020 ), .force_11(1'b0), .Q(n40398) );
  \**FFGEN**  \filter_0/pre_oi_10_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10023 ), .force_10(
        \filter_0/n10024 ), .force_11(1'b0), .Q(n40640) );
  \**FFGEN**  \filter_0/pre_oi_10_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10027 ), .force_10(
        \filter_0/n10028 ), .force_11(1'b0), .Q(n40366) );
  \**FFGEN**  \filter_0/pre_oi_10_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10031 ), .force_10(
        \filter_0/n10032 ), .force_11(1'b0), .Q(n40332) );
  \**FFGEN**  \filter_0/pre_oi_10_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10035 ), .force_10(
        \filter_0/n10036 ), .force_11(1'b0), .Q(n40639) );
  \**FFGEN**  \filter_0/pre_oi_10_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10039 ), .force_10(
        \filter_0/n10040 ), .force_11(1'b0), .Q(n40638) );
  \**FFGEN**  \filter_0/pre_oi_10_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10043 ), .force_10(
        \filter_0/n10044 ), .force_11(1'b0), .Q(n40298) );
  \**FFGEN**  \filter_0/pre_oi_10_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10047 ), .force_10(
        \filter_0/n10048 ), .force_11(1'b0), .Q(n40265) );
  \**FFGEN**  \filter_0/pre_oi_9_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10051 ), .force_10(
        \filter_0/n10052 ), .force_11(1'b0), .Q(n40661) );
  \**FFGEN**  \filter_0/pre_oi_9_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10055 ), .force_10(
        \filter_0/n10056 ), .force_11(1'b0), .Q(n40660) );
  \**FFGEN**  \filter_0/pre_oi_9_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10059 ), .force_10(
        \filter_0/n10060 ), .force_11(1'b0), .Q(n40659) );
  \**FFGEN**  \filter_0/pre_oi_9_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10063 ), .force_10(
        \filter_0/n10064 ), .force_11(1'b0), .Q(n40658) );
  \**FFGEN**  \filter_0/pre_oi_9_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10067 ), .force_10(
        \filter_0/n10068 ), .force_11(1'b0), .Q(n40657) );
  \**FFGEN**  \filter_0/pre_oi_9_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10071 ), .force_10(
        \filter_0/n10072 ), .force_11(1'b0), .Q(n40656) );
  \**FFGEN**  \filter_0/pre_oi_9_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10075 ), .force_10(
        \filter_0/n10076 ), .force_11(1'b0), .Q(n40655) );
  \**FFGEN**  \filter_0/pre_oi_9_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10079 ), .force_10(
        \filter_0/n10080 ), .force_11(1'b0), .Q(n40654) );
  \**FFGEN**  \filter_0/pre_oi_9_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10083 ), .force_10(
        \filter_0/n10084 ), .force_11(1'b0), .Q(n40653) );
  \**FFGEN**  \filter_0/pre_oi_9_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10087 ), .force_10(
        \filter_0/n10088 ), .force_11(1'b0), .Q(n40493) );
  \**FFGEN**  \filter_0/pre_oi_9_reg[9]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10091 ), .force_10(\filter_0/n10092 ), 
        .force_11(1'b0), .Q(n40461) );
  \**FFGEN**  \filter_0/pre_oi_9_reg[8]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10095 ), .force_10(\filter_0/n10096 ), 
        .force_11(1'b0), .Q(n40430) );
  \**FFGEN**  \filter_0/pre_oi_9_reg[7]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10099 ), .force_10(\filter_0/n10100 ), 
        .force_11(1'b0), .Q(n40397) );
  \**FFGEN**  \filter_0/pre_oi_9_reg[6]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10103 ), .force_10(\filter_0/n10104 ), 
        .force_11(1'b0), .Q(n40652) );
  \**FFGEN**  \filter_0/pre_oi_9_reg[5]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10107 ), .force_10(\filter_0/n10108 ), 
        .force_11(1'b0), .Q(n40365) );
  \**FFGEN**  \filter_0/pre_oi_9_reg[4]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10111 ), .force_10(\filter_0/n10112 ), 
        .force_11(1'b0), .Q(n40331) );
  \**FFGEN**  \filter_0/pre_oi_9_reg[3]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10115 ), .force_10(\filter_0/n10116 ), 
        .force_11(1'b0), .Q(n40651) );
  \**FFGEN**  \filter_0/pre_oi_9_reg[2]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10119 ), .force_10(\filter_0/n10120 ), 
        .force_11(1'b0), .Q(n40650) );
  \**FFGEN**  \filter_0/pre_oi_9_reg[1]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10123 ), .force_10(\filter_0/n10124 ), 
        .force_11(1'b0), .Q(n40297) );
  \**FFGEN**  \filter_0/pre_oi_9_reg[0]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10127 ), .force_10(\filter_0/n10128 ), 
        .force_11(1'b0), .Q(n40264) );
  \**FFGEN**  \filter_0/pre_oi_8_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10131 ), .force_10(
        \filter_0/n10132 ), .force_11(1'b0), .Q(n40673) );
  \**FFGEN**  \filter_0/pre_oi_8_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10135 ), .force_10(
        \filter_0/n10136 ), .force_11(1'b0), .Q(n40672) );
  \**FFGEN**  \filter_0/pre_oi_8_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10139 ), .force_10(
        \filter_0/n10140 ), .force_11(1'b0), .Q(n40671) );
  \**FFGEN**  \filter_0/pre_oi_8_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10143 ), .force_10(
        \filter_0/n10144 ), .force_11(1'b0), .Q(n40670) );
  \**FFGEN**  \filter_0/pre_oi_8_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10147 ), .force_10(
        \filter_0/n10148 ), .force_11(1'b0), .Q(n40669) );
  \**FFGEN**  \filter_0/pre_oi_8_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10151 ), .force_10(
        \filter_0/n10152 ), .force_11(1'b0), .Q(n40668) );
  \**FFGEN**  \filter_0/pre_oi_8_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10155 ), .force_10(
        \filter_0/n10156 ), .force_11(1'b0), .Q(n40667) );
  \**FFGEN**  \filter_0/pre_oi_8_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10159 ), .force_10(
        \filter_0/n10160 ), .force_11(1'b0), .Q(n40666) );
  \**FFGEN**  \filter_0/pre_oi_8_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10163 ), .force_10(
        \filter_0/n10164 ), .force_11(1'b0), .Q(n40665) );
  \**FFGEN**  \filter_0/pre_oi_8_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10167 ), .force_10(
        \filter_0/n10168 ), .force_11(1'b0), .Q(n40492) );
  \**FFGEN**  \filter_0/pre_oi_8_reg[9]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10171 ), .force_10(\filter_0/n10172 ), 
        .force_11(1'b0), .Q(n40460) );
  \**FFGEN**  \filter_0/pre_oi_8_reg[8]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10175 ), .force_10(\filter_0/n10176 ), 
        .force_11(1'b0), .Q(n40664) );
  \**FFGEN**  \filter_0/pre_oi_8_reg[7]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10179 ), .force_10(\filter_0/n10180 ), 
        .force_11(1'b0), .Q(n40429) );
  \**FFGEN**  \filter_0/pre_oi_8_reg[6]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10183 ), .force_10(\filter_0/n10184 ), 
        .force_11(1'b0), .Q(n40663) );
  \**FFGEN**  \filter_0/pre_oi_8_reg[5]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10187 ), .force_10(\filter_0/n10188 ), 
        .force_11(1'b0), .Q(n40396) );
  \**FFGEN**  \filter_0/pre_oi_8_reg[4]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10191 ), .force_10(\filter_0/n10192 ), 
        .force_11(1'b0), .Q(n40364) );
  \**FFGEN**  \filter_0/pre_oi_8_reg[3]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10195 ), .force_10(\filter_0/n10196 ), 
        .force_11(1'b0), .Q(n40662) );
  \**FFGEN**  \filter_0/pre_oi_8_reg[2]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10199 ), .force_10(\filter_0/n10200 ), 
        .force_11(1'b0), .Q(n40330) );
  \**FFGEN**  \filter_0/pre_oi_8_reg[1]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10203 ), .force_10(\filter_0/n10204 ), 
        .force_11(1'b0), .Q(n40296) );
  \**FFGEN**  \filter_0/pre_oi_8_reg[0]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10207 ), .force_10(\filter_0/n10208 ), 
        .force_11(1'b0), .Q(n40241) );
  \**FFGEN**  \filter_0/pre_oi_7_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10211 ), .force_10(
        \filter_0/n10212 ), .force_11(1'b0), .Q(n40589) );
  \**FFGEN**  \filter_0/pre_oi_7_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10215 ), .force_10(
        \filter_0/n10216 ), .force_11(1'b0), .Q(n40588) );
  \**FFGEN**  \filter_0/pre_oi_7_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10219 ), .force_10(
        \filter_0/n10220 ), .force_11(1'b0), .Q(n40587) );
  \**FFGEN**  \filter_0/pre_oi_7_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10223 ), .force_10(
        \filter_0/n10224 ), .force_11(1'b0), .Q(n40500) );
  \**FFGEN**  \filter_0/pre_oi_7_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10227 ), .force_10(
        \filter_0/n10228 ), .force_11(1'b0), .Q(n40586) );
  \**FFGEN**  \filter_0/pre_oi_7_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10231 ), .force_10(
        \filter_0/n10232 ), .force_11(1'b0), .Q(n40585) );
  \**FFGEN**  \filter_0/pre_oi_7_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10235 ), .force_10(
        \filter_0/n10236 ), .force_11(1'b0), .Q(n40468) );
  \**FFGEN**  \filter_0/pre_oi_7_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10239 ), .force_10(
        \filter_0/n10240 ), .force_11(1'b0), .Q(n40436) );
  \**FFGEN**  \filter_0/pre_oi_7_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10243 ), .force_10(
        \filter_0/n10244 ), .force_11(1'b0), .Q(n40584) );
  \**FFGEN**  \filter_0/pre_oi_7_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10247 ), .force_10(
        \filter_0/n10248 ), .force_11(1'b0), .Q(n40405) );
  \**FFGEN**  \filter_0/pre_oi_7_reg[9]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10251 ), .force_10(\filter_0/n10252 ), 
        .force_11(1'b0), .Q(n40583) );
  \**FFGEN**  \filter_0/pre_oi_7_reg[8]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10255 ), .force_10(\filter_0/n10256 ), 
        .force_11(1'b0), .Q(n40373) );
  \**FFGEN**  \filter_0/pre_oi_7_reg[7]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10259 ), .force_10(\filter_0/n10260 ), 
        .force_11(1'b0), .Q(n40582) );
  \**FFGEN**  \filter_0/pre_oi_7_reg[6]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10263 ), .force_10(\filter_0/n10264 ), 
        .force_11(1'b0), .Q(n40339) );
  \**FFGEN**  \filter_0/pre_oi_7_reg[5]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10267 ), .force_10(\filter_0/n10268 ), 
        .force_11(1'b0), .Q(n40581) );
  \**FFGEN**  \filter_0/pre_oi_7_reg[4]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10271 ), .force_10(\filter_0/n10272 ), 
        .force_11(1'b0), .Q(n40305) );
  \**FFGEN**  \filter_0/pre_oi_7_reg[3]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10275 ), .force_10(\filter_0/n10276 ), 
        .force_11(1'b0), .Q(n40580) );
  \**FFGEN**  \filter_0/pre_oi_7_reg[2]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10279 ), .force_10(\filter_0/n10280 ), 
        .force_11(1'b0), .Q(n40272) );
  \**FFGEN**  \filter_0/pre_oi_7_reg[1]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10283 ), .force_10(\filter_0/n10284 ), 
        .force_11(1'b0), .Q(n40579) );
  \**FFGEN**  \filter_0/pre_oi_7_reg[0]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10287 ), .force_10(\filter_0/n10288 ), 
        .force_11(1'b0), .Q(n40247) );
  \**FFGEN**  \filter_0/pre_oi_6_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10291 ), .force_10(
        \filter_0/n10292 ), .force_11(1'b0), .Q(n40578) );
  \**FFGEN**  \filter_0/pre_oi_6_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10295 ), .force_10(
        \filter_0/n10296 ), .force_11(1'b0), .Q(n40577) );
  \**FFGEN**  \filter_0/pre_oi_6_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10299 ), .force_10(
        \filter_0/n10300 ), .force_11(1'b0), .Q(n40576) );
  \**FFGEN**  \filter_0/pre_oi_6_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10303 ), .force_10(
        \filter_0/n10304 ), .force_11(1'b0), .Q(n40575) );
  \**FFGEN**  \filter_0/pre_oi_6_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10307 ), .force_10(
        \filter_0/n10308 ), .force_11(1'b0), .Q(n40574) );
  \**FFGEN**  \filter_0/pre_oi_6_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10311 ), .force_10(
        \filter_0/n10312 ), .force_11(1'b0), .Q(n40573) );
  \**FFGEN**  \filter_0/pre_oi_6_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10315 ), .force_10(
        \filter_0/n10316 ), .force_11(1'b0), .Q(n40572) );
  \**FFGEN**  \filter_0/pre_oi_6_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10319 ), .force_10(
        \filter_0/n10320 ), .force_11(1'b0), .Q(n40571) );
  \**FFGEN**  \filter_0/pre_oi_6_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10323 ), .force_10(
        \filter_0/n10324 ), .force_11(1'b0), .Q(n40570) );
  \**FFGEN**  \filter_0/pre_oi_6_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10327 ), .force_10(
        \filter_0/n10328 ), .force_11(1'b0), .Q(n40501) );
  \**FFGEN**  \filter_0/pre_oi_6_reg[9]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10331 ), .force_10(\filter_0/n10332 ), 
        .force_11(1'b0), .Q(n40469) );
  \**FFGEN**  \filter_0/pre_oi_6_reg[8]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10335 ), .force_10(\filter_0/n10336 ), 
        .force_11(1'b0), .Q(n40569) );
  \**FFGEN**  \filter_0/pre_oi_6_reg[7]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10339 ), .force_10(\filter_0/n10340 ), 
        .force_11(1'b0), .Q(n40437) );
  \**FFGEN**  \filter_0/pre_oi_6_reg[6]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10343 ), .force_10(\filter_0/n10344 ), 
        .force_11(1'b0), .Q(n40568) );
  \**FFGEN**  \filter_0/pre_oi_6_reg[5]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10347 ), .force_10(\filter_0/n10348 ), 
        .force_11(1'b0), .Q(n40406) );
  \**FFGEN**  \filter_0/pre_oi_6_reg[4]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10351 ), .force_10(\filter_0/n10352 ), 
        .force_11(1'b0), .Q(n40374) );
  \**FFGEN**  \filter_0/pre_oi_6_reg[3]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10355 ), .force_10(\filter_0/n10356 ), 
        .force_11(1'b0), .Q(n40567) );
  \**FFGEN**  \filter_0/pre_oi_6_reg[2]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10359 ), .force_10(\filter_0/n10360 ), 
        .force_11(1'b0), .Q(n40340) );
  \**FFGEN**  \filter_0/pre_oi_6_reg[1]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10363 ), .force_10(\filter_0/n10364 ), 
        .force_11(1'b0), .Q(n40306) );
  \**FFGEN**  \filter_0/pre_oi_6_reg[0]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10367 ), .force_10(\filter_0/n10368 ), 
        .force_11(1'b0), .Q(n40273) );
  \**FFGEN**  \filter_0/pre_oi_5_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10371 ), .force_10(
        \filter_0/n10372 ), .force_11(1'b0), .Q(n40566) );
  \**FFGEN**  \filter_0/pre_oi_5_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10375 ), .force_10(
        \filter_0/n10376 ), .force_11(1'b0), .Q(n40565) );
  \**FFGEN**  \filter_0/pre_oi_5_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10379 ), .force_10(
        \filter_0/n10380 ), .force_11(1'b0), .Q(n40564) );
  \**FFGEN**  \filter_0/pre_oi_5_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10383 ), .force_10(
        \filter_0/n10384 ), .force_11(1'b0), .Q(n40563) );
  \**FFGEN**  \filter_0/pre_oi_5_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10387 ), .force_10(
        \filter_0/n10388 ), .force_11(1'b0), .Q(n40562) );
  \**FFGEN**  \filter_0/pre_oi_5_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10391 ), .force_10(
        \filter_0/n10392 ), .force_11(1'b0), .Q(n40561) );
  \**FFGEN**  \filter_0/pre_oi_5_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10395 ), .force_10(
        \filter_0/n10396 ), .force_11(1'b0), .Q(n40560) );
  \**FFGEN**  \filter_0/pre_oi_5_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10399 ), .force_10(
        \filter_0/n10400 ), .force_11(1'b0), .Q(n40559) );
  \**FFGEN**  \filter_0/pre_oi_5_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10403 ), .force_10(
        \filter_0/n10404 ), .force_11(1'b0), .Q(n40558) );
  \**FFGEN**  \filter_0/pre_oi_5_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10407 ), .force_10(
        \filter_0/n10408 ), .force_11(1'b0), .Q(n40502) );
  \**FFGEN**  \filter_0/pre_oi_5_reg[9]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10411 ), .force_10(\filter_0/n10412 ), 
        .force_11(1'b0), .Q(n40470) );
  \**FFGEN**  \filter_0/pre_oi_5_reg[8]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10415 ), .force_10(\filter_0/n10416 ), 
        .force_11(1'b0), .Q(n40438) );
  \**FFGEN**  \filter_0/pre_oi_5_reg[7]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10419 ), .force_10(\filter_0/n10420 ), 
        .force_11(1'b0), .Q(n40407) );
  \**FFGEN**  \filter_0/pre_oi_5_reg[6]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10423 ), .force_10(\filter_0/n10424 ), 
        .force_11(1'b0), .Q(n40557) );
  \**FFGEN**  \filter_0/pre_oi_5_reg[5]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10427 ), .force_10(\filter_0/n10428 ), 
        .force_11(1'b0), .Q(n40375) );
  \**FFGEN**  \filter_0/pre_oi_5_reg[4]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10431 ), .force_10(\filter_0/n10432 ), 
        .force_11(1'b0), .Q(n40341) );
  \**FFGEN**  \filter_0/pre_oi_5_reg[3]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10435 ), .force_10(\filter_0/n10436 ), 
        .force_11(1'b0), .Q(n40556) );
  \**FFGEN**  \filter_0/pre_oi_5_reg[2]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10439 ), .force_10(\filter_0/n10440 ), 
        .force_11(1'b0), .Q(n40555) );
  \**FFGEN**  \filter_0/pre_oi_5_reg[1]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10443 ), .force_10(\filter_0/n10444 ), 
        .force_11(1'b0), .Q(n40307) );
  \**FFGEN**  \filter_0/pre_oi_5_reg[0]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10447 ), .force_10(\filter_0/n10448 ), 
        .force_11(1'b0), .Q(n40274) );
  \**FFGEN**  \filter_0/pre_oi_4_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10451 ), .force_10(
        \filter_0/n10452 ), .force_11(1'b0), .Q(n40554) );
  \**FFGEN**  \filter_0/pre_oi_4_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10455 ), .force_10(
        \filter_0/n10456 ), .force_11(1'b0), .Q(n40553) );
  \**FFGEN**  \filter_0/pre_oi_4_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10459 ), .force_10(
        \filter_0/n10460 ), .force_11(1'b0), .Q(n40552) );
  \**FFGEN**  \filter_0/pre_oi_4_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10463 ), .force_10(
        \filter_0/n10464 ), .force_11(1'b0), .Q(n40551) );
  \**FFGEN**  \filter_0/pre_oi_4_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10467 ), .force_10(
        \filter_0/n10468 ), .force_11(1'b0), .Q(n40550) );
  \**FFGEN**  \filter_0/pre_oi_4_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10471 ), .force_10(
        \filter_0/n10472 ), .force_11(1'b0), .Q(n40549) );
  \**FFGEN**  \filter_0/pre_oi_4_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10475 ), .force_10(
        \filter_0/n10476 ), .force_11(1'b0), .Q(n40548) );
  \**FFGEN**  \filter_0/pre_oi_4_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10479 ), .force_10(
        \filter_0/n10480 ), .force_11(1'b0), .Q(n40547) );
  \**FFGEN**  \filter_0/pre_oi_4_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10483 ), .force_10(
        \filter_0/n10484 ), .force_11(1'b0), .Q(n40546) );
  \**FFGEN**  \filter_0/pre_oi_4_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10487 ), .force_10(
        \filter_0/n10488 ), .force_11(1'b0), .Q(n40503) );
  \**FFGEN**  \filter_0/pre_oi_4_reg[9]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10491 ), .force_10(\filter_0/n10492 ), 
        .force_11(1'b0), .Q(n40471) );
  \**FFGEN**  \filter_0/pre_oi_4_reg[8]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10495 ), .force_10(\filter_0/n10496 ), 
        .force_11(1'b0), .Q(n40439) );
  \**FFGEN**  \filter_0/pre_oi_4_reg[7]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10499 ), .force_10(\filter_0/n10500 ), 
        .force_11(1'b0), .Q(n40408) );
  \**FFGEN**  \filter_0/pre_oi_4_reg[6]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10503 ), .force_10(\filter_0/n10504 ), 
        .force_11(1'b0), .Q(n40545) );
  \**FFGEN**  \filter_0/pre_oi_4_reg[5]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10507 ), .force_10(\filter_0/n10508 ), 
        .force_11(1'b0), .Q(n40376) );
  \**FFGEN**  \filter_0/pre_oi_4_reg[4]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10511 ), .force_10(\filter_0/n10512 ), 
        .force_11(1'b0), .Q(n40342) );
  \**FFGEN**  \filter_0/pre_oi_4_reg[3]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10515 ), .force_10(\filter_0/n10516 ), 
        .force_11(1'b0), .Q(n40544) );
  \**FFGEN**  \filter_0/pre_oi_4_reg[2]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10519 ), .force_10(\filter_0/n10520 ), 
        .force_11(1'b0), .Q(n40543) );
  \**FFGEN**  \filter_0/pre_oi_4_reg[1]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10523 ), .force_10(\filter_0/n10524 ), 
        .force_11(1'b0), .Q(n40308) );
  \**FFGEN**  \filter_0/pre_oi_4_reg[0]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10527 ), .force_10(\filter_0/n10528 ), 
        .force_11(1'b0), .Q(n40248) );
  \**FFGEN**  \filter_0/pre_oi_3_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10531 ), .force_10(
        \filter_0/n10532 ), .force_11(1'b0), .Q(n40542) );
  \**FFGEN**  \filter_0/pre_oi_3_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10535 ), .force_10(
        \filter_0/n10536 ), .force_11(1'b0), .Q(n40541) );
  \**FFGEN**  \filter_0/pre_oi_3_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10539 ), .force_10(
        \filter_0/n10540 ), .force_11(1'b0), .Q(n40540) );
  \**FFGEN**  \filter_0/pre_oi_3_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10543 ), .force_10(
        \filter_0/n10544 ), .force_11(1'b0), .Q(n40539) );
  \**FFGEN**  \filter_0/pre_oi_3_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10547 ), .force_10(
        \filter_0/n10548 ), .force_11(1'b0), .Q(n40538) );
  \**FFGEN**  \filter_0/pre_oi_3_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10551 ), .force_10(
        \filter_0/n10552 ), .force_11(1'b0), .Q(n40537) );
  \**FFGEN**  \filter_0/pre_oi_3_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10555 ), .force_10(
        \filter_0/n10556 ), .force_11(1'b0), .Q(n40536) );
  \**FFGEN**  \filter_0/pre_oi_3_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10559 ), .force_10(
        \filter_0/n10560 ), .force_11(1'b0), .Q(n40535) );
  \**FFGEN**  \filter_0/pre_oi_3_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10563 ), .force_10(
        \filter_0/n10564 ), .force_11(1'b0), .Q(n40534) );
  \**FFGEN**  \filter_0/pre_oi_3_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10567 ), .force_10(
        \filter_0/n10568 ), .force_11(1'b0), .Q(n40504) );
  \**FFGEN**  \filter_0/pre_oi_3_reg[9]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10571 ), .force_10(\filter_0/n10572 ), 
        .force_11(1'b0), .Q(n40472) );
  \**FFGEN**  \filter_0/pre_oi_3_reg[8]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10575 ), .force_10(\filter_0/n10576 ), 
        .force_11(1'b0), .Q(n40440) );
  \**FFGEN**  \filter_0/pre_oi_3_reg[7]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10579 ), .force_10(\filter_0/n10580 ), 
        .force_11(1'b0), .Q(n40409) );
  \**FFGEN**  \filter_0/pre_oi_3_reg[6]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10583 ), .force_10(\filter_0/n10584 ), 
        .force_11(1'b0), .Q(n40377) );
  \**FFGEN**  \filter_0/pre_oi_3_reg[5]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10587 ), .force_10(\filter_0/n10588 ), 
        .force_11(1'b0), .Q(n40533) );
  \**FFGEN**  \filter_0/pre_oi_3_reg[4]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10591 ), .force_10(\filter_0/n10592 ), 
        .force_11(1'b0), .Q(n40343) );
  \**FFGEN**  \filter_0/pre_oi_3_reg[3]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10595 ), .force_10(\filter_0/n10596 ), 
        .force_11(1'b0), .Q(n40532) );
  \**FFGEN**  \filter_0/pre_oi_3_reg[2]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10599 ), .force_10(\filter_0/n10600 ), 
        .force_11(1'b0), .Q(n40309) );
  \**FFGEN**  \filter_0/pre_oi_3_reg[1]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10603 ), .force_10(\filter_0/n10604 ), 
        .force_11(1'b0), .Q(n40531) );
  \**FFGEN**  \filter_0/pre_oi_3_reg[0]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10607 ), .force_10(\filter_0/n10608 ), 
        .force_11(1'b0), .Q(n40275) );
  \**FFGEN**  \filter_0/pre_oi_2_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10611 ), .force_10(
        \filter_0/n10612 ), .force_11(1'b0), .Q(n40530) );
  \**FFGEN**  \filter_0/pre_oi_2_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10615 ), .force_10(
        \filter_0/n10616 ), .force_11(1'b0), .Q(n40529) );
  \**FFGEN**  \filter_0/pre_oi_2_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10619 ), .force_10(
        \filter_0/n10620 ), .force_11(1'b0), .Q(n40528) );
  \**FFGEN**  \filter_0/pre_oi_2_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10623 ), .force_10(
        \filter_0/n10624 ), .force_11(1'b0), .Q(n40527) );
  \**FFGEN**  \filter_0/pre_oi_2_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10627 ), .force_10(
        \filter_0/n10628 ), .force_11(1'b0), .Q(n40526) );
  \**FFGEN**  \filter_0/pre_oi_2_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10631 ), .force_10(
        \filter_0/n10632 ), .force_11(1'b0), .Q(n40525) );
  \**FFGEN**  \filter_0/pre_oi_2_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10635 ), .force_10(
        \filter_0/n10636 ), .force_11(1'b0), .Q(n40524) );
  \**FFGEN**  \filter_0/pre_oi_2_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10639 ), .force_10(
        \filter_0/n10640 ), .force_11(1'b0), .Q(n40523) );
  \**FFGEN**  \filter_0/pre_oi_2_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10643 ), .force_10(
        \filter_0/n10644 ), .force_11(1'b0), .Q(n40522) );
  \**FFGEN**  \filter_0/pre_oi_2_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10647 ), .force_10(
        \filter_0/n10648 ), .force_11(1'b0), .Q(n40505) );
  \**FFGEN**  \filter_0/pre_oi_2_reg[9]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10651 ), .force_10(\filter_0/n10652 ), 
        .force_11(1'b0), .Q(n40473) );
  \**FFGEN**  \filter_0/pre_oi_2_reg[8]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10655 ), .force_10(\filter_0/n10656 ), 
        .force_11(1'b0), .Q(n40441) );
  \**FFGEN**  \filter_0/pre_oi_2_reg[7]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10659 ), .force_10(\filter_0/n10660 ), 
        .force_11(1'b0), .Q(n40410) );
  \**FFGEN**  \filter_0/pre_oi_2_reg[6]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10663 ), .force_10(\filter_0/n10664 ), 
        .force_11(1'b0), .Q(n40521) );
  \**FFGEN**  \filter_0/pre_oi_2_reg[5]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10667 ), .force_10(\filter_0/n10668 ), 
        .force_11(1'b0), .Q(n40378) );
  \**FFGEN**  \filter_0/pre_oi_2_reg[4]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10671 ), .force_10(\filter_0/n10672 ), 
        .force_11(1'b0), .Q(n40344) );
  \**FFGEN**  \filter_0/pre_oi_2_reg[3]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10675 ), .force_10(\filter_0/n10676 ), 
        .force_11(1'b0), .Q(n40520) );
  \**FFGEN**  \filter_0/pre_oi_2_reg[2]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10679 ), .force_10(\filter_0/n10680 ), 
        .force_11(1'b0), .Q(n40519) );
  \**FFGEN**  \filter_0/pre_oi_2_reg[1]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10683 ), .force_10(\filter_0/n10684 ), 
        .force_11(1'b0), .Q(n40310) );
  \**FFGEN**  \filter_0/pre_oi_2_reg[0]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10687 ), .force_10(\filter_0/n10688 ), 
        .force_11(1'b0), .Q(n40276) );
  \**FFGEN**  \filter_0/pre_oi_1_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10691 ), .force_10(
        \filter_0/n10692 ), .force_11(1'b0), .Q(n40518) );
  \**FFGEN**  \filter_0/pre_oi_1_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10695 ), .force_10(
        \filter_0/n10696 ), .force_11(1'b0), .Q(n40517) );
  \**FFGEN**  \filter_0/pre_oi_1_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10699 ), .force_10(
        \filter_0/n10700 ), .force_11(1'b0), .Q(n40516) );
  \**FFGEN**  \filter_0/pre_oi_1_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10703 ), .force_10(
        \filter_0/n10704 ), .force_11(1'b0), .Q(n40515) );
  \**FFGEN**  \filter_0/pre_oi_1_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10707 ), .force_10(
        \filter_0/n10708 ), .force_11(1'b0), .Q(n40514) );
  \**FFGEN**  \filter_0/pre_oi_1_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10711 ), .force_10(
        \filter_0/n10712 ), .force_11(1'b0), .Q(n40513) );
  \**FFGEN**  \filter_0/pre_oi_1_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10715 ), .force_10(
        \filter_0/n10716 ), .force_11(1'b0), .Q(n40512) );
  \**FFGEN**  \filter_0/pre_oi_1_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10719 ), .force_10(
        \filter_0/n10720 ), .force_11(1'b0), .Q(n40511) );
  \**FFGEN**  \filter_0/pre_oi_1_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10723 ), .force_10(
        \filter_0/n10724 ), .force_11(1'b0), .Q(n40510) );
  \**FFGEN**  \filter_0/pre_oi_1_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10727 ), .force_10(
        \filter_0/n10728 ), .force_11(1'b0), .Q(n40506) );
  \**FFGEN**  \filter_0/pre_oi_1_reg[9]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10731 ), .force_10(\filter_0/n10732 ), 
        .force_11(1'b0), .Q(n40474) );
  \**FFGEN**  \filter_0/pre_oi_1_reg[8]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10735 ), .force_10(\filter_0/n10736 ), 
        .force_11(1'b0), .Q(n40442) );
  \**FFGEN**  \filter_0/pre_oi_1_reg[7]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10739 ), .force_10(\filter_0/n10740 ), 
        .force_11(1'b0), .Q(n40411) );
  \**FFGEN**  \filter_0/pre_oi_1_reg[6]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10743 ), .force_10(\filter_0/n10744 ), 
        .force_11(1'b0), .Q(n40509) );
  \**FFGEN**  \filter_0/pre_oi_1_reg[5]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10747 ), .force_10(\filter_0/n10748 ), 
        .force_11(1'b0), .Q(n40379) );
  \**FFGEN**  \filter_0/pre_oi_1_reg[4]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10751 ), .force_10(\filter_0/n10752 ), 
        .force_11(1'b0), .Q(n40345) );
  \**FFGEN**  \filter_0/pre_oi_1_reg[3]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10755 ), .force_10(\filter_0/n10756 ), 
        .force_11(1'b0), .Q(n40508) );
  \**FFGEN**  \filter_0/pre_oi_1_reg[2]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10759 ), .force_10(\filter_0/n10760 ), 
        .force_11(1'b0), .Q(n40507) );
  \**FFGEN**  \filter_0/pre_oi_1_reg[1]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10763 ), .force_10(\filter_0/n10764 ), 
        .force_11(1'b0), .Q(n40311) );
  \**FFGEN**  \filter_0/pre_oi_1_reg[0]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10767 ), .force_10(\filter_0/n10768 ), 
        .force_11(1'b0), .Q(n40277) );
  \**FFGEN**  \filter_0/pre_oi_0_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10771 ), .force_10(
        \filter_0/n10772 ), .force_11(1'b0), .Q(n40686) );
  \**FFGEN**  \filter_0/pre_oi_0_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10775 ), .force_10(
        \filter_0/n10776 ), .force_11(1'b0), .Q(n40685) );
  \**FFGEN**  \filter_0/pre_oi_0_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10779 ), .force_10(
        \filter_0/n10780 ), .force_11(1'b0), .Q(n40684) );
  \**FFGEN**  \filter_0/pre_oi_0_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10783 ), .force_10(
        \filter_0/n10784 ), .force_11(1'b0), .Q(n40683) );
  \**FFGEN**  \filter_0/pre_oi_0_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10787 ), .force_10(
        \filter_0/n10788 ), .force_11(1'b0), .Q(n40682) );
  \**FFGEN**  \filter_0/pre_oi_0_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10791 ), .force_10(
        \filter_0/n10792 ), .force_11(1'b0), .Q(n40681) );
  \**FFGEN**  \filter_0/pre_oi_0_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10795 ), .force_10(
        \filter_0/n10796 ), .force_11(1'b0), .Q(n40680) );
  \**FFGEN**  \filter_0/pre_oi_0_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10799 ), .force_10(
        \filter_0/n10800 ), .force_11(1'b0), .Q(n40679) );
  \**FFGEN**  \filter_0/pre_oi_0_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10803 ), .force_10(
        \filter_0/n10804 ), .force_11(1'b0), .Q(n40678) );
  \**FFGEN**  \filter_0/pre_oi_0_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\filter_0/n10807 ), .force_10(
        \filter_0/n10808 ), .force_11(1'b0), .Q(n40677) );
  \**FFGEN**  \filter_0/pre_oi_0_reg[9]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10811 ), .force_10(\filter_0/n10812 ), 
        .force_11(1'b0), .Q(n40491) );
  \**FFGEN**  \filter_0/pre_oi_0_reg[8]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10815 ), .force_10(\filter_0/n10816 ), 
        .force_11(1'b0), .Q(n40676) );
  \**FFGEN**  \filter_0/pre_oi_0_reg[7]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10819 ), .force_10(\filter_0/n10820 ), 
        .force_11(1'b0), .Q(n40459) );
  \**FFGEN**  \filter_0/pre_oi_0_reg[6]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10823 ), .force_10(\filter_0/n10824 ), 
        .force_11(1'b0), .Q(n40675) );
  \**FFGEN**  \filter_0/pre_oi_0_reg[5]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10827 ), .force_10(\filter_0/n10828 ), 
        .force_11(1'b0), .Q(n40428) );
  \**FFGEN**  \filter_0/pre_oi_0_reg[4]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10831 ), .force_10(\filter_0/n10832 ), 
        .force_11(1'b0), .Q(n40395) );
  \**FFGEN**  \filter_0/pre_oi_0_reg[3]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10835 ), .force_10(\filter_0/n10836 ), 
        .force_11(1'b0), .Q(n40674) );
  \**FFGEN**  \filter_0/pre_oi_0_reg[2]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10839 ), .force_10(\filter_0/n10840 ), 
        .force_11(1'b0), .Q(n40363) );
  \**FFGEN**  \filter_0/pre_oi_0_reg[1]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n10843 ), .force_10(\filter_0/n10844 ), 
        .force_11(1'b0), .Q(n40329) );
  \**FFGEN**  \filter_0/pre_oi_0_reg[0]  ( .next_state(1'b0), .clocked_on(1'b0), .force_00(1'b0), .force_01(\filter_0/n8235 ), .force_10(\filter_0/n8236 ), 
        .force_11(1'b0), .Q(n40295) );
  \**FFGEN**  \shifter_0/pre_ow_15_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10208 ), .force_10(
        \shifter_0/n10209 ), .force_11(1'b0), .QN(n46214) );
  \**FFGEN**  \shifter_0/pre_ow_15_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10212 ), .force_10(
        \shifter_0/n10213 ), .force_11(1'b0), .QN(n46215) );
  \**FFGEN**  \shifter_0/pre_ow_15_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10216 ), .force_10(
        \shifter_0/n10217 ), .force_11(1'b0), .QN(n46216) );
  \**FFGEN**  \shifter_0/pre_ow_15_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10220 ), .force_10(
        \shifter_0/n10221 ), .force_11(1'b0), .QN(n46217) );
  \**FFGEN**  \shifter_0/pre_ow_15_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10224 ), .force_10(
        \shifter_0/n10225 ), .force_11(1'b0), .QN(n46218) );
  \**FFGEN**  \shifter_0/pre_ow_15_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10228 ), .force_10(
        \shifter_0/n10229 ), .force_11(1'b0), .QN(n46219) );
  \**FFGEN**  \shifter_0/pre_ow_15_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10232 ), .force_10(
        \shifter_0/n10233 ), .force_11(1'b0), .QN(n46220) );
  \**FFGEN**  \shifter_0/pre_ow_15_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10236 ), .force_10(
        \shifter_0/n10237 ), .force_11(1'b0), .QN(n46221) );
  \**FFGEN**  \shifter_0/pre_ow_15_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10240 ), .force_10(
        \shifter_0/n10241 ), .force_11(1'b0), .QN(n46222) );
  \**FFGEN**  \shifter_0/pre_ow_15_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10244 ), .force_10(
        \shifter_0/n10245 ), .force_11(1'b0), .QN(n46223) );
  \**FFGEN**  \shifter_0/pre_ow_15_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10248 ), .force_10(
        \shifter_0/n10249 ), .force_11(1'b0), .QN(n46224) );
  \**FFGEN**  \shifter_0/pre_ow_15_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10252 ), .force_10(
        \shifter_0/n10253 ), .force_11(1'b0), .QN(n46225) );
  \**FFGEN**  \shifter_0/pre_ow_15_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10256 ), .force_10(
        \shifter_0/n10257 ), .force_11(1'b0), .QN(n46226) );
  \**FFGEN**  \shifter_0/pre_ow_15_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10260 ), .force_10(
        \shifter_0/n10261 ), .force_11(1'b0), .QN(n46227) );
  \**FFGEN**  \shifter_0/pre_ow_15_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10264 ), .force_10(
        \shifter_0/n10265 ), .force_11(1'b0), .QN(n46228) );
  \**FFGEN**  \shifter_0/pre_ow_15_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10268 ), .force_10(
        \shifter_0/n10269 ), .force_11(1'b0), .QN(n46229) );
  \**FFGEN**  \shifter_0/pre_ow_15_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10272 ), .force_10(
        \shifter_0/n10273 ), .force_11(1'b0), .QN(n46230) );
  \**FFGEN**  \shifter_0/pre_ow_15_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10276 ), .force_10(
        \shifter_0/n10277 ), .force_11(1'b0), .QN(n46231) );
  \**FFGEN**  \shifter_0/pre_ow_15_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10280 ), .force_10(
        \shifter_0/n10281 ), .force_11(1'b0), .QN(n46232) );
  \**FFGEN**  \shifter_0/pre_ow_15_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10284 ), .force_10(
        \shifter_0/n10285 ), .force_11(1'b0), .QN(n46853) );
  \**FFGEN**  \shifter_0/pre_oi_0_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10288 ), .force_10(
        \shifter_0/n10289 ), .force_11(1'b0), .QN(n46233) );
  \**FFGEN**  \shifter_0/pre_oi_0_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10292 ), .force_10(
        \shifter_0/n10293 ), .force_11(1'b0), .QN(n46234) );
  \**FFGEN**  \shifter_0/pre_oi_0_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10296 ), .force_10(
        \shifter_0/n10297 ), .force_11(1'b0), .QN(n46235) );
  \**FFGEN**  \shifter_0/pre_oi_0_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10300 ), .force_10(
        \shifter_0/n10301 ), .force_11(1'b0), .QN(n46236) );
  \**FFGEN**  \shifter_0/pre_oi_0_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10304 ), .force_10(
        \shifter_0/n10305 ), .force_11(1'b0), .QN(n46237) );
  \**FFGEN**  \shifter_0/pre_oi_0_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10308 ), .force_10(
        \shifter_0/n10309 ), .force_11(1'b0), .QN(n46238) );
  \**FFGEN**  \shifter_0/pre_oi_0_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10312 ), .force_10(
        \shifter_0/n10313 ), .force_11(1'b0), .QN(n46239) );
  \**FFGEN**  \shifter_0/pre_oi_0_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10316 ), .force_10(
        \shifter_0/n10317 ), .force_11(1'b0), .QN(n46240) );
  \**FFGEN**  \shifter_0/pre_oi_0_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10320 ), .force_10(
        \shifter_0/n10321 ), .force_11(1'b0), .QN(n46241) );
  \**FFGEN**  \shifter_0/pre_oi_0_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10324 ), .force_10(
        \shifter_0/n10325 ), .force_11(1'b0), .QN(n46242) );
  \**FFGEN**  \shifter_0/pre_oi_0_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10328 ), .force_10(
        \shifter_0/n10329 ), .force_11(1'b0), .QN(n46243) );
  \**FFGEN**  \shifter_0/pre_oi_0_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10332 ), .force_10(
        \shifter_0/n10333 ), .force_11(1'b0), .QN(n46244) );
  \**FFGEN**  \shifter_0/pre_oi_0_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10336 ), .force_10(
        \shifter_0/n10337 ), .force_11(1'b0), .QN(n46245) );
  \**FFGEN**  \shifter_0/pre_oi_0_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10340 ), .force_10(
        \shifter_0/n10341 ), .force_11(1'b0), .QN(n46246) );
  \**FFGEN**  \shifter_0/pre_oi_0_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10344 ), .force_10(
        \shifter_0/n10345 ), .force_11(1'b0), .QN(n46247) );
  \**FFGEN**  \shifter_0/pre_oi_0_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10348 ), .force_10(
        \shifter_0/n10349 ), .force_11(1'b0), .QN(n46248) );
  \**FFGEN**  \shifter_0/pre_oi_0_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10352 ), .force_10(
        \shifter_0/n10353 ), .force_11(1'b0), .QN(n46249) );
  \**FFGEN**  \shifter_0/pre_oi_0_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10356 ), .force_10(
        \shifter_0/n10357 ), .force_11(1'b0), .QN(n46250) );
  \**FFGEN**  \shifter_0/pre_oi_0_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10360 ), .force_10(
        \shifter_0/n10361 ), .force_11(1'b0), .QN(n46251) );
  \**FFGEN**  \shifter_0/pre_oi_0_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10364 ), .force_10(
        \shifter_0/n10365 ), .force_11(1'b0), .QN(n46252) );
  \**FFGEN**  \shifter_0/pre_ow_0_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10368 ), .force_10(
        \shifter_0/n10369 ), .force_11(1'b0), .QN(n46553) );
  \**FFGEN**  \shifter_0/pre_ow_0_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10372 ), .force_10(
        \shifter_0/n10373 ), .force_11(1'b0), .QN(n46554) );
  \**FFGEN**  \shifter_0/pre_ow_0_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10376 ), .force_10(
        \shifter_0/n10377 ), .force_11(1'b0), .QN(n46555) );
  \**FFGEN**  \shifter_0/pre_ow_0_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10380 ), .force_10(
        \shifter_0/n10381 ), .force_11(1'b0), .QN(n46556) );
  \**FFGEN**  \shifter_0/pre_ow_0_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10384 ), .force_10(
        \shifter_0/n10385 ), .force_11(1'b0), .QN(n46557) );
  \**FFGEN**  \shifter_0/pre_ow_0_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10388 ), .force_10(
        \shifter_0/n10389 ), .force_11(1'b0), .QN(n46558) );
  \**FFGEN**  \shifter_0/pre_ow_0_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10392 ), .force_10(
        \shifter_0/n10393 ), .force_11(1'b0), .QN(n46559) );
  \**FFGEN**  \shifter_0/pre_ow_0_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10396 ), .force_10(
        \shifter_0/n10397 ), .force_11(1'b0), .QN(n46560) );
  \**FFGEN**  \shifter_0/pre_ow_0_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10400 ), .force_10(
        \shifter_0/n10401 ), .force_11(1'b0), .QN(n46561) );
  \**FFGEN**  \shifter_0/pre_ow_0_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10404 ), .force_10(
        \shifter_0/n10405 ), .force_11(1'b0), .QN(n46562) );
  \**FFGEN**  \shifter_0/pre_ow_0_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10408 ), .force_10(
        \shifter_0/n10409 ), .force_11(1'b0), .QN(n46563) );
  \**FFGEN**  \shifter_0/pre_ow_0_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10412 ), .force_10(
        \shifter_0/n10413 ), .force_11(1'b0), .QN(n46564) );
  \**FFGEN**  \shifter_0/pre_ow_0_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10416 ), .force_10(
        \shifter_0/n10417 ), .force_11(1'b0), .QN(n46565) );
  \**FFGEN**  \shifter_0/pre_ow_0_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10420 ), .force_10(
        \shifter_0/n10421 ), .force_11(1'b0), .QN(n46566) );
  \**FFGEN**  \shifter_0/pre_ow_0_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10424 ), .force_10(
        \shifter_0/n10425 ), .force_11(1'b0), .QN(n46567) );
  \**FFGEN**  \shifter_0/pre_ow_0_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10428 ), .force_10(
        \shifter_0/n10429 ), .force_11(1'b0), .QN(n46568) );
  \**FFGEN**  \shifter_0/pre_ow_0_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10432 ), .force_10(
        \shifter_0/n10433 ), .force_11(1'b0), .QN(n46569) );
  \**FFGEN**  \shifter_0/pre_ow_0_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10436 ), .force_10(
        \shifter_0/n10437 ), .force_11(1'b0), .QN(n46570) );
  \**FFGEN**  \shifter_0/pre_ow_0_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10440 ), .force_10(
        \shifter_0/n10441 ), .force_11(1'b0), .QN(n46571) );
  \**FFGEN**  \shifter_0/pre_ow_0_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10444 ), .force_10(
        \shifter_0/n10445 ), .force_11(1'b0), .QN(n46572) );
  \**FFGEN**  \shifter_0/pre_oi_1_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10448 ), .force_10(
        \shifter_0/n10449 ), .force_11(1'b0), .QN(n46253) );
  \**FFGEN**  \shifter_0/pre_oi_1_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10452 ), .force_10(
        \shifter_0/n10453 ), .force_11(1'b0), .QN(n46254) );
  \**FFGEN**  \shifter_0/pre_oi_1_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10456 ), .force_10(
        \shifter_0/n10457 ), .force_11(1'b0), .QN(n46255) );
  \**FFGEN**  \shifter_0/pre_oi_1_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10460 ), .force_10(
        \shifter_0/n10461 ), .force_11(1'b0), .QN(n46256) );
  \**FFGEN**  \shifter_0/pre_oi_1_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10464 ), .force_10(
        \shifter_0/n10465 ), .force_11(1'b0), .QN(n46257) );
  \**FFGEN**  \shifter_0/pre_oi_1_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10468 ), .force_10(
        \shifter_0/n10469 ), .force_11(1'b0), .QN(n46258) );
  \**FFGEN**  \shifter_0/pre_oi_1_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10472 ), .force_10(
        \shifter_0/n10473 ), .force_11(1'b0), .QN(n46259) );
  \**FFGEN**  \shifter_0/pre_oi_1_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10476 ), .force_10(
        \shifter_0/n10477 ), .force_11(1'b0), .QN(n46260) );
  \**FFGEN**  \shifter_0/pre_oi_1_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10480 ), .force_10(
        \shifter_0/n10481 ), .force_11(1'b0), .QN(n46261) );
  \**FFGEN**  \shifter_0/pre_oi_1_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10484 ), .force_10(
        \shifter_0/n10485 ), .force_11(1'b0), .QN(n46262) );
  \**FFGEN**  \shifter_0/pre_oi_1_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10488 ), .force_10(
        \shifter_0/n10489 ), .force_11(1'b0), .QN(n46263) );
  \**FFGEN**  \shifter_0/pre_oi_1_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10492 ), .force_10(
        \shifter_0/n10493 ), .force_11(1'b0), .QN(n46264) );
  \**FFGEN**  \shifter_0/pre_oi_1_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10496 ), .force_10(
        \shifter_0/n10497 ), .force_11(1'b0), .QN(n46265) );
  \**FFGEN**  \shifter_0/pre_oi_1_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10500 ), .force_10(
        \shifter_0/n10501 ), .force_11(1'b0), .QN(n46266) );
  \**FFGEN**  \shifter_0/pre_oi_1_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10504 ), .force_10(
        \shifter_0/n10505 ), .force_11(1'b0), .QN(n46267) );
  \**FFGEN**  \shifter_0/pre_oi_1_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10508 ), .force_10(
        \shifter_0/n10509 ), .force_11(1'b0), .QN(n46268) );
  \**FFGEN**  \shifter_0/pre_oi_1_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10512 ), .force_10(
        \shifter_0/n10513 ), .force_11(1'b0), .QN(n46269) );
  \**FFGEN**  \shifter_0/pre_oi_1_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10516 ), .force_10(
        \shifter_0/n10517 ), .force_11(1'b0), .QN(n46270) );
  \**FFGEN**  \shifter_0/pre_oi_1_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10520 ), .force_10(
        \shifter_0/n10521 ), .force_11(1'b0), .QN(n46271) );
  \**FFGEN**  \shifter_0/pre_oi_1_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10524 ), .force_10(
        \shifter_0/n10525 ), .force_11(1'b0), .QN(n46272) );
  \**FFGEN**  \shifter_0/pre_ow_1_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10528 ), .force_10(
        \shifter_0/n10529 ), .force_11(1'b0), .QN(n46573) );
  \**FFGEN**  \shifter_0/pre_ow_1_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10532 ), .force_10(
        \shifter_0/n10533 ), .force_11(1'b0), .QN(n46574) );
  \**FFGEN**  \shifter_0/pre_ow_1_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10536 ), .force_10(
        \shifter_0/n10537 ), .force_11(1'b0), .QN(n46575) );
  \**FFGEN**  \shifter_0/pre_ow_1_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10540 ), .force_10(
        \shifter_0/n10541 ), .force_11(1'b0), .QN(n46576) );
  \**FFGEN**  \shifter_0/pre_ow_1_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10544 ), .force_10(
        \shifter_0/n10545 ), .force_11(1'b0), .QN(n46577) );
  \**FFGEN**  \shifter_0/pre_ow_1_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10548 ), .force_10(
        \shifter_0/n10549 ), .force_11(1'b0), .QN(n46578) );
  \**FFGEN**  \shifter_0/pre_ow_1_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10552 ), .force_10(
        \shifter_0/n10553 ), .force_11(1'b0), .QN(n46579) );
  \**FFGEN**  \shifter_0/pre_ow_1_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10556 ), .force_10(
        \shifter_0/n10557 ), .force_11(1'b0), .QN(n46580) );
  \**FFGEN**  \shifter_0/pre_ow_1_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10560 ), .force_10(
        \shifter_0/n10561 ), .force_11(1'b0), .QN(n46581) );
  \**FFGEN**  \shifter_0/pre_ow_1_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10564 ), .force_10(
        \shifter_0/n10565 ), .force_11(1'b0), .QN(n46582) );
  \**FFGEN**  \shifter_0/pre_ow_1_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10568 ), .force_10(
        \shifter_0/n10569 ), .force_11(1'b0), .QN(n46583) );
  \**FFGEN**  \shifter_0/pre_ow_1_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10572 ), .force_10(
        \shifter_0/n10573 ), .force_11(1'b0), .QN(n46584) );
  \**FFGEN**  \shifter_0/pre_ow_1_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10576 ), .force_10(
        \shifter_0/n10577 ), .force_11(1'b0), .QN(n46585) );
  \**FFGEN**  \shifter_0/pre_ow_1_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10580 ), .force_10(
        \shifter_0/n10581 ), .force_11(1'b0), .QN(n46586) );
  \**FFGEN**  \shifter_0/pre_ow_1_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10584 ), .force_10(
        \shifter_0/n10585 ), .force_11(1'b0), .QN(n46587) );
  \**FFGEN**  \shifter_0/pre_ow_1_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10588 ), .force_10(
        \shifter_0/n10589 ), .force_11(1'b0), .QN(n46588) );
  \**FFGEN**  \shifter_0/pre_ow_1_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10592 ), .force_10(
        \shifter_0/n10593 ), .force_11(1'b0), .QN(n46589) );
  \**FFGEN**  \shifter_0/pre_ow_1_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10596 ), .force_10(
        \shifter_0/n10597 ), .force_11(1'b0), .QN(n46590) );
  \**FFGEN**  \shifter_0/pre_ow_1_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10600 ), .force_10(
        \shifter_0/n10601 ), .force_11(1'b0), .QN(n46591) );
  \**FFGEN**  \shifter_0/pre_ow_1_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10604 ), .force_10(
        \shifter_0/n10605 ), .force_11(1'b0), .QN(n46592) );
  \**FFGEN**  \shifter_0/pre_oi_2_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10608 ), .force_10(
        \shifter_0/n10609 ), .force_11(1'b0), .QN(n46273) );
  \**FFGEN**  \shifter_0/pre_oi_2_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10612 ), .force_10(
        \shifter_0/n10613 ), .force_11(1'b0), .QN(n46274) );
  \**FFGEN**  \shifter_0/pre_oi_2_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10616 ), .force_10(
        \shifter_0/n10617 ), .force_11(1'b0), .QN(n46275) );
  \**FFGEN**  \shifter_0/pre_oi_2_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10620 ), .force_10(
        \shifter_0/n10621 ), .force_11(1'b0), .QN(n46276) );
  \**FFGEN**  \shifter_0/pre_oi_2_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10624 ), .force_10(
        \shifter_0/n10625 ), .force_11(1'b0), .QN(n46277) );
  \**FFGEN**  \shifter_0/pre_oi_2_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10628 ), .force_10(
        \shifter_0/n10629 ), .force_11(1'b0), .QN(n46278) );
  \**FFGEN**  \shifter_0/pre_oi_2_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10632 ), .force_10(
        \shifter_0/n10633 ), .force_11(1'b0), .QN(n46279) );
  \**FFGEN**  \shifter_0/pre_oi_2_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10636 ), .force_10(
        \shifter_0/n10637 ), .force_11(1'b0), .QN(n46280) );
  \**FFGEN**  \shifter_0/pre_oi_2_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10640 ), .force_10(
        \shifter_0/n10641 ), .force_11(1'b0), .QN(n46281) );
  \**FFGEN**  \shifter_0/pre_oi_2_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10644 ), .force_10(
        \shifter_0/n10645 ), .force_11(1'b0), .QN(n46282) );
  \**FFGEN**  \shifter_0/pre_oi_2_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10648 ), .force_10(
        \shifter_0/n10649 ), .force_11(1'b0), .QN(n46283) );
  \**FFGEN**  \shifter_0/pre_oi_2_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10652 ), .force_10(
        \shifter_0/n10653 ), .force_11(1'b0), .QN(n46284) );
  \**FFGEN**  \shifter_0/pre_oi_2_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10656 ), .force_10(
        \shifter_0/n10657 ), .force_11(1'b0), .QN(n46285) );
  \**FFGEN**  \shifter_0/pre_oi_2_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10660 ), .force_10(
        \shifter_0/n10661 ), .force_11(1'b0), .QN(n46286) );
  \**FFGEN**  \shifter_0/pre_oi_2_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10664 ), .force_10(
        \shifter_0/n10665 ), .force_11(1'b0), .QN(n46287) );
  \**FFGEN**  \shifter_0/pre_oi_2_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10668 ), .force_10(
        \shifter_0/n10669 ), .force_11(1'b0), .QN(n46288) );
  \**FFGEN**  \shifter_0/pre_oi_2_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10672 ), .force_10(
        \shifter_0/n10673 ), .force_11(1'b0), .QN(n46289) );
  \**FFGEN**  \shifter_0/pre_oi_2_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10676 ), .force_10(
        \shifter_0/n10677 ), .force_11(1'b0), .QN(n46290) );
  \**FFGEN**  \shifter_0/pre_oi_2_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10680 ), .force_10(
        \shifter_0/n10681 ), .force_11(1'b0), .QN(n46291) );
  \**FFGEN**  \shifter_0/pre_oi_2_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10684 ), .force_10(
        \shifter_0/n10685 ), .force_11(1'b0), .QN(n46292) );
  \**FFGEN**  \shifter_0/pre_ow_2_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10688 ), .force_10(
        \shifter_0/n10689 ), .force_11(1'b0), .QN(n46593) );
  \**FFGEN**  \shifter_0/pre_ow_2_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10692 ), .force_10(
        \shifter_0/n10693 ), .force_11(1'b0), .QN(n46594) );
  \**FFGEN**  \shifter_0/pre_ow_2_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10696 ), .force_10(
        \shifter_0/n10697 ), .force_11(1'b0), .QN(n46595) );
  \**FFGEN**  \shifter_0/pre_ow_2_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10700 ), .force_10(
        \shifter_0/n10701 ), .force_11(1'b0), .QN(n46596) );
  \**FFGEN**  \shifter_0/pre_ow_2_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10704 ), .force_10(
        \shifter_0/n10705 ), .force_11(1'b0), .QN(n46597) );
  \**FFGEN**  \shifter_0/pre_ow_2_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10708 ), .force_10(
        \shifter_0/n10709 ), .force_11(1'b0), .QN(n46598) );
  \**FFGEN**  \shifter_0/pre_ow_2_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10712 ), .force_10(
        \shifter_0/n10713 ), .force_11(1'b0), .QN(n46599) );
  \**FFGEN**  \shifter_0/pre_ow_2_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10716 ), .force_10(
        \shifter_0/n10717 ), .force_11(1'b0), .QN(n46600) );
  \**FFGEN**  \shifter_0/pre_ow_2_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10720 ), .force_10(
        \shifter_0/n10721 ), .force_11(1'b0), .QN(n46601) );
  \**FFGEN**  \shifter_0/pre_ow_2_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10724 ), .force_10(
        \shifter_0/n10725 ), .force_11(1'b0), .QN(n46602) );
  \**FFGEN**  \shifter_0/pre_ow_2_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10728 ), .force_10(
        \shifter_0/n10729 ), .force_11(1'b0), .QN(n46603) );
  \**FFGEN**  \shifter_0/pre_ow_2_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10732 ), .force_10(
        \shifter_0/n10733 ), .force_11(1'b0), .QN(n46604) );
  \**FFGEN**  \shifter_0/pre_ow_2_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10736 ), .force_10(
        \shifter_0/n10737 ), .force_11(1'b0), .QN(n46605) );
  \**FFGEN**  \shifter_0/pre_ow_2_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10740 ), .force_10(
        \shifter_0/n10741 ), .force_11(1'b0), .QN(n46606) );
  \**FFGEN**  \shifter_0/pre_ow_2_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10744 ), .force_10(
        \shifter_0/n10745 ), .force_11(1'b0), .QN(n46607) );
  \**FFGEN**  \shifter_0/pre_ow_2_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10748 ), .force_10(
        \shifter_0/n10749 ), .force_11(1'b0), .QN(n46608) );
  \**FFGEN**  \shifter_0/pre_ow_2_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10752 ), .force_10(
        \shifter_0/n10753 ), .force_11(1'b0), .QN(n46609) );
  \**FFGEN**  \shifter_0/pre_ow_2_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10756 ), .force_10(
        \shifter_0/n10757 ), .force_11(1'b0), .QN(n46610) );
  \**FFGEN**  \shifter_0/pre_ow_2_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10760 ), .force_10(
        \shifter_0/n10761 ), .force_11(1'b0), .QN(n46611) );
  \**FFGEN**  \shifter_0/pre_ow_2_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10764 ), .force_10(
        \shifter_0/n10765 ), .force_11(1'b0), .QN(n46612) );
  \**FFGEN**  \shifter_0/pre_oi_3_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10768 ), .force_10(
        \shifter_0/n10769 ), .force_11(1'b0), .QN(n46293) );
  \**FFGEN**  \shifter_0/pre_oi_3_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10772 ), .force_10(
        \shifter_0/n10773 ), .force_11(1'b0), .QN(n46294) );
  \**FFGEN**  \shifter_0/pre_oi_3_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10776 ), .force_10(
        \shifter_0/n10777 ), .force_11(1'b0), .QN(n46295) );
  \**FFGEN**  \shifter_0/pre_oi_3_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10780 ), .force_10(
        \shifter_0/n10781 ), .force_11(1'b0), .QN(n46296) );
  \**FFGEN**  \shifter_0/pre_oi_3_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10784 ), .force_10(
        \shifter_0/n10785 ), .force_11(1'b0), .QN(n46297) );
  \**FFGEN**  \shifter_0/pre_oi_3_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10788 ), .force_10(
        \shifter_0/n10789 ), .force_11(1'b0), .QN(n46298) );
  \**FFGEN**  \shifter_0/pre_oi_3_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10792 ), .force_10(
        \shifter_0/n10793 ), .force_11(1'b0), .QN(n46299) );
  \**FFGEN**  \shifter_0/pre_oi_3_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10796 ), .force_10(
        \shifter_0/n10797 ), .force_11(1'b0), .QN(n46300) );
  \**FFGEN**  \shifter_0/pre_oi_3_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10800 ), .force_10(
        \shifter_0/n10801 ), .force_11(1'b0), .QN(n46301) );
  \**FFGEN**  \shifter_0/pre_oi_3_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10804 ), .force_10(
        \shifter_0/n10805 ), .force_11(1'b0), .QN(n46302) );
  \**FFGEN**  \shifter_0/pre_oi_3_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10808 ), .force_10(
        \shifter_0/n10809 ), .force_11(1'b0), .QN(n46303) );
  \**FFGEN**  \shifter_0/pre_oi_3_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10812 ), .force_10(
        \shifter_0/n10813 ), .force_11(1'b0), .QN(n46304) );
  \**FFGEN**  \shifter_0/pre_oi_3_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10816 ), .force_10(
        \shifter_0/n10817 ), .force_11(1'b0), .QN(n46305) );
  \**FFGEN**  \shifter_0/pre_oi_3_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10820 ), .force_10(
        \shifter_0/n10821 ), .force_11(1'b0), .QN(n46306) );
  \**FFGEN**  \shifter_0/pre_oi_3_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10824 ), .force_10(
        \shifter_0/n10825 ), .force_11(1'b0), .QN(n46307) );
  \**FFGEN**  \shifter_0/pre_oi_3_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10828 ), .force_10(
        \shifter_0/n10829 ), .force_11(1'b0), .QN(n46308) );
  \**FFGEN**  \shifter_0/pre_oi_3_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10832 ), .force_10(
        \shifter_0/n10833 ), .force_11(1'b0), .QN(n46309) );
  \**FFGEN**  \shifter_0/pre_oi_3_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10836 ), .force_10(
        \shifter_0/n10837 ), .force_11(1'b0), .QN(n46310) );
  \**FFGEN**  \shifter_0/pre_oi_3_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10840 ), .force_10(
        \shifter_0/n10841 ), .force_11(1'b0), .QN(n46311) );
  \**FFGEN**  \shifter_0/pre_oi_3_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10844 ), .force_10(
        \shifter_0/n10845 ), .force_11(1'b0), .QN(n46312) );
  \**FFGEN**  \shifter_0/pre_ow_3_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10848 ), .force_10(
        \shifter_0/n10849 ), .force_11(1'b0), .QN(n46613) );
  \**FFGEN**  \shifter_0/pre_ow_3_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10852 ), .force_10(
        \shifter_0/n10853 ), .force_11(1'b0), .QN(n46614) );
  \**FFGEN**  \shifter_0/pre_ow_3_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10856 ), .force_10(
        \shifter_0/n10857 ), .force_11(1'b0), .QN(n46615) );
  \**FFGEN**  \shifter_0/pre_ow_3_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10860 ), .force_10(
        \shifter_0/n10861 ), .force_11(1'b0), .QN(n46616) );
  \**FFGEN**  \shifter_0/pre_ow_3_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10864 ), .force_10(
        \shifter_0/n10865 ), .force_11(1'b0), .QN(n46617) );
  \**FFGEN**  \shifter_0/pre_ow_3_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10868 ), .force_10(
        \shifter_0/n10869 ), .force_11(1'b0), .QN(n46618) );
  \**FFGEN**  \shifter_0/pre_ow_3_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10872 ), .force_10(
        \shifter_0/n10873 ), .force_11(1'b0), .QN(n46619) );
  \**FFGEN**  \shifter_0/pre_ow_3_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10876 ), .force_10(
        \shifter_0/n10877 ), .force_11(1'b0), .QN(n46620) );
  \**FFGEN**  \shifter_0/pre_ow_3_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10880 ), .force_10(
        \shifter_0/n10881 ), .force_11(1'b0), .QN(n46621) );
  \**FFGEN**  \shifter_0/pre_ow_3_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10884 ), .force_10(
        \shifter_0/n10885 ), .force_11(1'b0), .QN(n46622) );
  \**FFGEN**  \shifter_0/pre_ow_3_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10888 ), .force_10(
        \shifter_0/n10889 ), .force_11(1'b0), .QN(n46623) );
  \**FFGEN**  \shifter_0/pre_ow_3_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10892 ), .force_10(
        \shifter_0/n10893 ), .force_11(1'b0), .QN(n46624) );
  \**FFGEN**  \shifter_0/pre_ow_3_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10896 ), .force_10(
        \shifter_0/n10897 ), .force_11(1'b0), .QN(n46625) );
  \**FFGEN**  \shifter_0/pre_ow_3_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10900 ), .force_10(
        \shifter_0/n10901 ), .force_11(1'b0), .QN(n46626) );
  \**FFGEN**  \shifter_0/pre_ow_3_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10904 ), .force_10(
        \shifter_0/n10905 ), .force_11(1'b0), .QN(n46627) );
  \**FFGEN**  \shifter_0/pre_ow_3_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10908 ), .force_10(
        \shifter_0/n10909 ), .force_11(1'b0), .QN(n46628) );
  \**FFGEN**  \shifter_0/pre_ow_3_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10912 ), .force_10(
        \shifter_0/n10913 ), .force_11(1'b0), .QN(n46629) );
  \**FFGEN**  \shifter_0/pre_ow_3_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10916 ), .force_10(
        \shifter_0/n10917 ), .force_11(1'b0), .QN(n46630) );
  \**FFGEN**  \shifter_0/pre_ow_3_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10920 ), .force_10(
        \shifter_0/n10921 ), .force_11(1'b0), .QN(n46631) );
  \**FFGEN**  \shifter_0/pre_ow_3_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10924 ), .force_10(
        \shifter_0/n10925 ), .force_11(1'b0), .QN(n46632) );
  \**FFGEN**  \shifter_0/pre_oi_4_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10928 ), .force_10(
        \shifter_0/n10929 ), .force_11(1'b0), .QN(n46313) );
  \**FFGEN**  \shifter_0/pre_oi_4_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10932 ), .force_10(
        \shifter_0/n10933 ), .force_11(1'b0), .QN(n46314) );
  \**FFGEN**  \shifter_0/pre_oi_4_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10936 ), .force_10(
        \shifter_0/n10937 ), .force_11(1'b0), .QN(n46315) );
  \**FFGEN**  \shifter_0/pre_oi_4_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10940 ), .force_10(
        \shifter_0/n10941 ), .force_11(1'b0), .QN(n46316) );
  \**FFGEN**  \shifter_0/pre_oi_4_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10944 ), .force_10(
        \shifter_0/n10945 ), .force_11(1'b0), .QN(n46317) );
  \**FFGEN**  \shifter_0/pre_oi_4_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10948 ), .force_10(
        \shifter_0/n10949 ), .force_11(1'b0), .QN(n46318) );
  \**FFGEN**  \shifter_0/pre_oi_4_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10952 ), .force_10(
        \shifter_0/n10953 ), .force_11(1'b0), .QN(n46319) );
  \**FFGEN**  \shifter_0/pre_oi_4_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10956 ), .force_10(
        \shifter_0/n10957 ), .force_11(1'b0), .QN(n46320) );
  \**FFGEN**  \shifter_0/pre_oi_4_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10960 ), .force_10(
        \shifter_0/n10961 ), .force_11(1'b0), .QN(n46321) );
  \**FFGEN**  \shifter_0/pre_oi_4_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10964 ), .force_10(
        \shifter_0/n10965 ), .force_11(1'b0), .QN(n46322) );
  \**FFGEN**  \shifter_0/pre_oi_4_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10968 ), .force_10(
        \shifter_0/n10969 ), .force_11(1'b0), .QN(n46323) );
  \**FFGEN**  \shifter_0/pre_oi_4_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10972 ), .force_10(
        \shifter_0/n10973 ), .force_11(1'b0), .QN(n46324) );
  \**FFGEN**  \shifter_0/pre_oi_4_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10976 ), .force_10(
        \shifter_0/n10977 ), .force_11(1'b0), .QN(n46325) );
  \**FFGEN**  \shifter_0/pre_oi_4_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10980 ), .force_10(
        \shifter_0/n10981 ), .force_11(1'b0), .QN(n46326) );
  \**FFGEN**  \shifter_0/pre_oi_4_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10984 ), .force_10(
        \shifter_0/n10985 ), .force_11(1'b0), .QN(n46327) );
  \**FFGEN**  \shifter_0/pre_oi_4_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10988 ), .force_10(
        \shifter_0/n10989 ), .force_11(1'b0), .QN(n46328) );
  \**FFGEN**  \shifter_0/pre_oi_4_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10992 ), .force_10(
        \shifter_0/n10993 ), .force_11(1'b0), .QN(n46329) );
  \**FFGEN**  \shifter_0/pre_oi_4_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10996 ), .force_10(
        \shifter_0/n10997 ), .force_11(1'b0), .QN(n46330) );
  \**FFGEN**  \shifter_0/pre_oi_4_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11000 ), .force_10(
        \shifter_0/n11001 ), .force_11(1'b0), .QN(n46331) );
  \**FFGEN**  \shifter_0/pre_oi_4_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11004 ), .force_10(
        \shifter_0/n11005 ), .force_11(1'b0), .QN(n46332) );
  \**FFGEN**  \shifter_0/pre_ow_4_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11008 ), .force_10(
        \shifter_0/n11009 ), .force_11(1'b0), .QN(n46633) );
  \**FFGEN**  \shifter_0/pre_ow_4_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11012 ), .force_10(
        \shifter_0/n11013 ), .force_11(1'b0), .QN(n46634) );
  \**FFGEN**  \shifter_0/pre_ow_4_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11016 ), .force_10(
        \shifter_0/n11017 ), .force_11(1'b0), .QN(n46635) );
  \**FFGEN**  \shifter_0/pre_ow_4_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11020 ), .force_10(
        \shifter_0/n11021 ), .force_11(1'b0), .QN(n46636) );
  \**FFGEN**  \shifter_0/pre_ow_4_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11024 ), .force_10(
        \shifter_0/n11025 ), .force_11(1'b0), .QN(n46637) );
  \**FFGEN**  \shifter_0/pre_ow_4_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11028 ), .force_10(
        \shifter_0/n11029 ), .force_11(1'b0), .QN(n46638) );
  \**FFGEN**  \shifter_0/pre_ow_4_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11032 ), .force_10(
        \shifter_0/n11033 ), .force_11(1'b0), .QN(n46639) );
  \**FFGEN**  \shifter_0/pre_ow_4_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11036 ), .force_10(
        \shifter_0/n11037 ), .force_11(1'b0), .QN(n46640) );
  \**FFGEN**  \shifter_0/pre_ow_4_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11040 ), .force_10(
        \shifter_0/n11041 ), .force_11(1'b0), .QN(n46641) );
  \**FFGEN**  \shifter_0/pre_ow_4_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11044 ), .force_10(
        \shifter_0/n11045 ), .force_11(1'b0), .QN(n46642) );
  \**FFGEN**  \shifter_0/pre_ow_4_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11048 ), .force_10(
        \shifter_0/n11049 ), .force_11(1'b0), .QN(n46643) );
  \**FFGEN**  \shifter_0/pre_ow_4_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11052 ), .force_10(
        \shifter_0/n11053 ), .force_11(1'b0), .QN(n46644) );
  \**FFGEN**  \shifter_0/pre_ow_4_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11056 ), .force_10(
        \shifter_0/n11057 ), .force_11(1'b0), .QN(n46645) );
  \**FFGEN**  \shifter_0/pre_ow_4_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11060 ), .force_10(
        \shifter_0/n11061 ), .force_11(1'b0), .QN(n46646) );
  \**FFGEN**  \shifter_0/pre_ow_4_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11064 ), .force_10(
        \shifter_0/n11065 ), .force_11(1'b0), .QN(n46647) );
  \**FFGEN**  \shifter_0/pre_ow_4_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11068 ), .force_10(
        \shifter_0/n11069 ), .force_11(1'b0), .QN(n46648) );
  \**FFGEN**  \shifter_0/pre_ow_4_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11072 ), .force_10(
        \shifter_0/n11073 ), .force_11(1'b0), .QN(n46649) );
  \**FFGEN**  \shifter_0/pre_ow_4_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11076 ), .force_10(
        \shifter_0/n11077 ), .force_11(1'b0), .QN(n46650) );
  \**FFGEN**  \shifter_0/pre_ow_4_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11080 ), .force_10(
        \shifter_0/n11081 ), .force_11(1'b0), .QN(n46651) );
  \**FFGEN**  \shifter_0/pre_ow_4_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11084 ), .force_10(
        \shifter_0/n11085 ), .force_11(1'b0), .QN(n46652) );
  \**FFGEN**  \shifter_0/pre_oi_5_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11088 ), .force_10(
        \shifter_0/n11089 ), .force_11(1'b0), .QN(n46333) );
  \**FFGEN**  \shifter_0/pre_oi_5_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11092 ), .force_10(
        \shifter_0/n11093 ), .force_11(1'b0), .QN(n46334) );
  \**FFGEN**  \shifter_0/pre_oi_5_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11096 ), .force_10(
        \shifter_0/n11097 ), .force_11(1'b0), .QN(n46335) );
  \**FFGEN**  \shifter_0/pre_oi_5_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11100 ), .force_10(
        \shifter_0/n11101 ), .force_11(1'b0), .QN(n46336) );
  \**FFGEN**  \shifter_0/pre_oi_5_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11104 ), .force_10(
        \shifter_0/n11105 ), .force_11(1'b0), .QN(n46337) );
  \**FFGEN**  \shifter_0/pre_oi_5_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11108 ), .force_10(
        \shifter_0/n11109 ), .force_11(1'b0), .QN(n46338) );
  \**FFGEN**  \shifter_0/pre_oi_5_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11112 ), .force_10(
        \shifter_0/n11113 ), .force_11(1'b0), .QN(n46339) );
  \**FFGEN**  \shifter_0/pre_oi_5_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11116 ), .force_10(
        \shifter_0/n11117 ), .force_11(1'b0), .QN(n46340) );
  \**FFGEN**  \shifter_0/pre_oi_5_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11120 ), .force_10(
        \shifter_0/n11121 ), .force_11(1'b0), .QN(n46341) );
  \**FFGEN**  \shifter_0/pre_oi_5_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11124 ), .force_10(
        \shifter_0/n11125 ), .force_11(1'b0), .QN(n46342) );
  \**FFGEN**  \shifter_0/pre_oi_5_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11128 ), .force_10(
        \shifter_0/n11129 ), .force_11(1'b0), .QN(n46343) );
  \**FFGEN**  \shifter_0/pre_oi_5_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11132 ), .force_10(
        \shifter_0/n11133 ), .force_11(1'b0), .QN(n46344) );
  \**FFGEN**  \shifter_0/pre_oi_5_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11136 ), .force_10(
        \shifter_0/n11137 ), .force_11(1'b0), .QN(n46345) );
  \**FFGEN**  \shifter_0/pre_oi_5_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11140 ), .force_10(
        \shifter_0/n11141 ), .force_11(1'b0), .QN(n46346) );
  \**FFGEN**  \shifter_0/pre_oi_5_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11144 ), .force_10(
        \shifter_0/n11145 ), .force_11(1'b0), .QN(n46347) );
  \**FFGEN**  \shifter_0/pre_oi_5_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11148 ), .force_10(
        \shifter_0/n11149 ), .force_11(1'b0), .QN(n46348) );
  \**FFGEN**  \shifter_0/pre_oi_5_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11152 ), .force_10(
        \shifter_0/n11153 ), .force_11(1'b0), .QN(n46349) );
  \**FFGEN**  \shifter_0/pre_oi_5_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11156 ), .force_10(
        \shifter_0/n11157 ), .force_11(1'b0), .QN(n46350) );
  \**FFGEN**  \shifter_0/pre_oi_5_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11160 ), .force_10(
        \shifter_0/n11161 ), .force_11(1'b0), .QN(n46351) );
  \**FFGEN**  \shifter_0/pre_oi_5_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11164 ), .force_10(
        \shifter_0/n11165 ), .force_11(1'b0), .QN(n46352) );
  \**FFGEN**  \shifter_0/pre_ow_5_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11168 ), .force_10(
        \shifter_0/n11169 ), .force_11(1'b0), .QN(n46653) );
  \**FFGEN**  \shifter_0/pre_ow_5_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11172 ), .force_10(
        \shifter_0/n11173 ), .force_11(1'b0), .QN(n46654) );
  \**FFGEN**  \shifter_0/pre_ow_5_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11176 ), .force_10(
        \shifter_0/n11177 ), .force_11(1'b0), .QN(n46655) );
  \**FFGEN**  \shifter_0/pre_ow_5_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11180 ), .force_10(
        \shifter_0/n11181 ), .force_11(1'b0), .QN(n46656) );
  \**FFGEN**  \shifter_0/pre_ow_5_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11184 ), .force_10(
        \shifter_0/n11185 ), .force_11(1'b0), .QN(n46657) );
  \**FFGEN**  \shifter_0/pre_ow_5_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11188 ), .force_10(
        \shifter_0/n11189 ), .force_11(1'b0), .QN(n46658) );
  \**FFGEN**  \shifter_0/pre_ow_5_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11192 ), .force_10(
        \shifter_0/n11193 ), .force_11(1'b0), .QN(n46659) );
  \**FFGEN**  \shifter_0/pre_ow_5_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11196 ), .force_10(
        \shifter_0/n11197 ), .force_11(1'b0), .QN(n46660) );
  \**FFGEN**  \shifter_0/pre_ow_5_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11200 ), .force_10(
        \shifter_0/n11201 ), .force_11(1'b0), .QN(n46661) );
  \**FFGEN**  \shifter_0/pre_ow_5_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11204 ), .force_10(
        \shifter_0/n11205 ), .force_11(1'b0), .QN(n46662) );
  \**FFGEN**  \shifter_0/pre_ow_5_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11208 ), .force_10(
        \shifter_0/n11209 ), .force_11(1'b0), .QN(n46663) );
  \**FFGEN**  \shifter_0/pre_ow_5_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11212 ), .force_10(
        \shifter_0/n11213 ), .force_11(1'b0), .QN(n46664) );
  \**FFGEN**  \shifter_0/pre_ow_5_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11216 ), .force_10(
        \shifter_0/n11217 ), .force_11(1'b0), .QN(n46665) );
  \**FFGEN**  \shifter_0/pre_ow_5_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11220 ), .force_10(
        \shifter_0/n11221 ), .force_11(1'b0), .QN(n46666) );
  \**FFGEN**  \shifter_0/pre_ow_5_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11224 ), .force_10(
        \shifter_0/n11225 ), .force_11(1'b0), .QN(n46667) );
  \**FFGEN**  \shifter_0/pre_ow_5_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11228 ), .force_10(
        \shifter_0/n11229 ), .force_11(1'b0), .QN(n46668) );
  \**FFGEN**  \shifter_0/pre_ow_5_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11232 ), .force_10(
        \shifter_0/n11233 ), .force_11(1'b0), .QN(n46669) );
  \**FFGEN**  \shifter_0/pre_ow_5_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11236 ), .force_10(
        \shifter_0/n11237 ), .force_11(1'b0), .QN(n46670) );
  \**FFGEN**  \shifter_0/pre_ow_5_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11240 ), .force_10(
        \shifter_0/n11241 ), .force_11(1'b0), .QN(n46671) );
  \**FFGEN**  \shifter_0/pre_ow_5_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11244 ), .force_10(
        \shifter_0/n11245 ), .force_11(1'b0), .QN(n46672) );
  \**FFGEN**  \shifter_0/pre_oi_6_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11248 ), .force_10(
        \shifter_0/n11249 ), .force_11(1'b0), .QN(n46353) );
  \**FFGEN**  \shifter_0/pre_oi_6_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11252 ), .force_10(
        \shifter_0/n11253 ), .force_11(1'b0), .QN(n46354) );
  \**FFGEN**  \shifter_0/pre_oi_6_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11256 ), .force_10(
        \shifter_0/n11257 ), .force_11(1'b0), .QN(n46355) );
  \**FFGEN**  \shifter_0/pre_oi_6_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11260 ), .force_10(
        \shifter_0/n11261 ), .force_11(1'b0), .QN(n46356) );
  \**FFGEN**  \shifter_0/pre_oi_6_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11264 ), .force_10(
        \shifter_0/n11265 ), .force_11(1'b0), .QN(n46357) );
  \**FFGEN**  \shifter_0/pre_oi_6_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11268 ), .force_10(
        \shifter_0/n11269 ), .force_11(1'b0), .QN(n46358) );
  \**FFGEN**  \shifter_0/pre_oi_6_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11272 ), .force_10(
        \shifter_0/n11273 ), .force_11(1'b0), .QN(n46359) );
  \**FFGEN**  \shifter_0/pre_oi_6_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11276 ), .force_10(
        \shifter_0/n11277 ), .force_11(1'b0), .QN(n46360) );
  \**FFGEN**  \shifter_0/pre_oi_6_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11280 ), .force_10(
        \shifter_0/n11281 ), .force_11(1'b0), .QN(n46361) );
  \**FFGEN**  \shifter_0/pre_oi_6_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11284 ), .force_10(
        \shifter_0/n11285 ), .force_11(1'b0), .QN(n46362) );
  \**FFGEN**  \shifter_0/pre_oi_6_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11288 ), .force_10(
        \shifter_0/n11289 ), .force_11(1'b0), .QN(n46363) );
  \**FFGEN**  \shifter_0/pre_oi_6_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11292 ), .force_10(
        \shifter_0/n11293 ), .force_11(1'b0), .QN(n46364) );
  \**FFGEN**  \shifter_0/pre_oi_6_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11296 ), .force_10(
        \shifter_0/n11297 ), .force_11(1'b0), .QN(n46365) );
  \**FFGEN**  \shifter_0/pre_oi_6_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11300 ), .force_10(
        \shifter_0/n11301 ), .force_11(1'b0), .QN(n46366) );
  \**FFGEN**  \shifter_0/pre_oi_6_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11304 ), .force_10(
        \shifter_0/n11305 ), .force_11(1'b0), .QN(n46367) );
  \**FFGEN**  \shifter_0/pre_oi_6_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11308 ), .force_10(
        \shifter_0/n11309 ), .force_11(1'b0), .QN(n46368) );
  \**FFGEN**  \shifter_0/pre_oi_6_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11312 ), .force_10(
        \shifter_0/n11313 ), .force_11(1'b0), .QN(n46369) );
  \**FFGEN**  \shifter_0/pre_oi_6_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11316 ), .force_10(
        \shifter_0/n11317 ), .force_11(1'b0), .QN(n46370) );
  \**FFGEN**  \shifter_0/pre_oi_6_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11320 ), .force_10(
        \shifter_0/n11321 ), .force_11(1'b0), .QN(n46371) );
  \**FFGEN**  \shifter_0/pre_oi_6_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11324 ), .force_10(
        \shifter_0/n11325 ), .force_11(1'b0), .QN(n46372) );
  \**FFGEN**  \shifter_0/pre_ow_6_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11328 ), .force_10(
        \shifter_0/n11329 ), .force_11(1'b0), .QN(n46673) );
  \**FFGEN**  \shifter_0/pre_ow_6_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11332 ), .force_10(
        \shifter_0/n11333 ), .force_11(1'b0), .QN(n46674) );
  \**FFGEN**  \shifter_0/pre_ow_6_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11336 ), .force_10(
        \shifter_0/n11337 ), .force_11(1'b0), .QN(n46675) );
  \**FFGEN**  \shifter_0/pre_ow_6_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11340 ), .force_10(
        \shifter_0/n11341 ), .force_11(1'b0), .QN(n46676) );
  \**FFGEN**  \shifter_0/pre_ow_6_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11344 ), .force_10(
        \shifter_0/n11345 ), .force_11(1'b0), .QN(n46677) );
  \**FFGEN**  \shifter_0/pre_ow_6_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11348 ), .force_10(
        \shifter_0/n11349 ), .force_11(1'b0), .QN(n46678) );
  \**FFGEN**  \shifter_0/pre_ow_6_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11352 ), .force_10(
        \shifter_0/n11353 ), .force_11(1'b0), .QN(n46679) );
  \**FFGEN**  \shifter_0/pre_ow_6_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11356 ), .force_10(
        \shifter_0/n11357 ), .force_11(1'b0), .QN(n46680) );
  \**FFGEN**  \shifter_0/pre_ow_6_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11360 ), .force_10(
        \shifter_0/n11361 ), .force_11(1'b0), .QN(n46681) );
  \**FFGEN**  \shifter_0/pre_ow_6_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11364 ), .force_10(
        \shifter_0/n11365 ), .force_11(1'b0), .QN(n46682) );
  \**FFGEN**  \shifter_0/pre_ow_6_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11368 ), .force_10(
        \shifter_0/n11369 ), .force_11(1'b0), .QN(n46683) );
  \**FFGEN**  \shifter_0/pre_ow_6_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11372 ), .force_10(
        \shifter_0/n11373 ), .force_11(1'b0), .QN(n46684) );
  \**FFGEN**  \shifter_0/pre_ow_6_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11376 ), .force_10(
        \shifter_0/n11377 ), .force_11(1'b0), .QN(n46685) );
  \**FFGEN**  \shifter_0/pre_ow_6_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11380 ), .force_10(
        \shifter_0/n11381 ), .force_11(1'b0), .QN(n46686) );
  \**FFGEN**  \shifter_0/pre_ow_6_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11384 ), .force_10(
        \shifter_0/n11385 ), .force_11(1'b0), .QN(n46687) );
  \**FFGEN**  \shifter_0/pre_ow_6_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11388 ), .force_10(
        \shifter_0/n11389 ), .force_11(1'b0), .QN(n46688) );
  \**FFGEN**  \shifter_0/pre_ow_6_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11392 ), .force_10(
        \shifter_0/n11393 ), .force_11(1'b0), .QN(n46689) );
  \**FFGEN**  \shifter_0/pre_ow_6_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11396 ), .force_10(
        \shifter_0/n11397 ), .force_11(1'b0), .QN(n46690) );
  \**FFGEN**  \shifter_0/pre_ow_6_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11400 ), .force_10(
        \shifter_0/n11401 ), .force_11(1'b0), .QN(n46691) );
  \**FFGEN**  \shifter_0/pre_ow_6_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11404 ), .force_10(
        \shifter_0/n11405 ), .force_11(1'b0), .QN(n46692) );
  \**FFGEN**  \shifter_0/pre_oi_7_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11408 ), .force_10(
        \shifter_0/n11409 ), .force_11(1'b0), .QN(n46373) );
  \**FFGEN**  \shifter_0/pre_oi_7_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11412 ), .force_10(
        \shifter_0/n11413 ), .force_11(1'b0), .QN(n46374) );
  \**FFGEN**  \shifter_0/pre_oi_7_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11416 ), .force_10(
        \shifter_0/n11417 ), .force_11(1'b0), .QN(n46375) );
  \**FFGEN**  \shifter_0/pre_oi_7_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11420 ), .force_10(
        \shifter_0/n11421 ), .force_11(1'b0), .QN(n46376) );
  \**FFGEN**  \shifter_0/pre_oi_7_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11424 ), .force_10(
        \shifter_0/n11425 ), .force_11(1'b0), .QN(n46377) );
  \**FFGEN**  \shifter_0/pre_oi_7_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11428 ), .force_10(
        \shifter_0/n11429 ), .force_11(1'b0), .QN(n46378) );
  \**FFGEN**  \shifter_0/pre_oi_7_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11432 ), .force_10(
        \shifter_0/n11433 ), .force_11(1'b0), .QN(n46379) );
  \**FFGEN**  \shifter_0/pre_oi_7_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11436 ), .force_10(
        \shifter_0/n11437 ), .force_11(1'b0), .QN(n46380) );
  \**FFGEN**  \shifter_0/pre_oi_7_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11440 ), .force_10(
        \shifter_0/n11441 ), .force_11(1'b0), .QN(n46381) );
  \**FFGEN**  \shifter_0/pre_oi_7_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11444 ), .force_10(
        \shifter_0/n11445 ), .force_11(1'b0), .QN(n46382) );
  \**FFGEN**  \shifter_0/pre_oi_7_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11448 ), .force_10(
        \shifter_0/n11449 ), .force_11(1'b0), .QN(n46383) );
  \**FFGEN**  \shifter_0/pre_oi_7_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11452 ), .force_10(
        \shifter_0/n11453 ), .force_11(1'b0), .QN(n46384) );
  \**FFGEN**  \shifter_0/pre_oi_7_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11456 ), .force_10(
        \shifter_0/n11457 ), .force_11(1'b0), .QN(n46385) );
  \**FFGEN**  \shifter_0/pre_oi_7_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11460 ), .force_10(
        \shifter_0/n11461 ), .force_11(1'b0), .QN(n46386) );
  \**FFGEN**  \shifter_0/pre_oi_7_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11464 ), .force_10(
        \shifter_0/n11465 ), .force_11(1'b0), .QN(n46387) );
  \**FFGEN**  \shifter_0/pre_oi_7_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11468 ), .force_10(
        \shifter_0/n11469 ), .force_11(1'b0), .QN(n46388) );
  \**FFGEN**  \shifter_0/pre_oi_7_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11472 ), .force_10(
        \shifter_0/n11473 ), .force_11(1'b0), .QN(n46389) );
  \**FFGEN**  \shifter_0/pre_oi_7_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11476 ), .force_10(
        \shifter_0/n11477 ), .force_11(1'b0), .QN(n46390) );
  \**FFGEN**  \shifter_0/pre_oi_7_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11480 ), .force_10(
        \shifter_0/n11481 ), .force_11(1'b0), .QN(n46391) );
  \**FFGEN**  \shifter_0/pre_oi_7_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11484 ), .force_10(
        \shifter_0/n11485 ), .force_11(1'b0), .QN(n46392) );
  \**FFGEN**  \shifter_0/pre_ow_7_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11488 ), .force_10(
        \shifter_0/n11489 ), .force_11(1'b0), .QN(n46693) );
  \**FFGEN**  \shifter_0/pre_ow_7_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11492 ), .force_10(
        \shifter_0/n11493 ), .force_11(1'b0), .QN(n46694) );
  \**FFGEN**  \shifter_0/pre_ow_7_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11496 ), .force_10(
        \shifter_0/n11497 ), .force_11(1'b0), .QN(n46695) );
  \**FFGEN**  \shifter_0/pre_ow_7_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11500 ), .force_10(
        \shifter_0/n11501 ), .force_11(1'b0), .QN(n46696) );
  \**FFGEN**  \shifter_0/pre_ow_7_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11504 ), .force_10(
        \shifter_0/n11505 ), .force_11(1'b0), .QN(n46697) );
  \**FFGEN**  \shifter_0/pre_ow_7_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11508 ), .force_10(
        \shifter_0/n11509 ), .force_11(1'b0), .QN(n46698) );
  \**FFGEN**  \shifter_0/pre_ow_7_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11512 ), .force_10(
        \shifter_0/n11513 ), .force_11(1'b0), .QN(n46699) );
  \**FFGEN**  \shifter_0/pre_ow_7_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11516 ), .force_10(
        \shifter_0/n11517 ), .force_11(1'b0), .QN(n46700) );
  \**FFGEN**  \shifter_0/pre_ow_7_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11520 ), .force_10(
        \shifter_0/n11521 ), .force_11(1'b0), .QN(n46701) );
  \**FFGEN**  \shifter_0/pre_ow_7_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11524 ), .force_10(
        \shifter_0/n11525 ), .force_11(1'b0), .QN(n46702) );
  \**FFGEN**  \shifter_0/pre_ow_7_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11528 ), .force_10(
        \shifter_0/n11529 ), .force_11(1'b0), .QN(n46703) );
  \**FFGEN**  \shifter_0/pre_ow_7_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11532 ), .force_10(
        \shifter_0/n11533 ), .force_11(1'b0), .QN(n46704) );
  \**FFGEN**  \shifter_0/pre_ow_7_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11536 ), .force_10(
        \shifter_0/n11537 ), .force_11(1'b0), .QN(n46705) );
  \**FFGEN**  \shifter_0/pre_ow_7_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11540 ), .force_10(
        \shifter_0/n11541 ), .force_11(1'b0), .QN(n46706) );
  \**FFGEN**  \shifter_0/pre_ow_7_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11544 ), .force_10(
        \shifter_0/n11545 ), .force_11(1'b0), .QN(n46707) );
  \**FFGEN**  \shifter_0/pre_ow_7_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11548 ), .force_10(
        \shifter_0/n11549 ), .force_11(1'b0), .QN(n46708) );
  \**FFGEN**  \shifter_0/pre_ow_7_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11552 ), .force_10(
        \shifter_0/n11553 ), .force_11(1'b0), .QN(n46709) );
  \**FFGEN**  \shifter_0/pre_ow_7_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11556 ), .force_10(
        \shifter_0/n11557 ), .force_11(1'b0), .QN(n46710) );
  \**FFGEN**  \shifter_0/pre_ow_7_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11560 ), .force_10(
        \shifter_0/n11561 ), .force_11(1'b0), .QN(n46711) );
  \**FFGEN**  \shifter_0/pre_ow_7_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11564 ), .force_10(
        \shifter_0/n11565 ), .force_11(1'b0), .QN(n46712) );
  \**FFGEN**  \shifter_0/pre_oi_8_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11568 ), .force_10(
        \shifter_0/n11569 ), .force_11(1'b0), .QN(n46393) );
  \**FFGEN**  \shifter_0/pre_oi_8_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11572 ), .force_10(
        \shifter_0/n11573 ), .force_11(1'b0), .QN(n46394) );
  \**FFGEN**  \shifter_0/pre_oi_8_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11576 ), .force_10(
        \shifter_0/n11577 ), .force_11(1'b0), .QN(n46395) );
  \**FFGEN**  \shifter_0/pre_oi_8_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11580 ), .force_10(
        \shifter_0/n11581 ), .force_11(1'b0), .QN(n46396) );
  \**FFGEN**  \shifter_0/pre_oi_8_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11584 ), .force_10(
        \shifter_0/n11585 ), .force_11(1'b0), .QN(n46397) );
  \**FFGEN**  \shifter_0/pre_oi_8_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11588 ), .force_10(
        \shifter_0/n11589 ), .force_11(1'b0), .QN(n46398) );
  \**FFGEN**  \shifter_0/pre_oi_8_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11592 ), .force_10(
        \shifter_0/n11593 ), .force_11(1'b0), .QN(n46399) );
  \**FFGEN**  \shifter_0/pre_oi_8_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11596 ), .force_10(
        \shifter_0/n11597 ), .force_11(1'b0), .QN(n46400) );
  \**FFGEN**  \shifter_0/pre_oi_8_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11600 ), .force_10(
        \shifter_0/n11601 ), .force_11(1'b0), .QN(n46401) );
  \**FFGEN**  \shifter_0/pre_oi_8_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11604 ), .force_10(
        \shifter_0/n11605 ), .force_11(1'b0), .QN(n46402) );
  \**FFGEN**  \shifter_0/pre_oi_8_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11608 ), .force_10(
        \shifter_0/n11609 ), .force_11(1'b0), .QN(n46403) );
  \**FFGEN**  \shifter_0/pre_oi_8_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11612 ), .force_10(
        \shifter_0/n11613 ), .force_11(1'b0), .QN(n46404) );
  \**FFGEN**  \shifter_0/pre_oi_8_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11616 ), .force_10(
        \shifter_0/n11617 ), .force_11(1'b0), .QN(n46405) );
  \**FFGEN**  \shifter_0/pre_oi_8_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11620 ), .force_10(
        \shifter_0/n11621 ), .force_11(1'b0), .QN(n46406) );
  \**FFGEN**  \shifter_0/pre_oi_8_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11624 ), .force_10(
        \shifter_0/n11625 ), .force_11(1'b0), .QN(n46407) );
  \**FFGEN**  \shifter_0/pre_oi_8_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11628 ), .force_10(
        \shifter_0/n11629 ), .force_11(1'b0), .QN(n46408) );
  \**FFGEN**  \shifter_0/pre_oi_8_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11632 ), .force_10(
        \shifter_0/n11633 ), .force_11(1'b0), .QN(n46409) );
  \**FFGEN**  \shifter_0/pre_oi_8_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11636 ), .force_10(
        \shifter_0/n11637 ), .force_11(1'b0), .QN(n46410) );
  \**FFGEN**  \shifter_0/pre_oi_8_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11640 ), .force_10(
        \shifter_0/n11641 ), .force_11(1'b0), .QN(n46411) );
  \**FFGEN**  \shifter_0/pre_oi_8_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11644 ), .force_10(
        \shifter_0/n11645 ), .force_11(1'b0), .QN(n46412) );
  \**FFGEN**  \shifter_0/pre_ow_8_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11648 ), .force_10(
        \shifter_0/n11649 ), .force_11(1'b0), .QN(n46713) );
  \**FFGEN**  \shifter_0/pre_ow_8_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11652 ), .force_10(
        \shifter_0/n11653 ), .force_11(1'b0), .QN(n46714) );
  \**FFGEN**  \shifter_0/pre_ow_8_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11656 ), .force_10(
        \shifter_0/n11657 ), .force_11(1'b0), .QN(n46715) );
  \**FFGEN**  \shifter_0/pre_ow_8_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11660 ), .force_10(
        \shifter_0/n11661 ), .force_11(1'b0), .QN(n46716) );
  \**FFGEN**  \shifter_0/pre_ow_8_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11664 ), .force_10(
        \shifter_0/n11665 ), .force_11(1'b0), .QN(n46717) );
  \**FFGEN**  \shifter_0/pre_ow_8_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11668 ), .force_10(
        \shifter_0/n11669 ), .force_11(1'b0), .QN(n46718) );
  \**FFGEN**  \shifter_0/pre_ow_8_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11672 ), .force_10(
        \shifter_0/n11673 ), .force_11(1'b0), .QN(n46719) );
  \**FFGEN**  \shifter_0/pre_ow_8_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11676 ), .force_10(
        \shifter_0/n11677 ), .force_11(1'b0), .QN(n46720) );
  \**FFGEN**  \shifter_0/pre_ow_8_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11680 ), .force_10(
        \shifter_0/n11681 ), .force_11(1'b0), .QN(n46721) );
  \**FFGEN**  \shifter_0/pre_ow_8_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11684 ), .force_10(
        \shifter_0/n11685 ), .force_11(1'b0), .QN(n46722) );
  \**FFGEN**  \shifter_0/pre_ow_8_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11688 ), .force_10(
        \shifter_0/n11689 ), .force_11(1'b0), .QN(n46723) );
  \**FFGEN**  \shifter_0/pre_ow_8_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11692 ), .force_10(
        \shifter_0/n11693 ), .force_11(1'b0), .QN(n46724) );
  \**FFGEN**  \shifter_0/pre_ow_8_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11696 ), .force_10(
        \shifter_0/n11697 ), .force_11(1'b0), .QN(n46725) );
  \**FFGEN**  \shifter_0/pre_ow_8_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11700 ), .force_10(
        \shifter_0/n11701 ), .force_11(1'b0), .QN(n46726) );
  \**FFGEN**  \shifter_0/pre_ow_8_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11704 ), .force_10(
        \shifter_0/n11705 ), .force_11(1'b0), .QN(n46727) );
  \**FFGEN**  \shifter_0/pre_ow_8_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11708 ), .force_10(
        \shifter_0/n11709 ), .force_11(1'b0), .QN(n46728) );
  \**FFGEN**  \shifter_0/pre_ow_8_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11712 ), .force_10(
        \shifter_0/n11713 ), .force_11(1'b0), .QN(n46729) );
  \**FFGEN**  \shifter_0/pre_ow_8_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11716 ), .force_10(
        \shifter_0/n11717 ), .force_11(1'b0), .QN(n46730) );
  \**FFGEN**  \shifter_0/pre_ow_8_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11720 ), .force_10(
        \shifter_0/n11721 ), .force_11(1'b0), .QN(n46731) );
  \**FFGEN**  \shifter_0/pre_ow_8_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11724 ), .force_10(
        \shifter_0/n11725 ), .force_11(1'b0), .QN(n46732) );
  \**FFGEN**  \shifter_0/pre_oi_9_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11728 ), .force_10(
        n67522), .force_11(1'b0), .QN(n46413) );
  \**FFGEN**  \shifter_0/pre_oi_9_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11732 ), .force_10(
        n67521), .force_11(1'b0), .QN(n46414) );
  \**FFGEN**  \shifter_0/pre_oi_9_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11736 ), .force_10(
        n67520), .force_11(1'b0), .QN(n46415) );
  \**FFGEN**  \shifter_0/pre_oi_9_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11740 ), .force_10(
        n67519), .force_11(1'b0), .QN(n46416) );
  \**FFGEN**  \shifter_0/pre_oi_9_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11744 ), .force_10(
        n67518), .force_11(1'b0), .QN(n46417) );
  \**FFGEN**  \shifter_0/pre_oi_9_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11748 ), .force_10(
        n67517), .force_11(1'b0), .QN(n46418) );
  \**FFGEN**  \shifter_0/pre_oi_9_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11752 ), .force_10(
        n67516), .force_11(1'b0), .QN(n46419) );
  \**FFGEN**  \shifter_0/pre_oi_9_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11756 ), .force_10(
        n67515), .force_11(1'b0), .QN(n46420) );
  \**FFGEN**  \shifter_0/pre_oi_9_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11760 ), .force_10(
        n67514), .force_11(1'b0), .QN(n46421) );
  \**FFGEN**  \shifter_0/pre_oi_9_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11764 ), .force_10(
        n67513), .force_11(1'b0), .QN(n46422) );
  \**FFGEN**  \shifter_0/pre_oi_9_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11768 ), .force_10(
        n67512), .force_11(1'b0), .QN(n46423) );
  \**FFGEN**  \shifter_0/pre_oi_9_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11772 ), .force_10(
        n67511), .force_11(1'b0), .QN(n46424) );
  \**FFGEN**  \shifter_0/pre_oi_9_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11776 ), .force_10(
        n67510), .force_11(1'b0), .QN(n46425) );
  \**FFGEN**  \shifter_0/pre_oi_9_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11780 ), .force_10(
        n67509), .force_11(1'b0), .QN(n46426) );
  \**FFGEN**  \shifter_0/pre_oi_9_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11784 ), .force_10(
        n67508), .force_11(1'b0), .QN(n46427) );
  \**FFGEN**  \shifter_0/pre_oi_9_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11788 ), .force_10(
        n67507), .force_11(1'b0), .QN(n46428) );
  \**FFGEN**  \shifter_0/pre_oi_9_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11792 ), .force_10(
        n67506), .force_11(1'b0), .QN(n46429) );
  \**FFGEN**  \shifter_0/pre_oi_9_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11796 ), .force_10(
        n67505), .force_11(1'b0), .QN(n46430) );
  \**FFGEN**  \shifter_0/pre_oi_9_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11800 ), .force_10(
        n67504), .force_11(1'b0), .QN(n46431) );
  \**FFGEN**  \shifter_0/pre_oi_9_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11804 ), .force_10(
        n67503), .force_11(1'b0), .QN(n46432) );
  \**FFGEN**  \shifter_0/pre_ow_9_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11808 ), .force_10(
        n67182), .force_11(1'b0), .QN(n46733) );
  \**FFGEN**  \shifter_0/pre_ow_9_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11812 ), .force_10(
        n67183), .force_11(1'b0), .QN(n46734) );
  \**FFGEN**  \shifter_0/pre_ow_9_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11816 ), .force_10(
        n67184), .force_11(1'b0), .QN(n46735) );
  \**FFGEN**  \shifter_0/pre_ow_9_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11820 ), .force_10(
        n67185), .force_11(1'b0), .QN(n46736) );
  \**FFGEN**  \shifter_0/pre_ow_9_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11824 ), .force_10(
        n67186), .force_11(1'b0), .QN(n46737) );
  \**FFGEN**  \shifter_0/pre_ow_9_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11828 ), .force_10(
        n67187), .force_11(1'b0), .QN(n46738) );
  \**FFGEN**  \shifter_0/pre_ow_9_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11832 ), .force_10(
        n67188), .force_11(1'b0), .QN(n46739) );
  \**FFGEN**  \shifter_0/pre_ow_9_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11836 ), .force_10(
        n67189), .force_11(1'b0), .QN(n46740) );
  \**FFGEN**  \shifter_0/pre_ow_9_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11840 ), .force_10(
        n67190), .force_11(1'b0), .QN(n46741) );
  \**FFGEN**  \shifter_0/pre_ow_9_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11844 ), .force_10(
        n67191), .force_11(1'b0), .QN(n46742) );
  \**FFGEN**  \shifter_0/pre_ow_9_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11848 ), .force_10(
        n67192), .force_11(1'b0), .QN(n46743) );
  \**FFGEN**  \shifter_0/pre_ow_9_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11852 ), .force_10(
        n67193), .force_11(1'b0), .QN(n46744) );
  \**FFGEN**  \shifter_0/pre_ow_9_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11856 ), .force_10(
        n67194), .force_11(1'b0), .QN(n46745) );
  \**FFGEN**  \shifter_0/pre_ow_9_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11860 ), .force_10(
        n67195), .force_11(1'b0), .QN(n46746) );
  \**FFGEN**  \shifter_0/pre_ow_9_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11864 ), .force_10(
        n67196), .force_11(1'b0), .QN(n46747) );
  \**FFGEN**  \shifter_0/pre_ow_9_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11868 ), .force_10(
        n67197), .force_11(1'b0), .QN(n46748) );
  \**FFGEN**  \shifter_0/pre_ow_9_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11872 ), .force_10(
        n67198), .force_11(1'b0), .QN(n46749) );
  \**FFGEN**  \shifter_0/pre_ow_9_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11876 ), .force_10(
        n67199), .force_11(1'b0), .QN(n46750) );
  \**FFGEN**  \shifter_0/pre_ow_9_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11880 ), .force_10(
        n67200), .force_11(1'b0), .QN(n46751) );
  \**FFGEN**  \shifter_0/pre_ow_9_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11884 ), .force_10(
        n67201), .force_11(1'b0), .QN(n46752) );
  \**FFGEN**  \shifter_0/pre_oi_10_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11888 ), .force_10(
        \shifter_0/n11889 ), .force_11(1'b0), .QN(n46433) );
  \**FFGEN**  \shifter_0/pre_oi_10_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11892 ), .force_10(
        \shifter_0/n11893 ), .force_11(1'b0), .QN(n46434) );
  \**FFGEN**  \shifter_0/pre_oi_10_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11896 ), .force_10(
        \shifter_0/n11897 ), .force_11(1'b0), .QN(n46435) );
  \**FFGEN**  \shifter_0/pre_oi_10_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11900 ), .force_10(
        \shifter_0/n11901 ), .force_11(1'b0), .QN(n46436) );
  \**FFGEN**  \shifter_0/pre_oi_10_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11904 ), .force_10(
        \shifter_0/n11905 ), .force_11(1'b0), .QN(n46437) );
  \**FFGEN**  \shifter_0/pre_oi_10_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11908 ), .force_10(
        \shifter_0/n11909 ), .force_11(1'b0), .QN(n46438) );
  \**FFGEN**  \shifter_0/pre_oi_10_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11912 ), .force_10(
        \shifter_0/n11913 ), .force_11(1'b0), .QN(n46439) );
  \**FFGEN**  \shifter_0/pre_oi_10_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11916 ), .force_10(
        \shifter_0/n11917 ), .force_11(1'b0), .QN(n46440) );
  \**FFGEN**  \shifter_0/pre_oi_10_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11920 ), .force_10(
        \shifter_0/n11921 ), .force_11(1'b0), .QN(n46441) );
  \**FFGEN**  \shifter_0/pre_oi_10_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11924 ), .force_10(
        \shifter_0/n11925 ), .force_11(1'b0), .QN(n46442) );
  \**FFGEN**  \shifter_0/pre_oi_10_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11928 ), .force_10(
        \shifter_0/n11929 ), .force_11(1'b0), .QN(n46443) );
  \**FFGEN**  \shifter_0/pre_oi_10_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11932 ), .force_10(
        \shifter_0/n11933 ), .force_11(1'b0), .QN(n46444) );
  \**FFGEN**  \shifter_0/pre_oi_10_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11936 ), .force_10(
        \shifter_0/n11937 ), .force_11(1'b0), .QN(n46445) );
  \**FFGEN**  \shifter_0/pre_oi_10_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11940 ), .force_10(
        \shifter_0/n11941 ), .force_11(1'b0), .QN(n46446) );
  \**FFGEN**  \shifter_0/pre_oi_10_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11944 ), .force_10(
        \shifter_0/n11945 ), .force_11(1'b0), .QN(n46447) );
  \**FFGEN**  \shifter_0/pre_oi_10_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11948 ), .force_10(
        \shifter_0/n11949 ), .force_11(1'b0), .QN(n46448) );
  \**FFGEN**  \shifter_0/pre_oi_10_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11952 ), .force_10(
        \shifter_0/n11953 ), .force_11(1'b0), .QN(n46449) );
  \**FFGEN**  \shifter_0/pre_oi_10_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11956 ), .force_10(
        \shifter_0/n11957 ), .force_11(1'b0), .QN(n46450) );
  \**FFGEN**  \shifter_0/pre_oi_10_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11960 ), .force_10(
        \shifter_0/n11961 ), .force_11(1'b0), .QN(n46451) );
  \**FFGEN**  \shifter_0/pre_oi_10_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11964 ), .force_10(
        \shifter_0/n11965 ), .force_11(1'b0), .QN(n46452) );
  \**FFGEN**  \shifter_0/pre_ow_10_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11968 ), .force_10(
        \shifter_0/n11969 ), .force_11(1'b0), .QN(n46753) );
  \**FFGEN**  \shifter_0/pre_ow_10_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11972 ), .force_10(
        \shifter_0/n11973 ), .force_11(1'b0), .QN(n46754) );
  \**FFGEN**  \shifter_0/pre_ow_10_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11976 ), .force_10(
        \shifter_0/n11977 ), .force_11(1'b0), .QN(n46755) );
  \**FFGEN**  \shifter_0/pre_ow_10_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11980 ), .force_10(
        \shifter_0/n11981 ), .force_11(1'b0), .QN(n46756) );
  \**FFGEN**  \shifter_0/pre_ow_10_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11984 ), .force_10(
        \shifter_0/n11985 ), .force_11(1'b0), .QN(n46757) );
  \**FFGEN**  \shifter_0/pre_ow_10_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11988 ), .force_10(
        \shifter_0/n11989 ), .force_11(1'b0), .QN(n46758) );
  \**FFGEN**  \shifter_0/pre_ow_10_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11992 ), .force_10(
        \shifter_0/n11993 ), .force_11(1'b0), .QN(n46759) );
  \**FFGEN**  \shifter_0/pre_ow_10_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n11996 ), .force_10(
        \shifter_0/n11997 ), .force_11(1'b0), .QN(n46760) );
  \**FFGEN**  \shifter_0/pre_ow_10_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12000 ), .force_10(
        \shifter_0/n12001 ), .force_11(1'b0), .QN(n46761) );
  \**FFGEN**  \shifter_0/pre_ow_10_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12004 ), .force_10(
        \shifter_0/n12005 ), .force_11(1'b0), .QN(n46762) );
  \**FFGEN**  \shifter_0/pre_ow_10_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12008 ), .force_10(
        \shifter_0/n12009 ), .force_11(1'b0), .QN(n46763) );
  \**FFGEN**  \shifter_0/pre_ow_10_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12012 ), .force_10(
        \shifter_0/n12013 ), .force_11(1'b0), .QN(n46764) );
  \**FFGEN**  \shifter_0/pre_ow_10_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12016 ), .force_10(
        \shifter_0/n12017 ), .force_11(1'b0), .QN(n46765) );
  \**FFGEN**  \shifter_0/pre_ow_10_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12020 ), .force_10(
        \shifter_0/n12021 ), .force_11(1'b0), .QN(n46766) );
  \**FFGEN**  \shifter_0/pre_ow_10_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12024 ), .force_10(
        \shifter_0/n12025 ), .force_11(1'b0), .QN(n46767) );
  \**FFGEN**  \shifter_0/pre_ow_10_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12028 ), .force_10(
        \shifter_0/n12029 ), .force_11(1'b0), .QN(n46768) );
  \**FFGEN**  \shifter_0/pre_ow_10_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12032 ), .force_10(
        \shifter_0/n12033 ), .force_11(1'b0), .QN(n46769) );
  \**FFGEN**  \shifter_0/pre_ow_10_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12036 ), .force_10(
        \shifter_0/n12037 ), .force_11(1'b0), .QN(n46770) );
  \**FFGEN**  \shifter_0/pre_ow_10_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12040 ), .force_10(
        \shifter_0/n12041 ), .force_11(1'b0), .QN(n46771) );
  \**FFGEN**  \shifter_0/pre_ow_10_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12044 ), .force_10(
        \shifter_0/n12045 ), .force_11(1'b0), .QN(n46772) );
  \**FFGEN**  \shifter_0/pre_oi_11_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12048 ), .force_10(
        \shifter_0/n12049 ), .force_11(1'b0), .QN(n46453) );
  \**FFGEN**  \shifter_0/pre_oi_11_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12052 ), .force_10(
        \shifter_0/n12053 ), .force_11(1'b0), .QN(n46454) );
  \**FFGEN**  \shifter_0/pre_oi_11_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12056 ), .force_10(
        \shifter_0/n12057 ), .force_11(1'b0), .QN(n46455) );
  \**FFGEN**  \shifter_0/pre_oi_11_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12060 ), .force_10(
        \shifter_0/n12061 ), .force_11(1'b0), .QN(n46456) );
  \**FFGEN**  \shifter_0/pre_oi_11_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12064 ), .force_10(
        \shifter_0/n12065 ), .force_11(1'b0), .QN(n46457) );
  \**FFGEN**  \shifter_0/pre_oi_11_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12068 ), .force_10(
        \shifter_0/n12069 ), .force_11(1'b0), .QN(n46458) );
  \**FFGEN**  \shifter_0/pre_oi_11_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12072 ), .force_10(
        \shifter_0/n12073 ), .force_11(1'b0), .QN(n46459) );
  \**FFGEN**  \shifter_0/pre_oi_11_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12076 ), .force_10(
        \shifter_0/n12077 ), .force_11(1'b0), .QN(n46460) );
  \**FFGEN**  \shifter_0/pre_oi_11_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12080 ), .force_10(
        \shifter_0/n12081 ), .force_11(1'b0), .QN(n46461) );
  \**FFGEN**  \shifter_0/pre_oi_11_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12084 ), .force_10(
        \shifter_0/n12085 ), .force_11(1'b0), .QN(n46462) );
  \**FFGEN**  \shifter_0/pre_oi_11_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12088 ), .force_10(
        \shifter_0/n12089 ), .force_11(1'b0), .QN(n46463) );
  \**FFGEN**  \shifter_0/pre_oi_11_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12092 ), .force_10(
        \shifter_0/n12093 ), .force_11(1'b0), .QN(n46464) );
  \**FFGEN**  \shifter_0/pre_oi_11_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12096 ), .force_10(
        \shifter_0/n12097 ), .force_11(1'b0), .QN(n46465) );
  \**FFGEN**  \shifter_0/pre_oi_11_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12100 ), .force_10(
        \shifter_0/n12101 ), .force_11(1'b0), .QN(n46466) );
  \**FFGEN**  \shifter_0/pre_oi_11_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12104 ), .force_10(
        \shifter_0/n12105 ), .force_11(1'b0), .QN(n46467) );
  \**FFGEN**  \shifter_0/pre_oi_11_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12108 ), .force_10(
        \shifter_0/n12109 ), .force_11(1'b0), .QN(n46468) );
  \**FFGEN**  \shifter_0/pre_oi_11_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12112 ), .force_10(
        \shifter_0/n12113 ), .force_11(1'b0), .QN(n46469) );
  \**FFGEN**  \shifter_0/pre_oi_11_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12116 ), .force_10(
        \shifter_0/n12117 ), .force_11(1'b0), .QN(n46470) );
  \**FFGEN**  \shifter_0/pre_oi_11_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12120 ), .force_10(
        \shifter_0/n12121 ), .force_11(1'b0), .QN(n46471) );
  \**FFGEN**  \shifter_0/pre_oi_11_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12124 ), .force_10(
        \shifter_0/n12125 ), .force_11(1'b0), .QN(n46472) );
  \**FFGEN**  \shifter_0/pre_ow_11_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12128 ), .force_10(
        \shifter_0/n12129 ), .force_11(1'b0), .QN(n46773) );
  \**FFGEN**  \shifter_0/pre_ow_11_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12132 ), .force_10(
        \shifter_0/n12133 ), .force_11(1'b0), .QN(n46774) );
  \**FFGEN**  \shifter_0/pre_ow_11_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12136 ), .force_10(
        \shifter_0/n12137 ), .force_11(1'b0), .QN(n46775) );
  \**FFGEN**  \shifter_0/pre_ow_11_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12140 ), .force_10(
        \shifter_0/n12141 ), .force_11(1'b0), .QN(n46776) );
  \**FFGEN**  \shifter_0/pre_ow_11_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12144 ), .force_10(
        \shifter_0/n12145 ), .force_11(1'b0), .QN(n46777) );
  \**FFGEN**  \shifter_0/pre_ow_11_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12148 ), .force_10(
        \shifter_0/n12149 ), .force_11(1'b0), .QN(n46778) );
  \**FFGEN**  \shifter_0/pre_ow_11_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12152 ), .force_10(
        \shifter_0/n12153 ), .force_11(1'b0), .QN(n46779) );
  \**FFGEN**  \shifter_0/pre_ow_11_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12156 ), .force_10(
        \shifter_0/n12157 ), .force_11(1'b0), .QN(n46780) );
  \**FFGEN**  \shifter_0/pre_ow_11_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12160 ), .force_10(
        \shifter_0/n12161 ), .force_11(1'b0), .QN(n46781) );
  \**FFGEN**  \shifter_0/pre_ow_11_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12164 ), .force_10(
        \shifter_0/n12165 ), .force_11(1'b0), .QN(n46782) );
  \**FFGEN**  \shifter_0/pre_ow_11_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12168 ), .force_10(
        \shifter_0/n12169 ), .force_11(1'b0), .QN(n46783) );
  \**FFGEN**  \shifter_0/pre_ow_11_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12172 ), .force_10(
        \shifter_0/n12173 ), .force_11(1'b0), .QN(n46784) );
  \**FFGEN**  \shifter_0/pre_ow_11_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12176 ), .force_10(
        \shifter_0/n12177 ), .force_11(1'b0), .QN(n46785) );
  \**FFGEN**  \shifter_0/pre_ow_11_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12180 ), .force_10(
        \shifter_0/n12181 ), .force_11(1'b0), .QN(n46786) );
  \**FFGEN**  \shifter_0/pre_ow_11_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12184 ), .force_10(
        \shifter_0/n12185 ), .force_11(1'b0), .QN(n46787) );
  \**FFGEN**  \shifter_0/pre_ow_11_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12188 ), .force_10(
        \shifter_0/n12189 ), .force_11(1'b0), .QN(n46788) );
  \**FFGEN**  \shifter_0/pre_ow_11_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12192 ), .force_10(
        \shifter_0/n12193 ), .force_11(1'b0), .QN(n46789) );
  \**FFGEN**  \shifter_0/pre_ow_11_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12196 ), .force_10(
        \shifter_0/n12197 ), .force_11(1'b0), .QN(n46790) );
  \**FFGEN**  \shifter_0/pre_ow_11_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12200 ), .force_10(
        \shifter_0/n12201 ), .force_11(1'b0), .QN(n46791) );
  \**FFGEN**  \shifter_0/pre_ow_11_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12204 ), .force_10(
        \shifter_0/n12205 ), .force_11(1'b0), .QN(n46792) );
  \**FFGEN**  \shifter_0/pre_oi_12_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12208 ), .force_10(
        \shifter_0/n12209 ), .force_11(1'b0), .QN(n46473) );
  \**FFGEN**  \shifter_0/pre_oi_12_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12212 ), .force_10(
        \shifter_0/n12213 ), .force_11(1'b0), .QN(n46474) );
  \**FFGEN**  \shifter_0/pre_oi_12_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12216 ), .force_10(
        \shifter_0/n12217 ), .force_11(1'b0), .QN(n46475) );
  \**FFGEN**  \shifter_0/pre_oi_12_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12220 ), .force_10(
        \shifter_0/n12221 ), .force_11(1'b0), .QN(n46476) );
  \**FFGEN**  \shifter_0/pre_oi_12_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12224 ), .force_10(
        \shifter_0/n12225 ), .force_11(1'b0), .QN(n46477) );
  \**FFGEN**  \shifter_0/pre_oi_12_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12228 ), .force_10(
        \shifter_0/n12229 ), .force_11(1'b0), .QN(n46478) );
  \**FFGEN**  \shifter_0/pre_oi_12_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12232 ), .force_10(
        \shifter_0/n12233 ), .force_11(1'b0), .QN(n46479) );
  \**FFGEN**  \shifter_0/pre_oi_12_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12236 ), .force_10(
        \shifter_0/n12237 ), .force_11(1'b0), .QN(n46480) );
  \**FFGEN**  \shifter_0/pre_oi_12_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12240 ), .force_10(
        \shifter_0/n12241 ), .force_11(1'b0), .QN(n46481) );
  \**FFGEN**  \shifter_0/pre_oi_12_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12244 ), .force_10(
        \shifter_0/n12245 ), .force_11(1'b0), .QN(n46482) );
  \**FFGEN**  \shifter_0/pre_oi_12_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12248 ), .force_10(
        \shifter_0/n12249 ), .force_11(1'b0), .QN(n46483) );
  \**FFGEN**  \shifter_0/pre_oi_12_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12252 ), .force_10(
        \shifter_0/n12253 ), .force_11(1'b0), .QN(n46484) );
  \**FFGEN**  \shifter_0/pre_oi_12_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12256 ), .force_10(
        \shifter_0/n12257 ), .force_11(1'b0), .QN(n46485) );
  \**FFGEN**  \shifter_0/pre_oi_12_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12260 ), .force_10(
        \shifter_0/n12261 ), .force_11(1'b0), .QN(n46486) );
  \**FFGEN**  \shifter_0/pre_oi_12_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12264 ), .force_10(
        \shifter_0/n12265 ), .force_11(1'b0), .QN(n46487) );
  \**FFGEN**  \shifter_0/pre_oi_12_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12268 ), .force_10(
        \shifter_0/n12269 ), .force_11(1'b0), .QN(n46488) );
  \**FFGEN**  \shifter_0/pre_oi_12_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12272 ), .force_10(
        \shifter_0/n12273 ), .force_11(1'b0), .QN(n46489) );
  \**FFGEN**  \shifter_0/pre_oi_12_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12276 ), .force_10(
        \shifter_0/n12277 ), .force_11(1'b0), .QN(n46490) );
  \**FFGEN**  \shifter_0/pre_oi_12_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12280 ), .force_10(
        \shifter_0/n12281 ), .force_11(1'b0), .QN(n46491) );
  \**FFGEN**  \shifter_0/pre_oi_12_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12284 ), .force_10(
        \shifter_0/n12285 ), .force_11(1'b0), .QN(n46492) );
  \**FFGEN**  \shifter_0/pre_ow_12_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12288 ), .force_10(
        \shifter_0/n12289 ), .force_11(1'b0), .QN(n46793) );
  \**FFGEN**  \shifter_0/pre_ow_12_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12292 ), .force_10(
        \shifter_0/n12293 ), .force_11(1'b0), .QN(n46794) );
  \**FFGEN**  \shifter_0/pre_ow_12_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12296 ), .force_10(
        \shifter_0/n12297 ), .force_11(1'b0), .QN(n46795) );
  \**FFGEN**  \shifter_0/pre_ow_12_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12300 ), .force_10(
        \shifter_0/n12301 ), .force_11(1'b0), .QN(n46796) );
  \**FFGEN**  \shifter_0/pre_ow_12_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12304 ), .force_10(
        \shifter_0/n12305 ), .force_11(1'b0), .QN(n46797) );
  \**FFGEN**  \shifter_0/pre_ow_12_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12308 ), .force_10(
        \shifter_0/n12309 ), .force_11(1'b0), .QN(n46798) );
  \**FFGEN**  \shifter_0/pre_ow_12_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12312 ), .force_10(
        \shifter_0/n12313 ), .force_11(1'b0), .QN(n46799) );
  \**FFGEN**  \shifter_0/pre_ow_12_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12316 ), .force_10(
        \shifter_0/n12317 ), .force_11(1'b0), .QN(n46800) );
  \**FFGEN**  \shifter_0/pre_ow_12_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12320 ), .force_10(
        \shifter_0/n12321 ), .force_11(1'b0), .QN(n46801) );
  \**FFGEN**  \shifter_0/pre_ow_12_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12324 ), .force_10(
        \shifter_0/n12325 ), .force_11(1'b0), .QN(n46802) );
  \**FFGEN**  \shifter_0/pre_ow_12_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12328 ), .force_10(
        \shifter_0/n12329 ), .force_11(1'b0), .QN(n46803) );
  \**FFGEN**  \shifter_0/pre_ow_12_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12332 ), .force_10(
        \shifter_0/n12333 ), .force_11(1'b0), .QN(n46804) );
  \**FFGEN**  \shifter_0/pre_ow_12_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12336 ), .force_10(
        \shifter_0/n12337 ), .force_11(1'b0), .QN(n46805) );
  \**FFGEN**  \shifter_0/pre_ow_12_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12340 ), .force_10(
        \shifter_0/n12341 ), .force_11(1'b0), .QN(n46806) );
  \**FFGEN**  \shifter_0/pre_ow_12_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12344 ), .force_10(
        \shifter_0/n12345 ), .force_11(1'b0), .QN(n46807) );
  \**FFGEN**  \shifter_0/pre_ow_12_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12348 ), .force_10(
        \shifter_0/n12349 ), .force_11(1'b0), .QN(n46808) );
  \**FFGEN**  \shifter_0/pre_ow_12_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12352 ), .force_10(
        \shifter_0/n12353 ), .force_11(1'b0), .QN(n46809) );
  \**FFGEN**  \shifter_0/pre_ow_12_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12356 ), .force_10(
        \shifter_0/n12357 ), .force_11(1'b0), .QN(n46810) );
  \**FFGEN**  \shifter_0/pre_ow_12_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12360 ), .force_10(
        \shifter_0/n12361 ), .force_11(1'b0), .QN(n46811) );
  \**FFGEN**  \shifter_0/pre_ow_12_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12364 ), .force_10(
        \shifter_0/n12365 ), .force_11(1'b0), .QN(n46812) );
  \**FFGEN**  \shifter_0/pre_oi_13_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12368 ), .force_10(
        \shifter_0/n12369 ), .force_11(1'b0), .QN(n46493) );
  \**FFGEN**  \shifter_0/pre_oi_13_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12372 ), .force_10(
        \shifter_0/n12373 ), .force_11(1'b0), .QN(n46494) );
  \**FFGEN**  \shifter_0/pre_oi_13_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12376 ), .force_10(
        \shifter_0/n12377 ), .force_11(1'b0), .QN(n46495) );
  \**FFGEN**  \shifter_0/pre_oi_13_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12380 ), .force_10(
        \shifter_0/n12381 ), .force_11(1'b0), .QN(n46496) );
  \**FFGEN**  \shifter_0/pre_oi_13_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12384 ), .force_10(
        \shifter_0/n12385 ), .force_11(1'b0), .QN(n46497) );
  \**FFGEN**  \shifter_0/pre_oi_13_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12388 ), .force_10(
        \shifter_0/n12389 ), .force_11(1'b0), .QN(n46498) );
  \**FFGEN**  \shifter_0/pre_oi_13_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12392 ), .force_10(
        \shifter_0/n12393 ), .force_11(1'b0), .QN(n46499) );
  \**FFGEN**  \shifter_0/pre_oi_13_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12396 ), .force_10(
        \shifter_0/n12397 ), .force_11(1'b0), .QN(n46500) );
  \**FFGEN**  \shifter_0/pre_oi_13_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12400 ), .force_10(
        \shifter_0/n12401 ), .force_11(1'b0), .QN(n46501) );
  \**FFGEN**  \shifter_0/pre_oi_13_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12404 ), .force_10(
        \shifter_0/n12405 ), .force_11(1'b0), .QN(n46502) );
  \**FFGEN**  \shifter_0/pre_oi_13_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12408 ), .force_10(
        \shifter_0/n12409 ), .force_11(1'b0), .QN(n46503) );
  \**FFGEN**  \shifter_0/pre_oi_13_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12412 ), .force_10(
        \shifter_0/n12413 ), .force_11(1'b0), .QN(n46504) );
  \**FFGEN**  \shifter_0/pre_oi_13_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12416 ), .force_10(
        \shifter_0/n12417 ), .force_11(1'b0), .QN(n46505) );
  \**FFGEN**  \shifter_0/pre_oi_13_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12420 ), .force_10(
        \shifter_0/n12421 ), .force_11(1'b0), .QN(n46506) );
  \**FFGEN**  \shifter_0/pre_oi_13_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12424 ), .force_10(
        \shifter_0/n12425 ), .force_11(1'b0), .QN(n46507) );
  \**FFGEN**  \shifter_0/pre_oi_13_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12428 ), .force_10(
        \shifter_0/n12429 ), .force_11(1'b0), .QN(n46508) );
  \**FFGEN**  \shifter_0/pre_oi_13_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12432 ), .force_10(
        \shifter_0/n12433 ), .force_11(1'b0), .QN(n46509) );
  \**FFGEN**  \shifter_0/pre_oi_13_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12436 ), .force_10(
        \shifter_0/n12437 ), .force_11(1'b0), .QN(n46510) );
  \**FFGEN**  \shifter_0/pre_oi_13_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12440 ), .force_10(
        \shifter_0/n12441 ), .force_11(1'b0), .QN(n46511) );
  \**FFGEN**  \shifter_0/pre_oi_13_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12444 ), .force_10(
        \shifter_0/n12445 ), .force_11(1'b0), .QN(n46512) );
  \**FFGEN**  \shifter_0/pre_ow_13_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12448 ), .force_10(
        \shifter_0/n12449 ), .force_11(1'b0), .QN(n46813) );
  \**FFGEN**  \shifter_0/pre_ow_13_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12452 ), .force_10(
        \shifter_0/n12453 ), .force_11(1'b0), .QN(n46814) );
  \**FFGEN**  \shifter_0/pre_ow_13_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12456 ), .force_10(
        \shifter_0/n12457 ), .force_11(1'b0), .QN(n46815) );
  \**FFGEN**  \shifter_0/pre_ow_13_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12460 ), .force_10(
        \shifter_0/n12461 ), .force_11(1'b0), .QN(n46816) );
  \**FFGEN**  \shifter_0/pre_ow_13_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12464 ), .force_10(
        \shifter_0/n12465 ), .force_11(1'b0), .QN(n46817) );
  \**FFGEN**  \shifter_0/pre_ow_13_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12468 ), .force_10(
        \shifter_0/n12469 ), .force_11(1'b0), .QN(n46818) );
  \**FFGEN**  \shifter_0/pre_ow_13_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12472 ), .force_10(
        \shifter_0/n12473 ), .force_11(1'b0), .QN(n46819) );
  \**FFGEN**  \shifter_0/pre_ow_13_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12476 ), .force_10(
        \shifter_0/n12477 ), .force_11(1'b0), .QN(n46820) );
  \**FFGEN**  \shifter_0/pre_ow_13_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12480 ), .force_10(
        \shifter_0/n12481 ), .force_11(1'b0), .QN(n46821) );
  \**FFGEN**  \shifter_0/pre_ow_13_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12484 ), .force_10(
        \shifter_0/n12485 ), .force_11(1'b0), .QN(n46822) );
  \**FFGEN**  \shifter_0/pre_ow_13_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12488 ), .force_10(
        \shifter_0/n12489 ), .force_11(1'b0), .QN(n46823) );
  \**FFGEN**  \shifter_0/pre_ow_13_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12492 ), .force_10(
        \shifter_0/n12493 ), .force_11(1'b0), .QN(n46824) );
  \**FFGEN**  \shifter_0/pre_ow_13_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12496 ), .force_10(
        \shifter_0/n12497 ), .force_11(1'b0), .QN(n46825) );
  \**FFGEN**  \shifter_0/pre_ow_13_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12500 ), .force_10(
        \shifter_0/n12501 ), .force_11(1'b0), .QN(n46826) );
  \**FFGEN**  \shifter_0/pre_ow_13_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12504 ), .force_10(
        \shifter_0/n12505 ), .force_11(1'b0), .QN(n46827) );
  \**FFGEN**  \shifter_0/pre_ow_13_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12508 ), .force_10(
        \shifter_0/n12509 ), .force_11(1'b0), .QN(n46828) );
  \**FFGEN**  \shifter_0/pre_ow_13_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12512 ), .force_10(
        \shifter_0/n12513 ), .force_11(1'b0), .QN(n46829) );
  \**FFGEN**  \shifter_0/pre_ow_13_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12516 ), .force_10(
        \shifter_0/n12517 ), .force_11(1'b0), .QN(n46830) );
  \**FFGEN**  \shifter_0/pre_ow_13_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12520 ), .force_10(
        \shifter_0/n12521 ), .force_11(1'b0), .QN(n46831) );
  \**FFGEN**  \shifter_0/pre_ow_13_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12524 ), .force_10(
        \shifter_0/n12525 ), .force_11(1'b0), .QN(n46832) );
  \**FFGEN**  \shifter_0/pre_oi_14_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12528 ), .force_10(
        \shifter_0/n12529 ), .force_11(1'b0), .QN(n46513) );
  \**FFGEN**  \shifter_0/pre_oi_14_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12532 ), .force_10(
        \shifter_0/n12533 ), .force_11(1'b0), .QN(n46514) );
  \**FFGEN**  \shifter_0/pre_oi_14_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12536 ), .force_10(
        \shifter_0/n12537 ), .force_11(1'b0), .QN(n46515) );
  \**FFGEN**  \shifter_0/pre_oi_14_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12540 ), .force_10(
        \shifter_0/n12541 ), .force_11(1'b0), .QN(n46516) );
  \**FFGEN**  \shifter_0/pre_oi_14_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12544 ), .force_10(
        \shifter_0/n12545 ), .force_11(1'b0), .QN(n46517) );
  \**FFGEN**  \shifter_0/pre_oi_14_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12548 ), .force_10(
        \shifter_0/n12549 ), .force_11(1'b0), .QN(n46518) );
  \**FFGEN**  \shifter_0/pre_oi_14_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12552 ), .force_10(
        \shifter_0/n12553 ), .force_11(1'b0), .QN(n46519) );
  \**FFGEN**  \shifter_0/pre_oi_14_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12556 ), .force_10(
        \shifter_0/n12557 ), .force_11(1'b0), .QN(n46520) );
  \**FFGEN**  \shifter_0/pre_oi_14_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12560 ), .force_10(
        \shifter_0/n12561 ), .force_11(1'b0), .QN(n46521) );
  \**FFGEN**  \shifter_0/pre_oi_14_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12564 ), .force_10(
        \shifter_0/n12565 ), .force_11(1'b0), .QN(n46522) );
  \**FFGEN**  \shifter_0/pre_oi_14_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12568 ), .force_10(
        \shifter_0/n12569 ), .force_11(1'b0), .QN(n46523) );
  \**FFGEN**  \shifter_0/pre_oi_14_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12572 ), .force_10(
        \shifter_0/n12573 ), .force_11(1'b0), .QN(n46524) );
  \**FFGEN**  \shifter_0/pre_oi_14_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12576 ), .force_10(
        \shifter_0/n12577 ), .force_11(1'b0), .QN(n46525) );
  \**FFGEN**  \shifter_0/pre_oi_14_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12580 ), .force_10(
        \shifter_0/n12581 ), .force_11(1'b0), .QN(n46526) );
  \**FFGEN**  \shifter_0/pre_oi_14_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12584 ), .force_10(
        \shifter_0/n12585 ), .force_11(1'b0), .QN(n46527) );
  \**FFGEN**  \shifter_0/pre_oi_14_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12588 ), .force_10(
        \shifter_0/n12589 ), .force_11(1'b0), .QN(n46528) );
  \**FFGEN**  \shifter_0/pre_oi_14_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12592 ), .force_10(
        \shifter_0/n12593 ), .force_11(1'b0), .QN(n46529) );
  \**FFGEN**  \shifter_0/pre_oi_14_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12596 ), .force_10(
        \shifter_0/n12597 ), .force_11(1'b0), .QN(n46530) );
  \**FFGEN**  \shifter_0/pre_oi_14_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12600 ), .force_10(
        \shifter_0/n12601 ), .force_11(1'b0), .QN(n46531) );
  \**FFGEN**  \shifter_0/pre_oi_14_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12604 ), .force_10(
        \shifter_0/n12605 ), .force_11(1'b0), .QN(n46532) );
  \**FFGEN**  \shifter_0/pre_ow_14_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12608 ), .force_10(
        \shifter_0/n12609 ), .force_11(1'b0), .QN(n46833) );
  \**FFGEN**  \shifter_0/pre_ow_14_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12612 ), .force_10(
        \shifter_0/n12613 ), .force_11(1'b0), .QN(n46834) );
  \**FFGEN**  \shifter_0/pre_ow_14_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12616 ), .force_10(
        \shifter_0/n12617 ), .force_11(1'b0), .QN(n46835) );
  \**FFGEN**  \shifter_0/pre_ow_14_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12620 ), .force_10(
        \shifter_0/n12621 ), .force_11(1'b0), .QN(n46836) );
  \**FFGEN**  \shifter_0/pre_ow_14_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12624 ), .force_10(
        \shifter_0/n12625 ), .force_11(1'b0), .QN(n46837) );
  \**FFGEN**  \shifter_0/pre_ow_14_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12628 ), .force_10(
        \shifter_0/n12629 ), .force_11(1'b0), .QN(n46838) );
  \**FFGEN**  \shifter_0/pre_ow_14_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12632 ), .force_10(
        \shifter_0/n12633 ), .force_11(1'b0), .QN(n46839) );
  \**FFGEN**  \shifter_0/pre_ow_14_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12636 ), .force_10(
        \shifter_0/n12637 ), .force_11(1'b0), .QN(n46840) );
  \**FFGEN**  \shifter_0/pre_ow_14_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12640 ), .force_10(
        \shifter_0/n12641 ), .force_11(1'b0), .QN(n46841) );
  \**FFGEN**  \shifter_0/pre_ow_14_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12644 ), .force_10(
        \shifter_0/n12645 ), .force_11(1'b0), .QN(n46842) );
  \**FFGEN**  \shifter_0/pre_ow_14_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12648 ), .force_10(
        \shifter_0/n12649 ), .force_11(1'b0), .QN(n46843) );
  \**FFGEN**  \shifter_0/pre_ow_14_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12652 ), .force_10(
        \shifter_0/n12653 ), .force_11(1'b0), .QN(n46844) );
  \**FFGEN**  \shifter_0/pre_ow_14_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12656 ), .force_10(
        \shifter_0/n12657 ), .force_11(1'b0), .QN(n46845) );
  \**FFGEN**  \shifter_0/pre_ow_14_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12660 ), .force_10(
        \shifter_0/n12661 ), .force_11(1'b0), .QN(n46846) );
  \**FFGEN**  \shifter_0/pre_ow_14_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12664 ), .force_10(
        \shifter_0/n12665 ), .force_11(1'b0), .QN(n46847) );
  \**FFGEN**  \shifter_0/pre_ow_14_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12668 ), .force_10(
        \shifter_0/n12669 ), .force_11(1'b0), .QN(n46848) );
  \**FFGEN**  \shifter_0/pre_ow_14_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12672 ), .force_10(
        \shifter_0/n12673 ), .force_11(1'b0), .QN(n46849) );
  \**FFGEN**  \shifter_0/pre_ow_14_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12676 ), .force_10(
        \shifter_0/n12677 ), .force_11(1'b0), .QN(n46850) );
  \**FFGEN**  \shifter_0/pre_ow_14_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12680 ), .force_10(
        \shifter_0/n12681 ), .force_11(1'b0), .QN(n46851) );
  \**FFGEN**  \shifter_0/pre_ow_14_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12684 ), .force_10(
        \shifter_0/n12685 ), .force_11(1'b0), .QN(n46852) );
  \**FFGEN**  \shifter_0/pre_oi_15_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12688 ), .force_10(
        \shifter_0/n12689 ), .force_11(1'b0), .QN(n46533) );
  \**FFGEN**  \shifter_0/pre_oi_15_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12692 ), .force_10(
        \shifter_0/n12693 ), .force_11(1'b0), .QN(n46534) );
  \**FFGEN**  \shifter_0/pre_oi_15_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12696 ), .force_10(
        \shifter_0/n12697 ), .force_11(1'b0), .QN(n46535) );
  \**FFGEN**  \shifter_0/pre_oi_15_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12700 ), .force_10(
        \shifter_0/n12701 ), .force_11(1'b0), .QN(n46536) );
  \**FFGEN**  \shifter_0/pre_oi_15_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12704 ), .force_10(
        \shifter_0/n12705 ), .force_11(1'b0), .QN(n46537) );
  \**FFGEN**  \shifter_0/pre_oi_15_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12708 ), .force_10(
        \shifter_0/n12709 ), .force_11(1'b0), .QN(n46538) );
  \**FFGEN**  \shifter_0/pre_oi_15_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12712 ), .force_10(
        \shifter_0/n12713 ), .force_11(1'b0), .QN(n46539) );
  \**FFGEN**  \shifter_0/pre_oi_15_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12716 ), .force_10(
        \shifter_0/n12717 ), .force_11(1'b0), .QN(n46540) );
  \**FFGEN**  \shifter_0/pre_oi_15_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12720 ), .force_10(
        \shifter_0/n12721 ), .force_11(1'b0), .QN(n46541) );
  \**FFGEN**  \shifter_0/pre_oi_15_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12724 ), .force_10(
        \shifter_0/n12725 ), .force_11(1'b0), .QN(n46542) );
  \**FFGEN**  \shifter_0/pre_oi_15_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12728 ), .force_10(
        \shifter_0/n12729 ), .force_11(1'b0), .QN(n46543) );
  \**FFGEN**  \shifter_0/pre_oi_15_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12732 ), .force_10(
        \shifter_0/n12733 ), .force_11(1'b0), .QN(n46544) );
  \**FFGEN**  \shifter_0/pre_oi_15_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12736 ), .force_10(
        \shifter_0/n12737 ), .force_11(1'b0), .QN(n46545) );
  \**FFGEN**  \shifter_0/pre_oi_15_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12740 ), .force_10(
        \shifter_0/n12741 ), .force_11(1'b0), .QN(n46546) );
  \**FFGEN**  \shifter_0/pre_oi_15_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12744 ), .force_10(
        \shifter_0/n12745 ), .force_11(1'b0), .QN(n46547) );
  \**FFGEN**  \shifter_0/pre_oi_15_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12748 ), .force_10(
        \shifter_0/n12749 ), .force_11(1'b0), .QN(n46548) );
  \**FFGEN**  \shifter_0/pre_oi_15_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12752 ), .force_10(
        \shifter_0/n12753 ), .force_11(1'b0), .QN(n46549) );
  \**FFGEN**  \shifter_0/pre_oi_15_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12756 ), .force_10(
        \shifter_0/n12757 ), .force_11(1'b0), .QN(n46550) );
  \**FFGEN**  \shifter_0/pre_oi_15_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n12760 ), .force_10(
        \shifter_0/n12761 ), .force_11(1'b0), .QN(n46551) );
  \**FFGEN**  \shifter_0/pre_oi_15_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\shifter_0/n10204 ), .force_10(
        \shifter_0/n10205 ), .force_11(1'b0), .QN(n46552) );
  nand_x8_sg U15742 ( .A(n22417), .B(n22418), .X(n22396) );
  nand_x8_sg U15786 ( .A(n22442), .B(n22443), .X(n22421) );
  nand_x8_sg U15830 ( .A(n22467), .B(n22468), .X(n22446) );
  nand_x8_sg U15875 ( .A(n67499), .B(n22494), .X(n22473) );
  nand_x8_sg U15918 ( .A(n22467), .B(n22519), .X(n22498) );
  nand_x8_sg U15962 ( .A(n67499), .B(n22544), .X(n22523) );
  nor_x2_sg U16096 ( .A(n22624), .B(n57864), .X(n22623) );
  nor_x2_sg U16095 ( .A(n57298), .B(n57300), .X(n22624) );
  nor_x2_sg U16144 ( .A(n22651), .B(n57864), .X(n22650) );
  nor_x2_sg U16143 ( .A(n57304), .B(n57306), .X(n22651) );
  nand_x8_sg U16217 ( .A(n22693), .B(n22694), .X(n22653) );
  nand_x8_sg U16311 ( .A(n67181), .B(n22751), .X(n22654) );
  nand_x8_sg U16335 ( .A(n67180), .B(n22765), .X(n22656) );
  nand_x8_sg U16359 ( .A(n67179), .B(n22776), .X(n22658) );
  nand_x8_sg U16383 ( .A(n67178), .B(n22787), .X(n22660) );
  nand_x8_sg U16407 ( .A(n67177), .B(n22798), .X(n22662) );
  nand_x8_sg U16431 ( .A(n67176), .B(n22809), .X(n22664) );
  nand_x8_sg U16455 ( .A(n67175), .B(n22820), .X(n22666) );
  nand_x8_sg U16479 ( .A(n67174), .B(n22831), .X(n22668) );
  nand_x8_sg U16503 ( .A(n67173), .B(n22842), .X(n22670) );
  nand_x8_sg U16527 ( .A(n67172), .B(n22853), .X(n22672) );
  nand_x8_sg U16551 ( .A(n67171), .B(n22864), .X(n22674) );
  nand_x8_sg U16575 ( .A(n67170), .B(n22875), .X(n22676) );
  nand_x8_sg U16599 ( .A(n67169), .B(n22886), .X(n22678) );
  nand_x8_sg U16623 ( .A(n67168), .B(n22897), .X(n22680) );
  nand_x8_sg U16647 ( .A(n67167), .B(n22908), .X(n22682) );
  nand_x8_sg U16671 ( .A(n67166), .B(n22919), .X(n22684) );
  nand_x8_sg U16695 ( .A(n67165), .B(n22930), .X(n22686) );
  nand_x8_sg U16719 ( .A(n67164), .B(n22941), .X(n22688) );
  nand_x8_sg U16743 ( .A(n67163), .B(n22952), .X(n22690) );
  nand_x8_sg U16769 ( .A(n67162), .B(n22963), .X(n22692) );
  nand_x8_sg U16288 ( .A(n22740), .B(n22741), .X(n22700) );
  nand_x8_sg U16284 ( .A(n57302), .B(n22742), .X(n22741) );
  nand_x8_sg U16798 ( .A(n67394), .B(n22979), .X(n22701) );
  nand_x8_sg U16822 ( .A(n67393), .B(n22992), .X(n22703) );
  nand_x8_sg U16846 ( .A(n67392), .B(n23003), .X(n22705) );
  nand_x8_sg U16870 ( .A(n67391), .B(n23014), .X(n22707) );
  nand_x8_sg U16894 ( .A(n67390), .B(n23025), .X(n22709) );
  nand_x8_sg U16918 ( .A(n67389), .B(n23036), .X(n22711) );
  nand_x8_sg U16942 ( .A(n67388), .B(n23047), .X(n22713) );
  nand_x8_sg U16966 ( .A(n67387), .B(n23058), .X(n22715) );
  nand_x8_sg U16990 ( .A(n67386), .B(n23069), .X(n22717) );
  nand_x8_sg U17014 ( .A(n67385), .B(n23080), .X(n22719) );
  nand_x8_sg U17038 ( .A(n67384), .B(n23091), .X(n22721) );
  nand_x8_sg U17062 ( .A(n67383), .B(n23102), .X(n22723) );
  nand_x8_sg U17086 ( .A(n67382), .B(n23113), .X(n22725) );
  nand_x8_sg U17110 ( .A(n67381), .B(n23124), .X(n22727) );
  nand_x8_sg U17134 ( .A(n67380), .B(n23135), .X(n22729) );
  nand_x8_sg U17158 ( .A(n67379), .B(n23146), .X(n22731) );
  nand_x8_sg U17182 ( .A(n67378), .B(n23157), .X(n22733) );
  nand_x8_sg U17206 ( .A(n67377), .B(n23168), .X(n22735) );
  nand_x8_sg U17230 ( .A(n67376), .B(n23179), .X(n22737) );
  nand_x8_sg U17256 ( .A(n67375), .B(n23190), .X(n22739) );
  nor_x2_sg U16313 ( .A(n22759), .B(n57157), .X(n22750) );
  nand_x8_sg U16774 ( .A(n57097), .B(n22971), .X(n22761) );
  nand_x8_sg U16773 ( .A(n68588), .B(n22972), .X(n22971) );
  nor_x2_sg U16337 ( .A(n22772), .B(n57157), .X(n22764) );
  nor_x2_sg U16361 ( .A(n22783), .B(n57157), .X(n22775) );
  nor_x2_sg U16385 ( .A(n22794), .B(n57157), .X(n22786) );
  nor_x2_sg U16409 ( .A(n22805), .B(n57157), .X(n22797) );
  nor_x2_sg U16433 ( .A(n22816), .B(n57157), .X(n22808) );
  nor_x2_sg U16457 ( .A(n22827), .B(n57157), .X(n22819) );
  nor_x2_sg U16481 ( .A(n22838), .B(n57157), .X(n22830) );
  nor_x2_sg U16505 ( .A(n22849), .B(n57157), .X(n22841) );
  nor_x2_sg U16529 ( .A(n22860), .B(n57157), .X(n22852) );
  nor_x2_sg U16553 ( .A(n22871), .B(n57157), .X(n22863) );
  nor_x2_sg U16577 ( .A(n22882), .B(n57157), .X(n22874) );
  nor_x2_sg U16601 ( .A(n22893), .B(n57157), .X(n22885) );
  nor_x2_sg U16625 ( .A(n22904), .B(n57157), .X(n22896) );
  nor_x2_sg U16649 ( .A(n22915), .B(n57157), .X(n22907) );
  nor_x2_sg U16673 ( .A(n22926), .B(n57157), .X(n22918) );
  nor_x2_sg U16697 ( .A(n22937), .B(n57157), .X(n22929) );
  nor_x2_sg U16721 ( .A(n22948), .B(n57157), .X(n22940) );
  nor_x2_sg U16800 ( .A(n22986), .B(n57151), .X(n22978) );
  nand_x8_sg U17282 ( .A(n57302), .B(n23198), .X(n22988) );
  nand_x8_sg U17281 ( .A(n68588), .B(n23199), .X(n23198) );
  nor_x2_sg U16824 ( .A(n22999), .B(n57151), .X(n22991) );
  nor_x2_sg U16848 ( .A(n23010), .B(n57151), .X(n23002) );
  nor_x2_sg U16872 ( .A(n23021), .B(n57151), .X(n23013) );
  nor_x2_sg U16896 ( .A(n23032), .B(n57151), .X(n23024) );
  nor_x2_sg U16920 ( .A(n23043), .B(n57151), .X(n23035) );
  nor_x2_sg U16944 ( .A(n23054), .B(n57151), .X(n23046) );
  nor_x2_sg U16968 ( .A(n23065), .B(n57151), .X(n23057) );
  nor_x2_sg U16992 ( .A(n23076), .B(n57151), .X(n23068) );
  nor_x2_sg U17016 ( .A(n23087), .B(n57151), .X(n23079) );
  nor_x2_sg U17040 ( .A(n23098), .B(n57151), .X(n23090) );
  nor_x2_sg U17064 ( .A(n23109), .B(n57151), .X(n23101) );
  nor_x2_sg U17088 ( .A(n23120), .B(n57151), .X(n23112) );
  nor_x2_sg U17112 ( .A(n23131), .B(n57151), .X(n23123) );
  nor_x2_sg U17136 ( .A(n23142), .B(n57151), .X(n23134) );
  nor_x2_sg U17160 ( .A(n23153), .B(n57151), .X(n23145) );
  nor_x2_sg U17184 ( .A(n23164), .B(n57151), .X(n23156) );
  nor_x2_sg U17208 ( .A(n23175), .B(n57151), .X(n23167) );
  nand_x8_sg U18336 ( .A(n57298), .B(n68576), .X(n23543) );
  nand_x8_sg U18487 ( .A(n57304), .B(n68397), .X(n23675) );
  nand_x8_sg U17730 ( .A(n23539), .B(n23540), .X(n23422) );
  nand_x8_sg U17723 ( .A(n23541), .B(n23542), .X(n23540) );
  nor_x2_sg U17721 ( .A(n57300), .B(n57918), .X(n23542) );
  nand_x8_sg U17882 ( .A(n23671), .B(n23672), .X(n23556) );
  nand_x8_sg U17874 ( .A(n23673), .B(n23674), .X(n23672) );
  nor_x2_sg U17872 ( .A(n57306), .B(n57918), .X(n23674) );
  nand_x8_sg U18035 ( .A(n23802), .B(n23803), .X(n23686) );
  nand_x8_sg U18034 ( .A(n23809), .B(n57917), .X(n23802) );
  nand_x8_sg U18031 ( .A(n23804), .B(n23805), .X(n23803) );
  nand_x8_sg U18187 ( .A(n23931), .B(n23932), .X(n23816) );
  nand_x8_sg U18186 ( .A(n23938), .B(n57917), .X(n23931) );
  nand_x8_sg U18183 ( .A(n23933), .B(n23934), .X(n23932) );
  nand_x8_sg U18621 ( .A(n24259), .B(n24260), .X(n24163) );
  nand_x8_sg U18620 ( .A(n57918), .B(n24262), .X(n24259) );
  nand_x8_sg U18754 ( .A(n24368), .B(n24369), .X(n24272) );
  nand_x8_sg U18887 ( .A(n24477), .B(n24478), .X(n24381) );
  nand_x8_sg U18886 ( .A(n57918), .B(n24480), .X(n24477) );
  nand_x8_sg U18876 ( .A(n24479), .B(n57920), .X(n24478) );
  nand_x8_sg U19020 ( .A(n24589), .B(n24590), .X(n24493) );
  nand_x8_sg U19019 ( .A(n57918), .B(n24592), .X(n24589) );
  nand_x8_sg U19009 ( .A(n24591), .B(n57917), .X(n24590) );
  nand_x8_sg U19155 ( .A(n24683), .B(n24684), .X(n24605) );
  nand_x8_sg U19154 ( .A(n57918), .B(n24685), .X(n24683) );
  nand_x8_sg U19142 ( .A(n67101), .B(n57920), .X(n24684) );
  nand_x8_sg U19291 ( .A(n24777), .B(n24778), .X(n24700) );
  nand_x8_sg U19290 ( .A(n57919), .B(n24779), .X(n24777) );
  nand_x8_sg U19277 ( .A(n67523), .B(n57920), .X(n24778) );
  nor_x2_sg U19338 ( .A(n24829), .B(n67305), .X(n24827) );
  nor_x2_sg U19383 ( .A(n24829), .B(n67304), .X(n24858) );
  nor_x2_sg U19428 ( .A(n24829), .B(n67303), .X(n24888) );
  nor_x2_sg U19563 ( .A(n24829), .B(n67302), .X(n24978) );
  nor_x2_sg U19608 ( .A(n24829), .B(n67301), .X(n25008) );
  nor_x2_sg U19653 ( .A(n24829), .B(n67300), .X(n25038) );
  nor_x2_sg U19788 ( .A(n24829), .B(n67299), .X(n25128) );
  nor_x2_sg U19833 ( .A(n24829), .B(n67298), .X(n25158) );
  nor_x2_sg U19968 ( .A(n24829), .B(n67297), .X(n25248) );
  nor_x2_sg U20013 ( .A(n24829), .B(n67296), .X(n25278) );
  nor_x2_sg U20058 ( .A(n24829), .B(n67295), .X(n25308) );
  nor_x2_sg U20200 ( .A(n24829), .B(n67294), .X(n25399) );
  nor_x2_sg U20245 ( .A(n24829), .B(n67498), .X(n25430) );
  nor_x2_sg U20290 ( .A(n24829), .B(n67497), .X(n25460) );
  nor_x2_sg U20335 ( .A(n24829), .B(n67496), .X(n25490) );
  nor_x2_sg U20470 ( .A(n24829), .B(n67495), .X(n25580) );
  nor_x2_sg U20515 ( .A(n24829), .B(n67494), .X(n25610) );
  nor_x2_sg U20560 ( .A(n24829), .B(n67493), .X(n25640) );
  nor_x2_sg U20695 ( .A(n24829), .B(n67492), .X(n25730) );
  nor_x2_sg U20740 ( .A(n24829), .B(n67491), .X(n25760) );
  nor_x2_sg U20875 ( .A(n24829), .B(n67490), .X(n25850) );
  nor_x2_sg U20920 ( .A(n24829), .B(n67489), .X(n25880) );
  nor_x2_sg U20965 ( .A(n24829), .B(n67488), .X(n25910) );
  nor_x2_sg U21129 ( .A(n24829), .B(n67487), .X(n26001) );
  nand_x8_sg U21271 ( .A(n34174), .B(n26010), .X(n26249) );
  nand_x8_sg U23181 ( .A(n57114), .B(n34222), .X(n26034) );
  nand_x8_sg U23449 ( .A(n26261), .B(n26262), .X(n34222) );
  nor_x2_sg U23445 ( .A(n26317), .B(n57310), .X(n26306) );
  nor_x2_sg U23444 ( .A(n26318), .B(n26319), .X(n26317) );
  nor_x2_sg U23433 ( .A(n67572), .B(n26330), .X(n26328) );
  nor_x2_sg U23430 ( .A(n26052), .B(n67571), .X(n26329) );
  nand_x8_sg U23530 ( .A(n57109), .B(n57308), .X(n26047) );
  nand_x8_sg U23538 ( .A(n57106), .B(n57308), .X(n26051) );
  nor_x2_sg U23401 ( .A(n57310), .B(n26281), .X(n26270) );
  nor_x2_sg U23400 ( .A(n26282), .B(n26283), .X(n26281) );
  nor_x2_sg U23397 ( .A(n26114), .B(n67567), .X(n26295) );
  nand_x8_sg U23523 ( .A(n57107), .B(n57308), .X(n26114) );
  nor_x2_sg U23391 ( .A(n26289), .B(n26290), .X(n26288) );
  nand_x8_sg U21332 ( .A(n34174), .B(n26012), .X(n26250) );
  nand_x8_sg U21393 ( .A(n34174), .B(n26014), .X(n26251) );
  nand_x8_sg U21455 ( .A(n34174), .B(n26008), .X(n26252) );
  nand_x8_sg U21516 ( .A(n33738), .B(n26010), .X(n26253) );
  nand_x8_sg U21577 ( .A(n33738), .B(n26012), .X(n26254) );
  nand_x8_sg U21638 ( .A(n33738), .B(n26014), .X(n26255) );
  nand_x8_sg U21699 ( .A(n33738), .B(n26008), .X(n26256) );
  nand_x8_sg U21760 ( .A(n26010), .B(n33868), .X(n26257) );
  nand_x8_sg U21821 ( .A(n26012), .B(n33868), .X(n26259) );
  nand_x8_sg U21882 ( .A(n26014), .B(n33868), .X(n26006) );
  nand_x8_sg U21944 ( .A(n26008), .B(n33868), .X(n26007) );
  nand_x8_sg U22007 ( .A(n26010), .B(n33266), .X(n26009) );
  nand_x8_sg U22070 ( .A(n26012), .B(n33266), .X(n26011) );
  nand_x8_sg U22133 ( .A(n26014), .B(n33266), .X(n26013) );
  nand_x8_sg U22196 ( .A(n26008), .B(n33266), .X(n26015) );
  nand_x8_sg U22257 ( .A(n33998), .B(n26017), .X(n26016) );
  nand_x8_sg U22318 ( .A(n26019), .B(n33998), .X(n26018) );
  nand_x8_sg U22379 ( .A(n26021), .B(n33998), .X(n26020) );
  nand_x8_sg U22441 ( .A(n26023), .B(n33998), .X(n26022) );
  nand_x8_sg U22502 ( .A(n34219), .B(n26017), .X(n26024) );
  nand_x8_sg U22563 ( .A(n34219), .B(n26019), .X(n26025) );
  nand_x8_sg U22624 ( .A(n34219), .B(n26021), .X(n26026) );
  nand_x8_sg U22685 ( .A(n34219), .B(n26023), .X(n26027) );
  nand_x8_sg U22746 ( .A(n34086), .B(n26017), .X(n26028) );
  nand_x8_sg U22807 ( .A(n34086), .B(n26019), .X(n26029) );
  nand_x8_sg U22868 ( .A(n34086), .B(n26021), .X(n26030) );
  nand_x8_sg U22930 ( .A(n34086), .B(n26023), .X(n26031) );
  nand_x8_sg U22993 ( .A(n26017), .B(n34131), .X(n26032) );
  nand_x8_sg U23056 ( .A(n26019), .B(n34131), .X(n26035) );
  nand_x8_sg U23119 ( .A(n26021), .B(n34131), .X(n26037) );
  nand_x8_sg U23183 ( .A(n26023), .B(n34131), .X(n26038) );
  nor_x2_sg U23318 ( .A(n26124), .B(n26125), .X(n26123) );
  nor_x2_sg U23307 ( .A(n57310), .B(n26136), .X(n26135) );
  nor_x2_sg U23306 ( .A(n26137), .B(n26138), .X(n26136) );
  nor_x2_sg U23303 ( .A(n26114), .B(n67562), .X(n26150) );
  nor_x2_sg U23297 ( .A(n26144), .B(n26145), .X(n26143) );
  nor_x2_sg U23277 ( .A(n26081), .B(n26082), .X(n26080) );
  nor_x2_sg U23266 ( .A(n57310), .B(n26097), .X(n26096) );
  nor_x2_sg U23265 ( .A(n26098), .B(n26099), .X(n26097) );
  nor_x2_sg U23262 ( .A(n26114), .B(n67556), .X(n26111) );
  nor_x2_sg U23256 ( .A(n26105), .B(n26106), .X(n26104) );
  nor_x2_sg U23554 ( .A(n26216), .B(n26217), .X(n26215) );
  nor_x2_sg U23528 ( .A(n57310), .B(n26228), .X(n26227) );
  nor_x2_sg U23527 ( .A(n26229), .B(n26230), .X(n26228) );
  nor_x2_sg U23524 ( .A(n26114), .B(n67550), .X(n26242) );
  nor_x2_sg U23514 ( .A(n26236), .B(n26237), .X(n26235) );
  nor_x2_sg U23491 ( .A(n26182), .B(n26183), .X(n26181) );
  nor_x2_sg U23480 ( .A(n57310), .B(n26194), .X(n26193) );
  nor_x2_sg U23479 ( .A(n26195), .B(n26196), .X(n26194) );
  nor_x2_sg U23476 ( .A(n26114), .B(n67544), .X(n26208) );
  nor_x2_sg U23470 ( .A(n26202), .B(n26203), .X(n26201) );
  inv_x4_sg U39564 ( .A(n57914), .X(n57913) );
  inv_x2_sg U39565 ( .A(n57915), .X(n57914) );
  inv_x4_sg U39566 ( .A(n57881), .X(n57869) );
  inv_x4_sg U39567 ( .A(n57881), .X(n57879) );
  inv_x4_sg U39568 ( .A(n57853), .X(n57852) );
  inv_x2_sg U39569 ( .A(n34232), .X(n57853) );
  inv_x2_sg U39570 ( .A(n51555), .X(n57723) );
  nor_x1_sg U39571 ( .A(n30624), .B(n57882), .X(n29327) );
  inv_x8_sg U39572 ( .A(n57772), .X(n46196) );
  inv_x8_sg U39573 ( .A(n46196), .X(n46197) );
  inv_x8_sg U39574 ( .A(n46196), .X(n46198) );
  inv_x8_sg U39575 ( .A(n57763), .X(n46199) );
  inv_x8_sg U39576 ( .A(n46199), .X(n46200) );
  inv_x8_sg U39577 ( .A(n46199), .X(n46201) );
  inv_x8_sg U39578 ( .A(n57852), .X(n46202) );
  inv_x4_sg U39579 ( .A(n46202), .X(n46203) );
  inv_x8_sg U39580 ( .A(n46202), .X(n46204) );
  inv_x8_sg U39581 ( .A(n57913), .X(n46205) );
  inv_x4_sg U39582 ( .A(n46205), .X(n46206) );
  inv_x8_sg U39583 ( .A(n46205), .X(n46207) );
  inv_x8_sg U39584 ( .A(n57869), .X(n46208) );
  inv_x8_sg U39585 ( .A(n46208), .X(n46209) );
  inv_x8_sg U39586 ( .A(n46208), .X(n46210) );
  inv_x8_sg U39587 ( .A(n57879), .X(n46211) );
  inv_x8_sg U39588 ( .A(n46211), .X(n46212) );
  inv_x8_sg U39589 ( .A(n46211), .X(n46213) );
  inv_x2_sg U39590 ( .A(n29327), .X(n57916) );
  inv_x2_sg U39591 ( .A(n57949), .X(n57947) );
  inv_x4_sg U39592 ( .A(n57884), .X(n57883) );
  inv_x2_sg U39593 ( .A(n29328), .X(n57885) );
  inv_x4_sg U39594 ( .A(n38414), .X(n57633) );
  inv_x4_sg U39595 ( .A(n57916), .X(n57915) );
  inv_x4_sg U39596 ( .A(n57845), .X(n57829) );
  inv_x2_sg U39597 ( .A(n57721), .X(n57714) );
  inv_x4_sg U39598 ( .A(n57723), .X(n57722) );
  nor_x1_sg U39599 ( .A(n57917), .B(n57296), .X(n61903) );
  nor_x1_sg U39600 ( .A(n68227), .B(n57714), .X(n35847) );
  inv_x2_sg U39601 ( .A(n61903), .X(n57458) );
  nand_x2_sg U39602 ( .A(n57348), .B(n57457), .X(n67084) );
  nor_x2_sg U39603 ( .A(n57917), .B(n57100), .X(n61904) );
  inv_x4_sg U39604 ( .A(n57777), .X(n57776) );
  inv_x2_sg U39605 ( .A(n57778), .X(n57777) );
  inv_x1_sg U39606 ( .A(n35847), .X(n57778) );
  inv_x2_sg U39607 ( .A(n29329), .X(n57868) );
  inv_x1_sg U39608 ( .A(n47523), .X(n47388) );
  inv_x1_sg U39609 ( .A(n51259), .X(n47386) );
  inv_x1_sg U39610 ( .A(n47525), .X(n47303) );
  inv_x1_sg U39611 ( .A(n56813), .X(n47384) );
  inv_x1_sg U39612 ( .A(n51367), .X(n47324) );
  inv_x1_sg U39613 ( .A(n51307), .X(n47301) );
  inv_x1_sg U39614 ( .A(n47555), .X(n47322) );
  inv_x1_sg U39615 ( .A(n47539), .X(n47382) );
  inv_x1_sg U39616 ( .A(n56793), .X(n47380) );
  inv_x1_sg U39617 ( .A(n51345), .X(n47320) );
  inv_x1_sg U39618 ( .A(n56745), .X(n47307) );
  inv_x1_sg U39619 ( .A(n51281), .X(n47290) );
  inv_x1_sg U39620 ( .A(n51415), .X(n47378) );
  inv_x1_sg U39621 ( .A(n47553), .X(n47376) );
  inv_x1_sg U39622 ( .A(n56851), .X(n47326) );
  inv_x1_sg U39623 ( .A(n51321), .X(n47305) );
  nand_x2_sg U39624 ( .A(n24234), .B(n25239), .X(n25238) );
  nand_x2_sg U39625 ( .A(n24239), .B(n25269), .X(n25268) );
  nand_x2_sg U39626 ( .A(n24328), .B(n25751), .X(n25750) );
  nand_x2_sg U39627 ( .A(n24376), .B(n25992), .X(n25991) );
  inv_x2_sg U39628 ( .A(n32353), .X(n47334) );
  nor_x1_sg U39629 ( .A(n68576), .B(n32354), .X(n32353) );
  inv_x2_sg U39630 ( .A(n35552), .X(n47296) );
  nor_x1_sg U39631 ( .A(n68370), .B(n35705), .X(n35552) );
  nand_x2_sg U39632 ( .A(n68272), .B(output_taken), .X(n39838) );
  inv_x2_sg U39633 ( .A(n22567), .X(n57512) );
  nand_x1_sg U39634 ( .A(n22568), .B(n22569), .X(n22567) );
  inv_x2_sg U39635 ( .A(n22593), .X(n57518) );
  nand_x1_sg U39636 ( .A(n22594), .B(n22595), .X(n22593) );
  inv_x2_sg U39637 ( .A(n22618), .X(n57509) );
  nand_x1_sg U39638 ( .A(n22619), .B(n22620), .X(n22618) );
  inv_x2_sg U39639 ( .A(n22645), .X(n57515) );
  nand_x1_sg U39640 ( .A(n22646), .B(n22647), .X(n22645) );
  nor_x2_sg U39641 ( .A(n57159), .B(n61902), .X(n22760) );
  nor_x2_sg U39642 ( .A(n57153), .B(n61902), .X(n22987) );
  nand_x2_sg U39643 ( .A(n47437), .B(n68387), .X(n34223) );
  inv_x2_sg U39644 ( .A(n53712), .X(n53713) );
  inv_x1_sg U39645 ( .A(\shifter_0/w_pointer [2]), .X(n53712) );
  inv_x2_sg U39646 ( .A(n51054), .X(n51055) );
  inv_x1_sg U39647 ( .A(\shifter_0/i_pointer [3]), .X(n51054) );
  inv_x2_sg U39648 ( .A(n32798), .X(n47330) );
  nor_x1_sg U39649 ( .A(n68397), .B(n32799), .X(n32798) );
  nand_x2_sg U39650 ( .A(n40227), .B(n61908), .X(n32831) );
  inv_x2_sg U39651 ( .A(n47314), .X(n47315) );
  inv_x1_sg U39652 ( .A(\filter_0/N15 ), .X(n47314) );
  inv_x2_sg U39653 ( .A(n32920), .X(n47294) );
  nor_x1_sg U39654 ( .A(n32921), .B(n68376), .X(n32920) );
  inv_x2_sg U39655 ( .A(n32875), .X(n47311) );
  nor_x1_sg U39656 ( .A(n32876), .B(n68381), .X(n32875) );
  inv_x2_sg U39657 ( .A(n35514), .X(n57794) );
  nor_x1_sg U39658 ( .A(n35705), .B(n57786), .X(n35514) );
  nor_x2_sg U39659 ( .A(n39838), .B(n68271), .X(n39837) );
  inv_x2_sg U39660 ( .A(n38410), .X(n47298) );
  nor_x1_sg U39661 ( .A(n38416), .B(n68272), .X(n38410) );
  inv_x4_sg U39662 ( .A(n57393), .X(n57389) );
  inv_x4_sg U39663 ( .A(n57392), .X(n57391) );
  inv_x4_sg U39664 ( .A(n47505), .X(n57921) );
  inv_x4_sg U39665 ( .A(n57794), .X(n57793) );
  inv_x4_sg U39666 ( .A(n57324), .X(n57323) );
  inv_x4_sg U39667 ( .A(n57458), .X(n57457) );
  inv_x4_sg U39668 ( .A(n29332), .X(n57863) );
  inv_x4_sg U39669 ( .A(n57347), .X(n57346) );
  inv_x1_sg U39670 ( .A(n58656), .X(n58481) );
  inv_x4_sg U39671 ( .A(n57482), .X(n57481) );
  inv_x4_sg U39672 ( .A(n58387), .X(n57319) );
  inv_x4_sg U39673 ( .A(n58388), .X(n57321) );
  inv_x4_sg U39674 ( .A(n58376), .X(n57317) );
  inv_x4_sg U39675 ( .A(n57784), .X(n57783) );
  inv_x4_sg U39676 ( .A(n57515), .X(n57514) );
  inv_x4_sg U39677 ( .A(n57512), .X(n57511) );
  inv_x4_sg U39678 ( .A(n57509), .X(n57508) );
  inv_x4_sg U39679 ( .A(n57518), .X(n57517) );
  inv_x4_sg U39680 ( .A(n57474), .X(n57473) );
  inv_x4_sg U39681 ( .A(n57466), .X(n57465) );
  inv_x4_sg U39682 ( .A(n57490), .X(n57489) );
  inv_x4_sg U39683 ( .A(n57486), .X(n57485) );
  inv_x4_sg U39684 ( .A(n57494), .X(n57493) );
  inv_x4_sg U39685 ( .A(n57501), .X(n57500) );
  inv_x4_sg U39686 ( .A(n57504), .X(n57503) );
  inv_x4_sg U39687 ( .A(n57470), .X(n57469) );
  inv_x4_sg U39688 ( .A(n57478), .X(n57477) );
  inv_x4_sg U39689 ( .A(n57498), .X(n57497) );
  inv_x4_sg U39690 ( .A(n58374), .X(n57315) );
  inv_x4_sg U39691 ( .A(n57313), .X(n57312) );
  inv_x4_sg U39692 ( .A(n47297), .X(n57787) );
  inv_x4_sg U39693 ( .A(n24829), .X(n57506) );
  inv_x4_sg U39694 ( .A(n67084), .X(n57101) );
  inv_x4_sg U39695 ( .A(n32831), .X(n57167) );
  inv_x4_sg U39696 ( .A(n32880), .X(n57287) );
  inv_x4_sg U39697 ( .A(n34223), .X(n57112) );
  inv_x4_sg U39698 ( .A(n33182), .X(n57259) );
  inv_x4_sg U39699 ( .A(n33011), .X(n57275) );
  inv_x4_sg U39700 ( .A(n33139), .X(n57263) );
  inv_x4_sg U39701 ( .A(n32968), .X(n57279) );
  inv_x4_sg U39702 ( .A(n33097), .X(n57267) );
  inv_x4_sg U39703 ( .A(n32925), .X(n57283) );
  inv_x4_sg U39704 ( .A(n33054), .X(n57271) );
  inv_x4_sg U39705 ( .A(n32881), .X(n57285) );
  inv_x4_sg U39706 ( .A(n32834), .X(n57291) );
  inv_x4_sg U39707 ( .A(n32835), .X(n57289) );
  inv_x4_sg U39708 ( .A(n57559), .X(n57555) );
  inv_x4_sg U39709 ( .A(n24829), .X(n57505) );
  inv_x4_sg U39710 ( .A(n57462), .X(n57461) );
  inv_x4_sg U39711 ( .A(n34180), .X(n57171) );
  inv_x4_sg U39712 ( .A(n33872), .X(n57198) );
  inv_x4_sg U39713 ( .A(n34135), .X(n57175) );
  inv_x4_sg U39714 ( .A(n34047), .X(n57182) );
  inv_x4_sg U39715 ( .A(n33871), .X(n57200) );
  inv_x4_sg U39716 ( .A(n34002), .X(n57186) );
  inv_x4_sg U39717 ( .A(n33742), .X(n57208) );
  inv_x4_sg U39718 ( .A(n33741), .X(n57210) );
  inv_x4_sg U39719 ( .A(n34179), .X(n57173) );
  inv_x4_sg U39720 ( .A(n34134), .X(n57177) );
  inv_x4_sg U39721 ( .A(n34046), .X(n57184) );
  inv_x4_sg U39722 ( .A(n33527), .X(n57228) );
  inv_x4_sg U39723 ( .A(n33786), .X(n57206) );
  inv_x4_sg U39724 ( .A(n33828), .X(n57203) );
  inv_x4_sg U39725 ( .A(n34001), .X(n57188) );
  inv_x4_sg U39726 ( .A(n33569), .X(n57225) );
  inv_x4_sg U39727 ( .A(n33484), .X(n57231) );
  inv_x4_sg U39728 ( .A(n34091), .X(n57180) );
  nand_x4_sg U39729 ( .A(n57170), .B(n34222), .X(n32874) );
  inv_x4_sg U39730 ( .A(n33400), .X(n57239) );
  inv_x4_sg U39731 ( .A(n33269), .X(n57251) );
  inv_x4_sg U39732 ( .A(n33225), .X(n57255) );
  inv_x4_sg U39733 ( .A(n33656), .X(n57218) );
  inv_x4_sg U39734 ( .A(n33698), .X(n57214) );
  inv_x4_sg U39735 ( .A(n33958), .X(n57192) );
  inv_x4_sg U39736 ( .A(n33915), .X(n57196) );
  inv_x4_sg U39737 ( .A(n33442), .X(n57235) );
  inv_x4_sg U39738 ( .A(n33355), .X(n57243) );
  inv_x4_sg U39739 ( .A(n33313), .X(n57247) );
  inv_x4_sg U39740 ( .A(n33612), .X(n57222) );
  inv_x4_sg U39741 ( .A(n53715), .X(n57295) );
  inv_x4_sg U39742 ( .A(n56950), .X(n56951) );
  inv_x4_sg U39743 ( .A(n56938), .X(n56939) );
  inv_x4_sg U39744 ( .A(n56942), .X(n56943) );
  inv_x4_sg U39745 ( .A(n56946), .X(n56947) );
  inv_x4_sg U39746 ( .A(n56966), .X(n56967) );
  inv_x4_sg U39747 ( .A(n56954), .X(n56955) );
  inv_x4_sg U39748 ( .A(n56958), .X(n56959) );
  inv_x4_sg U39749 ( .A(n56962), .X(n56963) );
  inv_x2_sg U39750 ( .A(n35708), .X(n57785) );
  inv_x4_sg U39751 ( .A(n32803), .X(n57169) );
  inv_x4_sg U39752 ( .A(n22987), .X(n57150) );
  inv_x4_sg U39753 ( .A(n22760), .X(n57156) );
  inv_x4_sg U39754 ( .A(n57867), .X(n57866) );
  inv_x4_sg U39755 ( .A(n61904), .X(n57462) );
  inv_x4_sg U39756 ( .A(n29333), .X(n57861) );
  inv_x4_sg U39757 ( .A(n26091), .X(n57108) );
  inv_x4_sg U39758 ( .A(n26092), .X(n57105) );
  inv_x4_sg U39759 ( .A(n26095), .X(n57110) );
  inv_x4_sg U39760 ( .A(n58644), .X(n57098) );
  inv_x4_sg U39761 ( .A(n47315), .X(n57309) );
  inv_x4_sg U39762 ( .A(n56964), .X(n56965) );
  inv_x4_sg U39763 ( .A(n56948), .X(n56949) );
  inv_x4_sg U39764 ( .A(n56952), .X(n56953) );
  inv_x4_sg U39765 ( .A(n56956), .X(n56957) );
  inv_x4_sg U39766 ( .A(n56960), .X(n56961) );
  inv_x4_sg U39767 ( .A(n56936), .X(n56937) );
  inv_x4_sg U39768 ( .A(n56940), .X(n56941) );
  inv_x4_sg U39769 ( .A(n56944), .X(n56945) );
  inv_x4_sg U39770 ( .A(n57785), .X(n57784) );
  inv_x4_sg U39771 ( .A(n47415), .X(n57299) );
  inv_x4_sg U39772 ( .A(n32802), .X(n57293) );
  inv_x4_sg U39773 ( .A(n47413), .X(n57305) );
  inv_x4_sg U39774 ( .A(n56928), .X(n56929) );
  inv_x4_sg U39775 ( .A(n51055), .X(n57301) );
  inv_x4_sg U39776 ( .A(n53713), .X(n57297) );
  inv_x2_sg U39777 ( .A(n22467), .X(n67097) );
  inv_x2_sg U39778 ( .A(n23946), .X(n57487) );
  inv_x2_sg U39779 ( .A(n24056), .X(n57495) );
  inv_x2_sg U39780 ( .A(n23205), .X(n57471) );
  inv_x2_sg U39781 ( .A(n23313), .X(n57479) );
  inv_x2_sg U39782 ( .A(n23204), .X(n57467) );
  inv_x2_sg U39783 ( .A(n23944), .X(n57483) );
  inv_x2_sg U39784 ( .A(n24054), .X(n57491) );
  inv_x2_sg U39785 ( .A(n23312), .X(n57475) );
  inv_x4_sg U39786 ( .A(n47364), .X(n47365) );
  inv_x4_sg U39787 ( .A(n47366), .X(n47367) );
  inv_x4_sg U39788 ( .A(n56922), .X(n56923) );
  inv_x4_sg U39789 ( .A(n47368), .X(n47369) );
  inv_x4_sg U39790 ( .A(n47428), .X(n47429) );
  inv_x4_sg U39791 ( .A(n56924), .X(n56925) );
  inv_x4_sg U39792 ( .A(n47430), .X(n47431) );
  inv_x4_sg U39793 ( .A(n56926), .X(n56927) );
  inv_x4_sg U39794 ( .A(n47370), .X(n47371) );
  inv_x4_sg U39795 ( .A(n47432), .X(n47433) );
  inv_x4_sg U39796 ( .A(n56932), .X(n56933) );
  inv_x4_sg U39797 ( .A(n47434), .X(n47435) );
  inv_x4_sg U39798 ( .A(n47356), .X(n47357) );
  inv_x4_sg U39799 ( .A(n47358), .X(n47359) );
  inv_x4_sg U39800 ( .A(n56916), .X(n56917) );
  inv_x4_sg U39801 ( .A(n47360), .X(n47361) );
  inv_x4_sg U39802 ( .A(n47420), .X(n47421) );
  inv_x4_sg U39803 ( .A(n56918), .X(n56919) );
  inv_x4_sg U39804 ( .A(n47422), .X(n47423) );
  inv_x4_sg U39805 ( .A(n56920), .X(n56921) );
  inv_x4_sg U39806 ( .A(n47362), .X(n47363) );
  inv_x4_sg U39807 ( .A(n47424), .X(n47425) );
  inv_x4_sg U39808 ( .A(n56930), .X(n56931) );
  inv_x4_sg U39809 ( .A(n47426), .X(n47427) );
  inv_x1_sg U39810 ( .A(n30626), .X(n46854) );
  inv_x2_sg U39811 ( .A(n46854), .X(n46855) );
  inv_x1_sg U39812 ( .A(n31972), .X(n46856) );
  inv_x2_sg U39813 ( .A(n46856), .X(n46857) );
  inv_x1_sg U39814 ( .A(n31986), .X(n46858) );
  inv_x2_sg U39815 ( .A(n46858), .X(n46859) );
  inv_x1_sg U39816 ( .A(n31985), .X(n46860) );
  inv_x2_sg U39817 ( .A(n46860), .X(n46861) );
  inv_x1_sg U39818 ( .A(n32508), .X(n46862) );
  inv_x2_sg U39819 ( .A(n46862), .X(n46863) );
  inv_x1_sg U39820 ( .A(n32507), .X(n46864) );
  inv_x2_sg U39821 ( .A(n46864), .X(n46865) );
  inv_x1_sg U39822 ( .A(n32385), .X(n46866) );
  inv_x2_sg U39823 ( .A(n46866), .X(n46867) );
  inv_x1_sg U39824 ( .A(n32384), .X(n46868) );
  inv_x2_sg U39825 ( .A(n46868), .X(n46869) );
  inv_x1_sg U39826 ( .A(n31983), .X(n46870) );
  inv_x2_sg U39827 ( .A(n46870), .X(n46871) );
  nor_x2_sg U39828 ( .A(n23530), .B(n24470), .X(n24469) );
  nor_x2_sg U39829 ( .A(n23536), .B(n24475), .X(n24474) );
  nand_x2_sg U39830 ( .A(n67396), .B(n57126), .X(n24588) );
  nand_x2_sg U39831 ( .A(n67396), .B(n57115), .X(n25974) );
  nand_x2_sg U39832 ( .A(n67223), .B(n57117), .X(n25072) );
  nand_x2_sg U39833 ( .A(n67221), .B(n57117), .X(n25102) );
  nand_x2_sg U39834 ( .A(n67219), .B(n57117), .X(n25132) );
  nand_x2_sg U39835 ( .A(n67410), .B(n57115), .X(n25764) );
  inv_x1_sg U39836 ( .A(n31977), .X(n46872) );
  inv_x2_sg U39837 ( .A(n46872), .X(n46873) );
  inv_x1_sg U39838 ( .A(n31976), .X(n46874) );
  inv_x2_sg U39839 ( .A(n46874), .X(n46875) );
  inv_x1_sg U39840 ( .A(n32062), .X(n46876) );
  inv_x2_sg U39841 ( .A(n46876), .X(n46877) );
  inv_x1_sg U39842 ( .A(n32061), .X(n46878) );
  inv_x2_sg U39843 ( .A(n46878), .X(n46879) );
  inv_x1_sg U39844 ( .A(n32376), .X(n46880) );
  inv_x2_sg U39845 ( .A(n46880), .X(n46881) );
  inv_x1_sg U39846 ( .A(n32375), .X(n46882) );
  inv_x2_sg U39847 ( .A(n46882), .X(n46883) );
  nor_x2_sg U39848 ( .A(n23530), .B(n24677), .X(n24676) );
  nor_x2_sg U39849 ( .A(n23536), .B(n24681), .X(n24680) );
  nand_x2_sg U39850 ( .A(n67402), .B(n57132), .X(n24352) );
  nand_x2_sg U39851 ( .A(n67400), .B(n24272), .X(n24357) );
  nand_x2_sg U39852 ( .A(n67203), .B(n57134), .X(n24258) );
  nand_x2_sg U39853 ( .A(n67406), .B(n24700), .X(n24756) );
  inv_x1_sg U39854 ( .A(n31997), .X(n46884) );
  inv_x2_sg U39855 ( .A(n46884), .X(n46885) );
  inv_x1_sg U39856 ( .A(n58130), .X(n46886) );
  inv_x2_sg U39857 ( .A(n46886), .X(n46887) );
  inv_x1_sg U39858 ( .A(n58128), .X(n46888) );
  inv_x2_sg U39859 ( .A(n46888), .X(n46889) );
  inv_x1_sg U39860 ( .A(\shifter_0/pointer [0]), .X(n46890) );
  inv_x2_sg U39861 ( .A(n46890), .X(n46891) );
  inv_x1_sg U39862 ( .A(\shifter_0/n27115 ), .X(n46892) );
  inv_x2_sg U39863 ( .A(n46892), .X(n46893) );
  inv_x1_sg U39864 ( .A(\shifter_0/reg_w_15 [19]), .X(n46894) );
  inv_x2_sg U39865 ( .A(n46894), .X(n46895) );
  inv_x1_sg U39866 ( .A(\shifter_0/reg_w_15 [18]), .X(n46896) );
  inv_x2_sg U39867 ( .A(n46896), .X(n46897) );
  inv_x1_sg U39868 ( .A(\shifter_0/reg_w_15 [17]), .X(n46898) );
  inv_x2_sg U39869 ( .A(n46898), .X(n46899) );
  inv_x1_sg U39870 ( .A(\shifter_0/reg_w_15 [16]), .X(n46900) );
  inv_x2_sg U39871 ( .A(n46900), .X(n46901) );
  inv_x1_sg U39872 ( .A(\shifter_0/reg_w_15 [15]), .X(n46902) );
  inv_x2_sg U39873 ( .A(n46902), .X(n46903) );
  inv_x1_sg U39874 ( .A(\shifter_0/reg_w_15 [14]), .X(n46904) );
  inv_x2_sg U39875 ( .A(n46904), .X(n46905) );
  inv_x1_sg U39876 ( .A(\shifter_0/reg_w_15 [13]), .X(n46906) );
  inv_x2_sg U39877 ( .A(n46906), .X(n46907) );
  inv_x1_sg U39878 ( .A(\shifter_0/reg_w_15 [12]), .X(n46908) );
  inv_x2_sg U39879 ( .A(n46908), .X(n46909) );
  inv_x1_sg U39880 ( .A(\shifter_0/reg_w_15 [11]), .X(n46910) );
  inv_x2_sg U39881 ( .A(n46910), .X(n46911) );
  inv_x1_sg U39882 ( .A(\shifter_0/reg_w_15 [10]), .X(n46912) );
  inv_x2_sg U39883 ( .A(n46912), .X(n46913) );
  inv_x1_sg U39884 ( .A(\shifter_0/reg_w_15 [9]), .X(n46914) );
  inv_x2_sg U39885 ( .A(n46914), .X(n46915) );
  inv_x1_sg U39886 ( .A(\shifter_0/reg_w_15 [8]), .X(n46916) );
  inv_x2_sg U39887 ( .A(n46916), .X(n46917) );
  inv_x1_sg U39888 ( .A(\shifter_0/reg_w_15 [7]), .X(n46918) );
  inv_x2_sg U39889 ( .A(n46918), .X(n46919) );
  inv_x1_sg U39890 ( .A(\shifter_0/reg_w_15 [6]), .X(n46920) );
  inv_x2_sg U39891 ( .A(n46920), .X(n46921) );
  inv_x1_sg U39892 ( .A(\shifter_0/reg_w_15 [5]), .X(n46922) );
  inv_x2_sg U39893 ( .A(n46922), .X(n46923) );
  inv_x1_sg U39894 ( .A(\shifter_0/reg_w_15 [4]), .X(n46924) );
  inv_x2_sg U39895 ( .A(n46924), .X(n46925) );
  inv_x1_sg U39896 ( .A(\shifter_0/reg_w_15 [3]), .X(n46926) );
  inv_x2_sg U39897 ( .A(n46926), .X(n46927) );
  inv_x1_sg U39898 ( .A(\shifter_0/reg_w_15 [2]), .X(n46928) );
  inv_x2_sg U39899 ( .A(n46928), .X(n46929) );
  inv_x1_sg U39900 ( .A(\shifter_0/reg_w_15 [1]), .X(n46930) );
  inv_x2_sg U39901 ( .A(n46930), .X(n46931) );
  inv_x1_sg U39902 ( .A(\shifter_0/reg_w_15 [0]), .X(n46932) );
  inv_x2_sg U39903 ( .A(n46932), .X(n46933) );
  inv_x1_sg U39904 ( .A(\shifter_0/w_pointer [3]), .X(n46934) );
  inv_x2_sg U39905 ( .A(n46934), .X(n46935) );
  inv_x1_sg U39906 ( .A(\shifter_0/w_pointer [1]), .X(n46936) );
  inv_x2_sg U39907 ( .A(n46936), .X(n46937) );
  inv_x1_sg U39908 ( .A(\shifter_0/reg_w_8 [19]), .X(n46938) );
  inv_x2_sg U39909 ( .A(n46938), .X(n46939) );
  inv_x1_sg U39910 ( .A(\shifter_0/reg_w_8 [18]), .X(n46940) );
  inv_x2_sg U39911 ( .A(n46940), .X(n46941) );
  inv_x1_sg U39912 ( .A(\shifter_0/reg_w_8 [17]), .X(n46942) );
  inv_x2_sg U39913 ( .A(n46942), .X(n46943) );
  inv_x1_sg U39914 ( .A(\shifter_0/reg_w_8 [16]), .X(n46944) );
  inv_x2_sg U39915 ( .A(n46944), .X(n46945) );
  inv_x1_sg U39916 ( .A(\shifter_0/reg_w_8 [15]), .X(n46946) );
  inv_x2_sg U39917 ( .A(n46946), .X(n46947) );
  inv_x1_sg U39918 ( .A(\shifter_0/reg_w_8 [14]), .X(n46948) );
  inv_x2_sg U39919 ( .A(n46948), .X(n46949) );
  inv_x1_sg U39920 ( .A(\shifter_0/reg_w_8 [13]), .X(n46950) );
  inv_x2_sg U39921 ( .A(n46950), .X(n46951) );
  inv_x1_sg U39922 ( .A(\shifter_0/reg_w_8 [12]), .X(n46952) );
  inv_x2_sg U39923 ( .A(n46952), .X(n46953) );
  inv_x1_sg U39924 ( .A(\shifter_0/reg_w_8 [11]), .X(n46954) );
  inv_x2_sg U39925 ( .A(n46954), .X(n46955) );
  inv_x1_sg U39926 ( .A(\shifter_0/reg_w_8 [10]), .X(n46956) );
  inv_x2_sg U39927 ( .A(n46956), .X(n46957) );
  inv_x1_sg U39928 ( .A(\shifter_0/reg_w_8 [9]), .X(n46958) );
  inv_x2_sg U39929 ( .A(n46958), .X(n46959) );
  inv_x1_sg U39930 ( .A(\shifter_0/reg_w_8 [8]), .X(n46960) );
  inv_x2_sg U39931 ( .A(n46960), .X(n46961) );
  inv_x1_sg U39932 ( .A(\shifter_0/reg_w_8 [7]), .X(n46962) );
  inv_x2_sg U39933 ( .A(n46962), .X(n46963) );
  inv_x1_sg U39934 ( .A(\shifter_0/reg_w_8 [6]), .X(n46964) );
  inv_x2_sg U39935 ( .A(n46964), .X(n46965) );
  inv_x1_sg U39936 ( .A(\shifter_0/reg_w_8 [5]), .X(n46966) );
  inv_x2_sg U39937 ( .A(n46966), .X(n46967) );
  inv_x1_sg U39938 ( .A(\shifter_0/reg_w_8 [4]), .X(n46968) );
  inv_x2_sg U39939 ( .A(n46968), .X(n46969) );
  inv_x1_sg U39940 ( .A(\shifter_0/reg_w_8 [3]), .X(n46970) );
  inv_x2_sg U39941 ( .A(n46970), .X(n46971) );
  inv_x1_sg U39942 ( .A(\shifter_0/reg_w_8 [2]), .X(n46972) );
  inv_x2_sg U39943 ( .A(n46972), .X(n46973) );
  inv_x1_sg U39944 ( .A(\shifter_0/reg_w_8 [1]), .X(n46974) );
  inv_x2_sg U39945 ( .A(n46974), .X(n46975) );
  inv_x1_sg U39946 ( .A(\shifter_0/reg_w_8 [0]), .X(n46976) );
  inv_x2_sg U39947 ( .A(n46976), .X(n46977) );
  inv_x1_sg U39948 ( .A(\shifter_0/reg_w_7 [19]), .X(n46978) );
  inv_x2_sg U39949 ( .A(n46978), .X(n46979) );
  inv_x1_sg U39950 ( .A(\shifter_0/reg_w_7 [18]), .X(n46980) );
  inv_x2_sg U39951 ( .A(n46980), .X(n46981) );
  inv_x1_sg U39952 ( .A(\shifter_0/reg_w_7 [17]), .X(n46982) );
  inv_x2_sg U39953 ( .A(n46982), .X(n46983) );
  inv_x1_sg U39954 ( .A(\shifter_0/reg_w_7 [16]), .X(n46984) );
  inv_x2_sg U39955 ( .A(n46984), .X(n46985) );
  inv_x1_sg U39956 ( .A(\shifter_0/reg_w_7 [15]), .X(n46986) );
  inv_x2_sg U39957 ( .A(n46986), .X(n46987) );
  inv_x1_sg U39958 ( .A(\shifter_0/reg_w_7 [14]), .X(n46988) );
  inv_x2_sg U39959 ( .A(n46988), .X(n46989) );
  inv_x1_sg U39960 ( .A(\shifter_0/reg_w_7 [13]), .X(n46990) );
  inv_x2_sg U39961 ( .A(n46990), .X(n46991) );
  inv_x1_sg U39962 ( .A(\shifter_0/reg_w_7 [12]), .X(n46992) );
  inv_x2_sg U39963 ( .A(n46992), .X(n46993) );
  inv_x1_sg U39964 ( .A(\shifter_0/reg_w_7 [11]), .X(n46994) );
  inv_x2_sg U39965 ( .A(n46994), .X(n46995) );
  inv_x1_sg U39966 ( .A(\shifter_0/reg_w_7 [10]), .X(n46996) );
  inv_x2_sg U39967 ( .A(n46996), .X(n46997) );
  inv_x1_sg U39968 ( .A(\shifter_0/reg_w_7 [9]), .X(n46998) );
  inv_x2_sg U39969 ( .A(n46998), .X(n46999) );
  inv_x1_sg U39970 ( .A(\shifter_0/reg_w_7 [8]), .X(n47000) );
  inv_x2_sg U39971 ( .A(n47000), .X(n47001) );
  inv_x1_sg U39972 ( .A(\shifter_0/reg_w_7 [7]), .X(n47002) );
  inv_x2_sg U39973 ( .A(n47002), .X(n47003) );
  inv_x1_sg U39974 ( .A(\shifter_0/reg_w_7 [6]), .X(n47004) );
  inv_x2_sg U39975 ( .A(n47004), .X(n47005) );
  inv_x1_sg U39976 ( .A(\shifter_0/reg_w_7 [5]), .X(n47006) );
  inv_x2_sg U39977 ( .A(n47006), .X(n47007) );
  inv_x1_sg U39978 ( .A(\shifter_0/reg_w_7 [4]), .X(n47008) );
  inv_x2_sg U39979 ( .A(n47008), .X(n47009) );
  inv_x1_sg U39980 ( .A(\shifter_0/reg_w_7 [3]), .X(n47010) );
  inv_x2_sg U39981 ( .A(n47010), .X(n47011) );
  inv_x1_sg U39982 ( .A(\shifter_0/reg_w_7 [2]), .X(n47012) );
  inv_x2_sg U39983 ( .A(n47012), .X(n47013) );
  inv_x1_sg U39984 ( .A(\shifter_0/reg_w_7 [1]), .X(n47014) );
  inv_x2_sg U39985 ( .A(n47014), .X(n47015) );
  inv_x1_sg U39986 ( .A(\shifter_0/reg_w_7 [0]), .X(n47016) );
  inv_x2_sg U39987 ( .A(n47016), .X(n47017) );
  inv_x1_sg U39988 ( .A(\shifter_0/reg_w_1 [19]), .X(n47018) );
  inv_x2_sg U39989 ( .A(n47018), .X(n47019) );
  inv_x1_sg U39990 ( .A(\shifter_0/reg_w_1 [16]), .X(n47020) );
  inv_x2_sg U39991 ( .A(n47020), .X(n47021) );
  inv_x1_sg U39992 ( .A(\shifter_0/reg_w_1 [15]), .X(n47022) );
  inv_x2_sg U39993 ( .A(n47022), .X(n47023) );
  inv_x1_sg U39994 ( .A(\shifter_0/reg_w_1 [14]), .X(n47024) );
  inv_x2_sg U39995 ( .A(n47024), .X(n47025) );
  inv_x1_sg U39996 ( .A(\shifter_0/reg_w_1 [11]), .X(n47026) );
  inv_x2_sg U39997 ( .A(n47026), .X(n47027) );
  inv_x1_sg U39998 ( .A(\shifter_0/reg_w_1 [10]), .X(n47028) );
  inv_x2_sg U39999 ( .A(n47028), .X(n47029) );
  inv_x1_sg U40000 ( .A(\shifter_0/reg_w_1 [7]), .X(n47030) );
  inv_x2_sg U40001 ( .A(n47030), .X(n47031) );
  inv_x1_sg U40002 ( .A(\shifter_0/reg_w_1 [6]), .X(n47032) );
  inv_x2_sg U40003 ( .A(n47032), .X(n47033) );
  inv_x1_sg U40004 ( .A(\shifter_0/reg_w_1 [5]), .X(n47034) );
  inv_x2_sg U40005 ( .A(n47034), .X(n47035) );
  inv_x1_sg U40006 ( .A(\shifter_0/reg_w_1 [2]), .X(n47036) );
  inv_x2_sg U40007 ( .A(n47036), .X(n47037) );
  inv_x1_sg U40008 ( .A(\shifter_0/reg_w_1 [1]), .X(n47038) );
  inv_x2_sg U40009 ( .A(n47038), .X(n47039) );
  inv_x1_sg U40010 ( .A(\shifter_0/reg_w_1 [0]), .X(n47040) );
  inv_x2_sg U40011 ( .A(n47040), .X(n47041) );
  inv_x1_sg U40012 ( .A(\shifter_0/reg_i_15 [19]), .X(n47042) );
  inv_x2_sg U40013 ( .A(n47042), .X(n47043) );
  inv_x1_sg U40014 ( .A(\shifter_0/reg_i_15 [18]), .X(n47044) );
  inv_x2_sg U40015 ( .A(n47044), .X(n47045) );
  inv_x1_sg U40016 ( .A(\shifter_0/reg_i_15 [17]), .X(n47046) );
  inv_x2_sg U40017 ( .A(n47046), .X(n47047) );
  inv_x1_sg U40018 ( .A(\shifter_0/reg_i_15 [16]), .X(n47048) );
  inv_x2_sg U40019 ( .A(n47048), .X(n47049) );
  inv_x1_sg U40020 ( .A(\shifter_0/reg_i_15 [15]), .X(n47050) );
  inv_x2_sg U40021 ( .A(n47050), .X(n47051) );
  inv_x1_sg U40022 ( .A(\shifter_0/reg_i_15 [14]), .X(n47052) );
  inv_x2_sg U40023 ( .A(n47052), .X(n47053) );
  inv_x1_sg U40024 ( .A(\shifter_0/reg_i_15 [13]), .X(n47054) );
  inv_x2_sg U40025 ( .A(n47054), .X(n47055) );
  inv_x1_sg U40026 ( .A(\shifter_0/reg_i_15 [12]), .X(n47056) );
  inv_x2_sg U40027 ( .A(n47056), .X(n47057) );
  inv_x1_sg U40028 ( .A(\shifter_0/reg_i_15 [11]), .X(n47058) );
  inv_x2_sg U40029 ( .A(n47058), .X(n47059) );
  inv_x1_sg U40030 ( .A(\shifter_0/reg_i_15 [10]), .X(n47060) );
  inv_x2_sg U40031 ( .A(n47060), .X(n47061) );
  inv_x1_sg U40032 ( .A(\shifter_0/reg_i_15 [9]), .X(n47062) );
  inv_x2_sg U40033 ( .A(n47062), .X(n47063) );
  inv_x1_sg U40034 ( .A(\shifter_0/reg_i_15 [8]), .X(n47064) );
  inv_x2_sg U40035 ( .A(n47064), .X(n47065) );
  inv_x1_sg U40036 ( .A(\shifter_0/reg_i_15 [7]), .X(n47066) );
  inv_x2_sg U40037 ( .A(n47066), .X(n47067) );
  inv_x1_sg U40038 ( .A(\shifter_0/reg_i_15 [6]), .X(n47068) );
  inv_x2_sg U40039 ( .A(n47068), .X(n47069) );
  inv_x1_sg U40040 ( .A(\shifter_0/reg_i_15 [5]), .X(n47070) );
  inv_x2_sg U40041 ( .A(n47070), .X(n47071) );
  inv_x1_sg U40042 ( .A(\shifter_0/reg_i_15 [4]), .X(n47072) );
  inv_x2_sg U40043 ( .A(n47072), .X(n47073) );
  inv_x1_sg U40044 ( .A(\shifter_0/reg_i_15 [3]), .X(n47074) );
  inv_x2_sg U40045 ( .A(n47074), .X(n47075) );
  inv_x1_sg U40046 ( .A(\shifter_0/reg_i_15 [2]), .X(n47076) );
  inv_x2_sg U40047 ( .A(n47076), .X(n47077) );
  inv_x1_sg U40048 ( .A(\shifter_0/reg_i_15 [1]), .X(n47078) );
  inv_x2_sg U40049 ( .A(n47078), .X(n47079) );
  inv_x1_sg U40050 ( .A(\shifter_0/reg_i_15 [0]), .X(n47080) );
  inv_x2_sg U40051 ( .A(n47080), .X(n47081) );
  inv_x1_sg U40052 ( .A(\shifter_0/reg_i_8 [19]), .X(n47082) );
  inv_x2_sg U40053 ( .A(n47082), .X(n47083) );
  inv_x1_sg U40054 ( .A(\shifter_0/reg_i_8 [18]), .X(n47084) );
  inv_x2_sg U40055 ( .A(n47084), .X(n47085) );
  inv_x1_sg U40056 ( .A(\shifter_0/reg_i_8 [17]), .X(n47086) );
  inv_x2_sg U40057 ( .A(n47086), .X(n47087) );
  inv_x1_sg U40058 ( .A(\shifter_0/reg_i_8 [16]), .X(n47088) );
  inv_x2_sg U40059 ( .A(n47088), .X(n47089) );
  inv_x1_sg U40060 ( .A(\shifter_0/reg_i_8 [15]), .X(n47090) );
  inv_x2_sg U40061 ( .A(n47090), .X(n47091) );
  inv_x1_sg U40062 ( .A(\shifter_0/reg_i_8 [14]), .X(n47092) );
  inv_x2_sg U40063 ( .A(n47092), .X(n47093) );
  inv_x1_sg U40064 ( .A(\shifter_0/reg_i_8 [13]), .X(n47094) );
  inv_x2_sg U40065 ( .A(n47094), .X(n47095) );
  inv_x1_sg U40066 ( .A(\shifter_0/reg_i_8 [12]), .X(n47096) );
  inv_x2_sg U40067 ( .A(n47096), .X(n47097) );
  inv_x1_sg U40068 ( .A(\shifter_0/reg_i_8 [11]), .X(n47098) );
  inv_x2_sg U40069 ( .A(n47098), .X(n47099) );
  inv_x1_sg U40070 ( .A(\shifter_0/reg_i_8 [10]), .X(n47100) );
  inv_x2_sg U40071 ( .A(n47100), .X(n47101) );
  inv_x1_sg U40072 ( .A(\shifter_0/reg_i_8 [9]), .X(n47102) );
  inv_x2_sg U40073 ( .A(n47102), .X(n47103) );
  inv_x1_sg U40074 ( .A(\shifter_0/reg_i_8 [8]), .X(n47104) );
  inv_x2_sg U40075 ( .A(n47104), .X(n47105) );
  inv_x1_sg U40076 ( .A(\shifter_0/reg_i_8 [7]), .X(n47106) );
  inv_x2_sg U40077 ( .A(n47106), .X(n47107) );
  inv_x1_sg U40078 ( .A(\shifter_0/reg_i_8 [6]), .X(n47108) );
  inv_x2_sg U40079 ( .A(n47108), .X(n47109) );
  inv_x1_sg U40080 ( .A(\shifter_0/reg_i_8 [5]), .X(n47110) );
  inv_x2_sg U40081 ( .A(n47110), .X(n47111) );
  inv_x1_sg U40082 ( .A(\shifter_0/reg_i_8 [4]), .X(n47112) );
  inv_x2_sg U40083 ( .A(n47112), .X(n47113) );
  inv_x1_sg U40084 ( .A(\shifter_0/reg_i_8 [3]), .X(n47114) );
  inv_x2_sg U40085 ( .A(n47114), .X(n47115) );
  inv_x1_sg U40086 ( .A(\shifter_0/reg_i_8 [2]), .X(n47116) );
  inv_x2_sg U40087 ( .A(n47116), .X(n47117) );
  inv_x1_sg U40088 ( .A(\shifter_0/reg_i_8 [1]), .X(n47118) );
  inv_x2_sg U40089 ( .A(n47118), .X(n47119) );
  inv_x1_sg U40090 ( .A(\shifter_0/reg_i_8 [0]), .X(n47120) );
  inv_x2_sg U40091 ( .A(n47120), .X(n47121) );
  inv_x1_sg U40092 ( .A(\shifter_0/reg_i_7 [19]), .X(n47122) );
  inv_x2_sg U40093 ( .A(n47122), .X(n47123) );
  inv_x1_sg U40094 ( .A(\shifter_0/reg_i_7 [18]), .X(n47124) );
  inv_x2_sg U40095 ( .A(n47124), .X(n47125) );
  inv_x1_sg U40096 ( .A(\shifter_0/reg_i_7 [17]), .X(n47126) );
  inv_x2_sg U40097 ( .A(n47126), .X(n47127) );
  inv_x1_sg U40098 ( .A(\shifter_0/reg_i_7 [16]), .X(n47128) );
  inv_x2_sg U40099 ( .A(n47128), .X(n47129) );
  inv_x1_sg U40100 ( .A(\shifter_0/reg_i_7 [15]), .X(n47130) );
  inv_x2_sg U40101 ( .A(n47130), .X(n47131) );
  inv_x1_sg U40102 ( .A(\shifter_0/reg_i_7 [14]), .X(n47132) );
  inv_x2_sg U40103 ( .A(n47132), .X(n47133) );
  inv_x1_sg U40104 ( .A(\shifter_0/reg_i_7 [13]), .X(n47134) );
  inv_x2_sg U40105 ( .A(n47134), .X(n47135) );
  inv_x1_sg U40106 ( .A(\shifter_0/reg_i_7 [12]), .X(n47136) );
  inv_x2_sg U40107 ( .A(n47136), .X(n47137) );
  inv_x1_sg U40108 ( .A(\shifter_0/reg_i_7 [11]), .X(n47138) );
  inv_x2_sg U40109 ( .A(n47138), .X(n47139) );
  inv_x1_sg U40110 ( .A(\shifter_0/reg_i_7 [10]), .X(n47140) );
  inv_x2_sg U40111 ( .A(n47140), .X(n47141) );
  inv_x1_sg U40112 ( .A(\shifter_0/reg_i_7 [9]), .X(n47142) );
  inv_x2_sg U40113 ( .A(n47142), .X(n47143) );
  inv_x1_sg U40114 ( .A(\shifter_0/reg_i_7 [8]), .X(n47144) );
  inv_x2_sg U40115 ( .A(n47144), .X(n47145) );
  inv_x1_sg U40116 ( .A(\shifter_0/reg_i_7 [7]), .X(n47146) );
  inv_x2_sg U40117 ( .A(n47146), .X(n47147) );
  inv_x1_sg U40118 ( .A(\shifter_0/reg_i_7 [6]), .X(n47148) );
  inv_x2_sg U40119 ( .A(n47148), .X(n47149) );
  inv_x1_sg U40120 ( .A(\shifter_0/reg_i_7 [5]), .X(n47150) );
  inv_x2_sg U40121 ( .A(n47150), .X(n47151) );
  inv_x1_sg U40122 ( .A(\shifter_0/reg_i_7 [4]), .X(n47152) );
  inv_x2_sg U40123 ( .A(n47152), .X(n47153) );
  inv_x1_sg U40124 ( .A(\shifter_0/reg_i_7 [3]), .X(n47154) );
  inv_x2_sg U40125 ( .A(n47154), .X(n47155) );
  inv_x1_sg U40126 ( .A(\shifter_0/reg_i_7 [2]), .X(n47156) );
  inv_x2_sg U40127 ( .A(n47156), .X(n47157) );
  inv_x1_sg U40128 ( .A(\shifter_0/reg_i_7 [1]), .X(n47158) );
  inv_x2_sg U40129 ( .A(n47158), .X(n47159) );
  inv_x1_sg U40130 ( .A(\shifter_0/reg_i_7 [0]), .X(n47160) );
  inv_x2_sg U40131 ( .A(n47160), .X(n47161) );
  inv_x1_sg U40132 ( .A(\shifter_0/reg_i_1 [19]), .X(n47162) );
  inv_x2_sg U40133 ( .A(n47162), .X(n47163) );
  inv_x1_sg U40134 ( .A(\shifter_0/reg_i_1 [16]), .X(n47164) );
  inv_x2_sg U40135 ( .A(n47164), .X(n47165) );
  inv_x1_sg U40136 ( .A(\shifter_0/reg_i_1 [15]), .X(n47166) );
  inv_x2_sg U40137 ( .A(n47166), .X(n47167) );
  inv_x1_sg U40138 ( .A(\shifter_0/reg_i_1 [14]), .X(n47168) );
  inv_x2_sg U40139 ( .A(n47168), .X(n47169) );
  inv_x1_sg U40140 ( .A(\shifter_0/reg_i_1 [11]), .X(n47170) );
  inv_x2_sg U40141 ( .A(n47170), .X(n47171) );
  inv_x1_sg U40142 ( .A(\shifter_0/reg_i_1 [10]), .X(n47172) );
  inv_x2_sg U40143 ( .A(n47172), .X(n47173) );
  inv_x1_sg U40144 ( .A(\shifter_0/reg_i_1 [7]), .X(n47174) );
  inv_x2_sg U40145 ( .A(n47174), .X(n47175) );
  inv_x1_sg U40146 ( .A(\shifter_0/reg_i_1 [6]), .X(n47176) );
  inv_x2_sg U40147 ( .A(n47176), .X(n47177) );
  inv_x1_sg U40148 ( .A(\shifter_0/reg_i_1 [5]), .X(n47178) );
  inv_x2_sg U40149 ( .A(n47178), .X(n47179) );
  inv_x1_sg U40150 ( .A(\shifter_0/reg_i_1 [2]), .X(n47180) );
  inv_x2_sg U40151 ( .A(n47180), .X(n47181) );
  inv_x1_sg U40152 ( .A(\shifter_0/reg_i_1 [1]), .X(n47182) );
  inv_x2_sg U40153 ( .A(n47182), .X(n47183) );
  inv_x1_sg U40154 ( .A(\shifter_0/reg_i_1 [0]), .X(n47184) );
  inv_x2_sg U40155 ( .A(n47184), .X(n47185) );
  inv_x1_sg U40156 ( .A(\shifter_0/i_pointer [1]), .X(n47186) );
  inv_x2_sg U40157 ( .A(n47186), .X(n47187) );
  inv_x1_sg U40158 ( .A(\filter_0/n17949 ), .X(n47188) );
  inv_x2_sg U40159 ( .A(n47188), .X(n47189) );
  inv_x1_sg U40160 ( .A(\filter_0/n17950 ), .X(n47190) );
  inv_x2_sg U40161 ( .A(n47190), .X(n47191) );
  inv_x1_sg U40162 ( .A(\filter_0/w_pointer [0]), .X(n47192) );
  inv_x2_sg U40163 ( .A(n47192), .X(n47193) );
  inv_x1_sg U40164 ( .A(\filter_0/w_pointer [1]), .X(n47194) );
  inv_x2_sg U40165 ( .A(n47194), .X(n47195) );
  inv_x1_sg U40166 ( .A(\filter_0/w_pointer [2]), .X(n47196) );
  inv_x2_sg U40167 ( .A(n47196), .X(n47197) );
  inv_x1_sg U40168 ( .A(\filter_0/w_pointer [3]), .X(n47198) );
  inv_x2_sg U40169 ( .A(n47198), .X(n47199) );
  inv_x1_sg U40170 ( .A(\filter_0/i_pointer [0]), .X(n47200) );
  inv_x2_sg U40171 ( .A(n47200), .X(n47201) );
  inv_x1_sg U40172 ( .A(\filter_0/i_pointer [1]), .X(n47202) );
  inv_x2_sg U40173 ( .A(n47202), .X(n47203) );
  inv_x1_sg U40174 ( .A(\filter_0/i_pointer [2]), .X(n47204) );
  inv_x2_sg U40175 ( .A(n47204), .X(n47205) );
  inv_x1_sg U40176 ( .A(\filter_0/i_pointer [3]), .X(n47206) );
  inv_x2_sg U40177 ( .A(n47206), .X(n47207) );
  inv_x1_sg U40178 ( .A(\filter_0/N12 ), .X(n47208) );
  inv_x2_sg U40179 ( .A(n47208), .X(n47209) );
  inv_x1_sg U40180 ( .A(\filter_0/N14 ), .X(n47210) );
  inv_x2_sg U40181 ( .A(n47210), .X(n47211) );
  inv_x1_sg U40182 ( .A(\filter_0/N16 ), .X(n47212) );
  inv_x2_sg U40183 ( .A(n47212), .X(n47213) );
  inv_x1_sg U40184 ( .A(\mask_0/counter [0]), .X(n47214) );
  inv_x2_sg U40185 ( .A(n47214), .X(n47215) );
  inv_x1_sg U40186 ( .A(\mask_0/n1654 ), .X(n47216) );
  inv_x2_sg U40187 ( .A(n47216), .X(n47217) );
  inv_x1_sg U40188 ( .A(\mask_0/n1655 ), .X(n47218) );
  inv_x2_sg U40189 ( .A(n47218), .X(n47219) );
  inv_x1_sg U40190 ( .A(n69232), .X(n47220) );
  inv_x2_sg U40191 ( .A(n47220), .X(n47221) );
  inv_x1_sg U40192 ( .A(n69233), .X(n47222) );
  inv_x2_sg U40193 ( .A(n47222), .X(n47223) );
  inv_x1_sg U40194 ( .A(n69234), .X(n47224) );
  inv_x2_sg U40195 ( .A(n47224), .X(n47225) );
  inv_x1_sg U40196 ( .A(n69235), .X(n47226) );
  inv_x2_sg U40197 ( .A(n47226), .X(n47227) );
  inv_x1_sg U40198 ( .A(n69236), .X(n47228) );
  inv_x2_sg U40199 ( .A(n47228), .X(n47229) );
  inv_x1_sg U40200 ( .A(n69237), .X(n47230) );
  inv_x2_sg U40201 ( .A(n47230), .X(n47231) );
  inv_x1_sg U40202 ( .A(n69238), .X(n47232) );
  inv_x2_sg U40203 ( .A(n47232), .X(n47233) );
  inv_x1_sg U40204 ( .A(n69239), .X(n47234) );
  inv_x2_sg U40205 ( .A(n47234), .X(n47235) );
  inv_x1_sg U40206 ( .A(n69240), .X(n47236) );
  inv_x2_sg U40207 ( .A(n47236), .X(n47237) );
  inv_x1_sg U40208 ( .A(n69241), .X(n47238) );
  inv_x2_sg U40209 ( .A(n47238), .X(n47239) );
  inv_x1_sg U40210 ( .A(n69242), .X(n47240) );
  inv_x2_sg U40211 ( .A(n47240), .X(n47241) );
  inv_x1_sg U40212 ( .A(n69243), .X(n47242) );
  inv_x2_sg U40213 ( .A(n47242), .X(n47243) );
  inv_x1_sg U40214 ( .A(n69244), .X(n47244) );
  inv_x2_sg U40215 ( .A(n47244), .X(n47245) );
  inv_x1_sg U40216 ( .A(n69245), .X(n47246) );
  inv_x2_sg U40217 ( .A(n47246), .X(n47247) );
  inv_x1_sg U40218 ( .A(n69246), .X(n47248) );
  inv_x2_sg U40219 ( .A(n47248), .X(n47249) );
  inv_x1_sg U40220 ( .A(n69247), .X(n47250) );
  inv_x2_sg U40221 ( .A(n47250), .X(n47251) );
  inv_x1_sg U40222 ( .A(n69248), .X(n47252) );
  inv_x2_sg U40223 ( .A(n47252), .X(n47253) );
  inv_x1_sg U40224 ( .A(n69249), .X(n47254) );
  inv_x2_sg U40225 ( .A(n47254), .X(n47255) );
  inv_x1_sg U40226 ( .A(n69250), .X(n47256) );
  inv_x2_sg U40227 ( .A(n47256), .X(n47257) );
  inv_x1_sg U40228 ( .A(n69251), .X(n47258) );
  inv_x2_sg U40229 ( .A(n47258), .X(n47259) );
  inv_x1_sg U40230 ( .A(n69252), .X(n47260) );
  inv_x2_sg U40231 ( .A(n47260), .X(n47261) );
  inv_x1_sg U40232 ( .A(n69253), .X(n47262) );
  inv_x2_sg U40233 ( .A(n47262), .X(n47263) );
  inv_x1_sg U40234 ( .A(n69254), .X(n47264) );
  inv_x2_sg U40235 ( .A(n47264), .X(n47265) );
  inv_x1_sg U40236 ( .A(n69255), .X(n47266) );
  inv_x2_sg U40237 ( .A(n47266), .X(n47267) );
  inv_x1_sg U40238 ( .A(n69256), .X(n47268) );
  inv_x2_sg U40239 ( .A(n47268), .X(n47269) );
  inv_x1_sg U40240 ( .A(n69257), .X(n47270) );
  inv_x2_sg U40241 ( .A(n47270), .X(n47271) );
  inv_x1_sg U40242 ( .A(n69258), .X(n47272) );
  inv_x2_sg U40243 ( .A(n47272), .X(n47273) );
  inv_x1_sg U40244 ( .A(n69259), .X(n47274) );
  inv_x2_sg U40245 ( .A(n47274), .X(n47275) );
  inv_x1_sg U40246 ( .A(n69260), .X(n47276) );
  inv_x2_sg U40247 ( .A(n47276), .X(n47277) );
  inv_x1_sg U40248 ( .A(n69261), .X(n47278) );
  inv_x2_sg U40249 ( .A(n47278), .X(n47279) );
  inv_x1_sg U40250 ( .A(n69262), .X(n47280) );
  inv_x2_sg U40251 ( .A(n47280), .X(n47281) );
  inv_x1_sg U40252 ( .A(n69263), .X(n47282) );
  inv_x2_sg U40253 ( .A(n47282), .X(n47283) );
  inv_x1_sg U40254 ( .A(n69265), .X(n47284) );
  inv_x2_sg U40255 ( .A(n47284), .X(n47285) );
  inv_x1_sg U40256 ( .A(n69264), .X(n47286) );
  inv_x2_sg U40257 ( .A(n47286), .X(n47287) );
  nand_x2_sg U40258 ( .A(n67414), .B(n57115), .X(n25704) );
  nand_x2_sg U40259 ( .A(n67416), .B(n57115), .X(n25674) );
  nor_x2_sg U40260 ( .A(n23602), .B(n25643), .X(n25642) );
  nor_x2_sg U40261 ( .A(n23596), .B(n25613), .X(n25612) );
  nor_x2_sg U40262 ( .A(n23590), .B(n25583), .X(n25582) );
  nand_x2_sg U40263 ( .A(n67424), .B(n57115), .X(n25554) );
  nor_x2_sg U40264 ( .A(n23488), .B(n25131), .X(n25130) );
  nor_x2_sg U40265 ( .A(n23482), .B(n25101), .X(n25100) );
  nor_x2_sg U40266 ( .A(n23476), .B(n25071), .X(n25070) );
  nor_x2_sg U40267 ( .A(n23620), .B(n24743), .X(n24742) );
  nor_x2_sg U40268 ( .A(n23614), .B(n24739), .X(n24738) );
  nor_x2_sg U40269 ( .A(n23608), .B(n24735), .X(n24734) );
  nand_x2_sg U40270 ( .A(n67420), .B(n57120), .X(n24728) );
  nor_x2_sg U40271 ( .A(n23512), .B(n24665), .X(n24664) );
  nand_x2_sg U40272 ( .A(n67213), .B(n24605), .X(n24662) );
  nand_x2_sg U40273 ( .A(n67215), .B(n57123), .X(n24658) );
  nand_x2_sg U40274 ( .A(n67217), .B(n57124), .X(n24654) );
  nand_x2_sg U40275 ( .A(n67398), .B(n57127), .X(n24583) );
  nor_x2_sg U40276 ( .A(n23638), .B(n24562), .X(n24561) );
  nor_x2_sg U40277 ( .A(n23632), .B(n24557), .X(n24556) );
  nand_x2_sg U40278 ( .A(n67207), .B(n24381), .X(n24466) );
  nand_x2_sg U40279 ( .A(n67209), .B(n57129), .X(n24461) );
  nand_x2_sg U40280 ( .A(n67211), .B(n57130), .X(n24456) );
  nor_x2_sg U40281 ( .A(n23656), .B(n24356), .X(n24355) );
  nor_x2_sg U40282 ( .A(n23650), .B(n24351), .X(n24350) );
  nor_x2_sg U40283 ( .A(n23644), .B(n24346), .X(n24345) );
  nand_x2_sg U40284 ( .A(n67406), .B(n24272), .X(n24342) );
  nand_x2_sg U40285 ( .A(n67408), .B(n57132), .X(n24337) );
  nor_x2_sg U40286 ( .A(n23536), .B(n24257), .X(n24256) );
  nor_x2_sg U40287 ( .A(n23530), .B(n24252), .X(n24251) );
  nor_x2_sg U40288 ( .A(n23668), .B(n23929), .X(n23928) );
  nor_x2_sg U40289 ( .A(n23662), .B(n23923), .X(n23922) );
  nand_x2_sg U40290 ( .A(n67396), .B(n57143), .X(n23670) );
  nor_x2_sg U40291 ( .A(n68443), .B(n68588), .X(n58598) );
  nor_x2_sg U40292 ( .A(n23620), .B(n25733), .X(n25732) );
  nor_x2_sg U40293 ( .A(n23614), .B(n25703), .X(n25702) );
  nor_x2_sg U40294 ( .A(n23608), .B(n25673), .X(n25672) );
  nand_x2_sg U40295 ( .A(n67420), .B(n57115), .X(n25614) );
  nand_x2_sg U40296 ( .A(n67430), .B(n57115), .X(n25464) );
  nand_x2_sg U40297 ( .A(n67213), .B(n57117), .X(n25222) );
  nand_x2_sg U40298 ( .A(n67215), .B(n57117), .X(n25192) );
  nand_x2_sg U40299 ( .A(n67217), .B(n57117), .X(n25162) );
  nor_x2_sg U40300 ( .A(n23452), .B(n24951), .X(n24950) );
  nor_x2_sg U40301 ( .A(n23428), .B(n24831), .X(n24830) );
  nor_x2_sg U40302 ( .A(n23419), .B(n24792), .X(n24791) );
  nand_x2_sg U40303 ( .A(n67410), .B(n57121), .X(n24748) );
  nand_x2_sg U40304 ( .A(n67414), .B(n57120), .X(n24740) );
  nor_x2_sg U40305 ( .A(n23602), .B(n24731), .X(n24730) );
  nor_x2_sg U40306 ( .A(n23596), .B(n24727), .X(n24726) );
  nor_x2_sg U40307 ( .A(n23590), .B(n24723), .X(n24722) );
  nor_x2_sg U40308 ( .A(n23506), .B(n24661), .X(n24660) );
  nand_x2_sg U40309 ( .A(n67219), .B(n24605), .X(n24650) );
  nand_x2_sg U40310 ( .A(n67221), .B(n57123), .X(n24646) );
  nand_x2_sg U40311 ( .A(n67223), .B(n57124), .X(n24642) );
  nor_x2_sg U40312 ( .A(n23656), .B(n24577), .X(n24576) );
  nor_x2_sg U40313 ( .A(n23650), .B(n24572), .X(n24571) );
  nor_x2_sg U40314 ( .A(n23644), .B(n24567), .X(n24566) );
  nand_x2_sg U40315 ( .A(n67406), .B(n24493), .X(n24563) );
  nand_x2_sg U40316 ( .A(n67408), .B(n57126), .X(n24558) );
  nand_x2_sg U40317 ( .A(n67203), .B(n57129), .X(n24476) );
  nand_x2_sg U40318 ( .A(n67398), .B(n57132), .X(n24362) );
  nor_x2_sg U40319 ( .A(n23638), .B(n24341), .X(n24340) );
  nor_x2_sg U40320 ( .A(n23632), .B(n24336), .X(n24335) );
  nor_x2_sg U40321 ( .A(n23626), .B(n24331), .X(n24330) );
  nand_x2_sg U40322 ( .A(n67412), .B(n24272), .X(n24327) );
  nand_x2_sg U40323 ( .A(n67207), .B(n24163), .X(n24248) );
  nand_x2_sg U40324 ( .A(n67209), .B(n57134), .X(n24243) );
  nand_x2_sg U40325 ( .A(n67211), .B(n57135), .X(n24238) );
  nand_x2_sg U40326 ( .A(n67396), .B(n57137), .X(n23930) );
  nor_x2_sg U40327 ( .A(n23524), .B(n23788), .X(n23787) );
  nor_x2_sg U40328 ( .A(n23518), .B(n23782), .X(n23781) );
  nor_x2_sg U40329 ( .A(n23512), .B(n23776), .X(n23775) );
  nor_x2_sg U40330 ( .A(n23668), .B(n23669), .X(n23667) );
  nor_x2_sg U40331 ( .A(n23662), .B(n23663), .X(n23661) );
  nand_x2_sg U40332 ( .A(n67400), .B(n23556), .X(n23658) );
  nand_x2_sg U40333 ( .A(n67402), .B(n57143), .X(n23652) );
  nor_x2_sg U40334 ( .A(n23536), .B(n23537), .X(n23535) );
  nor_x2_sg U40335 ( .A(n23530), .B(n23531), .X(n23529) );
  inv_x1_sg U40336 ( .A(n32373), .X(n47288) );
  nor_x8_sg U40337 ( .A(n26034), .B(n68385), .X(n26023) );
  nor_x2_sg U40338 ( .A(n35838), .B(n57779), .X(n35837) );
  nor_x2_sg U40339 ( .A(n68372), .B(n35705), .X(n35838) );
  nand_x2_sg U40340 ( .A(n67418), .B(n57115), .X(n25644) );
  nand_x2_sg U40341 ( .A(n67426), .B(n57115), .X(n25524) );
  nand_x2_sg U40342 ( .A(n67428), .B(n57115), .X(n25494) );
  nor_x2_sg U40343 ( .A(n23566), .B(n25463), .X(n25462) );
  nor_x2_sg U40344 ( .A(n23560), .B(n25433), .X(n25432) );
  nor_x2_sg U40345 ( .A(n23553), .B(n25403), .X(n25402) );
  nand_x2_sg U40346 ( .A(n67225), .B(n57117), .X(n25042) );
  nand_x2_sg U40347 ( .A(n67227), .B(n57117), .X(n25012) );
  nand_x2_sg U40348 ( .A(n67229), .B(n57117), .X(n24982) );
  nor_x2_sg U40349 ( .A(n23446), .B(n24921), .X(n24920) );
  nor_x2_sg U40350 ( .A(n23440), .B(n24891), .X(n24890) );
  nor_x2_sg U40351 ( .A(n23434), .B(n24861), .X(n24860) );
  nor_x2_sg U40352 ( .A(n23584), .B(n24719), .X(n24718) );
  nor_x2_sg U40353 ( .A(n23578), .B(n24715), .X(n24714) );
  nor_x2_sg U40354 ( .A(n23572), .B(n24711), .X(n24710) );
  nand_x2_sg U40355 ( .A(n67432), .B(n57120), .X(n24704) );
  nand_x2_sg U40356 ( .A(n67434), .B(n57121), .X(n24699) );
  nor_x2_sg U40357 ( .A(n23452), .B(n24625), .X(n24624) );
  nand_x2_sg U40358 ( .A(n67233), .B(n57123), .X(n24622) );
  nand_x2_sg U40359 ( .A(n67235), .B(n57124), .X(n24618) );
  nand_x2_sg U40360 ( .A(n67237), .B(n24605), .X(n24614) );
  nor_x2_sg U40361 ( .A(n23428), .B(n24609), .X(n24608) );
  nor_x2_sg U40362 ( .A(n23419), .B(n24603), .X(n24602) );
  nor_x2_sg U40363 ( .A(n23668), .B(n24587), .X(n24586) );
  nor_x2_sg U40364 ( .A(n23662), .B(n24582), .X(n24581) );
  nor_x2_sg U40365 ( .A(n23470), .B(n24420), .X(n24419) );
  nor_x2_sg U40366 ( .A(n23464), .B(n24415), .X(n24414) );
  nor_x2_sg U40367 ( .A(n23458), .B(n24410), .X(n24409) );
  nand_x2_sg U40368 ( .A(n67396), .B(n57132), .X(n24367) );
  nand_x2_sg U40369 ( .A(n67424), .B(n24272), .X(n24297) );
  nor_x2_sg U40370 ( .A(n23506), .B(n24232), .X(n24231) );
  nor_x2_sg U40371 ( .A(n23500), .B(n24227), .X(n24226) );
  nor_x2_sg U40372 ( .A(n23494), .B(n24222), .X(n24221) );
  nand_x2_sg U40373 ( .A(n67400), .B(n23816), .X(n23918) );
  nand_x2_sg U40374 ( .A(n67402), .B(n57137), .X(n23912) );
  nor_x2_sg U40375 ( .A(n23638), .B(n23899), .X(n23898) );
  nor_x2_sg U40376 ( .A(n23632), .B(n23893), .X(n23892) );
  nor_x2_sg U40377 ( .A(n23626), .B(n23887), .X(n23886) );
  nor_x2_sg U40378 ( .A(n23536), .B(n23800), .X(n23799) );
  nor_x2_sg U40379 ( .A(n23530), .B(n23794), .X(n23793) );
  nand_x2_sg U40380 ( .A(n67207), .B(n23686), .X(n23789) );
  nand_x2_sg U40381 ( .A(n67209), .B(n57140), .X(n23783) );
  nand_x2_sg U40382 ( .A(n67211), .B(n57141), .X(n23777) );
  nand_x2_sg U40383 ( .A(n67398), .B(n57144), .X(n23664) );
  nor_x2_sg U40384 ( .A(n23656), .B(n23657), .X(n23655) );
  nor_x2_sg U40385 ( .A(n23650), .B(n23651), .X(n23649) );
  nor_x2_sg U40386 ( .A(n23644), .B(n23645), .X(n23643) );
  nand_x2_sg U40387 ( .A(n67406), .B(n23556), .X(n23640) );
  nand_x2_sg U40388 ( .A(n67408), .B(n57143), .X(n23634) );
  nand_x2_sg U40389 ( .A(n67203), .B(n57146), .X(n23538) );
  nor_x2_sg U40390 ( .A(n23524), .B(n23525), .X(n23523) );
  nor_x2_sg U40391 ( .A(n23518), .B(n23519), .X(n23517) );
  nor_x2_sg U40392 ( .A(n23512), .B(n23513), .X(n23511) );
  nor_x2_sg U40393 ( .A(n68536), .B(n68588), .X(n58633) );
  inv_x1_sg U40394 ( .A(n32383), .X(n47292) );
  nor_x8_sg U40395 ( .A(n26036), .B(n26034), .X(n26019) );
  nand_x8_sg U40396 ( .A(n67524), .B(n51525), .X(n26036) );
  nor_x2_sg U40397 ( .A(n47439), .B(n68369), .X(n35836) );
  nand_x2_sg U40398 ( .A(n67412), .B(n57115), .X(n25734) );
  nor_x2_sg U40399 ( .A(n23584), .B(n25553), .X(n25552) );
  nor_x2_sg U40400 ( .A(n23578), .B(n25523), .X(n25522) );
  nor_x2_sg U40401 ( .A(n23572), .B(n25493), .X(n25492) );
  nand_x2_sg U40402 ( .A(n67432), .B(n57115), .X(n25434) );
  nand_x2_sg U40403 ( .A(n67434), .B(n57115), .X(n25404) );
  nor_x2_sg U40404 ( .A(n23470), .B(n25041), .X(n25040) );
  nor_x2_sg U40405 ( .A(n23464), .B(n25011), .X(n25010) );
  nor_x2_sg U40406 ( .A(n23458), .B(n24981), .X(n24980) );
  nand_x2_sg U40407 ( .A(n67233), .B(n57117), .X(n24922) );
  nand_x2_sg U40408 ( .A(n67235), .B(n57117), .X(n24892) );
  nand_x2_sg U40409 ( .A(n67237), .B(n57117), .X(n24862) );
  nand_x2_sg U40410 ( .A(n67418), .B(n24700), .X(n24732) );
  nand_x2_sg U40411 ( .A(n67426), .B(n57120), .X(n24716) );
  nand_x2_sg U40412 ( .A(n67428), .B(n57121), .X(n24712) );
  nor_x2_sg U40413 ( .A(n23566), .B(n24707), .X(n24706) );
  nor_x2_sg U40414 ( .A(n23560), .B(n24703), .X(n24702) );
  nor_x2_sg U40415 ( .A(n23553), .B(n24698), .X(n24697) );
  nand_x2_sg U40416 ( .A(n67225), .B(n24605), .X(n24638) );
  nand_x2_sg U40417 ( .A(n67227), .B(n57123), .X(n24634) );
  nand_x2_sg U40418 ( .A(n67229), .B(n57124), .X(n24630) );
  nor_x2_sg U40419 ( .A(n23446), .B(n24621), .X(n24620) );
  nor_x2_sg U40420 ( .A(n23440), .B(n24617), .X(n24616) );
  nor_x2_sg U40421 ( .A(n23434), .B(n24613), .X(n24612) );
  nand_x2_sg U40422 ( .A(n67400), .B(n24493), .X(n24578) );
  nand_x2_sg U40423 ( .A(n67402), .B(n57126), .X(n24573) );
  nor_x2_sg U40424 ( .A(n23590), .B(n24522), .X(n24521) );
  nor_x2_sg U40425 ( .A(n23452), .B(n24405), .X(n24404) );
  nor_x2_sg U40426 ( .A(n23428), .B(n24385), .X(n24384) );
  nor_x2_sg U40427 ( .A(n23419), .B(n24379), .X(n24378) );
  nor_x2_sg U40428 ( .A(n23668), .B(n24366), .X(n24365) );
  nor_x2_sg U40429 ( .A(n23662), .B(n24361), .X(n24360) );
  nand_x2_sg U40430 ( .A(n67416), .B(n57132), .X(n24317) );
  nand_x2_sg U40431 ( .A(n67430), .B(n24272), .X(n24282) );
  nor_x2_sg U40432 ( .A(n23524), .B(n24247), .X(n24246) );
  nor_x2_sg U40433 ( .A(n23518), .B(n24242), .X(n24241) );
  nor_x2_sg U40434 ( .A(n23512), .B(n24237), .X(n24236) );
  nand_x2_sg U40435 ( .A(n67398), .B(n57138), .X(n23924) );
  nor_x2_sg U40436 ( .A(n23656), .B(n23917), .X(n23916) );
  nor_x2_sg U40437 ( .A(n23650), .B(n23911), .X(n23910) );
  nor_x2_sg U40438 ( .A(n23644), .B(n23905), .X(n23904) );
  nand_x2_sg U40439 ( .A(n67406), .B(n23816), .X(n23900) );
  nand_x2_sg U40440 ( .A(n67408), .B(n57137), .X(n23894) );
  nand_x2_sg U40441 ( .A(n67203), .B(n57140), .X(n23801) );
  nor_x2_sg U40442 ( .A(n23488), .B(n23752), .X(n23751) );
  nor_x2_sg U40443 ( .A(n23482), .B(n23746), .X(n23745) );
  nor_x2_sg U40444 ( .A(n23476), .B(n23740), .X(n23739) );
  nor_x2_sg U40445 ( .A(n23638), .B(n23639), .X(n23637) );
  nor_x2_sg U40446 ( .A(n23632), .B(n23633), .X(n23631) );
  nor_x2_sg U40447 ( .A(n23626), .B(n23627), .X(n23625) );
  nand_x2_sg U40448 ( .A(n67207), .B(n23422), .X(n23526) );
  nand_x2_sg U40449 ( .A(n67209), .B(n57146), .X(n23520) );
  nand_x2_sg U40450 ( .A(n67211), .B(n57147), .X(n23514) );
  nor_x2_sg U40451 ( .A(n23506), .B(n23507), .X(n23505) );
  nor_x2_sg U40452 ( .A(n23500), .B(n23501), .X(n23499) );
  nor_x2_sg U40453 ( .A(n23494), .B(n23495), .X(n23493) );
  nor_x2_sg U40454 ( .A(n23935), .B(n23936), .X(n23934) );
  nor_x2_sg U40455 ( .A(n57302), .B(n68391), .X(n23935) );
  nor_x2_sg U40456 ( .A(n68396), .B(n23675), .X(n23673) );
  inv_x1_sg U40457 ( .A(n32481), .X(n47390) );
  inv_x1_sg U40458 ( .A(n31975), .X(n47328) );
  nor_x8_sg U40459 ( .A(n26033), .B(n26034), .X(n26017) );
  nand_x8_sg U40460 ( .A(n67524), .B(n68386), .X(n26033) );
  nor_x2_sg U40461 ( .A(n23668), .B(n25973), .X(n25972) );
  nor_x2_sg U40462 ( .A(n23662), .B(n25943), .X(n25942) );
  nand_x2_sg U40463 ( .A(n67400), .B(n57115), .X(n25914) );
  nor_x2_sg U40464 ( .A(n23530), .B(n25341), .X(n25340) );
  nor_x2_sg U40465 ( .A(n23524), .B(n25311), .X(n25310) );
  nand_x2_sg U40466 ( .A(n67396), .B(n57120), .X(n24776) );
  nor_x2_sg U40467 ( .A(n23644), .B(n24759), .X(n24758) );
  nand_x2_sg U40468 ( .A(n67430), .B(n24700), .X(n24708) );
  nor_x2_sg U40469 ( .A(n23470), .B(n24637), .X(n24636) );
  nor_x2_sg U40470 ( .A(n23464), .B(n24633), .X(n24632) );
  nor_x2_sg U40471 ( .A(n23458), .B(n24629), .X(n24628) );
  nand_x2_sg U40472 ( .A(n67424), .B(n24493), .X(n24518) );
  nand_x2_sg U40473 ( .A(n67426), .B(n57126), .X(n24513) );
  nand_x2_sg U40474 ( .A(n67428), .B(n57127), .X(n24508) );
  nor_x2_sg U40475 ( .A(n23566), .B(n24502), .X(n24501) );
  nor_x2_sg U40476 ( .A(n23560), .B(n24497), .X(n24496) );
  nor_x2_sg U40477 ( .A(n23553), .B(n24491), .X(n24490) );
  nand_x2_sg U40478 ( .A(n67225), .B(n24381), .X(n24421) );
  nand_x2_sg U40479 ( .A(n67227), .B(n57129), .X(n24416) );
  nand_x2_sg U40480 ( .A(n67229), .B(n57130), .X(n24411) );
  nor_x2_sg U40481 ( .A(n23446), .B(n24400), .X(n24399) );
  nor_x2_sg U40482 ( .A(n23440), .B(n24395), .X(n24394) );
  nor_x2_sg U40483 ( .A(n23434), .B(n24390), .X(n24389) );
  nor_x2_sg U40484 ( .A(n23584), .B(n24296), .X(n24295) );
  nor_x2_sg U40485 ( .A(n23578), .B(n24291), .X(n24290) );
  nor_x2_sg U40486 ( .A(n23572), .B(n24286), .X(n24285) );
  nand_x2_sg U40487 ( .A(n67432), .B(n24272), .X(n24277) );
  nand_x2_sg U40488 ( .A(n67434), .B(n57132), .X(n24271) );
  nor_x2_sg U40489 ( .A(n23452), .B(n24187), .X(n24186) );
  nand_x2_sg U40490 ( .A(n67233), .B(n57134), .X(n24183) );
  nand_x2_sg U40491 ( .A(n67235), .B(n57135), .X(n24178) );
  nand_x2_sg U40492 ( .A(n67237), .B(n24163), .X(n24173) );
  nor_x2_sg U40493 ( .A(n23428), .B(n24167), .X(n24166) );
  nor_x2_sg U40494 ( .A(n23419), .B(n24161), .X(n24160) );
  nand_x2_sg U40495 ( .A(n67412), .B(n23816), .X(n23882) );
  nand_x2_sg U40496 ( .A(n67414), .B(n57137), .X(n23876) );
  nand_x2_sg U40497 ( .A(n67416), .B(n57138), .X(n23870) );
  nor_x2_sg U40498 ( .A(n23602), .B(n23863), .X(n23862) );
  nor_x2_sg U40499 ( .A(n23596), .B(n23857), .X(n23856) );
  nor_x2_sg U40500 ( .A(n23590), .B(n23851), .X(n23850) );
  nor_x2_sg U40501 ( .A(n23506), .B(n23770), .X(n23769) );
  nor_x2_sg U40502 ( .A(n23500), .B(n23764), .X(n23763) );
  nor_x2_sg U40503 ( .A(n23494), .B(n23758), .X(n23757) );
  nand_x2_sg U40504 ( .A(n67219), .B(n23686), .X(n23753) );
  nand_x2_sg U40505 ( .A(n67221), .B(n57140), .X(n23747) );
  nand_x2_sg U40506 ( .A(n67223), .B(n57141), .X(n23741) );
  nand_x2_sg U40507 ( .A(n67410), .B(n57144), .X(n23628) );
  nor_x2_sg U40508 ( .A(n23620), .B(n23621), .X(n23619) );
  nor_x2_sg U40509 ( .A(n23614), .B(n23615), .X(n23613) );
  nor_x2_sg U40510 ( .A(n23608), .B(n23609), .X(n23607) );
  nand_x2_sg U40511 ( .A(n67418), .B(n23556), .X(n23604) );
  nand_x2_sg U40512 ( .A(n67420), .B(n57143), .X(n23598) );
  nand_x2_sg U40513 ( .A(n67213), .B(n23422), .X(n23508) );
  nand_x2_sg U40514 ( .A(n67215), .B(n57146), .X(n23502) );
  nand_x2_sg U40515 ( .A(n67217), .B(n57147), .X(n23496) );
  nor_x2_sg U40516 ( .A(n23488), .B(n23489), .X(n23487) );
  nor_x2_sg U40517 ( .A(n23482), .B(n23483), .X(n23481) );
  nor_x2_sg U40518 ( .A(n23476), .B(n23477), .X(n23475) );
  nor_x2_sg U40519 ( .A(n23677), .B(n58379), .X(n58380) );
  nor_x2_sg U40520 ( .A(n57302), .B(n47445), .X(n23677) );
  nand_x2_sg U40521 ( .A(n68371), .B(n47439), .X(n35840) );
  nand_x4_sg U40522 ( .A(n68374), .B(n26046), .X(n26044) );
  inv_x1_sg U40523 ( .A(n31984), .X(n47392) );
  inv_x2_sg U40524 ( .A(n47288), .X(n47289) );
  nor_x8_sg U40525 ( .A(n26034), .B(n68379), .X(n26008) );
  nor_x2_sg U40526 ( .A(n32440), .B(n32372), .X(n32439) );
  nor_x2_sg U40527 ( .A(n23656), .B(n25913), .X(n25912) );
  nor_x2_sg U40528 ( .A(n23650), .B(n25883), .X(n25882) );
  nand_x2_sg U40529 ( .A(n67406), .B(n57115), .X(n25824) );
  nand_x2_sg U40530 ( .A(n67408), .B(n57115), .X(n25794) );
  nor_x2_sg U40531 ( .A(n23626), .B(n25763), .X(n25762) );
  nand_x2_sg U40532 ( .A(n67211), .B(n57117), .X(n25252) );
  nor_x2_sg U40533 ( .A(n23500), .B(n25191), .X(n25190) );
  nor_x2_sg U40534 ( .A(n23494), .B(n25161), .X(n25160) );
  nor_x2_sg U40535 ( .A(n23668), .B(n24775), .X(n24774) );
  nand_x2_sg U40536 ( .A(n67398), .B(n57121), .X(n24772) );
  nor_x2_sg U40537 ( .A(n23638), .B(n24755), .X(n24754) );
  nand_x2_sg U40538 ( .A(n67424), .B(n24700), .X(n24720) );
  nand_x2_sg U40539 ( .A(n67203), .B(n57123), .X(n24682) );
  nor_x2_sg U40540 ( .A(n23488), .B(n24649), .X(n24648) );
  nor_x2_sg U40541 ( .A(n23482), .B(n24645), .X(n24644) );
  nor_x2_sg U40542 ( .A(n23476), .B(n24641), .X(n24640) );
  nor_x2_sg U40543 ( .A(n23584), .B(n24517), .X(n24516) );
  nor_x2_sg U40544 ( .A(n23578), .B(n24512), .X(n24511) );
  nor_x2_sg U40545 ( .A(n23572), .B(n24507), .X(n24506) );
  nand_x2_sg U40546 ( .A(n67430), .B(n24493), .X(n24503) );
  nand_x2_sg U40547 ( .A(n67432), .B(n57126), .X(n24498) );
  nand_x2_sg U40548 ( .A(n67434), .B(n57127), .X(n24492) );
  nor_x2_sg U40549 ( .A(n23524), .B(n24465), .X(n24464) );
  nor_x2_sg U40550 ( .A(n23518), .B(n24460), .X(n24459) );
  nor_x2_sg U40551 ( .A(n23512), .B(n24455), .X(n24454) );
  nand_x2_sg U40552 ( .A(n67233), .B(n57129), .X(n24401) );
  nand_x2_sg U40553 ( .A(n67235), .B(n57130), .X(n24396) );
  nand_x2_sg U40554 ( .A(n67237), .B(n24381), .X(n24391) );
  nand_x2_sg U40555 ( .A(n67426), .B(n24272), .X(n24292) );
  nand_x2_sg U40556 ( .A(n67428), .B(n57132), .X(n24287) );
  nor_x2_sg U40557 ( .A(n23566), .B(n24281), .X(n24280) );
  nor_x2_sg U40558 ( .A(n23560), .B(n24276), .X(n24275) );
  nor_x2_sg U40559 ( .A(n23553), .B(n24270), .X(n24269) );
  nand_x2_sg U40560 ( .A(n67225), .B(n24163), .X(n24203) );
  nand_x2_sg U40561 ( .A(n67227), .B(n57134), .X(n24198) );
  nand_x2_sg U40562 ( .A(n67229), .B(n57135), .X(n24193) );
  nor_x2_sg U40563 ( .A(n23446), .B(n24182), .X(n24181) );
  nor_x2_sg U40564 ( .A(n23440), .B(n24177), .X(n24176) );
  nor_x2_sg U40565 ( .A(n23434), .B(n24172), .X(n24171) );
  nand_x2_sg U40566 ( .A(n67410), .B(n57138), .X(n23888) );
  nor_x2_sg U40567 ( .A(n23620), .B(n23881), .X(n23880) );
  nor_x2_sg U40568 ( .A(n23614), .B(n23875), .X(n23874) );
  nor_x2_sg U40569 ( .A(n23608), .B(n23869), .X(n23868) );
  nand_x2_sg U40570 ( .A(n67418), .B(n23816), .X(n23864) );
  nand_x2_sg U40571 ( .A(n67420), .B(n57137), .X(n23858) );
  nand_x2_sg U40572 ( .A(n67213), .B(n23686), .X(n23771) );
  nand_x2_sg U40573 ( .A(n67215), .B(n57140), .X(n23765) );
  nand_x2_sg U40574 ( .A(n67217), .B(n57141), .X(n23759) );
  nor_x2_sg U40575 ( .A(n23452), .B(n23716), .X(n23715) );
  nor_x2_sg U40576 ( .A(n23428), .B(n23692), .X(n23691) );
  nor_x2_sg U40577 ( .A(n23419), .B(n23684), .X(n23683) );
  nand_x2_sg U40578 ( .A(n67412), .B(n23556), .X(n23622) );
  nand_x2_sg U40579 ( .A(n67414), .B(n57143), .X(n23616) );
  nand_x2_sg U40580 ( .A(n67416), .B(n57144), .X(n23610) );
  nor_x2_sg U40581 ( .A(n23602), .B(n23603), .X(n23601) );
  nor_x2_sg U40582 ( .A(n23596), .B(n23597), .X(n23595) );
  nor_x2_sg U40583 ( .A(n23590), .B(n23591), .X(n23589) );
  nand_x2_sg U40584 ( .A(n67219), .B(n23422), .X(n23490) );
  nand_x2_sg U40585 ( .A(n67221), .B(n57146), .X(n23484) );
  nand_x2_sg U40586 ( .A(n67223), .B(n57147), .X(n23478) );
  nor_x2_sg U40587 ( .A(n23470), .B(n23471), .X(n23469) );
  nor_x2_sg U40588 ( .A(n23464), .B(n23465), .X(n23463) );
  nor_x2_sg U40589 ( .A(n23458), .B(n23459), .X(n23457) );
  nor_x2_sg U40590 ( .A(n47445), .B(n67500), .X(n24597) );
  inv_x2_sg U40591 ( .A(n33998), .X(n68383) );
  inv_x2_sg U40592 ( .A(n47290), .X(n47291) );
  inv_x1_sg U40593 ( .A(n32039), .X(n47309) );
  inv_x1_sg U40594 ( .A(\filter_0/done ), .X(n47410) );
  inv_x2_sg U40595 ( .A(\shifter_0/i_pointer [0]), .X(n47412) );
  inv_x2_sg U40596 ( .A(\shifter_0/w_pointer [0]), .X(n47414) );
  inv_x2_sg U40597 ( .A(\shifter_0/n27114 ), .X(n47354) );
  inv_x2_sg U40598 ( .A(n47292), .X(n47293) );
  inv_x4_sg U40599 ( .A(n47294), .X(n47295) );
  inv_x4_sg U40600 ( .A(n47296), .X(n47297) );
  inv_x4_sg U40601 ( .A(n35842), .X(n68369) );
  nand_x2_sg U40602 ( .A(n35843), .B(n35844), .X(n35842) );
  nor_x2_sg U40603 ( .A(n32371), .B(n32372), .X(n32370) );
  nand_x4_sg U40604 ( .A(n68389), .B(n68391), .X(n32371) );
  nor_x8_sg U40605 ( .A(n33783), .B(n26034), .X(n26014) );
  nand_x8_sg U40606 ( .A(n68380), .B(n56969), .X(n33783) );
  nor_x8_sg U40607 ( .A(n26260), .B(n26034), .X(n26012) );
  nand_x8_sg U40608 ( .A(n67527), .B(n51523), .X(n26260) );
  nand_x2_sg U40609 ( .A(n67398), .B(n57115), .X(n25944) );
  nand_x2_sg U40610 ( .A(n67402), .B(n57115), .X(n25884) );
  nor_x2_sg U40611 ( .A(n23644), .B(n25853), .X(n25852) );
  nor_x2_sg U40612 ( .A(n23638), .B(n25823), .X(n25822) );
  nor_x2_sg U40613 ( .A(n23632), .B(n25793), .X(n25792) );
  nand_x2_sg U40614 ( .A(n67203), .B(n57117), .X(n25372) );
  nor_x2_sg U40615 ( .A(n23518), .B(n25281), .X(n25280) );
  nor_x2_sg U40616 ( .A(n23512), .B(n25251), .X(n25250) );
  nor_x2_sg U40617 ( .A(n23506), .B(n25221), .X(n25220) );
  nand_x2_sg U40618 ( .A(n67400), .B(n24700), .X(n24768) );
  nor_x2_sg U40619 ( .A(n23650), .B(n24763), .X(n24762) );
  nand_x2_sg U40620 ( .A(n67408), .B(n57120), .X(n24752) );
  nor_x2_sg U40621 ( .A(n23626), .B(n24747), .X(n24746) );
  nand_x2_sg U40622 ( .A(n67416), .B(n57121), .X(n24736) );
  nand_x2_sg U40623 ( .A(n67207), .B(n24605), .X(n24674) );
  nand_x2_sg U40624 ( .A(n67209), .B(n57123), .X(n24670) );
  nand_x2_sg U40625 ( .A(n67211), .B(n57124), .X(n24666) );
  nor_x2_sg U40626 ( .A(n23500), .B(n24657), .X(n24656) );
  nor_x2_sg U40627 ( .A(n23494), .B(n24653), .X(n24652) );
  nand_x2_sg U40628 ( .A(n67410), .B(n57127), .X(n24553) );
  nand_x2_sg U40629 ( .A(n67412), .B(n24493), .X(n24548) );
  nand_x2_sg U40630 ( .A(n67414), .B(n57126), .X(n24543) );
  nor_x2_sg U40631 ( .A(n23608), .B(n24537), .X(n24536) );
  nor_x2_sg U40632 ( .A(n23602), .B(n24532), .X(n24531) );
  nor_x2_sg U40633 ( .A(n23596), .B(n24527), .X(n24526) );
  nand_x2_sg U40634 ( .A(n67213), .B(n24381), .X(n24451) );
  nand_x2_sg U40635 ( .A(n67215), .B(n57129), .X(n24446) );
  nand_x2_sg U40636 ( .A(n67217), .B(n57130), .X(n24441) );
  nor_x2_sg U40637 ( .A(n23488), .B(n24435), .X(n24434) );
  nor_x2_sg U40638 ( .A(n23482), .B(n24430), .X(n24429) );
  nor_x2_sg U40639 ( .A(n23476), .B(n24425), .X(n24424) );
  nor_x2_sg U40640 ( .A(n23620), .B(n24326), .X(n24325) );
  nor_x2_sg U40641 ( .A(n23614), .B(n24321), .X(n24320) );
  nand_x2_sg U40642 ( .A(n67418), .B(n24272), .X(n24312) );
  nand_x2_sg U40643 ( .A(n67420), .B(n57132), .X(n24307) );
  nor_x2_sg U40644 ( .A(n23590), .B(n24301), .X(n24300) );
  nand_x2_sg U40645 ( .A(n67219), .B(n24163), .X(n24218) );
  nand_x2_sg U40646 ( .A(n67221), .B(n57134), .X(n24213) );
  nand_x2_sg U40647 ( .A(n67223), .B(n57135), .X(n24208) );
  nor_x2_sg U40648 ( .A(n23470), .B(n24202), .X(n24201) );
  nor_x2_sg U40649 ( .A(n23464), .B(n24197), .X(n24196) );
  nor_x2_sg U40650 ( .A(n23458), .B(n24192), .X(n24191) );
  nand_x2_sg U40651 ( .A(n67424), .B(n23816), .X(n23846) );
  nand_x2_sg U40652 ( .A(n67426), .B(n57137), .X(n23840) );
  nand_x2_sg U40653 ( .A(n67428), .B(n57138), .X(n23834) );
  nor_x2_sg U40654 ( .A(n23566), .B(n23827), .X(n23826) );
  nor_x2_sg U40655 ( .A(n23560), .B(n23821), .X(n23820) );
  nor_x2_sg U40656 ( .A(n23553), .B(n23814), .X(n23813) );
  nand_x2_sg U40657 ( .A(n67225), .B(n23686), .X(n23735) );
  nand_x2_sg U40658 ( .A(n67227), .B(n57140), .X(n23729) );
  nand_x2_sg U40659 ( .A(n67229), .B(n57141), .X(n23723) );
  nor_x2_sg U40660 ( .A(n23446), .B(n23710), .X(n23709) );
  nor_x2_sg U40661 ( .A(n23440), .B(n23704), .X(n23703) );
  nor_x2_sg U40662 ( .A(n23434), .B(n23698), .X(n23697) );
  nor_x2_sg U40663 ( .A(n23584), .B(n23585), .X(n23583) );
  nor_x2_sg U40664 ( .A(n23578), .B(n23579), .X(n23577) );
  nor_x2_sg U40665 ( .A(n23572), .B(n23573), .X(n23571) );
  nand_x2_sg U40666 ( .A(n67430), .B(n23556), .X(n23568) );
  nand_x2_sg U40667 ( .A(n67432), .B(n57143), .X(n23562) );
  nand_x2_sg U40668 ( .A(n67434), .B(n57144), .X(n23555) );
  nor_x2_sg U40669 ( .A(n23452), .B(n23453), .X(n23451) );
  nand_x2_sg U40670 ( .A(n67233), .B(n57146), .X(n23448) );
  nand_x2_sg U40671 ( .A(n67235), .B(n57147), .X(n23442) );
  nand_x2_sg U40672 ( .A(n67237), .B(n23422), .X(n23436) );
  nor_x2_sg U40673 ( .A(n23428), .B(n23429), .X(n23427) );
  nor_x2_sg U40674 ( .A(n23419), .B(n23420), .X(n23418) );
  nor_x2_sg U40675 ( .A(n23186), .B(n57151), .X(n23178) );
  nor_x2_sg U40676 ( .A(n57037), .B(n57152), .X(n23186) );
  nor_x2_sg U40677 ( .A(n24788), .B(n58639), .X(n58052) );
  nor_x8_sg U40678 ( .A(n67500), .B(n68391), .X(n24788) );
  nand_x2_sg U40679 ( .A(n47291), .B(n57862), .X(n23102) );
  nor_x2_sg U40680 ( .A(n25947), .B(n25948), .X(n25946) );
  nor_x2_sg U40681 ( .A(n25953), .B(n25954), .X(n25945) );
  nor_x2_sg U40682 ( .A(n25677), .B(n25678), .X(n25676) );
  nor_x2_sg U40683 ( .A(n25683), .B(n25684), .X(n25675) );
  nor_x2_sg U40684 ( .A(n25315), .B(n25316), .X(n25314) );
  nor_x2_sg U40685 ( .A(n25321), .B(n25322), .X(n25313) );
  nor_x2_sg U40686 ( .A(n25195), .B(n25196), .X(n25194) );
  nor_x2_sg U40687 ( .A(n25201), .B(n25202), .X(n25193) );
  inv_x2_sg U40688 ( .A(n33738), .X(n68378) );
  inv_x2_sg U40689 ( .A(n34219), .X(n68384) );
  inv_x4_sg U40690 ( .A(n47298), .X(n47299) );
  inv_x1_sg U40691 ( .A(n32721), .X(n47300) );
  nand_x4_sg U40692 ( .A(n32722), .B(n32723), .X(n32721) );
  inv_x2_sg U40693 ( .A(n47301), .X(n47302) );
  inv_x2_sg U40694 ( .A(n47303), .X(n47304) );
  inv_x2_sg U40695 ( .A(n47305), .X(n47306) );
  inv_x2_sg U40696 ( .A(n47307), .X(n47308) );
  inv_x1_sg U40697 ( .A(\filter_0/n17951 ), .X(n47336) );
  inv_x1_sg U40698 ( .A(\filter_0/reg_o_mask [15]), .X(n47338) );
  inv_x1_sg U40699 ( .A(\filter_0/reg_o_mask [31]), .X(n47340) );
  inv_x1_sg U40700 ( .A(\filter_0/reg_xor_i_mask [15]), .X(n47342) );
  inv_x1_sg U40701 ( .A(\filter_0/reg_xor_i_mask [31]), .X(n47344) );
  inv_x1_sg U40702 ( .A(\filter_0/reg_xor_w_mask [15]), .X(n47346) );
  inv_x1_sg U40703 ( .A(\filter_0/reg_xor_w_mask [31]), .X(n47348) );
  inv_x1_sg U40704 ( .A(\shifter_0/n27116 ), .X(n47408) );
  inv_x2_sg U40705 ( .A(n47309), .X(n47310) );
  inv_x4_sg U40706 ( .A(n47311), .X(n47312) );
  nand_x4_sg U40707 ( .A(n32510), .B(n32511), .X(n32509) );
  inv_x4_sg U40708 ( .A(n31987), .X(n68570) );
  nand_x2_sg U40709 ( .A(n31988), .B(n31989), .X(n31987) );
  nor_x8_sg U40710 ( .A(n34043), .B(n26034), .X(n26021) );
  nand_x8_sg U40711 ( .A(n68386), .B(n56971), .X(n34043) );
  nand_x4_sg U40712 ( .A(n68572), .B(n47775), .X(n24487) );
  inv_x4_sg U40713 ( .A(n22497), .X(n47313) );
  nor_x8_sg U40714 ( .A(n68390), .B(n47445), .X(n22497) );
  nand_x8_sg U40715 ( .A(n57097), .B(n22695), .X(n22694) );
  nand_x2_sg U40716 ( .A(n22696), .B(n22697), .X(n22695) );
  nor_x4_sg U40717 ( .A(n34228), .B(n57168), .X(n32820) );
  nand_x4_sg U40718 ( .A(n34227), .B(n34229), .X(n34228) );
  inv_x4_sg U40719 ( .A(n35844), .X(n68370) );
  inv_x4_sg U40720 ( .A(n57964), .X(n47316) );
  inv_x8_sg U40721 ( .A(n47316), .X(n47317) );
  nor_x8_sg U40722 ( .A(n57306), .B(n47445), .X(n22546) );
  nor_x8_sg U40723 ( .A(n26258), .B(n26034), .X(n26010) );
  nand_x8_sg U40724 ( .A(n67527), .B(n68380), .X(n26258) );
  nor_x2_sg U40725 ( .A(n38413), .B(n57619), .X(n38412) );
  nor_x2_sg U40726 ( .A(n68272), .B(n38415), .X(n38413) );
  nor_x2_sg U40727 ( .A(n23536), .B(n25371), .X(n25370) );
  nand_x2_sg U40728 ( .A(n67207), .B(n57117), .X(n25312) );
  nand_x2_sg U40729 ( .A(n67209), .B(n57117), .X(n25282) );
  nor_x2_sg U40730 ( .A(n23662), .B(n24771), .X(n24770) );
  nor_x2_sg U40731 ( .A(n23656), .B(n24767), .X(n24766) );
  nand_x2_sg U40732 ( .A(n67402), .B(n57120), .X(n24764) );
  nor_x2_sg U40733 ( .A(n23632), .B(n24751), .X(n24750) );
  nand_x2_sg U40734 ( .A(n67412), .B(n24700), .X(n24744) );
  nor_x2_sg U40735 ( .A(n23524), .B(n24673), .X(n24672) );
  nor_x2_sg U40736 ( .A(n23518), .B(n24669), .X(n24668) );
  nor_x2_sg U40737 ( .A(n23626), .B(n24552), .X(n24551) );
  nor_x2_sg U40738 ( .A(n23620), .B(n24547), .X(n24546) );
  nor_x2_sg U40739 ( .A(n23614), .B(n24542), .X(n24541) );
  nand_x2_sg U40740 ( .A(n67416), .B(n57127), .X(n24538) );
  nand_x2_sg U40741 ( .A(n67418), .B(n24493), .X(n24533) );
  nand_x2_sg U40742 ( .A(n67420), .B(n57126), .X(n24528) );
  nor_x2_sg U40743 ( .A(n23506), .B(n24450), .X(n24449) );
  nor_x2_sg U40744 ( .A(n23500), .B(n24445), .X(n24444) );
  nor_x2_sg U40745 ( .A(n23494), .B(n24440), .X(n24439) );
  nand_x2_sg U40746 ( .A(n67219), .B(n24381), .X(n24436) );
  nand_x2_sg U40747 ( .A(n67221), .B(n57129), .X(n24431) );
  nand_x2_sg U40748 ( .A(n67223), .B(n57130), .X(n24426) );
  nand_x2_sg U40749 ( .A(n67410), .B(n57132), .X(n24332) );
  nand_x2_sg U40750 ( .A(n67414), .B(n24272), .X(n24322) );
  nor_x2_sg U40751 ( .A(n23608), .B(n24316), .X(n24315) );
  nor_x2_sg U40752 ( .A(n23602), .B(n24311), .X(n24310) );
  nor_x2_sg U40753 ( .A(n23596), .B(n24306), .X(n24305) );
  nand_x2_sg U40754 ( .A(n67213), .B(n24163), .X(n24233) );
  nand_x2_sg U40755 ( .A(n67215), .B(n57134), .X(n24228) );
  nand_x2_sg U40756 ( .A(n67217), .B(n57135), .X(n24223) );
  nor_x2_sg U40757 ( .A(n23488), .B(n24217), .X(n24216) );
  nor_x2_sg U40758 ( .A(n23482), .B(n24212), .X(n24211) );
  nor_x2_sg U40759 ( .A(n23476), .B(n24207), .X(n24206) );
  nor_x2_sg U40760 ( .A(n23584), .B(n23845), .X(n23844) );
  nor_x2_sg U40761 ( .A(n23578), .B(n23839), .X(n23838) );
  nor_x2_sg U40762 ( .A(n23572), .B(n23833), .X(n23832) );
  nand_x2_sg U40763 ( .A(n67430), .B(n23816), .X(n23828) );
  nand_x2_sg U40764 ( .A(n67432), .B(n57137), .X(n23822) );
  nand_x2_sg U40765 ( .A(n67434), .B(n57138), .X(n23815) );
  nor_x2_sg U40766 ( .A(n23470), .B(n23734), .X(n23733) );
  nor_x2_sg U40767 ( .A(n23464), .B(n23728), .X(n23727) );
  nor_x2_sg U40768 ( .A(n23458), .B(n23722), .X(n23721) );
  nand_x2_sg U40769 ( .A(n67233), .B(n57140), .X(n23711) );
  nand_x2_sg U40770 ( .A(n67235), .B(n57141), .X(n23705) );
  nand_x2_sg U40771 ( .A(n67237), .B(n23686), .X(n23699) );
  nand_x2_sg U40772 ( .A(n67424), .B(n23556), .X(n23586) );
  nand_x2_sg U40773 ( .A(n67426), .B(n57143), .X(n23580) );
  nand_x2_sg U40774 ( .A(n67428), .B(n57144), .X(n23574) );
  nor_x2_sg U40775 ( .A(n23566), .B(n23567), .X(n23565) );
  nor_x2_sg U40776 ( .A(n23560), .B(n23561), .X(n23559) );
  nor_x2_sg U40777 ( .A(n23553), .B(n23554), .X(n23552) );
  nand_x2_sg U40778 ( .A(n67225), .B(n23422), .X(n23472) );
  nand_x2_sg U40779 ( .A(n67227), .B(n57146), .X(n23466) );
  nand_x2_sg U40780 ( .A(n67229), .B(n57147), .X(n23460) );
  nor_x2_sg U40781 ( .A(n23446), .B(n23447), .X(n23445) );
  nor_x2_sg U40782 ( .A(n23440), .B(n23441), .X(n23439) );
  nor_x2_sg U40783 ( .A(n23434), .B(n23435), .X(n23433) );
  nor_x2_sg U40784 ( .A(n22970), .B(n57157), .X(n22962) );
  nor_x2_sg U40785 ( .A(n57029), .B(n57158), .X(n22970) );
  nor_x2_sg U40786 ( .A(n24829), .B(n68495), .X(n25368) );
  inv_x2_sg U40787 ( .A(n34227), .X(n47318) );
  nand_x4_sg U40788 ( .A(n47411), .B(n57114), .X(n34227) );
  nor_x2_sg U40789 ( .A(n24785), .B(n57099), .X(n58051) );
  nor_x2_sg U40790 ( .A(n24695), .B(n58639), .X(n58122) );
  nor_x8_sg U40791 ( .A(n67096), .B(n68573), .X(n24695) );
  nor_x2_sg U40792 ( .A(n57302), .B(n29338), .X(n23417) );
  nand_x2_sg U40793 ( .A(n47306), .B(n57862), .X(n23190) );
  nand_x2_sg U40794 ( .A(n47308), .B(n57862), .X(n23091) );
  nand_x2_sg U40795 ( .A(n47302), .B(n57862), .X(n22919) );
  nor_x2_sg U40796 ( .A(n25978), .B(n25979), .X(n25977) );
  nor_x2_sg U40797 ( .A(n25984), .B(n25985), .X(n25976) );
  nor_x2_sg U40798 ( .A(n25917), .B(n25918), .X(n25916) );
  nor_x2_sg U40799 ( .A(n25923), .B(n25924), .X(n25915) );
  nor_x2_sg U40800 ( .A(n25887), .B(n25888), .X(n25886) );
  nor_x2_sg U40801 ( .A(n25893), .B(n25894), .X(n25885) );
  nor_x2_sg U40802 ( .A(n25827), .B(n25828), .X(n25826) );
  nor_x2_sg U40803 ( .A(n25833), .B(n25834), .X(n25825) );
  nor_x2_sg U40804 ( .A(n25797), .B(n25798), .X(n25796) );
  nor_x2_sg U40805 ( .A(n25803), .B(n25804), .X(n25795) );
  nor_x2_sg U40806 ( .A(n25767), .B(n25768), .X(n25766) );
  nor_x2_sg U40807 ( .A(n25773), .B(n25774), .X(n25765) );
  nor_x2_sg U40808 ( .A(n25737), .B(n25738), .X(n25736) );
  nor_x2_sg U40809 ( .A(n25743), .B(n25744), .X(n25735) );
  nor_x2_sg U40810 ( .A(n25707), .B(n25708), .X(n25706) );
  nor_x2_sg U40811 ( .A(n25713), .B(n25714), .X(n25705) );
  nor_x2_sg U40812 ( .A(n25647), .B(n25648), .X(n25646) );
  nor_x2_sg U40813 ( .A(n25653), .B(n25654), .X(n25645) );
  nor_x2_sg U40814 ( .A(n25617), .B(n25618), .X(n25616) );
  nor_x2_sg U40815 ( .A(n25623), .B(n25624), .X(n25615) );
  nor_x2_sg U40816 ( .A(n25557), .B(n25558), .X(n25556) );
  nor_x2_sg U40817 ( .A(n25563), .B(n25564), .X(n25555) );
  nor_x2_sg U40818 ( .A(n25527), .B(n25528), .X(n25526) );
  nor_x2_sg U40819 ( .A(n25533), .B(n25534), .X(n25525) );
  nor_x2_sg U40820 ( .A(n25497), .B(n25498), .X(n25496) );
  nor_x2_sg U40821 ( .A(n25503), .B(n25504), .X(n25495) );
  nor_x2_sg U40822 ( .A(n25467), .B(n25468), .X(n25466) );
  nor_x2_sg U40823 ( .A(n25473), .B(n25474), .X(n25465) );
  nor_x2_sg U40824 ( .A(n25437), .B(n25438), .X(n25436) );
  nor_x2_sg U40825 ( .A(n25443), .B(n25444), .X(n25435) );
  nor_x2_sg U40826 ( .A(n25407), .B(n25408), .X(n25406) );
  nor_x2_sg U40827 ( .A(n25413), .B(n25414), .X(n25405) );
  nor_x2_sg U40828 ( .A(n25376), .B(n25377), .X(n25375) );
  nor_x2_sg U40829 ( .A(n25382), .B(n25383), .X(n25374) );
  nor_x2_sg U40830 ( .A(n25285), .B(n25286), .X(n25284) );
  nor_x2_sg U40831 ( .A(n25291), .B(n25292), .X(n25283) );
  nor_x2_sg U40832 ( .A(n25255), .B(n25256), .X(n25254) );
  nor_x2_sg U40833 ( .A(n25261), .B(n25262), .X(n25253) );
  nor_x2_sg U40834 ( .A(n25225), .B(n25226), .X(n25224) );
  nor_x2_sg U40835 ( .A(n25231), .B(n25232), .X(n25223) );
  nor_x2_sg U40836 ( .A(n25165), .B(n25166), .X(n25164) );
  nor_x2_sg U40837 ( .A(n25171), .B(n25172), .X(n25163) );
  nor_x2_sg U40838 ( .A(n25135), .B(n25136), .X(n25134) );
  nor_x2_sg U40839 ( .A(n25141), .B(n25142), .X(n25133) );
  nor_x2_sg U40840 ( .A(n25105), .B(n25106), .X(n25104) );
  nor_x2_sg U40841 ( .A(n25111), .B(n25112), .X(n25103) );
  nor_x2_sg U40842 ( .A(n25075), .B(n25076), .X(n25074) );
  nor_x2_sg U40843 ( .A(n25081), .B(n25082), .X(n25073) );
  nor_x2_sg U40844 ( .A(n25045), .B(n25046), .X(n25044) );
  nor_x2_sg U40845 ( .A(n25051), .B(n25052), .X(n25043) );
  nor_x2_sg U40846 ( .A(n25015), .B(n25016), .X(n25014) );
  nor_x2_sg U40847 ( .A(n25021), .B(n25022), .X(n25013) );
  nor_x2_sg U40848 ( .A(n24985), .B(n24986), .X(n24984) );
  nor_x2_sg U40849 ( .A(n24991), .B(n24992), .X(n24983) );
  nor_x2_sg U40850 ( .A(n24925), .B(n24926), .X(n24924) );
  nor_x2_sg U40851 ( .A(n24931), .B(n24932), .X(n24923) );
  nor_x2_sg U40852 ( .A(n24895), .B(n24896), .X(n24894) );
  nor_x2_sg U40853 ( .A(n24901), .B(n24902), .X(n24893) );
  nor_x2_sg U40854 ( .A(n24865), .B(n24866), .X(n24864) );
  nor_x2_sg U40855 ( .A(n24871), .B(n24872), .X(n24863) );
  inv_x2_sg U40856 ( .A(n34086), .X(n68382) );
  inv_x1_sg U40857 ( .A(n32276), .X(n47319) );
  nand_x4_sg U40858 ( .A(n32277), .B(n32278), .X(n32276) );
  inv_x2_sg U40859 ( .A(n47320), .X(n47321) );
  inv_x2_sg U40860 ( .A(n47322), .X(n47323) );
  inv_x2_sg U40861 ( .A(n47324), .X(n47325) );
  inv_x2_sg U40862 ( .A(n47326), .X(n47327) );
  nor_x8_sg U40863 ( .A(n67085), .B(n22522), .X(n22572) );
  nand_x8_sg U40864 ( .A(n58480), .B(n58483), .X(n67085) );
  inv_x1_sg U40865 ( .A(\filter_0/reg_o_mask [11]), .X(n47396) );
  inv_x1_sg U40866 ( .A(\filter_0/reg_o_mask [27]), .X(n47398) );
  inv_x1_sg U40867 ( .A(\filter_0/reg_xor_i_mask [11]), .X(n47400) );
  inv_x1_sg U40868 ( .A(\filter_0/reg_xor_i_mask [27]), .X(n47402) );
  inv_x1_sg U40869 ( .A(\filter_0/reg_xor_w_mask [11]), .X(n47404) );
  inv_x1_sg U40870 ( .A(\filter_0/reg_xor_w_mask [27]), .X(n47406) );
  inv_x2_sg U40871 ( .A(n47328), .X(n47329) );
  inv_x4_sg U40872 ( .A(n47330), .X(n47331) );
  inv_x4_sg U40873 ( .A(n22471), .X(n67100) );
  nor_x8_sg U40874 ( .A(n68572), .B(n47775), .X(n22471) );
  inv_x1_sg U40875 ( .A(n25991), .X(n47332) );
  inv_x1_sg U40876 ( .A(n25991), .X(n67455) );
  inv_x1_sg U40877 ( .A(n25268), .X(n47333) );
  inv_x1_sg U40878 ( .A(n25268), .X(n67266) );
  nor_x4_sg U40879 ( .A(n57506), .B(n24788), .X(n25401) );
  nand_x8_sg U40880 ( .A(n32517), .B(n32518), .X(n32420) );
  nor_x2_sg U40881 ( .A(n32519), .B(n68463), .X(n32518) );
  nor_x2_sg U40882 ( .A(n32528), .B(n32529), .X(n32517) );
  inv_x4_sg U40883 ( .A(n47334), .X(n47335) );
  nor_x4_sg U40884 ( .A(n47335), .B(n29337), .X(n31998) );
  nor_x2_sg U40885 ( .A(n68571), .B(n68575), .X(n32354) );
  inv_x2_sg U40886 ( .A(n47336), .X(n47337) );
  inv_x2_sg U40887 ( .A(n47338), .X(n47339) );
  inv_x2_sg U40888 ( .A(n47340), .X(n47341) );
  inv_x2_sg U40889 ( .A(n47342), .X(n47343) );
  inv_x2_sg U40890 ( .A(n47344), .X(n47345) );
  inv_x2_sg U40891 ( .A(n47346), .X(n47347) );
  inv_x2_sg U40892 ( .A(n47348), .X(n47349) );
  inv_x8_sg U40893 ( .A(n56971), .X(n67524) );
  inv_x8_sg U40894 ( .A(n56969), .X(n67527) );
  nand_x8_sg U40895 ( .A(n25855), .B(n25856), .X(n23389) );
  nor_x2_sg U40896 ( .A(n25863), .B(n25864), .X(n25855) );
  nor_x2_sg U40897 ( .A(n25857), .B(n25858), .X(n25856) );
  nand_x8_sg U40898 ( .A(n25585), .B(n25586), .X(n23344) );
  nor_x2_sg U40899 ( .A(n25593), .B(n25594), .X(n25585) );
  nor_x2_sg U40900 ( .A(n25587), .B(n25588), .X(n25586) );
  nand_x8_sg U40901 ( .A(n25343), .B(n25344), .X(n23296) );
  nor_x2_sg U40902 ( .A(n25351), .B(n25352), .X(n25343) );
  nor_x2_sg U40903 ( .A(n25345), .B(n25346), .X(n25344) );
  nand_x8_sg U40904 ( .A(n24953), .B(n24954), .X(n23231) );
  nor_x2_sg U40905 ( .A(n24961), .B(n24962), .X(n24953) );
  nor_x2_sg U40906 ( .A(n24955), .B(n24956), .X(n24954) );
  nand_x8_sg U40907 ( .A(n24833), .B(n24834), .X(n23211) );
  nor_x2_sg U40908 ( .A(n24841), .B(n24842), .X(n24833) );
  nor_x2_sg U40909 ( .A(n24835), .B(n24836), .X(n24834) );
  nand_x8_sg U40910 ( .A(n24794), .B(n24795), .X(n23206) );
  nor_x2_sg U40911 ( .A(n24805), .B(n24806), .X(n24794) );
  nor_x2_sg U40912 ( .A(n24796), .B(n24797), .X(n24795) );
  nor_x2_sg U40913 ( .A(n24159), .B(n57328), .X(n24158) );
  nor_x4_sg U40914 ( .A(n23675), .B(n68391), .X(n24159) );
  inv_x4_sg U40915 ( .A(n47219), .X(n47350) );
  inv_x8_sg U40916 ( .A(n47350), .X(n47351) );
  nand_x2_sg U40917 ( .A(n30627), .B(n61905), .X(n30625) );
  nor_x4_sg U40918 ( .A(n68387), .B(n47437), .X(n30627) );
  nor_x4_sg U40919 ( .A(n24599), .B(n67500), .X(n24591) );
  nand_x4_sg U40920 ( .A(n68390), .B(n47445), .X(n24599) );
  inv_x4_sg U40921 ( .A(n47189), .X(n47352) );
  inv_x4_sg U40922 ( .A(n47352), .X(n47353) );
  inv_x4_sg U40923 ( .A(n47353), .X(n68387) );
  nor_x4_sg U40924 ( .A(n68385), .B(n67581), .X(n26162) );
  inv_x8_sg U40925 ( .A(n26177), .X(n67581) );
  nor_x4_sg U40926 ( .A(n68379), .B(n67575), .X(n26066) );
  inv_x8_sg U40927 ( .A(n26060), .X(n67575) );
  inv_x4_sg U40928 ( .A(n47354), .X(n47355) );
  nor_x8_sg U40929 ( .A(n57300), .B(n47775), .X(n22521) );
  nor_x8_sg U40930 ( .A(n68372), .B(n47439), .X(n35844) );
  inv_x8_sg U40931 ( .A(n47351), .X(n68372) );
  inv_x4_sg U40932 ( .A(n47185), .X(n47356) );
  inv_x4_sg U40933 ( .A(n47183), .X(n47358) );
  inv_x4_sg U40934 ( .A(n47179), .X(n47360) );
  inv_x4_sg U40935 ( .A(n47169), .X(n47362) );
  inv_x4_sg U40936 ( .A(n47041), .X(n47364) );
  inv_x4_sg U40937 ( .A(n47039), .X(n47366) );
  inv_x4_sg U40938 ( .A(n47035), .X(n47368) );
  inv_x4_sg U40939 ( .A(n47025), .X(n47370) );
  nand_x2_sg U40940 ( .A(n67404), .B(n57121), .X(n24760) );
  nand_x2_sg U40941 ( .A(n67404), .B(n57132), .X(n24347) );
  nand_x2_sg U40942 ( .A(n67404), .B(n57138), .X(n23906) );
  nand_x2_sg U40943 ( .A(n67404), .B(n57144), .X(n23646) );
  nand_x2_sg U40944 ( .A(n67404), .B(n57115), .X(n25854) );
  nand_x2_sg U40945 ( .A(n67404), .B(n57127), .X(n24568) );
  inv_x8_sg U40946 ( .A(n23644), .X(n67404) );
  nand_x2_sg U40947 ( .A(n67422), .B(n57121), .X(n24724) );
  nand_x2_sg U40948 ( .A(n67422), .B(n57132), .X(n24302) );
  nand_x2_sg U40949 ( .A(n67422), .B(n57138), .X(n23852) );
  nand_x2_sg U40950 ( .A(n67422), .B(n57144), .X(n23592) );
  nand_x2_sg U40951 ( .A(n67422), .B(n57115), .X(n25584) );
  nand_x2_sg U40952 ( .A(n67422), .B(n57127), .X(n24523) );
  inv_x8_sg U40953 ( .A(n23590), .X(n67422) );
  nand_x2_sg U40954 ( .A(n67205), .B(n57124), .X(n24678) );
  nand_x2_sg U40955 ( .A(n67205), .B(n57135), .X(n24253) );
  nand_x2_sg U40956 ( .A(n67205), .B(n57141), .X(n23795) );
  nand_x2_sg U40957 ( .A(n67205), .B(n57147), .X(n23532) );
  nand_x2_sg U40958 ( .A(n67205), .B(n57117), .X(n25342) );
  nand_x2_sg U40959 ( .A(n67205), .B(n57130), .X(n24471) );
  inv_x8_sg U40960 ( .A(n23530), .X(n67205) );
  nand_x2_sg U40961 ( .A(n67231), .B(n24605), .X(n24626) );
  nand_x2_sg U40962 ( .A(n67231), .B(n24163), .X(n24188) );
  nand_x2_sg U40963 ( .A(n67231), .B(n23686), .X(n23717) );
  nand_x2_sg U40964 ( .A(n67231), .B(n23422), .X(n23454) );
  nand_x2_sg U40965 ( .A(n67231), .B(n57117), .X(n24952) );
  nand_x2_sg U40966 ( .A(n67231), .B(n24381), .X(n24406) );
  inv_x8_sg U40967 ( .A(n23452), .X(n67231) );
  nand_x2_sg U40968 ( .A(n67239), .B(n57123), .X(n24610) );
  nand_x2_sg U40969 ( .A(n67239), .B(n57134), .X(n24168) );
  nand_x2_sg U40970 ( .A(n67239), .B(n57140), .X(n23693) );
  nand_x2_sg U40971 ( .A(n67239), .B(n57146), .X(n23430) );
  nand_x2_sg U40972 ( .A(n67239), .B(n57117), .X(n24832) );
  nand_x2_sg U40973 ( .A(n67239), .B(n57129), .X(n24386) );
  inv_x8_sg U40974 ( .A(n23428), .X(n67239) );
  nand_x2_sg U40975 ( .A(n67241), .B(n57124), .X(n24604) );
  nand_x2_sg U40976 ( .A(n67241), .B(n57135), .X(n24162) );
  nand_x2_sg U40977 ( .A(n67241), .B(n57141), .X(n23685) );
  nand_x2_sg U40978 ( .A(n67241), .B(n57147), .X(n23421) );
  nand_x2_sg U40979 ( .A(n67241), .B(n57117), .X(n24793) );
  nand_x2_sg U40980 ( .A(n67241), .B(n57130), .X(n24380) );
  inv_x8_sg U40981 ( .A(n23419), .X(n67241) );
  inv_x4_sg U40982 ( .A(n34131), .X(n68381) );
  nor_x8_sg U40983 ( .A(n67525), .B(n67526), .X(n34131) );
  inv_x4_sg U40984 ( .A(n33266), .X(n68376) );
  nor_x8_sg U40985 ( .A(n67529), .B(n67528), .X(n33266) );
  nor_x8_sg U40986 ( .A(n67537), .B(n57308), .X(n26085) );
  nor_x8_sg U40987 ( .A(n26051), .B(n67537), .X(n26117) );
  inv_x8_sg U40988 ( .A(n57310), .X(n67537) );
  nor_x8_sg U40989 ( .A(n68396), .B(n68390), .X(n29338) );
  nor_x2_sg U40990 ( .A(n32419), .B(n68390), .X(n32418) );
  inv_x8_sg U40991 ( .A(n57306), .X(n68390) );
  inv_x4_sg U40992 ( .A(n47207), .X(n47372) );
  inv_x8_sg U40993 ( .A(n47372), .X(n47373) );
  inv_x8_sg U40994 ( .A(n47373), .X(n67529) );
  inv_x4_sg U40995 ( .A(n47199), .X(n47374) );
  inv_x8_sg U40996 ( .A(n47374), .X(n47375) );
  inv_x8_sg U40997 ( .A(n47375), .X(n67526) );
  nor_x2_sg U40998 ( .A(n23197), .B(n57151), .X(n23189) );
  nor_x2_sg U40999 ( .A(n57025), .B(n57152), .X(n23197) );
  nor_x2_sg U41000 ( .A(n22959), .B(n57157), .X(n22951) );
  nor_x2_sg U41001 ( .A(n57043), .B(n57158), .X(n22959) );
  nor_x2_sg U41002 ( .A(n26181), .B(n68373), .X(n26180) );
  nor_x2_sg U41003 ( .A(n57069), .B(n26215), .X(n26179) );
  nor_x2_sg U41004 ( .A(n24050), .B(n57328), .X(n24049) );
  nand_x2_sg U41005 ( .A(n47327), .B(n57862), .X(n23179) );
  nand_x2_sg U41006 ( .A(n47321), .B(n57862), .X(n23080) );
  nand_x2_sg U41007 ( .A(n47323), .B(n57862), .X(n22941) );
  nand_x2_sg U41008 ( .A(n47325), .B(n57862), .X(n22897) );
  nand_x2_sg U41009 ( .A(n47304), .B(n57862), .X(n22809) );
  nand_x2_sg U41010 ( .A(n67500), .B(n57103), .X(n23936) );
  nor_x2_sg U41011 ( .A(n23938), .B(n57925), .X(n58352) );
  nor_x4_sg U41012 ( .A(n23675), .B(n47313), .X(n23938) );
  nor_x2_sg U41013 ( .A(n58352), .B(n57460), .X(n23933) );
  nor_x2_sg U41014 ( .A(n23806), .B(n23807), .X(n23805) );
  nor_x2_sg U41015 ( .A(n23809), .B(n57925), .X(n58373) );
  nor_x4_sg U41016 ( .A(n23543), .B(n67100), .X(n23809) );
  nor_x2_sg U41017 ( .A(n58373), .B(n57460), .X(n23804) );
  nor_x2_sg U41018 ( .A(n68396), .B(n22445), .X(n22442) );
  nand_x8_sg U41019 ( .A(n57302), .B(n57304), .X(n22445) );
  inv_x2_sg U41020 ( .A(n34174), .X(n68377) );
  inv_x2_sg U41021 ( .A(n33868), .X(n68375) );
  inv_x2_sg U41022 ( .A(n47376), .X(n47377) );
  inv_x2_sg U41023 ( .A(n47378), .X(n47379) );
  inv_x2_sg U41024 ( .A(n47380), .X(n47381) );
  inv_x2_sg U41025 ( .A(n47382), .X(n47383) );
  inv_x2_sg U41026 ( .A(n47384), .X(n47385) );
  inv_x2_sg U41027 ( .A(n47386), .X(n47387) );
  inv_x2_sg U41028 ( .A(n47388), .X(n47389) );
  inv_x2_sg U41029 ( .A(\shifter_0/reg_i_2 [19]), .X(n47612) );
  inv_x2_sg U41030 ( .A(n47390), .X(n47391) );
  nor_x4_sg U41031 ( .A(n32420), .B(n32509), .X(n32377) );
  inv_x2_sg U41032 ( .A(n47392), .X(n47393) );
  inv_x1_sg U41033 ( .A(n25750), .X(n47394) );
  inv_x1_sg U41034 ( .A(n25750), .X(n67463) );
  inv_x1_sg U41035 ( .A(n25238), .X(n47395) );
  inv_x1_sg U41036 ( .A(n25238), .X(n67267) );
  nor_x4_sg U41037 ( .A(n57505), .B(n24695), .X(n24790) );
  nor_x4_sg U41038 ( .A(n47331), .B(n29339), .X(n32440) );
  nor_x4_sg U41039 ( .A(n23675), .B(n68389), .X(n29339) );
  inv_x2_sg U41040 ( .A(n47396), .X(n47397) );
  inv_x2_sg U41041 ( .A(n47398), .X(n47399) );
  inv_x2_sg U41042 ( .A(n47400), .X(n47401) );
  inv_x2_sg U41043 ( .A(n47402), .X(n47403) );
  inv_x2_sg U41044 ( .A(n47404), .X(n47405) );
  inv_x2_sg U41045 ( .A(n47406), .X(n47407) );
  inv_x2_sg U41046 ( .A(n47408), .X(n47409) );
  inv_x2_sg U41047 ( .A(n47410), .X(n47411) );
  inv_x4_sg U41048 ( .A(n47412), .X(n47413) );
  inv_x4_sg U41049 ( .A(n47414), .X(n47415) );
  nor_x4_sg U41050 ( .A(n23543), .B(n68571), .X(n29337) );
  inv_x4_sg U41051 ( .A(n24785), .X(n67523) );
  inv_x8_sg U41052 ( .A(n22546), .X(n68391) );
  inv_x8_sg U41053 ( .A(n23409), .X(n67395) );
  nand_x8_sg U41054 ( .A(n25976), .B(n25977), .X(n23409) );
  inv_x8_sg U41055 ( .A(n23404), .X(n67397) );
  nand_x8_sg U41056 ( .A(n25945), .B(n25946), .X(n23404) );
  inv_x8_sg U41057 ( .A(n23399), .X(n67399) );
  nand_x8_sg U41058 ( .A(n25915), .B(n25916), .X(n23399) );
  inv_x8_sg U41059 ( .A(n23394), .X(n67401) );
  nand_x8_sg U41060 ( .A(n25885), .B(n25886), .X(n23394) );
  inv_x8_sg U41061 ( .A(n23384), .X(n67405) );
  nand_x8_sg U41062 ( .A(n25825), .B(n25826), .X(n23384) );
  inv_x8_sg U41063 ( .A(n23379), .X(n67407) );
  nand_x8_sg U41064 ( .A(n25795), .B(n25796), .X(n23379) );
  inv_x8_sg U41065 ( .A(n23374), .X(n67409) );
  nand_x8_sg U41066 ( .A(n25765), .B(n25766), .X(n23374) );
  inv_x8_sg U41067 ( .A(n23369), .X(n67411) );
  nand_x8_sg U41068 ( .A(n25735), .B(n25736), .X(n23369) );
  inv_x8_sg U41069 ( .A(n23364), .X(n67413) );
  nand_x8_sg U41070 ( .A(n25705), .B(n25706), .X(n23364) );
  inv_x8_sg U41071 ( .A(n23359), .X(n67415) );
  nand_x8_sg U41072 ( .A(n25675), .B(n25676), .X(n23359) );
  inv_x8_sg U41073 ( .A(n23354), .X(n67417) );
  nand_x8_sg U41074 ( .A(n25645), .B(n25646), .X(n23354) );
  inv_x8_sg U41075 ( .A(n23349), .X(n67419) );
  nand_x8_sg U41076 ( .A(n25615), .B(n25616), .X(n23349) );
  inv_x8_sg U41077 ( .A(n23339), .X(n67423) );
  nand_x8_sg U41078 ( .A(n25555), .B(n25556), .X(n23339) );
  inv_x8_sg U41079 ( .A(n23334), .X(n67425) );
  nand_x8_sg U41080 ( .A(n25525), .B(n25526), .X(n23334) );
  inv_x8_sg U41081 ( .A(n23329), .X(n67427) );
  nand_x8_sg U41082 ( .A(n25495), .B(n25496), .X(n23329) );
  inv_x8_sg U41083 ( .A(n23324), .X(n67429) );
  nand_x8_sg U41084 ( .A(n25465), .B(n25466), .X(n23324) );
  inv_x8_sg U41085 ( .A(n23319), .X(n67431) );
  nand_x8_sg U41086 ( .A(n25435), .B(n25436), .X(n23319) );
  inv_x8_sg U41087 ( .A(n23314), .X(n67433) );
  nand_x8_sg U41088 ( .A(n25405), .B(n25406), .X(n23314) );
  inv_x8_sg U41089 ( .A(n23301), .X(n67202) );
  nand_x8_sg U41090 ( .A(n25374), .B(n25375), .X(n23301) );
  inv_x8_sg U41091 ( .A(n23291), .X(n67206) );
  nand_x8_sg U41092 ( .A(n25313), .B(n25314), .X(n23291) );
  inv_x8_sg U41093 ( .A(n23286), .X(n67208) );
  nand_x8_sg U41094 ( .A(n25283), .B(n25284), .X(n23286) );
  inv_x8_sg U41095 ( .A(n23281), .X(n67210) );
  nand_x8_sg U41096 ( .A(n25253), .B(n25254), .X(n23281) );
  inv_x8_sg U41097 ( .A(n23276), .X(n67212) );
  nand_x8_sg U41098 ( .A(n25223), .B(n25224), .X(n23276) );
  inv_x8_sg U41099 ( .A(n23271), .X(n67214) );
  nand_x8_sg U41100 ( .A(n25193), .B(n25194), .X(n23271) );
  inv_x8_sg U41101 ( .A(n23266), .X(n67216) );
  nand_x8_sg U41102 ( .A(n25163), .B(n25164), .X(n23266) );
  inv_x8_sg U41103 ( .A(n23261), .X(n67218) );
  nand_x8_sg U41104 ( .A(n25133), .B(n25134), .X(n23261) );
  inv_x8_sg U41105 ( .A(n23256), .X(n67220) );
  nand_x8_sg U41106 ( .A(n25103), .B(n25104), .X(n23256) );
  inv_x8_sg U41107 ( .A(n23251), .X(n67222) );
  nand_x8_sg U41108 ( .A(n25073), .B(n25074), .X(n23251) );
  inv_x8_sg U41109 ( .A(n23246), .X(n67224) );
  nand_x8_sg U41110 ( .A(n25043), .B(n25044), .X(n23246) );
  inv_x8_sg U41111 ( .A(n23241), .X(n67226) );
  nand_x8_sg U41112 ( .A(n25013), .B(n25014), .X(n23241) );
  inv_x8_sg U41113 ( .A(n23236), .X(n67228) );
  nand_x8_sg U41114 ( .A(n24983), .B(n24984), .X(n23236) );
  inv_x8_sg U41115 ( .A(n23226), .X(n67232) );
  nand_x8_sg U41116 ( .A(n24923), .B(n24924), .X(n23226) );
  inv_x8_sg U41117 ( .A(n23221), .X(n67234) );
  nand_x8_sg U41118 ( .A(n24893), .B(n24894), .X(n23221) );
  inv_x8_sg U41119 ( .A(n23216), .X(n67236) );
  nand_x8_sg U41120 ( .A(n24863), .B(n24864), .X(n23216) );
  inv_x2_sg U41121 ( .A(n68385), .X(n47416) );
  inv_x8_sg U41122 ( .A(n32877), .X(n68385) );
  nor_x4_sg U41123 ( .A(n67524), .B(n68386), .X(n32877) );
  inv_x2_sg U41124 ( .A(n68379), .X(n47417) );
  inv_x8_sg U41125 ( .A(n32922), .X(n68379) );
  nor_x4_sg U41126 ( .A(n68380), .B(n67527), .X(n32922) );
  inv_x4_sg U41127 ( .A(n47355), .X(n61907) );
  inv_x4_sg U41128 ( .A(n39837), .X(n47418) );
  inv_x8_sg U41129 ( .A(n47418), .X(n47419) );
  nor_x8_sg U41130 ( .A(reset), .B(n47419), .X(n38411) );
  inv_x8_sg U41131 ( .A(n68588), .X(n61902) );
  inv_x4_sg U41132 ( .A(n47177), .X(n47420) );
  inv_x4_sg U41133 ( .A(n47173), .X(n47422) );
  inv_x4_sg U41134 ( .A(n47167), .X(n47424) );
  inv_x4_sg U41135 ( .A(n47163), .X(n47426) );
  inv_x4_sg U41136 ( .A(n47033), .X(n47428) );
  inv_x4_sg U41137 ( .A(n47029), .X(n47430) );
  inv_x4_sg U41138 ( .A(n47023), .X(n47432) );
  inv_x4_sg U41139 ( .A(n47019), .X(n47434) );
  inv_x8_sg U41140 ( .A(n22746), .X(n67086) );
  nand_x8_sg U41141 ( .A(n22572), .B(n68589), .X(n22746) );
  inv_x4_sg U41142 ( .A(n47191), .X(n47436) );
  inv_x8_sg U41143 ( .A(n47436), .X(n47437) );
  inv_x4_sg U41144 ( .A(n47217), .X(n47438) );
  inv_x8_sg U41145 ( .A(n47438), .X(n47439) );
  inv_x8_sg U41146 ( .A(n23668), .X(n67396) );
  nor_x8_sg U41147 ( .A(n57918), .B(n67395), .X(n23668) );
  inv_x8_sg U41148 ( .A(n23662), .X(n67398) );
  nor_x8_sg U41149 ( .A(n57918), .B(n67397), .X(n23662) );
  inv_x8_sg U41150 ( .A(n23656), .X(n67400) );
  nor_x8_sg U41151 ( .A(n57918), .B(n67399), .X(n23656) );
  inv_x8_sg U41152 ( .A(n23650), .X(n67402) );
  nor_x8_sg U41153 ( .A(n57918), .B(n67401), .X(n23650) );
  inv_x8_sg U41154 ( .A(n23638), .X(n67406) );
  nor_x8_sg U41155 ( .A(n57918), .B(n67405), .X(n23638) );
  inv_x8_sg U41156 ( .A(n23632), .X(n67408) );
  nor_x8_sg U41157 ( .A(n57918), .B(n67407), .X(n23632) );
  inv_x8_sg U41158 ( .A(n23626), .X(n67410) );
  nor_x8_sg U41159 ( .A(n57918), .B(n67409), .X(n23626) );
  inv_x8_sg U41160 ( .A(n23620), .X(n67412) );
  nor_x8_sg U41161 ( .A(n57918), .B(n67411), .X(n23620) );
  inv_x8_sg U41162 ( .A(n23614), .X(n67414) );
  nor_x8_sg U41163 ( .A(n57918), .B(n67413), .X(n23614) );
  inv_x8_sg U41164 ( .A(n23608), .X(n67416) );
  nor_x8_sg U41165 ( .A(n57918), .B(n67415), .X(n23608) );
  inv_x8_sg U41166 ( .A(n23602), .X(n67418) );
  nor_x8_sg U41167 ( .A(n57918), .B(n67417), .X(n23602) );
  inv_x8_sg U41168 ( .A(n23596), .X(n67420) );
  nor_x8_sg U41169 ( .A(n57918), .B(n67419), .X(n23596) );
  inv_x8_sg U41170 ( .A(n23584), .X(n67424) );
  nor_x8_sg U41171 ( .A(n57918), .B(n67423), .X(n23584) );
  inv_x8_sg U41172 ( .A(n23578), .X(n67426) );
  nor_x8_sg U41173 ( .A(n57918), .B(n67425), .X(n23578) );
  inv_x8_sg U41174 ( .A(n23572), .X(n67428) );
  nor_x8_sg U41175 ( .A(n57918), .B(n67427), .X(n23572) );
  inv_x8_sg U41176 ( .A(n23566), .X(n67430) );
  nor_x8_sg U41177 ( .A(n57918), .B(n67429), .X(n23566) );
  inv_x8_sg U41178 ( .A(n23560), .X(n67432) );
  nor_x8_sg U41179 ( .A(n57918), .B(n67431), .X(n23560) );
  inv_x8_sg U41180 ( .A(n23553), .X(n67434) );
  nor_x8_sg U41181 ( .A(n57918), .B(n67433), .X(n23553) );
  inv_x8_sg U41182 ( .A(n23536), .X(n67203) );
  nor_x8_sg U41183 ( .A(n57918), .B(n67202), .X(n23536) );
  inv_x8_sg U41184 ( .A(n23524), .X(n67207) );
  nor_x8_sg U41185 ( .A(n57918), .B(n67206), .X(n23524) );
  inv_x8_sg U41186 ( .A(n23518), .X(n67209) );
  nor_x8_sg U41187 ( .A(n57918), .B(n67208), .X(n23518) );
  inv_x8_sg U41188 ( .A(n23512), .X(n67211) );
  nor_x8_sg U41189 ( .A(n57918), .B(n67210), .X(n23512) );
  inv_x8_sg U41190 ( .A(n23506), .X(n67213) );
  nor_x8_sg U41191 ( .A(n57918), .B(n67212), .X(n23506) );
  inv_x8_sg U41192 ( .A(n23500), .X(n67215) );
  nor_x8_sg U41193 ( .A(n57918), .B(n67214), .X(n23500) );
  inv_x8_sg U41194 ( .A(n23494), .X(n67217) );
  nor_x8_sg U41195 ( .A(n57918), .B(n67216), .X(n23494) );
  inv_x8_sg U41196 ( .A(n23488), .X(n67219) );
  nor_x8_sg U41197 ( .A(n57919), .B(n67218), .X(n23488) );
  inv_x8_sg U41198 ( .A(n23482), .X(n67221) );
  nor_x8_sg U41199 ( .A(n57918), .B(n67220), .X(n23482) );
  inv_x8_sg U41200 ( .A(n23476), .X(n67223) );
  nor_x8_sg U41201 ( .A(n57919), .B(n67222), .X(n23476) );
  inv_x8_sg U41202 ( .A(n23470), .X(n67225) );
  nor_x8_sg U41203 ( .A(n57918), .B(n67224), .X(n23470) );
  inv_x8_sg U41204 ( .A(n23464), .X(n67227) );
  nor_x8_sg U41205 ( .A(n57919), .B(n67226), .X(n23464) );
  inv_x8_sg U41206 ( .A(n23458), .X(n67229) );
  nor_x8_sg U41207 ( .A(n57918), .B(n67228), .X(n23458) );
  inv_x8_sg U41208 ( .A(n23446), .X(n67233) );
  nor_x8_sg U41209 ( .A(n57918), .B(n67232), .X(n23446) );
  inv_x8_sg U41210 ( .A(n23440), .X(n67235) );
  nor_x8_sg U41211 ( .A(n57918), .B(n67234), .X(n23440) );
  inv_x8_sg U41212 ( .A(n23434), .X(n67237) );
  nor_x8_sg U41213 ( .A(n57918), .B(n67236), .X(n23434) );
  nor_x2_sg U41214 ( .A(n57097), .B(n68573), .X(n23806) );
  nor_x4_sg U41215 ( .A(n23543), .B(n68573), .X(n24050) );
  nand_x4_sg U41216 ( .A(n68573), .B(n68571), .X(n31973) );
  inv_x8_sg U41217 ( .A(n22521), .X(n68573) );
  inv_x4_sg U41218 ( .A(n47205), .X(n47440) );
  inv_x8_sg U41219 ( .A(n47440), .X(n47441) );
  nor_x8_sg U41220 ( .A(n47373), .B(n47441), .X(n34174) );
  nor_x8_sg U41221 ( .A(n67529), .B(n47441), .X(n33868) );
  inv_x4_sg U41222 ( .A(n47197), .X(n47442) );
  inv_x8_sg U41223 ( .A(n47442), .X(n47443) );
  nor_x8_sg U41224 ( .A(n47375), .B(n47443), .X(n33998) );
  nor_x8_sg U41225 ( .A(n67526), .B(n47443), .X(n34086) );
  inv_x8_sg U41226 ( .A(n23416), .X(n67500) );
  nand_x4_sg U41227 ( .A(n23416), .B(n22497), .X(n24785) );
  nor_x8_sg U41228 ( .A(n57304), .B(n57302), .X(n23416) );
  inv_x4_sg U41229 ( .A(n26043), .X(n68374) );
  nor_x8_sg U41230 ( .A(n26047), .B(n67537), .X(n26043) );
  nor_x8_sg U41231 ( .A(n57918), .B(n67403), .X(n23644) );
  inv_x8_sg U41232 ( .A(n23389), .X(n67403) );
  nor_x8_sg U41233 ( .A(n57918), .B(n67421), .X(n23590) );
  inv_x8_sg U41234 ( .A(n23344), .X(n67421) );
  nor_x8_sg U41235 ( .A(n57918), .B(n67204), .X(n23530) );
  inv_x8_sg U41236 ( .A(n23296), .X(n67204) );
  nor_x8_sg U41237 ( .A(n57918), .B(n67230), .X(n23452) );
  inv_x8_sg U41238 ( .A(n23231), .X(n67230) );
  nor_x8_sg U41239 ( .A(n57919), .B(n67238), .X(n23428) );
  inv_x8_sg U41240 ( .A(n23211), .X(n67238) );
  nor_x8_sg U41241 ( .A(n57919), .B(n67240), .X(n23419) );
  inv_x8_sg U41242 ( .A(n23206), .X(n67240) );
  nor_x8_sg U41243 ( .A(n67525), .B(n47375), .X(n34219) );
  inv_x8_sg U41244 ( .A(n47443), .X(n67525) );
  nor_x8_sg U41245 ( .A(n67528), .B(n47373), .X(n33738) );
  inv_x8_sg U41246 ( .A(n47441), .X(n67528) );
  inv_x4_sg U41247 ( .A(n47187), .X(n47444) );
  inv_x8_sg U41248 ( .A(n47444), .X(n47445) );
  inv_x8_sg U41249 ( .A(n47445), .X(n68396) );
  nand_x1_sg U41250 ( .A(n26325), .B(n67573), .X(n26324) );
  inv_x1_sg U41251 ( .A(n26326), .X(n67573) );
  nor_x1_sg U41252 ( .A(n26295), .B(n67566), .X(n26286) );
  inv_x1_sg U41253 ( .A(n26287), .X(n67568) );
  nor_x1_sg U41254 ( .A(n68227), .B(n51557), .X(n35848) );
  inv_x2_sg U41255 ( .A(n51556), .X(n51557) );
  inv_x1_sg U41256 ( .A(n38407), .X(n51556) );
  nor_x1_sg U41257 ( .A(n68272), .B(state[1]), .X(n38407) );
  nand_x1_sg U41258 ( .A(n26334), .B(n26335), .X(n26333) );
  nand_x1_sg U41259 ( .A(n26323), .B(n26324), .X(n26322) );
  inv_x1_sg U41260 ( .A(n26310), .X(n67570) );
  inv_x1_sg U41261 ( .A(n26274), .X(n67565) );
  nand_x1_sg U41262 ( .A(n61911), .B(n61907), .X(n30626) );
  inv_x1_sg U41263 ( .A(n35848), .X(n51554) );
  nor_x1_sg U41264 ( .A(n57460), .B(n58472), .X(n58473) );
  nor_x1_sg U41265 ( .A(n57460), .B(n58430), .X(n58431) );
  inv_x1_sg U41266 ( .A(n26142), .X(n67563) );
  inv_x1_sg U41267 ( .A(n26103), .X(n67557) );
  inv_x1_sg U41268 ( .A(n26234), .X(n67551) );
  inv_x1_sg U41269 ( .A(n26200), .X(n67545) );
  nor_x1_sg U41270 ( .A(n67569), .B(n26300), .X(n26299) );
  nand_x1_sg U41271 ( .A(n26264), .B(n26265), .X(n26263) );
  nand_x1_sg U41272 ( .A(n58625), .B(n58624), .X(n58626) );
  nand_x1_sg U41273 ( .A(n32087), .B(n57924), .X(n58624) );
  nand_x1_sg U41274 ( .A(n32079), .B(n57927), .X(n58625) );
  inv_x1_sg U41275 ( .A(n58623), .X(n58628) );
  nand_x2_sg U41276 ( .A(n32240), .B(n32241), .X(n32087) );
  nor_x1_sg U41277 ( .A(n30625), .B(n46855), .X(n29328) );
  nand_x1_sg U41278 ( .A(n58591), .B(n58590), .X(n58592) );
  nand_x1_sg U41279 ( .A(n32532), .B(n57924), .X(n58590) );
  nand_x1_sg U41280 ( .A(n32524), .B(n57928), .X(n58591) );
  inv_x1_sg U41281 ( .A(n58589), .X(n58594) );
  nand_x2_sg U41282 ( .A(n32685), .B(n32686), .X(n32532) );
  nand_x1_sg U41283 ( .A(n24047), .B(n57459), .X(n24046) );
  nand_x1_sg U41284 ( .A(n24157), .B(n57459), .X(n24156) );
  nand_x1_sg U41285 ( .A(n26155), .B(n26156), .X(n26154) );
  inv_x1_sg U41286 ( .A(n26128), .X(n67560) );
  nand_x1_sg U41287 ( .A(n26119), .B(n26120), .X(n26118) );
  inv_x1_sg U41288 ( .A(n26086), .X(n67554) );
  nand_x1_sg U41289 ( .A(n26247), .B(n26248), .X(n26246) );
  inv_x1_sg U41290 ( .A(n26220), .X(n67548) );
  nand_x1_sg U41291 ( .A(n26213), .B(n26214), .X(n26212) );
  inv_x1_sg U41292 ( .A(n26186), .X(n67542) );
  nand_x1_sg U41293 ( .A(n26298), .B(n26299), .X(n26297) );
  nand_x1_sg U41294 ( .A(n57862), .B(n32082), .X(n32297) );
  nand_x1_sg U41295 ( .A(n57858), .B(n32078), .X(n32296) );
  nand_x1_sg U41296 ( .A(n32089), .B(n57864), .X(n32334) );
  nand_x1_sg U41297 ( .A(n58629), .B(n47505), .X(n58631) );
  nand_x1_sg U41298 ( .A(n58628), .B(n58627), .X(n58629) );
  nand_x1_sg U41299 ( .A(n58626), .B(n57296), .X(n58627) );
  nand_x2_sg U41300 ( .A(n32298), .B(n32299), .X(n32082) );
  inv_x1_sg U41301 ( .A(n32087), .X(n68565) );
  nand_x1_sg U41302 ( .A(n29332), .B(n32527), .X(n32742) );
  nand_x1_sg U41303 ( .A(n57858), .B(n32523), .X(n32741) );
  nand_x1_sg U41304 ( .A(n32534), .B(n57864), .X(n32779) );
  nand_x1_sg U41305 ( .A(n58595), .B(n57917), .X(n58596) );
  nand_x1_sg U41306 ( .A(n58594), .B(n58593), .X(n58595) );
  nand_x1_sg U41307 ( .A(n58592), .B(n53715), .X(n58593) );
  nand_x2_sg U41308 ( .A(n32743), .B(n32744), .X(n32527) );
  inv_x1_sg U41309 ( .A(n32532), .X(n68472) );
  inv_x2_sg U41310 ( .A(n35709), .X(n47572) );
  nor_x1_sg U41311 ( .A(n35839), .B(n35705), .X(n35709) );
  inv_x1_sg U41312 ( .A(n22420), .X(n58584) );
  inv_x1_sg U41313 ( .A(n22444), .X(n58582) );
  nand_x1_sg U41314 ( .A(n22570), .B(n22571), .X(n22569) );
  nand_x1_sg U41315 ( .A(n22596), .B(n22597), .X(n22595) );
  nand_x1_sg U41316 ( .A(n22621), .B(n22622), .X(n22620) );
  nand_x1_sg U41317 ( .A(n22648), .B(n22649), .X(n22647) );
  nor_x1_sg U41318 ( .A(n57919), .B(n67099), .X(n23205) );
  nor_x1_sg U41319 ( .A(n67099), .B(n57917), .X(n23204) );
  nor_x1_sg U41320 ( .A(n57919), .B(n67502), .X(n23313) );
  nor_x1_sg U41321 ( .A(n67502), .B(n57920), .X(n23312) );
  nand_x1_sg U41322 ( .A(n23549), .B(n57928), .X(n58383) );
  nand_x1_sg U41323 ( .A(n23680), .B(n57928), .X(n58378) );
  nor_x1_sg U41324 ( .A(n57918), .B(n67098), .X(n23946) );
  nor_x1_sg U41325 ( .A(n67098), .B(n47505), .X(n23944) );
  nor_x1_sg U41326 ( .A(n57919), .B(n67501), .X(n24056) );
  nor_x1_sg U41327 ( .A(n67501), .B(n57920), .X(n24054) );
  nand_x1_sg U41328 ( .A(n57923), .B(n57100), .X(n58127) );
  nor_x1_sg U41329 ( .A(n24597), .B(n46889), .X(n58129) );
  nand_x1_sg U41330 ( .A(n24689), .B(n24690), .X(n24688) );
  nand_x1_sg U41331 ( .A(n24783), .B(n24784), .X(n24782) );
  inv_x1_sg U41332 ( .A(n26154), .X(n67559) );
  inv_x1_sg U41333 ( .A(n26118), .X(n67553) );
  inv_x1_sg U41334 ( .A(n26246), .X(n67547) );
  inv_x1_sg U41335 ( .A(n26212), .X(n67541) );
  nor_x1_sg U41336 ( .A(n32067), .B(n57100), .X(n32093) );
  nand_x1_sg U41337 ( .A(n58637), .B(n58636), .X(n32172) );
  inv_x1_sg U41338 ( .A(n58635), .X(n58636) );
  nand_x1_sg U41339 ( .A(n31961), .B(n57349), .X(n58637) );
  nor_x1_sg U41340 ( .A(n57100), .B(n68514), .X(n32066) );
  nand_x1_sg U41341 ( .A(n58647), .B(n58646), .X(n32068) );
  inv_x1_sg U41342 ( .A(n58645), .X(n58646) );
  nand_x1_sg U41343 ( .A(n68541), .B(n57862), .X(n32080) );
  inv_x1_sg U41344 ( .A(n32082), .X(n68541) );
  nand_x1_sg U41345 ( .A(n68551), .B(n57345), .X(n32085) );
  nand_x1_sg U41346 ( .A(n68565), .B(n29329), .X(n32086) );
  inv_x1_sg U41347 ( .A(n32088), .X(n68551) );
  inv_x1_sg U41348 ( .A(n31962), .X(n68535) );
  nand_x1_sg U41349 ( .A(n57857), .B(n31961), .X(n31960) );
  nand_x4_sg U41350 ( .A(n32136), .B(n32137), .X(n31943) );
  nor_x1_sg U41351 ( .A(n32146), .B(n32147), .X(n32136) );
  nor_x1_sg U41352 ( .A(n32138), .B(n32139), .X(n32137) );
  nand_x4_sg U41353 ( .A(n32154), .B(n32155), .X(n31947) );
  nor_x1_sg U41354 ( .A(n32164), .B(n32165), .X(n32154) );
  nor_x1_sg U41355 ( .A(n32156), .B(n32157), .X(n32155) );
  nand_x4_sg U41356 ( .A(n32098), .B(n32099), .X(n31933) );
  nor_x1_sg U41357 ( .A(n32108), .B(n32109), .X(n32098) );
  nor_x1_sg U41358 ( .A(n32100), .B(n32101), .X(n32099) );
  nand_x4_sg U41359 ( .A(n32116), .B(n32117), .X(n31937) );
  nor_x1_sg U41360 ( .A(n32126), .B(n32127), .X(n32116) );
  nor_x1_sg U41361 ( .A(n32118), .B(n32119), .X(n32117) );
  nand_x1_sg U41362 ( .A(n32021), .B(n32022), .X(n32020) );
  nor_x1_sg U41363 ( .A(n32031), .B(n32032), .X(n32021) );
  nor_x1_sg U41364 ( .A(n32023), .B(n32024), .X(n32022) );
  nand_x1_sg U41365 ( .A(n32042), .B(n32043), .X(n32041) );
  nor_x1_sg U41366 ( .A(n32053), .B(n32054), .X(n32042) );
  nor_x1_sg U41367 ( .A(n57100), .B(n68425), .X(n32512) );
  nand_x1_sg U41368 ( .A(n58608), .B(n58607), .X(n32514) );
  inv_x1_sg U41369 ( .A(n58606), .X(n58607) );
  nor_x1_sg U41370 ( .A(n32513), .B(n57100), .X(n32538) );
  nand_x1_sg U41371 ( .A(n58602), .B(n58601), .X(n32617) );
  inv_x1_sg U41372 ( .A(n58600), .X(n58601) );
  nand_x1_sg U41373 ( .A(n32428), .B(n57349), .X(n58602) );
  nand_x1_sg U41374 ( .A(n68448), .B(n57862), .X(n32525) );
  inv_x1_sg U41375 ( .A(n32527), .X(n68448) );
  nand_x1_sg U41376 ( .A(n68458), .B(n57347), .X(n32530) );
  nand_x1_sg U41377 ( .A(n68472), .B(n57865), .X(n32531) );
  inv_x1_sg U41378 ( .A(n32533), .X(n68458) );
  inv_x1_sg U41379 ( .A(n32429), .X(n68442) );
  nand_x1_sg U41380 ( .A(n57857), .B(n32428), .X(n32427) );
  nand_x4_sg U41381 ( .A(n32581), .B(n32582), .X(n32411) );
  nor_x1_sg U41382 ( .A(n32591), .B(n32592), .X(n32581) );
  nor_x1_sg U41383 ( .A(n32583), .B(n32584), .X(n32582) );
  nand_x4_sg U41384 ( .A(n32599), .B(n32600), .X(n32415) );
  nor_x1_sg U41385 ( .A(n32609), .B(n32610), .X(n32599) );
  nor_x1_sg U41386 ( .A(n32601), .B(n32602), .X(n32600) );
  nand_x4_sg U41387 ( .A(n32543), .B(n32544), .X(n32401) );
  nor_x1_sg U41388 ( .A(n32553), .B(n32554), .X(n32543) );
  nor_x1_sg U41389 ( .A(n32545), .B(n32546), .X(n32544) );
  nand_x4_sg U41390 ( .A(n32561), .B(n32562), .X(n32405) );
  nor_x1_sg U41391 ( .A(n32571), .B(n32572), .X(n32561) );
  nor_x1_sg U41392 ( .A(n32563), .B(n32564), .X(n32562) );
  nand_x1_sg U41393 ( .A(n32463), .B(n32464), .X(n32462) );
  nor_x1_sg U41394 ( .A(n32473), .B(n32474), .X(n32463) );
  nor_x1_sg U41395 ( .A(n32465), .B(n32466), .X(n32464) );
  nor_x1_sg U41396 ( .A(n32496), .B(n32497), .X(n32485) );
  nand_x1_sg U41397 ( .A(n58585), .B(n58584), .X(n58586) );
  nand_x1_sg U41398 ( .A(n58585), .B(n58582), .X(n58583) );
  inv_x1_sg U41399 ( .A(n47521), .X(n47474) );
  inv_x1_sg U41400 ( .A(n56675), .X(n47446) );
  inv_x1_sg U41401 ( .A(n56721), .X(n47476) );
  inv_x1_sg U41402 ( .A(n56677), .X(n47482) );
  inv_x1_sg U41403 ( .A(n51215), .X(n47454) );
  inv_x1_sg U41404 ( .A(n56811), .X(n47486) );
  inv_x1_sg U41405 ( .A(n51365), .X(n47466) );
  inv_x1_sg U41406 ( .A(n56763), .X(n47462) );
  inv_x1_sg U41407 ( .A(n51305), .X(n47452) );
  inv_x1_sg U41408 ( .A(n56765), .X(n47494) );
  inv_x1_sg U41409 ( .A(n51419), .X(n47472) );
  inv_x1_sg U41410 ( .A(n56855), .X(n47488) );
  inv_x1_sg U41411 ( .A(n51325), .X(n47464) );
  inv_x1_sg U41412 ( .A(n47537), .X(n47448) );
  inv_x1_sg U41413 ( .A(n56741), .X(n47456) );
  inv_x1_sg U41414 ( .A(n56791), .X(n47478) );
  inv_x1_sg U41415 ( .A(n51343), .X(n47468) );
  inv_x1_sg U41416 ( .A(n47541), .X(n47450) );
  inv_x1_sg U41417 ( .A(n56743), .X(n47484) );
  inv_x1_sg U41418 ( .A(n51279), .X(n47458) );
  inv_x1_sg U41419 ( .A(n56795), .X(n47480) );
  inv_x1_sg U41420 ( .A(n51347), .X(n47470) );
  inv_x1_sg U41421 ( .A(n56747), .X(n47492) );
  inv_x1_sg U41422 ( .A(n51283), .X(n47460) );
  nand_x1_sg U41423 ( .A(n57922), .B(n58375), .X(n58331) );
  nand_x1_sg U41424 ( .A(n57922), .B(n58372), .X(n58326) );
  nand_x1_sg U41425 ( .A(n57922), .B(n58371), .X(n58321) );
  nand_x1_sg U41426 ( .A(n57922), .B(n58370), .X(n58315) );
  nand_x1_sg U41427 ( .A(n57922), .B(n58369), .X(n58310) );
  nand_x1_sg U41428 ( .A(n57923), .B(n58368), .X(n58306) );
  nand_x1_sg U41429 ( .A(n57922), .B(n58367), .X(n58301) );
  nand_x1_sg U41430 ( .A(n57922), .B(n58366), .X(n58296) );
  nand_x1_sg U41431 ( .A(n57924), .B(n58365), .X(n58290) );
  nand_x1_sg U41432 ( .A(n57924), .B(n58364), .X(n58285) );
  nand_x1_sg U41433 ( .A(n57923), .B(n58363), .X(n58281) );
  nand_x1_sg U41434 ( .A(n57924), .B(n58362), .X(n58276) );
  nand_x1_sg U41435 ( .A(n57924), .B(n58361), .X(n58270) );
  nand_x1_sg U41436 ( .A(n57924), .B(n58360), .X(n58265) );
  nand_x1_sg U41437 ( .A(n57922), .B(n58359), .X(n58261) );
  nand_x1_sg U41438 ( .A(n53717), .B(n58358), .X(n58256) );
  nand_x1_sg U41439 ( .A(n57923), .B(n58357), .X(n58251) );
  nand_x1_sg U41440 ( .A(n57923), .B(n58356), .X(n58245) );
  nand_x1_sg U41441 ( .A(n57924), .B(n58355), .X(n58240) );
  nand_x1_sg U41442 ( .A(n57923), .B(n58354), .X(n58236) );
  nand_x1_sg U41443 ( .A(n57923), .B(n58353), .X(n58231) );
  nand_x1_sg U41444 ( .A(n57923), .B(n58351), .X(n58226) );
  nand_x1_sg U41445 ( .A(n57924), .B(n58350), .X(n58221) );
  nand_x1_sg U41446 ( .A(n57923), .B(n58349), .X(n58215) );
  nand_x1_sg U41447 ( .A(n57923), .B(n58348), .X(n58210) );
  nand_x1_sg U41448 ( .A(n57923), .B(n58347), .X(n58206) );
  nand_x1_sg U41449 ( .A(n57924), .B(n58346), .X(n58201) );
  nand_x1_sg U41450 ( .A(n57923), .B(n58345), .X(n58196) );
  nand_x1_sg U41451 ( .A(n57924), .B(n58344), .X(n58190) );
  nand_x1_sg U41452 ( .A(n57923), .B(n58343), .X(n58185) );
  nand_x1_sg U41453 ( .A(n57924), .B(n58342), .X(n58181) );
  nand_x1_sg U41454 ( .A(n57923), .B(n58341), .X(n58176) );
  nand_x1_sg U41455 ( .A(n57924), .B(n58340), .X(n58170) );
  nand_x1_sg U41456 ( .A(n57923), .B(n58339), .X(n58165) );
  nand_x1_sg U41457 ( .A(n57923), .B(n58338), .X(n58161) );
  nand_x1_sg U41458 ( .A(n57923), .B(n58337), .X(n58156) );
  nand_x1_sg U41459 ( .A(n57923), .B(n58336), .X(n58151) );
  nand_x1_sg U41460 ( .A(n57923), .B(n58335), .X(n58145) );
  nand_x1_sg U41461 ( .A(n57923), .B(n58334), .X(n58140) );
  nand_x1_sg U41462 ( .A(n57923), .B(n58333), .X(n58136) );
  nand_x1_sg U41463 ( .A(n24266), .B(n57322), .X(n24263) );
  nand_x4_sg U41464 ( .A(n57918), .B(n24371), .X(n24368) );
  nand_x1_sg U41465 ( .A(n24372), .B(n24373), .X(n24371) );
  nand_x1_sg U41466 ( .A(n24375), .B(n57322), .X(n24372) );
  nand_x1_sg U41467 ( .A(n58132), .B(n58131), .X(n24481) );
  nand_x1_sg U41468 ( .A(n57100), .B(n24688), .X(n24686) );
  nand_x1_sg U41469 ( .A(n57100), .B(n24782), .X(n24780) );
  nand_x1_sg U41470 ( .A(n24383), .B(n57311), .X(n24817) );
  nand_x1_sg U41471 ( .A(n57311), .B(n24388), .X(n24849) );
  nand_x1_sg U41472 ( .A(n57311), .B(n24393), .X(n24879) );
  nand_x1_sg U41473 ( .A(n57311), .B(n24398), .X(n24909) );
  nand_x1_sg U41474 ( .A(n57311), .B(n24403), .X(n24939) );
  nand_x1_sg U41475 ( .A(n57311), .B(n24408), .X(n24969) );
  nand_x1_sg U41476 ( .A(n57311), .B(n24413), .X(n24999) );
  nand_x1_sg U41477 ( .A(n57311), .B(n24418), .X(n25029) );
  nand_x1_sg U41478 ( .A(n57311), .B(n24423), .X(n25059) );
  nand_x1_sg U41479 ( .A(n57311), .B(n24428), .X(n25089) );
  nand_x1_sg U41480 ( .A(n57311), .B(n24433), .X(n25119) );
  nand_x1_sg U41481 ( .A(n57311), .B(n24438), .X(n25149) );
  nand_x1_sg U41482 ( .A(n57311), .B(n24443), .X(n25179) );
  nand_x1_sg U41483 ( .A(n57311), .B(n24448), .X(n25209) );
  nand_x1_sg U41484 ( .A(n57311), .B(n24453), .X(n25239) );
  nand_x1_sg U41485 ( .A(n57311), .B(n24458), .X(n25269) );
  nand_x1_sg U41486 ( .A(n57311), .B(n24463), .X(n25299) );
  nand_x1_sg U41487 ( .A(n57311), .B(n24468), .X(n25329) );
  nand_x1_sg U41488 ( .A(n57311), .B(n24473), .X(n25359) );
  nand_x1_sg U41489 ( .A(n57311), .B(n24489), .X(n25390) );
  nand_x1_sg U41490 ( .A(n57311), .B(n24495), .X(n25421) );
  nand_x1_sg U41491 ( .A(n57311), .B(n24500), .X(n25451) );
  nand_x1_sg U41492 ( .A(n57311), .B(n24505), .X(n25481) );
  nand_x1_sg U41493 ( .A(n57311), .B(n24510), .X(n25511) );
  nand_x1_sg U41494 ( .A(n57311), .B(n24515), .X(n25541) );
  nand_x1_sg U41495 ( .A(n57311), .B(n24520), .X(n25571) );
  nand_x1_sg U41496 ( .A(n57311), .B(n24525), .X(n25601) );
  nand_x1_sg U41497 ( .A(n57311), .B(n24530), .X(n25631) );
  nand_x1_sg U41498 ( .A(n57311), .B(n24535), .X(n25661) );
  nand_x1_sg U41499 ( .A(n57311), .B(n24540), .X(n25691) );
  nand_x1_sg U41500 ( .A(n57311), .B(n24545), .X(n25721) );
  nand_x1_sg U41501 ( .A(n57311), .B(n24550), .X(n25751) );
  nand_x1_sg U41502 ( .A(n57313), .B(n24555), .X(n25781) );
  nand_x1_sg U41503 ( .A(n57311), .B(n24560), .X(n25811) );
  nand_x1_sg U41504 ( .A(n57311), .B(n24565), .X(n25841) );
  nand_x1_sg U41505 ( .A(n57311), .B(n24570), .X(n25871) );
  nand_x1_sg U41506 ( .A(n57311), .B(n24575), .X(n25901) );
  nand_x1_sg U41507 ( .A(n57311), .B(n24580), .X(n25931) );
  nand_x1_sg U41508 ( .A(n57311), .B(n24585), .X(n25961) );
  nand_x1_sg U41509 ( .A(n57311), .B(n24601), .X(n25992) );
  nand_x1_sg U41510 ( .A(n57455), .B(n32172), .X(n32091) );
  nand_x1_sg U41511 ( .A(n32093), .B(n57918), .X(n32092) );
  nand_x1_sg U41512 ( .A(n57454), .B(n32068), .X(n32064) );
  nand_x1_sg U41513 ( .A(n32066), .B(n57918), .X(n32065) );
  nand_x1_sg U41514 ( .A(n68496), .B(n57857), .X(n31954) );
  inv_x1_sg U41515 ( .A(n58654), .X(n31964) );
  nand_x1_sg U41516 ( .A(n57300), .B(n31943), .X(n31942) );
  inv_x1_sg U41517 ( .A(n31944), .X(n68524) );
  nand_x1_sg U41518 ( .A(n57300), .B(n31947), .X(n31946) );
  inv_x1_sg U41519 ( .A(n31948), .X(n68515) );
  nand_x1_sg U41520 ( .A(n57300), .B(n31933), .X(n31932) );
  inv_x1_sg U41521 ( .A(n31934), .X(n68534) );
  nand_x1_sg U41522 ( .A(n47415), .B(n31937), .X(n31936) );
  inv_x1_sg U41523 ( .A(n31938), .X(n68529) );
  nand_x4_sg U41524 ( .A(n58652), .B(n58651), .X(n31995) );
  nand_x1_sg U41525 ( .A(n32001), .B(n57924), .X(n58652) );
  nand_x1_sg U41526 ( .A(n32020), .B(n57925), .X(n58651) );
  nand_x1_sg U41527 ( .A(n32002), .B(n32003), .X(n32001) );
  inv_x2_sg U41528 ( .A(n31992), .X(n47490) );
  nor_x1_sg U41529 ( .A(n68267), .B(n61909), .X(n31992) );
  nand_x1_sg U41530 ( .A(n57454), .B(n32514), .X(n32510) );
  nand_x1_sg U41531 ( .A(n32512), .B(n57919), .X(n32511) );
  nand_x1_sg U41532 ( .A(n57455), .B(n32617), .X(n32536) );
  nand_x1_sg U41533 ( .A(n32538), .B(n57918), .X(n32537) );
  nand_x1_sg U41534 ( .A(n68407), .B(n57857), .X(n32422) );
  inv_x1_sg U41535 ( .A(n58619), .X(n32431) );
  nand_x1_sg U41536 ( .A(n47413), .B(n32411), .X(n32410) );
  inv_x1_sg U41537 ( .A(n32412), .X(n68393) );
  nand_x1_sg U41538 ( .A(n57306), .B(n32415), .X(n32414) );
  inv_x1_sg U41539 ( .A(n32416), .X(n68392) );
  nand_x1_sg U41540 ( .A(n57306), .B(n32401), .X(n32400) );
  inv_x1_sg U41541 ( .A(n32402), .X(n68395) );
  nand_x1_sg U41542 ( .A(n57306), .B(n32405), .X(n32404) );
  inv_x1_sg U41543 ( .A(n32406), .X(n68394) );
  nand_x4_sg U41544 ( .A(n58615), .B(n58614), .X(n32437) );
  nand_x1_sg U41545 ( .A(n32443), .B(n57924), .X(n58615) );
  nand_x1_sg U41546 ( .A(n32462), .B(n57925), .X(n58614) );
  nand_x1_sg U41547 ( .A(n32444), .B(n32445), .X(n32443) );
  nand_x1_sg U41548 ( .A(n32485), .B(n32486), .X(n32483) );
  inv_x1_sg U41549 ( .A(n58579), .X(n58580) );
  inv_x1_sg U41550 ( .A(n58577), .X(n58578) );
  inv_x1_sg U41551 ( .A(n58574), .X(n58575) );
  inv_x1_sg U41552 ( .A(n58572), .X(n58573) );
  inv_x1_sg U41553 ( .A(n58570), .X(n58571) );
  inv_x1_sg U41554 ( .A(n58567), .X(n58568) );
  inv_x1_sg U41555 ( .A(n58565), .X(n58566) );
  inv_x1_sg U41556 ( .A(n58563), .X(n58564) );
  inv_x1_sg U41557 ( .A(n58560), .X(n58561) );
  inv_x1_sg U41558 ( .A(n58558), .X(n58559) );
  inv_x1_sg U41559 ( .A(n58556), .X(n58557) );
  inv_x1_sg U41560 ( .A(n58553), .X(n58554) );
  inv_x1_sg U41561 ( .A(n58551), .X(n58552) );
  inv_x1_sg U41562 ( .A(n58549), .X(n58550) );
  inv_x1_sg U41563 ( .A(n58546), .X(n58547) );
  inv_x1_sg U41564 ( .A(n58543), .X(n58544) );
  inv_x1_sg U41565 ( .A(n58540), .X(n58541) );
  inv_x1_sg U41566 ( .A(n58538), .X(n58539) );
  inv_x1_sg U41567 ( .A(n58536), .X(n58537) );
  inv_x1_sg U41568 ( .A(n58533), .X(n58534) );
  inv_x1_sg U41569 ( .A(n58530), .X(n58531) );
  inv_x1_sg U41570 ( .A(n58528), .X(n58529) );
  inv_x1_sg U41571 ( .A(n58525), .X(n58526) );
  inv_x1_sg U41572 ( .A(n58523), .X(n58524) );
  inv_x1_sg U41573 ( .A(n58521), .X(n58522) );
  inv_x1_sg U41574 ( .A(n58518), .X(n58519) );
  inv_x1_sg U41575 ( .A(n58516), .X(n58517) );
  inv_x1_sg U41576 ( .A(n58514), .X(n58515) );
  inv_x1_sg U41577 ( .A(n58511), .X(n58512) );
  inv_x1_sg U41578 ( .A(n58509), .X(n58510) );
  inv_x1_sg U41579 ( .A(n58507), .X(n58508) );
  inv_x1_sg U41580 ( .A(n58504), .X(n58505) );
  inv_x1_sg U41581 ( .A(n58502), .X(n58503) );
  inv_x1_sg U41582 ( .A(n58500), .X(n58501) );
  inv_x1_sg U41583 ( .A(n58497), .X(n58498) );
  inv_x1_sg U41584 ( .A(n58494), .X(n58495) );
  inv_x1_sg U41585 ( .A(n58491), .X(n58492) );
  inv_x1_sg U41586 ( .A(n58489), .X(n58490) );
  inv_x1_sg U41587 ( .A(n58487), .X(n58488) );
  inv_x1_sg U41588 ( .A(n58485), .X(n58486) );
  nand_x1_sg U41589 ( .A(n58375), .B(n57314), .X(n23687) );
  nand_x1_sg U41590 ( .A(n57314), .B(n58372), .X(n23694) );
  nand_x1_sg U41591 ( .A(n57314), .B(n58371), .X(n23700) );
  nand_x1_sg U41592 ( .A(n57314), .B(n58370), .X(n23706) );
  nand_x1_sg U41593 ( .A(n57314), .B(n58369), .X(n23712) );
  nand_x1_sg U41594 ( .A(n57314), .B(n58368), .X(n23718) );
  nand_x1_sg U41595 ( .A(n57314), .B(n58367), .X(n23724) );
  nand_x1_sg U41596 ( .A(n57314), .B(n58366), .X(n23730) );
  nand_x1_sg U41597 ( .A(n57314), .B(n58365), .X(n23736) );
  nand_x1_sg U41598 ( .A(n57314), .B(n58364), .X(n23742) );
  nand_x1_sg U41599 ( .A(n57314), .B(n58363), .X(n23748) );
  nand_x1_sg U41600 ( .A(n57314), .B(n58362), .X(n23754) );
  nand_x1_sg U41601 ( .A(n57314), .B(n58361), .X(n23760) );
  nand_x1_sg U41602 ( .A(n57314), .B(n58360), .X(n23766) );
  nand_x1_sg U41603 ( .A(n57314), .B(n58359), .X(n23772) );
  nand_x1_sg U41604 ( .A(n57314), .B(n58358), .X(n23778) );
  nand_x1_sg U41605 ( .A(n57314), .B(n58357), .X(n23784) );
  nand_x1_sg U41606 ( .A(n57314), .B(n58356), .X(n23790) );
  nand_x1_sg U41607 ( .A(n57314), .B(n58355), .X(n23796) );
  nand_x1_sg U41608 ( .A(n57314), .B(n58354), .X(n23810) );
  nand_x1_sg U41609 ( .A(n57314), .B(n58353), .X(n23817) );
  nand_x1_sg U41610 ( .A(n57314), .B(n58351), .X(n23823) );
  nand_x1_sg U41611 ( .A(n57314), .B(n58350), .X(n23829) );
  nand_x1_sg U41612 ( .A(n57314), .B(n58349), .X(n23835) );
  nand_x1_sg U41613 ( .A(n57314), .B(n58348), .X(n23841) );
  nand_x1_sg U41614 ( .A(n57314), .B(n58347), .X(n23847) );
  nand_x1_sg U41615 ( .A(n57314), .B(n58346), .X(n23853) );
  nand_x1_sg U41616 ( .A(n57314), .B(n58345), .X(n23859) );
  nand_x1_sg U41617 ( .A(n57314), .B(n58344), .X(n23865) );
  nand_x1_sg U41618 ( .A(n57314), .B(n58343), .X(n23871) );
  nand_x1_sg U41619 ( .A(n57314), .B(n58342), .X(n23877) );
  nand_x1_sg U41620 ( .A(n57314), .B(n58341), .X(n23883) );
  nand_x1_sg U41621 ( .A(n58374), .B(n58340), .X(n23889) );
  nand_x1_sg U41622 ( .A(n57314), .B(n58339), .X(n23895) );
  nand_x1_sg U41623 ( .A(n57314), .B(n58338), .X(n23901) );
  nand_x1_sg U41624 ( .A(n57314), .B(n58337), .X(n23907) );
  nand_x1_sg U41625 ( .A(n57314), .B(n58336), .X(n23913) );
  nand_x1_sg U41626 ( .A(n57314), .B(n58335), .X(n23919) );
  nand_x1_sg U41627 ( .A(n57314), .B(n58334), .X(n23925) );
  nand_x1_sg U41628 ( .A(n57314), .B(n58333), .X(n23939) );
  inv_x1_sg U41629 ( .A(n58332), .X(n24821) );
  nand_x1_sg U41630 ( .A(n58331), .B(n58330), .X(n58332) );
  inv_x1_sg U41631 ( .A(n58327), .X(n24852) );
  nand_x1_sg U41632 ( .A(n58326), .B(n58325), .X(n58327) );
  inv_x1_sg U41633 ( .A(n58322), .X(n24882) );
  nand_x1_sg U41634 ( .A(n58321), .B(n58320), .X(n58322) );
  nor_x1_sg U41635 ( .A(n58317), .B(n58316), .X(n24912) );
  nor_x1_sg U41636 ( .A(n58312), .B(n58311), .X(n24942) );
  inv_x1_sg U41637 ( .A(n58307), .X(n24972) );
  nand_x1_sg U41638 ( .A(n58306), .B(n58305), .X(n58307) );
  inv_x1_sg U41639 ( .A(n58302), .X(n25002) );
  nand_x1_sg U41640 ( .A(n58301), .B(n58300), .X(n58302) );
  inv_x1_sg U41641 ( .A(n58297), .X(n25032) );
  nand_x1_sg U41642 ( .A(n58296), .B(n58295), .X(n58297) );
  nor_x1_sg U41643 ( .A(n58292), .B(n58291), .X(n25062) );
  nor_x1_sg U41644 ( .A(n58287), .B(n58286), .X(n25092) );
  inv_x1_sg U41645 ( .A(n58282), .X(n25122) );
  nand_x1_sg U41646 ( .A(n58281), .B(n58280), .X(n58282) );
  inv_x1_sg U41647 ( .A(n58277), .X(n25152) );
  nand_x1_sg U41648 ( .A(n58276), .B(n58275), .X(n58277) );
  nor_x1_sg U41649 ( .A(n58272), .B(n58271), .X(n25182) );
  nor_x1_sg U41650 ( .A(n58267), .B(n58266), .X(n25212) );
  inv_x1_sg U41651 ( .A(n58262), .X(n25242) );
  nand_x1_sg U41652 ( .A(n58261), .B(n58260), .X(n58262) );
  inv_x1_sg U41653 ( .A(n58257), .X(n25272) );
  nand_x1_sg U41654 ( .A(n58256), .B(n58255), .X(n58257) );
  inv_x1_sg U41655 ( .A(n58252), .X(n25302) );
  nand_x1_sg U41656 ( .A(n58251), .B(n58250), .X(n58252) );
  nor_x1_sg U41657 ( .A(n58247), .B(n58246), .X(n25332) );
  nor_x1_sg U41658 ( .A(n58242), .B(n58241), .X(n25362) );
  inv_x1_sg U41659 ( .A(n58237), .X(n25393) );
  nand_x1_sg U41660 ( .A(n58236), .B(n58235), .X(n58237) );
  inv_x1_sg U41661 ( .A(n58232), .X(n25424) );
  nand_x1_sg U41662 ( .A(n58231), .B(n58230), .X(n58232) );
  inv_x1_sg U41663 ( .A(n58227), .X(n25454) );
  nand_x1_sg U41664 ( .A(n58226), .B(n58225), .X(n58227) );
  inv_x1_sg U41665 ( .A(n58222), .X(n25484) );
  nand_x1_sg U41666 ( .A(n58221), .B(n58220), .X(n58222) );
  nor_x1_sg U41667 ( .A(n58217), .B(n58216), .X(n25514) );
  nor_x1_sg U41668 ( .A(n58212), .B(n58211), .X(n25544) );
  inv_x1_sg U41669 ( .A(n58207), .X(n25574) );
  nand_x1_sg U41670 ( .A(n58206), .B(n58205), .X(n58207) );
  inv_x1_sg U41671 ( .A(n58202), .X(n25604) );
  nand_x1_sg U41672 ( .A(n58201), .B(n58200), .X(n58202) );
  inv_x1_sg U41673 ( .A(n58197), .X(n25634) );
  nand_x1_sg U41674 ( .A(n58196), .B(n58195), .X(n58197) );
  nor_x1_sg U41675 ( .A(n58192), .B(n58191), .X(n25664) );
  nor_x1_sg U41676 ( .A(n58187), .B(n58186), .X(n25694) );
  inv_x1_sg U41677 ( .A(n58182), .X(n25724) );
  nand_x1_sg U41678 ( .A(n58181), .B(n58180), .X(n58182) );
  inv_x1_sg U41679 ( .A(n58177), .X(n25754) );
  nand_x1_sg U41680 ( .A(n58176), .B(n58175), .X(n58177) );
  nor_x1_sg U41681 ( .A(n58172), .B(n58171), .X(n25784) );
  nor_x1_sg U41682 ( .A(n58167), .B(n58166), .X(n25814) );
  inv_x1_sg U41683 ( .A(n58162), .X(n25844) );
  nand_x1_sg U41684 ( .A(n58161), .B(n58160), .X(n58162) );
  inv_x1_sg U41685 ( .A(n58157), .X(n25874) );
  nand_x1_sg U41686 ( .A(n58156), .B(n58155), .X(n58157) );
  inv_x1_sg U41687 ( .A(n58152), .X(n25904) );
  nand_x1_sg U41688 ( .A(n58151), .B(n58150), .X(n58152) );
  nor_x1_sg U41689 ( .A(n58147), .B(n58146), .X(n25934) );
  nor_x1_sg U41690 ( .A(n58142), .B(n58141), .X(n25964) );
  inv_x1_sg U41691 ( .A(n58137), .X(n25995) );
  nand_x1_sg U41692 ( .A(n58136), .B(n58135), .X(n58137) );
  nand_x1_sg U41693 ( .A(n57455), .B(n24383), .X(n24382) );
  nand_x1_sg U41694 ( .A(n57454), .B(n24388), .X(n24387) );
  nand_x1_sg U41695 ( .A(n57455), .B(n24393), .X(n24392) );
  nand_x1_sg U41696 ( .A(n57455), .B(n24398), .X(n24397) );
  nand_x1_sg U41697 ( .A(n57454), .B(n24403), .X(n24402) );
  nand_x1_sg U41698 ( .A(n57454), .B(n24408), .X(n24407) );
  nand_x1_sg U41699 ( .A(n57454), .B(n24413), .X(n24412) );
  nand_x1_sg U41700 ( .A(n57454), .B(n24418), .X(n24417) );
  nand_x1_sg U41701 ( .A(n57454), .B(n24423), .X(n24422) );
  nand_x1_sg U41702 ( .A(n57454), .B(n24428), .X(n24427) );
  nand_x1_sg U41703 ( .A(n57454), .B(n24433), .X(n24432) );
  nand_x1_sg U41704 ( .A(n57454), .B(n24438), .X(n24437) );
  nand_x1_sg U41705 ( .A(n57455), .B(n24443), .X(n24442) );
  nand_x1_sg U41706 ( .A(n57455), .B(n24448), .X(n24447) );
  nand_x1_sg U41707 ( .A(n57455), .B(n24453), .X(n24452) );
  nand_x1_sg U41708 ( .A(n57455), .B(n24458), .X(n24457) );
  nand_x1_sg U41709 ( .A(n57455), .B(n24463), .X(n24462) );
  nand_x1_sg U41710 ( .A(n57455), .B(n24468), .X(n24467) );
  nand_x1_sg U41711 ( .A(n57455), .B(n24473), .X(n24472) );
  nand_x1_sg U41712 ( .A(n57455), .B(n24489), .X(n24488) );
  nand_x1_sg U41713 ( .A(n57454), .B(n24495), .X(n24494) );
  nand_x1_sg U41714 ( .A(n57455), .B(n24500), .X(n24499) );
  nand_x1_sg U41715 ( .A(n57454), .B(n24505), .X(n24504) );
  nand_x1_sg U41716 ( .A(n57455), .B(n24510), .X(n24509) );
  nand_x1_sg U41717 ( .A(n57454), .B(n24515), .X(n24514) );
  nand_x1_sg U41718 ( .A(n57455), .B(n24520), .X(n24519) );
  nand_x1_sg U41719 ( .A(n57454), .B(n24525), .X(n24524) );
  nand_x1_sg U41720 ( .A(n57455), .B(n24530), .X(n24529) );
  nand_x1_sg U41721 ( .A(n57454), .B(n24535), .X(n24534) );
  nand_x1_sg U41722 ( .A(n57455), .B(n24540), .X(n24539) );
  nand_x1_sg U41723 ( .A(n57454), .B(n24545), .X(n24544) );
  nand_x1_sg U41724 ( .A(n57455), .B(n24550), .X(n24549) );
  nand_x1_sg U41725 ( .A(n57455), .B(n24555), .X(n24554) );
  nand_x1_sg U41726 ( .A(n57454), .B(n24560), .X(n24559) );
  nand_x1_sg U41727 ( .A(n57454), .B(n24565), .X(n24564) );
  nand_x1_sg U41728 ( .A(n57455), .B(n24570), .X(n24569) );
  nand_x1_sg U41729 ( .A(n57454), .B(n24575), .X(n24574) );
  nand_x1_sg U41730 ( .A(n57455), .B(n24580), .X(n24579) );
  nand_x1_sg U41731 ( .A(n57454), .B(n24585), .X(n24584) );
  nand_x1_sg U41732 ( .A(n57455), .B(n24601), .X(n24600) );
  inv_x1_sg U41733 ( .A(n58126), .X(n24606) );
  inv_x1_sg U41734 ( .A(n58120), .X(n24611) );
  inv_x1_sg U41735 ( .A(n58117), .X(n24615) );
  inv_x1_sg U41736 ( .A(n58114), .X(n24619) );
  inv_x1_sg U41737 ( .A(n58110), .X(n24623) );
  inv_x1_sg U41738 ( .A(n58106), .X(n24627) );
  inv_x1_sg U41739 ( .A(n58103), .X(n24631) );
  inv_x1_sg U41740 ( .A(n58100), .X(n24635) );
  inv_x1_sg U41741 ( .A(n58097), .X(n24639) );
  inv_x1_sg U41742 ( .A(n58093), .X(n24643) );
  inv_x1_sg U41743 ( .A(n58089), .X(n24647) );
  inv_x1_sg U41744 ( .A(n58086), .X(n24651) );
  inv_x1_sg U41745 ( .A(n58083), .X(n24655) );
  inv_x1_sg U41746 ( .A(n58079), .X(n24659) );
  inv_x1_sg U41747 ( .A(n58075), .X(n24663) );
  inv_x1_sg U41748 ( .A(n58072), .X(n24667) );
  inv_x1_sg U41749 ( .A(n58069), .X(n24671) );
  inv_x1_sg U41750 ( .A(n58066), .X(n24675) );
  inv_x1_sg U41751 ( .A(n58062), .X(n24679) );
  inv_x1_sg U41752 ( .A(n58058), .X(n24696) );
  inv_x1_sg U41753 ( .A(n58055), .X(n24701) );
  inv_x1_sg U41754 ( .A(n58050), .X(n24705) );
  inv_x1_sg U41755 ( .A(n58047), .X(n24709) );
  inv_x1_sg U41756 ( .A(n58044), .X(n24713) );
  inv_x1_sg U41757 ( .A(n58040), .X(n24717) );
  inv_x1_sg U41758 ( .A(n58036), .X(n24721) );
  inv_x1_sg U41759 ( .A(n58033), .X(n24725) );
  inv_x1_sg U41760 ( .A(n58030), .X(n24729) );
  inv_x1_sg U41761 ( .A(n58027), .X(n24733) );
  inv_x1_sg U41762 ( .A(n58023), .X(n24737) );
  inv_x1_sg U41763 ( .A(n58019), .X(n24741) );
  inv_x1_sg U41764 ( .A(n58016), .X(n24745) );
  inv_x1_sg U41765 ( .A(n58013), .X(n24749) );
  inv_x1_sg U41766 ( .A(n58009), .X(n24753) );
  inv_x1_sg U41767 ( .A(n58005), .X(n24757) );
  inv_x1_sg U41768 ( .A(n58002), .X(n24761) );
  inv_x1_sg U41769 ( .A(n57999), .X(n24765) );
  inv_x1_sg U41770 ( .A(n57996), .X(n24769) );
  inv_x1_sg U41771 ( .A(n57992), .X(n24773) );
  inv_x1_sg U41772 ( .A(n57988), .X(n24789) );
  nor_x1_sg U41773 ( .A(n46879), .B(n46877), .X(n32039) );
  nor_x1_sg U41774 ( .A(n46861), .B(n46859), .X(n31984) );
  nand_x4_sg U41775 ( .A(n31994), .B(n31995), .X(n31974) );
  nor_x1_sg U41776 ( .A(n46875), .B(n46873), .X(n31975) );
  nand_x1_sg U41777 ( .A(n31926), .B(n57918), .X(n31925) );
  nand_x1_sg U41778 ( .A(n31927), .B(n31928), .X(n31926) );
  inv_x1_sg U41779 ( .A(n31995), .X(n68487) );
  inv_x1_sg U41780 ( .A(n31967), .X(n68266) );
  nor_x1_sg U41781 ( .A(n46865), .B(n46863), .X(n32481) );
  nand_x1_sg U41782 ( .A(n57304), .B(n68389), .X(n32388) );
  nor_x1_sg U41783 ( .A(n46869), .B(n46867), .X(n32383) );
  nor_x1_sg U41784 ( .A(n46883), .B(n46881), .X(n32373) );
  nand_x1_sg U41785 ( .A(n32394), .B(n57918), .X(n32393) );
  nand_x1_sg U41786 ( .A(n32395), .B(n32396), .X(n32394) );
  inv_x1_sg U41787 ( .A(n32437), .X(n68398) );
  inv_x1_sg U41788 ( .A(n32374), .X(n68264) );
  inv_x1_sg U41789 ( .A(n40224), .X(n68336) );
  inv_x1_sg U41790 ( .A(n40219), .X(n68335) );
  inv_x1_sg U41791 ( .A(\filter_0/reg_xor_w_mask [30]), .X(n51042) );
  inv_x1_sg U41792 ( .A(n40214), .X(n68334) );
  inv_x1_sg U41793 ( .A(\filter_0/reg_xor_w_mask [29]), .X(n53638) );
  inv_x1_sg U41794 ( .A(n40209), .X(n68333) );
  inv_x1_sg U41795 ( .A(\filter_0/reg_xor_w_mask [28]), .X(n53636) );
  inv_x1_sg U41796 ( .A(n40204), .X(n68332) );
  inv_x1_sg U41797 ( .A(n40199), .X(n68331) );
  inv_x1_sg U41798 ( .A(\filter_0/reg_xor_w_mask [26]), .X(n47582) );
  inv_x1_sg U41799 ( .A(n40194), .X(n68330) );
  inv_x1_sg U41800 ( .A(\filter_0/reg_xor_w_mask [25]), .X(n51040) );
  inv_x1_sg U41801 ( .A(n40189), .X(n68329) );
  inv_x1_sg U41802 ( .A(\filter_0/reg_xor_w_mask [24]), .X(n53634) );
  inv_x1_sg U41803 ( .A(n40184), .X(n68328) );
  inv_x1_sg U41804 ( .A(\filter_0/reg_xor_w_mask [23]), .X(n47594) );
  inv_x1_sg U41805 ( .A(n40179), .X(n68327) );
  inv_x1_sg U41806 ( .A(\filter_0/reg_xor_w_mask [22]), .X(n53632) );
  inv_x1_sg U41807 ( .A(n40174), .X(n68326) );
  inv_x1_sg U41808 ( .A(\filter_0/reg_xor_w_mask [21]), .X(n53630) );
  inv_x1_sg U41809 ( .A(n40169), .X(n68325) );
  inv_x1_sg U41810 ( .A(\filter_0/reg_xor_w_mask [20]), .X(n53628) );
  inv_x1_sg U41811 ( .A(n40164), .X(n68324) );
  inv_x1_sg U41812 ( .A(\filter_0/reg_xor_w_mask [19]), .X(n47502) );
  inv_x1_sg U41813 ( .A(n40159), .X(n68323) );
  inv_x1_sg U41814 ( .A(n40154), .X(n68322) );
  inv_x1_sg U41815 ( .A(\filter_0/reg_xor_w_mask [17]), .X(n53626) );
  inv_x1_sg U41816 ( .A(n40149), .X(n68321) );
  inv_x1_sg U41817 ( .A(\filter_0/reg_xor_w_mask [16]), .X(n53646) );
  inv_x1_sg U41818 ( .A(n40144), .X(n68320) );
  inv_x1_sg U41819 ( .A(n40139), .X(n68319) );
  inv_x1_sg U41820 ( .A(\filter_0/reg_xor_w_mask [14]), .X(n51038) );
  inv_x1_sg U41821 ( .A(n40134), .X(n68318) );
  inv_x1_sg U41822 ( .A(\filter_0/reg_xor_w_mask [13]), .X(n53624) );
  inv_x1_sg U41823 ( .A(n40129), .X(n68317) );
  inv_x1_sg U41824 ( .A(\filter_0/reg_xor_w_mask [12]), .X(n53622) );
  inv_x1_sg U41825 ( .A(n40124), .X(n68316) );
  inv_x1_sg U41826 ( .A(n40119), .X(n68315) );
  inv_x1_sg U41827 ( .A(\filter_0/reg_xor_w_mask [10]), .X(n47580) );
  inv_x1_sg U41828 ( .A(n40114), .X(n68314) );
  inv_x1_sg U41829 ( .A(\filter_0/reg_xor_w_mask [9]), .X(n51036) );
  inv_x1_sg U41830 ( .A(n40109), .X(n68313) );
  inv_x1_sg U41831 ( .A(\filter_0/reg_xor_w_mask [8]), .X(n53620) );
  inv_x1_sg U41832 ( .A(n40104), .X(n68312) );
  inv_x1_sg U41833 ( .A(\filter_0/reg_xor_w_mask [7]), .X(n47592) );
  inv_x1_sg U41834 ( .A(n40099), .X(n68311) );
  inv_x1_sg U41835 ( .A(\filter_0/reg_xor_w_mask [6]), .X(n53618) );
  inv_x1_sg U41836 ( .A(n40094), .X(n68310) );
  inv_x1_sg U41837 ( .A(\filter_0/reg_xor_w_mask [5]), .X(n53616) );
  inv_x1_sg U41838 ( .A(n40089), .X(n68309) );
  inv_x1_sg U41839 ( .A(\filter_0/reg_xor_w_mask [4]), .X(n53614) );
  inv_x1_sg U41840 ( .A(n40084), .X(n68308) );
  inv_x1_sg U41841 ( .A(\filter_0/reg_xor_w_mask [3]), .X(n47500) );
  inv_x1_sg U41842 ( .A(n40079), .X(n68307) );
  inv_x1_sg U41843 ( .A(n40074), .X(n68306) );
  inv_x1_sg U41844 ( .A(\filter_0/reg_xor_w_mask [1]), .X(n53612) );
  inv_x1_sg U41845 ( .A(n40069), .X(n68305) );
  inv_x1_sg U41846 ( .A(\filter_0/reg_xor_w_mask [0]), .X(n53644) );
  inv_x1_sg U41847 ( .A(n40064), .X(n68304) );
  inv_x1_sg U41848 ( .A(n40059), .X(n68303) );
  inv_x1_sg U41849 ( .A(\filter_0/reg_xor_i_mask [30]), .X(n51034) );
  inv_x1_sg U41850 ( .A(n40054), .X(n68302) );
  inv_x1_sg U41851 ( .A(\filter_0/reg_xor_i_mask [29]), .X(n53610) );
  inv_x1_sg U41852 ( .A(n40049), .X(n68301) );
  inv_x1_sg U41853 ( .A(\filter_0/reg_xor_i_mask [28]), .X(n53608) );
  inv_x1_sg U41854 ( .A(n40044), .X(n68300) );
  inv_x1_sg U41855 ( .A(n40039), .X(n68299) );
  inv_x1_sg U41856 ( .A(\filter_0/reg_xor_i_mask [26]), .X(n47578) );
  inv_x1_sg U41857 ( .A(n40034), .X(n68298) );
  inv_x1_sg U41858 ( .A(\filter_0/reg_xor_i_mask [25]), .X(n51032) );
  inv_x1_sg U41859 ( .A(n40029), .X(n68297) );
  inv_x1_sg U41860 ( .A(\filter_0/reg_xor_i_mask [24]), .X(n53606) );
  inv_x1_sg U41861 ( .A(n40024), .X(n68296) );
  inv_x1_sg U41862 ( .A(\filter_0/reg_xor_i_mask [23]), .X(n47590) );
  inv_x1_sg U41863 ( .A(n40019), .X(n68295) );
  inv_x1_sg U41864 ( .A(\filter_0/reg_xor_i_mask [22]), .X(n53604) );
  inv_x1_sg U41865 ( .A(n40014), .X(n68294) );
  inv_x1_sg U41866 ( .A(\filter_0/reg_xor_i_mask [21]), .X(n53602) );
  inv_x1_sg U41867 ( .A(n40009), .X(n68293) );
  inv_x1_sg U41868 ( .A(\filter_0/reg_xor_i_mask [20]), .X(n53600) );
  inv_x1_sg U41869 ( .A(n40004), .X(n68292) );
  inv_x1_sg U41870 ( .A(\filter_0/reg_xor_i_mask [19]), .X(n47498) );
  inv_x1_sg U41871 ( .A(n39999), .X(n68291) );
  inv_x1_sg U41872 ( .A(n39994), .X(n68290) );
  inv_x1_sg U41873 ( .A(\filter_0/reg_xor_i_mask [17]), .X(n53598) );
  inv_x1_sg U41874 ( .A(n39989), .X(n68289) );
  inv_x1_sg U41875 ( .A(\filter_0/reg_xor_i_mask [16]), .X(n53642) );
  inv_x1_sg U41876 ( .A(n39984), .X(n68288) );
  inv_x1_sg U41877 ( .A(n39979), .X(n68287) );
  inv_x1_sg U41878 ( .A(\filter_0/reg_xor_i_mask [14]), .X(n51030) );
  inv_x1_sg U41879 ( .A(n39974), .X(n68286) );
  inv_x1_sg U41880 ( .A(\filter_0/reg_xor_i_mask [13]), .X(n53596) );
  inv_x1_sg U41881 ( .A(n39969), .X(n68285) );
  inv_x1_sg U41882 ( .A(\filter_0/reg_xor_i_mask [12]), .X(n53594) );
  inv_x1_sg U41883 ( .A(n39964), .X(n68284) );
  inv_x1_sg U41884 ( .A(n39959), .X(n68283) );
  inv_x1_sg U41885 ( .A(\filter_0/reg_xor_i_mask [10]), .X(n47576) );
  inv_x1_sg U41886 ( .A(n39954), .X(n68282) );
  inv_x1_sg U41887 ( .A(\filter_0/reg_xor_i_mask [9]), .X(n51028) );
  inv_x1_sg U41888 ( .A(n39949), .X(n68281) );
  inv_x1_sg U41889 ( .A(\filter_0/reg_xor_i_mask [8]), .X(n53592) );
  inv_x1_sg U41890 ( .A(n39944), .X(n68280) );
  inv_x1_sg U41891 ( .A(\filter_0/reg_xor_i_mask [7]), .X(n47588) );
  inv_x1_sg U41892 ( .A(n39939), .X(n68279) );
  inv_x1_sg U41893 ( .A(\filter_0/reg_xor_i_mask [6]), .X(n53590) );
  inv_x1_sg U41894 ( .A(n39934), .X(n68278) );
  inv_x1_sg U41895 ( .A(\filter_0/reg_xor_i_mask [5]), .X(n53588) );
  inv_x1_sg U41896 ( .A(n39929), .X(n68277) );
  inv_x1_sg U41897 ( .A(\filter_0/reg_xor_i_mask [4]), .X(n53586) );
  inv_x1_sg U41898 ( .A(n39924), .X(n68276) );
  inv_x1_sg U41899 ( .A(\filter_0/reg_xor_i_mask [3]), .X(n47496) );
  inv_x1_sg U41900 ( .A(n39919), .X(n68275) );
  inv_x1_sg U41901 ( .A(n39914), .X(n68274) );
  inv_x1_sg U41902 ( .A(\filter_0/reg_xor_i_mask [1]), .X(n53584) );
  inv_x1_sg U41903 ( .A(n39909), .X(n68273) );
  inv_x1_sg U41904 ( .A(\filter_0/reg_xor_i_mask [0]), .X(n53640) );
  inv_x1_sg U41905 ( .A(\filter_0/reg_o_mask [30]), .X(n51048) );
  inv_x1_sg U41906 ( .A(\filter_0/reg_o_mask [29]), .X(n51026) );
  inv_x1_sg U41907 ( .A(\filter_0/reg_o_mask [28]), .X(n51024) );
  inv_x1_sg U41908 ( .A(\filter_0/reg_o_mask [26]), .X(n47596) );
  inv_x1_sg U41909 ( .A(\filter_0/reg_o_mask [25]), .X(n51022) );
  inv_x1_sg U41910 ( .A(\filter_0/reg_o_mask [24]), .X(n51020) );
  inv_x1_sg U41911 ( .A(\filter_0/reg_o_mask [23]), .X(n51050) );
  inv_x1_sg U41912 ( .A(\filter_0/reg_o_mask [22]), .X(n51018) );
  inv_x1_sg U41913 ( .A(\filter_0/reg_o_mask [21]), .X(n51044) );
  inv_x1_sg U41914 ( .A(\filter_0/reg_o_mask [20]), .X(n51016) );
  inv_x1_sg U41915 ( .A(\filter_0/reg_o_mask [19]), .X(n47598) );
  inv_x1_sg U41916 ( .A(\filter_0/reg_o_mask [17]), .X(n47584) );
  inv_x1_sg U41917 ( .A(\filter_0/reg_o_mask [16]), .X(n51014) );
  inv_x1_sg U41918 ( .A(\filter_0/reg_o_mask [14]), .X(n51012) );
  inv_x1_sg U41919 ( .A(\filter_0/reg_o_mask [13]), .X(n51010) );
  inv_x1_sg U41920 ( .A(\filter_0/reg_o_mask [12]), .X(n51008) );
  inv_x1_sg U41921 ( .A(\filter_0/reg_o_mask [10]), .X(n47574) );
  inv_x1_sg U41922 ( .A(\filter_0/reg_o_mask [9]), .X(n51006) );
  inv_x1_sg U41923 ( .A(\filter_0/reg_o_mask [8]), .X(n51004) );
  inv_x1_sg U41924 ( .A(\filter_0/reg_o_mask [7]), .X(n51002) );
  inv_x1_sg U41925 ( .A(\filter_0/reg_o_mask [6]), .X(n51000) );
  inv_x1_sg U41926 ( .A(\filter_0/reg_o_mask [5]), .X(n51046) );
  inv_x1_sg U41927 ( .A(\filter_0/reg_o_mask [4]), .X(n47586) );
  inv_x1_sg U41928 ( .A(\filter_0/n17329 ), .X(n53582) );
  inv_x1_sg U41929 ( .A(\filter_0/n17330 ), .X(n50998) );
  inv_x1_sg U41930 ( .A(\filter_0/n17331 ), .X(n50996) );
  inv_x1_sg U41931 ( .A(\filter_0/n17332 ), .X(n50994) );
  inv_x1_sg U41932 ( .A(\filter_0/n17333 ), .X(n53580) );
  inv_x1_sg U41933 ( .A(\filter_0/n17334 ), .X(n53578) );
  inv_x1_sg U41934 ( .A(\filter_0/n17335 ), .X(n50992) );
  inv_x1_sg U41935 ( .A(\filter_0/n17336 ), .X(n50990) );
  inv_x1_sg U41936 ( .A(\filter_0/n17337 ), .X(n50988) );
  inv_x1_sg U41937 ( .A(\filter_0/n17338 ), .X(n53576) );
  inv_x1_sg U41938 ( .A(\filter_0/n17339 ), .X(n50986) );
  inv_x1_sg U41939 ( .A(\filter_0/n17340 ), .X(n50984) );
  inv_x1_sg U41940 ( .A(\filter_0/n17341 ), .X(n50982) );
  inv_x1_sg U41941 ( .A(\filter_0/n17342 ), .X(n53574) );
  inv_x1_sg U41942 ( .A(\filter_0/n17343 ), .X(n53572) );
  inv_x1_sg U41943 ( .A(\filter_0/n17344 ), .X(n50980) );
  inv_x1_sg U41944 ( .A(\filter_0/n17345 ), .X(n50978) );
  inv_x1_sg U41945 ( .A(\filter_0/n17346 ), .X(n50976) );
  inv_x1_sg U41946 ( .A(\filter_0/n17347 ), .X(n53570) );
  inv_x1_sg U41947 ( .A(\filter_0/n17348 ), .X(n53568) );
  inv_x1_sg U41948 ( .A(\filter_0/n17349 ), .X(n53566) );
  inv_x1_sg U41949 ( .A(\filter_0/n17350 ), .X(n53564) );
  inv_x1_sg U41950 ( .A(\filter_0/n17351 ), .X(n50974) );
  inv_x1_sg U41951 ( .A(\filter_0/n17352 ), .X(n53562) );
  inv_x1_sg U41952 ( .A(\filter_0/n17353 ), .X(n53560) );
  inv_x1_sg U41953 ( .A(\filter_0/n17354 ), .X(n50972) );
  inv_x1_sg U41954 ( .A(\filter_0/n17355 ), .X(n53558) );
  inv_x1_sg U41955 ( .A(\filter_0/n17356 ), .X(n50970) );
  inv_x1_sg U41956 ( .A(\filter_0/n17357 ), .X(n53556) );
  inv_x1_sg U41957 ( .A(\filter_0/n17358 ), .X(n50968) );
  inv_x1_sg U41958 ( .A(\filter_0/n17359 ), .X(n53554) );
  inv_x1_sg U41959 ( .A(\filter_0/n17360 ), .X(n50966) );
  inv_x1_sg U41960 ( .A(\filter_0/n17361 ), .X(n53552) );
  inv_x1_sg U41961 ( .A(\filter_0/n17362 ), .X(n50964) );
  inv_x1_sg U41962 ( .A(\filter_0/n17363 ), .X(n53550) );
  inv_x1_sg U41963 ( .A(\filter_0/n17364 ), .X(n53548) );
  inv_x1_sg U41964 ( .A(\filter_0/n17365 ), .X(n50962) );
  inv_x1_sg U41965 ( .A(\filter_0/n17366 ), .X(n50960) );
  inv_x1_sg U41966 ( .A(\filter_0/n17367 ), .X(n53546) );
  inv_x1_sg U41967 ( .A(\filter_0/n17368 ), .X(n53544) );
  inv_x1_sg U41968 ( .A(\filter_0/n17369 ), .X(n50958) );
  inv_x1_sg U41969 ( .A(\filter_0/n17370 ), .X(n50956) );
  inv_x1_sg U41970 ( .A(\filter_0/n17371 ), .X(n53542) );
  inv_x1_sg U41971 ( .A(\filter_0/n17372 ), .X(n53540) );
  inv_x1_sg U41972 ( .A(\filter_0/n17373 ), .X(n50954) );
  inv_x1_sg U41973 ( .A(\filter_0/n17374 ), .X(n53538) );
  inv_x1_sg U41974 ( .A(\filter_0/n17375 ), .X(n50952) );
  inv_x1_sg U41975 ( .A(\filter_0/n17376 ), .X(n53536) );
  inv_x1_sg U41976 ( .A(\filter_0/n17377 ), .X(n50950) );
  inv_x1_sg U41977 ( .A(\filter_0/n17378 ), .X(n53534) );
  inv_x1_sg U41978 ( .A(\filter_0/n17379 ), .X(n50948) );
  inv_x1_sg U41979 ( .A(\filter_0/n17380 ), .X(n53532) );
  inv_x1_sg U41980 ( .A(\filter_0/n17381 ), .X(n50946) );
  inv_x1_sg U41981 ( .A(\filter_0/n17382 ), .X(n53530) );
  inv_x1_sg U41982 ( .A(\filter_0/n17383 ), .X(n53528) );
  inv_x1_sg U41983 ( .A(\filter_0/n17384 ), .X(n50944) );
  inv_x1_sg U41984 ( .A(\filter_0/n17385 ), .X(n53526) );
  inv_x1_sg U41985 ( .A(\filter_0/n17386 ), .X(n53524) );
  inv_x1_sg U41986 ( .A(\filter_0/n17387 ), .X(n53522) );
  inv_x1_sg U41987 ( .A(\filter_0/n17388 ), .X(n53520) );
  inv_x1_sg U41988 ( .A(\filter_0/n17389 ), .X(n50942) );
  inv_x1_sg U41989 ( .A(\filter_0/n17390 ), .X(n50940) );
  inv_x1_sg U41990 ( .A(\filter_0/n17391 ), .X(n50938) );
  inv_x1_sg U41991 ( .A(\filter_0/n17392 ), .X(n50936) );
  inv_x1_sg U41992 ( .A(\filter_0/n17393 ), .X(n50934) );
  inv_x1_sg U41993 ( .A(\filter_0/n17394 ), .X(n53518) );
  inv_x1_sg U41994 ( .A(\filter_0/n17395 ), .X(n50932) );
  inv_x1_sg U41995 ( .A(\filter_0/n17396 ), .X(n50930) );
  inv_x1_sg U41996 ( .A(\filter_0/n17397 ), .X(n50928) );
  inv_x1_sg U41997 ( .A(\filter_0/n17398 ), .X(n53516) );
  inv_x1_sg U41998 ( .A(\filter_0/n17399 ), .X(n50926) );
  inv_x1_sg U41999 ( .A(\filter_0/n17400 ), .X(n50924) );
  inv_x1_sg U42000 ( .A(\filter_0/n17401 ), .X(n50922) );
  inv_x1_sg U42001 ( .A(\filter_0/n17402 ), .X(n53514) );
  inv_x1_sg U42002 ( .A(\filter_0/n17403 ), .X(n53512) );
  inv_x1_sg U42003 ( .A(\filter_0/n17404 ), .X(n50920) );
  inv_x1_sg U42004 ( .A(\filter_0/n17405 ), .X(n50918) );
  inv_x1_sg U42005 ( .A(\filter_0/n17406 ), .X(n53510) );
  inv_x1_sg U42006 ( .A(\filter_0/n17407 ), .X(n53508) );
  inv_x1_sg U42007 ( .A(\filter_0/n17408 ), .X(n53506) );
  inv_x1_sg U42008 ( .A(\filter_0/n17409 ), .X(n50916) );
  inv_x1_sg U42009 ( .A(\filter_0/n17410 ), .X(n53504) );
  inv_x1_sg U42010 ( .A(\filter_0/n17411 ), .X(n53502) );
  inv_x1_sg U42011 ( .A(\filter_0/n17412 ), .X(n50914) );
  inv_x1_sg U42012 ( .A(\filter_0/n17413 ), .X(n50912) );
  inv_x1_sg U42013 ( .A(\filter_0/n17414 ), .X(n53500) );
  inv_x1_sg U42014 ( .A(\filter_0/n17415 ), .X(n50910) );
  inv_x1_sg U42015 ( .A(\filter_0/n17416 ), .X(n53498) );
  inv_x1_sg U42016 ( .A(\filter_0/n17417 ), .X(n50908) );
  inv_x1_sg U42017 ( .A(\filter_0/n17418 ), .X(n53496) );
  inv_x1_sg U42018 ( .A(\filter_0/n17419 ), .X(n50906) );
  inv_x1_sg U42019 ( .A(\filter_0/n17420 ), .X(n53494) );
  inv_x1_sg U42020 ( .A(\filter_0/n17421 ), .X(n50904) );
  inv_x1_sg U42021 ( .A(\filter_0/n17422 ), .X(n53492) );
  inv_x1_sg U42022 ( .A(\filter_0/n17423 ), .X(n53490) );
  inv_x1_sg U42023 ( .A(\filter_0/n17424 ), .X(n50902) );
  inv_x1_sg U42024 ( .A(\filter_0/n17425 ), .X(n53488) );
  inv_x1_sg U42025 ( .A(\filter_0/n17426 ), .X(n53486) );
  inv_x1_sg U42026 ( .A(\filter_0/n17427 ), .X(n53484) );
  inv_x1_sg U42027 ( .A(\filter_0/n17428 ), .X(n53482) );
  inv_x1_sg U42028 ( .A(\filter_0/n17429 ), .X(n53480) );
  inv_x1_sg U42029 ( .A(\filter_0/n17430 ), .X(n53478) );
  inv_x1_sg U42030 ( .A(\filter_0/n17431 ), .X(n53476) );
  inv_x1_sg U42031 ( .A(\filter_0/n17432 ), .X(n53474) );
  inv_x1_sg U42032 ( .A(\filter_0/n17433 ), .X(n53472) );
  inv_x1_sg U42033 ( .A(\filter_0/n17434 ), .X(n50900) );
  inv_x1_sg U42034 ( .A(\filter_0/n17435 ), .X(n53470) );
  inv_x1_sg U42035 ( .A(\filter_0/n17436 ), .X(n53468) );
  inv_x1_sg U42036 ( .A(\filter_0/n17437 ), .X(n53466) );
  inv_x1_sg U42037 ( .A(\filter_0/n17438 ), .X(n50898) );
  inv_x1_sg U42038 ( .A(\filter_0/n17439 ), .X(n53464) );
  inv_x1_sg U42039 ( .A(\filter_0/n17440 ), .X(n53462) );
  inv_x1_sg U42040 ( .A(\filter_0/n17441 ), .X(n53460) );
  inv_x1_sg U42041 ( .A(\filter_0/n17442 ), .X(n50896) );
  inv_x1_sg U42042 ( .A(\filter_0/n17443 ), .X(n53458) );
  inv_x1_sg U42043 ( .A(\filter_0/n17444 ), .X(n53456) );
  inv_x1_sg U42044 ( .A(\filter_0/n17445 ), .X(n53454) );
  inv_x1_sg U42045 ( .A(\filter_0/n17446 ), .X(n50894) );
  inv_x1_sg U42046 ( .A(\filter_0/n17447 ), .X(n53452) );
  inv_x1_sg U42047 ( .A(\filter_0/n17448 ), .X(n53450) );
  inv_x1_sg U42048 ( .A(\filter_0/n17449 ), .X(n50892) );
  inv_x1_sg U42049 ( .A(\filter_0/n17450 ), .X(n50890) );
  inv_x1_sg U42050 ( .A(\filter_0/n17451 ), .X(n50888) );
  inv_x1_sg U42051 ( .A(\filter_0/n17452 ), .X(n50886) );
  inv_x1_sg U42052 ( .A(\filter_0/n17453 ), .X(n50884) );
  inv_x1_sg U42053 ( .A(\filter_0/n17454 ), .X(n53448) );
  inv_x1_sg U42054 ( .A(\filter_0/n17455 ), .X(n50882) );
  inv_x1_sg U42055 ( .A(\filter_0/n17456 ), .X(n50880) );
  inv_x1_sg U42056 ( .A(\filter_0/n17457 ), .X(n50878) );
  inv_x1_sg U42057 ( .A(\filter_0/n17458 ), .X(n53446) );
  inv_x1_sg U42058 ( .A(\filter_0/n17459 ), .X(n50876) );
  inv_x1_sg U42059 ( .A(\filter_0/n17460 ), .X(n50874) );
  inv_x1_sg U42060 ( .A(\filter_0/n17461 ), .X(n50872) );
  inv_x1_sg U42061 ( .A(\filter_0/n17462 ), .X(n53444) );
  inv_x1_sg U42062 ( .A(\filter_0/n17463 ), .X(n53442) );
  inv_x1_sg U42063 ( .A(\filter_0/n17464 ), .X(n50870) );
  inv_x1_sg U42064 ( .A(\filter_0/n17465 ), .X(n50868) );
  inv_x1_sg U42065 ( .A(\filter_0/n17466 ), .X(n53440) );
  inv_x1_sg U42066 ( .A(\filter_0/n17467 ), .X(n53438) );
  inv_x1_sg U42067 ( .A(\filter_0/n17468 ), .X(n53436) );
  inv_x1_sg U42068 ( .A(\filter_0/n17609 ), .X(n53434) );
  inv_x1_sg U42069 ( .A(\filter_0/n17610 ), .X(n53432) );
  inv_x1_sg U42070 ( .A(\filter_0/n17611 ), .X(n50866) );
  inv_x1_sg U42071 ( .A(\filter_0/n17612 ), .X(n50864) );
  inv_x1_sg U42072 ( .A(\filter_0/n17613 ), .X(n50862) );
  inv_x1_sg U42073 ( .A(\filter_0/n17614 ), .X(n50860) );
  inv_x1_sg U42074 ( .A(\filter_0/n17615 ), .X(n53430) );
  inv_x1_sg U42075 ( .A(\filter_0/n17616 ), .X(n50858) );
  inv_x1_sg U42076 ( .A(\filter_0/n17617 ), .X(n50856) );
  inv_x1_sg U42077 ( .A(\filter_0/n17618 ), .X(n50854) );
  inv_x1_sg U42078 ( .A(\filter_0/n17619 ), .X(n50852) );
  inv_x1_sg U42079 ( .A(\filter_0/n17620 ), .X(n50850) );
  inv_x1_sg U42080 ( .A(\filter_0/n17621 ), .X(n50848) );
  inv_x1_sg U42081 ( .A(\filter_0/n17622 ), .X(n50846) );
  inv_x1_sg U42082 ( .A(\filter_0/n17623 ), .X(n50844) );
  inv_x1_sg U42083 ( .A(\filter_0/n17624 ), .X(n53428) );
  inv_x1_sg U42084 ( .A(\filter_0/n17625 ), .X(n50842) );
  inv_x1_sg U42085 ( .A(\filter_0/n17626 ), .X(n50840) );
  inv_x1_sg U42086 ( .A(\filter_0/n17627 ), .X(n50838) );
  inv_x1_sg U42087 ( .A(\filter_0/n17628 ), .X(n50836) );
  inv_x1_sg U42088 ( .A(\filter_0/n17589 ), .X(n50834) );
  inv_x1_sg U42089 ( .A(\filter_0/n17590 ), .X(n50832) );
  inv_x1_sg U42090 ( .A(\filter_0/n17591 ), .X(n53426) );
  inv_x1_sg U42091 ( .A(\filter_0/n17592 ), .X(n53424) );
  inv_x1_sg U42092 ( .A(\filter_0/n17593 ), .X(n53422) );
  inv_x1_sg U42093 ( .A(\filter_0/n17594 ), .X(n53420) );
  inv_x1_sg U42094 ( .A(\filter_0/n17595 ), .X(n50830) );
  inv_x1_sg U42095 ( .A(\filter_0/n17596 ), .X(n53418) );
  inv_x1_sg U42096 ( .A(\filter_0/n17597 ), .X(n53416) );
  inv_x1_sg U42097 ( .A(\filter_0/n17598 ), .X(n53414) );
  inv_x1_sg U42098 ( .A(\filter_0/n17599 ), .X(n53412) );
  inv_x1_sg U42099 ( .A(\filter_0/n17600 ), .X(n53410) );
  inv_x1_sg U42100 ( .A(\filter_0/n17601 ), .X(n53408) );
  inv_x1_sg U42101 ( .A(\filter_0/n17602 ), .X(n53406) );
  inv_x1_sg U42102 ( .A(\filter_0/n17603 ), .X(n53404) );
  inv_x1_sg U42103 ( .A(\filter_0/n17604 ), .X(n50828) );
  inv_x1_sg U42104 ( .A(\filter_0/n17605 ), .X(n53402) );
  inv_x1_sg U42105 ( .A(\filter_0/n17606 ), .X(n53400) );
  inv_x1_sg U42106 ( .A(\filter_0/n17607 ), .X(n53398) );
  inv_x1_sg U42107 ( .A(\filter_0/n17608 ), .X(n53396) );
  inv_x1_sg U42108 ( .A(\filter_0/n17569 ), .X(n50826) );
  inv_x1_sg U42109 ( .A(\filter_0/n17570 ), .X(n50824) );
  inv_x1_sg U42110 ( .A(\filter_0/n17571 ), .X(n53394) );
  inv_x1_sg U42111 ( .A(\filter_0/n17572 ), .X(n53392) );
  inv_x1_sg U42112 ( .A(\filter_0/n17573 ), .X(n50822) );
  inv_x1_sg U42113 ( .A(\filter_0/n17574 ), .X(n53390) );
  inv_x1_sg U42114 ( .A(\filter_0/n17575 ), .X(n50820) );
  inv_x1_sg U42115 ( .A(\filter_0/n17576 ), .X(n53388) );
  inv_x1_sg U42116 ( .A(\filter_0/n17577 ), .X(n50818) );
  inv_x1_sg U42117 ( .A(\filter_0/n17578 ), .X(n53386) );
  inv_x1_sg U42118 ( .A(\filter_0/n17579 ), .X(n50816) );
  inv_x1_sg U42119 ( .A(\filter_0/n17580 ), .X(n53384) );
  inv_x1_sg U42120 ( .A(\filter_0/n17581 ), .X(n50814) );
  inv_x1_sg U42121 ( .A(\filter_0/n17582 ), .X(n53382) );
  inv_x1_sg U42122 ( .A(\filter_0/n17583 ), .X(n53380) );
  inv_x1_sg U42123 ( .A(\filter_0/n17584 ), .X(n50812) );
  inv_x1_sg U42124 ( .A(\filter_0/n17585 ), .X(n53378) );
  inv_x1_sg U42125 ( .A(\filter_0/n17586 ), .X(n53376) );
  inv_x1_sg U42126 ( .A(\filter_0/n17587 ), .X(n53374) );
  inv_x1_sg U42127 ( .A(\filter_0/n17588 ), .X(n53372) );
  inv_x1_sg U42128 ( .A(\filter_0/n17549 ), .X(n50810) );
  inv_x1_sg U42129 ( .A(\filter_0/n17550 ), .X(n50808) );
  inv_x1_sg U42130 ( .A(\filter_0/n17551 ), .X(n53370) );
  inv_x1_sg U42131 ( .A(\filter_0/n17552 ), .X(n53368) );
  inv_x1_sg U42132 ( .A(\filter_0/n17553 ), .X(n50806) );
  inv_x1_sg U42133 ( .A(\filter_0/n17554 ), .X(n53366) );
  inv_x1_sg U42134 ( .A(\filter_0/n17555 ), .X(n50804) );
  inv_x1_sg U42135 ( .A(\filter_0/n17556 ), .X(n53364) );
  inv_x1_sg U42136 ( .A(\filter_0/n17557 ), .X(n50802) );
  inv_x1_sg U42137 ( .A(\filter_0/n17558 ), .X(n53362) );
  inv_x1_sg U42138 ( .A(\filter_0/n17559 ), .X(n50800) );
  inv_x1_sg U42139 ( .A(\filter_0/n17560 ), .X(n53360) );
  inv_x1_sg U42140 ( .A(\filter_0/n17561 ), .X(n50798) );
  inv_x1_sg U42141 ( .A(\filter_0/n17562 ), .X(n53358) );
  inv_x1_sg U42142 ( .A(\filter_0/n17563 ), .X(n53356) );
  inv_x1_sg U42143 ( .A(\filter_0/n17564 ), .X(n50796) );
  inv_x1_sg U42144 ( .A(\filter_0/n17565 ), .X(n53354) );
  inv_x1_sg U42145 ( .A(\filter_0/n17566 ), .X(n53352) );
  inv_x1_sg U42146 ( .A(\filter_0/n17567 ), .X(n53350) );
  inv_x1_sg U42147 ( .A(\filter_0/n17568 ), .X(n53348) );
  inv_x1_sg U42148 ( .A(\filter_0/n17529 ), .X(n50794) );
  inv_x1_sg U42149 ( .A(\filter_0/n17530 ), .X(n53346) );
  inv_x1_sg U42150 ( .A(\filter_0/n17531 ), .X(n53344) );
  inv_x1_sg U42151 ( .A(\filter_0/n17532 ), .X(n50792) );
  inv_x1_sg U42152 ( .A(\filter_0/n17533 ), .X(n50790) );
  inv_x1_sg U42153 ( .A(\filter_0/n17534 ), .X(n53342) );
  inv_x1_sg U42154 ( .A(\filter_0/n17535 ), .X(n50788) );
  inv_x1_sg U42155 ( .A(\filter_0/n17536 ), .X(n53340) );
  inv_x1_sg U42156 ( .A(\filter_0/n17537 ), .X(n50786) );
  inv_x1_sg U42157 ( .A(\filter_0/n17538 ), .X(n53338) );
  inv_x1_sg U42158 ( .A(\filter_0/n17539 ), .X(n50784) );
  inv_x1_sg U42159 ( .A(\filter_0/n17540 ), .X(n53336) );
  inv_x1_sg U42160 ( .A(\filter_0/n17541 ), .X(n50782) );
  inv_x1_sg U42161 ( .A(\filter_0/n17542 ), .X(n53334) );
  inv_x1_sg U42162 ( .A(\filter_0/n17543 ), .X(n53332) );
  inv_x1_sg U42163 ( .A(\filter_0/n17544 ), .X(n50780) );
  inv_x1_sg U42164 ( .A(\filter_0/n17545 ), .X(n53330) );
  inv_x1_sg U42165 ( .A(\filter_0/n17546 ), .X(n53328) );
  inv_x1_sg U42166 ( .A(\filter_0/n17547 ), .X(n53326) );
  inv_x1_sg U42167 ( .A(\filter_0/n17548 ), .X(n53324) );
  inv_x1_sg U42168 ( .A(\filter_0/n17509 ), .X(n53322) );
  inv_x1_sg U42169 ( .A(\filter_0/n17510 ), .X(n53320) );
  inv_x1_sg U42170 ( .A(\filter_0/n17511 ), .X(n50778) );
  inv_x1_sg U42171 ( .A(\filter_0/n17512 ), .X(n53318) );
  inv_x1_sg U42172 ( .A(\filter_0/n17513 ), .X(n50776) );
  inv_x1_sg U42173 ( .A(\filter_0/n17514 ), .X(n53316) );
  inv_x1_sg U42174 ( .A(\filter_0/n17515 ), .X(n53314) );
  inv_x1_sg U42175 ( .A(\filter_0/n17516 ), .X(n50774) );
  inv_x1_sg U42176 ( .A(\filter_0/n17517 ), .X(n53312) );
  inv_x1_sg U42177 ( .A(\filter_0/n17518 ), .X(n50772) );
  inv_x1_sg U42178 ( .A(\filter_0/n17519 ), .X(n53310) );
  inv_x1_sg U42179 ( .A(\filter_0/n17520 ), .X(n50770) );
  inv_x1_sg U42180 ( .A(\filter_0/n17521 ), .X(n53308) );
  inv_x1_sg U42181 ( .A(\filter_0/n17522 ), .X(n50768) );
  inv_x1_sg U42182 ( .A(\filter_0/n17523 ), .X(n53306) );
  inv_x1_sg U42183 ( .A(\filter_0/n17524 ), .X(n53304) );
  inv_x1_sg U42184 ( .A(\filter_0/n17525 ), .X(n50766) );
  inv_x1_sg U42185 ( .A(\filter_0/n17526 ), .X(n50764) );
  inv_x1_sg U42186 ( .A(\filter_0/n17527 ), .X(n53302) );
  inv_x1_sg U42187 ( .A(\filter_0/n17528 ), .X(n53300) );
  inv_x1_sg U42188 ( .A(\filter_0/n17489 ), .X(n53298) );
  inv_x1_sg U42189 ( .A(\filter_0/n17490 ), .X(n50762) );
  inv_x1_sg U42190 ( .A(\filter_0/n17491 ), .X(n53296) );
  inv_x1_sg U42191 ( .A(\filter_0/n17492 ), .X(n53294) );
  inv_x1_sg U42192 ( .A(\filter_0/n17493 ), .X(n53292) );
  inv_x1_sg U42193 ( .A(\filter_0/n17494 ), .X(n50760) );
  inv_x1_sg U42194 ( .A(\filter_0/n17495 ), .X(n53290) );
  inv_x1_sg U42195 ( .A(\filter_0/n17496 ), .X(n50758) );
  inv_x1_sg U42196 ( .A(\filter_0/n17497 ), .X(n53288) );
  inv_x1_sg U42197 ( .A(\filter_0/n17498 ), .X(n50756) );
  inv_x1_sg U42198 ( .A(\filter_0/n17499 ), .X(n53286) );
  inv_x1_sg U42199 ( .A(\filter_0/n17500 ), .X(n50754) );
  inv_x1_sg U42200 ( .A(\filter_0/n17501 ), .X(n53284) );
  inv_x1_sg U42201 ( .A(\filter_0/n17502 ), .X(n50752) );
  inv_x1_sg U42202 ( .A(\filter_0/n17503 ), .X(n53282) );
  inv_x1_sg U42203 ( .A(\filter_0/n17504 ), .X(n53280) );
  inv_x1_sg U42204 ( .A(\filter_0/n17505 ), .X(n50750) );
  inv_x1_sg U42205 ( .A(\filter_0/n17506 ), .X(n50748) );
  inv_x1_sg U42206 ( .A(\filter_0/n17507 ), .X(n53278) );
  inv_x1_sg U42207 ( .A(\filter_0/n17508 ), .X(n53276) );
  inv_x1_sg U42208 ( .A(\filter_0/n17469 ), .X(n50746) );
  inv_x1_sg U42209 ( .A(\filter_0/n17470 ), .X(n50744) );
  inv_x1_sg U42210 ( .A(\filter_0/n17471 ), .X(n53274) );
  inv_x1_sg U42211 ( .A(\filter_0/n17472 ), .X(n50742) );
  inv_x1_sg U42212 ( .A(\filter_0/n17473 ), .X(n53272) );
  inv_x1_sg U42213 ( .A(\filter_0/n17474 ), .X(n53270) );
  inv_x1_sg U42214 ( .A(\filter_0/n17475 ), .X(n50740) );
  inv_x1_sg U42215 ( .A(\filter_0/n17476 ), .X(n53268) );
  inv_x1_sg U42216 ( .A(\filter_0/n17477 ), .X(n50738) );
  inv_x1_sg U42217 ( .A(\filter_0/n17478 ), .X(n53266) );
  inv_x1_sg U42218 ( .A(\filter_0/n17479 ), .X(n50736) );
  inv_x1_sg U42219 ( .A(\filter_0/n17480 ), .X(n53264) );
  inv_x1_sg U42220 ( .A(\filter_0/n17481 ), .X(n50734) );
  inv_x1_sg U42221 ( .A(\filter_0/n17482 ), .X(n53262) );
  inv_x1_sg U42222 ( .A(\filter_0/n17483 ), .X(n53260) );
  inv_x1_sg U42223 ( .A(\filter_0/n17484 ), .X(n50732) );
  inv_x1_sg U42224 ( .A(\filter_0/n17485 ), .X(n53258) );
  inv_x1_sg U42225 ( .A(\filter_0/n17486 ), .X(n53256) );
  inv_x1_sg U42226 ( .A(\filter_0/n17487 ), .X(n53254) );
  inv_x1_sg U42227 ( .A(\filter_0/n17488 ), .X(n53252) );
  inv_x1_sg U42228 ( .A(\filter_0/n17309 ), .X(n50730) );
  inv_x1_sg U42229 ( .A(\filter_0/n17310 ), .X(n50728) );
  inv_x1_sg U42230 ( .A(\filter_0/n17311 ), .X(n50726) );
  inv_x1_sg U42231 ( .A(\filter_0/n17312 ), .X(n50724) );
  inv_x1_sg U42232 ( .A(\filter_0/n17313 ), .X(n50722) );
  inv_x1_sg U42233 ( .A(\filter_0/n17314 ), .X(n53250) );
  inv_x1_sg U42234 ( .A(\filter_0/n17315 ), .X(n50720) );
  inv_x1_sg U42235 ( .A(\filter_0/n17316 ), .X(n50718) );
  inv_x1_sg U42236 ( .A(\filter_0/n17317 ), .X(n50716) );
  inv_x1_sg U42237 ( .A(\filter_0/n17318 ), .X(n50714) );
  inv_x1_sg U42238 ( .A(\filter_0/n17319 ), .X(n50712) );
  inv_x1_sg U42239 ( .A(\filter_0/n17320 ), .X(n50710) );
  inv_x1_sg U42240 ( .A(\filter_0/n17321 ), .X(n50708) );
  inv_x1_sg U42241 ( .A(\filter_0/n17322 ), .X(n50706) );
  inv_x1_sg U42242 ( .A(\filter_0/n17323 ), .X(n53248) );
  inv_x1_sg U42243 ( .A(\filter_0/n17324 ), .X(n50704) );
  inv_x1_sg U42244 ( .A(\filter_0/n17325 ), .X(n50702) );
  inv_x1_sg U42245 ( .A(\filter_0/n17326 ), .X(n50700) );
  inv_x1_sg U42246 ( .A(\filter_0/n17327 ), .X(n53246) );
  inv_x1_sg U42247 ( .A(\filter_0/n17328 ), .X(n53244) );
  inv_x1_sg U42248 ( .A(\filter_0/n17649 ), .X(n53242) );
  inv_x1_sg U42249 ( .A(\filter_0/n17650 ), .X(n50698) );
  inv_x1_sg U42250 ( .A(\filter_0/n17651 ), .X(n50696) );
  inv_x1_sg U42251 ( .A(\filter_0/n17652 ), .X(n50694) );
  inv_x1_sg U42252 ( .A(\filter_0/n17653 ), .X(n53240) );
  inv_x1_sg U42253 ( .A(\filter_0/n17654 ), .X(n53238) );
  inv_x1_sg U42254 ( .A(\filter_0/n17655 ), .X(n50692) );
  inv_x1_sg U42255 ( .A(\filter_0/n17656 ), .X(n50690) );
  inv_x1_sg U42256 ( .A(\filter_0/n17657 ), .X(n50688) );
  inv_x1_sg U42257 ( .A(\filter_0/n17658 ), .X(n53236) );
  inv_x1_sg U42258 ( .A(\filter_0/n17659 ), .X(n50686) );
  inv_x1_sg U42259 ( .A(\filter_0/n17660 ), .X(n50684) );
  inv_x1_sg U42260 ( .A(\filter_0/n17661 ), .X(n50682) );
  inv_x1_sg U42261 ( .A(\filter_0/n17662 ), .X(n53234) );
  inv_x1_sg U42262 ( .A(\filter_0/n17663 ), .X(n53232) );
  inv_x1_sg U42263 ( .A(\filter_0/n17664 ), .X(n50680) );
  inv_x1_sg U42264 ( .A(\filter_0/n17665 ), .X(n50678) );
  inv_x1_sg U42265 ( .A(\filter_0/n17666 ), .X(n50676) );
  inv_x1_sg U42266 ( .A(\filter_0/n17667 ), .X(n53230) );
  inv_x1_sg U42267 ( .A(\filter_0/n17668 ), .X(n53228) );
  inv_x1_sg U42268 ( .A(\filter_0/n17669 ), .X(n53226) );
  inv_x1_sg U42269 ( .A(\filter_0/n17670 ), .X(n53224) );
  inv_x1_sg U42270 ( .A(\filter_0/n17671 ), .X(n50674) );
  inv_x1_sg U42271 ( .A(\filter_0/n17672 ), .X(n53222) );
  inv_x1_sg U42272 ( .A(\filter_0/n17673 ), .X(n53220) );
  inv_x1_sg U42273 ( .A(\filter_0/n17674 ), .X(n50672) );
  inv_x1_sg U42274 ( .A(\filter_0/n17675 ), .X(n53218) );
  inv_x1_sg U42275 ( .A(\filter_0/n17676 ), .X(n50670) );
  inv_x1_sg U42276 ( .A(\filter_0/n17677 ), .X(n53216) );
  inv_x1_sg U42277 ( .A(\filter_0/n17678 ), .X(n50668) );
  inv_x1_sg U42278 ( .A(\filter_0/n17679 ), .X(n53214) );
  inv_x1_sg U42279 ( .A(\filter_0/n17680 ), .X(n50666) );
  inv_x1_sg U42280 ( .A(\filter_0/n17681 ), .X(n53212) );
  inv_x1_sg U42281 ( .A(\filter_0/n17682 ), .X(n50664) );
  inv_x1_sg U42282 ( .A(\filter_0/n17683 ), .X(n53210) );
  inv_x1_sg U42283 ( .A(\filter_0/n17684 ), .X(n53208) );
  inv_x1_sg U42284 ( .A(\filter_0/n17685 ), .X(n50662) );
  inv_x1_sg U42285 ( .A(\filter_0/n17686 ), .X(n50660) );
  inv_x1_sg U42286 ( .A(\filter_0/n17687 ), .X(n53206) );
  inv_x1_sg U42287 ( .A(\filter_0/n17688 ), .X(n53204) );
  inv_x1_sg U42288 ( .A(\filter_0/n17689 ), .X(n50658) );
  inv_x1_sg U42289 ( .A(\filter_0/n17690 ), .X(n50656) );
  inv_x1_sg U42290 ( .A(\filter_0/n17691 ), .X(n53202) );
  inv_x1_sg U42291 ( .A(\filter_0/n17692 ), .X(n53200) );
  inv_x1_sg U42292 ( .A(\filter_0/n17693 ), .X(n50654) );
  inv_x1_sg U42293 ( .A(\filter_0/n17694 ), .X(n53198) );
  inv_x1_sg U42294 ( .A(\filter_0/n17695 ), .X(n50652) );
  inv_x1_sg U42295 ( .A(\filter_0/n17696 ), .X(n53196) );
  inv_x1_sg U42296 ( .A(\filter_0/n17697 ), .X(n50650) );
  inv_x1_sg U42297 ( .A(\filter_0/n17698 ), .X(n53194) );
  inv_x1_sg U42298 ( .A(\filter_0/n17699 ), .X(n50648) );
  inv_x1_sg U42299 ( .A(\filter_0/n17700 ), .X(n53192) );
  inv_x1_sg U42300 ( .A(\filter_0/n17701 ), .X(n50646) );
  inv_x1_sg U42301 ( .A(\filter_0/n17702 ), .X(n53190) );
  inv_x1_sg U42302 ( .A(\filter_0/n17703 ), .X(n53188) );
  inv_x1_sg U42303 ( .A(\filter_0/n17704 ), .X(n50644) );
  inv_x1_sg U42304 ( .A(\filter_0/n17705 ), .X(n53186) );
  inv_x1_sg U42305 ( .A(\filter_0/n17706 ), .X(n53184) );
  inv_x1_sg U42306 ( .A(\filter_0/n17707 ), .X(n53182) );
  inv_x1_sg U42307 ( .A(\filter_0/n17708 ), .X(n53180) );
  inv_x1_sg U42308 ( .A(\filter_0/n17709 ), .X(n50642) );
  inv_x1_sg U42309 ( .A(\filter_0/n17710 ), .X(n50640) );
  inv_x1_sg U42310 ( .A(\filter_0/n17711 ), .X(n50638) );
  inv_x1_sg U42311 ( .A(\filter_0/n17712 ), .X(n50636) );
  inv_x1_sg U42312 ( .A(\filter_0/n17713 ), .X(n50634) );
  inv_x1_sg U42313 ( .A(\filter_0/n17714 ), .X(n53178) );
  inv_x1_sg U42314 ( .A(\filter_0/n17715 ), .X(n50632) );
  inv_x1_sg U42315 ( .A(\filter_0/n17716 ), .X(n50630) );
  inv_x1_sg U42316 ( .A(\filter_0/n17717 ), .X(n50628) );
  inv_x1_sg U42317 ( .A(\filter_0/n17718 ), .X(n53176) );
  inv_x1_sg U42318 ( .A(\filter_0/n17719 ), .X(n50626) );
  inv_x1_sg U42319 ( .A(\filter_0/n17720 ), .X(n50624) );
  inv_x1_sg U42320 ( .A(\filter_0/n17721 ), .X(n50622) );
  inv_x1_sg U42321 ( .A(\filter_0/n17722 ), .X(n53174) );
  inv_x1_sg U42322 ( .A(\filter_0/n17723 ), .X(n53172) );
  inv_x1_sg U42323 ( .A(\filter_0/n17724 ), .X(n50620) );
  inv_x1_sg U42324 ( .A(\filter_0/n17725 ), .X(n50618) );
  inv_x1_sg U42325 ( .A(\filter_0/n17726 ), .X(n53170) );
  inv_x1_sg U42326 ( .A(\filter_0/n17727 ), .X(n53168) );
  inv_x1_sg U42327 ( .A(\filter_0/n17728 ), .X(n53166) );
  inv_x1_sg U42328 ( .A(\filter_0/n17729 ), .X(n50616) );
  inv_x1_sg U42329 ( .A(\filter_0/n17730 ), .X(n53164) );
  inv_x1_sg U42330 ( .A(\filter_0/n17731 ), .X(n53162) );
  inv_x1_sg U42331 ( .A(\filter_0/n17732 ), .X(n50614) );
  inv_x1_sg U42332 ( .A(\filter_0/n17733 ), .X(n50612) );
  inv_x1_sg U42333 ( .A(\filter_0/n17734 ), .X(n53160) );
  inv_x1_sg U42334 ( .A(\filter_0/n17735 ), .X(n50610) );
  inv_x1_sg U42335 ( .A(\filter_0/n17736 ), .X(n53158) );
  inv_x1_sg U42336 ( .A(\filter_0/n17737 ), .X(n50608) );
  inv_x1_sg U42337 ( .A(\filter_0/n17738 ), .X(n53156) );
  inv_x1_sg U42338 ( .A(\filter_0/n17739 ), .X(n50606) );
  inv_x1_sg U42339 ( .A(\filter_0/n17740 ), .X(n53154) );
  inv_x1_sg U42340 ( .A(\filter_0/n17741 ), .X(n50604) );
  inv_x1_sg U42341 ( .A(\filter_0/n17742 ), .X(n53152) );
  inv_x1_sg U42342 ( .A(\filter_0/n17743 ), .X(n53150) );
  inv_x1_sg U42343 ( .A(\filter_0/n17744 ), .X(n50602) );
  inv_x1_sg U42344 ( .A(\filter_0/n17745 ), .X(n53148) );
  inv_x1_sg U42345 ( .A(\filter_0/n17746 ), .X(n53146) );
  inv_x1_sg U42346 ( .A(\filter_0/n17747 ), .X(n53144) );
  inv_x1_sg U42347 ( .A(\filter_0/n17748 ), .X(n53142) );
  inv_x1_sg U42348 ( .A(\filter_0/n17749 ), .X(n53140) );
  inv_x1_sg U42349 ( .A(\filter_0/n17750 ), .X(n53138) );
  inv_x1_sg U42350 ( .A(\filter_0/n17751 ), .X(n53136) );
  inv_x1_sg U42351 ( .A(\filter_0/n17752 ), .X(n53134) );
  inv_x1_sg U42352 ( .A(\filter_0/n17753 ), .X(n53132) );
  inv_x1_sg U42353 ( .A(\filter_0/n17754 ), .X(n50600) );
  inv_x1_sg U42354 ( .A(\filter_0/n17755 ), .X(n53130) );
  inv_x1_sg U42355 ( .A(\filter_0/n17756 ), .X(n53128) );
  inv_x1_sg U42356 ( .A(\filter_0/n17757 ), .X(n53126) );
  inv_x1_sg U42357 ( .A(\filter_0/n17758 ), .X(n50598) );
  inv_x1_sg U42358 ( .A(\filter_0/n17759 ), .X(n53124) );
  inv_x1_sg U42359 ( .A(\filter_0/n17760 ), .X(n53122) );
  inv_x1_sg U42360 ( .A(\filter_0/n17761 ), .X(n53120) );
  inv_x1_sg U42361 ( .A(\filter_0/n17762 ), .X(n50596) );
  inv_x1_sg U42362 ( .A(\filter_0/n17763 ), .X(n53118) );
  inv_x1_sg U42363 ( .A(\filter_0/n17764 ), .X(n53116) );
  inv_x1_sg U42364 ( .A(\filter_0/n17765 ), .X(n53114) );
  inv_x1_sg U42365 ( .A(\filter_0/n17766 ), .X(n50594) );
  inv_x1_sg U42366 ( .A(\filter_0/n17767 ), .X(n53112) );
  inv_x1_sg U42367 ( .A(\filter_0/n17768 ), .X(n53110) );
  inv_x1_sg U42368 ( .A(\filter_0/n17769 ), .X(n50592) );
  inv_x1_sg U42369 ( .A(\filter_0/n17770 ), .X(n50590) );
  inv_x1_sg U42370 ( .A(\filter_0/n17771 ), .X(n50588) );
  inv_x1_sg U42371 ( .A(\filter_0/n17772 ), .X(n50586) );
  inv_x1_sg U42372 ( .A(\filter_0/n17773 ), .X(n50584) );
  inv_x1_sg U42373 ( .A(\filter_0/n17774 ), .X(n53108) );
  inv_x1_sg U42374 ( .A(\filter_0/n17775 ), .X(n50582) );
  inv_x1_sg U42375 ( .A(\filter_0/n17776 ), .X(n50580) );
  inv_x1_sg U42376 ( .A(\filter_0/n17777 ), .X(n50578) );
  inv_x1_sg U42377 ( .A(\filter_0/n17778 ), .X(n53106) );
  inv_x1_sg U42378 ( .A(\filter_0/n17779 ), .X(n50576) );
  inv_x1_sg U42379 ( .A(\filter_0/n17780 ), .X(n50574) );
  inv_x1_sg U42380 ( .A(\filter_0/n17781 ), .X(n50572) );
  inv_x1_sg U42381 ( .A(\filter_0/n17782 ), .X(n53104) );
  inv_x1_sg U42382 ( .A(\filter_0/n17783 ), .X(n53102) );
  inv_x1_sg U42383 ( .A(\filter_0/n17784 ), .X(n50570) );
  inv_x1_sg U42384 ( .A(\filter_0/n17785 ), .X(n50568) );
  inv_x1_sg U42385 ( .A(\filter_0/n17786 ), .X(n53100) );
  inv_x1_sg U42386 ( .A(\filter_0/n17787 ), .X(n53098) );
  inv_x1_sg U42387 ( .A(\filter_0/n17788 ), .X(n53096) );
  inv_x1_sg U42388 ( .A(\filter_0/n17929 ), .X(n50566) );
  inv_x1_sg U42389 ( .A(\filter_0/n17930 ), .X(n53094) );
  inv_x1_sg U42390 ( .A(\filter_0/n17931 ), .X(n50564) );
  inv_x1_sg U42391 ( .A(\filter_0/n17932 ), .X(n50562) );
  inv_x1_sg U42392 ( .A(\filter_0/n17933 ), .X(n50560) );
  inv_x1_sg U42393 ( .A(\filter_0/n17934 ), .X(n50558) );
  inv_x1_sg U42394 ( .A(\filter_0/n17935 ), .X(n53092) );
  inv_x1_sg U42395 ( .A(\filter_0/n17936 ), .X(n50556) );
  inv_x1_sg U42396 ( .A(\filter_0/n17937 ), .X(n50554) );
  inv_x1_sg U42397 ( .A(\filter_0/n17938 ), .X(n50552) );
  inv_x1_sg U42398 ( .A(\filter_0/n17939 ), .X(n50550) );
  inv_x1_sg U42399 ( .A(\filter_0/n17940 ), .X(n50548) );
  inv_x1_sg U42400 ( .A(\filter_0/n17941 ), .X(n50546) );
  inv_x1_sg U42401 ( .A(\filter_0/n17942 ), .X(n50544) );
  inv_x1_sg U42402 ( .A(\filter_0/n17943 ), .X(n50542) );
  inv_x1_sg U42403 ( .A(\filter_0/n17944 ), .X(n53090) );
  inv_x1_sg U42404 ( .A(\filter_0/n17945 ), .X(n50540) );
  inv_x1_sg U42405 ( .A(\filter_0/n17946 ), .X(n50538) );
  inv_x1_sg U42406 ( .A(\filter_0/n17947 ), .X(n53088) );
  inv_x1_sg U42407 ( .A(\filter_0/n17948 ), .X(n50536) );
  inv_x1_sg U42408 ( .A(\filter_0/n17909 ), .X(n53086) );
  inv_x1_sg U42409 ( .A(\filter_0/n17910 ), .X(n50534) );
  inv_x1_sg U42410 ( .A(\filter_0/n17911 ), .X(n53084) );
  inv_x1_sg U42411 ( .A(\filter_0/n17912 ), .X(n53082) );
  inv_x1_sg U42412 ( .A(\filter_0/n17913 ), .X(n53080) );
  inv_x1_sg U42413 ( .A(\filter_0/n17914 ), .X(n53078) );
  inv_x1_sg U42414 ( .A(\filter_0/n17915 ), .X(n50532) );
  inv_x1_sg U42415 ( .A(\filter_0/n17916 ), .X(n53076) );
  inv_x1_sg U42416 ( .A(\filter_0/n17917 ), .X(n53074) );
  inv_x1_sg U42417 ( .A(\filter_0/n17918 ), .X(n53072) );
  inv_x1_sg U42418 ( .A(\filter_0/n17919 ), .X(n53070) );
  inv_x1_sg U42419 ( .A(\filter_0/n17920 ), .X(n53068) );
  inv_x1_sg U42420 ( .A(\filter_0/n17921 ), .X(n53066) );
  inv_x1_sg U42421 ( .A(\filter_0/n17922 ), .X(n53064) );
  inv_x1_sg U42422 ( .A(\filter_0/n17923 ), .X(n53062) );
  inv_x1_sg U42423 ( .A(\filter_0/n17924 ), .X(n50530) );
  inv_x1_sg U42424 ( .A(\filter_0/n17925 ), .X(n53060) );
  inv_x1_sg U42425 ( .A(\filter_0/n17926 ), .X(n53058) );
  inv_x1_sg U42426 ( .A(\filter_0/n17927 ), .X(n50528) );
  inv_x1_sg U42427 ( .A(\filter_0/n17928 ), .X(n53056) );
  inv_x1_sg U42428 ( .A(\filter_0/n17889 ), .X(n50526) );
  inv_x1_sg U42429 ( .A(\filter_0/n17890 ), .X(n50524) );
  inv_x1_sg U42430 ( .A(\filter_0/n17891 ), .X(n53054) );
  inv_x1_sg U42431 ( .A(\filter_0/n17892 ), .X(n53052) );
  inv_x1_sg U42432 ( .A(\filter_0/n17893 ), .X(n50522) );
  inv_x1_sg U42433 ( .A(\filter_0/n17894 ), .X(n53050) );
  inv_x1_sg U42434 ( .A(\filter_0/n17895 ), .X(n50520) );
  inv_x1_sg U42435 ( .A(\filter_0/n17896 ), .X(n53048) );
  inv_x1_sg U42436 ( .A(\filter_0/n17897 ), .X(n50518) );
  inv_x1_sg U42437 ( .A(\filter_0/n17898 ), .X(n53046) );
  inv_x1_sg U42438 ( .A(\filter_0/n17899 ), .X(n50516) );
  inv_x1_sg U42439 ( .A(\filter_0/n17900 ), .X(n53044) );
  inv_x1_sg U42440 ( .A(\filter_0/n17901 ), .X(n50514) );
  inv_x1_sg U42441 ( .A(\filter_0/n17902 ), .X(n53042) );
  inv_x1_sg U42442 ( .A(\filter_0/n17903 ), .X(n53040) );
  inv_x1_sg U42443 ( .A(\filter_0/n17904 ), .X(n50512) );
  inv_x1_sg U42444 ( .A(\filter_0/n17905 ), .X(n53038) );
  inv_x1_sg U42445 ( .A(\filter_0/n17906 ), .X(n53036) );
  inv_x1_sg U42446 ( .A(\filter_0/n17907 ), .X(n53034) );
  inv_x1_sg U42447 ( .A(\filter_0/n17908 ), .X(n53032) );
  inv_x1_sg U42448 ( .A(\filter_0/n17869 ), .X(n50510) );
  inv_x1_sg U42449 ( .A(\filter_0/n17870 ), .X(n50508) );
  inv_x1_sg U42450 ( .A(\filter_0/n17871 ), .X(n53030) );
  inv_x1_sg U42451 ( .A(\filter_0/n17872 ), .X(n53028) );
  inv_x1_sg U42452 ( .A(\filter_0/n17873 ), .X(n50506) );
  inv_x1_sg U42453 ( .A(\filter_0/n17874 ), .X(n53026) );
  inv_x1_sg U42454 ( .A(\filter_0/n17875 ), .X(n50504) );
  inv_x1_sg U42455 ( .A(\filter_0/n17876 ), .X(n53024) );
  inv_x1_sg U42456 ( .A(\filter_0/n17877 ), .X(n50502) );
  inv_x1_sg U42457 ( .A(\filter_0/n17878 ), .X(n53022) );
  inv_x1_sg U42458 ( .A(\filter_0/n17879 ), .X(n50500) );
  inv_x1_sg U42459 ( .A(\filter_0/n17880 ), .X(n53020) );
  inv_x1_sg U42460 ( .A(\filter_0/n17881 ), .X(n50498) );
  inv_x1_sg U42461 ( .A(\filter_0/n17882 ), .X(n53018) );
  inv_x1_sg U42462 ( .A(\filter_0/n17883 ), .X(n53016) );
  inv_x1_sg U42463 ( .A(\filter_0/n17884 ), .X(n50496) );
  inv_x1_sg U42464 ( .A(\filter_0/n17885 ), .X(n53014) );
  inv_x1_sg U42465 ( .A(\filter_0/n17886 ), .X(n53012) );
  inv_x1_sg U42466 ( .A(\filter_0/n17887 ), .X(n53010) );
  inv_x1_sg U42467 ( .A(\filter_0/n17888 ), .X(n53008) );
  inv_x1_sg U42468 ( .A(\filter_0/n17849 ), .X(n50494) );
  inv_x1_sg U42469 ( .A(\filter_0/n17850 ), .X(n53006) );
  inv_x1_sg U42470 ( .A(\filter_0/n17851 ), .X(n53004) );
  inv_x1_sg U42471 ( .A(\filter_0/n17852 ), .X(n50492) );
  inv_x1_sg U42472 ( .A(\filter_0/n17853 ), .X(n50490) );
  inv_x1_sg U42473 ( .A(\filter_0/n17854 ), .X(n53002) );
  inv_x1_sg U42474 ( .A(\filter_0/n17855 ), .X(n50488) );
  inv_x1_sg U42475 ( .A(\filter_0/n17856 ), .X(n53000) );
  inv_x1_sg U42476 ( .A(\filter_0/n17857 ), .X(n50486) );
  inv_x1_sg U42477 ( .A(\filter_0/n17858 ), .X(n52998) );
  inv_x1_sg U42478 ( .A(\filter_0/n17859 ), .X(n50484) );
  inv_x1_sg U42479 ( .A(\filter_0/n17860 ), .X(n52996) );
  inv_x1_sg U42480 ( .A(\filter_0/n17861 ), .X(n50482) );
  inv_x1_sg U42481 ( .A(\filter_0/n17862 ), .X(n52994) );
  inv_x1_sg U42482 ( .A(\filter_0/n17863 ), .X(n52992) );
  inv_x1_sg U42483 ( .A(\filter_0/n17864 ), .X(n50480) );
  inv_x1_sg U42484 ( .A(\filter_0/n17865 ), .X(n52990) );
  inv_x1_sg U42485 ( .A(\filter_0/n17866 ), .X(n52988) );
  inv_x1_sg U42486 ( .A(\filter_0/n17867 ), .X(n52986) );
  inv_x1_sg U42487 ( .A(\filter_0/n17868 ), .X(n52984) );
  inv_x1_sg U42488 ( .A(\filter_0/n17829 ), .X(n52982) );
  inv_x1_sg U42489 ( .A(\filter_0/n17830 ), .X(n52980) );
  inv_x1_sg U42490 ( .A(\filter_0/n17831 ), .X(n50478) );
  inv_x1_sg U42491 ( .A(\filter_0/n17832 ), .X(n52978) );
  inv_x1_sg U42492 ( .A(\filter_0/n17833 ), .X(n50476) );
  inv_x1_sg U42493 ( .A(\filter_0/n17834 ), .X(n52976) );
  inv_x1_sg U42494 ( .A(\filter_0/n17835 ), .X(n52974) );
  inv_x1_sg U42495 ( .A(\filter_0/n17836 ), .X(n50474) );
  inv_x1_sg U42496 ( .A(\filter_0/n17837 ), .X(n52972) );
  inv_x1_sg U42497 ( .A(\filter_0/n17838 ), .X(n50472) );
  inv_x1_sg U42498 ( .A(\filter_0/n17839 ), .X(n52970) );
  inv_x1_sg U42499 ( .A(\filter_0/n17840 ), .X(n50470) );
  inv_x1_sg U42500 ( .A(\filter_0/n17841 ), .X(n52968) );
  inv_x1_sg U42501 ( .A(\filter_0/n17842 ), .X(n50468) );
  inv_x1_sg U42502 ( .A(\filter_0/n17843 ), .X(n52966) );
  inv_x1_sg U42503 ( .A(\filter_0/n17844 ), .X(n52964) );
  inv_x1_sg U42504 ( .A(\filter_0/n17845 ), .X(n50466) );
  inv_x1_sg U42505 ( .A(\filter_0/n17846 ), .X(n50464) );
  inv_x1_sg U42506 ( .A(\filter_0/n17847 ), .X(n52962) );
  inv_x1_sg U42507 ( .A(\filter_0/n17848 ), .X(n52960) );
  inv_x1_sg U42508 ( .A(\filter_0/n17809 ), .X(n52958) );
  inv_x1_sg U42509 ( .A(\filter_0/n17810 ), .X(n50462) );
  inv_x1_sg U42510 ( .A(\filter_0/n17811 ), .X(n52956) );
  inv_x1_sg U42511 ( .A(\filter_0/n17812 ), .X(n52954) );
  inv_x1_sg U42512 ( .A(\filter_0/n17813 ), .X(n52952) );
  inv_x1_sg U42513 ( .A(\filter_0/n17814 ), .X(n50460) );
  inv_x1_sg U42514 ( .A(\filter_0/n17815 ), .X(n52950) );
  inv_x1_sg U42515 ( .A(\filter_0/n17816 ), .X(n50458) );
  inv_x1_sg U42516 ( .A(\filter_0/n17817 ), .X(n52948) );
  inv_x1_sg U42517 ( .A(\filter_0/n17818 ), .X(n50456) );
  inv_x1_sg U42518 ( .A(\filter_0/n17819 ), .X(n52946) );
  inv_x1_sg U42519 ( .A(\filter_0/n17820 ), .X(n50454) );
  inv_x1_sg U42520 ( .A(\filter_0/n17821 ), .X(n52944) );
  inv_x1_sg U42521 ( .A(\filter_0/n17822 ), .X(n50452) );
  inv_x1_sg U42522 ( .A(\filter_0/n17823 ), .X(n52942) );
  inv_x1_sg U42523 ( .A(\filter_0/n17824 ), .X(n52940) );
  inv_x1_sg U42524 ( .A(\filter_0/n17825 ), .X(n50450) );
  inv_x1_sg U42525 ( .A(\filter_0/n17826 ), .X(n50448) );
  inv_x1_sg U42526 ( .A(\filter_0/n17827 ), .X(n52938) );
  inv_x1_sg U42527 ( .A(\filter_0/n17828 ), .X(n52936) );
  inv_x1_sg U42528 ( .A(\filter_0/n17789 ), .X(n50446) );
  inv_x1_sg U42529 ( .A(\filter_0/n17790 ), .X(n50444) );
  inv_x1_sg U42530 ( .A(\filter_0/n17791 ), .X(n52934) );
  inv_x1_sg U42531 ( .A(\filter_0/n17792 ), .X(n50442) );
  inv_x1_sg U42532 ( .A(\filter_0/n17793 ), .X(n52932) );
  inv_x1_sg U42533 ( .A(\filter_0/n17794 ), .X(n52930) );
  inv_x1_sg U42534 ( .A(\filter_0/n17795 ), .X(n50440) );
  inv_x1_sg U42535 ( .A(\filter_0/n17796 ), .X(n52928) );
  inv_x1_sg U42536 ( .A(\filter_0/n17797 ), .X(n50438) );
  inv_x1_sg U42537 ( .A(\filter_0/n17798 ), .X(n52926) );
  inv_x1_sg U42538 ( .A(\filter_0/n17799 ), .X(n50436) );
  inv_x1_sg U42539 ( .A(\filter_0/n17800 ), .X(n52924) );
  inv_x1_sg U42540 ( .A(\filter_0/n17801 ), .X(n50434) );
  inv_x1_sg U42541 ( .A(\filter_0/n17802 ), .X(n52922) );
  inv_x1_sg U42542 ( .A(\filter_0/n17803 ), .X(n52920) );
  inv_x1_sg U42543 ( .A(\filter_0/n17804 ), .X(n50432) );
  inv_x1_sg U42544 ( .A(\filter_0/n17805 ), .X(n52918) );
  inv_x1_sg U42545 ( .A(\filter_0/n17806 ), .X(n52916) );
  inv_x1_sg U42546 ( .A(\filter_0/n17807 ), .X(n52914) );
  inv_x1_sg U42547 ( .A(\filter_0/n17808 ), .X(n52912) );
  inv_x1_sg U42548 ( .A(\filter_0/n17629 ), .X(n50430) );
  inv_x1_sg U42549 ( .A(\filter_0/n17630 ), .X(n50428) );
  inv_x1_sg U42550 ( .A(\filter_0/n17631 ), .X(n50426) );
  inv_x1_sg U42551 ( .A(\filter_0/n17632 ), .X(n50424) );
  inv_x1_sg U42552 ( .A(\filter_0/n17633 ), .X(n50422) );
  inv_x1_sg U42553 ( .A(\filter_0/n17634 ), .X(n52910) );
  inv_x1_sg U42554 ( .A(\filter_0/n17635 ), .X(n50420) );
  inv_x1_sg U42555 ( .A(\filter_0/n17636 ), .X(n50418) );
  inv_x1_sg U42556 ( .A(\filter_0/n17637 ), .X(n50416) );
  inv_x1_sg U42557 ( .A(\filter_0/n17638 ), .X(n50414) );
  inv_x1_sg U42558 ( .A(\filter_0/n17639 ), .X(n50412) );
  inv_x1_sg U42559 ( .A(\filter_0/n17640 ), .X(n50410) );
  inv_x1_sg U42560 ( .A(\filter_0/n17641 ), .X(n50408) );
  inv_x1_sg U42561 ( .A(\filter_0/n17642 ), .X(n50406) );
  inv_x1_sg U42562 ( .A(\filter_0/n17643 ), .X(n52908) );
  inv_x1_sg U42563 ( .A(\filter_0/n17644 ), .X(n50404) );
  inv_x1_sg U42564 ( .A(\filter_0/n17645 ), .X(n50402) );
  inv_x1_sg U42565 ( .A(\filter_0/n17646 ), .X(n50400) );
  inv_x1_sg U42566 ( .A(\filter_0/n17647 ), .X(n52906) );
  inv_x1_sg U42567 ( .A(\filter_0/n17648 ), .X(n52904) );
  nand_x1_sg U42568 ( .A(n39701), .B(n39702), .X(n39700) );
  inv_x1_sg U42569 ( .A(n35841), .X(n68371) );
  inv_x1_sg U42570 ( .A(\mask_0/reg_w_mask [27]), .X(n53710) );
  inv_x1_sg U42571 ( .A(\mask_0/reg_w_mask [26]), .X(n53708) );
  inv_x1_sg U42572 ( .A(\mask_0/reg_w_mask [25]), .X(n53706) );
  inv_x1_sg U42573 ( .A(\mask_0/reg_w_mask [24]), .X(n53704) );
  inv_x1_sg U42574 ( .A(\mask_0/reg_w_mask [23]), .X(n53702) );
  inv_x1_sg U42575 ( .A(\mask_0/reg_w_mask [22]), .X(n53700) );
  inv_x1_sg U42576 ( .A(\mask_0/reg_w_mask [21]), .X(n53698) );
  inv_x1_sg U42577 ( .A(\mask_0/reg_w_mask [20]), .X(n53696) );
  inv_x1_sg U42578 ( .A(\mask_0/reg_w_mask [19]), .X(n53694) );
  inv_x1_sg U42579 ( .A(\mask_0/reg_w_mask [18]), .X(n53692) );
  inv_x1_sg U42580 ( .A(\mask_0/reg_w_mask [16]), .X(n53690) );
  inv_x1_sg U42581 ( .A(\mask_0/reg_w_mask [15]), .X(n53688) );
  inv_x1_sg U42582 ( .A(\mask_0/reg_w_mask [14]), .X(n53686) );
  inv_x1_sg U42583 ( .A(\mask_0/reg_w_mask [13]), .X(n53684) );
  inv_x1_sg U42584 ( .A(\mask_0/reg_w_mask [12]), .X(n53682) );
  inv_x1_sg U42585 ( .A(\mask_0/reg_w_mask [11]), .X(n53680) );
  inv_x1_sg U42586 ( .A(\mask_0/reg_w_mask [10]), .X(n53678) );
  inv_x1_sg U42587 ( .A(\mask_0/reg_w_mask [9]), .X(n53676) );
  inv_x1_sg U42588 ( .A(\mask_0/reg_w_mask [8]), .X(n53674) );
  inv_x1_sg U42589 ( .A(\mask_0/reg_w_mask [7]), .X(n53672) );
  inv_x1_sg U42590 ( .A(\mask_0/reg_w_mask [6]), .X(n53670) );
  inv_x1_sg U42591 ( .A(\mask_0/reg_w_mask [3]), .X(n53668) );
  inv_x1_sg U42592 ( .A(\mask_0/reg_w_mask [2]), .X(n53666) );
  inv_x1_sg U42593 ( .A(\mask_0/reg_w_mask [1]), .X(n53664) );
  inv_x1_sg U42594 ( .A(\mask_0/reg_i_mask [31]), .X(n53662) );
  inv_x1_sg U42595 ( .A(\mask_0/reg_i_mask [30]), .X(n53660) );
  inv_x1_sg U42596 ( .A(\mask_0/reg_i_mask [29]), .X(n53658) );
  inv_x1_sg U42597 ( .A(\mask_0/reg_i_mask [28]), .X(n53656) );
  inv_x1_sg U42598 ( .A(\mask_0/reg_i_mask [17]), .X(n53654) );
  inv_x1_sg U42599 ( .A(\mask_0/reg_i_mask [5]), .X(n53652) );
  inv_x1_sg U42600 ( .A(\mask_0/reg_i_mask [4]), .X(n53650) );
  inv_x1_sg U42601 ( .A(\mask_0/reg_i_mask [0]), .X(n53648) );
  inv_x1_sg U42602 ( .A(reg_www_13[14]), .X(n50398) );
  inv_x1_sg U42603 ( .A(reg_ww_13[14]), .X(n52902) );
  inv_x1_sg U42604 ( .A(reg_www_13[15]), .X(n50396) );
  inv_x1_sg U42605 ( .A(reg_ww_13[15]), .X(n52900) );
  inv_x1_sg U42606 ( .A(reg_www_13[16]), .X(n50394) );
  inv_x1_sg U42607 ( .A(reg_ww_13[16]), .X(n52898) );
  inv_x1_sg U42608 ( .A(reg_www_13[17]), .X(n50392) );
  inv_x1_sg U42609 ( .A(reg_ww_13[17]), .X(n52896) );
  inv_x1_sg U42610 ( .A(reg_www_13[18]), .X(n50390) );
  inv_x1_sg U42611 ( .A(reg_ww_13[18]), .X(n52894) );
  inv_x1_sg U42612 ( .A(reg_www_13[19]), .X(n50388) );
  inv_x1_sg U42613 ( .A(reg_ww_13[19]), .X(n52892) );
  inv_x1_sg U42614 ( .A(reg_www_14[0]), .X(n50386) );
  inv_x1_sg U42615 ( .A(reg_ww_14[0]), .X(n52890) );
  inv_x1_sg U42616 ( .A(reg_www_14[1]), .X(n50384) );
  inv_x1_sg U42617 ( .A(reg_ww_14[1]), .X(n52888) );
  inv_x1_sg U42618 ( .A(reg_www_14[2]), .X(n50382) );
  inv_x1_sg U42619 ( .A(reg_ww_14[2]), .X(n52886) );
  inv_x1_sg U42620 ( .A(reg_www_14[3]), .X(n50380) );
  inv_x1_sg U42621 ( .A(reg_ww_14[3]), .X(n52884) );
  inv_x1_sg U42622 ( .A(reg_www_14[4]), .X(n50378) );
  inv_x1_sg U42623 ( .A(reg_ww_14[4]), .X(n52882) );
  inv_x1_sg U42624 ( .A(reg_www_14[5]), .X(n50376) );
  inv_x1_sg U42625 ( .A(reg_ww_14[5]), .X(n52880) );
  inv_x1_sg U42626 ( .A(reg_www_14[6]), .X(n50374) );
  inv_x1_sg U42627 ( .A(reg_ww_14[6]), .X(n52878) );
  inv_x1_sg U42628 ( .A(reg_www_14[7]), .X(n50372) );
  inv_x1_sg U42629 ( .A(reg_ww_14[7]), .X(n52876) );
  inv_x1_sg U42630 ( .A(reg_www_14[8]), .X(n50370) );
  inv_x1_sg U42631 ( .A(reg_ww_14[8]), .X(n52874) );
  inv_x1_sg U42632 ( .A(reg_www_14[9]), .X(n50368) );
  inv_x1_sg U42633 ( .A(reg_ww_14[9]), .X(n52872) );
  inv_x1_sg U42634 ( .A(reg_www_14[10]), .X(n50366) );
  inv_x1_sg U42635 ( .A(reg_ww_14[10]), .X(n52870) );
  inv_x1_sg U42636 ( .A(reg_www_14[11]), .X(n50364) );
  inv_x1_sg U42637 ( .A(reg_ww_14[11]), .X(n52868) );
  inv_x1_sg U42638 ( .A(reg_www_14[12]), .X(n50362) );
  inv_x1_sg U42639 ( .A(reg_ww_14[12]), .X(n52866) );
  inv_x1_sg U42640 ( .A(reg_www_14[13]), .X(n50360) );
  inv_x1_sg U42641 ( .A(reg_ww_14[13]), .X(n52864) );
  inv_x1_sg U42642 ( .A(reg_www_14[14]), .X(n50358) );
  inv_x1_sg U42643 ( .A(reg_ww_14[14]), .X(n52862) );
  inv_x1_sg U42644 ( .A(reg_www_14[15]), .X(n50356) );
  inv_x1_sg U42645 ( .A(reg_ww_14[15]), .X(n52860) );
  inv_x1_sg U42646 ( .A(reg_www_14[16]), .X(n50354) );
  inv_x1_sg U42647 ( .A(reg_ww_14[16]), .X(n52858) );
  inv_x1_sg U42648 ( .A(reg_www_14[17]), .X(n50352) );
  inv_x1_sg U42649 ( .A(reg_ww_14[17]), .X(n52856) );
  inv_x1_sg U42650 ( .A(reg_www_14[18]), .X(n50350) );
  inv_x1_sg U42651 ( .A(reg_ww_14[18]), .X(n52854) );
  inv_x1_sg U42652 ( .A(reg_www_14[19]), .X(n50348) );
  inv_x1_sg U42653 ( .A(reg_ww_14[19]), .X(n52852) );
  inv_x1_sg U42654 ( .A(reg_www_15[0]), .X(n50346) );
  inv_x1_sg U42655 ( .A(reg_ww_15[0]), .X(n52850) );
  inv_x1_sg U42656 ( .A(reg_www_15[1]), .X(n50344) );
  inv_x1_sg U42657 ( .A(reg_ww_15[1]), .X(n52848) );
  inv_x1_sg U42658 ( .A(reg_www_15[2]), .X(n50342) );
  inv_x1_sg U42659 ( .A(reg_ww_15[2]), .X(n52846) );
  inv_x1_sg U42660 ( .A(reg_www_15[3]), .X(n50340) );
  inv_x1_sg U42661 ( .A(reg_ww_15[3]), .X(n52844) );
  inv_x1_sg U42662 ( .A(reg_www_15[4]), .X(n50338) );
  inv_x1_sg U42663 ( .A(reg_ww_15[4]), .X(n52842) );
  inv_x1_sg U42664 ( .A(reg_www_15[5]), .X(n50336) );
  inv_x1_sg U42665 ( .A(reg_ww_15[5]), .X(n52840) );
  inv_x1_sg U42666 ( .A(reg_www_15[6]), .X(n50334) );
  inv_x1_sg U42667 ( .A(reg_ww_15[6]), .X(n52838) );
  inv_x1_sg U42668 ( .A(reg_www_15[7]), .X(n50332) );
  inv_x1_sg U42669 ( .A(reg_ww_15[7]), .X(n52836) );
  inv_x1_sg U42670 ( .A(reg_www_15[8]), .X(n50330) );
  inv_x1_sg U42671 ( .A(reg_ww_15[8]), .X(n52834) );
  inv_x1_sg U42672 ( .A(reg_www_15[9]), .X(n50328) );
  inv_x1_sg U42673 ( .A(reg_ww_15[9]), .X(n52832) );
  inv_x1_sg U42674 ( .A(reg_www_15[10]), .X(n50326) );
  inv_x1_sg U42675 ( .A(reg_ww_15[10]), .X(n52830) );
  inv_x1_sg U42676 ( .A(reg_www_15[11]), .X(n50324) );
  inv_x1_sg U42677 ( .A(reg_ww_15[11]), .X(n52828) );
  inv_x1_sg U42678 ( .A(reg_www_15[12]), .X(n50322) );
  inv_x1_sg U42679 ( .A(reg_ww_15[12]), .X(n52826) );
  inv_x1_sg U42680 ( .A(reg_www_15[13]), .X(n50320) );
  inv_x1_sg U42681 ( .A(reg_ww_15[13]), .X(n52824) );
  inv_x1_sg U42682 ( .A(reg_www_15[14]), .X(n50318) );
  inv_x1_sg U42683 ( .A(reg_ww_15[14]), .X(n52822) );
  inv_x1_sg U42684 ( .A(reg_www_15[15]), .X(n50316) );
  inv_x1_sg U42685 ( .A(reg_ww_15[15]), .X(n52820) );
  inv_x1_sg U42686 ( .A(reg_www_15[16]), .X(n50314) );
  inv_x1_sg U42687 ( .A(reg_ww_15[16]), .X(n52818) );
  inv_x1_sg U42688 ( .A(reg_www_15[17]), .X(n50312) );
  inv_x1_sg U42689 ( .A(reg_ww_15[17]), .X(n52816) );
  inv_x1_sg U42690 ( .A(reg_www_15[18]), .X(n50310) );
  inv_x1_sg U42691 ( .A(reg_ww_15[18]), .X(n52814) );
  inv_x1_sg U42692 ( .A(reg_www_15[19]), .X(n50308) );
  inv_x1_sg U42693 ( .A(reg_ww_15[19]), .X(n52812) );
  inv_x1_sg U42694 ( .A(reg_www_8[15]), .X(n50306) );
  inv_x1_sg U42695 ( .A(reg_ww_8[15]), .X(n52810) );
  inv_x1_sg U42696 ( .A(reg_www_8[16]), .X(n50304) );
  inv_x1_sg U42697 ( .A(reg_ww_8[16]), .X(n52808) );
  inv_x1_sg U42698 ( .A(reg_www_8[17]), .X(n50302) );
  inv_x1_sg U42699 ( .A(reg_ww_8[17]), .X(n52806) );
  inv_x1_sg U42700 ( .A(reg_www_8[18]), .X(n50300) );
  inv_x1_sg U42701 ( .A(reg_ww_8[18]), .X(n52804) );
  inv_x1_sg U42702 ( .A(reg_www_8[19]), .X(n50298) );
  inv_x1_sg U42703 ( .A(reg_ww_8[19]), .X(n52802) );
  inv_x1_sg U42704 ( .A(reg_www_9[0]), .X(n50296) );
  inv_x1_sg U42705 ( .A(reg_ww_9[0]), .X(n52800) );
  inv_x1_sg U42706 ( .A(reg_www_9[1]), .X(n50294) );
  inv_x1_sg U42707 ( .A(reg_ww_9[1]), .X(n52798) );
  inv_x1_sg U42708 ( .A(reg_www_9[2]), .X(n50292) );
  inv_x1_sg U42709 ( .A(reg_ww_9[2]), .X(n52796) );
  inv_x1_sg U42710 ( .A(reg_www_9[3]), .X(n50290) );
  inv_x1_sg U42711 ( .A(reg_ww_9[3]), .X(n52794) );
  inv_x1_sg U42712 ( .A(reg_www_9[4]), .X(n50288) );
  inv_x1_sg U42713 ( .A(reg_ww_9[4]), .X(n52792) );
  inv_x1_sg U42714 ( .A(reg_www_9[5]), .X(n50286) );
  inv_x1_sg U42715 ( .A(reg_ww_9[5]), .X(n52790) );
  inv_x1_sg U42716 ( .A(reg_www_9[6]), .X(n50284) );
  inv_x1_sg U42717 ( .A(reg_ww_9[6]), .X(n52788) );
  inv_x1_sg U42718 ( .A(reg_www_9[7]), .X(n50282) );
  inv_x1_sg U42719 ( .A(reg_ww_9[7]), .X(n52786) );
  inv_x1_sg U42720 ( .A(reg_www_9[8]), .X(n50280) );
  inv_x1_sg U42721 ( .A(reg_ww_9[8]), .X(n52784) );
  inv_x1_sg U42722 ( .A(reg_www_9[9]), .X(n50278) );
  inv_x1_sg U42723 ( .A(reg_ww_9[9]), .X(n52782) );
  inv_x1_sg U42724 ( .A(reg_www_9[10]), .X(n50276) );
  inv_x1_sg U42725 ( .A(reg_ww_9[10]), .X(n52780) );
  inv_x1_sg U42726 ( .A(reg_www_9[11]), .X(n50274) );
  inv_x1_sg U42727 ( .A(reg_ww_9[11]), .X(n52778) );
  inv_x1_sg U42728 ( .A(reg_www_9[12]), .X(n50272) );
  inv_x1_sg U42729 ( .A(reg_ww_9[12]), .X(n52776) );
  inv_x1_sg U42730 ( .A(reg_www_9[13]), .X(n50270) );
  inv_x1_sg U42731 ( .A(reg_ww_9[13]), .X(n52774) );
  inv_x1_sg U42732 ( .A(reg_www_9[14]), .X(n50268) );
  inv_x1_sg U42733 ( .A(reg_ww_9[14]), .X(n52772) );
  inv_x1_sg U42734 ( .A(reg_www_9[15]), .X(n50266) );
  inv_x1_sg U42735 ( .A(reg_ww_9[15]), .X(n52770) );
  inv_x1_sg U42736 ( .A(reg_www_9[16]), .X(n50264) );
  inv_x1_sg U42737 ( .A(reg_ww_9[16]), .X(n52768) );
  inv_x1_sg U42738 ( .A(reg_www_9[17]), .X(n50262) );
  inv_x1_sg U42739 ( .A(reg_ww_9[17]), .X(n52766) );
  inv_x1_sg U42740 ( .A(reg_www_9[18]), .X(n50260) );
  inv_x1_sg U42741 ( .A(reg_ww_9[18]), .X(n52764) );
  inv_x1_sg U42742 ( .A(reg_www_9[19]), .X(n50258) );
  inv_x1_sg U42743 ( .A(reg_ww_9[19]), .X(n52762) );
  inv_x1_sg U42744 ( .A(reg_www_10[0]), .X(n50256) );
  inv_x1_sg U42745 ( .A(reg_ww_10[0]), .X(n52760) );
  inv_x1_sg U42746 ( .A(reg_www_10[1]), .X(n50254) );
  inv_x1_sg U42747 ( .A(reg_ww_10[1]), .X(n52758) );
  inv_x1_sg U42748 ( .A(reg_www_10[2]), .X(n50252) );
  inv_x1_sg U42749 ( .A(reg_ww_10[2]), .X(n52756) );
  inv_x1_sg U42750 ( .A(reg_www_10[3]), .X(n50250) );
  inv_x1_sg U42751 ( .A(reg_ww_10[3]), .X(n52754) );
  inv_x1_sg U42752 ( .A(reg_www_10[4]), .X(n50248) );
  inv_x1_sg U42753 ( .A(reg_ww_10[4]), .X(n52752) );
  inv_x1_sg U42754 ( .A(reg_www_10[5]), .X(n50246) );
  inv_x1_sg U42755 ( .A(reg_ww_10[5]), .X(n52750) );
  inv_x1_sg U42756 ( .A(reg_www_10[6]), .X(n50244) );
  inv_x1_sg U42757 ( .A(reg_ww_10[6]), .X(n52748) );
  inv_x1_sg U42758 ( .A(reg_www_10[7]), .X(n50242) );
  inv_x1_sg U42759 ( .A(reg_ww_10[7]), .X(n52746) );
  inv_x1_sg U42760 ( .A(reg_www_10[8]), .X(n50240) );
  inv_x1_sg U42761 ( .A(reg_ww_10[8]), .X(n52744) );
  inv_x1_sg U42762 ( .A(reg_www_10[9]), .X(n50238) );
  inv_x1_sg U42763 ( .A(reg_ww_10[9]), .X(n52742) );
  inv_x1_sg U42764 ( .A(reg_www_10[10]), .X(n50236) );
  inv_x1_sg U42765 ( .A(reg_ww_10[10]), .X(n52740) );
  inv_x1_sg U42766 ( .A(reg_www_10[11]), .X(n50234) );
  inv_x1_sg U42767 ( .A(reg_ww_10[11]), .X(n52738) );
  inv_x1_sg U42768 ( .A(reg_www_10[12]), .X(n50232) );
  inv_x1_sg U42769 ( .A(reg_ww_10[12]), .X(n52736) );
  inv_x1_sg U42770 ( .A(reg_www_10[13]), .X(n50230) );
  inv_x1_sg U42771 ( .A(reg_ww_10[13]), .X(n52734) );
  inv_x1_sg U42772 ( .A(reg_www_10[14]), .X(n50228) );
  inv_x1_sg U42773 ( .A(reg_ww_10[14]), .X(n52732) );
  inv_x1_sg U42774 ( .A(reg_www_10[15]), .X(n50226) );
  inv_x1_sg U42775 ( .A(reg_ww_10[15]), .X(n52730) );
  inv_x1_sg U42776 ( .A(reg_www_10[16]), .X(n50224) );
  inv_x1_sg U42777 ( .A(reg_ww_10[16]), .X(n52728) );
  inv_x1_sg U42778 ( .A(reg_www_10[17]), .X(n50222) );
  inv_x1_sg U42779 ( .A(reg_ww_10[17]), .X(n52726) );
  inv_x1_sg U42780 ( .A(reg_www_10[18]), .X(n50220) );
  inv_x1_sg U42781 ( .A(reg_ww_10[18]), .X(n52724) );
  inv_x1_sg U42782 ( .A(reg_www_10[19]), .X(n50218) );
  inv_x1_sg U42783 ( .A(reg_ww_10[19]), .X(n52722) );
  inv_x1_sg U42784 ( .A(reg_www_11[0]), .X(n50216) );
  inv_x1_sg U42785 ( .A(reg_ww_11[0]), .X(n52720) );
  inv_x1_sg U42786 ( .A(reg_www_11[1]), .X(n50214) );
  inv_x1_sg U42787 ( .A(reg_ww_11[1]), .X(n52718) );
  inv_x1_sg U42788 ( .A(reg_www_11[2]), .X(n50212) );
  inv_x1_sg U42789 ( .A(reg_ww_11[2]), .X(n52716) );
  inv_x1_sg U42790 ( .A(reg_www_11[3]), .X(n50210) );
  inv_x1_sg U42791 ( .A(reg_ww_11[3]), .X(n52714) );
  inv_x1_sg U42792 ( .A(reg_www_11[4]), .X(n50208) );
  inv_x1_sg U42793 ( .A(reg_ww_11[4]), .X(n52712) );
  inv_x1_sg U42794 ( .A(reg_www_11[5]), .X(n50206) );
  inv_x1_sg U42795 ( .A(reg_ww_11[5]), .X(n52710) );
  inv_x1_sg U42796 ( .A(reg_www_11[6]), .X(n50204) );
  inv_x1_sg U42797 ( .A(reg_ww_11[6]), .X(n52708) );
  inv_x1_sg U42798 ( .A(reg_www_11[7]), .X(n50202) );
  inv_x1_sg U42799 ( .A(reg_ww_11[7]), .X(n52706) );
  inv_x1_sg U42800 ( .A(reg_www_11[8]), .X(n50200) );
  inv_x1_sg U42801 ( .A(reg_ww_11[8]), .X(n52704) );
  inv_x1_sg U42802 ( .A(reg_www_11[9]), .X(n50198) );
  inv_x1_sg U42803 ( .A(reg_ww_11[9]), .X(n52702) );
  inv_x1_sg U42804 ( .A(reg_www_11[10]), .X(n50196) );
  inv_x1_sg U42805 ( .A(reg_ww_11[10]), .X(n52700) );
  inv_x1_sg U42806 ( .A(reg_www_11[11]), .X(n50194) );
  inv_x1_sg U42807 ( .A(reg_ww_11[11]), .X(n52698) );
  inv_x1_sg U42808 ( .A(reg_www_11[12]), .X(n50192) );
  inv_x1_sg U42809 ( .A(reg_ww_11[12]), .X(n52696) );
  inv_x1_sg U42810 ( .A(reg_www_11[13]), .X(n50190) );
  inv_x1_sg U42811 ( .A(reg_ww_11[13]), .X(n52694) );
  inv_x1_sg U42812 ( .A(reg_www_11[14]), .X(n50188) );
  inv_x1_sg U42813 ( .A(reg_ww_11[14]), .X(n52692) );
  inv_x1_sg U42814 ( .A(reg_www_11[15]), .X(n50186) );
  inv_x1_sg U42815 ( .A(reg_ww_11[15]), .X(n52690) );
  inv_x1_sg U42816 ( .A(reg_www_11[16]), .X(n50184) );
  inv_x1_sg U42817 ( .A(reg_ww_11[16]), .X(n52688) );
  inv_x1_sg U42818 ( .A(reg_www_11[17]), .X(n50182) );
  inv_x1_sg U42819 ( .A(reg_ww_11[17]), .X(n52686) );
  inv_x1_sg U42820 ( .A(reg_www_11[18]), .X(n50180) );
  inv_x1_sg U42821 ( .A(reg_ww_11[18]), .X(n52684) );
  inv_x1_sg U42822 ( .A(reg_www_11[19]), .X(n50178) );
  inv_x1_sg U42823 ( .A(reg_ww_11[19]), .X(n52682) );
  inv_x1_sg U42824 ( .A(reg_www_12[0]), .X(n50176) );
  inv_x1_sg U42825 ( .A(reg_ww_12[0]), .X(n52680) );
  inv_x1_sg U42826 ( .A(reg_www_12[1]), .X(n50174) );
  inv_x1_sg U42827 ( .A(reg_ww_12[1]), .X(n52678) );
  inv_x1_sg U42828 ( .A(reg_www_12[2]), .X(n50172) );
  inv_x1_sg U42829 ( .A(reg_ww_12[2]), .X(n52676) );
  inv_x1_sg U42830 ( .A(reg_www_12[3]), .X(n50170) );
  inv_x1_sg U42831 ( .A(reg_ww_12[3]), .X(n52674) );
  inv_x1_sg U42832 ( .A(reg_www_12[4]), .X(n50168) );
  inv_x1_sg U42833 ( .A(reg_ww_12[4]), .X(n52672) );
  inv_x1_sg U42834 ( .A(reg_www_12[5]), .X(n50166) );
  inv_x1_sg U42835 ( .A(reg_ww_12[5]), .X(n52670) );
  inv_x1_sg U42836 ( .A(reg_www_12[6]), .X(n50164) );
  inv_x1_sg U42837 ( .A(reg_ww_12[6]), .X(n52668) );
  inv_x1_sg U42838 ( .A(reg_www_12[7]), .X(n50162) );
  inv_x1_sg U42839 ( .A(reg_ww_12[7]), .X(n52666) );
  inv_x1_sg U42840 ( .A(reg_www_12[8]), .X(n50160) );
  inv_x1_sg U42841 ( .A(reg_ww_12[8]), .X(n52664) );
  inv_x1_sg U42842 ( .A(reg_www_12[9]), .X(n50158) );
  inv_x1_sg U42843 ( .A(reg_ww_12[9]), .X(n52662) );
  inv_x1_sg U42844 ( .A(reg_www_12[10]), .X(n50156) );
  inv_x1_sg U42845 ( .A(reg_ww_12[10]), .X(n52660) );
  inv_x1_sg U42846 ( .A(reg_www_12[11]), .X(n50154) );
  inv_x1_sg U42847 ( .A(reg_ww_12[11]), .X(n52658) );
  inv_x1_sg U42848 ( .A(reg_www_12[12]), .X(n50152) );
  inv_x1_sg U42849 ( .A(reg_ww_12[12]), .X(n52656) );
  inv_x1_sg U42850 ( .A(reg_www_12[13]), .X(n50150) );
  inv_x1_sg U42851 ( .A(reg_ww_12[13]), .X(n52654) );
  inv_x1_sg U42852 ( .A(reg_www_12[14]), .X(n50148) );
  inv_x1_sg U42853 ( .A(reg_ww_12[14]), .X(n52652) );
  inv_x1_sg U42854 ( .A(reg_www_12[15]), .X(n50146) );
  inv_x1_sg U42855 ( .A(reg_ww_12[15]), .X(n52650) );
  inv_x1_sg U42856 ( .A(reg_www_12[16]), .X(n50144) );
  inv_x1_sg U42857 ( .A(reg_ww_12[16]), .X(n52648) );
  inv_x1_sg U42858 ( .A(reg_www_12[17]), .X(n50142) );
  inv_x1_sg U42859 ( .A(reg_ww_12[17]), .X(n52646) );
  inv_x1_sg U42860 ( .A(reg_www_12[18]), .X(n50140) );
  inv_x1_sg U42861 ( .A(reg_ww_12[18]), .X(n52644) );
  inv_x1_sg U42862 ( .A(reg_www_12[19]), .X(n50138) );
  inv_x1_sg U42863 ( .A(reg_ww_12[19]), .X(n52642) );
  inv_x1_sg U42864 ( .A(reg_www_13[0]), .X(n50136) );
  inv_x1_sg U42865 ( .A(reg_ww_13[0]), .X(n52640) );
  inv_x1_sg U42866 ( .A(reg_www_13[1]), .X(n50134) );
  inv_x1_sg U42867 ( .A(reg_ww_13[1]), .X(n52638) );
  inv_x1_sg U42868 ( .A(reg_www_13[2]), .X(n50132) );
  inv_x1_sg U42869 ( .A(reg_ww_13[2]), .X(n52636) );
  inv_x1_sg U42870 ( .A(reg_www_13[3]), .X(n50130) );
  inv_x1_sg U42871 ( .A(reg_ww_13[3]), .X(n52634) );
  inv_x1_sg U42872 ( .A(reg_www_13[4]), .X(n50128) );
  inv_x1_sg U42873 ( .A(reg_ww_13[4]), .X(n52632) );
  inv_x1_sg U42874 ( .A(reg_www_13[5]), .X(n50126) );
  inv_x1_sg U42875 ( .A(reg_ww_13[5]), .X(n52630) );
  inv_x1_sg U42876 ( .A(reg_www_13[6]), .X(n50124) );
  inv_x1_sg U42877 ( .A(reg_ww_13[6]), .X(n52628) );
  inv_x1_sg U42878 ( .A(reg_www_13[7]), .X(n50122) );
  inv_x1_sg U42879 ( .A(reg_ww_13[7]), .X(n52626) );
  inv_x1_sg U42880 ( .A(reg_www_13[8]), .X(n50120) );
  inv_x1_sg U42881 ( .A(reg_ww_13[8]), .X(n52624) );
  inv_x1_sg U42882 ( .A(reg_www_13[9]), .X(n50118) );
  inv_x1_sg U42883 ( .A(reg_ww_13[9]), .X(n52622) );
  inv_x1_sg U42884 ( .A(reg_www_13[10]), .X(n50116) );
  inv_x1_sg U42885 ( .A(reg_ww_13[10]), .X(n52620) );
  inv_x1_sg U42886 ( .A(reg_www_13[11]), .X(n50114) );
  inv_x1_sg U42887 ( .A(reg_ww_13[11]), .X(n52618) );
  inv_x1_sg U42888 ( .A(reg_www_13[12]), .X(n50112) );
  inv_x1_sg U42889 ( .A(reg_ww_13[12]), .X(n52616) );
  inv_x1_sg U42890 ( .A(reg_www_13[13]), .X(n50110) );
  inv_x1_sg U42891 ( .A(reg_ww_13[13]), .X(n52614) );
  inv_x1_sg U42892 ( .A(reg_www_3[16]), .X(n50108) );
  inv_x1_sg U42893 ( .A(reg_ww_3[16]), .X(n52612) );
  inv_x1_sg U42894 ( .A(reg_www_3[17]), .X(n50106) );
  inv_x1_sg U42895 ( .A(reg_ww_3[17]), .X(n52610) );
  inv_x1_sg U42896 ( .A(reg_www_3[18]), .X(n50104) );
  inv_x1_sg U42897 ( .A(reg_ww_3[18]), .X(n52608) );
  inv_x1_sg U42898 ( .A(reg_www_3[19]), .X(n50102) );
  inv_x1_sg U42899 ( .A(reg_ww_3[19]), .X(n52606) );
  inv_x1_sg U42900 ( .A(reg_www_4[0]), .X(n50100) );
  inv_x1_sg U42901 ( .A(reg_ww_4[0]), .X(n52604) );
  inv_x1_sg U42902 ( .A(reg_www_4[1]), .X(n50098) );
  inv_x1_sg U42903 ( .A(reg_ww_4[1]), .X(n52602) );
  inv_x1_sg U42904 ( .A(reg_www_4[2]), .X(n50096) );
  inv_x1_sg U42905 ( .A(reg_ww_4[2]), .X(n52600) );
  inv_x1_sg U42906 ( .A(reg_www_4[3]), .X(n50094) );
  inv_x1_sg U42907 ( .A(reg_ww_4[3]), .X(n52598) );
  inv_x1_sg U42908 ( .A(reg_www_4[4]), .X(n50092) );
  inv_x1_sg U42909 ( .A(reg_ww_4[4]), .X(n52596) );
  inv_x1_sg U42910 ( .A(reg_www_4[5]), .X(n50090) );
  inv_x1_sg U42911 ( .A(reg_ww_4[5]), .X(n52594) );
  inv_x1_sg U42912 ( .A(reg_www_4[6]), .X(n50088) );
  inv_x1_sg U42913 ( .A(reg_ww_4[6]), .X(n52592) );
  inv_x1_sg U42914 ( .A(reg_www_4[7]), .X(n50086) );
  inv_x1_sg U42915 ( .A(reg_ww_4[7]), .X(n52590) );
  inv_x1_sg U42916 ( .A(reg_www_4[8]), .X(n50084) );
  inv_x1_sg U42917 ( .A(reg_ww_4[8]), .X(n52588) );
  inv_x1_sg U42918 ( .A(reg_www_4[9]), .X(n50082) );
  inv_x1_sg U42919 ( .A(reg_ww_4[9]), .X(n52586) );
  inv_x1_sg U42920 ( .A(reg_www_4[10]), .X(n50080) );
  inv_x1_sg U42921 ( .A(reg_ww_4[10]), .X(n52584) );
  inv_x1_sg U42922 ( .A(reg_www_4[11]), .X(n50078) );
  inv_x1_sg U42923 ( .A(reg_ww_4[11]), .X(n52582) );
  inv_x1_sg U42924 ( .A(reg_www_4[12]), .X(n50076) );
  inv_x1_sg U42925 ( .A(reg_ww_4[12]), .X(n52580) );
  inv_x1_sg U42926 ( .A(reg_www_4[13]), .X(n50074) );
  inv_x1_sg U42927 ( .A(reg_ww_4[13]), .X(n52578) );
  inv_x1_sg U42928 ( .A(reg_www_4[14]), .X(n50072) );
  inv_x1_sg U42929 ( .A(reg_ww_4[14]), .X(n52576) );
  inv_x1_sg U42930 ( .A(reg_www_4[15]), .X(n50070) );
  inv_x1_sg U42931 ( .A(reg_ww_4[15]), .X(n52574) );
  inv_x1_sg U42932 ( .A(reg_www_4[16]), .X(n50068) );
  inv_x1_sg U42933 ( .A(reg_ww_4[16]), .X(n52572) );
  inv_x1_sg U42934 ( .A(reg_www_4[17]), .X(n50066) );
  inv_x1_sg U42935 ( .A(reg_ww_4[17]), .X(n52570) );
  inv_x1_sg U42936 ( .A(reg_www_4[18]), .X(n50064) );
  inv_x1_sg U42937 ( .A(reg_ww_4[18]), .X(n52568) );
  inv_x1_sg U42938 ( .A(reg_www_4[19]), .X(n50062) );
  inv_x1_sg U42939 ( .A(reg_ww_4[19]), .X(n52566) );
  inv_x1_sg U42940 ( .A(reg_www_5[0]), .X(n50060) );
  inv_x1_sg U42941 ( .A(reg_ww_5[0]), .X(n52564) );
  inv_x1_sg U42942 ( .A(reg_www_5[1]), .X(n50058) );
  inv_x1_sg U42943 ( .A(reg_ww_5[1]), .X(n52562) );
  inv_x1_sg U42944 ( .A(reg_www_5[2]), .X(n50056) );
  inv_x1_sg U42945 ( .A(reg_ww_5[2]), .X(n52560) );
  inv_x1_sg U42946 ( .A(reg_www_5[3]), .X(n50054) );
  inv_x1_sg U42947 ( .A(reg_ww_5[3]), .X(n52558) );
  inv_x1_sg U42948 ( .A(reg_www_5[4]), .X(n50052) );
  inv_x1_sg U42949 ( .A(reg_ww_5[4]), .X(n52556) );
  inv_x1_sg U42950 ( .A(reg_www_5[5]), .X(n50050) );
  inv_x1_sg U42951 ( .A(reg_ww_5[5]), .X(n52554) );
  inv_x1_sg U42952 ( .A(reg_www_5[6]), .X(n50048) );
  inv_x1_sg U42953 ( .A(reg_ww_5[6]), .X(n52552) );
  inv_x1_sg U42954 ( .A(reg_www_5[7]), .X(n50046) );
  inv_x1_sg U42955 ( .A(reg_ww_5[7]), .X(n52550) );
  inv_x1_sg U42956 ( .A(reg_www_5[8]), .X(n50044) );
  inv_x1_sg U42957 ( .A(reg_ww_5[8]), .X(n52548) );
  inv_x1_sg U42958 ( .A(reg_www_5[9]), .X(n50042) );
  inv_x1_sg U42959 ( .A(reg_ww_5[9]), .X(n52546) );
  inv_x1_sg U42960 ( .A(reg_www_5[10]), .X(n50040) );
  inv_x1_sg U42961 ( .A(reg_ww_5[10]), .X(n52544) );
  inv_x1_sg U42962 ( .A(reg_www_5[11]), .X(n50038) );
  inv_x1_sg U42963 ( .A(reg_ww_5[11]), .X(n52542) );
  inv_x1_sg U42964 ( .A(reg_www_5[12]), .X(n50036) );
  inv_x1_sg U42965 ( .A(reg_ww_5[12]), .X(n52540) );
  inv_x1_sg U42966 ( .A(reg_www_5[13]), .X(n50034) );
  inv_x1_sg U42967 ( .A(reg_ww_5[13]), .X(n52538) );
  inv_x1_sg U42968 ( .A(reg_www_5[14]), .X(n50032) );
  inv_x1_sg U42969 ( .A(reg_ww_5[14]), .X(n52536) );
  inv_x1_sg U42970 ( .A(reg_www_5[15]), .X(n50030) );
  inv_x1_sg U42971 ( .A(reg_ww_5[15]), .X(n52534) );
  inv_x1_sg U42972 ( .A(reg_www_5[16]), .X(n50028) );
  inv_x1_sg U42973 ( .A(reg_ww_5[16]), .X(n52532) );
  inv_x1_sg U42974 ( .A(reg_www_5[17]), .X(n50026) );
  inv_x1_sg U42975 ( .A(reg_ww_5[17]), .X(n52530) );
  inv_x1_sg U42976 ( .A(reg_www_5[18]), .X(n50024) );
  inv_x1_sg U42977 ( .A(reg_ww_5[18]), .X(n52528) );
  inv_x1_sg U42978 ( .A(reg_www_5[19]), .X(n50022) );
  inv_x1_sg U42979 ( .A(reg_ww_5[19]), .X(n52526) );
  inv_x1_sg U42980 ( .A(reg_www_6[0]), .X(n50020) );
  inv_x1_sg U42981 ( .A(reg_ww_6[0]), .X(n52524) );
  inv_x1_sg U42982 ( .A(reg_www_6[1]), .X(n50018) );
  inv_x1_sg U42983 ( .A(reg_ww_6[1]), .X(n52522) );
  inv_x1_sg U42984 ( .A(reg_www_6[2]), .X(n50016) );
  inv_x1_sg U42985 ( .A(reg_ww_6[2]), .X(n52520) );
  inv_x1_sg U42986 ( .A(reg_www_6[3]), .X(n50014) );
  inv_x1_sg U42987 ( .A(reg_ww_6[3]), .X(n52518) );
  inv_x1_sg U42988 ( .A(reg_www_6[4]), .X(n50012) );
  inv_x1_sg U42989 ( .A(reg_ww_6[4]), .X(n52516) );
  inv_x1_sg U42990 ( .A(reg_www_6[5]), .X(n50010) );
  inv_x1_sg U42991 ( .A(reg_ww_6[5]), .X(n52514) );
  inv_x1_sg U42992 ( .A(reg_www_6[6]), .X(n50008) );
  inv_x1_sg U42993 ( .A(reg_ww_6[6]), .X(n52512) );
  inv_x1_sg U42994 ( .A(reg_www_6[7]), .X(n50006) );
  inv_x1_sg U42995 ( .A(reg_ww_6[7]), .X(n52510) );
  inv_x1_sg U42996 ( .A(reg_www_6[8]), .X(n50004) );
  inv_x1_sg U42997 ( .A(reg_ww_6[8]), .X(n52508) );
  inv_x1_sg U42998 ( .A(reg_www_6[9]), .X(n50002) );
  inv_x1_sg U42999 ( .A(reg_ww_6[9]), .X(n52506) );
  inv_x1_sg U43000 ( .A(reg_www_6[10]), .X(n50000) );
  inv_x1_sg U43001 ( .A(reg_ww_6[10]), .X(n52504) );
  inv_x1_sg U43002 ( .A(reg_www_6[11]), .X(n49998) );
  inv_x1_sg U43003 ( .A(reg_ww_6[11]), .X(n52502) );
  inv_x1_sg U43004 ( .A(reg_www_6[12]), .X(n49996) );
  inv_x1_sg U43005 ( .A(reg_ww_6[12]), .X(n52500) );
  inv_x1_sg U43006 ( .A(reg_www_6[13]), .X(n49994) );
  inv_x1_sg U43007 ( .A(reg_ww_6[13]), .X(n52498) );
  inv_x1_sg U43008 ( .A(reg_www_6[14]), .X(n49992) );
  inv_x1_sg U43009 ( .A(reg_ww_6[14]), .X(n52496) );
  inv_x1_sg U43010 ( .A(reg_www_6[15]), .X(n49990) );
  inv_x1_sg U43011 ( .A(reg_ww_6[15]), .X(n52494) );
  inv_x1_sg U43012 ( .A(reg_www_6[16]), .X(n49988) );
  inv_x1_sg U43013 ( .A(reg_ww_6[16]), .X(n52492) );
  inv_x1_sg U43014 ( .A(reg_www_6[17]), .X(n49986) );
  inv_x1_sg U43015 ( .A(reg_ww_6[17]), .X(n52490) );
  inv_x1_sg U43016 ( .A(reg_www_6[18]), .X(n49984) );
  inv_x1_sg U43017 ( .A(reg_ww_6[18]), .X(n52488) );
  inv_x1_sg U43018 ( .A(reg_www_6[19]), .X(n49982) );
  inv_x1_sg U43019 ( .A(reg_ww_6[19]), .X(n52486) );
  inv_x1_sg U43020 ( .A(reg_www_7[0]), .X(n49980) );
  inv_x1_sg U43021 ( .A(reg_ww_7[0]), .X(n52484) );
  inv_x1_sg U43022 ( .A(reg_www_7[1]), .X(n49978) );
  inv_x1_sg U43023 ( .A(reg_ww_7[1]), .X(n52482) );
  inv_x1_sg U43024 ( .A(reg_www_7[2]), .X(n49976) );
  inv_x1_sg U43025 ( .A(reg_ww_7[2]), .X(n52480) );
  inv_x1_sg U43026 ( .A(reg_www_7[3]), .X(n49974) );
  inv_x1_sg U43027 ( .A(reg_ww_7[3]), .X(n52478) );
  inv_x1_sg U43028 ( .A(reg_www_7[4]), .X(n49972) );
  inv_x1_sg U43029 ( .A(reg_ww_7[4]), .X(n52476) );
  inv_x1_sg U43030 ( .A(reg_www_7[5]), .X(n49970) );
  inv_x1_sg U43031 ( .A(reg_ww_7[5]), .X(n52474) );
  inv_x1_sg U43032 ( .A(reg_www_7[6]), .X(n49968) );
  inv_x1_sg U43033 ( .A(reg_ww_7[6]), .X(n52472) );
  inv_x1_sg U43034 ( .A(reg_www_7[7]), .X(n49966) );
  inv_x1_sg U43035 ( .A(reg_ww_7[7]), .X(n52470) );
  inv_x1_sg U43036 ( .A(reg_www_7[8]), .X(n49964) );
  inv_x1_sg U43037 ( .A(reg_ww_7[8]), .X(n52468) );
  inv_x1_sg U43038 ( .A(reg_www_7[9]), .X(n49962) );
  inv_x1_sg U43039 ( .A(reg_ww_7[9]), .X(n52466) );
  inv_x1_sg U43040 ( .A(reg_www_7[10]), .X(n49960) );
  inv_x1_sg U43041 ( .A(reg_ww_7[10]), .X(n52464) );
  inv_x1_sg U43042 ( .A(reg_www_7[11]), .X(n49958) );
  inv_x1_sg U43043 ( .A(reg_ww_7[11]), .X(n52462) );
  inv_x1_sg U43044 ( .A(reg_www_7[12]), .X(n49956) );
  inv_x1_sg U43045 ( .A(reg_ww_7[12]), .X(n52460) );
  inv_x1_sg U43046 ( .A(reg_www_7[13]), .X(n49954) );
  inv_x1_sg U43047 ( .A(reg_ww_7[13]), .X(n52458) );
  inv_x1_sg U43048 ( .A(reg_www_7[14]), .X(n49952) );
  inv_x1_sg U43049 ( .A(reg_ww_7[14]), .X(n52456) );
  inv_x1_sg U43050 ( .A(reg_www_7[15]), .X(n49950) );
  inv_x1_sg U43051 ( .A(reg_ww_7[15]), .X(n52454) );
  inv_x1_sg U43052 ( .A(reg_www_7[16]), .X(n49948) );
  inv_x1_sg U43053 ( .A(reg_ww_7[16]), .X(n52452) );
  inv_x1_sg U43054 ( .A(reg_www_7[17]), .X(n49946) );
  inv_x1_sg U43055 ( .A(reg_ww_7[17]), .X(n52450) );
  inv_x1_sg U43056 ( .A(reg_www_7[18]), .X(n49944) );
  inv_x1_sg U43057 ( .A(reg_ww_7[18]), .X(n52448) );
  inv_x1_sg U43058 ( .A(reg_www_7[19]), .X(n49942) );
  inv_x1_sg U43059 ( .A(reg_ww_7[19]), .X(n52446) );
  inv_x1_sg U43060 ( .A(reg_www_8[0]), .X(n49940) );
  inv_x1_sg U43061 ( .A(reg_ww_8[0]), .X(n52444) );
  inv_x1_sg U43062 ( .A(reg_www_8[1]), .X(n49938) );
  inv_x1_sg U43063 ( .A(reg_ww_8[1]), .X(n52442) );
  inv_x1_sg U43064 ( .A(reg_www_8[2]), .X(n49936) );
  inv_x1_sg U43065 ( .A(reg_ww_8[2]), .X(n52440) );
  inv_x1_sg U43066 ( .A(reg_www_8[3]), .X(n49934) );
  inv_x1_sg U43067 ( .A(reg_ww_8[3]), .X(n52438) );
  inv_x1_sg U43068 ( .A(reg_www_8[4]), .X(n49932) );
  inv_x1_sg U43069 ( .A(reg_ww_8[4]), .X(n52436) );
  inv_x1_sg U43070 ( .A(reg_www_8[5]), .X(n49930) );
  inv_x1_sg U43071 ( .A(reg_ww_8[5]), .X(n52434) );
  inv_x1_sg U43072 ( .A(reg_www_8[6]), .X(n49928) );
  inv_x1_sg U43073 ( .A(reg_ww_8[6]), .X(n52432) );
  inv_x1_sg U43074 ( .A(reg_www_8[7]), .X(n49926) );
  inv_x1_sg U43075 ( .A(reg_ww_8[7]), .X(n52430) );
  inv_x1_sg U43076 ( .A(reg_www_8[8]), .X(n49924) );
  inv_x1_sg U43077 ( .A(reg_ww_8[8]), .X(n52428) );
  inv_x1_sg U43078 ( .A(reg_www_8[9]), .X(n49922) );
  inv_x1_sg U43079 ( .A(reg_ww_8[9]), .X(n52426) );
  inv_x1_sg U43080 ( .A(reg_www_8[10]), .X(n49920) );
  inv_x1_sg U43081 ( .A(reg_ww_8[10]), .X(n52424) );
  inv_x1_sg U43082 ( .A(reg_www_8[11]), .X(n49918) );
  inv_x1_sg U43083 ( .A(reg_ww_8[11]), .X(n52422) );
  inv_x1_sg U43084 ( .A(reg_www_8[12]), .X(n49916) );
  inv_x1_sg U43085 ( .A(reg_ww_8[12]), .X(n52420) );
  inv_x1_sg U43086 ( .A(reg_www_8[13]), .X(n49914) );
  inv_x1_sg U43087 ( .A(reg_ww_8[13]), .X(n52418) );
  inv_x1_sg U43088 ( .A(reg_www_8[14]), .X(n49912) );
  inv_x1_sg U43089 ( .A(reg_ww_8[14]), .X(n52416) );
  inv_x1_sg U43090 ( .A(reg_iii_14[17]), .X(n49910) );
  inv_x1_sg U43091 ( .A(reg_ii_14[17]), .X(n52414) );
  inv_x1_sg U43092 ( .A(reg_iii_14[18]), .X(n49908) );
  inv_x1_sg U43093 ( .A(reg_ii_14[18]), .X(n52412) );
  inv_x1_sg U43094 ( .A(reg_iii_14[19]), .X(n49906) );
  inv_x1_sg U43095 ( .A(reg_ii_14[19]), .X(n52410) );
  inv_x1_sg U43096 ( .A(reg_iii_15[0]), .X(n49904) );
  inv_x1_sg U43097 ( .A(reg_ii_15[0]), .X(n52408) );
  inv_x1_sg U43098 ( .A(reg_iii_15[1]), .X(n49902) );
  inv_x1_sg U43099 ( .A(reg_ii_15[1]), .X(n52406) );
  inv_x1_sg U43100 ( .A(reg_iii_15[2]), .X(n49900) );
  inv_x1_sg U43101 ( .A(reg_ii_15[2]), .X(n52404) );
  inv_x1_sg U43102 ( .A(reg_iii_15[3]), .X(n49898) );
  inv_x1_sg U43103 ( .A(reg_ii_15[3]), .X(n52402) );
  inv_x1_sg U43104 ( .A(reg_iii_15[4]), .X(n49896) );
  inv_x1_sg U43105 ( .A(reg_ii_15[4]), .X(n52400) );
  inv_x1_sg U43106 ( .A(reg_iii_15[5]), .X(n49894) );
  inv_x1_sg U43107 ( .A(reg_ii_15[5]), .X(n52398) );
  inv_x1_sg U43108 ( .A(reg_iii_15[6]), .X(n49892) );
  inv_x1_sg U43109 ( .A(reg_ii_15[6]), .X(n52396) );
  inv_x1_sg U43110 ( .A(reg_iii_15[7]), .X(n49890) );
  inv_x1_sg U43111 ( .A(reg_ii_15[7]), .X(n52394) );
  inv_x1_sg U43112 ( .A(reg_iii_15[8]), .X(n49888) );
  inv_x1_sg U43113 ( .A(reg_ii_15[8]), .X(n52392) );
  inv_x1_sg U43114 ( .A(reg_iii_15[9]), .X(n49886) );
  inv_x1_sg U43115 ( .A(reg_ii_15[9]), .X(n52390) );
  inv_x1_sg U43116 ( .A(reg_iii_15[10]), .X(n49884) );
  inv_x1_sg U43117 ( .A(reg_ii_15[10]), .X(n52388) );
  inv_x1_sg U43118 ( .A(reg_iii_15[11]), .X(n49882) );
  inv_x1_sg U43119 ( .A(reg_ii_15[11]), .X(n52386) );
  inv_x1_sg U43120 ( .A(reg_iii_15[12]), .X(n49880) );
  inv_x1_sg U43121 ( .A(reg_ii_15[12]), .X(n52384) );
  inv_x1_sg U43122 ( .A(reg_iii_15[13]), .X(n49878) );
  inv_x1_sg U43123 ( .A(reg_ii_15[13]), .X(n52382) );
  inv_x1_sg U43124 ( .A(reg_iii_15[14]), .X(n49876) );
  inv_x1_sg U43125 ( .A(reg_ii_15[14]), .X(n52380) );
  inv_x1_sg U43126 ( .A(reg_iii_15[15]), .X(n49874) );
  inv_x1_sg U43127 ( .A(reg_ii_15[15]), .X(n52378) );
  inv_x1_sg U43128 ( .A(reg_iii_15[16]), .X(n49872) );
  inv_x1_sg U43129 ( .A(reg_ii_15[16]), .X(n52376) );
  inv_x1_sg U43130 ( .A(reg_iii_15[17]), .X(n49870) );
  inv_x1_sg U43131 ( .A(reg_ii_15[17]), .X(n52374) );
  inv_x1_sg U43132 ( .A(reg_iii_15[18]), .X(n49868) );
  inv_x1_sg U43133 ( .A(reg_ii_15[18]), .X(n52372) );
  inv_x1_sg U43134 ( .A(reg_iii_15[19]), .X(n49866) );
  inv_x1_sg U43135 ( .A(reg_ii_15[19]), .X(n52370) );
  inv_x1_sg U43136 ( .A(reg_www_0[0]), .X(n49864) );
  inv_x1_sg U43137 ( .A(reg_ww_0[0]), .X(n52368) );
  inv_x1_sg U43138 ( .A(reg_www_0[1]), .X(n49862) );
  inv_x1_sg U43139 ( .A(reg_ww_0[1]), .X(n52366) );
  inv_x1_sg U43140 ( .A(reg_www_0[2]), .X(n49860) );
  inv_x1_sg U43141 ( .A(reg_ww_0[2]), .X(n52364) );
  inv_x1_sg U43142 ( .A(reg_www_0[3]), .X(n49858) );
  inv_x1_sg U43143 ( .A(reg_ww_0[3]), .X(n52362) );
  inv_x1_sg U43144 ( .A(reg_www_0[4]), .X(n49856) );
  inv_x1_sg U43145 ( .A(reg_ww_0[4]), .X(n52360) );
  inv_x1_sg U43146 ( .A(reg_www_0[5]), .X(n49854) );
  inv_x1_sg U43147 ( .A(reg_ww_0[5]), .X(n52358) );
  inv_x1_sg U43148 ( .A(reg_www_0[6]), .X(n49852) );
  inv_x1_sg U43149 ( .A(reg_ww_0[6]), .X(n52356) );
  inv_x1_sg U43150 ( .A(reg_www_0[7]), .X(n49850) );
  inv_x1_sg U43151 ( .A(reg_ww_0[7]), .X(n52354) );
  inv_x1_sg U43152 ( .A(reg_www_0[8]), .X(n49848) );
  inv_x1_sg U43153 ( .A(reg_ww_0[8]), .X(n52352) );
  inv_x1_sg U43154 ( .A(reg_www_0[9]), .X(n49846) );
  inv_x1_sg U43155 ( .A(reg_ww_0[9]), .X(n52350) );
  inv_x1_sg U43156 ( .A(reg_www_0[10]), .X(n49844) );
  inv_x1_sg U43157 ( .A(reg_ww_0[10]), .X(n52348) );
  inv_x1_sg U43158 ( .A(reg_www_0[11]), .X(n49842) );
  inv_x1_sg U43159 ( .A(reg_ww_0[11]), .X(n52346) );
  inv_x1_sg U43160 ( .A(reg_www_0[12]), .X(n49840) );
  inv_x1_sg U43161 ( .A(reg_ww_0[12]), .X(n52344) );
  inv_x1_sg U43162 ( .A(reg_www_0[13]), .X(n49838) );
  inv_x1_sg U43163 ( .A(reg_ww_0[13]), .X(n52342) );
  inv_x1_sg U43164 ( .A(reg_www_0[14]), .X(n49836) );
  inv_x1_sg U43165 ( .A(reg_ww_0[14]), .X(n52340) );
  inv_x1_sg U43166 ( .A(reg_www_0[15]), .X(n49834) );
  inv_x1_sg U43167 ( .A(reg_ww_0[15]), .X(n52338) );
  inv_x1_sg U43168 ( .A(reg_www_0[16]), .X(n49832) );
  inv_x1_sg U43169 ( .A(reg_ww_0[16]), .X(n52336) );
  inv_x1_sg U43170 ( .A(reg_www_0[17]), .X(n49830) );
  inv_x1_sg U43171 ( .A(reg_ww_0[17]), .X(n52334) );
  inv_x1_sg U43172 ( .A(reg_www_0[18]), .X(n49828) );
  inv_x1_sg U43173 ( .A(reg_ww_0[18]), .X(n52332) );
  inv_x1_sg U43174 ( .A(reg_www_0[19]), .X(n49826) );
  inv_x1_sg U43175 ( .A(reg_ww_0[19]), .X(n52330) );
  inv_x1_sg U43176 ( .A(reg_www_1[0]), .X(n49824) );
  inv_x1_sg U43177 ( .A(reg_ww_1[0]), .X(n52328) );
  inv_x1_sg U43178 ( .A(reg_www_1[1]), .X(n49822) );
  inv_x1_sg U43179 ( .A(reg_ww_1[1]), .X(n52326) );
  inv_x1_sg U43180 ( .A(reg_www_1[2]), .X(n49820) );
  inv_x1_sg U43181 ( .A(reg_ww_1[2]), .X(n52324) );
  inv_x1_sg U43182 ( .A(reg_www_1[3]), .X(n49818) );
  inv_x1_sg U43183 ( .A(reg_ww_1[3]), .X(n52322) );
  inv_x1_sg U43184 ( .A(reg_www_1[4]), .X(n49816) );
  inv_x1_sg U43185 ( .A(reg_ww_1[4]), .X(n52320) );
  inv_x1_sg U43186 ( .A(reg_www_1[5]), .X(n49814) );
  inv_x1_sg U43187 ( .A(reg_ww_1[5]), .X(n52318) );
  inv_x1_sg U43188 ( .A(reg_www_1[6]), .X(n49812) );
  inv_x1_sg U43189 ( .A(reg_ww_1[6]), .X(n52316) );
  inv_x1_sg U43190 ( .A(reg_www_1[7]), .X(n49810) );
  inv_x1_sg U43191 ( .A(reg_ww_1[7]), .X(n52314) );
  inv_x1_sg U43192 ( .A(reg_www_1[8]), .X(n49808) );
  inv_x1_sg U43193 ( .A(reg_ww_1[8]), .X(n52312) );
  inv_x1_sg U43194 ( .A(reg_www_1[9]), .X(n49806) );
  inv_x1_sg U43195 ( .A(reg_ww_1[9]), .X(n52310) );
  inv_x1_sg U43196 ( .A(reg_www_1[10]), .X(n49804) );
  inv_x1_sg U43197 ( .A(reg_ww_1[10]), .X(n52308) );
  inv_x1_sg U43198 ( .A(reg_www_1[11]), .X(n49802) );
  inv_x1_sg U43199 ( .A(reg_ww_1[11]), .X(n52306) );
  inv_x1_sg U43200 ( .A(reg_www_1[12]), .X(n49800) );
  inv_x1_sg U43201 ( .A(reg_ww_1[12]), .X(n52304) );
  inv_x1_sg U43202 ( .A(reg_www_1[13]), .X(n49798) );
  inv_x1_sg U43203 ( .A(reg_ww_1[13]), .X(n52302) );
  inv_x1_sg U43204 ( .A(reg_www_1[14]), .X(n49796) );
  inv_x1_sg U43205 ( .A(reg_ww_1[14]), .X(n52300) );
  inv_x1_sg U43206 ( .A(reg_www_1[15]), .X(n49794) );
  inv_x1_sg U43207 ( .A(reg_ww_1[15]), .X(n52298) );
  inv_x1_sg U43208 ( .A(reg_www_1[16]), .X(n49792) );
  inv_x1_sg U43209 ( .A(reg_ww_1[16]), .X(n52296) );
  inv_x1_sg U43210 ( .A(reg_www_1[17]), .X(n49790) );
  inv_x1_sg U43211 ( .A(reg_ww_1[17]), .X(n52294) );
  inv_x1_sg U43212 ( .A(reg_www_1[18]), .X(n49788) );
  inv_x1_sg U43213 ( .A(reg_ww_1[18]), .X(n52292) );
  inv_x1_sg U43214 ( .A(reg_www_1[19]), .X(n49786) );
  inv_x1_sg U43215 ( .A(reg_ww_1[19]), .X(n52290) );
  inv_x1_sg U43216 ( .A(reg_www_2[0]), .X(n49784) );
  inv_x1_sg U43217 ( .A(reg_ww_2[0]), .X(n52288) );
  inv_x1_sg U43218 ( .A(reg_www_2[1]), .X(n49782) );
  inv_x1_sg U43219 ( .A(reg_ww_2[1]), .X(n52286) );
  inv_x1_sg U43220 ( .A(reg_www_2[2]), .X(n49780) );
  inv_x1_sg U43221 ( .A(reg_ww_2[2]), .X(n52284) );
  inv_x1_sg U43222 ( .A(reg_www_2[3]), .X(n49778) );
  inv_x1_sg U43223 ( .A(reg_ww_2[3]), .X(n52282) );
  inv_x1_sg U43224 ( .A(reg_www_2[4]), .X(n49776) );
  inv_x1_sg U43225 ( .A(reg_ww_2[4]), .X(n52280) );
  inv_x1_sg U43226 ( .A(reg_www_2[5]), .X(n49774) );
  inv_x1_sg U43227 ( .A(reg_ww_2[5]), .X(n52278) );
  inv_x1_sg U43228 ( .A(reg_www_2[6]), .X(n49772) );
  inv_x1_sg U43229 ( .A(reg_ww_2[6]), .X(n52276) );
  inv_x1_sg U43230 ( .A(reg_www_2[7]), .X(n49770) );
  inv_x1_sg U43231 ( .A(reg_ww_2[7]), .X(n52274) );
  inv_x1_sg U43232 ( .A(reg_www_2[8]), .X(n49768) );
  inv_x1_sg U43233 ( .A(reg_ww_2[8]), .X(n52272) );
  inv_x1_sg U43234 ( .A(reg_www_2[9]), .X(n49766) );
  inv_x1_sg U43235 ( .A(reg_ww_2[9]), .X(n52270) );
  inv_x1_sg U43236 ( .A(reg_www_2[10]), .X(n49764) );
  inv_x1_sg U43237 ( .A(reg_ww_2[10]), .X(n52268) );
  inv_x1_sg U43238 ( .A(reg_www_2[11]), .X(n49762) );
  inv_x1_sg U43239 ( .A(reg_ww_2[11]), .X(n52266) );
  inv_x1_sg U43240 ( .A(reg_www_2[12]), .X(n49760) );
  inv_x1_sg U43241 ( .A(reg_ww_2[12]), .X(n52264) );
  inv_x1_sg U43242 ( .A(reg_www_2[13]), .X(n49758) );
  inv_x1_sg U43243 ( .A(reg_ww_2[13]), .X(n52262) );
  inv_x1_sg U43244 ( .A(reg_www_2[14]), .X(n49756) );
  inv_x1_sg U43245 ( .A(reg_ww_2[14]), .X(n52260) );
  inv_x1_sg U43246 ( .A(reg_www_2[15]), .X(n49754) );
  inv_x1_sg U43247 ( .A(reg_ww_2[15]), .X(n52258) );
  inv_x1_sg U43248 ( .A(reg_www_2[16]), .X(n49752) );
  inv_x1_sg U43249 ( .A(reg_ww_2[16]), .X(n52256) );
  inv_x1_sg U43250 ( .A(reg_www_2[17]), .X(n49750) );
  inv_x1_sg U43251 ( .A(reg_ww_2[17]), .X(n52254) );
  inv_x1_sg U43252 ( .A(reg_www_2[18]), .X(n49748) );
  inv_x1_sg U43253 ( .A(reg_ww_2[18]), .X(n52252) );
  inv_x1_sg U43254 ( .A(reg_www_2[19]), .X(n49746) );
  inv_x1_sg U43255 ( .A(reg_ww_2[19]), .X(n52250) );
  inv_x1_sg U43256 ( .A(reg_www_3[0]), .X(n49744) );
  inv_x1_sg U43257 ( .A(reg_ww_3[0]), .X(n52248) );
  inv_x1_sg U43258 ( .A(reg_www_3[1]), .X(n49742) );
  inv_x1_sg U43259 ( .A(reg_ww_3[1]), .X(n52246) );
  inv_x1_sg U43260 ( .A(reg_www_3[2]), .X(n49740) );
  inv_x1_sg U43261 ( .A(reg_ww_3[2]), .X(n52244) );
  inv_x1_sg U43262 ( .A(reg_www_3[3]), .X(n49738) );
  inv_x1_sg U43263 ( .A(reg_ww_3[3]), .X(n52242) );
  inv_x1_sg U43264 ( .A(reg_www_3[4]), .X(n49736) );
  inv_x1_sg U43265 ( .A(reg_ww_3[4]), .X(n52240) );
  inv_x1_sg U43266 ( .A(reg_www_3[5]), .X(n49734) );
  inv_x1_sg U43267 ( .A(reg_ww_3[5]), .X(n52238) );
  inv_x1_sg U43268 ( .A(reg_www_3[6]), .X(n49732) );
  inv_x1_sg U43269 ( .A(reg_ww_3[6]), .X(n52236) );
  inv_x1_sg U43270 ( .A(reg_www_3[7]), .X(n49730) );
  inv_x1_sg U43271 ( .A(reg_ww_3[7]), .X(n52234) );
  inv_x1_sg U43272 ( .A(reg_www_3[8]), .X(n49728) );
  inv_x1_sg U43273 ( .A(reg_ww_3[8]), .X(n52232) );
  inv_x1_sg U43274 ( .A(reg_www_3[9]), .X(n49726) );
  inv_x1_sg U43275 ( .A(reg_ww_3[9]), .X(n52230) );
  inv_x1_sg U43276 ( .A(reg_www_3[10]), .X(n49724) );
  inv_x1_sg U43277 ( .A(reg_ww_3[10]), .X(n52228) );
  inv_x1_sg U43278 ( .A(reg_www_3[11]), .X(n49722) );
  inv_x1_sg U43279 ( .A(reg_ww_3[11]), .X(n52226) );
  inv_x1_sg U43280 ( .A(reg_www_3[12]), .X(n49720) );
  inv_x1_sg U43281 ( .A(reg_ww_3[12]), .X(n52224) );
  inv_x1_sg U43282 ( .A(reg_www_3[13]), .X(n49718) );
  inv_x1_sg U43283 ( .A(reg_ww_3[13]), .X(n52222) );
  inv_x1_sg U43284 ( .A(reg_www_3[14]), .X(n49716) );
  inv_x1_sg U43285 ( .A(reg_ww_3[14]), .X(n52220) );
  inv_x1_sg U43286 ( .A(reg_www_3[15]), .X(n49714) );
  inv_x1_sg U43287 ( .A(reg_ww_3[15]), .X(n52218) );
  inv_x1_sg U43288 ( .A(reg_iii_9[18]), .X(n49712) );
  inv_x1_sg U43289 ( .A(reg_ii_9[18]), .X(n52216) );
  inv_x1_sg U43290 ( .A(reg_iii_9[19]), .X(n49710) );
  inv_x1_sg U43291 ( .A(reg_ii_9[19]), .X(n52214) );
  inv_x1_sg U43292 ( .A(reg_iii_10[0]), .X(n49708) );
  inv_x1_sg U43293 ( .A(reg_ii_10[0]), .X(n52212) );
  inv_x1_sg U43294 ( .A(reg_iii_10[1]), .X(n49706) );
  inv_x1_sg U43295 ( .A(reg_ii_10[1]), .X(n52210) );
  inv_x1_sg U43296 ( .A(reg_iii_10[2]), .X(n49704) );
  inv_x1_sg U43297 ( .A(reg_ii_10[2]), .X(n52208) );
  inv_x1_sg U43298 ( .A(reg_iii_10[3]), .X(n49702) );
  inv_x1_sg U43299 ( .A(reg_ii_10[3]), .X(n52206) );
  inv_x1_sg U43300 ( .A(reg_iii_10[4]), .X(n49700) );
  inv_x1_sg U43301 ( .A(reg_ii_10[4]), .X(n52204) );
  inv_x1_sg U43302 ( .A(reg_iii_10[5]), .X(n49698) );
  inv_x1_sg U43303 ( .A(reg_ii_10[5]), .X(n52202) );
  inv_x1_sg U43304 ( .A(reg_iii_10[6]), .X(n49696) );
  inv_x1_sg U43305 ( .A(reg_ii_10[6]), .X(n52200) );
  inv_x1_sg U43306 ( .A(reg_iii_10[7]), .X(n49694) );
  inv_x1_sg U43307 ( .A(reg_ii_10[7]), .X(n52198) );
  inv_x1_sg U43308 ( .A(reg_iii_10[8]), .X(n49692) );
  inv_x1_sg U43309 ( .A(reg_ii_10[8]), .X(n52196) );
  inv_x1_sg U43310 ( .A(reg_iii_10[9]), .X(n49690) );
  inv_x1_sg U43311 ( .A(reg_ii_10[9]), .X(n52194) );
  inv_x1_sg U43312 ( .A(reg_iii_10[10]), .X(n49688) );
  inv_x1_sg U43313 ( .A(reg_ii_10[10]), .X(n52192) );
  inv_x1_sg U43314 ( .A(reg_iii_10[11]), .X(n49686) );
  inv_x1_sg U43315 ( .A(reg_ii_10[11]), .X(n52190) );
  inv_x1_sg U43316 ( .A(reg_iii_10[12]), .X(n49684) );
  inv_x1_sg U43317 ( .A(reg_ii_10[12]), .X(n52188) );
  inv_x1_sg U43318 ( .A(reg_iii_10[13]), .X(n49682) );
  inv_x1_sg U43319 ( .A(reg_ii_10[13]), .X(n52186) );
  inv_x1_sg U43320 ( .A(reg_iii_10[14]), .X(n49680) );
  inv_x1_sg U43321 ( .A(reg_ii_10[14]), .X(n52184) );
  inv_x1_sg U43322 ( .A(reg_iii_10[15]), .X(n49678) );
  inv_x1_sg U43323 ( .A(reg_ii_10[15]), .X(n52182) );
  inv_x1_sg U43324 ( .A(reg_iii_10[16]), .X(n49676) );
  inv_x1_sg U43325 ( .A(reg_ii_10[16]), .X(n52180) );
  inv_x1_sg U43326 ( .A(reg_iii_10[17]), .X(n49674) );
  inv_x1_sg U43327 ( .A(reg_ii_10[17]), .X(n52178) );
  inv_x1_sg U43328 ( .A(reg_iii_10[18]), .X(n49672) );
  inv_x1_sg U43329 ( .A(reg_ii_10[18]), .X(n52176) );
  inv_x1_sg U43330 ( .A(reg_iii_10[19]), .X(n49670) );
  inv_x1_sg U43331 ( .A(reg_ii_10[19]), .X(n52174) );
  inv_x1_sg U43332 ( .A(reg_iii_11[0]), .X(n49668) );
  inv_x1_sg U43333 ( .A(reg_ii_11[0]), .X(n52172) );
  inv_x1_sg U43334 ( .A(reg_iii_11[1]), .X(n49666) );
  inv_x1_sg U43335 ( .A(reg_ii_11[1]), .X(n52170) );
  inv_x1_sg U43336 ( .A(reg_iii_11[2]), .X(n49664) );
  inv_x1_sg U43337 ( .A(reg_ii_11[2]), .X(n52168) );
  inv_x1_sg U43338 ( .A(reg_iii_11[3]), .X(n49662) );
  inv_x1_sg U43339 ( .A(reg_ii_11[3]), .X(n52166) );
  inv_x1_sg U43340 ( .A(reg_iii_11[4]), .X(n49660) );
  inv_x1_sg U43341 ( .A(reg_ii_11[4]), .X(n52164) );
  inv_x1_sg U43342 ( .A(reg_iii_11[5]), .X(n49658) );
  inv_x1_sg U43343 ( .A(reg_ii_11[5]), .X(n52162) );
  inv_x1_sg U43344 ( .A(reg_iii_11[6]), .X(n49656) );
  inv_x1_sg U43345 ( .A(reg_ii_11[6]), .X(n52160) );
  inv_x1_sg U43346 ( .A(reg_iii_11[7]), .X(n49654) );
  inv_x1_sg U43347 ( .A(reg_ii_11[7]), .X(n52158) );
  inv_x1_sg U43348 ( .A(reg_iii_11[8]), .X(n49652) );
  inv_x1_sg U43349 ( .A(reg_ii_11[8]), .X(n52156) );
  inv_x1_sg U43350 ( .A(reg_iii_11[9]), .X(n49650) );
  inv_x1_sg U43351 ( .A(reg_ii_11[9]), .X(n52154) );
  inv_x1_sg U43352 ( .A(reg_iii_11[10]), .X(n49648) );
  inv_x1_sg U43353 ( .A(reg_ii_11[10]), .X(n52152) );
  inv_x1_sg U43354 ( .A(reg_iii_11[11]), .X(n49646) );
  inv_x1_sg U43355 ( .A(reg_ii_11[11]), .X(n52150) );
  inv_x1_sg U43356 ( .A(reg_iii_11[12]), .X(n49644) );
  inv_x1_sg U43357 ( .A(reg_ii_11[12]), .X(n52148) );
  inv_x1_sg U43358 ( .A(reg_iii_11[13]), .X(n49642) );
  inv_x1_sg U43359 ( .A(reg_ii_11[13]), .X(n52146) );
  inv_x1_sg U43360 ( .A(reg_iii_11[14]), .X(n49640) );
  inv_x1_sg U43361 ( .A(reg_ii_11[14]), .X(n52144) );
  inv_x1_sg U43362 ( .A(reg_iii_11[15]), .X(n49638) );
  inv_x1_sg U43363 ( .A(reg_ii_11[15]), .X(n52142) );
  inv_x1_sg U43364 ( .A(reg_iii_11[16]), .X(n49636) );
  inv_x1_sg U43365 ( .A(reg_ii_11[16]), .X(n52140) );
  inv_x1_sg U43366 ( .A(reg_iii_11[17]), .X(n49634) );
  inv_x1_sg U43367 ( .A(reg_ii_11[17]), .X(n52138) );
  inv_x1_sg U43368 ( .A(reg_iii_11[18]), .X(n49632) );
  inv_x1_sg U43369 ( .A(reg_ii_11[18]), .X(n52136) );
  inv_x1_sg U43370 ( .A(reg_iii_11[19]), .X(n49630) );
  inv_x1_sg U43371 ( .A(reg_ii_11[19]), .X(n52134) );
  inv_x1_sg U43372 ( .A(reg_iii_12[0]), .X(n49628) );
  inv_x1_sg U43373 ( .A(reg_ii_12[0]), .X(n52132) );
  inv_x1_sg U43374 ( .A(reg_iii_12[1]), .X(n49626) );
  inv_x1_sg U43375 ( .A(reg_ii_12[1]), .X(n52130) );
  inv_x1_sg U43376 ( .A(reg_iii_12[2]), .X(n49624) );
  inv_x1_sg U43377 ( .A(reg_ii_12[2]), .X(n52128) );
  inv_x1_sg U43378 ( .A(reg_iii_12[3]), .X(n49622) );
  inv_x1_sg U43379 ( .A(reg_ii_12[3]), .X(n52126) );
  inv_x1_sg U43380 ( .A(reg_iii_12[4]), .X(n49620) );
  inv_x1_sg U43381 ( .A(reg_ii_12[4]), .X(n52124) );
  inv_x1_sg U43382 ( .A(reg_iii_12[5]), .X(n49618) );
  inv_x1_sg U43383 ( .A(reg_ii_12[5]), .X(n52122) );
  inv_x1_sg U43384 ( .A(reg_iii_12[6]), .X(n49616) );
  inv_x1_sg U43385 ( .A(reg_ii_12[6]), .X(n52120) );
  inv_x1_sg U43386 ( .A(reg_iii_12[7]), .X(n49614) );
  inv_x1_sg U43387 ( .A(reg_ii_12[7]), .X(n52118) );
  inv_x1_sg U43388 ( .A(reg_iii_12[8]), .X(n49612) );
  inv_x1_sg U43389 ( .A(reg_ii_12[8]), .X(n52116) );
  inv_x1_sg U43390 ( .A(reg_iii_12[9]), .X(n49610) );
  inv_x1_sg U43391 ( .A(reg_ii_12[9]), .X(n52114) );
  inv_x1_sg U43392 ( .A(reg_iii_12[10]), .X(n49608) );
  inv_x1_sg U43393 ( .A(reg_ii_12[10]), .X(n52112) );
  inv_x1_sg U43394 ( .A(reg_iii_12[11]), .X(n49606) );
  inv_x1_sg U43395 ( .A(reg_ii_12[11]), .X(n52110) );
  inv_x1_sg U43396 ( .A(reg_iii_12[12]), .X(n49604) );
  inv_x1_sg U43397 ( .A(reg_ii_12[12]), .X(n52108) );
  inv_x1_sg U43398 ( .A(reg_iii_12[13]), .X(n49602) );
  inv_x1_sg U43399 ( .A(reg_ii_12[13]), .X(n52106) );
  inv_x1_sg U43400 ( .A(reg_iii_12[14]), .X(n49600) );
  inv_x1_sg U43401 ( .A(reg_ii_12[14]), .X(n52104) );
  inv_x1_sg U43402 ( .A(reg_iii_12[15]), .X(n49598) );
  inv_x1_sg U43403 ( .A(reg_ii_12[15]), .X(n52102) );
  inv_x1_sg U43404 ( .A(reg_iii_12[16]), .X(n49596) );
  inv_x1_sg U43405 ( .A(reg_ii_12[16]), .X(n52100) );
  inv_x1_sg U43406 ( .A(reg_iii_12[17]), .X(n49594) );
  inv_x1_sg U43407 ( .A(reg_ii_12[17]), .X(n52098) );
  inv_x1_sg U43408 ( .A(reg_iii_12[18]), .X(n49592) );
  inv_x1_sg U43409 ( .A(reg_ii_12[18]), .X(n52096) );
  inv_x1_sg U43410 ( .A(reg_iii_12[19]), .X(n49590) );
  inv_x1_sg U43411 ( .A(reg_ii_12[19]), .X(n52094) );
  inv_x1_sg U43412 ( .A(reg_iii_13[0]), .X(n49588) );
  inv_x1_sg U43413 ( .A(reg_ii_13[0]), .X(n52092) );
  inv_x1_sg U43414 ( .A(reg_iii_13[1]), .X(n49586) );
  inv_x1_sg U43415 ( .A(reg_ii_13[1]), .X(n52090) );
  inv_x1_sg U43416 ( .A(reg_iii_13[2]), .X(n49584) );
  inv_x1_sg U43417 ( .A(reg_ii_13[2]), .X(n52088) );
  inv_x1_sg U43418 ( .A(reg_iii_13[3]), .X(n49582) );
  inv_x1_sg U43419 ( .A(reg_ii_13[3]), .X(n52086) );
  inv_x1_sg U43420 ( .A(reg_iii_13[4]), .X(n49580) );
  inv_x1_sg U43421 ( .A(reg_ii_13[4]), .X(n52084) );
  inv_x1_sg U43422 ( .A(reg_iii_13[5]), .X(n49578) );
  inv_x1_sg U43423 ( .A(reg_ii_13[5]), .X(n52082) );
  inv_x1_sg U43424 ( .A(reg_iii_13[6]), .X(n49576) );
  inv_x1_sg U43425 ( .A(reg_ii_13[6]), .X(n52080) );
  inv_x1_sg U43426 ( .A(reg_iii_13[7]), .X(n49574) );
  inv_x1_sg U43427 ( .A(reg_ii_13[7]), .X(n52078) );
  inv_x1_sg U43428 ( .A(reg_iii_13[8]), .X(n49572) );
  inv_x1_sg U43429 ( .A(reg_ii_13[8]), .X(n52076) );
  inv_x1_sg U43430 ( .A(reg_iii_13[9]), .X(n49570) );
  inv_x1_sg U43431 ( .A(reg_ii_13[9]), .X(n52074) );
  inv_x1_sg U43432 ( .A(reg_iii_13[10]), .X(n49568) );
  inv_x1_sg U43433 ( .A(reg_ii_13[10]), .X(n52072) );
  inv_x1_sg U43434 ( .A(reg_iii_13[11]), .X(n49566) );
  inv_x1_sg U43435 ( .A(reg_ii_13[11]), .X(n52070) );
  inv_x1_sg U43436 ( .A(reg_iii_13[12]), .X(n49564) );
  inv_x1_sg U43437 ( .A(reg_ii_13[12]), .X(n52068) );
  inv_x1_sg U43438 ( .A(reg_iii_13[13]), .X(n49562) );
  inv_x1_sg U43439 ( .A(reg_ii_13[13]), .X(n52066) );
  inv_x1_sg U43440 ( .A(reg_iii_13[14]), .X(n49560) );
  inv_x1_sg U43441 ( .A(reg_ii_13[14]), .X(n52064) );
  inv_x1_sg U43442 ( .A(reg_iii_13[15]), .X(n49558) );
  inv_x1_sg U43443 ( .A(reg_ii_13[15]), .X(n52062) );
  inv_x1_sg U43444 ( .A(reg_iii_13[16]), .X(n49556) );
  inv_x1_sg U43445 ( .A(reg_ii_13[16]), .X(n52060) );
  inv_x1_sg U43446 ( .A(reg_iii_13[17]), .X(n49554) );
  inv_x1_sg U43447 ( .A(reg_ii_13[17]), .X(n52058) );
  inv_x1_sg U43448 ( .A(reg_iii_13[18]), .X(n49552) );
  inv_x1_sg U43449 ( .A(reg_ii_13[18]), .X(n52056) );
  inv_x1_sg U43450 ( .A(reg_iii_13[19]), .X(n49550) );
  inv_x1_sg U43451 ( .A(reg_ii_13[19]), .X(n52054) );
  inv_x1_sg U43452 ( .A(reg_iii_14[0]), .X(n49548) );
  inv_x1_sg U43453 ( .A(reg_ii_14[0]), .X(n52052) );
  inv_x1_sg U43454 ( .A(reg_iii_14[1]), .X(n49546) );
  inv_x1_sg U43455 ( .A(reg_ii_14[1]), .X(n52050) );
  inv_x1_sg U43456 ( .A(reg_iii_14[2]), .X(n49544) );
  inv_x1_sg U43457 ( .A(reg_ii_14[2]), .X(n52048) );
  inv_x1_sg U43458 ( .A(reg_iii_14[3]), .X(n49542) );
  inv_x1_sg U43459 ( .A(reg_ii_14[3]), .X(n52046) );
  inv_x1_sg U43460 ( .A(reg_iii_14[4]), .X(n49540) );
  inv_x1_sg U43461 ( .A(reg_ii_14[4]), .X(n52044) );
  inv_x1_sg U43462 ( .A(reg_iii_14[5]), .X(n49538) );
  inv_x1_sg U43463 ( .A(reg_ii_14[5]), .X(n52042) );
  inv_x1_sg U43464 ( .A(reg_iii_14[6]), .X(n49536) );
  inv_x1_sg U43465 ( .A(reg_ii_14[6]), .X(n52040) );
  inv_x1_sg U43466 ( .A(reg_iii_14[7]), .X(n49534) );
  inv_x1_sg U43467 ( .A(reg_ii_14[7]), .X(n52038) );
  inv_x1_sg U43468 ( .A(reg_iii_14[8]), .X(n49532) );
  inv_x1_sg U43469 ( .A(reg_ii_14[8]), .X(n52036) );
  inv_x1_sg U43470 ( .A(reg_iii_14[9]), .X(n49530) );
  inv_x1_sg U43471 ( .A(reg_ii_14[9]), .X(n52034) );
  inv_x1_sg U43472 ( .A(reg_iii_14[10]), .X(n49528) );
  inv_x1_sg U43473 ( .A(reg_ii_14[10]), .X(n52032) );
  inv_x1_sg U43474 ( .A(reg_iii_14[11]), .X(n49526) );
  inv_x1_sg U43475 ( .A(reg_ii_14[11]), .X(n52030) );
  inv_x1_sg U43476 ( .A(reg_iii_14[12]), .X(n49524) );
  inv_x1_sg U43477 ( .A(reg_ii_14[12]), .X(n52028) );
  inv_x1_sg U43478 ( .A(reg_iii_14[13]), .X(n49522) );
  inv_x1_sg U43479 ( .A(reg_ii_14[13]), .X(n52026) );
  inv_x1_sg U43480 ( .A(reg_iii_14[14]), .X(n49520) );
  inv_x1_sg U43481 ( .A(reg_ii_14[14]), .X(n52024) );
  inv_x1_sg U43482 ( .A(reg_iii_14[15]), .X(n49518) );
  inv_x1_sg U43483 ( .A(reg_ii_14[15]), .X(n52022) );
  inv_x1_sg U43484 ( .A(reg_iii_14[16]), .X(n49516) );
  inv_x1_sg U43485 ( .A(reg_ii_14[16]), .X(n52020) );
  inv_x1_sg U43486 ( .A(reg_iii_4[19]), .X(n49514) );
  inv_x1_sg U43487 ( .A(reg_ii_4[19]), .X(n52018) );
  inv_x1_sg U43488 ( .A(reg_iii_5[0]), .X(n49512) );
  inv_x1_sg U43489 ( .A(reg_ii_5[0]), .X(n52016) );
  inv_x1_sg U43490 ( .A(reg_iii_5[1]), .X(n49510) );
  inv_x1_sg U43491 ( .A(reg_ii_5[1]), .X(n52014) );
  inv_x1_sg U43492 ( .A(reg_iii_5[2]), .X(n49508) );
  inv_x1_sg U43493 ( .A(reg_ii_5[2]), .X(n52012) );
  inv_x1_sg U43494 ( .A(reg_iii_5[3]), .X(n49506) );
  inv_x1_sg U43495 ( .A(reg_ii_5[3]), .X(n52010) );
  inv_x1_sg U43496 ( .A(reg_iii_5[4]), .X(n49504) );
  inv_x1_sg U43497 ( .A(reg_ii_5[4]), .X(n52008) );
  inv_x1_sg U43498 ( .A(reg_iii_5[5]), .X(n49502) );
  inv_x1_sg U43499 ( .A(reg_ii_5[5]), .X(n52006) );
  inv_x1_sg U43500 ( .A(reg_iii_5[6]), .X(n49500) );
  inv_x1_sg U43501 ( .A(reg_ii_5[6]), .X(n52004) );
  inv_x1_sg U43502 ( .A(reg_iii_5[7]), .X(n49498) );
  inv_x1_sg U43503 ( .A(reg_ii_5[7]), .X(n52002) );
  inv_x1_sg U43504 ( .A(reg_iii_5[8]), .X(n49496) );
  inv_x1_sg U43505 ( .A(reg_ii_5[8]), .X(n52000) );
  inv_x1_sg U43506 ( .A(reg_iii_5[9]), .X(n49494) );
  inv_x1_sg U43507 ( .A(reg_ii_5[9]), .X(n51998) );
  inv_x1_sg U43508 ( .A(reg_iii_5[10]), .X(n49492) );
  inv_x1_sg U43509 ( .A(reg_ii_5[10]), .X(n51996) );
  inv_x1_sg U43510 ( .A(reg_iii_5[11]), .X(n49490) );
  inv_x1_sg U43511 ( .A(reg_ii_5[11]), .X(n51994) );
  inv_x1_sg U43512 ( .A(reg_iii_5[12]), .X(n49488) );
  inv_x1_sg U43513 ( .A(reg_ii_5[12]), .X(n51992) );
  inv_x1_sg U43514 ( .A(reg_iii_5[13]), .X(n49486) );
  inv_x1_sg U43515 ( .A(reg_ii_5[13]), .X(n51990) );
  inv_x1_sg U43516 ( .A(reg_iii_5[14]), .X(n49484) );
  inv_x1_sg U43517 ( .A(reg_ii_5[14]), .X(n51988) );
  inv_x1_sg U43518 ( .A(reg_iii_5[15]), .X(n49482) );
  inv_x1_sg U43519 ( .A(reg_ii_5[15]), .X(n51986) );
  inv_x1_sg U43520 ( .A(reg_iii_5[16]), .X(n49480) );
  inv_x1_sg U43521 ( .A(reg_ii_5[16]), .X(n51984) );
  inv_x1_sg U43522 ( .A(reg_iii_5[17]), .X(n49478) );
  inv_x1_sg U43523 ( .A(reg_ii_5[17]), .X(n51982) );
  inv_x1_sg U43524 ( .A(reg_iii_5[18]), .X(n49476) );
  inv_x1_sg U43525 ( .A(reg_ii_5[18]), .X(n51980) );
  inv_x1_sg U43526 ( .A(reg_iii_5[19]), .X(n49474) );
  inv_x1_sg U43527 ( .A(reg_ii_5[19]), .X(n51978) );
  inv_x1_sg U43528 ( .A(reg_iii_6[0]), .X(n49472) );
  inv_x1_sg U43529 ( .A(reg_ii_6[0]), .X(n51976) );
  inv_x1_sg U43530 ( .A(reg_iii_6[1]), .X(n49470) );
  inv_x1_sg U43531 ( .A(reg_ii_6[1]), .X(n51974) );
  inv_x1_sg U43532 ( .A(reg_iii_6[2]), .X(n49468) );
  inv_x1_sg U43533 ( .A(reg_ii_6[2]), .X(n51972) );
  inv_x1_sg U43534 ( .A(reg_iii_6[3]), .X(n49466) );
  inv_x1_sg U43535 ( .A(reg_ii_6[3]), .X(n51970) );
  inv_x1_sg U43536 ( .A(reg_iii_6[4]), .X(n49464) );
  inv_x1_sg U43537 ( .A(reg_ii_6[4]), .X(n51968) );
  inv_x1_sg U43538 ( .A(reg_iii_6[5]), .X(n49462) );
  inv_x1_sg U43539 ( .A(reg_ii_6[5]), .X(n51966) );
  inv_x1_sg U43540 ( .A(reg_iii_6[6]), .X(n49460) );
  inv_x1_sg U43541 ( .A(reg_ii_6[6]), .X(n51964) );
  inv_x1_sg U43542 ( .A(reg_iii_6[7]), .X(n49458) );
  inv_x1_sg U43543 ( .A(reg_ii_6[7]), .X(n51962) );
  inv_x1_sg U43544 ( .A(reg_iii_6[8]), .X(n49456) );
  inv_x1_sg U43545 ( .A(reg_ii_6[8]), .X(n51960) );
  inv_x1_sg U43546 ( .A(reg_iii_6[9]), .X(n49454) );
  inv_x1_sg U43547 ( .A(reg_ii_6[9]), .X(n51958) );
  inv_x1_sg U43548 ( .A(reg_iii_6[10]), .X(n49452) );
  inv_x1_sg U43549 ( .A(reg_ii_6[10]), .X(n51956) );
  inv_x1_sg U43550 ( .A(reg_iii_6[11]), .X(n49450) );
  inv_x1_sg U43551 ( .A(reg_ii_6[11]), .X(n51954) );
  inv_x1_sg U43552 ( .A(reg_iii_6[12]), .X(n49448) );
  inv_x1_sg U43553 ( .A(reg_ii_6[12]), .X(n51952) );
  inv_x1_sg U43554 ( .A(reg_iii_6[13]), .X(n49446) );
  inv_x1_sg U43555 ( .A(reg_ii_6[13]), .X(n51950) );
  inv_x1_sg U43556 ( .A(reg_iii_6[14]), .X(n49444) );
  inv_x1_sg U43557 ( .A(reg_ii_6[14]), .X(n51948) );
  inv_x1_sg U43558 ( .A(reg_iii_6[15]), .X(n49442) );
  inv_x1_sg U43559 ( .A(reg_ii_6[15]), .X(n51946) );
  inv_x1_sg U43560 ( .A(reg_iii_6[16]), .X(n49440) );
  inv_x1_sg U43561 ( .A(reg_ii_6[16]), .X(n51944) );
  inv_x1_sg U43562 ( .A(reg_iii_6[17]), .X(n49438) );
  inv_x1_sg U43563 ( .A(reg_ii_6[17]), .X(n51942) );
  inv_x1_sg U43564 ( .A(reg_iii_6[18]), .X(n49436) );
  inv_x1_sg U43565 ( .A(reg_ii_6[18]), .X(n51940) );
  inv_x1_sg U43566 ( .A(reg_iii_6[19]), .X(n49434) );
  inv_x1_sg U43567 ( .A(reg_ii_6[19]), .X(n51938) );
  inv_x1_sg U43568 ( .A(reg_iii_7[0]), .X(n49432) );
  inv_x1_sg U43569 ( .A(reg_ii_7[0]), .X(n51936) );
  inv_x1_sg U43570 ( .A(reg_iii_7[1]), .X(n49430) );
  inv_x1_sg U43571 ( .A(reg_ii_7[1]), .X(n51934) );
  inv_x1_sg U43572 ( .A(reg_iii_7[2]), .X(n49428) );
  inv_x1_sg U43573 ( .A(reg_ii_7[2]), .X(n51932) );
  inv_x1_sg U43574 ( .A(reg_iii_7[3]), .X(n49426) );
  inv_x1_sg U43575 ( .A(reg_ii_7[3]), .X(n51930) );
  inv_x1_sg U43576 ( .A(reg_iii_7[4]), .X(n49424) );
  inv_x1_sg U43577 ( .A(reg_ii_7[4]), .X(n51928) );
  inv_x1_sg U43578 ( .A(reg_iii_7[5]), .X(n49422) );
  inv_x1_sg U43579 ( .A(reg_ii_7[5]), .X(n51926) );
  inv_x1_sg U43580 ( .A(reg_iii_7[6]), .X(n49420) );
  inv_x1_sg U43581 ( .A(reg_ii_7[6]), .X(n51924) );
  inv_x1_sg U43582 ( .A(reg_iii_7[7]), .X(n49418) );
  inv_x1_sg U43583 ( .A(reg_ii_7[7]), .X(n51922) );
  inv_x1_sg U43584 ( .A(reg_iii_7[8]), .X(n49416) );
  inv_x1_sg U43585 ( .A(reg_ii_7[8]), .X(n51920) );
  inv_x1_sg U43586 ( .A(reg_iii_7[9]), .X(n49414) );
  inv_x1_sg U43587 ( .A(reg_ii_7[9]), .X(n51918) );
  inv_x1_sg U43588 ( .A(reg_iii_7[10]), .X(n49412) );
  inv_x1_sg U43589 ( .A(reg_ii_7[10]), .X(n51916) );
  inv_x1_sg U43590 ( .A(reg_iii_7[11]), .X(n49410) );
  inv_x1_sg U43591 ( .A(reg_ii_7[11]), .X(n51914) );
  inv_x1_sg U43592 ( .A(reg_iii_7[12]), .X(n49408) );
  inv_x1_sg U43593 ( .A(reg_ii_7[12]), .X(n51912) );
  inv_x1_sg U43594 ( .A(reg_iii_7[13]), .X(n49406) );
  inv_x1_sg U43595 ( .A(reg_ii_7[13]), .X(n51910) );
  inv_x1_sg U43596 ( .A(reg_iii_7[14]), .X(n49404) );
  inv_x1_sg U43597 ( .A(reg_ii_7[14]), .X(n51908) );
  inv_x1_sg U43598 ( .A(reg_iii_7[15]), .X(n49402) );
  inv_x1_sg U43599 ( .A(reg_ii_7[15]), .X(n51906) );
  inv_x1_sg U43600 ( .A(reg_iii_7[16]), .X(n49400) );
  inv_x1_sg U43601 ( .A(reg_ii_7[16]), .X(n51904) );
  inv_x1_sg U43602 ( .A(reg_iii_7[17]), .X(n49398) );
  inv_x1_sg U43603 ( .A(reg_ii_7[17]), .X(n51902) );
  inv_x1_sg U43604 ( .A(reg_iii_7[18]), .X(n49396) );
  inv_x1_sg U43605 ( .A(reg_ii_7[18]), .X(n51900) );
  inv_x1_sg U43606 ( .A(reg_iii_7[19]), .X(n49394) );
  inv_x1_sg U43607 ( .A(reg_ii_7[19]), .X(n51898) );
  inv_x1_sg U43608 ( .A(reg_iii_8[0]), .X(n49392) );
  inv_x1_sg U43609 ( .A(reg_ii_8[0]), .X(n51896) );
  inv_x1_sg U43610 ( .A(reg_iii_8[1]), .X(n49390) );
  inv_x1_sg U43611 ( .A(reg_ii_8[1]), .X(n51894) );
  inv_x1_sg U43612 ( .A(reg_iii_8[2]), .X(n49388) );
  inv_x1_sg U43613 ( .A(reg_ii_8[2]), .X(n51892) );
  inv_x1_sg U43614 ( .A(reg_iii_8[3]), .X(n49386) );
  inv_x1_sg U43615 ( .A(reg_ii_8[3]), .X(n51890) );
  inv_x1_sg U43616 ( .A(reg_iii_8[4]), .X(n49384) );
  inv_x1_sg U43617 ( .A(reg_ii_8[4]), .X(n51888) );
  inv_x1_sg U43618 ( .A(reg_iii_8[5]), .X(n49382) );
  inv_x1_sg U43619 ( .A(reg_ii_8[5]), .X(n51886) );
  inv_x1_sg U43620 ( .A(reg_iii_8[6]), .X(n49380) );
  inv_x1_sg U43621 ( .A(reg_ii_8[6]), .X(n51884) );
  inv_x1_sg U43622 ( .A(reg_iii_8[7]), .X(n49378) );
  inv_x1_sg U43623 ( .A(reg_ii_8[7]), .X(n51882) );
  inv_x1_sg U43624 ( .A(reg_iii_8[8]), .X(n49376) );
  inv_x1_sg U43625 ( .A(reg_ii_8[8]), .X(n51880) );
  inv_x1_sg U43626 ( .A(reg_iii_8[9]), .X(n49374) );
  inv_x1_sg U43627 ( .A(reg_ii_8[9]), .X(n51878) );
  inv_x1_sg U43628 ( .A(reg_iii_8[10]), .X(n49372) );
  inv_x1_sg U43629 ( .A(reg_ii_8[10]), .X(n51876) );
  inv_x1_sg U43630 ( .A(reg_iii_8[11]), .X(n49370) );
  inv_x1_sg U43631 ( .A(reg_ii_8[11]), .X(n51874) );
  inv_x1_sg U43632 ( .A(reg_iii_8[12]), .X(n49368) );
  inv_x1_sg U43633 ( .A(reg_ii_8[12]), .X(n51872) );
  inv_x1_sg U43634 ( .A(reg_iii_8[13]), .X(n49366) );
  inv_x1_sg U43635 ( .A(reg_ii_8[13]), .X(n51870) );
  inv_x1_sg U43636 ( .A(reg_iii_8[14]), .X(n49364) );
  inv_x1_sg U43637 ( .A(reg_ii_8[14]), .X(n51868) );
  inv_x1_sg U43638 ( .A(reg_iii_8[15]), .X(n49362) );
  inv_x1_sg U43639 ( .A(reg_ii_8[15]), .X(n51866) );
  inv_x1_sg U43640 ( .A(reg_iii_8[16]), .X(n49360) );
  inv_x1_sg U43641 ( .A(reg_ii_8[16]), .X(n51864) );
  inv_x1_sg U43642 ( .A(reg_iii_8[17]), .X(n49358) );
  inv_x1_sg U43643 ( .A(reg_ii_8[17]), .X(n51862) );
  inv_x1_sg U43644 ( .A(reg_iii_8[18]), .X(n49356) );
  inv_x1_sg U43645 ( .A(reg_ii_8[18]), .X(n51860) );
  inv_x1_sg U43646 ( .A(reg_iii_8[19]), .X(n49354) );
  inv_x1_sg U43647 ( .A(reg_ii_8[19]), .X(n51858) );
  inv_x1_sg U43648 ( .A(reg_iii_9[0]), .X(n49352) );
  inv_x1_sg U43649 ( .A(reg_ii_9[0]), .X(n51856) );
  inv_x1_sg U43650 ( .A(reg_iii_9[1]), .X(n49350) );
  inv_x1_sg U43651 ( .A(reg_ii_9[1]), .X(n51854) );
  inv_x1_sg U43652 ( .A(reg_iii_9[2]), .X(n49348) );
  inv_x1_sg U43653 ( .A(reg_ii_9[2]), .X(n51852) );
  inv_x1_sg U43654 ( .A(reg_iii_9[3]), .X(n49346) );
  inv_x1_sg U43655 ( .A(reg_ii_9[3]), .X(n51850) );
  inv_x1_sg U43656 ( .A(reg_iii_9[4]), .X(n49344) );
  inv_x1_sg U43657 ( .A(reg_ii_9[4]), .X(n51848) );
  inv_x1_sg U43658 ( .A(reg_iii_9[5]), .X(n49342) );
  inv_x1_sg U43659 ( .A(reg_ii_9[5]), .X(n51846) );
  inv_x1_sg U43660 ( .A(reg_iii_9[6]), .X(n49340) );
  inv_x1_sg U43661 ( .A(reg_ii_9[6]), .X(n51844) );
  inv_x1_sg U43662 ( .A(reg_iii_9[7]), .X(n49338) );
  inv_x1_sg U43663 ( .A(reg_ii_9[7]), .X(n51842) );
  inv_x1_sg U43664 ( .A(reg_iii_9[8]), .X(n49336) );
  inv_x1_sg U43665 ( .A(reg_ii_9[8]), .X(n51840) );
  inv_x1_sg U43666 ( .A(reg_iii_9[9]), .X(n49334) );
  inv_x1_sg U43667 ( .A(reg_ii_9[9]), .X(n51838) );
  inv_x1_sg U43668 ( .A(reg_iii_9[10]), .X(n49332) );
  inv_x1_sg U43669 ( .A(reg_ii_9[10]), .X(n51836) );
  inv_x1_sg U43670 ( .A(reg_iii_9[11]), .X(n49330) );
  inv_x1_sg U43671 ( .A(reg_ii_9[11]), .X(n51834) );
  inv_x1_sg U43672 ( .A(reg_iii_9[12]), .X(n49328) );
  inv_x1_sg U43673 ( .A(reg_ii_9[12]), .X(n51832) );
  inv_x1_sg U43674 ( .A(reg_iii_9[13]), .X(n49326) );
  inv_x1_sg U43675 ( .A(reg_ii_9[13]), .X(n51830) );
  inv_x1_sg U43676 ( .A(reg_iii_9[14]), .X(n49324) );
  inv_x1_sg U43677 ( .A(reg_ii_9[14]), .X(n51828) );
  inv_x1_sg U43678 ( .A(reg_iii_9[15]), .X(n49322) );
  inv_x1_sg U43679 ( .A(reg_ii_9[15]), .X(n51826) );
  inv_x1_sg U43680 ( .A(reg_iii_9[16]), .X(n49320) );
  inv_x1_sg U43681 ( .A(reg_ii_9[16]), .X(n51824) );
  inv_x1_sg U43682 ( .A(reg_iii_9[17]), .X(n49318) );
  inv_x1_sg U43683 ( .A(reg_ii_9[17]), .X(n51822) );
  inv_x1_sg U43684 ( .A(reg_iii_0[0]), .X(n49316) );
  inv_x1_sg U43685 ( .A(reg_ii_0[0]), .X(n51820) );
  inv_x1_sg U43686 ( .A(reg_iii_0[1]), .X(n49314) );
  inv_x1_sg U43687 ( .A(reg_ii_0[1]), .X(n51818) );
  inv_x1_sg U43688 ( .A(reg_iii_0[2]), .X(n49312) );
  inv_x1_sg U43689 ( .A(reg_ii_0[2]), .X(n51816) );
  inv_x1_sg U43690 ( .A(reg_iii_0[3]), .X(n49310) );
  inv_x1_sg U43691 ( .A(reg_ii_0[3]), .X(n51814) );
  inv_x1_sg U43692 ( .A(reg_iii_0[4]), .X(n49308) );
  inv_x1_sg U43693 ( .A(reg_ii_0[4]), .X(n51812) );
  inv_x1_sg U43694 ( .A(reg_iii_0[5]), .X(n49306) );
  inv_x1_sg U43695 ( .A(reg_ii_0[5]), .X(n51810) );
  inv_x1_sg U43696 ( .A(reg_iii_0[6]), .X(n49304) );
  inv_x1_sg U43697 ( .A(reg_ii_0[6]), .X(n51808) );
  inv_x1_sg U43698 ( .A(reg_iii_0[7]), .X(n49302) );
  inv_x1_sg U43699 ( .A(reg_ii_0[7]), .X(n51806) );
  inv_x1_sg U43700 ( .A(reg_iii_0[8]), .X(n49300) );
  inv_x1_sg U43701 ( .A(reg_ii_0[8]), .X(n51804) );
  inv_x1_sg U43702 ( .A(reg_iii_0[9]), .X(n49298) );
  inv_x1_sg U43703 ( .A(reg_ii_0[9]), .X(n51802) );
  inv_x1_sg U43704 ( .A(reg_iii_0[10]), .X(n49296) );
  inv_x1_sg U43705 ( .A(reg_ii_0[10]), .X(n51800) );
  inv_x1_sg U43706 ( .A(reg_iii_0[11]), .X(n49294) );
  inv_x1_sg U43707 ( .A(reg_ii_0[11]), .X(n51798) );
  inv_x1_sg U43708 ( .A(reg_iii_0[12]), .X(n49292) );
  inv_x1_sg U43709 ( .A(reg_ii_0[12]), .X(n51796) );
  inv_x1_sg U43710 ( .A(reg_iii_0[13]), .X(n49290) );
  inv_x1_sg U43711 ( .A(reg_ii_0[13]), .X(n51794) );
  inv_x1_sg U43712 ( .A(reg_iii_0[14]), .X(n49288) );
  inv_x1_sg U43713 ( .A(reg_ii_0[14]), .X(n51792) );
  inv_x1_sg U43714 ( .A(reg_iii_0[15]), .X(n49286) );
  inv_x1_sg U43715 ( .A(reg_ii_0[15]), .X(n51790) );
  inv_x1_sg U43716 ( .A(reg_iii_0[16]), .X(n49284) );
  inv_x1_sg U43717 ( .A(reg_ii_0[16]), .X(n51788) );
  inv_x1_sg U43718 ( .A(reg_iii_0[17]), .X(n49282) );
  inv_x1_sg U43719 ( .A(reg_ii_0[17]), .X(n51786) );
  inv_x1_sg U43720 ( .A(reg_iii_0[18]), .X(n49280) );
  inv_x1_sg U43721 ( .A(reg_ii_0[18]), .X(n51784) );
  inv_x1_sg U43722 ( .A(reg_iii_0[19]), .X(n49278) );
  inv_x1_sg U43723 ( .A(reg_ii_0[19]), .X(n51782) );
  inv_x1_sg U43724 ( .A(reg_iii_1[0]), .X(n49276) );
  inv_x1_sg U43725 ( .A(reg_ii_1[0]), .X(n51780) );
  inv_x1_sg U43726 ( .A(reg_iii_1[1]), .X(n49274) );
  inv_x1_sg U43727 ( .A(reg_ii_1[1]), .X(n51778) );
  inv_x1_sg U43728 ( .A(reg_iii_1[2]), .X(n49272) );
  inv_x1_sg U43729 ( .A(reg_ii_1[2]), .X(n51776) );
  inv_x1_sg U43730 ( .A(reg_iii_1[3]), .X(n49270) );
  inv_x1_sg U43731 ( .A(reg_ii_1[3]), .X(n51774) );
  inv_x1_sg U43732 ( .A(reg_iii_1[4]), .X(n49268) );
  inv_x1_sg U43733 ( .A(reg_ii_1[4]), .X(n51772) );
  inv_x1_sg U43734 ( .A(reg_iii_1[5]), .X(n49266) );
  inv_x1_sg U43735 ( .A(reg_ii_1[5]), .X(n51770) );
  inv_x1_sg U43736 ( .A(reg_iii_1[6]), .X(n49264) );
  inv_x1_sg U43737 ( .A(reg_ii_1[6]), .X(n51768) );
  inv_x1_sg U43738 ( .A(reg_iii_1[7]), .X(n49262) );
  inv_x1_sg U43739 ( .A(reg_ii_1[7]), .X(n51766) );
  inv_x1_sg U43740 ( .A(reg_iii_1[8]), .X(n49260) );
  inv_x1_sg U43741 ( .A(reg_ii_1[8]), .X(n51764) );
  inv_x1_sg U43742 ( .A(reg_iii_1[9]), .X(n49258) );
  inv_x1_sg U43743 ( .A(reg_ii_1[9]), .X(n51762) );
  inv_x1_sg U43744 ( .A(reg_iii_1[10]), .X(n49256) );
  inv_x1_sg U43745 ( .A(reg_ii_1[10]), .X(n51760) );
  inv_x1_sg U43746 ( .A(reg_iii_1[11]), .X(n49254) );
  inv_x1_sg U43747 ( .A(reg_ii_1[11]), .X(n51758) );
  inv_x1_sg U43748 ( .A(reg_iii_1[12]), .X(n49252) );
  inv_x1_sg U43749 ( .A(reg_ii_1[12]), .X(n51756) );
  inv_x1_sg U43750 ( .A(reg_iii_1[13]), .X(n49250) );
  inv_x1_sg U43751 ( .A(reg_ii_1[13]), .X(n51754) );
  inv_x1_sg U43752 ( .A(reg_iii_1[14]), .X(n49248) );
  inv_x1_sg U43753 ( .A(reg_ii_1[14]), .X(n51752) );
  inv_x1_sg U43754 ( .A(reg_iii_1[15]), .X(n49246) );
  inv_x1_sg U43755 ( .A(reg_ii_1[15]), .X(n51750) );
  inv_x1_sg U43756 ( .A(reg_iii_1[16]), .X(n49244) );
  inv_x1_sg U43757 ( .A(reg_ii_1[16]), .X(n51748) );
  inv_x1_sg U43758 ( .A(reg_iii_1[17]), .X(n49242) );
  inv_x1_sg U43759 ( .A(reg_ii_1[17]), .X(n51746) );
  inv_x1_sg U43760 ( .A(reg_iii_1[18]), .X(n49240) );
  inv_x1_sg U43761 ( .A(reg_ii_1[18]), .X(n51744) );
  inv_x1_sg U43762 ( .A(reg_iii_1[19]), .X(n49238) );
  inv_x1_sg U43763 ( .A(reg_ii_1[19]), .X(n51742) );
  inv_x1_sg U43764 ( .A(reg_iii_2[0]), .X(n49236) );
  inv_x1_sg U43765 ( .A(reg_ii_2[0]), .X(n51740) );
  inv_x1_sg U43766 ( .A(reg_iii_2[1]), .X(n49234) );
  inv_x1_sg U43767 ( .A(reg_ii_2[1]), .X(n51738) );
  inv_x1_sg U43768 ( .A(reg_iii_2[2]), .X(n49232) );
  inv_x1_sg U43769 ( .A(reg_ii_2[2]), .X(n51736) );
  inv_x1_sg U43770 ( .A(reg_iii_2[3]), .X(n49230) );
  inv_x1_sg U43771 ( .A(reg_ii_2[3]), .X(n51734) );
  inv_x1_sg U43772 ( .A(reg_iii_2[4]), .X(n49228) );
  inv_x1_sg U43773 ( .A(reg_ii_2[4]), .X(n51732) );
  inv_x1_sg U43774 ( .A(reg_iii_2[5]), .X(n49226) );
  inv_x1_sg U43775 ( .A(reg_ii_2[5]), .X(n51730) );
  inv_x1_sg U43776 ( .A(reg_iii_2[6]), .X(n49224) );
  inv_x1_sg U43777 ( .A(reg_ii_2[6]), .X(n51728) );
  inv_x1_sg U43778 ( .A(reg_iii_2[7]), .X(n49222) );
  inv_x1_sg U43779 ( .A(reg_ii_2[7]), .X(n51726) );
  inv_x1_sg U43780 ( .A(reg_iii_2[8]), .X(n49220) );
  inv_x1_sg U43781 ( .A(reg_ii_2[8]), .X(n51724) );
  inv_x1_sg U43782 ( .A(reg_iii_2[9]), .X(n49218) );
  inv_x1_sg U43783 ( .A(reg_ii_2[9]), .X(n51722) );
  inv_x1_sg U43784 ( .A(reg_iii_2[10]), .X(n49216) );
  inv_x1_sg U43785 ( .A(reg_ii_2[10]), .X(n51720) );
  inv_x1_sg U43786 ( .A(reg_iii_2[11]), .X(n49214) );
  inv_x1_sg U43787 ( .A(reg_ii_2[11]), .X(n51718) );
  inv_x1_sg U43788 ( .A(reg_iii_2[12]), .X(n49212) );
  inv_x1_sg U43789 ( .A(reg_ii_2[12]), .X(n51716) );
  inv_x1_sg U43790 ( .A(reg_iii_2[13]), .X(n49210) );
  inv_x1_sg U43791 ( .A(reg_ii_2[13]), .X(n51714) );
  inv_x1_sg U43792 ( .A(reg_iii_2[14]), .X(n49208) );
  inv_x1_sg U43793 ( .A(reg_ii_2[14]), .X(n51712) );
  inv_x1_sg U43794 ( .A(reg_iii_2[15]), .X(n49206) );
  inv_x1_sg U43795 ( .A(reg_ii_2[15]), .X(n51710) );
  inv_x1_sg U43796 ( .A(reg_iii_2[16]), .X(n49204) );
  inv_x1_sg U43797 ( .A(reg_ii_2[16]), .X(n51708) );
  inv_x1_sg U43798 ( .A(reg_iii_2[17]), .X(n49202) );
  inv_x1_sg U43799 ( .A(reg_ii_2[17]), .X(n51706) );
  inv_x1_sg U43800 ( .A(reg_iii_2[18]), .X(n49200) );
  inv_x1_sg U43801 ( .A(reg_ii_2[18]), .X(n51704) );
  inv_x1_sg U43802 ( .A(reg_iii_2[19]), .X(n49198) );
  inv_x1_sg U43803 ( .A(reg_ii_2[19]), .X(n51702) );
  inv_x1_sg U43804 ( .A(reg_iii_3[0]), .X(n49196) );
  inv_x1_sg U43805 ( .A(reg_ii_3[0]), .X(n51700) );
  inv_x1_sg U43806 ( .A(reg_iii_3[1]), .X(n49194) );
  inv_x1_sg U43807 ( .A(reg_ii_3[1]), .X(n51698) );
  inv_x1_sg U43808 ( .A(reg_iii_3[2]), .X(n49192) );
  inv_x1_sg U43809 ( .A(reg_ii_3[2]), .X(n51696) );
  inv_x1_sg U43810 ( .A(reg_iii_3[3]), .X(n49190) );
  inv_x1_sg U43811 ( .A(reg_ii_3[3]), .X(n51694) );
  inv_x1_sg U43812 ( .A(reg_iii_3[4]), .X(n49188) );
  inv_x1_sg U43813 ( .A(reg_ii_3[4]), .X(n51692) );
  inv_x1_sg U43814 ( .A(reg_iii_3[5]), .X(n49186) );
  inv_x1_sg U43815 ( .A(reg_ii_3[5]), .X(n51690) );
  inv_x1_sg U43816 ( .A(reg_iii_3[6]), .X(n49184) );
  inv_x1_sg U43817 ( .A(reg_ii_3[6]), .X(n51688) );
  inv_x1_sg U43818 ( .A(reg_iii_3[7]), .X(n49182) );
  inv_x1_sg U43819 ( .A(reg_ii_3[7]), .X(n51686) );
  inv_x1_sg U43820 ( .A(reg_iii_3[8]), .X(n49180) );
  inv_x1_sg U43821 ( .A(reg_ii_3[8]), .X(n51684) );
  inv_x1_sg U43822 ( .A(reg_iii_3[9]), .X(n49178) );
  inv_x1_sg U43823 ( .A(reg_ii_3[9]), .X(n51682) );
  inv_x1_sg U43824 ( .A(reg_iii_3[10]), .X(n49176) );
  inv_x1_sg U43825 ( .A(reg_ii_3[10]), .X(n51680) );
  inv_x1_sg U43826 ( .A(reg_iii_3[11]), .X(n49174) );
  inv_x1_sg U43827 ( .A(reg_ii_3[11]), .X(n51678) );
  inv_x1_sg U43828 ( .A(reg_iii_3[12]), .X(n49172) );
  inv_x1_sg U43829 ( .A(reg_ii_3[12]), .X(n51676) );
  inv_x1_sg U43830 ( .A(reg_iii_3[13]), .X(n49170) );
  inv_x1_sg U43831 ( .A(reg_ii_3[13]), .X(n51674) );
  inv_x1_sg U43832 ( .A(reg_iii_3[14]), .X(n49168) );
  inv_x1_sg U43833 ( .A(reg_ii_3[14]), .X(n51672) );
  inv_x1_sg U43834 ( .A(reg_iii_3[15]), .X(n49166) );
  inv_x1_sg U43835 ( .A(reg_ii_3[15]), .X(n51670) );
  inv_x1_sg U43836 ( .A(reg_iii_3[16]), .X(n49164) );
  inv_x1_sg U43837 ( .A(reg_ii_3[16]), .X(n51668) );
  inv_x1_sg U43838 ( .A(reg_iii_3[17]), .X(n49162) );
  inv_x1_sg U43839 ( .A(reg_ii_3[17]), .X(n51666) );
  inv_x1_sg U43840 ( .A(reg_iii_3[18]), .X(n49160) );
  inv_x1_sg U43841 ( .A(reg_ii_3[18]), .X(n51664) );
  inv_x1_sg U43842 ( .A(reg_iii_3[19]), .X(n49158) );
  inv_x1_sg U43843 ( .A(reg_ii_3[19]), .X(n51662) );
  inv_x1_sg U43844 ( .A(reg_iii_4[0]), .X(n49156) );
  inv_x1_sg U43845 ( .A(reg_ii_4[0]), .X(n51660) );
  inv_x1_sg U43846 ( .A(reg_iii_4[1]), .X(n49154) );
  inv_x1_sg U43847 ( .A(reg_ii_4[1]), .X(n51658) );
  inv_x1_sg U43848 ( .A(reg_iii_4[2]), .X(n49152) );
  inv_x1_sg U43849 ( .A(reg_ii_4[2]), .X(n51656) );
  inv_x1_sg U43850 ( .A(reg_iii_4[3]), .X(n49150) );
  inv_x1_sg U43851 ( .A(reg_ii_4[3]), .X(n51654) );
  inv_x1_sg U43852 ( .A(reg_iii_4[4]), .X(n49148) );
  inv_x1_sg U43853 ( .A(reg_ii_4[4]), .X(n51652) );
  inv_x1_sg U43854 ( .A(reg_iii_4[5]), .X(n49146) );
  inv_x1_sg U43855 ( .A(reg_ii_4[5]), .X(n51650) );
  inv_x1_sg U43856 ( .A(reg_iii_4[6]), .X(n49144) );
  inv_x1_sg U43857 ( .A(reg_ii_4[6]), .X(n51648) );
  inv_x1_sg U43858 ( .A(reg_iii_4[7]), .X(n49142) );
  inv_x1_sg U43859 ( .A(reg_ii_4[7]), .X(n51646) );
  inv_x1_sg U43860 ( .A(reg_iii_4[8]), .X(n49140) );
  inv_x1_sg U43861 ( .A(reg_ii_4[8]), .X(n51644) );
  inv_x1_sg U43862 ( .A(reg_iii_4[9]), .X(n49138) );
  inv_x1_sg U43863 ( .A(reg_ii_4[9]), .X(n51642) );
  inv_x1_sg U43864 ( .A(reg_iii_4[10]), .X(n49136) );
  inv_x1_sg U43865 ( .A(reg_ii_4[10]), .X(n51640) );
  inv_x1_sg U43866 ( .A(reg_iii_4[11]), .X(n49134) );
  inv_x1_sg U43867 ( .A(reg_ii_4[11]), .X(n51638) );
  inv_x1_sg U43868 ( .A(reg_iii_4[12]), .X(n49132) );
  inv_x1_sg U43869 ( .A(reg_ii_4[12]), .X(n51636) );
  inv_x1_sg U43870 ( .A(reg_iii_4[13]), .X(n49130) );
  inv_x1_sg U43871 ( .A(reg_ii_4[13]), .X(n51634) );
  inv_x1_sg U43872 ( .A(reg_iii_4[14]), .X(n49128) );
  inv_x1_sg U43873 ( .A(reg_ii_4[14]), .X(n51632) );
  inv_x1_sg U43874 ( .A(reg_iii_4[15]), .X(n49126) );
  inv_x1_sg U43875 ( .A(reg_ii_4[15]), .X(n51630) );
  inv_x1_sg U43876 ( .A(reg_iii_4[16]), .X(n49124) );
  inv_x1_sg U43877 ( .A(reg_ii_4[16]), .X(n51628) );
  inv_x1_sg U43878 ( .A(reg_iii_4[17]), .X(n49122) );
  inv_x1_sg U43879 ( .A(reg_ii_4[17]), .X(n51626) );
  inv_x1_sg U43880 ( .A(reg_iii_4[18]), .X(n49120) );
  inv_x1_sg U43881 ( .A(reg_ii_4[18]), .X(n51624) );
  inv_x1_sg U43882 ( .A(reg_w_15[19]), .X(n49118) );
  inv_x1_sg U43883 ( .A(reg_w_15[18]), .X(n49116) );
  inv_x1_sg U43884 ( .A(reg_w_15[17]), .X(n49114) );
  inv_x1_sg U43885 ( .A(reg_w_15[16]), .X(n49112) );
  inv_x1_sg U43886 ( .A(reg_w_15[15]), .X(n49110) );
  inv_x1_sg U43887 ( .A(reg_w_15[14]), .X(n49108) );
  inv_x1_sg U43888 ( .A(reg_w_15[13]), .X(n49106) );
  inv_x1_sg U43889 ( .A(reg_w_15[12]), .X(n49104) );
  inv_x1_sg U43890 ( .A(reg_w_15[11]), .X(n49102) );
  inv_x1_sg U43891 ( .A(reg_w_15[10]), .X(n49100) );
  inv_x1_sg U43892 ( .A(reg_w_15[9]), .X(n49098) );
  inv_x1_sg U43893 ( .A(reg_w_15[8]), .X(n49096) );
  inv_x1_sg U43894 ( .A(reg_w_15[7]), .X(n49094) );
  inv_x1_sg U43895 ( .A(reg_w_15[6]), .X(n49092) );
  inv_x1_sg U43896 ( .A(reg_w_15[5]), .X(n49090) );
  inv_x1_sg U43897 ( .A(reg_w_15[4]), .X(n49088) );
  inv_x1_sg U43898 ( .A(reg_w_15[3]), .X(n49086) );
  inv_x1_sg U43899 ( .A(reg_w_15[2]), .X(n49084) );
  inv_x1_sg U43900 ( .A(reg_w_15[1]), .X(n49082) );
  inv_x1_sg U43901 ( .A(reg_w_15[0]), .X(n49080) );
  inv_x1_sg U43902 ( .A(reg_w_14[19]), .X(n49078) );
  inv_x1_sg U43903 ( .A(reg_w_14[18]), .X(n49076) );
  inv_x1_sg U43904 ( .A(reg_w_14[17]), .X(n49074) );
  inv_x1_sg U43905 ( .A(reg_w_14[16]), .X(n49072) );
  inv_x1_sg U43906 ( .A(reg_w_14[15]), .X(n49070) );
  inv_x1_sg U43907 ( .A(reg_w_14[14]), .X(n49068) );
  inv_x1_sg U43908 ( .A(reg_w_14[13]), .X(n49066) );
  inv_x1_sg U43909 ( .A(reg_w_14[12]), .X(n49064) );
  inv_x1_sg U43910 ( .A(reg_w_14[11]), .X(n49062) );
  inv_x1_sg U43911 ( .A(reg_w_14[10]), .X(n49060) );
  inv_x1_sg U43912 ( .A(reg_w_14[9]), .X(n49058) );
  inv_x1_sg U43913 ( .A(reg_w_14[8]), .X(n49056) );
  inv_x1_sg U43914 ( .A(reg_w_14[7]), .X(n49054) );
  inv_x1_sg U43915 ( .A(reg_w_14[6]), .X(n49052) );
  inv_x1_sg U43916 ( .A(reg_w_14[5]), .X(n49050) );
  inv_x1_sg U43917 ( .A(reg_w_14[4]), .X(n49048) );
  inv_x1_sg U43918 ( .A(reg_w_14[3]), .X(n49046) );
  inv_x1_sg U43919 ( .A(reg_w_14[2]), .X(n49044) );
  inv_x1_sg U43920 ( .A(reg_w_14[1]), .X(n49042) );
  inv_x1_sg U43921 ( .A(reg_w_14[0]), .X(n49040) );
  inv_x1_sg U43922 ( .A(reg_w_13[19]), .X(n49038) );
  inv_x1_sg U43923 ( .A(reg_w_13[18]), .X(n49036) );
  inv_x1_sg U43924 ( .A(reg_w_13[17]), .X(n49034) );
  inv_x1_sg U43925 ( .A(reg_w_13[16]), .X(n49032) );
  inv_x1_sg U43926 ( .A(reg_w_13[15]), .X(n49030) );
  inv_x1_sg U43927 ( .A(reg_w_13[14]), .X(n49028) );
  inv_x1_sg U43928 ( .A(reg_w_13[13]), .X(n49026) );
  inv_x1_sg U43929 ( .A(reg_w_13[12]), .X(n49024) );
  inv_x1_sg U43930 ( .A(reg_w_13[11]), .X(n49022) );
  inv_x1_sg U43931 ( .A(reg_w_13[10]), .X(n49020) );
  inv_x1_sg U43932 ( .A(reg_w_13[9]), .X(n49018) );
  inv_x1_sg U43933 ( .A(reg_w_13[8]), .X(n49016) );
  inv_x1_sg U43934 ( .A(reg_w_13[7]), .X(n49014) );
  inv_x1_sg U43935 ( .A(reg_w_13[6]), .X(n49012) );
  inv_x1_sg U43936 ( .A(reg_w_13[5]), .X(n49010) );
  inv_x1_sg U43937 ( .A(reg_w_13[4]), .X(n49008) );
  inv_x1_sg U43938 ( .A(reg_w_13[3]), .X(n49006) );
  inv_x1_sg U43939 ( .A(reg_w_13[2]), .X(n49004) );
  inv_x1_sg U43940 ( .A(reg_w_13[1]), .X(n49002) );
  inv_x1_sg U43941 ( .A(reg_w_13[0]), .X(n49000) );
  inv_x1_sg U43942 ( .A(reg_w_12[19]), .X(n48998) );
  inv_x1_sg U43943 ( .A(reg_w_12[18]), .X(n48996) );
  inv_x1_sg U43944 ( .A(reg_w_12[17]), .X(n48994) );
  inv_x1_sg U43945 ( .A(reg_w_12[16]), .X(n48992) );
  inv_x1_sg U43946 ( .A(reg_w_12[15]), .X(n48990) );
  inv_x1_sg U43947 ( .A(reg_w_12[14]), .X(n48988) );
  inv_x1_sg U43948 ( .A(reg_w_12[13]), .X(n48986) );
  inv_x1_sg U43949 ( .A(reg_w_12[12]), .X(n48984) );
  inv_x1_sg U43950 ( .A(reg_w_12[11]), .X(n48982) );
  inv_x1_sg U43951 ( .A(reg_w_12[10]), .X(n48980) );
  inv_x1_sg U43952 ( .A(reg_w_12[9]), .X(n48978) );
  inv_x1_sg U43953 ( .A(reg_w_12[8]), .X(n48976) );
  inv_x1_sg U43954 ( .A(reg_w_12[7]), .X(n48974) );
  inv_x1_sg U43955 ( .A(reg_w_12[6]), .X(n48972) );
  inv_x1_sg U43956 ( .A(reg_w_12[5]), .X(n48970) );
  inv_x1_sg U43957 ( .A(reg_w_12[4]), .X(n48968) );
  inv_x1_sg U43958 ( .A(reg_w_12[3]), .X(n48966) );
  inv_x1_sg U43959 ( .A(reg_w_12[2]), .X(n48964) );
  inv_x1_sg U43960 ( .A(reg_w_12[1]), .X(n48962) );
  inv_x1_sg U43961 ( .A(reg_w_12[0]), .X(n48960) );
  inv_x1_sg U43962 ( .A(reg_w_11[19]), .X(n48958) );
  inv_x1_sg U43963 ( .A(reg_w_11[18]), .X(n48956) );
  inv_x1_sg U43964 ( .A(reg_w_11[17]), .X(n48954) );
  inv_x1_sg U43965 ( .A(reg_w_11[16]), .X(n48952) );
  inv_x1_sg U43966 ( .A(reg_w_11[15]), .X(n48950) );
  inv_x1_sg U43967 ( .A(reg_w_11[14]), .X(n48948) );
  inv_x1_sg U43968 ( .A(reg_w_11[13]), .X(n48946) );
  inv_x1_sg U43969 ( .A(reg_w_11[12]), .X(n48944) );
  inv_x1_sg U43970 ( .A(reg_w_11[11]), .X(n48942) );
  inv_x1_sg U43971 ( .A(reg_w_11[10]), .X(n48940) );
  inv_x1_sg U43972 ( .A(reg_w_11[9]), .X(n48938) );
  inv_x1_sg U43973 ( .A(reg_w_11[8]), .X(n48936) );
  inv_x1_sg U43974 ( .A(reg_w_11[7]), .X(n48934) );
  inv_x1_sg U43975 ( .A(reg_w_11[6]), .X(n48932) );
  inv_x1_sg U43976 ( .A(reg_w_11[5]), .X(n48930) );
  inv_x1_sg U43977 ( .A(reg_w_11[4]), .X(n48928) );
  inv_x1_sg U43978 ( .A(reg_w_11[3]), .X(n48926) );
  inv_x1_sg U43979 ( .A(reg_w_11[2]), .X(n48924) );
  inv_x1_sg U43980 ( .A(reg_w_11[1]), .X(n48922) );
  inv_x1_sg U43981 ( .A(reg_w_11[0]), .X(n48920) );
  inv_x1_sg U43982 ( .A(reg_w_10[19]), .X(n48918) );
  inv_x1_sg U43983 ( .A(reg_w_10[18]), .X(n48916) );
  inv_x1_sg U43984 ( .A(reg_w_10[17]), .X(n48914) );
  inv_x1_sg U43985 ( .A(reg_w_10[16]), .X(n48912) );
  inv_x1_sg U43986 ( .A(reg_w_10[15]), .X(n48910) );
  inv_x1_sg U43987 ( .A(reg_w_10[14]), .X(n48908) );
  inv_x1_sg U43988 ( .A(reg_w_10[13]), .X(n48906) );
  inv_x1_sg U43989 ( .A(reg_w_10[12]), .X(n48904) );
  inv_x1_sg U43990 ( .A(reg_w_10[11]), .X(n48902) );
  inv_x1_sg U43991 ( .A(reg_w_10[10]), .X(n48900) );
  inv_x1_sg U43992 ( .A(reg_w_10[9]), .X(n48898) );
  inv_x1_sg U43993 ( .A(reg_w_10[8]), .X(n48896) );
  inv_x1_sg U43994 ( .A(reg_w_10[7]), .X(n48894) );
  inv_x1_sg U43995 ( .A(reg_w_10[6]), .X(n48892) );
  inv_x1_sg U43996 ( .A(reg_w_10[5]), .X(n48890) );
  inv_x1_sg U43997 ( .A(reg_w_10[4]), .X(n48888) );
  inv_x1_sg U43998 ( .A(reg_w_10[3]), .X(n48886) );
  inv_x1_sg U43999 ( .A(reg_w_10[2]), .X(n48884) );
  inv_x1_sg U44000 ( .A(reg_w_10[1]), .X(n48882) );
  inv_x1_sg U44001 ( .A(reg_w_10[0]), .X(n48880) );
  inv_x1_sg U44002 ( .A(reg_w_9[19]), .X(n48878) );
  inv_x1_sg U44003 ( .A(reg_w_9[18]), .X(n48876) );
  inv_x1_sg U44004 ( .A(reg_w_9[17]), .X(n48874) );
  inv_x1_sg U44005 ( .A(reg_w_9[16]), .X(n48872) );
  inv_x1_sg U44006 ( .A(reg_w_9[15]), .X(n48870) );
  inv_x1_sg U44007 ( .A(reg_w_9[14]), .X(n48868) );
  inv_x1_sg U44008 ( .A(reg_w_9[13]), .X(n48866) );
  inv_x1_sg U44009 ( .A(reg_w_9[12]), .X(n48864) );
  inv_x1_sg U44010 ( .A(reg_w_9[11]), .X(n48862) );
  inv_x1_sg U44011 ( .A(reg_w_9[10]), .X(n48860) );
  inv_x1_sg U44012 ( .A(reg_w_9[9]), .X(n48858) );
  inv_x1_sg U44013 ( .A(reg_w_9[8]), .X(n48856) );
  inv_x1_sg U44014 ( .A(reg_w_9[7]), .X(n48854) );
  inv_x1_sg U44015 ( .A(reg_w_9[6]), .X(n48852) );
  inv_x1_sg U44016 ( .A(reg_w_9[5]), .X(n48850) );
  inv_x1_sg U44017 ( .A(reg_w_9[4]), .X(n48848) );
  inv_x1_sg U44018 ( .A(reg_w_9[3]), .X(n48846) );
  inv_x1_sg U44019 ( .A(reg_w_9[2]), .X(n48844) );
  inv_x1_sg U44020 ( .A(reg_w_9[1]), .X(n48842) );
  inv_x1_sg U44021 ( .A(reg_w_9[0]), .X(n48840) );
  inv_x1_sg U44022 ( .A(reg_w_8[19]), .X(n48838) );
  inv_x1_sg U44023 ( .A(reg_w_8[18]), .X(n48836) );
  inv_x1_sg U44024 ( .A(reg_w_8[17]), .X(n48834) );
  inv_x1_sg U44025 ( .A(reg_w_8[16]), .X(n48832) );
  inv_x1_sg U44026 ( .A(reg_w_8[15]), .X(n48830) );
  inv_x1_sg U44027 ( .A(reg_w_8[14]), .X(n48828) );
  inv_x1_sg U44028 ( .A(reg_w_8[13]), .X(n48826) );
  inv_x1_sg U44029 ( .A(reg_w_8[12]), .X(n48824) );
  inv_x1_sg U44030 ( .A(reg_w_8[11]), .X(n48822) );
  inv_x1_sg U44031 ( .A(reg_w_8[10]), .X(n48820) );
  inv_x1_sg U44032 ( .A(reg_w_8[9]), .X(n48818) );
  inv_x1_sg U44033 ( .A(reg_w_8[8]), .X(n48816) );
  inv_x1_sg U44034 ( .A(reg_w_8[7]), .X(n48814) );
  inv_x1_sg U44035 ( .A(reg_w_8[6]), .X(n48812) );
  inv_x1_sg U44036 ( .A(reg_w_8[5]), .X(n48810) );
  inv_x1_sg U44037 ( .A(reg_w_8[4]), .X(n48808) );
  inv_x1_sg U44038 ( .A(reg_w_8[3]), .X(n48806) );
  inv_x1_sg U44039 ( .A(reg_w_8[2]), .X(n48804) );
  inv_x1_sg U44040 ( .A(reg_w_8[1]), .X(n48802) );
  inv_x1_sg U44041 ( .A(reg_w_8[0]), .X(n48800) );
  inv_x1_sg U44042 ( .A(reg_w_7[19]), .X(n48798) );
  inv_x1_sg U44043 ( .A(reg_w_7[18]), .X(n48796) );
  inv_x1_sg U44044 ( .A(reg_w_7[17]), .X(n48794) );
  inv_x1_sg U44045 ( .A(reg_w_7[16]), .X(n48792) );
  inv_x1_sg U44046 ( .A(reg_w_7[15]), .X(n48790) );
  inv_x1_sg U44047 ( .A(reg_w_7[14]), .X(n48788) );
  inv_x1_sg U44048 ( .A(reg_w_7[13]), .X(n48786) );
  inv_x1_sg U44049 ( .A(reg_w_7[12]), .X(n48784) );
  inv_x1_sg U44050 ( .A(reg_w_7[11]), .X(n48782) );
  inv_x1_sg U44051 ( .A(reg_w_7[10]), .X(n48780) );
  inv_x1_sg U44052 ( .A(reg_w_7[9]), .X(n48778) );
  inv_x1_sg U44053 ( .A(reg_w_7[8]), .X(n48776) );
  inv_x1_sg U44054 ( .A(reg_w_7[7]), .X(n48774) );
  inv_x1_sg U44055 ( .A(reg_w_7[6]), .X(n48772) );
  inv_x1_sg U44056 ( .A(reg_w_7[5]), .X(n48770) );
  inv_x1_sg U44057 ( .A(reg_w_7[4]), .X(n48768) );
  inv_x1_sg U44058 ( .A(reg_w_7[3]), .X(n48766) );
  inv_x1_sg U44059 ( .A(reg_w_7[2]), .X(n48764) );
  inv_x1_sg U44060 ( .A(reg_w_7[1]), .X(n48762) );
  inv_x1_sg U44061 ( .A(reg_w_7[0]), .X(n48760) );
  inv_x1_sg U44062 ( .A(reg_w_6[19]), .X(n48758) );
  inv_x1_sg U44063 ( .A(reg_w_6[18]), .X(n48756) );
  inv_x1_sg U44064 ( .A(reg_w_6[17]), .X(n48754) );
  inv_x1_sg U44065 ( .A(reg_w_6[16]), .X(n48752) );
  inv_x1_sg U44066 ( .A(reg_w_6[15]), .X(n48750) );
  inv_x1_sg U44067 ( .A(reg_w_6[14]), .X(n48748) );
  inv_x1_sg U44068 ( .A(reg_w_6[13]), .X(n48746) );
  inv_x1_sg U44069 ( .A(reg_w_6[12]), .X(n48744) );
  inv_x1_sg U44070 ( .A(reg_w_6[11]), .X(n48742) );
  inv_x1_sg U44071 ( .A(reg_w_6[10]), .X(n48740) );
  inv_x1_sg U44072 ( .A(reg_w_6[9]), .X(n48738) );
  inv_x1_sg U44073 ( .A(reg_w_6[8]), .X(n48736) );
  inv_x1_sg U44074 ( .A(reg_w_6[7]), .X(n48734) );
  inv_x1_sg U44075 ( .A(reg_w_6[6]), .X(n48732) );
  inv_x1_sg U44076 ( .A(reg_w_6[5]), .X(n48730) );
  inv_x1_sg U44077 ( .A(reg_w_6[4]), .X(n48728) );
  inv_x1_sg U44078 ( .A(reg_w_6[3]), .X(n48726) );
  inv_x1_sg U44079 ( .A(reg_w_6[2]), .X(n48724) );
  inv_x1_sg U44080 ( .A(reg_w_6[1]), .X(n48722) );
  inv_x1_sg U44081 ( .A(reg_w_6[0]), .X(n48720) );
  inv_x1_sg U44082 ( .A(reg_w_5[19]), .X(n48718) );
  inv_x1_sg U44083 ( .A(reg_w_5[18]), .X(n48716) );
  inv_x1_sg U44084 ( .A(reg_w_5[17]), .X(n48714) );
  inv_x1_sg U44085 ( .A(reg_w_5[16]), .X(n48712) );
  inv_x1_sg U44086 ( .A(reg_w_5[15]), .X(n48710) );
  inv_x1_sg U44087 ( .A(reg_w_5[14]), .X(n48708) );
  inv_x1_sg U44088 ( .A(reg_w_5[13]), .X(n48706) );
  inv_x1_sg U44089 ( .A(reg_w_5[12]), .X(n48704) );
  inv_x1_sg U44090 ( .A(reg_w_5[11]), .X(n48702) );
  inv_x1_sg U44091 ( .A(reg_w_5[10]), .X(n48700) );
  inv_x1_sg U44092 ( .A(reg_w_5[9]), .X(n48698) );
  inv_x1_sg U44093 ( .A(reg_w_5[8]), .X(n48696) );
  inv_x1_sg U44094 ( .A(reg_w_5[7]), .X(n48694) );
  inv_x1_sg U44095 ( .A(reg_w_5[6]), .X(n48692) );
  inv_x1_sg U44096 ( .A(reg_w_5[5]), .X(n48690) );
  inv_x1_sg U44097 ( .A(reg_w_5[4]), .X(n48688) );
  inv_x1_sg U44098 ( .A(reg_w_5[3]), .X(n48686) );
  inv_x1_sg U44099 ( .A(reg_w_5[2]), .X(n48684) );
  inv_x1_sg U44100 ( .A(reg_w_5[1]), .X(n48682) );
  inv_x1_sg U44101 ( .A(reg_w_5[0]), .X(n48680) );
  inv_x1_sg U44102 ( .A(reg_w_4[19]), .X(n48678) );
  inv_x1_sg U44103 ( .A(reg_w_4[18]), .X(n48676) );
  inv_x1_sg U44104 ( .A(reg_w_4[17]), .X(n48674) );
  inv_x1_sg U44105 ( .A(reg_w_4[16]), .X(n48672) );
  inv_x1_sg U44106 ( .A(reg_w_4[15]), .X(n48670) );
  inv_x1_sg U44107 ( .A(reg_w_4[14]), .X(n48668) );
  inv_x1_sg U44108 ( .A(reg_w_4[13]), .X(n48666) );
  inv_x1_sg U44109 ( .A(reg_w_4[12]), .X(n48664) );
  inv_x1_sg U44110 ( .A(reg_w_4[11]), .X(n48662) );
  inv_x1_sg U44111 ( .A(reg_w_4[10]), .X(n48660) );
  inv_x1_sg U44112 ( .A(reg_w_4[9]), .X(n48658) );
  inv_x1_sg U44113 ( .A(reg_w_4[8]), .X(n48656) );
  inv_x1_sg U44114 ( .A(reg_w_4[7]), .X(n48654) );
  inv_x1_sg U44115 ( .A(reg_w_4[6]), .X(n48652) );
  inv_x1_sg U44116 ( .A(reg_w_4[5]), .X(n48650) );
  inv_x1_sg U44117 ( .A(reg_w_4[4]), .X(n48648) );
  inv_x1_sg U44118 ( .A(reg_w_4[3]), .X(n48646) );
  inv_x1_sg U44119 ( .A(reg_w_4[2]), .X(n48644) );
  inv_x1_sg U44120 ( .A(reg_w_4[1]), .X(n48642) );
  inv_x1_sg U44121 ( .A(reg_w_4[0]), .X(n48640) );
  inv_x1_sg U44122 ( .A(reg_w_3[19]), .X(n48638) );
  inv_x1_sg U44123 ( .A(reg_w_3[18]), .X(n48636) );
  inv_x1_sg U44124 ( .A(reg_w_3[17]), .X(n48634) );
  inv_x1_sg U44125 ( .A(reg_w_3[16]), .X(n48632) );
  inv_x1_sg U44126 ( .A(reg_w_3[15]), .X(n48630) );
  inv_x1_sg U44127 ( .A(reg_w_3[14]), .X(n48628) );
  inv_x1_sg U44128 ( .A(reg_w_3[13]), .X(n48626) );
  inv_x1_sg U44129 ( .A(reg_w_3[12]), .X(n48624) );
  inv_x1_sg U44130 ( .A(reg_w_3[11]), .X(n48622) );
  inv_x1_sg U44131 ( .A(reg_w_3[10]), .X(n48620) );
  inv_x1_sg U44132 ( .A(reg_w_3[9]), .X(n48618) );
  inv_x1_sg U44133 ( .A(reg_w_3[8]), .X(n48616) );
  inv_x1_sg U44134 ( .A(reg_w_3[7]), .X(n48614) );
  inv_x1_sg U44135 ( .A(reg_w_3[6]), .X(n48612) );
  inv_x1_sg U44136 ( .A(reg_w_3[5]), .X(n48610) );
  inv_x1_sg U44137 ( .A(reg_w_3[4]), .X(n48608) );
  inv_x1_sg U44138 ( .A(reg_w_3[3]), .X(n48606) );
  inv_x1_sg U44139 ( .A(reg_w_3[2]), .X(n48604) );
  inv_x1_sg U44140 ( .A(reg_w_3[1]), .X(n48602) );
  inv_x1_sg U44141 ( .A(reg_w_3[0]), .X(n48600) );
  inv_x1_sg U44142 ( .A(reg_w_2[19]), .X(n48598) );
  inv_x1_sg U44143 ( .A(reg_w_2[18]), .X(n48596) );
  inv_x1_sg U44144 ( .A(reg_w_2[17]), .X(n48594) );
  inv_x1_sg U44145 ( .A(reg_w_2[16]), .X(n48592) );
  inv_x1_sg U44146 ( .A(reg_w_2[15]), .X(n48590) );
  inv_x1_sg U44147 ( .A(reg_w_2[14]), .X(n48588) );
  inv_x1_sg U44148 ( .A(reg_w_2[13]), .X(n48586) );
  inv_x1_sg U44149 ( .A(reg_w_2[12]), .X(n48584) );
  inv_x1_sg U44150 ( .A(reg_w_2[11]), .X(n48582) );
  inv_x1_sg U44151 ( .A(reg_w_2[10]), .X(n48580) );
  inv_x1_sg U44152 ( .A(reg_w_2[9]), .X(n48578) );
  inv_x1_sg U44153 ( .A(reg_w_2[8]), .X(n48576) );
  inv_x1_sg U44154 ( .A(reg_w_2[7]), .X(n48574) );
  inv_x1_sg U44155 ( .A(reg_w_2[6]), .X(n48572) );
  inv_x1_sg U44156 ( .A(reg_w_2[5]), .X(n48570) );
  inv_x1_sg U44157 ( .A(reg_w_2[4]), .X(n48568) );
  inv_x1_sg U44158 ( .A(reg_w_2[3]), .X(n48566) );
  inv_x1_sg U44159 ( .A(reg_w_2[2]), .X(n48564) );
  inv_x1_sg U44160 ( .A(reg_w_2[1]), .X(n48562) );
  inv_x1_sg U44161 ( .A(reg_w_2[0]), .X(n48560) );
  inv_x1_sg U44162 ( .A(reg_w_1[19]), .X(n48558) );
  inv_x1_sg U44163 ( .A(reg_w_1[18]), .X(n48556) );
  inv_x1_sg U44164 ( .A(reg_w_1[17]), .X(n48554) );
  inv_x1_sg U44165 ( .A(reg_w_1[16]), .X(n48552) );
  inv_x1_sg U44166 ( .A(reg_w_1[15]), .X(n48550) );
  inv_x1_sg U44167 ( .A(reg_w_1[14]), .X(n48548) );
  inv_x1_sg U44168 ( .A(reg_w_1[13]), .X(n48546) );
  inv_x1_sg U44169 ( .A(reg_w_1[12]), .X(n48544) );
  inv_x1_sg U44170 ( .A(reg_w_1[11]), .X(n48542) );
  inv_x1_sg U44171 ( .A(reg_w_1[10]), .X(n48540) );
  inv_x1_sg U44172 ( .A(reg_w_1[9]), .X(n48538) );
  inv_x1_sg U44173 ( .A(reg_w_1[8]), .X(n48536) );
  inv_x1_sg U44174 ( .A(reg_w_1[7]), .X(n48534) );
  inv_x1_sg U44175 ( .A(reg_w_1[6]), .X(n48532) );
  inv_x1_sg U44176 ( .A(reg_w_1[5]), .X(n48530) );
  inv_x1_sg U44177 ( .A(reg_w_1[4]), .X(n48528) );
  inv_x1_sg U44178 ( .A(reg_w_1[3]), .X(n48526) );
  inv_x1_sg U44179 ( .A(reg_w_1[2]), .X(n48524) );
  inv_x1_sg U44180 ( .A(reg_w_1[1]), .X(n48522) );
  inv_x1_sg U44181 ( .A(reg_w_1[0]), .X(n48520) );
  inv_x1_sg U44182 ( .A(reg_w_0[19]), .X(n48518) );
  inv_x1_sg U44183 ( .A(reg_w_0[18]), .X(n48516) );
  inv_x1_sg U44184 ( .A(reg_w_0[17]), .X(n48514) );
  inv_x1_sg U44185 ( .A(reg_w_0[16]), .X(n48512) );
  inv_x1_sg U44186 ( .A(reg_w_0[15]), .X(n48510) );
  inv_x1_sg U44187 ( .A(reg_w_0[14]), .X(n48508) );
  inv_x1_sg U44188 ( .A(reg_w_0[13]), .X(n48506) );
  inv_x1_sg U44189 ( .A(reg_w_0[12]), .X(n48504) );
  inv_x1_sg U44190 ( .A(reg_w_0[11]), .X(n48502) );
  inv_x1_sg U44191 ( .A(reg_w_0[10]), .X(n48500) );
  inv_x1_sg U44192 ( .A(reg_w_0[9]), .X(n48498) );
  inv_x1_sg U44193 ( .A(reg_w_0[8]), .X(n48496) );
  inv_x1_sg U44194 ( .A(reg_w_0[7]), .X(n48494) );
  inv_x1_sg U44195 ( .A(reg_w_0[6]), .X(n48492) );
  inv_x1_sg U44196 ( .A(reg_w_0[5]), .X(n48490) );
  inv_x1_sg U44197 ( .A(reg_w_0[4]), .X(n48488) );
  inv_x1_sg U44198 ( .A(reg_w_0[3]), .X(n48486) );
  inv_x1_sg U44199 ( .A(reg_w_0[2]), .X(n48484) );
  inv_x1_sg U44200 ( .A(reg_w_0[1]), .X(n48482) );
  inv_x1_sg U44201 ( .A(reg_w_0[0]), .X(n48480) );
  inv_x1_sg U44202 ( .A(reg_i_15[19]), .X(n48478) );
  inv_x1_sg U44203 ( .A(reg_i_15[18]), .X(n48476) );
  inv_x1_sg U44204 ( .A(reg_i_15[17]), .X(n48474) );
  inv_x1_sg U44205 ( .A(reg_i_15[16]), .X(n48472) );
  inv_x1_sg U44206 ( .A(reg_i_15[15]), .X(n48470) );
  inv_x1_sg U44207 ( .A(reg_i_15[14]), .X(n48468) );
  inv_x1_sg U44208 ( .A(reg_i_15[13]), .X(n48466) );
  inv_x1_sg U44209 ( .A(reg_i_15[12]), .X(n48464) );
  inv_x1_sg U44210 ( .A(reg_i_15[11]), .X(n48462) );
  inv_x1_sg U44211 ( .A(reg_i_15[10]), .X(n48460) );
  inv_x1_sg U44212 ( .A(reg_i_15[9]), .X(n48458) );
  inv_x1_sg U44213 ( .A(reg_i_15[8]), .X(n48456) );
  inv_x1_sg U44214 ( .A(reg_i_15[7]), .X(n48454) );
  inv_x1_sg U44215 ( .A(reg_i_15[6]), .X(n48452) );
  inv_x1_sg U44216 ( .A(reg_i_15[5]), .X(n48450) );
  inv_x1_sg U44217 ( .A(reg_i_15[4]), .X(n48448) );
  inv_x1_sg U44218 ( .A(reg_i_15[3]), .X(n48446) );
  inv_x1_sg U44219 ( .A(reg_i_15[2]), .X(n48444) );
  inv_x1_sg U44220 ( .A(reg_i_15[1]), .X(n48442) );
  inv_x1_sg U44221 ( .A(reg_i_15[0]), .X(n48440) );
  inv_x1_sg U44222 ( .A(reg_i_14[19]), .X(n48438) );
  inv_x1_sg U44223 ( .A(reg_i_14[18]), .X(n48436) );
  inv_x1_sg U44224 ( .A(reg_i_14[17]), .X(n48434) );
  inv_x1_sg U44225 ( .A(reg_i_14[16]), .X(n48432) );
  inv_x1_sg U44226 ( .A(reg_i_14[15]), .X(n48430) );
  inv_x1_sg U44227 ( .A(reg_i_14[14]), .X(n48428) );
  inv_x1_sg U44228 ( .A(reg_i_14[13]), .X(n48426) );
  inv_x1_sg U44229 ( .A(reg_i_14[12]), .X(n48424) );
  inv_x1_sg U44230 ( .A(reg_i_14[11]), .X(n48422) );
  inv_x1_sg U44231 ( .A(reg_i_14[10]), .X(n48420) );
  inv_x1_sg U44232 ( .A(reg_i_14[9]), .X(n48418) );
  inv_x1_sg U44233 ( .A(reg_i_14[8]), .X(n48416) );
  inv_x1_sg U44234 ( .A(reg_i_14[7]), .X(n48414) );
  inv_x1_sg U44235 ( .A(reg_i_14[6]), .X(n48412) );
  inv_x1_sg U44236 ( .A(reg_i_14[5]), .X(n48410) );
  inv_x1_sg U44237 ( .A(reg_i_14[4]), .X(n48408) );
  inv_x1_sg U44238 ( .A(reg_i_14[3]), .X(n48406) );
  inv_x1_sg U44239 ( .A(reg_i_14[2]), .X(n48404) );
  inv_x1_sg U44240 ( .A(reg_i_14[1]), .X(n48402) );
  inv_x1_sg U44241 ( .A(reg_i_14[0]), .X(n48400) );
  inv_x1_sg U44242 ( .A(reg_i_13[19]), .X(n48398) );
  inv_x1_sg U44243 ( .A(reg_i_13[18]), .X(n48396) );
  inv_x1_sg U44244 ( .A(reg_i_13[17]), .X(n48394) );
  inv_x1_sg U44245 ( .A(reg_i_13[16]), .X(n48392) );
  inv_x1_sg U44246 ( .A(reg_i_13[15]), .X(n48390) );
  inv_x1_sg U44247 ( .A(reg_i_13[14]), .X(n48388) );
  inv_x1_sg U44248 ( .A(reg_i_13[13]), .X(n48386) );
  inv_x1_sg U44249 ( .A(reg_i_13[12]), .X(n48384) );
  inv_x1_sg U44250 ( .A(reg_i_13[11]), .X(n48382) );
  inv_x1_sg U44251 ( .A(reg_i_13[10]), .X(n48380) );
  inv_x1_sg U44252 ( .A(reg_i_13[9]), .X(n48378) );
  inv_x1_sg U44253 ( .A(reg_i_13[8]), .X(n48376) );
  inv_x1_sg U44254 ( .A(reg_i_13[7]), .X(n48374) );
  inv_x1_sg U44255 ( .A(reg_i_13[6]), .X(n48372) );
  inv_x1_sg U44256 ( .A(reg_i_13[5]), .X(n48370) );
  inv_x1_sg U44257 ( .A(reg_i_13[4]), .X(n48368) );
  inv_x1_sg U44258 ( .A(reg_i_13[3]), .X(n48366) );
  inv_x1_sg U44259 ( .A(reg_i_13[2]), .X(n48364) );
  inv_x1_sg U44260 ( .A(reg_i_13[1]), .X(n48362) );
  inv_x1_sg U44261 ( .A(reg_i_13[0]), .X(n48360) );
  inv_x1_sg U44262 ( .A(reg_i_12[19]), .X(n48358) );
  inv_x1_sg U44263 ( .A(reg_i_12[18]), .X(n48356) );
  inv_x1_sg U44264 ( .A(reg_i_12[17]), .X(n48354) );
  inv_x1_sg U44265 ( .A(reg_i_12[16]), .X(n48352) );
  inv_x1_sg U44266 ( .A(reg_i_12[15]), .X(n48350) );
  inv_x1_sg U44267 ( .A(reg_i_12[14]), .X(n48348) );
  inv_x1_sg U44268 ( .A(reg_i_12[13]), .X(n48346) );
  inv_x1_sg U44269 ( .A(reg_i_12[12]), .X(n48344) );
  inv_x1_sg U44270 ( .A(reg_i_12[11]), .X(n48342) );
  inv_x1_sg U44271 ( .A(reg_i_12[10]), .X(n48340) );
  inv_x1_sg U44272 ( .A(reg_i_12[9]), .X(n48338) );
  inv_x1_sg U44273 ( .A(reg_i_12[8]), .X(n48336) );
  inv_x1_sg U44274 ( .A(reg_i_12[7]), .X(n48334) );
  inv_x1_sg U44275 ( .A(reg_i_12[6]), .X(n48332) );
  inv_x1_sg U44276 ( .A(reg_i_12[5]), .X(n48330) );
  inv_x1_sg U44277 ( .A(reg_i_12[4]), .X(n48328) );
  inv_x1_sg U44278 ( .A(reg_i_12[3]), .X(n48326) );
  inv_x1_sg U44279 ( .A(reg_i_12[2]), .X(n48324) );
  inv_x1_sg U44280 ( .A(reg_i_12[1]), .X(n48322) );
  inv_x1_sg U44281 ( .A(reg_i_12[0]), .X(n48320) );
  inv_x1_sg U44282 ( .A(reg_i_11[19]), .X(n48318) );
  inv_x1_sg U44283 ( .A(reg_i_11[18]), .X(n48316) );
  inv_x1_sg U44284 ( .A(reg_i_11[17]), .X(n48314) );
  inv_x1_sg U44285 ( .A(reg_i_11[16]), .X(n48312) );
  inv_x1_sg U44286 ( .A(reg_i_11[15]), .X(n48310) );
  inv_x1_sg U44287 ( .A(reg_i_11[14]), .X(n48308) );
  inv_x1_sg U44288 ( .A(reg_i_11[13]), .X(n48306) );
  inv_x1_sg U44289 ( .A(reg_i_11[12]), .X(n48304) );
  inv_x1_sg U44290 ( .A(reg_i_11[11]), .X(n48302) );
  inv_x1_sg U44291 ( .A(reg_i_11[10]), .X(n48300) );
  inv_x1_sg U44292 ( .A(reg_i_11[9]), .X(n48298) );
  inv_x1_sg U44293 ( .A(reg_i_11[8]), .X(n48296) );
  inv_x1_sg U44294 ( .A(reg_i_11[7]), .X(n48294) );
  inv_x1_sg U44295 ( .A(reg_i_11[6]), .X(n48292) );
  inv_x1_sg U44296 ( .A(reg_i_11[5]), .X(n48290) );
  inv_x1_sg U44297 ( .A(reg_i_11[4]), .X(n48288) );
  inv_x1_sg U44298 ( .A(reg_i_11[3]), .X(n48286) );
  inv_x1_sg U44299 ( .A(reg_i_11[2]), .X(n48284) );
  inv_x1_sg U44300 ( .A(reg_i_11[1]), .X(n48282) );
  inv_x1_sg U44301 ( .A(reg_i_11[0]), .X(n48280) );
  inv_x1_sg U44302 ( .A(reg_i_10[19]), .X(n48278) );
  inv_x1_sg U44303 ( .A(reg_i_10[18]), .X(n48276) );
  inv_x1_sg U44304 ( .A(reg_i_10[17]), .X(n48274) );
  inv_x1_sg U44305 ( .A(reg_i_10[16]), .X(n48272) );
  inv_x1_sg U44306 ( .A(reg_i_10[15]), .X(n48270) );
  inv_x1_sg U44307 ( .A(reg_i_10[14]), .X(n48268) );
  inv_x1_sg U44308 ( .A(reg_i_10[13]), .X(n48266) );
  inv_x1_sg U44309 ( .A(reg_i_10[12]), .X(n48264) );
  inv_x1_sg U44310 ( .A(reg_i_10[11]), .X(n48262) );
  inv_x1_sg U44311 ( .A(reg_i_10[10]), .X(n48260) );
  inv_x1_sg U44312 ( .A(reg_i_10[9]), .X(n48258) );
  inv_x1_sg U44313 ( .A(reg_i_10[8]), .X(n48256) );
  inv_x1_sg U44314 ( .A(reg_i_10[7]), .X(n48254) );
  inv_x1_sg U44315 ( .A(reg_i_10[6]), .X(n48252) );
  inv_x1_sg U44316 ( .A(reg_i_10[5]), .X(n48250) );
  inv_x1_sg U44317 ( .A(reg_i_10[4]), .X(n48248) );
  inv_x1_sg U44318 ( .A(reg_i_10[3]), .X(n48246) );
  inv_x1_sg U44319 ( .A(reg_i_10[2]), .X(n48244) );
  inv_x1_sg U44320 ( .A(reg_i_10[1]), .X(n48242) );
  inv_x1_sg U44321 ( .A(reg_i_10[0]), .X(n48240) );
  inv_x1_sg U44322 ( .A(reg_i_9[19]), .X(n48238) );
  inv_x1_sg U44323 ( .A(reg_i_9[18]), .X(n48236) );
  inv_x1_sg U44324 ( .A(reg_i_9[17]), .X(n48234) );
  inv_x1_sg U44325 ( .A(reg_i_9[16]), .X(n48232) );
  inv_x1_sg U44326 ( .A(reg_i_9[15]), .X(n48230) );
  inv_x1_sg U44327 ( .A(reg_i_9[14]), .X(n48228) );
  inv_x1_sg U44328 ( .A(reg_i_9[13]), .X(n48226) );
  inv_x1_sg U44329 ( .A(reg_i_9[12]), .X(n48224) );
  inv_x1_sg U44330 ( .A(reg_i_9[11]), .X(n48222) );
  inv_x1_sg U44331 ( .A(reg_i_9[10]), .X(n48220) );
  inv_x1_sg U44332 ( .A(reg_i_9[9]), .X(n48218) );
  inv_x1_sg U44333 ( .A(reg_i_9[8]), .X(n48216) );
  inv_x1_sg U44334 ( .A(reg_i_9[7]), .X(n48214) );
  inv_x1_sg U44335 ( .A(reg_i_9[6]), .X(n48212) );
  inv_x1_sg U44336 ( .A(reg_i_9[5]), .X(n48210) );
  inv_x1_sg U44337 ( .A(reg_i_9[4]), .X(n48208) );
  inv_x1_sg U44338 ( .A(reg_i_9[3]), .X(n48206) );
  inv_x1_sg U44339 ( .A(reg_i_9[2]), .X(n48204) );
  inv_x1_sg U44340 ( .A(reg_i_9[1]), .X(n48202) );
  inv_x1_sg U44341 ( .A(reg_i_9[0]), .X(n48200) );
  inv_x1_sg U44342 ( .A(reg_i_8[19]), .X(n48198) );
  inv_x1_sg U44343 ( .A(reg_i_8[18]), .X(n48196) );
  inv_x1_sg U44344 ( .A(reg_i_8[17]), .X(n48194) );
  inv_x1_sg U44345 ( .A(reg_i_8[16]), .X(n48192) );
  inv_x1_sg U44346 ( .A(reg_i_8[15]), .X(n48190) );
  inv_x1_sg U44347 ( .A(reg_i_8[14]), .X(n48188) );
  inv_x1_sg U44348 ( .A(reg_i_8[13]), .X(n48186) );
  inv_x1_sg U44349 ( .A(reg_i_8[12]), .X(n48184) );
  inv_x1_sg U44350 ( .A(reg_i_8[11]), .X(n48182) );
  inv_x1_sg U44351 ( .A(reg_i_8[10]), .X(n48180) );
  inv_x1_sg U44352 ( .A(reg_i_8[9]), .X(n48178) );
  inv_x1_sg U44353 ( .A(reg_i_8[8]), .X(n48176) );
  inv_x1_sg U44354 ( .A(reg_i_8[7]), .X(n48174) );
  inv_x1_sg U44355 ( .A(reg_i_8[6]), .X(n48172) );
  inv_x1_sg U44356 ( .A(reg_i_8[5]), .X(n48170) );
  inv_x1_sg U44357 ( .A(reg_i_8[4]), .X(n48168) );
  inv_x1_sg U44358 ( .A(reg_i_8[3]), .X(n48166) );
  inv_x1_sg U44359 ( .A(reg_i_8[2]), .X(n48164) );
  inv_x1_sg U44360 ( .A(reg_i_8[1]), .X(n48162) );
  inv_x1_sg U44361 ( .A(reg_i_8[0]), .X(n48160) );
  inv_x1_sg U44362 ( .A(reg_i_7[19]), .X(n48158) );
  inv_x1_sg U44363 ( .A(reg_i_7[18]), .X(n48156) );
  inv_x1_sg U44364 ( .A(reg_i_7[17]), .X(n48154) );
  inv_x1_sg U44365 ( .A(reg_i_7[16]), .X(n48152) );
  inv_x1_sg U44366 ( .A(reg_i_7[15]), .X(n48150) );
  inv_x1_sg U44367 ( .A(reg_i_7[14]), .X(n48148) );
  inv_x1_sg U44368 ( .A(reg_i_7[13]), .X(n48146) );
  inv_x1_sg U44369 ( .A(reg_i_7[12]), .X(n48144) );
  inv_x1_sg U44370 ( .A(reg_i_7[11]), .X(n48142) );
  inv_x1_sg U44371 ( .A(reg_i_7[10]), .X(n48140) );
  inv_x1_sg U44372 ( .A(reg_i_7[9]), .X(n48138) );
  inv_x1_sg U44373 ( .A(reg_i_7[8]), .X(n48136) );
  inv_x1_sg U44374 ( .A(reg_i_7[7]), .X(n48134) );
  inv_x1_sg U44375 ( .A(reg_i_7[6]), .X(n48132) );
  inv_x1_sg U44376 ( .A(reg_i_7[5]), .X(n48130) );
  inv_x1_sg U44377 ( .A(reg_i_7[4]), .X(n48128) );
  inv_x1_sg U44378 ( .A(reg_i_7[3]), .X(n48126) );
  inv_x1_sg U44379 ( .A(reg_i_7[2]), .X(n48124) );
  inv_x1_sg U44380 ( .A(reg_i_7[1]), .X(n48122) );
  inv_x1_sg U44381 ( .A(reg_i_7[0]), .X(n48120) );
  inv_x1_sg U44382 ( .A(reg_i_6[19]), .X(n48118) );
  inv_x1_sg U44383 ( .A(reg_i_6[18]), .X(n48116) );
  inv_x1_sg U44384 ( .A(reg_i_6[17]), .X(n48114) );
  inv_x1_sg U44385 ( .A(reg_i_6[16]), .X(n48112) );
  inv_x1_sg U44386 ( .A(reg_i_6[15]), .X(n48110) );
  inv_x1_sg U44387 ( .A(reg_i_6[14]), .X(n48108) );
  inv_x1_sg U44388 ( .A(reg_i_6[13]), .X(n48106) );
  inv_x1_sg U44389 ( .A(reg_i_6[12]), .X(n48104) );
  inv_x1_sg U44390 ( .A(reg_i_6[11]), .X(n48102) );
  inv_x1_sg U44391 ( .A(reg_i_6[10]), .X(n48100) );
  inv_x1_sg U44392 ( .A(reg_i_6[9]), .X(n48098) );
  inv_x1_sg U44393 ( .A(reg_i_6[8]), .X(n48096) );
  inv_x1_sg U44394 ( .A(reg_i_6[7]), .X(n48094) );
  inv_x1_sg U44395 ( .A(reg_i_6[6]), .X(n48092) );
  inv_x1_sg U44396 ( .A(reg_i_6[5]), .X(n48090) );
  inv_x1_sg U44397 ( .A(reg_i_6[4]), .X(n48088) );
  inv_x1_sg U44398 ( .A(reg_i_6[3]), .X(n48086) );
  inv_x1_sg U44399 ( .A(reg_i_6[2]), .X(n48084) );
  inv_x1_sg U44400 ( .A(reg_i_6[1]), .X(n48082) );
  inv_x1_sg U44401 ( .A(reg_i_6[0]), .X(n48080) );
  inv_x1_sg U44402 ( .A(reg_i_5[19]), .X(n48078) );
  inv_x1_sg U44403 ( .A(reg_i_5[18]), .X(n48076) );
  inv_x1_sg U44404 ( .A(reg_i_5[17]), .X(n48074) );
  inv_x1_sg U44405 ( .A(reg_i_5[16]), .X(n48072) );
  inv_x1_sg U44406 ( .A(reg_i_5[15]), .X(n48070) );
  inv_x1_sg U44407 ( .A(reg_i_5[14]), .X(n48068) );
  inv_x1_sg U44408 ( .A(reg_i_5[13]), .X(n48066) );
  inv_x1_sg U44409 ( .A(reg_i_5[12]), .X(n48064) );
  inv_x1_sg U44410 ( .A(reg_i_5[11]), .X(n48062) );
  inv_x1_sg U44411 ( .A(reg_i_5[10]), .X(n48060) );
  inv_x1_sg U44412 ( .A(reg_i_5[9]), .X(n48058) );
  inv_x1_sg U44413 ( .A(reg_i_5[8]), .X(n48056) );
  inv_x1_sg U44414 ( .A(reg_i_5[7]), .X(n48054) );
  inv_x1_sg U44415 ( .A(reg_i_5[6]), .X(n48052) );
  inv_x1_sg U44416 ( .A(reg_i_5[5]), .X(n48050) );
  inv_x1_sg U44417 ( .A(reg_i_5[4]), .X(n48048) );
  inv_x1_sg U44418 ( .A(reg_i_5[3]), .X(n48046) );
  inv_x1_sg U44419 ( .A(reg_i_5[2]), .X(n48044) );
  inv_x1_sg U44420 ( .A(reg_i_5[1]), .X(n48042) );
  inv_x1_sg U44421 ( .A(reg_i_5[0]), .X(n48040) );
  inv_x1_sg U44422 ( .A(reg_i_4[19]), .X(n48038) );
  inv_x1_sg U44423 ( .A(reg_i_4[18]), .X(n48036) );
  inv_x1_sg U44424 ( .A(reg_i_4[17]), .X(n48034) );
  inv_x1_sg U44425 ( .A(reg_i_4[16]), .X(n48032) );
  inv_x1_sg U44426 ( .A(reg_i_4[15]), .X(n48030) );
  inv_x1_sg U44427 ( .A(reg_i_4[14]), .X(n48028) );
  inv_x1_sg U44428 ( .A(reg_i_4[13]), .X(n48026) );
  inv_x1_sg U44429 ( .A(reg_i_4[12]), .X(n48024) );
  inv_x1_sg U44430 ( .A(reg_i_4[11]), .X(n48022) );
  inv_x1_sg U44431 ( .A(reg_i_4[10]), .X(n48020) );
  inv_x1_sg U44432 ( .A(reg_i_4[9]), .X(n48018) );
  inv_x1_sg U44433 ( .A(reg_i_4[8]), .X(n48016) );
  inv_x1_sg U44434 ( .A(reg_i_4[7]), .X(n48014) );
  inv_x1_sg U44435 ( .A(reg_i_4[6]), .X(n48012) );
  inv_x1_sg U44436 ( .A(reg_i_4[5]), .X(n48010) );
  inv_x1_sg U44437 ( .A(reg_i_4[4]), .X(n48008) );
  inv_x1_sg U44438 ( .A(reg_i_4[3]), .X(n48006) );
  inv_x1_sg U44439 ( .A(reg_i_4[2]), .X(n48004) );
  inv_x1_sg U44440 ( .A(reg_i_4[1]), .X(n48002) );
  inv_x1_sg U44441 ( .A(reg_i_4[0]), .X(n48000) );
  inv_x1_sg U44442 ( .A(reg_i_3[19]), .X(n47998) );
  inv_x1_sg U44443 ( .A(reg_i_3[18]), .X(n47996) );
  inv_x1_sg U44444 ( .A(reg_i_3[17]), .X(n47994) );
  inv_x1_sg U44445 ( .A(reg_i_3[16]), .X(n47992) );
  inv_x1_sg U44446 ( .A(reg_i_3[15]), .X(n47990) );
  inv_x1_sg U44447 ( .A(reg_i_3[14]), .X(n47988) );
  inv_x1_sg U44448 ( .A(reg_i_3[13]), .X(n47986) );
  inv_x1_sg U44449 ( .A(reg_i_3[12]), .X(n47984) );
  inv_x1_sg U44450 ( .A(reg_i_3[11]), .X(n47982) );
  inv_x1_sg U44451 ( .A(reg_i_3[10]), .X(n47980) );
  inv_x1_sg U44452 ( .A(reg_i_3[9]), .X(n47978) );
  inv_x1_sg U44453 ( .A(reg_i_3[8]), .X(n47976) );
  inv_x1_sg U44454 ( .A(reg_i_3[7]), .X(n47974) );
  inv_x1_sg U44455 ( .A(reg_i_3[6]), .X(n47972) );
  inv_x1_sg U44456 ( .A(reg_i_3[5]), .X(n47970) );
  inv_x1_sg U44457 ( .A(reg_i_3[4]), .X(n47968) );
  inv_x1_sg U44458 ( .A(reg_i_3[3]), .X(n47966) );
  inv_x1_sg U44459 ( .A(reg_i_3[2]), .X(n47964) );
  inv_x1_sg U44460 ( .A(reg_i_3[1]), .X(n47962) );
  inv_x1_sg U44461 ( .A(reg_i_3[0]), .X(n47960) );
  inv_x1_sg U44462 ( .A(reg_i_2[19]), .X(n47958) );
  inv_x1_sg U44463 ( .A(reg_i_2[18]), .X(n47956) );
  inv_x1_sg U44464 ( .A(reg_i_2[17]), .X(n47954) );
  inv_x1_sg U44465 ( .A(reg_i_2[16]), .X(n47952) );
  inv_x1_sg U44466 ( .A(reg_i_2[15]), .X(n47950) );
  inv_x1_sg U44467 ( .A(reg_i_2[14]), .X(n47948) );
  inv_x1_sg U44468 ( .A(reg_i_2[13]), .X(n47946) );
  inv_x1_sg U44469 ( .A(reg_i_2[12]), .X(n47944) );
  inv_x1_sg U44470 ( .A(reg_i_2[11]), .X(n47942) );
  inv_x1_sg U44471 ( .A(reg_i_2[10]), .X(n47940) );
  inv_x1_sg U44472 ( .A(reg_i_2[9]), .X(n47938) );
  inv_x1_sg U44473 ( .A(reg_i_2[8]), .X(n47936) );
  inv_x1_sg U44474 ( .A(reg_i_2[7]), .X(n47934) );
  inv_x1_sg U44475 ( .A(reg_i_2[6]), .X(n47932) );
  inv_x1_sg U44476 ( .A(reg_i_2[5]), .X(n47930) );
  inv_x1_sg U44477 ( .A(reg_i_2[4]), .X(n47928) );
  inv_x1_sg U44478 ( .A(reg_i_2[3]), .X(n47926) );
  inv_x1_sg U44479 ( .A(reg_i_2[2]), .X(n47924) );
  inv_x1_sg U44480 ( .A(reg_i_2[1]), .X(n47922) );
  inv_x1_sg U44481 ( .A(reg_i_2[0]), .X(n47920) );
  inv_x1_sg U44482 ( .A(reg_i_1[19]), .X(n47918) );
  inv_x1_sg U44483 ( .A(reg_i_1[18]), .X(n47916) );
  inv_x1_sg U44484 ( .A(reg_i_1[17]), .X(n47914) );
  inv_x1_sg U44485 ( .A(reg_i_1[16]), .X(n47912) );
  inv_x1_sg U44486 ( .A(reg_i_1[15]), .X(n47910) );
  inv_x1_sg U44487 ( .A(reg_i_1[14]), .X(n47908) );
  inv_x1_sg U44488 ( .A(reg_i_1[13]), .X(n47906) );
  inv_x1_sg U44489 ( .A(reg_i_1[12]), .X(n47904) );
  inv_x1_sg U44490 ( .A(reg_i_1[11]), .X(n47902) );
  inv_x1_sg U44491 ( .A(reg_i_1[10]), .X(n47900) );
  inv_x1_sg U44492 ( .A(reg_i_1[9]), .X(n47898) );
  inv_x1_sg U44493 ( .A(reg_i_1[8]), .X(n47896) );
  inv_x1_sg U44494 ( .A(reg_i_1[7]), .X(n47894) );
  inv_x1_sg U44495 ( .A(reg_i_1[6]), .X(n47892) );
  inv_x1_sg U44496 ( .A(reg_i_1[5]), .X(n47890) );
  inv_x1_sg U44497 ( .A(reg_i_1[4]), .X(n47888) );
  inv_x1_sg U44498 ( .A(reg_i_1[3]), .X(n47886) );
  inv_x1_sg U44499 ( .A(reg_i_1[2]), .X(n47884) );
  inv_x1_sg U44500 ( .A(reg_i_1[1]), .X(n47882) );
  inv_x1_sg U44501 ( .A(reg_i_1[0]), .X(n47880) );
  inv_x1_sg U44502 ( .A(reg_i_0[19]), .X(n47878) );
  inv_x1_sg U44503 ( .A(reg_i_0[18]), .X(n47876) );
  inv_x1_sg U44504 ( .A(reg_i_0[17]), .X(n47874) );
  inv_x1_sg U44505 ( .A(reg_i_0[16]), .X(n47872) );
  inv_x1_sg U44506 ( .A(reg_i_0[15]), .X(n47870) );
  inv_x1_sg U44507 ( .A(reg_i_0[14]), .X(n47868) );
  inv_x1_sg U44508 ( .A(reg_i_0[13]), .X(n47866) );
  inv_x1_sg U44509 ( .A(reg_i_0[12]), .X(n47864) );
  inv_x1_sg U44510 ( .A(reg_i_0[11]), .X(n47862) );
  inv_x1_sg U44511 ( .A(reg_i_0[10]), .X(n47860) );
  inv_x1_sg U44512 ( .A(reg_i_0[9]), .X(n47858) );
  inv_x1_sg U44513 ( .A(reg_i_0[8]), .X(n47856) );
  inv_x1_sg U44514 ( .A(reg_i_0[7]), .X(n47854) );
  inv_x1_sg U44515 ( .A(reg_i_0[6]), .X(n47852) );
  inv_x1_sg U44516 ( .A(reg_i_0[5]), .X(n47850) );
  inv_x1_sg U44517 ( .A(reg_i_0[4]), .X(n47848) );
  inv_x1_sg U44518 ( .A(reg_i_0[3]), .X(n47846) );
  inv_x1_sg U44519 ( .A(reg_i_0[2]), .X(n47844) );
  inv_x1_sg U44520 ( .A(reg_i_0[1]), .X(n47842) );
  inv_x1_sg U44521 ( .A(reg_i_0[0]), .X(n47840) );
  inv_x1_sg U44522 ( .A(reg_i_mask[0]), .X(n47838) );
  inv_x1_sg U44523 ( .A(reg_i_mask[1]), .X(n51622) );
  inv_x1_sg U44524 ( .A(reg_i_mask[2]), .X(n51620) );
  inv_x1_sg U44525 ( .A(reg_i_mask[3]), .X(n51618) );
  inv_x1_sg U44526 ( .A(reg_i_mask[4]), .X(n47836) );
  inv_x1_sg U44527 ( .A(reg_i_mask[5]), .X(n47834) );
  inv_x1_sg U44528 ( .A(reg_i_mask[6]), .X(n51616) );
  inv_x1_sg U44529 ( .A(reg_i_mask[7]), .X(n51614) );
  inv_x1_sg U44530 ( .A(reg_i_mask[8]), .X(n51612) );
  inv_x1_sg U44531 ( .A(reg_i_mask[9]), .X(n51610) );
  inv_x1_sg U44532 ( .A(reg_i_mask[10]), .X(n51608) );
  inv_x1_sg U44533 ( .A(reg_i_mask[11]), .X(n51606) );
  inv_x1_sg U44534 ( .A(reg_i_mask[12]), .X(n51604) );
  inv_x1_sg U44535 ( .A(reg_i_mask[13]), .X(n51602) );
  inv_x1_sg U44536 ( .A(reg_i_mask[14]), .X(n51600) );
  inv_x1_sg U44537 ( .A(reg_i_mask[15]), .X(n51598) );
  inv_x1_sg U44538 ( .A(reg_i_mask[16]), .X(n51596) );
  inv_x1_sg U44539 ( .A(reg_i_mask[17]), .X(n47832) );
  inv_x1_sg U44540 ( .A(reg_i_mask[18]), .X(n51594) );
  inv_x1_sg U44541 ( .A(reg_i_mask[19]), .X(n51592) );
  inv_x1_sg U44542 ( .A(reg_i_mask[20]), .X(n51590) );
  inv_x1_sg U44543 ( .A(reg_i_mask[21]), .X(n51588) );
  inv_x1_sg U44544 ( .A(reg_i_mask[22]), .X(n51586) );
  inv_x1_sg U44545 ( .A(reg_i_mask[23]), .X(n51584) );
  inv_x1_sg U44546 ( .A(reg_i_mask[24]), .X(n51582) );
  inv_x1_sg U44547 ( .A(reg_i_mask[25]), .X(n51580) );
  inv_x1_sg U44548 ( .A(reg_i_mask[26]), .X(n51578) );
  inv_x1_sg U44549 ( .A(reg_i_mask[27]), .X(n51576) );
  inv_x1_sg U44550 ( .A(reg_i_mask[28]), .X(n47830) );
  inv_x1_sg U44551 ( .A(reg_i_mask[29]), .X(n47828) );
  inv_x1_sg U44552 ( .A(reg_i_mask[30]), .X(n47826) );
  inv_x1_sg U44553 ( .A(reg_i_mask[31]), .X(n47824) );
  inv_x1_sg U44554 ( .A(reg_w_mask[0]), .X(n51574) );
  inv_x1_sg U44555 ( .A(reg_w_mask[1]), .X(n47822) );
  inv_x1_sg U44556 ( .A(reg_w_mask[2]), .X(n47820) );
  inv_x1_sg U44557 ( .A(reg_w_mask[3]), .X(n47818) );
  inv_x1_sg U44558 ( .A(reg_w_mask[4]), .X(n51572) );
  inv_x1_sg U44559 ( .A(reg_w_mask[5]), .X(n51570) );
  inv_x1_sg U44560 ( .A(reg_w_mask[6]), .X(n47816) );
  inv_x1_sg U44561 ( .A(reg_w_mask[7]), .X(n47814) );
  inv_x1_sg U44562 ( .A(reg_w_mask[8]), .X(n47812) );
  inv_x1_sg U44563 ( .A(reg_w_mask[9]), .X(n47810) );
  inv_x1_sg U44564 ( .A(reg_w_mask[10]), .X(n47808) );
  inv_x1_sg U44565 ( .A(reg_w_mask[11]), .X(n47806) );
  inv_x1_sg U44566 ( .A(reg_w_mask[12]), .X(n47804) );
  inv_x1_sg U44567 ( .A(reg_w_mask[13]), .X(n47802) );
  inv_x1_sg U44568 ( .A(reg_w_mask[14]), .X(n47800) );
  inv_x1_sg U44569 ( .A(reg_w_mask[15]), .X(n47798) );
  inv_x1_sg U44570 ( .A(reg_w_mask[16]), .X(n47796) );
  inv_x1_sg U44571 ( .A(reg_w_mask[17]), .X(n51568) );
  inv_x1_sg U44572 ( .A(reg_w_mask[18]), .X(n47794) );
  inv_x1_sg U44573 ( .A(reg_w_mask[19]), .X(n47792) );
  inv_x1_sg U44574 ( .A(reg_w_mask[20]), .X(n47790) );
  inv_x1_sg U44575 ( .A(reg_w_mask[21]), .X(n47788) );
  inv_x1_sg U44576 ( .A(reg_w_mask[22]), .X(n47786) );
  inv_x1_sg U44577 ( .A(reg_w_mask[23]), .X(n47784) );
  inv_x1_sg U44578 ( .A(reg_w_mask[24]), .X(n47782) );
  inv_x1_sg U44579 ( .A(reg_w_mask[25]), .X(n47780) );
  inv_x1_sg U44580 ( .A(reg_w_mask[26]), .X(n47778) );
  inv_x1_sg U44581 ( .A(reg_w_mask[27]), .X(n47776) );
  inv_x1_sg U44582 ( .A(reg_w_mask[28]), .X(n51566) );
  inv_x1_sg U44583 ( .A(reg_w_mask[29]), .X(n51564) );
  inv_x1_sg U44584 ( .A(reg_w_mask[30]), .X(n51562) );
  inv_x1_sg U44585 ( .A(reg_w_mask[31]), .X(n51560) );
  nand_x1_sg U44586 ( .A(n39836), .B(input_ready), .X(n39835) );
  inv_x1_sg U44587 ( .A(n69266), .X(n51558) );
  inv_x1_sg U44588 ( .A(n69231), .X(n54996) );
  inv_x1_sg U44589 ( .A(n69230), .X(n54958) );
  inv_x1_sg U44590 ( .A(n69229), .X(n54960) );
  inv_x1_sg U44591 ( .A(n69228), .X(n54962) );
  inv_x1_sg U44592 ( .A(n69227), .X(n54964) );
  inv_x1_sg U44593 ( .A(n69226), .X(n54966) );
  inv_x1_sg U44594 ( .A(n69225), .X(n54968) );
  inv_x1_sg U44595 ( .A(n69224), .X(n54970) );
  inv_x1_sg U44596 ( .A(n69223), .X(n54972) );
  inv_x1_sg U44597 ( .A(n69222), .X(n54974) );
  inv_x1_sg U44598 ( .A(n69221), .X(n54976) );
  inv_x1_sg U44599 ( .A(n69220), .X(n54978) );
  inv_x1_sg U44600 ( .A(n69219), .X(n54980) );
  inv_x1_sg U44601 ( .A(n69218), .X(n54982) );
  inv_x1_sg U44602 ( .A(n69217), .X(n54984) );
  inv_x1_sg U44603 ( .A(n69216), .X(n54986) );
  inv_x1_sg U44604 ( .A(n69215), .X(n54988) );
  inv_x1_sg U44605 ( .A(n69214), .X(n54990) );
  inv_x1_sg U44606 ( .A(n69213), .X(n54992) );
  inv_x1_sg U44607 ( .A(n69212), .X(n54994) );
  inv_x1_sg U44608 ( .A(n69211), .X(n53718) );
  inv_x1_sg U44609 ( .A(n69210), .X(n53720) );
  inv_x1_sg U44610 ( .A(n69209), .X(n53722) );
  inv_x1_sg U44611 ( .A(n69208), .X(n53724) );
  inv_x1_sg U44612 ( .A(n69207), .X(n53726) );
  inv_x1_sg U44613 ( .A(n69206), .X(n53728) );
  inv_x1_sg U44614 ( .A(n69205), .X(n53730) );
  inv_x1_sg U44615 ( .A(n69204), .X(n53732) );
  inv_x1_sg U44616 ( .A(n69203), .X(n53734) );
  inv_x1_sg U44617 ( .A(n69202), .X(n53736) );
  inv_x1_sg U44618 ( .A(n69201), .X(n53738) );
  inv_x1_sg U44619 ( .A(n69200), .X(n53740) );
  inv_x1_sg U44620 ( .A(n69199), .X(n53742) );
  inv_x1_sg U44621 ( .A(n69198), .X(n53744) );
  inv_x1_sg U44622 ( .A(n69197), .X(n53746) );
  inv_x1_sg U44623 ( .A(n69196), .X(n53748) );
  inv_x1_sg U44624 ( .A(n69195), .X(n53750) );
  inv_x1_sg U44625 ( .A(n69194), .X(n53752) );
  inv_x1_sg U44626 ( .A(n69193), .X(n53754) );
  inv_x1_sg U44627 ( .A(n69192), .X(n53756) );
  inv_x1_sg U44628 ( .A(n69191), .X(n53758) );
  inv_x1_sg U44629 ( .A(n69190), .X(n53760) );
  inv_x1_sg U44630 ( .A(n69189), .X(n53762) );
  inv_x1_sg U44631 ( .A(n69188), .X(n53764) );
  inv_x1_sg U44632 ( .A(n69187), .X(n53766) );
  inv_x1_sg U44633 ( .A(n69186), .X(n53768) );
  inv_x1_sg U44634 ( .A(n69185), .X(n53770) );
  inv_x1_sg U44635 ( .A(n69184), .X(n53772) );
  inv_x1_sg U44636 ( .A(n69183), .X(n53774) );
  inv_x1_sg U44637 ( .A(n69182), .X(n53776) );
  inv_x1_sg U44638 ( .A(n69181), .X(n53778) );
  inv_x1_sg U44639 ( .A(n69180), .X(n53780) );
  inv_x1_sg U44640 ( .A(n69179), .X(n53782) );
  inv_x1_sg U44641 ( .A(n69178), .X(n53784) );
  inv_x1_sg U44642 ( .A(n69177), .X(n53786) );
  inv_x1_sg U44643 ( .A(n69176), .X(n53788) );
  inv_x1_sg U44644 ( .A(n69175), .X(n53790) );
  inv_x1_sg U44645 ( .A(n69174), .X(n53792) );
  inv_x1_sg U44646 ( .A(n69173), .X(n53794) );
  inv_x1_sg U44647 ( .A(n69172), .X(n53796) );
  inv_x1_sg U44648 ( .A(n69171), .X(n53798) );
  inv_x1_sg U44649 ( .A(n69170), .X(n53800) );
  inv_x1_sg U44650 ( .A(n69169), .X(n53802) );
  inv_x1_sg U44651 ( .A(n69168), .X(n53804) );
  inv_x1_sg U44652 ( .A(n69167), .X(n53806) );
  inv_x1_sg U44653 ( .A(n69166), .X(n53808) );
  inv_x1_sg U44654 ( .A(n69165), .X(n53810) );
  inv_x1_sg U44655 ( .A(n69164), .X(n53812) );
  inv_x1_sg U44656 ( .A(n69163), .X(n53814) );
  inv_x1_sg U44657 ( .A(n69162), .X(n53816) );
  inv_x1_sg U44658 ( .A(n69161), .X(n53818) );
  inv_x1_sg U44659 ( .A(n69160), .X(n53820) );
  inv_x1_sg U44660 ( .A(n69159), .X(n53822) );
  inv_x1_sg U44661 ( .A(n69158), .X(n53824) );
  inv_x1_sg U44662 ( .A(n69157), .X(n53826) );
  inv_x1_sg U44663 ( .A(n69156), .X(n53828) );
  inv_x1_sg U44664 ( .A(n69155), .X(n53830) );
  inv_x1_sg U44665 ( .A(n69154), .X(n53832) );
  inv_x1_sg U44666 ( .A(n69153), .X(n53834) );
  inv_x1_sg U44667 ( .A(n69152), .X(n53836) );
  inv_x1_sg U44668 ( .A(n69151), .X(n53838) );
  inv_x1_sg U44669 ( .A(n69150), .X(n53840) );
  inv_x1_sg U44670 ( .A(n69149), .X(n53842) );
  inv_x1_sg U44671 ( .A(n69148), .X(n53844) );
  inv_x1_sg U44672 ( .A(n69147), .X(n53846) );
  inv_x1_sg U44673 ( .A(n69146), .X(n53848) );
  inv_x1_sg U44674 ( .A(n69145), .X(n53850) );
  inv_x1_sg U44675 ( .A(n69144), .X(n53852) );
  inv_x1_sg U44676 ( .A(n69143), .X(n53854) );
  inv_x1_sg U44677 ( .A(n69142), .X(n53856) );
  inv_x1_sg U44678 ( .A(n69141), .X(n53858) );
  inv_x1_sg U44679 ( .A(n69140), .X(n53860) );
  inv_x1_sg U44680 ( .A(n69139), .X(n53862) );
  inv_x1_sg U44681 ( .A(n69138), .X(n53864) );
  inv_x1_sg U44682 ( .A(n69137), .X(n53866) );
  inv_x1_sg U44683 ( .A(n69136), .X(n53868) );
  inv_x1_sg U44684 ( .A(n69135), .X(n53870) );
  inv_x1_sg U44685 ( .A(n69134), .X(n53872) );
  inv_x1_sg U44686 ( .A(n69133), .X(n53874) );
  inv_x1_sg U44687 ( .A(n69132), .X(n53876) );
  inv_x1_sg U44688 ( .A(n69131), .X(n53878) );
  inv_x1_sg U44689 ( .A(n69130), .X(n53880) );
  inv_x1_sg U44690 ( .A(n69129), .X(n53882) );
  inv_x1_sg U44691 ( .A(n69128), .X(n53884) );
  inv_x1_sg U44692 ( .A(n69127), .X(n53886) );
  inv_x1_sg U44693 ( .A(n69126), .X(n53888) );
  inv_x1_sg U44694 ( .A(n69125), .X(n53890) );
  inv_x1_sg U44695 ( .A(n69124), .X(n53892) );
  inv_x1_sg U44696 ( .A(n69123), .X(n53894) );
  inv_x1_sg U44697 ( .A(n69122), .X(n53896) );
  inv_x1_sg U44698 ( .A(n69121), .X(n53898) );
  inv_x1_sg U44699 ( .A(n69120), .X(n53900) );
  inv_x1_sg U44700 ( .A(n69119), .X(n53902) );
  inv_x1_sg U44701 ( .A(n69118), .X(n53904) );
  inv_x1_sg U44702 ( .A(n69117), .X(n53906) );
  inv_x1_sg U44703 ( .A(n69116), .X(n53908) );
  inv_x1_sg U44704 ( .A(n69115), .X(n53910) );
  inv_x1_sg U44705 ( .A(n69114), .X(n53912) );
  inv_x1_sg U44706 ( .A(n69113), .X(n53914) );
  inv_x1_sg U44707 ( .A(n69112), .X(n53916) );
  inv_x1_sg U44708 ( .A(n69111), .X(n53918) );
  inv_x1_sg U44709 ( .A(n69110), .X(n53920) );
  inv_x1_sg U44710 ( .A(n69109), .X(n53922) );
  inv_x1_sg U44711 ( .A(n69108), .X(n53924) );
  inv_x1_sg U44712 ( .A(n69107), .X(n53926) );
  inv_x1_sg U44713 ( .A(n69106), .X(n53928) );
  inv_x1_sg U44714 ( .A(n69105), .X(n53930) );
  inv_x1_sg U44715 ( .A(n69104), .X(n53932) );
  inv_x1_sg U44716 ( .A(n69103), .X(n53934) );
  inv_x1_sg U44717 ( .A(n69102), .X(n53936) );
  inv_x1_sg U44718 ( .A(n69101), .X(n53938) );
  inv_x1_sg U44719 ( .A(n69100), .X(n53940) );
  inv_x1_sg U44720 ( .A(n69099), .X(n53942) );
  inv_x1_sg U44721 ( .A(n69098), .X(n53944) );
  inv_x1_sg U44722 ( .A(n69097), .X(n53946) );
  inv_x1_sg U44723 ( .A(n69096), .X(n53948) );
  inv_x1_sg U44724 ( .A(n69095), .X(n53950) );
  inv_x1_sg U44725 ( .A(n69094), .X(n53952) );
  inv_x1_sg U44726 ( .A(n69093), .X(n53954) );
  inv_x1_sg U44727 ( .A(n69092), .X(n53956) );
  inv_x1_sg U44728 ( .A(n69091), .X(n53958) );
  inv_x1_sg U44729 ( .A(n69090), .X(n53960) );
  inv_x1_sg U44730 ( .A(n69089), .X(n53962) );
  inv_x1_sg U44731 ( .A(n69088), .X(n53964) );
  inv_x1_sg U44732 ( .A(n69087), .X(n53966) );
  inv_x1_sg U44733 ( .A(n69086), .X(n53968) );
  inv_x1_sg U44734 ( .A(n69085), .X(n53970) );
  inv_x1_sg U44735 ( .A(n69084), .X(n53972) );
  inv_x1_sg U44736 ( .A(n69083), .X(n53974) );
  inv_x1_sg U44737 ( .A(n69082), .X(n53976) );
  inv_x1_sg U44738 ( .A(n69081), .X(n53978) );
  inv_x1_sg U44739 ( .A(n69080), .X(n53980) );
  inv_x1_sg U44740 ( .A(n69079), .X(n53982) );
  inv_x1_sg U44741 ( .A(n69078), .X(n53984) );
  inv_x1_sg U44742 ( .A(n69077), .X(n53986) );
  inv_x1_sg U44743 ( .A(n69076), .X(n53988) );
  inv_x1_sg U44744 ( .A(n69075), .X(n53990) );
  inv_x1_sg U44745 ( .A(n69074), .X(n53992) );
  inv_x1_sg U44746 ( .A(n69073), .X(n53994) );
  inv_x1_sg U44747 ( .A(n69072), .X(n53996) );
  inv_x1_sg U44748 ( .A(n69071), .X(n53998) );
  inv_x1_sg U44749 ( .A(n69070), .X(n54000) );
  inv_x1_sg U44750 ( .A(n69069), .X(n54002) );
  inv_x1_sg U44751 ( .A(n69068), .X(n54004) );
  inv_x1_sg U44752 ( .A(n69067), .X(n54006) );
  inv_x1_sg U44753 ( .A(n69066), .X(n54008) );
  inv_x1_sg U44754 ( .A(n69065), .X(n54010) );
  inv_x1_sg U44755 ( .A(n69064), .X(n54012) );
  inv_x1_sg U44756 ( .A(n69063), .X(n54014) );
  inv_x1_sg U44757 ( .A(n69062), .X(n54016) );
  inv_x1_sg U44758 ( .A(n69061), .X(n54018) );
  inv_x1_sg U44759 ( .A(n69060), .X(n54020) );
  inv_x1_sg U44760 ( .A(n69059), .X(n54022) );
  inv_x1_sg U44761 ( .A(n69058), .X(n54024) );
  inv_x1_sg U44762 ( .A(n69057), .X(n54026) );
  inv_x1_sg U44763 ( .A(n69056), .X(n54028) );
  inv_x1_sg U44764 ( .A(n69055), .X(n54030) );
  inv_x1_sg U44765 ( .A(n69054), .X(n54032) );
  inv_x1_sg U44766 ( .A(n69053), .X(n54034) );
  inv_x1_sg U44767 ( .A(n69052), .X(n54036) );
  inv_x1_sg U44768 ( .A(n69051), .X(n54038) );
  inv_x1_sg U44769 ( .A(n69050), .X(n54040) );
  inv_x1_sg U44770 ( .A(n69049), .X(n54042) );
  inv_x1_sg U44771 ( .A(n69048), .X(n54044) );
  inv_x1_sg U44772 ( .A(n69047), .X(n54046) );
  inv_x1_sg U44773 ( .A(n69046), .X(n54048) );
  inv_x1_sg U44774 ( .A(n69045), .X(n54050) );
  inv_x1_sg U44775 ( .A(n69044), .X(n54052) );
  inv_x1_sg U44776 ( .A(n69043), .X(n54054) );
  inv_x1_sg U44777 ( .A(n69042), .X(n54056) );
  inv_x1_sg U44778 ( .A(n69041), .X(n54058) );
  inv_x1_sg U44779 ( .A(n69040), .X(n54060) );
  inv_x1_sg U44780 ( .A(n69039), .X(n54062) );
  inv_x1_sg U44781 ( .A(n69038), .X(n54064) );
  inv_x1_sg U44782 ( .A(n69037), .X(n54066) );
  inv_x1_sg U44783 ( .A(n69036), .X(n54068) );
  inv_x1_sg U44784 ( .A(n69035), .X(n54070) );
  inv_x1_sg U44785 ( .A(n69034), .X(n54072) );
  inv_x1_sg U44786 ( .A(n69033), .X(n54074) );
  inv_x1_sg U44787 ( .A(n69032), .X(n54076) );
  inv_x1_sg U44788 ( .A(n69031), .X(n54078) );
  inv_x1_sg U44789 ( .A(n69030), .X(n54080) );
  inv_x1_sg U44790 ( .A(n69029), .X(n54082) );
  inv_x1_sg U44791 ( .A(n69028), .X(n54084) );
  inv_x1_sg U44792 ( .A(n69027), .X(n54086) );
  inv_x1_sg U44793 ( .A(n69026), .X(n54088) );
  inv_x1_sg U44794 ( .A(n69025), .X(n54090) );
  inv_x1_sg U44795 ( .A(n69024), .X(n54092) );
  inv_x1_sg U44796 ( .A(n69023), .X(n54094) );
  inv_x1_sg U44797 ( .A(n69022), .X(n54096) );
  inv_x1_sg U44798 ( .A(n69021), .X(n54098) );
  inv_x1_sg U44799 ( .A(n69020), .X(n54100) );
  inv_x1_sg U44800 ( .A(n69019), .X(n54102) );
  inv_x1_sg U44801 ( .A(n69018), .X(n54104) );
  inv_x1_sg U44802 ( .A(n69017), .X(n54106) );
  inv_x1_sg U44803 ( .A(n69016), .X(n54108) );
  inv_x1_sg U44804 ( .A(n69015), .X(n54110) );
  inv_x1_sg U44805 ( .A(n69014), .X(n54112) );
  inv_x1_sg U44806 ( .A(n69013), .X(n54114) );
  inv_x1_sg U44807 ( .A(n69012), .X(n54116) );
  inv_x1_sg U44808 ( .A(n69011), .X(n54118) );
  inv_x1_sg U44809 ( .A(n69010), .X(n54120) );
  inv_x1_sg U44810 ( .A(n69009), .X(n54122) );
  inv_x1_sg U44811 ( .A(n69008), .X(n54124) );
  inv_x1_sg U44812 ( .A(n69007), .X(n54126) );
  inv_x1_sg U44813 ( .A(n69006), .X(n54128) );
  inv_x1_sg U44814 ( .A(n69005), .X(n54130) );
  inv_x1_sg U44815 ( .A(n69004), .X(n54132) );
  inv_x1_sg U44816 ( .A(n69003), .X(n54134) );
  inv_x1_sg U44817 ( .A(n69002), .X(n54136) );
  inv_x1_sg U44818 ( .A(n69001), .X(n54138) );
  inv_x1_sg U44819 ( .A(n69000), .X(n54140) );
  inv_x1_sg U44820 ( .A(n68999), .X(n54142) );
  inv_x1_sg U44821 ( .A(n68998), .X(n54144) );
  inv_x1_sg U44822 ( .A(n68997), .X(n54146) );
  inv_x1_sg U44823 ( .A(n68996), .X(n54148) );
  inv_x1_sg U44824 ( .A(n68995), .X(n54150) );
  inv_x1_sg U44825 ( .A(n68994), .X(n54152) );
  inv_x1_sg U44826 ( .A(n68993), .X(n54154) );
  inv_x1_sg U44827 ( .A(n68992), .X(n54156) );
  inv_x1_sg U44828 ( .A(n68991), .X(n54158) );
  inv_x1_sg U44829 ( .A(n68990), .X(n54160) );
  inv_x1_sg U44830 ( .A(n68989), .X(n54162) );
  inv_x1_sg U44831 ( .A(n68988), .X(n54164) );
  inv_x1_sg U44832 ( .A(n68987), .X(n54166) );
  inv_x1_sg U44833 ( .A(n68986), .X(n54168) );
  inv_x1_sg U44834 ( .A(n68985), .X(n54170) );
  inv_x1_sg U44835 ( .A(n68984), .X(n54172) );
  inv_x1_sg U44836 ( .A(n68983), .X(n54174) );
  inv_x1_sg U44837 ( .A(n68982), .X(n54176) );
  inv_x1_sg U44838 ( .A(n68981), .X(n54178) );
  inv_x1_sg U44839 ( .A(n68980), .X(n54180) );
  inv_x1_sg U44840 ( .A(n68979), .X(n54182) );
  inv_x1_sg U44841 ( .A(n68978), .X(n54184) );
  inv_x1_sg U44842 ( .A(n68977), .X(n54186) );
  inv_x1_sg U44843 ( .A(n68976), .X(n54188) );
  inv_x1_sg U44844 ( .A(n68975), .X(n54190) );
  inv_x1_sg U44845 ( .A(n68974), .X(n54192) );
  inv_x1_sg U44846 ( .A(n68973), .X(n54194) );
  inv_x1_sg U44847 ( .A(n68972), .X(n54196) );
  inv_x1_sg U44848 ( .A(n68971), .X(n54198) );
  inv_x1_sg U44849 ( .A(n68970), .X(n54200) );
  inv_x1_sg U44850 ( .A(n68969), .X(n54202) );
  inv_x1_sg U44851 ( .A(n68968), .X(n54204) );
  inv_x1_sg U44852 ( .A(n68967), .X(n54206) );
  inv_x1_sg U44853 ( .A(n68966), .X(n54208) );
  inv_x1_sg U44854 ( .A(n68965), .X(n54210) );
  inv_x1_sg U44855 ( .A(n68964), .X(n54212) );
  inv_x1_sg U44856 ( .A(n68963), .X(n54214) );
  inv_x1_sg U44857 ( .A(n68962), .X(n54216) );
  inv_x1_sg U44858 ( .A(n68961), .X(n54218) );
  inv_x1_sg U44859 ( .A(n68960), .X(n54220) );
  inv_x1_sg U44860 ( .A(n68959), .X(n54222) );
  inv_x1_sg U44861 ( .A(n68958), .X(n54224) );
  inv_x1_sg U44862 ( .A(n68957), .X(n54226) );
  inv_x1_sg U44863 ( .A(n68956), .X(n54228) );
  inv_x1_sg U44864 ( .A(n68955), .X(n54230) );
  inv_x1_sg U44865 ( .A(n68954), .X(n54232) );
  inv_x1_sg U44866 ( .A(n68953), .X(n54234) );
  inv_x1_sg U44867 ( .A(n68952), .X(n54236) );
  inv_x1_sg U44868 ( .A(n68951), .X(n54238) );
  inv_x1_sg U44869 ( .A(n68950), .X(n54240) );
  inv_x1_sg U44870 ( .A(n68949), .X(n54242) );
  inv_x1_sg U44871 ( .A(n68948), .X(n54244) );
  inv_x1_sg U44872 ( .A(n68947), .X(n54246) );
  inv_x1_sg U44873 ( .A(n68946), .X(n54248) );
  inv_x1_sg U44874 ( .A(n68945), .X(n54250) );
  inv_x1_sg U44875 ( .A(n68944), .X(n54252) );
  inv_x1_sg U44876 ( .A(n68943), .X(n54254) );
  inv_x1_sg U44877 ( .A(n68942), .X(n54256) );
  inv_x1_sg U44878 ( .A(n68941), .X(n54258) );
  inv_x1_sg U44879 ( .A(n68940), .X(n54260) );
  inv_x1_sg U44880 ( .A(n68939), .X(n54262) );
  inv_x1_sg U44881 ( .A(n68938), .X(n54264) );
  inv_x1_sg U44882 ( .A(n68937), .X(n54266) );
  inv_x1_sg U44883 ( .A(n68936), .X(n54268) );
  inv_x1_sg U44884 ( .A(n68935), .X(n54270) );
  inv_x1_sg U44885 ( .A(n68934), .X(n54272) );
  inv_x1_sg U44886 ( .A(n68933), .X(n54274) );
  inv_x1_sg U44887 ( .A(n68932), .X(n54276) );
  inv_x1_sg U44888 ( .A(n68931), .X(n54278) );
  inv_x1_sg U44889 ( .A(n68930), .X(n54280) );
  inv_x1_sg U44890 ( .A(n68929), .X(n54282) );
  inv_x1_sg U44891 ( .A(n68928), .X(n54284) );
  inv_x1_sg U44892 ( .A(n68927), .X(n54286) );
  inv_x1_sg U44893 ( .A(n68926), .X(n54288) );
  inv_x1_sg U44894 ( .A(n68925), .X(n54290) );
  inv_x1_sg U44895 ( .A(n68924), .X(n54292) );
  inv_x1_sg U44896 ( .A(n68923), .X(n54294) );
  inv_x1_sg U44897 ( .A(n68922), .X(n54296) );
  inv_x1_sg U44898 ( .A(n68921), .X(n54298) );
  inv_x1_sg U44899 ( .A(n68920), .X(n54300) );
  inv_x1_sg U44900 ( .A(n68919), .X(n54302) );
  inv_x1_sg U44901 ( .A(n68918), .X(n54304) );
  inv_x1_sg U44902 ( .A(n68917), .X(n54306) );
  inv_x1_sg U44903 ( .A(n68916), .X(n54308) );
  inv_x1_sg U44904 ( .A(n68915), .X(n54310) );
  inv_x1_sg U44905 ( .A(n68914), .X(n54312) );
  inv_x1_sg U44906 ( .A(n68913), .X(n54314) );
  inv_x1_sg U44907 ( .A(n68912), .X(n54316) );
  inv_x1_sg U44908 ( .A(n68911), .X(n54318) );
  inv_x1_sg U44909 ( .A(n68910), .X(n54320) );
  inv_x1_sg U44910 ( .A(n68909), .X(n54322) );
  inv_x1_sg U44911 ( .A(n68908), .X(n54324) );
  inv_x1_sg U44912 ( .A(n68907), .X(n54326) );
  inv_x1_sg U44913 ( .A(n68906), .X(n54328) );
  inv_x1_sg U44914 ( .A(n68905), .X(n54330) );
  inv_x1_sg U44915 ( .A(n68904), .X(n54332) );
  inv_x1_sg U44916 ( .A(n68903), .X(n54334) );
  inv_x1_sg U44917 ( .A(n68902), .X(n54336) );
  inv_x1_sg U44918 ( .A(n68901), .X(n54338) );
  inv_x1_sg U44919 ( .A(n68900), .X(n54340) );
  inv_x1_sg U44920 ( .A(n68899), .X(n54342) );
  inv_x1_sg U44921 ( .A(n68898), .X(n54344) );
  inv_x1_sg U44922 ( .A(n68897), .X(n54346) );
  inv_x1_sg U44923 ( .A(n68896), .X(n54348) );
  inv_x1_sg U44924 ( .A(n68895), .X(n54350) );
  inv_x1_sg U44925 ( .A(n68894), .X(n54352) );
  inv_x1_sg U44926 ( .A(n68893), .X(n54354) );
  inv_x1_sg U44927 ( .A(n68892), .X(n54356) );
  inv_x1_sg U44928 ( .A(n68891), .X(n54358) );
  inv_x1_sg U44929 ( .A(n68890), .X(n54360) );
  inv_x1_sg U44930 ( .A(n68889), .X(n54362) );
  inv_x1_sg U44931 ( .A(n68888), .X(n54364) );
  inv_x1_sg U44932 ( .A(n68887), .X(n54366) );
  inv_x1_sg U44933 ( .A(n68886), .X(n54368) );
  inv_x1_sg U44934 ( .A(n68885), .X(n54370) );
  inv_x1_sg U44935 ( .A(n68884), .X(n54372) );
  inv_x1_sg U44936 ( .A(n68883), .X(n54374) );
  inv_x1_sg U44937 ( .A(n68882), .X(n54376) );
  inv_x1_sg U44938 ( .A(n68881), .X(n54378) );
  inv_x1_sg U44939 ( .A(n68880), .X(n54380) );
  inv_x1_sg U44940 ( .A(n68879), .X(n54382) );
  inv_x1_sg U44941 ( .A(n68878), .X(n54384) );
  inv_x1_sg U44942 ( .A(n68877), .X(n54386) );
  inv_x1_sg U44943 ( .A(n68876), .X(n54388) );
  inv_x1_sg U44944 ( .A(n68875), .X(n54390) );
  inv_x1_sg U44945 ( .A(n68874), .X(n54392) );
  inv_x1_sg U44946 ( .A(n68873), .X(n54394) );
  inv_x1_sg U44947 ( .A(n68872), .X(n54396) );
  inv_x1_sg U44948 ( .A(n68871), .X(n54398) );
  inv_x1_sg U44949 ( .A(n68870), .X(n54400) );
  inv_x1_sg U44950 ( .A(n68869), .X(n54402) );
  inv_x1_sg U44951 ( .A(n68868), .X(n54404) );
  inv_x1_sg U44952 ( .A(n68867), .X(n54406) );
  inv_x1_sg U44953 ( .A(n68866), .X(n54408) );
  inv_x1_sg U44954 ( .A(n68865), .X(n54410) );
  inv_x1_sg U44955 ( .A(n68864), .X(n54412) );
  inv_x1_sg U44956 ( .A(n68863), .X(n54414) );
  inv_x1_sg U44957 ( .A(n68862), .X(n54416) );
  inv_x1_sg U44958 ( .A(n68861), .X(n54418) );
  inv_x1_sg U44959 ( .A(n68860), .X(n54420) );
  inv_x1_sg U44960 ( .A(n68859), .X(n54422) );
  inv_x1_sg U44961 ( .A(n68858), .X(n54424) );
  inv_x1_sg U44962 ( .A(n68857), .X(n54426) );
  inv_x1_sg U44963 ( .A(n68856), .X(n54428) );
  inv_x1_sg U44964 ( .A(n68855), .X(n54430) );
  inv_x1_sg U44965 ( .A(n68854), .X(n54432) );
  inv_x1_sg U44966 ( .A(n68853), .X(n54434) );
  inv_x1_sg U44967 ( .A(n68852), .X(n54436) );
  inv_x1_sg U44968 ( .A(n68851), .X(n54438) );
  inv_x1_sg U44969 ( .A(n68850), .X(n54440) );
  inv_x1_sg U44970 ( .A(n68849), .X(n54442) );
  inv_x1_sg U44971 ( .A(n68848), .X(n54444) );
  inv_x1_sg U44972 ( .A(n68847), .X(n54446) );
  inv_x1_sg U44973 ( .A(n68846), .X(n54448) );
  inv_x1_sg U44974 ( .A(n68845), .X(n54450) );
  inv_x1_sg U44975 ( .A(n68844), .X(n54452) );
  inv_x1_sg U44976 ( .A(n68843), .X(n54454) );
  inv_x1_sg U44977 ( .A(n68842), .X(n54456) );
  inv_x1_sg U44978 ( .A(n68841), .X(n54458) );
  inv_x1_sg U44979 ( .A(n68840), .X(n54460) );
  inv_x1_sg U44980 ( .A(n68839), .X(n54462) );
  inv_x1_sg U44981 ( .A(n68838), .X(n54464) );
  inv_x1_sg U44982 ( .A(n68837), .X(n54466) );
  inv_x1_sg U44983 ( .A(n68836), .X(n54468) );
  inv_x1_sg U44984 ( .A(n68835), .X(n54470) );
  inv_x1_sg U44985 ( .A(n68834), .X(n54472) );
  inv_x1_sg U44986 ( .A(n68833), .X(n54474) );
  inv_x1_sg U44987 ( .A(n68832), .X(n54476) );
  inv_x1_sg U44988 ( .A(n68831), .X(n54478) );
  inv_x1_sg U44989 ( .A(n68830), .X(n54480) );
  inv_x1_sg U44990 ( .A(n68829), .X(n54482) );
  inv_x1_sg U44991 ( .A(n68828), .X(n54484) );
  inv_x1_sg U44992 ( .A(n68827), .X(n54486) );
  inv_x1_sg U44993 ( .A(n68826), .X(n54488) );
  inv_x1_sg U44994 ( .A(n68825), .X(n54490) );
  inv_x1_sg U44995 ( .A(n68824), .X(n54492) );
  inv_x1_sg U44996 ( .A(n68823), .X(n54494) );
  inv_x1_sg U44997 ( .A(n68822), .X(n54496) );
  inv_x1_sg U44998 ( .A(n68821), .X(n54498) );
  inv_x1_sg U44999 ( .A(n68820), .X(n54500) );
  inv_x1_sg U45000 ( .A(n68819), .X(n54502) );
  inv_x1_sg U45001 ( .A(n68818), .X(n54504) );
  inv_x1_sg U45002 ( .A(n68817), .X(n54506) );
  inv_x1_sg U45003 ( .A(n68816), .X(n54508) );
  inv_x1_sg U45004 ( .A(n68815), .X(n54510) );
  inv_x1_sg U45005 ( .A(n68814), .X(n54512) );
  inv_x1_sg U45006 ( .A(n68813), .X(n54514) );
  inv_x1_sg U45007 ( .A(n68812), .X(n54516) );
  inv_x1_sg U45008 ( .A(n68811), .X(n54518) );
  inv_x1_sg U45009 ( .A(n68810), .X(n54520) );
  inv_x1_sg U45010 ( .A(n68809), .X(n54522) );
  inv_x1_sg U45011 ( .A(n68808), .X(n54524) );
  inv_x1_sg U45012 ( .A(n68807), .X(n54526) );
  inv_x1_sg U45013 ( .A(n68806), .X(n54528) );
  inv_x1_sg U45014 ( .A(n68805), .X(n54530) );
  inv_x1_sg U45015 ( .A(n68804), .X(n54532) );
  inv_x1_sg U45016 ( .A(n68803), .X(n54534) );
  inv_x1_sg U45017 ( .A(n68802), .X(n54536) );
  inv_x1_sg U45018 ( .A(n68801), .X(n54538) );
  inv_x1_sg U45019 ( .A(n68800), .X(n54540) );
  inv_x1_sg U45020 ( .A(n68799), .X(n54542) );
  inv_x1_sg U45021 ( .A(n68798), .X(n54544) );
  inv_x1_sg U45022 ( .A(n68797), .X(n54546) );
  inv_x1_sg U45023 ( .A(n68796), .X(n54548) );
  inv_x1_sg U45024 ( .A(n68795), .X(n54550) );
  inv_x1_sg U45025 ( .A(n68794), .X(n54552) );
  inv_x1_sg U45026 ( .A(n68793), .X(n54554) );
  inv_x1_sg U45027 ( .A(n68792), .X(n54556) );
  inv_x1_sg U45028 ( .A(n68791), .X(n54558) );
  inv_x1_sg U45029 ( .A(n68790), .X(n54560) );
  inv_x1_sg U45030 ( .A(n68789), .X(n54562) );
  inv_x1_sg U45031 ( .A(n68788), .X(n54564) );
  inv_x1_sg U45032 ( .A(n68787), .X(n54566) );
  inv_x1_sg U45033 ( .A(n68786), .X(n54568) );
  inv_x1_sg U45034 ( .A(n68785), .X(n54570) );
  inv_x1_sg U45035 ( .A(n68784), .X(n54572) );
  inv_x1_sg U45036 ( .A(n68783), .X(n54574) );
  inv_x1_sg U45037 ( .A(n68782), .X(n54576) );
  inv_x1_sg U45038 ( .A(n68781), .X(n54578) );
  inv_x1_sg U45039 ( .A(n68780), .X(n54580) );
  inv_x1_sg U45040 ( .A(n68779), .X(n54582) );
  inv_x1_sg U45041 ( .A(n68778), .X(n54584) );
  inv_x1_sg U45042 ( .A(n68777), .X(n54586) );
  inv_x1_sg U45043 ( .A(n68776), .X(n54588) );
  inv_x1_sg U45044 ( .A(n68775), .X(n54590) );
  inv_x1_sg U45045 ( .A(n68774), .X(n54592) );
  inv_x1_sg U45046 ( .A(n68773), .X(n54594) );
  inv_x1_sg U45047 ( .A(n68772), .X(n54596) );
  inv_x1_sg U45048 ( .A(n68771), .X(n54598) );
  inv_x1_sg U45049 ( .A(n68770), .X(n54600) );
  inv_x1_sg U45050 ( .A(n68769), .X(n54602) );
  inv_x1_sg U45051 ( .A(n68768), .X(n54604) );
  inv_x1_sg U45052 ( .A(n68767), .X(n54606) );
  inv_x1_sg U45053 ( .A(n68766), .X(n54608) );
  inv_x1_sg U45054 ( .A(n68765), .X(n54610) );
  inv_x1_sg U45055 ( .A(n68764), .X(n54612) );
  inv_x1_sg U45056 ( .A(n68763), .X(n54614) );
  inv_x1_sg U45057 ( .A(n68762), .X(n54616) );
  inv_x1_sg U45058 ( .A(n68761), .X(n54618) );
  inv_x1_sg U45059 ( .A(n68760), .X(n54620) );
  inv_x1_sg U45060 ( .A(n68759), .X(n54622) );
  inv_x1_sg U45061 ( .A(n68758), .X(n54624) );
  inv_x1_sg U45062 ( .A(n68757), .X(n54626) );
  inv_x1_sg U45063 ( .A(n68756), .X(n54628) );
  inv_x1_sg U45064 ( .A(n68755), .X(n54630) );
  inv_x1_sg U45065 ( .A(n68754), .X(n54632) );
  inv_x1_sg U45066 ( .A(n68753), .X(n54634) );
  inv_x1_sg U45067 ( .A(n68752), .X(n54636) );
  inv_x1_sg U45068 ( .A(n68751), .X(n54638) );
  inv_x1_sg U45069 ( .A(n68750), .X(n54640) );
  inv_x1_sg U45070 ( .A(n68749), .X(n54642) );
  inv_x1_sg U45071 ( .A(n68748), .X(n54644) );
  inv_x1_sg U45072 ( .A(n68747), .X(n54646) );
  inv_x1_sg U45073 ( .A(n68746), .X(n54648) );
  inv_x1_sg U45074 ( .A(n68745), .X(n54650) );
  inv_x1_sg U45075 ( .A(n68744), .X(n54652) );
  inv_x1_sg U45076 ( .A(n68743), .X(n54654) );
  inv_x1_sg U45077 ( .A(n68742), .X(n54656) );
  inv_x1_sg U45078 ( .A(n68741), .X(n54658) );
  inv_x1_sg U45079 ( .A(n68740), .X(n54660) );
  inv_x1_sg U45080 ( .A(n68739), .X(n54662) );
  inv_x1_sg U45081 ( .A(n68738), .X(n54664) );
  inv_x1_sg U45082 ( .A(n68737), .X(n54666) );
  inv_x1_sg U45083 ( .A(n68736), .X(n54668) );
  inv_x1_sg U45084 ( .A(n68735), .X(n54670) );
  inv_x1_sg U45085 ( .A(n68734), .X(n54672) );
  inv_x1_sg U45086 ( .A(n68733), .X(n54674) );
  inv_x1_sg U45087 ( .A(n68732), .X(n54676) );
  inv_x1_sg U45088 ( .A(n68731), .X(n54678) );
  inv_x1_sg U45089 ( .A(n68730), .X(n54680) );
  inv_x1_sg U45090 ( .A(n68729), .X(n54682) );
  inv_x1_sg U45091 ( .A(n68728), .X(n54684) );
  inv_x1_sg U45092 ( .A(n68727), .X(n54686) );
  inv_x1_sg U45093 ( .A(n68726), .X(n54688) );
  inv_x1_sg U45094 ( .A(n68725), .X(n54690) );
  inv_x1_sg U45095 ( .A(n68724), .X(n54692) );
  inv_x1_sg U45096 ( .A(n68723), .X(n54694) );
  inv_x1_sg U45097 ( .A(n68722), .X(n54696) );
  inv_x1_sg U45098 ( .A(n68721), .X(n54698) );
  inv_x1_sg U45099 ( .A(n68720), .X(n54700) );
  inv_x1_sg U45100 ( .A(n68719), .X(n54702) );
  inv_x1_sg U45101 ( .A(n68718), .X(n54704) );
  inv_x1_sg U45102 ( .A(n68717), .X(n54706) );
  inv_x1_sg U45103 ( .A(n68716), .X(n54708) );
  inv_x1_sg U45104 ( .A(n68715), .X(n54710) );
  inv_x1_sg U45105 ( .A(n68714), .X(n54712) );
  inv_x1_sg U45106 ( .A(n68713), .X(n54714) );
  inv_x1_sg U45107 ( .A(n68712), .X(n54716) );
  inv_x1_sg U45108 ( .A(n68711), .X(n54718) );
  inv_x1_sg U45109 ( .A(n68710), .X(n54720) );
  inv_x1_sg U45110 ( .A(n68709), .X(n54722) );
  inv_x1_sg U45111 ( .A(n68708), .X(n54724) );
  inv_x1_sg U45112 ( .A(n68707), .X(n54726) );
  inv_x1_sg U45113 ( .A(n68706), .X(n54728) );
  inv_x1_sg U45114 ( .A(n68705), .X(n54730) );
  inv_x1_sg U45115 ( .A(n68704), .X(n54732) );
  inv_x1_sg U45116 ( .A(n68703), .X(n54734) );
  inv_x1_sg U45117 ( .A(n68702), .X(n54736) );
  inv_x1_sg U45118 ( .A(n68701), .X(n54738) );
  inv_x1_sg U45119 ( .A(n68700), .X(n54740) );
  inv_x1_sg U45120 ( .A(n68699), .X(n54742) );
  inv_x1_sg U45121 ( .A(n68698), .X(n54744) );
  inv_x1_sg U45122 ( .A(n68697), .X(n54746) );
  inv_x1_sg U45123 ( .A(n68696), .X(n54748) );
  inv_x1_sg U45124 ( .A(n68695), .X(n54750) );
  inv_x1_sg U45125 ( .A(n68694), .X(n54752) );
  inv_x1_sg U45126 ( .A(n68693), .X(n54754) );
  inv_x1_sg U45127 ( .A(n68692), .X(n54756) );
  inv_x1_sg U45128 ( .A(n68691), .X(n54758) );
  inv_x1_sg U45129 ( .A(n68690), .X(n54760) );
  inv_x1_sg U45130 ( .A(n68689), .X(n54762) );
  inv_x1_sg U45131 ( .A(n68688), .X(n54764) );
  inv_x1_sg U45132 ( .A(n68687), .X(n54766) );
  inv_x1_sg U45133 ( .A(n68686), .X(n54768) );
  inv_x1_sg U45134 ( .A(n68685), .X(n54770) );
  inv_x1_sg U45135 ( .A(n68684), .X(n54772) );
  inv_x1_sg U45136 ( .A(n68683), .X(n54774) );
  inv_x1_sg U45137 ( .A(n68682), .X(n54776) );
  inv_x1_sg U45138 ( .A(n68681), .X(n54778) );
  inv_x1_sg U45139 ( .A(n68680), .X(n54780) );
  inv_x1_sg U45140 ( .A(n68679), .X(n54782) );
  inv_x1_sg U45141 ( .A(n68678), .X(n54784) );
  inv_x1_sg U45142 ( .A(n68677), .X(n54786) );
  inv_x1_sg U45143 ( .A(n68676), .X(n54788) );
  inv_x1_sg U45144 ( .A(n68675), .X(n54790) );
  inv_x1_sg U45145 ( .A(n68674), .X(n54792) );
  inv_x1_sg U45146 ( .A(n68673), .X(n54794) );
  inv_x1_sg U45147 ( .A(n68672), .X(n54796) );
  inv_x1_sg U45148 ( .A(n68671), .X(n54798) );
  inv_x1_sg U45149 ( .A(n68670), .X(n54800) );
  inv_x1_sg U45150 ( .A(n68669), .X(n54802) );
  inv_x1_sg U45151 ( .A(n68668), .X(n54804) );
  inv_x1_sg U45152 ( .A(n68667), .X(n54806) );
  inv_x1_sg U45153 ( .A(n68666), .X(n54808) );
  inv_x1_sg U45154 ( .A(n68665), .X(n54810) );
  inv_x1_sg U45155 ( .A(n68664), .X(n54812) );
  inv_x1_sg U45156 ( .A(n68663), .X(n54814) );
  inv_x1_sg U45157 ( .A(n68662), .X(n54816) );
  inv_x1_sg U45158 ( .A(n68661), .X(n54818) );
  inv_x1_sg U45159 ( .A(n68660), .X(n54820) );
  inv_x1_sg U45160 ( .A(n68659), .X(n54822) );
  inv_x1_sg U45161 ( .A(n68658), .X(n54824) );
  inv_x1_sg U45162 ( .A(n68657), .X(n54826) );
  inv_x1_sg U45163 ( .A(n68656), .X(n54828) );
  inv_x1_sg U45164 ( .A(n68655), .X(n54830) );
  inv_x1_sg U45165 ( .A(n68654), .X(n54832) );
  inv_x1_sg U45166 ( .A(n68653), .X(n54834) );
  inv_x1_sg U45167 ( .A(n68652), .X(n54836) );
  inv_x1_sg U45168 ( .A(n68651), .X(n54838) );
  inv_x1_sg U45169 ( .A(n68650), .X(n54840) );
  inv_x1_sg U45170 ( .A(n68649), .X(n54842) );
  inv_x1_sg U45171 ( .A(n68648), .X(n54844) );
  inv_x1_sg U45172 ( .A(n68647), .X(n54846) );
  inv_x1_sg U45173 ( .A(n68646), .X(n54848) );
  inv_x1_sg U45174 ( .A(n68645), .X(n54850) );
  inv_x1_sg U45175 ( .A(n68644), .X(n54852) );
  inv_x1_sg U45176 ( .A(n68643), .X(n54854) );
  inv_x1_sg U45177 ( .A(n68642), .X(n54856) );
  inv_x1_sg U45178 ( .A(n68641), .X(n54858) );
  inv_x1_sg U45179 ( .A(n68640), .X(n54860) );
  inv_x1_sg U45180 ( .A(n68639), .X(n54862) );
  inv_x1_sg U45181 ( .A(n68638), .X(n54864) );
  inv_x1_sg U45182 ( .A(n68637), .X(n54866) );
  inv_x1_sg U45183 ( .A(n68636), .X(n54868) );
  inv_x1_sg U45184 ( .A(n68635), .X(n54870) );
  inv_x1_sg U45185 ( .A(n68634), .X(n54872) );
  inv_x1_sg U45186 ( .A(n68633), .X(n54874) );
  inv_x1_sg U45187 ( .A(n68632), .X(n54876) );
  inv_x1_sg U45188 ( .A(n68631), .X(n54878) );
  inv_x1_sg U45189 ( .A(n68630), .X(n54880) );
  inv_x1_sg U45190 ( .A(n68629), .X(n54882) );
  inv_x1_sg U45191 ( .A(n68628), .X(n54884) );
  inv_x1_sg U45192 ( .A(n68627), .X(n54886) );
  inv_x1_sg U45193 ( .A(n68626), .X(n54888) );
  inv_x1_sg U45194 ( .A(n68625), .X(n54890) );
  inv_x1_sg U45195 ( .A(n68624), .X(n54892) );
  inv_x1_sg U45196 ( .A(n68623), .X(n54894) );
  inv_x1_sg U45197 ( .A(n68622), .X(n54896) );
  inv_x1_sg U45198 ( .A(n68621), .X(n54898) );
  inv_x1_sg U45199 ( .A(n68620), .X(n54900) );
  inv_x1_sg U45200 ( .A(n68619), .X(n54902) );
  inv_x1_sg U45201 ( .A(n68618), .X(n54904) );
  inv_x1_sg U45202 ( .A(n68617), .X(n54906) );
  inv_x1_sg U45203 ( .A(n68616), .X(n54908) );
  inv_x1_sg U45204 ( .A(n68615), .X(n54910) );
  inv_x1_sg U45205 ( .A(n68614), .X(n54912) );
  inv_x1_sg U45206 ( .A(n68613), .X(n54914) );
  inv_x1_sg U45207 ( .A(n68612), .X(n54916) );
  inv_x1_sg U45208 ( .A(n68611), .X(n54918) );
  inv_x1_sg U45209 ( .A(n68610), .X(n54920) );
  inv_x1_sg U45210 ( .A(n68609), .X(n54922) );
  inv_x1_sg U45211 ( .A(n68608), .X(n54924) );
  inv_x1_sg U45212 ( .A(n68607), .X(n54926) );
  inv_x1_sg U45213 ( .A(n68606), .X(n54928) );
  inv_x1_sg U45214 ( .A(n68605), .X(n54930) );
  inv_x1_sg U45215 ( .A(n68604), .X(n54932) );
  inv_x1_sg U45216 ( .A(n68603), .X(n54934) );
  inv_x1_sg U45217 ( .A(n68602), .X(n54936) );
  inv_x1_sg U45218 ( .A(n68601), .X(n54938) );
  inv_x1_sg U45219 ( .A(n68600), .X(n54940) );
  inv_x1_sg U45220 ( .A(n68599), .X(n54942) );
  inv_x1_sg U45221 ( .A(n68598), .X(n54944) );
  inv_x1_sg U45222 ( .A(n68597), .X(n54946) );
  inv_x1_sg U45223 ( .A(n68596), .X(n54948) );
  inv_x1_sg U45224 ( .A(n68595), .X(n54950) );
  inv_x1_sg U45225 ( .A(n68594), .X(n54952) );
  inv_x1_sg U45226 ( .A(n68593), .X(n54954) );
  inv_x1_sg U45227 ( .A(n68592), .X(n54956) );
  inv_x1_sg U45228 ( .A(n22652), .X(n67201) );
  nand_x1_sg U45229 ( .A(n57164), .B(n22654), .X(n22652) );
  inv_x1_sg U45230 ( .A(n22655), .X(n67200) );
  nand_x1_sg U45231 ( .A(n57163), .B(n22656), .X(n22655) );
  inv_x1_sg U45232 ( .A(n22657), .X(n67199) );
  nand_x1_sg U45233 ( .A(n22653), .B(n22658), .X(n22657) );
  inv_x1_sg U45234 ( .A(n22659), .X(n67198) );
  nand_x1_sg U45235 ( .A(n57164), .B(n22660), .X(n22659) );
  inv_x1_sg U45236 ( .A(n22661), .X(n67197) );
  nand_x1_sg U45237 ( .A(n57163), .B(n22662), .X(n22661) );
  inv_x1_sg U45238 ( .A(n22663), .X(n67196) );
  nand_x1_sg U45239 ( .A(n22653), .B(n22664), .X(n22663) );
  inv_x1_sg U45240 ( .A(n22665), .X(n67195) );
  nand_x1_sg U45241 ( .A(n57164), .B(n22666), .X(n22665) );
  inv_x1_sg U45242 ( .A(n22667), .X(n67194) );
  nand_x1_sg U45243 ( .A(n57163), .B(n22668), .X(n22667) );
  inv_x1_sg U45244 ( .A(n22669), .X(n67193) );
  nand_x1_sg U45245 ( .A(n22653), .B(n22670), .X(n22669) );
  inv_x1_sg U45246 ( .A(n22671), .X(n67192) );
  nand_x1_sg U45247 ( .A(n57164), .B(n22672), .X(n22671) );
  inv_x1_sg U45248 ( .A(n22673), .X(n67191) );
  nand_x1_sg U45249 ( .A(n57163), .B(n22674), .X(n22673) );
  inv_x1_sg U45250 ( .A(n22675), .X(n67190) );
  nand_x1_sg U45251 ( .A(n22653), .B(n22676), .X(n22675) );
  inv_x1_sg U45252 ( .A(n22677), .X(n67189) );
  nand_x1_sg U45253 ( .A(n57164), .B(n22678), .X(n22677) );
  inv_x1_sg U45254 ( .A(n22679), .X(n67188) );
  nand_x1_sg U45255 ( .A(n57163), .B(n22680), .X(n22679) );
  inv_x1_sg U45256 ( .A(n22681), .X(n67187) );
  nand_x1_sg U45257 ( .A(n22653), .B(n22682), .X(n22681) );
  inv_x1_sg U45258 ( .A(n22683), .X(n67186) );
  nand_x1_sg U45259 ( .A(n57164), .B(n22684), .X(n22683) );
  inv_x1_sg U45260 ( .A(n22685), .X(n67185) );
  nand_x1_sg U45261 ( .A(n57163), .B(n22686), .X(n22685) );
  inv_x1_sg U45262 ( .A(n22687), .X(n67184) );
  nand_x1_sg U45263 ( .A(n22653), .B(n22688), .X(n22687) );
  inv_x1_sg U45264 ( .A(n22689), .X(n67183) );
  nand_x1_sg U45265 ( .A(n57164), .B(n22690), .X(n22689) );
  inv_x1_sg U45266 ( .A(n22691), .X(n67182) );
  nand_x1_sg U45267 ( .A(n57163), .B(n22692), .X(n22691) );
  inv_x1_sg U45268 ( .A(n22699), .X(n67503) );
  nand_x1_sg U45269 ( .A(n57161), .B(n22701), .X(n22699) );
  inv_x1_sg U45270 ( .A(n22702), .X(n67504) );
  nand_x1_sg U45271 ( .A(n57160), .B(n22703), .X(n22702) );
  inv_x1_sg U45272 ( .A(n22704), .X(n67505) );
  nand_x1_sg U45273 ( .A(n22700), .B(n22705), .X(n22704) );
  inv_x1_sg U45274 ( .A(n22706), .X(n67506) );
  nand_x1_sg U45275 ( .A(n57161), .B(n22707), .X(n22706) );
  inv_x1_sg U45276 ( .A(n22708), .X(n67507) );
  nand_x1_sg U45277 ( .A(n57160), .B(n22709), .X(n22708) );
  inv_x1_sg U45278 ( .A(n22710), .X(n67508) );
  nand_x1_sg U45279 ( .A(n22700), .B(n22711), .X(n22710) );
  inv_x1_sg U45280 ( .A(n22712), .X(n67509) );
  nand_x1_sg U45281 ( .A(n57161), .B(n22713), .X(n22712) );
  inv_x1_sg U45282 ( .A(n22714), .X(n67510) );
  nand_x1_sg U45283 ( .A(n57160), .B(n22715), .X(n22714) );
  inv_x1_sg U45284 ( .A(n22716), .X(n67511) );
  nand_x1_sg U45285 ( .A(n22700), .B(n22717), .X(n22716) );
  inv_x1_sg U45286 ( .A(n22718), .X(n67512) );
  nand_x1_sg U45287 ( .A(n57161), .B(n22719), .X(n22718) );
  inv_x1_sg U45288 ( .A(n22720), .X(n67513) );
  nand_x1_sg U45289 ( .A(n57160), .B(n22721), .X(n22720) );
  inv_x1_sg U45290 ( .A(n22722), .X(n67514) );
  nand_x1_sg U45291 ( .A(n22700), .B(n22723), .X(n22722) );
  inv_x1_sg U45292 ( .A(n22724), .X(n67515) );
  nand_x1_sg U45293 ( .A(n57161), .B(n22725), .X(n22724) );
  inv_x1_sg U45294 ( .A(n22726), .X(n67516) );
  nand_x1_sg U45295 ( .A(n57160), .B(n22727), .X(n22726) );
  inv_x1_sg U45296 ( .A(n22728), .X(n67517) );
  nand_x1_sg U45297 ( .A(n22700), .B(n22729), .X(n22728) );
  inv_x1_sg U45298 ( .A(n22730), .X(n67518) );
  nand_x1_sg U45299 ( .A(n57161), .B(n22731), .X(n22730) );
  inv_x1_sg U45300 ( .A(n22732), .X(n67519) );
  nand_x1_sg U45301 ( .A(n57160), .B(n22733), .X(n22732) );
  inv_x1_sg U45302 ( .A(n22734), .X(n67520) );
  nand_x1_sg U45303 ( .A(n22700), .B(n22735), .X(n22734) );
  inv_x1_sg U45304 ( .A(n22736), .X(n67521) );
  nand_x1_sg U45305 ( .A(n57161), .B(n22737), .X(n22736) );
  inv_x1_sg U45306 ( .A(n22738), .X(n67522) );
  nand_x1_sg U45307 ( .A(n57160), .B(n22739), .X(n22738) );
  nand_x1_sg U45308 ( .A(n22747), .B(n22748), .X(\shifter_0/n11725 ) );
  nand_x1_sg U45309 ( .A(n57155), .B(n22654), .X(n22747) );
  nand_x1_sg U45310 ( .A(n22762), .B(n22763), .X(\shifter_0/n11721 ) );
  nand_x1_sg U45311 ( .A(n57155), .B(n22656), .X(n22762) );
  nand_x1_sg U45312 ( .A(n22773), .B(n22774), .X(\shifter_0/n11717 ) );
  nand_x1_sg U45313 ( .A(n57155), .B(n22658), .X(n22773) );
  nand_x1_sg U45314 ( .A(n22784), .B(n22785), .X(\shifter_0/n11713 ) );
  nand_x1_sg U45315 ( .A(n57155), .B(n22660), .X(n22784) );
  nand_x1_sg U45316 ( .A(n22795), .B(n22796), .X(\shifter_0/n11709 ) );
  nand_x1_sg U45317 ( .A(n57155), .B(n22662), .X(n22795) );
  nand_x1_sg U45318 ( .A(n22806), .B(n22807), .X(\shifter_0/n11705 ) );
  nand_x1_sg U45319 ( .A(n57155), .B(n22664), .X(n22806) );
  nand_x1_sg U45320 ( .A(n22817), .B(n22818), .X(\shifter_0/n11701 ) );
  nand_x1_sg U45321 ( .A(n57155), .B(n22666), .X(n22817) );
  nand_x1_sg U45322 ( .A(n22828), .B(n22829), .X(\shifter_0/n11697 ) );
  nand_x1_sg U45323 ( .A(n57155), .B(n22668), .X(n22828) );
  nand_x1_sg U45324 ( .A(n22839), .B(n22840), .X(\shifter_0/n11693 ) );
  nand_x1_sg U45325 ( .A(n57155), .B(n22670), .X(n22839) );
  nand_x1_sg U45326 ( .A(n22850), .B(n22851), .X(\shifter_0/n11689 ) );
  nand_x1_sg U45327 ( .A(n57155), .B(n22672), .X(n22850) );
  nand_x1_sg U45328 ( .A(n22861), .B(n22862), .X(\shifter_0/n11685 ) );
  nand_x1_sg U45329 ( .A(n57155), .B(n22674), .X(n22861) );
  nand_x1_sg U45330 ( .A(n22872), .B(n22873), .X(\shifter_0/n11681 ) );
  nand_x1_sg U45331 ( .A(n57155), .B(n22676), .X(n22872) );
  nand_x1_sg U45332 ( .A(n22883), .B(n22884), .X(\shifter_0/n11677 ) );
  nand_x1_sg U45333 ( .A(n57155), .B(n22678), .X(n22883) );
  nand_x1_sg U45334 ( .A(n22894), .B(n22895), .X(\shifter_0/n11673 ) );
  nand_x1_sg U45335 ( .A(n57155), .B(n22680), .X(n22894) );
  nand_x1_sg U45336 ( .A(n22905), .B(n22906), .X(\shifter_0/n11669 ) );
  nand_x1_sg U45337 ( .A(n57155), .B(n22682), .X(n22905) );
  nand_x1_sg U45338 ( .A(n22916), .B(n22917), .X(\shifter_0/n11665 ) );
  nand_x1_sg U45339 ( .A(n57155), .B(n22684), .X(n22916) );
  nand_x1_sg U45340 ( .A(n22927), .B(n22928), .X(\shifter_0/n11661 ) );
  nand_x1_sg U45341 ( .A(n57155), .B(n22686), .X(n22927) );
  nand_x1_sg U45342 ( .A(n22938), .B(n22939), .X(\shifter_0/n11657 ) );
  nand_x1_sg U45343 ( .A(n57155), .B(n22688), .X(n22938) );
  nand_x1_sg U45344 ( .A(n22949), .B(n22950), .X(\shifter_0/n11653 ) );
  nand_x1_sg U45345 ( .A(n57155), .B(n22690), .X(n22949) );
  nand_x1_sg U45346 ( .A(n22960), .B(n22961), .X(\shifter_0/n11649 ) );
  nand_x1_sg U45347 ( .A(n57155), .B(n22692), .X(n22960) );
  nand_x1_sg U45348 ( .A(n22975), .B(n22976), .X(\shifter_0/n11645 ) );
  nand_x1_sg U45349 ( .A(n57149), .B(n22701), .X(n22975) );
  nand_x1_sg U45350 ( .A(n22989), .B(n22990), .X(\shifter_0/n11641 ) );
  nand_x1_sg U45351 ( .A(n57149), .B(n22703), .X(n22989) );
  nand_x1_sg U45352 ( .A(n23000), .B(n23001), .X(\shifter_0/n11637 ) );
  nand_x1_sg U45353 ( .A(n57149), .B(n22705), .X(n23000) );
  nand_x1_sg U45354 ( .A(n23011), .B(n23012), .X(\shifter_0/n11633 ) );
  nand_x1_sg U45355 ( .A(n57149), .B(n22707), .X(n23011) );
  nand_x1_sg U45356 ( .A(n23022), .B(n23023), .X(\shifter_0/n11629 ) );
  nand_x1_sg U45357 ( .A(n57149), .B(n22709), .X(n23022) );
  nand_x1_sg U45358 ( .A(n23033), .B(n23034), .X(\shifter_0/n11625 ) );
  nand_x1_sg U45359 ( .A(n57149), .B(n22711), .X(n23033) );
  nand_x1_sg U45360 ( .A(n23044), .B(n23045), .X(\shifter_0/n11621 ) );
  nand_x1_sg U45361 ( .A(n57149), .B(n22713), .X(n23044) );
  nand_x1_sg U45362 ( .A(n23055), .B(n23056), .X(\shifter_0/n11617 ) );
  nand_x1_sg U45363 ( .A(n57149), .B(n22715), .X(n23055) );
  nand_x1_sg U45364 ( .A(n23066), .B(n23067), .X(\shifter_0/n11613 ) );
  nand_x1_sg U45365 ( .A(n57149), .B(n22717), .X(n23066) );
  nand_x1_sg U45366 ( .A(n23077), .B(n23078), .X(\shifter_0/n11609 ) );
  nand_x1_sg U45367 ( .A(n57149), .B(n22719), .X(n23077) );
  nand_x1_sg U45368 ( .A(n23088), .B(n23089), .X(\shifter_0/n11605 ) );
  nand_x1_sg U45369 ( .A(n57149), .B(n22721), .X(n23088) );
  nand_x1_sg U45370 ( .A(n23099), .B(n23100), .X(\shifter_0/n11601 ) );
  nand_x1_sg U45371 ( .A(n57149), .B(n22723), .X(n23099) );
  nand_x1_sg U45372 ( .A(n23110), .B(n23111), .X(\shifter_0/n11597 ) );
  nand_x1_sg U45373 ( .A(n57149), .B(n22725), .X(n23110) );
  nand_x1_sg U45374 ( .A(n23121), .B(n23122), .X(\shifter_0/n11593 ) );
  nand_x1_sg U45375 ( .A(n57149), .B(n22727), .X(n23121) );
  nand_x1_sg U45376 ( .A(n23132), .B(n23133), .X(\shifter_0/n11589 ) );
  nand_x1_sg U45377 ( .A(n57149), .B(n22729), .X(n23132) );
  nand_x1_sg U45378 ( .A(n23143), .B(n23144), .X(\shifter_0/n11585 ) );
  nand_x1_sg U45379 ( .A(n57149), .B(n22731), .X(n23143) );
  nand_x1_sg U45380 ( .A(n23154), .B(n23155), .X(\shifter_0/n11581 ) );
  nand_x1_sg U45381 ( .A(n57149), .B(n22733), .X(n23154) );
  nand_x1_sg U45382 ( .A(n23165), .B(n23166), .X(\shifter_0/n11577 ) );
  nand_x1_sg U45383 ( .A(n57149), .B(n22735), .X(n23165) );
  nand_x1_sg U45384 ( .A(n23176), .B(n23177), .X(\shifter_0/n11573 ) );
  nand_x1_sg U45385 ( .A(n57149), .B(n22737), .X(n23176) );
  nand_x1_sg U45386 ( .A(n23187), .B(n23188), .X(\shifter_0/n11569 ) );
  nand_x1_sg U45387 ( .A(n57149), .B(n22739), .X(n23187) );
  nand_x1_sg U45388 ( .A(n23202), .B(n23203), .X(\shifter_0/n11565 ) );
  nand_x1_sg U45389 ( .A(n57468), .B(n23206), .X(n23202) );
  nand_x1_sg U45390 ( .A(n23207), .B(n23208), .X(\shifter_0/n11564 ) );
  nand_x1_sg U45391 ( .A(n57464), .B(n47766), .X(n23208) );
  nand_x1_sg U45392 ( .A(n23209), .B(n23210), .X(\shifter_0/n11561 ) );
  nand_x1_sg U45393 ( .A(n57468), .B(n23211), .X(n23209) );
  nand_x1_sg U45394 ( .A(n23212), .B(n23213), .X(\shifter_0/n11560 ) );
  nand_x1_sg U45395 ( .A(n57464), .B(n47768), .X(n23213) );
  nand_x1_sg U45396 ( .A(n23214), .B(n23215), .X(\shifter_0/n11557 ) );
  nand_x1_sg U45397 ( .A(n57468), .B(n23216), .X(n23214) );
  nand_x1_sg U45398 ( .A(n23217), .B(n23218), .X(\shifter_0/n11556 ) );
  nand_x1_sg U45399 ( .A(n57464), .B(n51534), .X(n23218) );
  nand_x1_sg U45400 ( .A(n23219), .B(n23220), .X(\shifter_0/n11553 ) );
  nand_x1_sg U45401 ( .A(n57468), .B(n23221), .X(n23219) );
  nand_x1_sg U45402 ( .A(n23222), .B(n23223), .X(\shifter_0/n11552 ) );
  nand_x1_sg U45403 ( .A(n57464), .B(n56952), .X(n23223) );
  nand_x1_sg U45404 ( .A(n23224), .B(n23225), .X(\shifter_0/n11549 ) );
  nand_x1_sg U45405 ( .A(n57468), .B(n23226), .X(n23224) );
  nand_x1_sg U45406 ( .A(n23227), .B(n23228), .X(\shifter_0/n11548 ) );
  nand_x1_sg U45407 ( .A(n57464), .B(n56954), .X(n23228) );
  nand_x1_sg U45408 ( .A(n23229), .B(n23230), .X(\shifter_0/n11545 ) );
  nand_x1_sg U45409 ( .A(n57468), .B(n23231), .X(n23229) );
  nand_x1_sg U45410 ( .A(n23232), .B(n23233), .X(\shifter_0/n11544 ) );
  nand_x1_sg U45411 ( .A(n57464), .B(n47770), .X(n23233) );
  nand_x1_sg U45412 ( .A(n23234), .B(n23235), .X(\shifter_0/n11541 ) );
  nand_x1_sg U45413 ( .A(n57468), .B(n23236), .X(n23234) );
  nand_x1_sg U45414 ( .A(n23237), .B(n23238), .X(\shifter_0/n11540 ) );
  nand_x1_sg U45415 ( .A(n57464), .B(n51536), .X(n23238) );
  nand_x1_sg U45416 ( .A(n23239), .B(n23240), .X(\shifter_0/n11537 ) );
  nand_x1_sg U45417 ( .A(n57468), .B(n23241), .X(n23239) );
  nand_x1_sg U45418 ( .A(n23242), .B(n23243), .X(\shifter_0/n11536 ) );
  nand_x1_sg U45419 ( .A(n57464), .B(n57056), .X(n23243) );
  nand_x1_sg U45420 ( .A(n23244), .B(n23245), .X(\shifter_0/n11533 ) );
  nand_x1_sg U45421 ( .A(n57468), .B(n23246), .X(n23244) );
  nand_x1_sg U45422 ( .A(n23247), .B(n23248), .X(\shifter_0/n11532 ) );
  nand_x1_sg U45423 ( .A(n57464), .B(n56956), .X(n23248) );
  nand_x1_sg U45424 ( .A(n23249), .B(n23250), .X(\shifter_0/n11529 ) );
  nand_x1_sg U45425 ( .A(n57468), .B(n23251), .X(n23249) );
  nand_x1_sg U45426 ( .A(n23252), .B(n23253), .X(\shifter_0/n11528 ) );
  nand_x1_sg U45427 ( .A(n57464), .B(n56958), .X(n23253) );
  nand_x1_sg U45428 ( .A(n23254), .B(n23255), .X(\shifter_0/n11525 ) );
  nand_x1_sg U45429 ( .A(n57468), .B(n23256), .X(n23254) );
  nand_x1_sg U45430 ( .A(n23257), .B(n23258), .X(\shifter_0/n11524 ) );
  nand_x1_sg U45431 ( .A(n57464), .B(n51538), .X(n23258) );
  nand_x1_sg U45432 ( .A(n23259), .B(n23260), .X(\shifter_0/n11521 ) );
  nand_x1_sg U45433 ( .A(n57468), .B(n23261), .X(n23259) );
  nand_x1_sg U45434 ( .A(n23262), .B(n23263), .X(\shifter_0/n11520 ) );
  nand_x1_sg U45435 ( .A(n57464), .B(n57058), .X(n23263) );
  nand_x1_sg U45436 ( .A(n23264), .B(n23265), .X(\shifter_0/n11517 ) );
  nand_x1_sg U45437 ( .A(n57468), .B(n23266), .X(n23264) );
  nand_x1_sg U45438 ( .A(n23267), .B(n23268), .X(\shifter_0/n11516 ) );
  nand_x1_sg U45439 ( .A(n57464), .B(n56960), .X(n23268) );
  nand_x1_sg U45440 ( .A(n23269), .B(n23270), .X(\shifter_0/n11513 ) );
  nand_x1_sg U45441 ( .A(n57468), .B(n23271), .X(n23269) );
  nand_x1_sg U45442 ( .A(n23272), .B(n23273), .X(\shifter_0/n11512 ) );
  nand_x1_sg U45443 ( .A(n57464), .B(n56962), .X(n23273) );
  nand_x1_sg U45444 ( .A(n23274), .B(n23275), .X(\shifter_0/n11509 ) );
  nand_x1_sg U45445 ( .A(n57468), .B(n23276), .X(n23274) );
  nand_x1_sg U45446 ( .A(n23277), .B(n23278), .X(\shifter_0/n11508 ) );
  nand_x1_sg U45447 ( .A(n57464), .B(n51540), .X(n23278) );
  nand_x1_sg U45448 ( .A(n23279), .B(n23280), .X(\shifter_0/n11505 ) );
  nand_x1_sg U45449 ( .A(n57468), .B(n23281), .X(n23279) );
  nand_x1_sg U45450 ( .A(n23282), .B(n23283), .X(\shifter_0/n11504 ) );
  nand_x1_sg U45451 ( .A(n57464), .B(n57060), .X(n23283) );
  nand_x1_sg U45452 ( .A(n23284), .B(n23285), .X(\shifter_0/n11501 ) );
  nand_x1_sg U45453 ( .A(n57470), .B(n23286), .X(n23284) );
  nand_x1_sg U45454 ( .A(n23287), .B(n23288), .X(\shifter_0/n11500 ) );
  nand_x1_sg U45455 ( .A(n57466), .B(n57066), .X(n23288) );
  nand_x1_sg U45456 ( .A(n23289), .B(n23290), .X(\shifter_0/n11497 ) );
  nand_x1_sg U45457 ( .A(n57468), .B(n23291), .X(n23289) );
  nand_x1_sg U45458 ( .A(n23292), .B(n23293), .X(\shifter_0/n11496 ) );
  nand_x1_sg U45459 ( .A(n57464), .B(n56964), .X(n23293) );
  nand_x1_sg U45460 ( .A(n23294), .B(n23295), .X(\shifter_0/n11493 ) );
  nand_x1_sg U45461 ( .A(n57468), .B(n23296), .X(n23294) );
  nand_x1_sg U45462 ( .A(n23297), .B(n23298), .X(\shifter_0/n11492 ) );
  nand_x1_sg U45463 ( .A(n57464), .B(n56966), .X(n23298) );
  nand_x1_sg U45464 ( .A(n23299), .B(n23300), .X(\shifter_0/n11489 ) );
  nand_x1_sg U45465 ( .A(n57468), .B(n23301), .X(n23299) );
  nand_x1_sg U45466 ( .A(n23302), .B(n23303), .X(\shifter_0/n11488 ) );
  nand_x1_sg U45467 ( .A(n57464), .B(n57062), .X(n23303) );
  nand_x1_sg U45468 ( .A(n23310), .B(n23311), .X(\shifter_0/n11485 ) );
  nand_x1_sg U45469 ( .A(n57476), .B(n23314), .X(n23310) );
  nand_x1_sg U45470 ( .A(n23315), .B(n23316), .X(\shifter_0/n11484 ) );
  nand_x1_sg U45471 ( .A(n57472), .B(n47760), .X(n23316) );
  nand_x1_sg U45472 ( .A(n23317), .B(n23318), .X(\shifter_0/n11481 ) );
  nand_x1_sg U45473 ( .A(n57476), .B(n23319), .X(n23317) );
  nand_x1_sg U45474 ( .A(n23320), .B(n23321), .X(\shifter_0/n11480 ) );
  nand_x1_sg U45475 ( .A(n57472), .B(n47762), .X(n23321) );
  nand_x1_sg U45476 ( .A(n23322), .B(n23323), .X(\shifter_0/n11477 ) );
  nand_x1_sg U45477 ( .A(n57476), .B(n23324), .X(n23322) );
  nand_x1_sg U45478 ( .A(n23325), .B(n23326), .X(\shifter_0/n11476 ) );
  nand_x1_sg U45479 ( .A(n57472), .B(n51526), .X(n23326) );
  nand_x1_sg U45480 ( .A(n23327), .B(n23328), .X(\shifter_0/n11473 ) );
  nand_x1_sg U45481 ( .A(n57476), .B(n23329), .X(n23327) );
  nand_x1_sg U45482 ( .A(n23330), .B(n23331), .X(\shifter_0/n11472 ) );
  nand_x1_sg U45483 ( .A(n57472), .B(n56936), .X(n23331) );
  nand_x1_sg U45484 ( .A(n23332), .B(n23333), .X(\shifter_0/n11469 ) );
  nand_x1_sg U45485 ( .A(n57476), .B(n23334), .X(n23332) );
  nand_x1_sg U45486 ( .A(n23335), .B(n23336), .X(\shifter_0/n11468 ) );
  nand_x1_sg U45487 ( .A(n57472), .B(n56938), .X(n23336) );
  nand_x1_sg U45488 ( .A(n23337), .B(n23338), .X(\shifter_0/n11465 ) );
  nand_x1_sg U45489 ( .A(n57476), .B(n23339), .X(n23337) );
  nand_x1_sg U45490 ( .A(n23340), .B(n23341), .X(\shifter_0/n11464 ) );
  nand_x1_sg U45491 ( .A(n57472), .B(n47764), .X(n23341) );
  nand_x1_sg U45492 ( .A(n23342), .B(n23343), .X(\shifter_0/n11461 ) );
  nand_x1_sg U45493 ( .A(n57476), .B(n23344), .X(n23342) );
  nand_x1_sg U45494 ( .A(n23345), .B(n23346), .X(\shifter_0/n11460 ) );
  nand_x1_sg U45495 ( .A(n57472), .B(n51528), .X(n23346) );
  nand_x1_sg U45496 ( .A(n23347), .B(n23348), .X(\shifter_0/n11457 ) );
  nand_x1_sg U45497 ( .A(n57476), .B(n23349), .X(n23347) );
  nand_x1_sg U45498 ( .A(n23350), .B(n23351), .X(\shifter_0/n11456 ) );
  nand_x1_sg U45499 ( .A(n57472), .B(n57048), .X(n23351) );
  nand_x1_sg U45500 ( .A(n23352), .B(n23353), .X(\shifter_0/n11453 ) );
  nand_x1_sg U45501 ( .A(n57476), .B(n23354), .X(n23352) );
  nand_x1_sg U45502 ( .A(n23355), .B(n23356), .X(\shifter_0/n11452 ) );
  nand_x1_sg U45503 ( .A(n57472), .B(n56940), .X(n23356) );
  nand_x1_sg U45504 ( .A(n23357), .B(n23358), .X(\shifter_0/n11449 ) );
  nand_x1_sg U45505 ( .A(n57476), .B(n23359), .X(n23357) );
  nand_x1_sg U45506 ( .A(n23360), .B(n23361), .X(\shifter_0/n11448 ) );
  nand_x1_sg U45507 ( .A(n57472), .B(n56942), .X(n23361) );
  nand_x1_sg U45508 ( .A(n23362), .B(n23363), .X(\shifter_0/n11445 ) );
  nand_x1_sg U45509 ( .A(n57476), .B(n23364), .X(n23362) );
  nand_x1_sg U45510 ( .A(n23365), .B(n23366), .X(\shifter_0/n11444 ) );
  nand_x1_sg U45511 ( .A(n57472), .B(n51530), .X(n23366) );
  nand_x1_sg U45512 ( .A(n23367), .B(n23368), .X(\shifter_0/n11441 ) );
  nand_x1_sg U45513 ( .A(n57476), .B(n23369), .X(n23367) );
  nand_x1_sg U45514 ( .A(n23370), .B(n23371), .X(\shifter_0/n11440 ) );
  nand_x1_sg U45515 ( .A(n57472), .B(n57050), .X(n23371) );
  nand_x1_sg U45516 ( .A(n23372), .B(n23373), .X(\shifter_0/n11437 ) );
  nand_x1_sg U45517 ( .A(n57476), .B(n23374), .X(n23372) );
  nand_x1_sg U45518 ( .A(n23375), .B(n23376), .X(\shifter_0/n11436 ) );
  nand_x1_sg U45519 ( .A(n57472), .B(n56944), .X(n23376) );
  nand_x1_sg U45520 ( .A(n23377), .B(n23378), .X(\shifter_0/n11433 ) );
  nand_x1_sg U45521 ( .A(n57476), .B(n23379), .X(n23377) );
  nand_x1_sg U45522 ( .A(n23380), .B(n23381), .X(\shifter_0/n11432 ) );
  nand_x1_sg U45523 ( .A(n57472), .B(n56946), .X(n23381) );
  nand_x1_sg U45524 ( .A(n23382), .B(n23383), .X(\shifter_0/n11429 ) );
  nand_x1_sg U45525 ( .A(n57476), .B(n23384), .X(n23382) );
  nand_x1_sg U45526 ( .A(n23385), .B(n23386), .X(\shifter_0/n11428 ) );
  nand_x1_sg U45527 ( .A(n57472), .B(n51532), .X(n23386) );
  nand_x1_sg U45528 ( .A(n23387), .B(n23388), .X(\shifter_0/n11425 ) );
  nand_x1_sg U45529 ( .A(n57476), .B(n23389), .X(n23387) );
  nand_x1_sg U45530 ( .A(n23390), .B(n23391), .X(\shifter_0/n11424 ) );
  nand_x1_sg U45531 ( .A(n57472), .B(n57052), .X(n23391) );
  nand_x1_sg U45532 ( .A(n23392), .B(n23393), .X(\shifter_0/n11421 ) );
  nand_x1_sg U45533 ( .A(n57478), .B(n23394), .X(n23392) );
  nand_x1_sg U45534 ( .A(n23395), .B(n23396), .X(\shifter_0/n11420 ) );
  nand_x1_sg U45535 ( .A(n57474), .B(n57064), .X(n23396) );
  nand_x1_sg U45536 ( .A(n23397), .B(n23398), .X(\shifter_0/n11417 ) );
  nand_x1_sg U45537 ( .A(n57476), .B(n23399), .X(n23397) );
  nand_x1_sg U45538 ( .A(n23400), .B(n23401), .X(\shifter_0/n11416 ) );
  nand_x1_sg U45539 ( .A(n57472), .B(n56948), .X(n23401) );
  nand_x1_sg U45540 ( .A(n23402), .B(n23403), .X(\shifter_0/n11413 ) );
  nand_x1_sg U45541 ( .A(n57476), .B(n23404), .X(n23402) );
  nand_x1_sg U45542 ( .A(n23405), .B(n23406), .X(\shifter_0/n11412 ) );
  nand_x1_sg U45543 ( .A(n57472), .B(n56950), .X(n23406) );
  nand_x1_sg U45544 ( .A(n23407), .B(n23408), .X(\shifter_0/n11409 ) );
  nand_x1_sg U45545 ( .A(n57476), .B(n23409), .X(n23407) );
  nand_x1_sg U45546 ( .A(n23410), .B(n23411), .X(\shifter_0/n11408 ) );
  nand_x1_sg U45547 ( .A(n57472), .B(n57054), .X(n23411) );
  nand_x1_sg U45548 ( .A(n23942), .B(n23943), .X(\shifter_0/n11085 ) );
  nand_x1_sg U45549 ( .A(n57484), .B(n23206), .X(n23942) );
  nand_x1_sg U45550 ( .A(n57480), .B(n23945), .X(n23943) );
  nand_x1_sg U45551 ( .A(n23947), .B(n23948), .X(\shifter_0/n11084 ) );
  nand_x1_sg U45552 ( .A(n67261), .B(n57480), .X(n23948) );
  inv_x1_sg U45553 ( .A(n23945), .X(n67261) );
  nand_x1_sg U45554 ( .A(n23949), .B(n23950), .X(\shifter_0/n11081 ) );
  nand_x1_sg U45555 ( .A(n57484), .B(n23211), .X(n23949) );
  nand_x1_sg U45556 ( .A(n57480), .B(n23951), .X(n23950) );
  nand_x1_sg U45557 ( .A(n23952), .B(n23953), .X(\shifter_0/n11080 ) );
  nand_x1_sg U45558 ( .A(n67260), .B(n57480), .X(n23953) );
  inv_x1_sg U45559 ( .A(n23951), .X(n67260) );
  nand_x1_sg U45560 ( .A(n23954), .B(n23955), .X(\shifter_0/n11077 ) );
  nand_x1_sg U45561 ( .A(n57484), .B(n23216), .X(n23954) );
  nand_x1_sg U45562 ( .A(n57480), .B(n23956), .X(n23955) );
  nand_x1_sg U45563 ( .A(n23957), .B(n23958), .X(\shifter_0/n11076 ) );
  nand_x1_sg U45564 ( .A(n67259), .B(n57480), .X(n23958) );
  inv_x1_sg U45565 ( .A(n23956), .X(n67259) );
  nand_x1_sg U45566 ( .A(n23959), .B(n23960), .X(\shifter_0/n11073 ) );
  nand_x1_sg U45567 ( .A(n57484), .B(n23221), .X(n23959) );
  nand_x1_sg U45568 ( .A(n57480), .B(n23961), .X(n23960) );
  nand_x1_sg U45569 ( .A(n23962), .B(n23963), .X(\shifter_0/n11072 ) );
  nand_x1_sg U45570 ( .A(n67258), .B(n57480), .X(n23963) );
  inv_x1_sg U45571 ( .A(n23961), .X(n67258) );
  nand_x1_sg U45572 ( .A(n23964), .B(n23965), .X(\shifter_0/n11069 ) );
  nand_x1_sg U45573 ( .A(n57484), .B(n23226), .X(n23964) );
  nand_x1_sg U45574 ( .A(n57480), .B(n23966), .X(n23965) );
  nand_x1_sg U45575 ( .A(n23967), .B(n23968), .X(\shifter_0/n11068 ) );
  nand_x1_sg U45576 ( .A(n67257), .B(n57480), .X(n23968) );
  inv_x1_sg U45577 ( .A(n23966), .X(n67257) );
  nand_x1_sg U45578 ( .A(n23969), .B(n23970), .X(\shifter_0/n11065 ) );
  nand_x1_sg U45579 ( .A(n57484), .B(n23231), .X(n23969) );
  nand_x1_sg U45580 ( .A(n57480), .B(n23971), .X(n23970) );
  nand_x1_sg U45581 ( .A(n23972), .B(n23973), .X(\shifter_0/n11064 ) );
  nand_x1_sg U45582 ( .A(n67256), .B(n57480), .X(n23973) );
  inv_x1_sg U45583 ( .A(n23971), .X(n67256) );
  nand_x1_sg U45584 ( .A(n23974), .B(n23975), .X(\shifter_0/n11061 ) );
  nand_x1_sg U45585 ( .A(n57484), .B(n23236), .X(n23974) );
  nand_x1_sg U45586 ( .A(n57480), .B(n23976), .X(n23975) );
  nand_x1_sg U45587 ( .A(n23977), .B(n23978), .X(\shifter_0/n11060 ) );
  nand_x1_sg U45588 ( .A(n67255), .B(n57480), .X(n23978) );
  inv_x1_sg U45589 ( .A(n23976), .X(n67255) );
  nand_x1_sg U45590 ( .A(n23979), .B(n23980), .X(\shifter_0/n11057 ) );
  nand_x1_sg U45591 ( .A(n57484), .B(n23241), .X(n23979) );
  nand_x1_sg U45592 ( .A(n57480), .B(n23981), .X(n23980) );
  nand_x1_sg U45593 ( .A(n23982), .B(n23983), .X(\shifter_0/n11056 ) );
  nand_x1_sg U45594 ( .A(n67254), .B(n57480), .X(n23983) );
  inv_x1_sg U45595 ( .A(n23981), .X(n67254) );
  nand_x1_sg U45596 ( .A(n23984), .B(n23985), .X(\shifter_0/n11053 ) );
  nand_x1_sg U45597 ( .A(n57484), .B(n23246), .X(n23984) );
  nand_x1_sg U45598 ( .A(n57480), .B(n23986), .X(n23985) );
  nand_x1_sg U45599 ( .A(n23987), .B(n23988), .X(\shifter_0/n11052 ) );
  nand_x1_sg U45600 ( .A(n67253), .B(n57480), .X(n23988) );
  inv_x1_sg U45601 ( .A(n23986), .X(n67253) );
  nand_x1_sg U45602 ( .A(n23989), .B(n23990), .X(\shifter_0/n11049 ) );
  nand_x1_sg U45603 ( .A(n57484), .B(n23251), .X(n23989) );
  nand_x1_sg U45604 ( .A(n57480), .B(n23991), .X(n23990) );
  nand_x1_sg U45605 ( .A(n23992), .B(n23993), .X(\shifter_0/n11048 ) );
  nand_x1_sg U45606 ( .A(n67252), .B(n57480), .X(n23993) );
  inv_x1_sg U45607 ( .A(n23991), .X(n67252) );
  nand_x1_sg U45608 ( .A(n23994), .B(n23995), .X(\shifter_0/n11045 ) );
  nand_x1_sg U45609 ( .A(n57484), .B(n23256), .X(n23994) );
  nand_x1_sg U45610 ( .A(n57480), .B(n23996), .X(n23995) );
  nand_x1_sg U45611 ( .A(n23997), .B(n23998), .X(\shifter_0/n11044 ) );
  nand_x1_sg U45612 ( .A(n67251), .B(n57480), .X(n23998) );
  inv_x1_sg U45613 ( .A(n23996), .X(n67251) );
  nand_x1_sg U45614 ( .A(n23999), .B(n24000), .X(\shifter_0/n11041 ) );
  nand_x1_sg U45615 ( .A(n57484), .B(n23261), .X(n23999) );
  nand_x1_sg U45616 ( .A(n57480), .B(n24001), .X(n24000) );
  nand_x1_sg U45617 ( .A(n24002), .B(n24003), .X(\shifter_0/n11040 ) );
  nand_x1_sg U45618 ( .A(n67250), .B(n57480), .X(n24003) );
  inv_x1_sg U45619 ( .A(n24001), .X(n67250) );
  nand_x1_sg U45620 ( .A(n24004), .B(n24005), .X(\shifter_0/n11037 ) );
  nand_x1_sg U45621 ( .A(n57484), .B(n23266), .X(n24004) );
  nand_x1_sg U45622 ( .A(n57480), .B(n24006), .X(n24005) );
  nand_x1_sg U45623 ( .A(n24007), .B(n24008), .X(\shifter_0/n11036 ) );
  nand_x1_sg U45624 ( .A(n67249), .B(n57480), .X(n24008) );
  inv_x1_sg U45625 ( .A(n24006), .X(n67249) );
  nand_x1_sg U45626 ( .A(n24009), .B(n24010), .X(\shifter_0/n11033 ) );
  nand_x1_sg U45627 ( .A(n57484), .B(n23271), .X(n24009) );
  nand_x1_sg U45628 ( .A(n57480), .B(n24011), .X(n24010) );
  nand_x1_sg U45629 ( .A(n24012), .B(n24013), .X(\shifter_0/n11032 ) );
  nand_x1_sg U45630 ( .A(n67248), .B(n57480), .X(n24013) );
  inv_x1_sg U45631 ( .A(n24011), .X(n67248) );
  nand_x1_sg U45632 ( .A(n24014), .B(n24015), .X(\shifter_0/n11029 ) );
  nand_x1_sg U45633 ( .A(n57484), .B(n23276), .X(n24014) );
  nand_x1_sg U45634 ( .A(n57480), .B(n24016), .X(n24015) );
  nand_x1_sg U45635 ( .A(n24017), .B(n24018), .X(\shifter_0/n11028 ) );
  nand_x1_sg U45636 ( .A(n67247), .B(n57480), .X(n24018) );
  inv_x1_sg U45637 ( .A(n24016), .X(n67247) );
  nand_x1_sg U45638 ( .A(n24019), .B(n24020), .X(\shifter_0/n11025 ) );
  nand_x1_sg U45639 ( .A(n57484), .B(n23281), .X(n24019) );
  nand_x1_sg U45640 ( .A(n57480), .B(n24021), .X(n24020) );
  nand_x1_sg U45641 ( .A(n24022), .B(n24023), .X(\shifter_0/n11024 ) );
  nand_x1_sg U45642 ( .A(n67246), .B(n57480), .X(n24023) );
  inv_x1_sg U45643 ( .A(n24021), .X(n67246) );
  nand_x1_sg U45644 ( .A(n24024), .B(n24025), .X(\shifter_0/n11021 ) );
  nand_x1_sg U45645 ( .A(n57486), .B(n23286), .X(n24024) );
  nand_x1_sg U45646 ( .A(n57482), .B(n24026), .X(n24025) );
  nand_x1_sg U45647 ( .A(n24027), .B(n24028), .X(\shifter_0/n11020 ) );
  nand_x1_sg U45648 ( .A(n67245), .B(n57480), .X(n24028) );
  inv_x1_sg U45649 ( .A(n24026), .X(n67245) );
  nand_x1_sg U45650 ( .A(n24029), .B(n24030), .X(\shifter_0/n11017 ) );
  nand_x1_sg U45651 ( .A(n57484), .B(n23291), .X(n24029) );
  nand_x1_sg U45652 ( .A(n57480), .B(n24031), .X(n24030) );
  nand_x1_sg U45653 ( .A(n24032), .B(n24033), .X(\shifter_0/n11016 ) );
  nand_x1_sg U45654 ( .A(n67244), .B(n57480), .X(n24033) );
  inv_x1_sg U45655 ( .A(n24031), .X(n67244) );
  nand_x1_sg U45656 ( .A(n24034), .B(n24035), .X(\shifter_0/n11013 ) );
  nand_x1_sg U45657 ( .A(n57484), .B(n23296), .X(n24034) );
  nand_x1_sg U45658 ( .A(n57480), .B(n24036), .X(n24035) );
  nand_x1_sg U45659 ( .A(n24037), .B(n24038), .X(\shifter_0/n11012 ) );
  nand_x1_sg U45660 ( .A(n67243), .B(n57480), .X(n24038) );
  inv_x1_sg U45661 ( .A(n24036), .X(n67243) );
  nand_x1_sg U45662 ( .A(n24039), .B(n24040), .X(\shifter_0/n11009 ) );
  nand_x1_sg U45663 ( .A(n57484), .B(n23301), .X(n24039) );
  nand_x1_sg U45664 ( .A(n57480), .B(n24041), .X(n24040) );
  nand_x1_sg U45665 ( .A(n24042), .B(n24043), .X(\shifter_0/n11008 ) );
  nand_x1_sg U45666 ( .A(n67242), .B(n57480), .X(n24043) );
  inv_x1_sg U45667 ( .A(n24041), .X(n67242) );
  nand_x1_sg U45668 ( .A(n24052), .B(n24053), .X(\shifter_0/n11005 ) );
  nand_x1_sg U45669 ( .A(n57492), .B(n23314), .X(n24052) );
  nand_x1_sg U45670 ( .A(n57488), .B(n24055), .X(n24053) );
  nand_x1_sg U45671 ( .A(n24057), .B(n24058), .X(\shifter_0/n11004 ) );
  nand_x1_sg U45672 ( .A(n67454), .B(n57488), .X(n24058) );
  inv_x1_sg U45673 ( .A(n24055), .X(n67454) );
  nand_x1_sg U45674 ( .A(n24059), .B(n24060), .X(\shifter_0/n11001 ) );
  nand_x1_sg U45675 ( .A(n57492), .B(n23319), .X(n24059) );
  nand_x1_sg U45676 ( .A(n57488), .B(n24061), .X(n24060) );
  nand_x1_sg U45677 ( .A(n24062), .B(n24063), .X(\shifter_0/n11000 ) );
  nand_x1_sg U45678 ( .A(n67453), .B(n57488), .X(n24063) );
  inv_x1_sg U45679 ( .A(n24061), .X(n67453) );
  nand_x1_sg U45680 ( .A(n24064), .B(n24065), .X(\shifter_0/n10997 ) );
  nand_x1_sg U45681 ( .A(n57492), .B(n23324), .X(n24064) );
  nand_x1_sg U45682 ( .A(n57488), .B(n24066), .X(n24065) );
  nand_x1_sg U45683 ( .A(n24067), .B(n24068), .X(\shifter_0/n10996 ) );
  nand_x1_sg U45684 ( .A(n67452), .B(n57488), .X(n24068) );
  inv_x1_sg U45685 ( .A(n24066), .X(n67452) );
  nand_x1_sg U45686 ( .A(n24069), .B(n24070), .X(\shifter_0/n10993 ) );
  nand_x1_sg U45687 ( .A(n57492), .B(n23329), .X(n24069) );
  nand_x1_sg U45688 ( .A(n57488), .B(n24071), .X(n24070) );
  nand_x1_sg U45689 ( .A(n24072), .B(n24073), .X(\shifter_0/n10992 ) );
  nand_x1_sg U45690 ( .A(n67451), .B(n57488), .X(n24073) );
  inv_x1_sg U45691 ( .A(n24071), .X(n67451) );
  nand_x1_sg U45692 ( .A(n24074), .B(n24075), .X(\shifter_0/n10989 ) );
  nand_x1_sg U45693 ( .A(n57492), .B(n23334), .X(n24074) );
  nand_x1_sg U45694 ( .A(n57488), .B(n24076), .X(n24075) );
  nand_x1_sg U45695 ( .A(n24077), .B(n24078), .X(\shifter_0/n10988 ) );
  nand_x1_sg U45696 ( .A(n67450), .B(n57488), .X(n24078) );
  inv_x1_sg U45697 ( .A(n24076), .X(n67450) );
  nand_x1_sg U45698 ( .A(n24079), .B(n24080), .X(\shifter_0/n10985 ) );
  nand_x1_sg U45699 ( .A(n57492), .B(n23339), .X(n24079) );
  nand_x1_sg U45700 ( .A(n57488), .B(n24081), .X(n24080) );
  nand_x1_sg U45701 ( .A(n24082), .B(n24083), .X(\shifter_0/n10984 ) );
  nand_x1_sg U45702 ( .A(n67449), .B(n57488), .X(n24083) );
  inv_x1_sg U45703 ( .A(n24081), .X(n67449) );
  nand_x1_sg U45704 ( .A(n24084), .B(n24085), .X(\shifter_0/n10981 ) );
  nand_x1_sg U45705 ( .A(n57492), .B(n23344), .X(n24084) );
  nand_x1_sg U45706 ( .A(n57488), .B(n24086), .X(n24085) );
  nand_x1_sg U45707 ( .A(n24087), .B(n24088), .X(\shifter_0/n10980 ) );
  nand_x1_sg U45708 ( .A(n67448), .B(n57488), .X(n24088) );
  inv_x1_sg U45709 ( .A(n24086), .X(n67448) );
  nand_x1_sg U45710 ( .A(n24089), .B(n24090), .X(\shifter_0/n10977 ) );
  nand_x1_sg U45711 ( .A(n57492), .B(n23349), .X(n24089) );
  nand_x1_sg U45712 ( .A(n57488), .B(n24091), .X(n24090) );
  nand_x1_sg U45713 ( .A(n24092), .B(n24093), .X(\shifter_0/n10976 ) );
  nand_x1_sg U45714 ( .A(n67447), .B(n57488), .X(n24093) );
  inv_x1_sg U45715 ( .A(n24091), .X(n67447) );
  nand_x1_sg U45716 ( .A(n24094), .B(n24095), .X(\shifter_0/n10973 ) );
  nand_x1_sg U45717 ( .A(n57492), .B(n23354), .X(n24094) );
  nand_x1_sg U45718 ( .A(n57488), .B(n24096), .X(n24095) );
  nand_x1_sg U45719 ( .A(n24097), .B(n24098), .X(\shifter_0/n10972 ) );
  nand_x1_sg U45720 ( .A(n67446), .B(n57488), .X(n24098) );
  inv_x1_sg U45721 ( .A(n24096), .X(n67446) );
  nand_x1_sg U45722 ( .A(n24099), .B(n24100), .X(\shifter_0/n10969 ) );
  nand_x1_sg U45723 ( .A(n57492), .B(n23359), .X(n24099) );
  nand_x1_sg U45724 ( .A(n57488), .B(n24101), .X(n24100) );
  nand_x1_sg U45725 ( .A(n24102), .B(n24103), .X(\shifter_0/n10968 ) );
  nand_x1_sg U45726 ( .A(n67445), .B(n57488), .X(n24103) );
  inv_x1_sg U45727 ( .A(n24101), .X(n67445) );
  nand_x1_sg U45728 ( .A(n24104), .B(n24105), .X(\shifter_0/n10965 ) );
  nand_x1_sg U45729 ( .A(n57492), .B(n23364), .X(n24104) );
  nand_x1_sg U45730 ( .A(n57488), .B(n24106), .X(n24105) );
  nand_x1_sg U45731 ( .A(n24107), .B(n24108), .X(\shifter_0/n10964 ) );
  nand_x1_sg U45732 ( .A(n67444), .B(n57488), .X(n24108) );
  inv_x1_sg U45733 ( .A(n24106), .X(n67444) );
  nand_x1_sg U45734 ( .A(n24109), .B(n24110), .X(\shifter_0/n10961 ) );
  nand_x1_sg U45735 ( .A(n57492), .B(n23369), .X(n24109) );
  nand_x1_sg U45736 ( .A(n57488), .B(n24111), .X(n24110) );
  nand_x1_sg U45737 ( .A(n24112), .B(n24113), .X(\shifter_0/n10960 ) );
  nand_x1_sg U45738 ( .A(n67443), .B(n57488), .X(n24113) );
  inv_x1_sg U45739 ( .A(n24111), .X(n67443) );
  nand_x1_sg U45740 ( .A(n24114), .B(n24115), .X(\shifter_0/n10957 ) );
  nand_x1_sg U45741 ( .A(n57492), .B(n23374), .X(n24114) );
  nand_x1_sg U45742 ( .A(n57488), .B(n24116), .X(n24115) );
  nand_x1_sg U45743 ( .A(n24117), .B(n24118), .X(\shifter_0/n10956 ) );
  nand_x1_sg U45744 ( .A(n67442), .B(n57488), .X(n24118) );
  inv_x1_sg U45745 ( .A(n24116), .X(n67442) );
  nand_x1_sg U45746 ( .A(n24119), .B(n24120), .X(\shifter_0/n10953 ) );
  nand_x1_sg U45747 ( .A(n57492), .B(n23379), .X(n24119) );
  nand_x1_sg U45748 ( .A(n57488), .B(n24121), .X(n24120) );
  nand_x1_sg U45749 ( .A(n24122), .B(n24123), .X(\shifter_0/n10952 ) );
  nand_x1_sg U45750 ( .A(n67441), .B(n57488), .X(n24123) );
  inv_x1_sg U45751 ( .A(n24121), .X(n67441) );
  nand_x1_sg U45752 ( .A(n24124), .B(n24125), .X(\shifter_0/n10949 ) );
  nand_x1_sg U45753 ( .A(n57492), .B(n23384), .X(n24124) );
  nand_x1_sg U45754 ( .A(n57488), .B(n24126), .X(n24125) );
  nand_x1_sg U45755 ( .A(n24127), .B(n24128), .X(\shifter_0/n10948 ) );
  nand_x1_sg U45756 ( .A(n67440), .B(n57488), .X(n24128) );
  inv_x1_sg U45757 ( .A(n24126), .X(n67440) );
  nand_x1_sg U45758 ( .A(n24129), .B(n24130), .X(\shifter_0/n10945 ) );
  nand_x1_sg U45759 ( .A(n57492), .B(n23389), .X(n24129) );
  nand_x1_sg U45760 ( .A(n57488), .B(n24131), .X(n24130) );
  nand_x1_sg U45761 ( .A(n24132), .B(n24133), .X(\shifter_0/n10944 ) );
  nand_x1_sg U45762 ( .A(n67439), .B(n57488), .X(n24133) );
  inv_x1_sg U45763 ( .A(n24131), .X(n67439) );
  nand_x1_sg U45764 ( .A(n24134), .B(n24135), .X(\shifter_0/n10941 ) );
  nand_x1_sg U45765 ( .A(n57494), .B(n23394), .X(n24134) );
  nand_x1_sg U45766 ( .A(n57490), .B(n24136), .X(n24135) );
  nand_x1_sg U45767 ( .A(n24137), .B(n24138), .X(\shifter_0/n10940 ) );
  nand_x1_sg U45768 ( .A(n67438), .B(n57488), .X(n24138) );
  inv_x1_sg U45769 ( .A(n24136), .X(n67438) );
  nand_x1_sg U45770 ( .A(n24139), .B(n24140), .X(\shifter_0/n10937 ) );
  nand_x1_sg U45771 ( .A(n57492), .B(n23399), .X(n24139) );
  nand_x1_sg U45772 ( .A(n57488), .B(n24141), .X(n24140) );
  nand_x1_sg U45773 ( .A(n24142), .B(n24143), .X(\shifter_0/n10936 ) );
  nand_x1_sg U45774 ( .A(n67437), .B(n57488), .X(n24143) );
  inv_x1_sg U45775 ( .A(n24141), .X(n67437) );
  nand_x1_sg U45776 ( .A(n24144), .B(n24145), .X(\shifter_0/n10933 ) );
  nand_x1_sg U45777 ( .A(n57492), .B(n23404), .X(n24144) );
  nand_x1_sg U45778 ( .A(n57488), .B(n24146), .X(n24145) );
  nand_x1_sg U45779 ( .A(n24147), .B(n24148), .X(\shifter_0/n10932 ) );
  nand_x1_sg U45780 ( .A(n67436), .B(n57488), .X(n24148) );
  inv_x1_sg U45781 ( .A(n24146), .X(n67436) );
  nand_x1_sg U45782 ( .A(n24149), .B(n24150), .X(\shifter_0/n10929 ) );
  nand_x1_sg U45783 ( .A(n57492), .B(n23409), .X(n24149) );
  nand_x1_sg U45784 ( .A(n57488), .B(n24151), .X(n24150) );
  nand_x1_sg U45785 ( .A(n24152), .B(n24153), .X(\shifter_0/n10928 ) );
  nand_x1_sg U45786 ( .A(n67435), .B(n57488), .X(n24153) );
  inv_x1_sg U45787 ( .A(n24151), .X(n67435) );
  inv_x1_sg U45788 ( .A(n26039), .X(n67539) );
  nand_x1_sg U45789 ( .A(n26040), .B(n57114), .X(n26039) );
  inv_x1_sg U45790 ( .A(n26045), .X(n67538) );
  inv_x1_sg U45791 ( .A(n26048), .X(n67533) );
  nand_x1_sg U45792 ( .A(n26049), .B(n57114), .X(n26048) );
  inv_x1_sg U45793 ( .A(n26054), .X(n67531) );
  nand_x1_sg U45794 ( .A(n26053), .B(n57114), .X(n26054) );
  inv_x1_sg U45795 ( .A(n26057), .X(n67580) );
  nand_x1_sg U45796 ( .A(n26056), .B(n57114), .X(n26057) );
  inv_x1_sg U45797 ( .A(n26062), .X(n67577) );
  nand_x1_sg U45798 ( .A(n26061), .B(n57114), .X(n26062) );
  inv_x1_sg U45799 ( .A(n26068), .X(n67578) );
  nand_x1_sg U45800 ( .A(n26069), .B(n57114), .X(n26068) );
  inv_x1_sg U45801 ( .A(n26072), .X(n67579) );
  nand_x1_sg U45802 ( .A(n26073), .B(n57114), .X(n26072) );
  inv_x1_sg U45803 ( .A(n26158), .X(n67583) );
  nand_x1_sg U45804 ( .A(n26157), .B(n57114), .X(n26158) );
  inv_x1_sg U45805 ( .A(n26164), .X(n67584) );
  nand_x1_sg U45806 ( .A(n26165), .B(n57114), .X(n26164) );
  inv_x1_sg U45807 ( .A(n26168), .X(n67585) );
  nand_x1_sg U45808 ( .A(n26169), .B(n57114), .X(n26168) );
  inv_x1_sg U45809 ( .A(n26174), .X(n67586) );
  nand_x1_sg U45810 ( .A(n26173), .B(n57114), .X(n26174) );
  nand_x1_sg U45811 ( .A(n57971), .B(n57970), .X(n42803) );
  inv_x1_sg U45812 ( .A(n57969), .X(n57971) );
  nand_x1_sg U45813 ( .A(n57978), .B(n57977), .X(n42809) );
  nand_x1_sg U45814 ( .A(n57981), .B(n57296), .X(n57978) );
  nand_x1_sg U45815 ( .A(n57430), .B(n57960), .X(n42802) );
  inv_x1_sg U45816 ( .A(n57959), .X(n57960) );
  nand_x1_sg U45817 ( .A(n57967), .B(n57966), .X(n42801) );
  inv_x1_sg U45818 ( .A(n57961), .X(n57967) );
  inv_x1_sg U45819 ( .A(n57965), .X(n57966) );
  nand_x1_sg U45820 ( .A(n57974), .B(n57973), .X(n42810) );
  nand_x1_sg U45821 ( .A(n58639), .B(n58640), .X(n57972) );
  nand_x1_sg U45822 ( .A(n57983), .B(n57982), .X(n42808) );
  nand_x1_sg U45823 ( .A(n57981), .B(n57920), .X(n57982) );
  nand_x1_sg U45824 ( .A(n57979), .B(n58476), .X(n57980) );
  nand_x1_sg U45825 ( .A(n30618), .B(n30619), .X(n42158) );
  nand_x1_sg U45826 ( .A(n30606), .B(n30607), .X(n42152) );
  nand_x1_sg U45827 ( .A(n30552), .B(n30553), .X(n42125) );
  nand_x1_sg U45828 ( .A(n30594), .B(n30595), .X(n42146) );
  nand_x1_sg U45829 ( .A(n29734), .B(n29735), .X(n41716) );
  nand_x1_sg U45830 ( .A(n29732), .B(n29733), .X(n41715) );
  nand_x1_sg U45831 ( .A(n29740), .B(n29741), .X(n41719) );
  nand_x1_sg U45832 ( .A(n29738), .B(n29739), .X(n41718) );
  nand_x1_sg U45833 ( .A(n29722), .B(n29723), .X(n41710) );
  nand_x1_sg U45834 ( .A(n29720), .B(n29721), .X(n41709) );
  nand_x1_sg U45835 ( .A(n29728), .B(n29729), .X(n41713) );
  nand_x1_sg U45836 ( .A(n29726), .B(n29727), .X(n41712) );
  nand_x1_sg U45837 ( .A(n29758), .B(n29759), .X(n41728) );
  nand_x1_sg U45838 ( .A(n29756), .B(n29757), .X(n41727) );
  nand_x1_sg U45839 ( .A(n29764), .B(n29765), .X(n41731) );
  nand_x1_sg U45840 ( .A(n29762), .B(n29763), .X(n41730) );
  nand_x1_sg U45841 ( .A(n29746), .B(n29747), .X(n41722) );
  nand_x1_sg U45842 ( .A(n29744), .B(n29745), .X(n41721) );
  nand_x1_sg U45843 ( .A(n29752), .B(n29753), .X(n41725) );
  nand_x1_sg U45844 ( .A(n29750), .B(n29751), .X(n41724) );
  nand_x1_sg U45845 ( .A(n31990), .B(n31991), .X(n42807) );
  nand_x1_sg U45846 ( .A(n31980), .B(n31981), .X(n42806) );
  nand_x1_sg U45847 ( .A(n57298), .B(n31968), .X(n31981) );
  nand_x1_sg U45848 ( .A(n31969), .B(n31970), .X(n42805) );
  nor_x1_sg U45849 ( .A(n31973), .B(n31974), .X(n31972) );
  nand_x1_sg U45850 ( .A(n31921), .B(n31922), .X(n42804) );
  nand_x1_sg U45851 ( .A(n68266), .B(n31923), .X(n31922) );
  nand_x1_sg U45852 ( .A(n57300), .B(n31968), .X(n31921) );
  nand_x1_sg U45853 ( .A(n31924), .B(n31925), .X(n31923) );
  nand_x1_sg U45854 ( .A(n29582), .B(n29583), .X(n41640) );
  nand_x1_sg U45855 ( .A(n29580), .B(n29581), .X(n41639) );
  nand_x1_sg U45856 ( .A(n29588), .B(n29589), .X(n41643) );
  nand_x1_sg U45857 ( .A(n29586), .B(n29587), .X(n41642) );
  nand_x1_sg U45858 ( .A(n29570), .B(n29571), .X(n41634) );
  nand_x1_sg U45859 ( .A(n29568), .B(n29569), .X(n41633) );
  nand_x1_sg U45860 ( .A(n29576), .B(n29577), .X(n41637) );
  nand_x1_sg U45861 ( .A(n29574), .B(n29575), .X(n41636) );
  nand_x1_sg U45862 ( .A(n29606), .B(n29607), .X(n41652) );
  nand_x1_sg U45863 ( .A(n29604), .B(n29605), .X(n41651) );
  nand_x1_sg U45864 ( .A(n29612), .B(n29613), .X(n41655) );
  nand_x1_sg U45865 ( .A(n29610), .B(n29611), .X(n41654) );
  nand_x1_sg U45866 ( .A(n29594), .B(n29595), .X(n41646) );
  nand_x1_sg U45867 ( .A(n29592), .B(n29593), .X(n41645) );
  nand_x1_sg U45868 ( .A(n29600), .B(n29601), .X(n41649) );
  nand_x1_sg U45869 ( .A(n29598), .B(n29599), .X(n41648) );
  nand_x1_sg U45870 ( .A(n29534), .B(n29535), .X(n41616) );
  nand_x1_sg U45871 ( .A(n29532), .B(n29533), .X(n41615) );
  nand_x1_sg U45872 ( .A(n29540), .B(n29541), .X(n41619) );
  nand_x1_sg U45873 ( .A(n29538), .B(n29539), .X(n41618) );
  nand_x1_sg U45874 ( .A(n29522), .B(n29523), .X(n41610) );
  nand_x1_sg U45875 ( .A(n29520), .B(n29521), .X(n41609) );
  nand_x1_sg U45876 ( .A(n29528), .B(n29529), .X(n41613) );
  nand_x1_sg U45877 ( .A(n29526), .B(n29527), .X(n41612) );
  nand_x1_sg U45878 ( .A(n29558), .B(n29559), .X(n41628) );
  nand_x1_sg U45879 ( .A(n29556), .B(n29557), .X(n41627) );
  nand_x1_sg U45880 ( .A(n29564), .B(n29565), .X(n41631) );
  nand_x1_sg U45881 ( .A(n29562), .B(n29563), .X(n41630) );
  nand_x1_sg U45882 ( .A(n29546), .B(n29547), .X(n41622) );
  nand_x1_sg U45883 ( .A(n29544), .B(n29545), .X(n41621) );
  nand_x1_sg U45884 ( .A(n29552), .B(n29553), .X(n41625) );
  nand_x1_sg U45885 ( .A(n29550), .B(n29551), .X(n41624) );
  nand_x1_sg U45886 ( .A(n29678), .B(n29679), .X(n41688) );
  nand_x1_sg U45887 ( .A(n29676), .B(n29677), .X(n41687) );
  nand_x1_sg U45888 ( .A(n29684), .B(n29685), .X(n41691) );
  nand_x1_sg U45889 ( .A(n29682), .B(n29683), .X(n41690) );
  nand_x1_sg U45890 ( .A(n29666), .B(n29667), .X(n41682) );
  nand_x1_sg U45891 ( .A(n29664), .B(n29665), .X(n41681) );
  nand_x1_sg U45892 ( .A(n29672), .B(n29673), .X(n41685) );
  nand_x1_sg U45893 ( .A(n29670), .B(n29671), .X(n41684) );
  nand_x1_sg U45894 ( .A(n29702), .B(n29703), .X(n41700) );
  nand_x1_sg U45895 ( .A(n29700), .B(n29701), .X(n41699) );
  nand_x1_sg U45896 ( .A(n29708), .B(n29709), .X(n41703) );
  nand_x1_sg U45897 ( .A(n29706), .B(n29707), .X(n41702) );
  nand_x1_sg U45898 ( .A(n29690), .B(n29691), .X(n41694) );
  nand_x1_sg U45899 ( .A(n29688), .B(n29689), .X(n41693) );
  nand_x1_sg U45900 ( .A(n29696), .B(n29697), .X(n41697) );
  nand_x1_sg U45901 ( .A(n29694), .B(n29695), .X(n41696) );
  nand_x1_sg U45902 ( .A(n29630), .B(n29631), .X(n41664) );
  nand_x1_sg U45903 ( .A(n29628), .B(n29629), .X(n41663) );
  nand_x1_sg U45904 ( .A(n29636), .B(n29637), .X(n41667) );
  nand_x1_sg U45905 ( .A(n29634), .B(n29635), .X(n41666) );
  nand_x1_sg U45906 ( .A(n29618), .B(n29619), .X(n41658) );
  nand_x1_sg U45907 ( .A(n29616), .B(n29617), .X(n41657) );
  nand_x1_sg U45908 ( .A(n29624), .B(n29625), .X(n41661) );
  nand_x1_sg U45909 ( .A(n29622), .B(n29623), .X(n41660) );
  nand_x1_sg U45910 ( .A(n29654), .B(n29655), .X(n41676) );
  nand_x1_sg U45911 ( .A(n29652), .B(n29653), .X(n41675) );
  nand_x1_sg U45912 ( .A(n29660), .B(n29661), .X(n41679) );
  nand_x1_sg U45913 ( .A(n29658), .B(n29659), .X(n41678) );
  nand_x1_sg U45914 ( .A(n29642), .B(n29643), .X(n41670) );
  nand_x1_sg U45915 ( .A(n29640), .B(n29641), .X(n41669) );
  nand_x1_sg U45916 ( .A(n29648), .B(n29649), .X(n41673) );
  nand_x1_sg U45917 ( .A(n29646), .B(n29647), .X(n41672) );
  nand_x1_sg U45918 ( .A(n30012), .B(n30013), .X(n41855) );
  nand_x1_sg U45919 ( .A(n30010), .B(n30011), .X(n41854) );
  nand_x1_sg U45920 ( .A(n30018), .B(n30019), .X(n41858) );
  nand_x1_sg U45921 ( .A(n30016), .B(n30017), .X(n41857) );
  nand_x1_sg U45922 ( .A(n30000), .B(n30001), .X(n41849) );
  nand_x1_sg U45923 ( .A(n29998), .B(n29999), .X(n41848) );
  nand_x1_sg U45924 ( .A(n30006), .B(n30007), .X(n41852) );
  nand_x1_sg U45925 ( .A(n30004), .B(n30005), .X(n41851) );
  nand_x1_sg U45926 ( .A(n30036), .B(n30037), .X(n41867) );
  nand_x1_sg U45927 ( .A(n30034), .B(n30035), .X(n41866) );
  nand_x1_sg U45928 ( .A(n30042), .B(n30043), .X(n41870) );
  nand_x1_sg U45929 ( .A(n30040), .B(n30041), .X(n41869) );
  nand_x1_sg U45930 ( .A(n30024), .B(n30025), .X(n41861) );
  nand_x1_sg U45931 ( .A(n30022), .B(n30023), .X(n41860) );
  nand_x1_sg U45932 ( .A(n30030), .B(n30031), .X(n41864) );
  nand_x1_sg U45933 ( .A(n30028), .B(n30029), .X(n41863) );
  nand_x1_sg U45934 ( .A(n29974), .B(n29975), .X(n41836) );
  nand_x1_sg U45935 ( .A(n29972), .B(n29973), .X(n41835) );
  nand_x1_sg U45936 ( .A(n29980), .B(n29981), .X(n41839) );
  nand_x1_sg U45937 ( .A(n29978), .B(n29979), .X(n41838) );
  nand_x1_sg U45938 ( .A(n29962), .B(n29963), .X(n41830) );
  nand_x1_sg U45939 ( .A(n29960), .B(n29961), .X(n41829) );
  nand_x1_sg U45940 ( .A(n29968), .B(n29969), .X(n41833) );
  nand_x1_sg U45941 ( .A(n29966), .B(n29967), .X(n41832) );
  nand_x1_sg U45942 ( .A(n29964), .B(n29965), .X(n41831) );
  nand_x1_sg U45943 ( .A(n29716), .B(n29717), .X(n41707) );
  nand_x1_sg U45944 ( .A(n30014), .B(n30015), .X(n41856) );
  nand_x1_sg U45945 ( .A(n30002), .B(n30003), .X(n41850) );
  nand_x1_sg U45946 ( .A(n29988), .B(n29989), .X(n41843) );
  nand_x1_sg U45947 ( .A(n29986), .B(n29987), .X(n41842) );
  nand_x1_sg U45948 ( .A(n29994), .B(n29995), .X(n41846) );
  nand_x1_sg U45949 ( .A(n29992), .B(n29993), .X(n41845) );
  nand_x1_sg U45950 ( .A(n30108), .B(n30109), .X(n41903) );
  nand_x1_sg U45951 ( .A(n30106), .B(n30107), .X(n41902) );
  nand_x1_sg U45952 ( .A(n30114), .B(n30115), .X(n41906) );
  nand_x1_sg U45953 ( .A(n30112), .B(n30113), .X(n41905) );
  nand_x1_sg U45954 ( .A(n30096), .B(n30097), .X(n41897) );
  nand_x1_sg U45955 ( .A(n30094), .B(n30095), .X(n41896) );
  nand_x1_sg U45956 ( .A(n30102), .B(n30103), .X(n41900) );
  nand_x1_sg U45957 ( .A(n30100), .B(n30101), .X(n41899) );
  nand_x1_sg U45958 ( .A(n30132), .B(n30133), .X(n41915) );
  nand_x1_sg U45959 ( .A(n30130), .B(n30131), .X(n41914) );
  nand_x1_sg U45960 ( .A(n30074), .B(n30075), .X(n41886) );
  nand_x1_sg U45961 ( .A(n30122), .B(n30123), .X(n41910) );
  nand_x1_sg U45962 ( .A(n30120), .B(n30121), .X(n41909) );
  nand_x1_sg U45963 ( .A(n30118), .B(n30119), .X(n41908) );
  nand_x1_sg U45964 ( .A(n30126), .B(n30127), .X(n41912) );
  nand_x1_sg U45965 ( .A(n30124), .B(n30125), .X(n41911) );
  nand_x1_sg U45966 ( .A(n30060), .B(n30061), .X(n41879) );
  nand_x1_sg U45967 ( .A(n30058), .B(n30059), .X(n41878) );
  nand_x1_sg U45968 ( .A(n30066), .B(n30067), .X(n41882) );
  nand_x1_sg U45969 ( .A(n30064), .B(n30065), .X(n41881) );
  nand_x1_sg U45970 ( .A(n30048), .B(n30049), .X(n41873) );
  nand_x1_sg U45971 ( .A(n30046), .B(n30047), .X(n41872) );
  nand_x1_sg U45972 ( .A(n30054), .B(n30055), .X(n41876) );
  nand_x1_sg U45973 ( .A(n30052), .B(n30053), .X(n41875) );
  nand_x1_sg U45974 ( .A(n30084), .B(n30085), .X(n41891) );
  nand_x1_sg U45975 ( .A(n30082), .B(n30083), .X(n41890) );
  nand_x1_sg U45976 ( .A(n30090), .B(n30091), .X(n41894) );
  nand_x1_sg U45977 ( .A(n30088), .B(n30089), .X(n41893) );
  nand_x1_sg U45978 ( .A(n30072), .B(n30073), .X(n41885) );
  nand_x1_sg U45979 ( .A(n30070), .B(n30071), .X(n41884) );
  nand_x1_sg U45980 ( .A(n30078), .B(n30079), .X(n41888) );
  nand_x1_sg U45981 ( .A(n30076), .B(n30077), .X(n41887) );
  nand_x1_sg U45982 ( .A(n29830), .B(n29831), .X(n41764) );
  nand_x1_sg U45983 ( .A(n29828), .B(n29829), .X(n41763) );
  nand_x1_sg U45984 ( .A(n29836), .B(n29837), .X(n41767) );
  nand_x1_sg U45985 ( .A(n29834), .B(n29835), .X(n41766) );
  nand_x1_sg U45986 ( .A(n29818), .B(n29819), .X(n41758) );
  nand_x1_sg U45987 ( .A(n29816), .B(n29817), .X(n41757) );
  nand_x1_sg U45988 ( .A(n29824), .B(n29825), .X(n41761) );
  nand_x1_sg U45989 ( .A(n29822), .B(n29823), .X(n41760) );
  nand_x1_sg U45990 ( .A(n29854), .B(n29855), .X(n41776) );
  nand_x1_sg U45991 ( .A(n29852), .B(n29853), .X(n41775) );
  nand_x1_sg U45992 ( .A(n29860), .B(n29861), .X(n41779) );
  nand_x1_sg U45993 ( .A(n29858), .B(n29859), .X(n41778) );
  nand_x1_sg U45994 ( .A(n29842), .B(n29843), .X(n41770) );
  nand_x1_sg U45995 ( .A(n29840), .B(n29841), .X(n41769) );
  nand_x1_sg U45996 ( .A(n29848), .B(n29849), .X(n41773) );
  nand_x1_sg U45997 ( .A(n29846), .B(n29847), .X(n41772) );
  nand_x1_sg U45998 ( .A(n29782), .B(n29783), .X(n41740) );
  nand_x1_sg U45999 ( .A(n29780), .B(n29781), .X(n41739) );
  nand_x1_sg U46000 ( .A(n29788), .B(n29789), .X(n41743) );
  nand_x1_sg U46001 ( .A(n29786), .B(n29787), .X(n41742) );
  nand_x1_sg U46002 ( .A(n29770), .B(n29771), .X(n41734) );
  nand_x1_sg U46003 ( .A(n29768), .B(n29769), .X(n41733) );
  nand_x1_sg U46004 ( .A(n29776), .B(n29777), .X(n41737) );
  nand_x1_sg U46005 ( .A(n29774), .B(n29775), .X(n41736) );
  nand_x1_sg U46006 ( .A(n29806), .B(n29807), .X(n41752) );
  nand_x1_sg U46007 ( .A(n29804), .B(n29805), .X(n41751) );
  nand_x1_sg U46008 ( .A(n29812), .B(n29813), .X(n41755) );
  nand_x1_sg U46009 ( .A(n29810), .B(n29811), .X(n41754) );
  nand_x1_sg U46010 ( .A(n29794), .B(n29795), .X(n41746) );
  nand_x1_sg U46011 ( .A(n29792), .B(n29793), .X(n41745) );
  nand_x1_sg U46012 ( .A(n29800), .B(n29801), .X(n41749) );
  nand_x1_sg U46013 ( .A(n29798), .B(n29799), .X(n41748) );
  nand_x1_sg U46014 ( .A(n29926), .B(n29927), .X(n41812) );
  nand_x1_sg U46015 ( .A(n29924), .B(n29925), .X(n41811) );
  nand_x1_sg U46016 ( .A(n29932), .B(n29933), .X(n41815) );
  nand_x1_sg U46017 ( .A(n29930), .B(n29931), .X(n41814) );
  nand_x1_sg U46018 ( .A(n29914), .B(n29915), .X(n41806) );
  nand_x1_sg U46019 ( .A(n29912), .B(n29913), .X(n41805) );
  nand_x1_sg U46020 ( .A(n29920), .B(n29921), .X(n41809) );
  nand_x1_sg U46021 ( .A(n29918), .B(n29919), .X(n41808) );
  nand_x1_sg U46022 ( .A(n29950), .B(n29951), .X(n41824) );
  nand_x1_sg U46023 ( .A(n29948), .B(n29949), .X(n41823) );
  nand_x1_sg U46024 ( .A(n29956), .B(n29957), .X(n41827) );
  nand_x1_sg U46025 ( .A(n29954), .B(n29955), .X(n41826) );
  nand_x1_sg U46026 ( .A(n29938), .B(n29939), .X(n41818) );
  nand_x1_sg U46027 ( .A(n29936), .B(n29937), .X(n41817) );
  nand_x1_sg U46028 ( .A(n29944), .B(n29945), .X(n41821) );
  nand_x1_sg U46029 ( .A(n29942), .B(n29943), .X(n41820) );
  nand_x1_sg U46030 ( .A(n29878), .B(n29879), .X(n41788) );
  nand_x1_sg U46031 ( .A(n29876), .B(n29877), .X(n41787) );
  nand_x1_sg U46032 ( .A(n29884), .B(n29885), .X(n41791) );
  nand_x1_sg U46033 ( .A(n29882), .B(n29883), .X(n41790) );
  nand_x1_sg U46034 ( .A(n29866), .B(n29867), .X(n41782) );
  nand_x1_sg U46035 ( .A(n29864), .B(n29865), .X(n41781) );
  nand_x1_sg U46036 ( .A(n29872), .B(n29873), .X(n41785) );
  nand_x1_sg U46037 ( .A(n29870), .B(n29871), .X(n41784) );
  nand_x1_sg U46038 ( .A(n29902), .B(n29903), .X(n41800) );
  nand_x1_sg U46039 ( .A(n29900), .B(n29901), .X(n41799) );
  nand_x1_sg U46040 ( .A(n29908), .B(n29909), .X(n41803) );
  nand_x1_sg U46041 ( .A(n29906), .B(n29907), .X(n41802) );
  nand_x1_sg U46042 ( .A(n29890), .B(n29891), .X(n41794) );
  nand_x1_sg U46043 ( .A(n29888), .B(n29889), .X(n41793) );
  nand_x1_sg U46044 ( .A(n29896), .B(n29897), .X(n41797) );
  nand_x1_sg U46045 ( .A(n29894), .B(n29895), .X(n41796) );
  nand_x1_sg U46046 ( .A(n29382), .B(n29383), .X(n41540) );
  nand_x1_sg U46047 ( .A(n29386), .B(n29387), .X(n41542) );
  nand_x1_sg U46048 ( .A(n30316), .B(n30317), .X(n42007) );
  nand_x1_sg U46049 ( .A(n30328), .B(n30329), .X(n42013) );
  nand_x1_sg U46050 ( .A(n30310), .B(n30311), .X(n42004) );
  nand_x1_sg U46051 ( .A(n30298), .B(n30299), .X(n41998) );
  nand_x1_sg U46052 ( .A(n30286), .B(n30287), .X(n41992) );
  nand_x1_sg U46053 ( .A(n30280), .B(n30281), .X(n41989) );
  nand_x1_sg U46054 ( .A(n30406), .B(n30407), .X(n42052) );
  nand_x1_sg U46055 ( .A(n30148), .B(n30149), .X(n41923) );
  nand_x1_sg U46056 ( .A(n30364), .B(n30365), .X(n42031) );
  nand_x1_sg U46057 ( .A(n30340), .B(n30341), .X(n42019) );
  nand_x1_sg U46058 ( .A(n29596), .B(n29597), .X(n41647) );
  nand_x1_sg U46059 ( .A(n29898), .B(n29899), .X(n41798) );
  nand_x1_sg U46060 ( .A(n29536), .B(n29537), .X(n41617) );
  nand_x1_sg U46061 ( .A(n29530), .B(n29531), .X(n41614) );
  nand_x1_sg U46062 ( .A(n30268), .B(n30269), .X(n41983) );
  nand_x1_sg U46063 ( .A(n30322), .B(n30323), .X(n42010) );
  nand_x1_sg U46064 ( .A(n29698), .B(n29699), .X(n41698) );
  nand_x1_sg U46065 ( .A(n30292), .B(n30293), .X(n41995) );
  nand_x1_sg U46066 ( .A(n30472), .B(n30473), .X(n42085) );
  nand_x1_sg U46067 ( .A(n30442), .B(n30443), .X(n42070) );
  nand_x1_sg U46068 ( .A(n29584), .B(n29585), .X(n41641) );
  nand_x1_sg U46069 ( .A(n29366), .B(n29367), .X(n41532) );
  nand_x1_sg U46070 ( .A(n29362), .B(n29363), .X(n41530) );
  nand_x1_sg U46071 ( .A(n29364), .B(n29365), .X(n41531) );
  nand_x1_sg U46072 ( .A(n30208), .B(n30209), .X(n41953) );
  nand_x1_sg U46073 ( .A(n30508), .B(n30509), .X(n42103) );
  nand_x1_sg U46074 ( .A(n30304), .B(n30305), .X(n42001) );
  nand_x1_sg U46075 ( .A(n29406), .B(n29407), .X(n41552) );
  nand_x1_sg U46076 ( .A(n29446), .B(n29447), .X(n41572) );
  nand_x1_sg U46077 ( .A(n29820), .B(n29821), .X(n41759) );
  nand_x1_sg U46078 ( .A(n29704), .B(n29705), .X(n41701) );
  nand_x1_sg U46079 ( .A(n29384), .B(n29385), .X(n41541) );
  nand_x1_sg U46080 ( .A(n29686), .B(n29687), .X(n41692) );
  nand_x1_sg U46081 ( .A(n29680), .B(n29681), .X(n41689) );
  nand_x1_sg U46082 ( .A(n29856), .B(n29857), .X(n41777) );
  nand_x1_sg U46083 ( .A(n29638), .B(n29639), .X(n41668) );
  nand_x1_sg U46084 ( .A(n29668), .B(n29669), .X(n41683) );
  nand_x1_sg U46085 ( .A(n29662), .B(n29663), .X(n41680) );
  nand_x1_sg U46086 ( .A(n29626), .B(n29627), .X(n41662) );
  nand_x1_sg U46087 ( .A(n29620), .B(n29621), .X(n41659) );
  nand_x1_sg U46088 ( .A(n29614), .B(n29615), .X(n41656) );
  nand_x1_sg U46089 ( .A(n29602), .B(n29603), .X(n41650) );
  nand_x1_sg U46090 ( .A(n29674), .B(n29675), .X(n41686) );
  nand_x1_sg U46091 ( .A(n29656), .B(n29657), .X(n41677) );
  nand_x1_sg U46092 ( .A(n29650), .B(n29651), .X(n41674) );
  nand_x1_sg U46093 ( .A(n29644), .B(n29645), .X(n41671) );
  nand_x1_sg U46094 ( .A(n29578), .B(n29579), .X(n41638) );
  nand_x1_sg U46095 ( .A(n29566), .B(n29567), .X(n41632) );
  nand_x1_sg U46096 ( .A(n30358), .B(n30359), .X(n42028) );
  nand_x1_sg U46097 ( .A(n29518), .B(n29519), .X(n41608) );
  nand_x1_sg U46098 ( .A(n29554), .B(n29555), .X(n41626) );
  nand_x1_sg U46099 ( .A(n29542), .B(n29543), .X(n41620) );
  nand_x1_sg U46100 ( .A(n29524), .B(n29525), .X(n41611) );
  nand_x1_sg U46101 ( .A(n29590), .B(n29591), .X(n41644) );
  nand_x1_sg U46102 ( .A(n29784), .B(n29785), .X(n41741) );
  nand_x1_sg U46103 ( .A(n29400), .B(n29401), .X(n41549) );
  nand_x1_sg U46104 ( .A(n29904), .B(n29905), .X(n41801) );
  nand_x1_sg U46105 ( .A(n29488), .B(n29489), .X(n41593) );
  nand_x1_sg U46106 ( .A(n30044), .B(n30045), .X(n41871) );
  nand_x1_sg U46107 ( .A(n29376), .B(n29377), .X(n41537) );
  nand_x1_sg U46108 ( .A(n29910), .B(n29911), .X(n41804) );
  nand_x1_sg U46109 ( .A(n29710), .B(n29711), .X(n41704) );
  nand_x1_sg U46110 ( .A(n29754), .B(n29755), .X(n41726) );
  nand_x1_sg U46111 ( .A(n29730), .B(n29731), .X(n41714) );
  nand_x1_sg U46112 ( .A(n30196), .B(n30197), .X(n41947) );
  nand_x1_sg U46113 ( .A(n30382), .B(n30383), .X(n42040) );
  nand_x1_sg U46114 ( .A(n30154), .B(n30155), .X(n41926) );
  nand_x1_sg U46115 ( .A(n30172), .B(n30173), .X(n41935) );
  nand_x1_sg U46116 ( .A(n30424), .B(n30425), .X(n42061) );
  nand_x1_sg U46117 ( .A(n29358), .B(n29359), .X(n41528) );
  nand_x1_sg U46118 ( .A(n30376), .B(n30377), .X(n42037) );
  nand_x1_sg U46119 ( .A(n30202), .B(n30203), .X(n41950) );
  nand_x1_sg U46120 ( .A(n30190), .B(n30191), .X(n41944) );
  nand_x1_sg U46121 ( .A(n30184), .B(n30185), .X(n41941) );
  nand_x1_sg U46122 ( .A(n29356), .B(n29357), .X(n41527) );
  nand_x1_sg U46123 ( .A(n29354), .B(n29355), .X(n41526) );
  nand_x1_sg U46124 ( .A(n29372), .B(n29373), .X(n41535) );
  nand_x1_sg U46125 ( .A(n30460), .B(n30461), .X(n42079) );
  nand_x1_sg U46126 ( .A(n29760), .B(n29761), .X(n41729) );
  nand_x1_sg U46127 ( .A(n29718), .B(n29719), .X(n41708) );
  nand_x1_sg U46128 ( .A(n30142), .B(n30143), .X(n41920) );
  nand_x1_sg U46129 ( .A(n30612), .B(n30613), .X(n42155) );
  nand_x1_sg U46130 ( .A(n30588), .B(n30589), .X(n42143) );
  nand_x1_sg U46131 ( .A(n30534), .B(n30535), .X(n42116) );
  nand_x1_sg U46132 ( .A(n29742), .B(n29743), .X(n41720) );
  nand_x1_sg U46133 ( .A(n29736), .B(n29737), .X(n41717) );
  nand_x1_sg U46134 ( .A(n29724), .B(n29725), .X(n41711) );
  nand_x1_sg U46135 ( .A(n29346), .B(n29347), .X(n41522) );
  nand_x1_sg U46136 ( .A(n30214), .B(n30215), .X(n41956) );
  nand_x1_sg U46137 ( .A(n30220), .B(n30221), .X(n41959) );
  nand_x1_sg U46138 ( .A(n30582), .B(n30583), .X(n42140) );
  nand_x1_sg U46139 ( .A(n30576), .B(n30577), .X(n42137) );
  nand_x1_sg U46140 ( .A(n30546), .B(n30547), .X(n42122) );
  nand_x1_sg U46141 ( .A(n30540), .B(n30541), .X(n42119) );
  nand_x1_sg U46142 ( .A(n30250), .B(n30251), .X(n41974) );
  nand_x1_sg U46143 ( .A(n30466), .B(n30467), .X(n42082) );
  nand_x1_sg U46144 ( .A(n30244), .B(n30245), .X(n41971) );
  nand_x1_sg U46145 ( .A(n30238), .B(n30239), .X(n41968) );
  nand_x1_sg U46146 ( .A(n30490), .B(n30491), .X(n42094) );
  nand_x1_sg U46147 ( .A(n29374), .B(n29375), .X(n41536) );
  nand_x1_sg U46148 ( .A(n30484), .B(n30485), .X(n42091) );
  nand_x1_sg U46149 ( .A(n30274), .B(n30275), .X(n41986) );
  nand_x1_sg U46150 ( .A(n30454), .B(n30455), .X(n42076) );
  nand_x1_sg U46151 ( .A(n30394), .B(n30395), .X(n42046) );
  nand_x1_sg U46152 ( .A(n30370), .B(n30371), .X(n42034) );
  nand_x1_sg U46153 ( .A(n30346), .B(n30347), .X(n42022) );
  nand_x1_sg U46154 ( .A(n30256), .B(n30257), .X(n41977) );
  nand_x1_sg U46155 ( .A(n30352), .B(n30353), .X(n42025) );
  nand_x1_sg U46156 ( .A(n30232), .B(n30233), .X(n41965) );
  nand_x1_sg U46157 ( .A(n30496), .B(n30497), .X(n42097) );
  nand_x1_sg U46158 ( .A(n29368), .B(n29369), .X(n41533) );
  nand_x1_sg U46159 ( .A(n29370), .B(n29371), .X(n41534) );
  nand_x1_sg U46160 ( .A(n30178), .B(n30179), .X(n41938) );
  nand_x1_sg U46161 ( .A(n30166), .B(n30167), .X(n41932) );
  nand_x1_sg U46162 ( .A(n30448), .B(n30449), .X(n42073) );
  nand_x1_sg U46163 ( .A(n30430), .B(n30431), .X(n42064) );
  nand_x1_sg U46164 ( .A(n30418), .B(n30419), .X(n42058) );
  nand_x1_sg U46165 ( .A(n30412), .B(n30413), .X(n42055) );
  nand_x1_sg U46166 ( .A(n30334), .B(n30335), .X(n42016) );
  nand_x1_sg U46167 ( .A(n30514), .B(n30515), .X(n42106) );
  nand_x1_sg U46168 ( .A(n30436), .B(n30437), .X(n42067) );
  nand_x1_sg U46169 ( .A(n29360), .B(n29361), .X(n41529) );
  nand_x1_sg U46170 ( .A(n30478), .B(n30479), .X(n42088) );
  nand_x1_sg U46171 ( .A(n30388), .B(n30389), .X(n42043) );
  nand_x1_sg U46172 ( .A(n30502), .B(n30503), .X(n42100) );
  nand_x1_sg U46173 ( .A(n30160), .B(n30161), .X(n41929) );
  nand_x1_sg U46174 ( .A(n29414), .B(n29415), .X(n41556) );
  nand_x1_sg U46175 ( .A(n29344), .B(n29345), .X(n41521) );
  nand_x1_sg U46176 ( .A(n29802), .B(n29803), .X(n41750) );
  nand_x1_sg U46177 ( .A(n29790), .B(n29791), .X(n41744) );
  nand_x1_sg U46178 ( .A(n30526), .B(n30527), .X(n42112) );
  nand_x1_sg U46179 ( .A(n30524), .B(n30525), .X(n42111) );
  nand_x1_sg U46180 ( .A(n29714), .B(n29715), .X(n41706) );
  nand_x1_sg U46181 ( .A(n29712), .B(n29713), .X(n41705) );
  nand_x1_sg U46182 ( .A(n29432), .B(n29433), .X(n41565) );
  nand_x1_sg U46183 ( .A(n29430), .B(n29431), .X(n41564) );
  nand_x1_sg U46184 ( .A(n29438), .B(n29439), .X(n41568) );
  nand_x1_sg U46185 ( .A(n29436), .B(n29437), .X(n41567) );
  nand_x1_sg U46186 ( .A(n29420), .B(n29421), .X(n41559) );
  nand_x1_sg U46187 ( .A(n29418), .B(n29419), .X(n41558) );
  nand_x1_sg U46188 ( .A(n29426), .B(n29427), .X(n41562) );
  nand_x1_sg U46189 ( .A(n29424), .B(n29425), .X(n41561) );
  nand_x1_sg U46190 ( .A(n30050), .B(n30051), .X(n41874) );
  nand_x1_sg U46191 ( .A(n29350), .B(n29351), .X(n41524) );
  nand_x1_sg U46192 ( .A(n30038), .B(n30039), .X(n41868) );
  nand_x1_sg U46193 ( .A(n30032), .B(n30033), .X(n41865) );
  nand_x1_sg U46194 ( .A(n29970), .B(n29971), .X(n41834) );
  nand_x1_sg U46195 ( .A(n29976), .B(n29977), .X(n41837) );
  nand_x1_sg U46196 ( .A(n29916), .B(n29917), .X(n41807) );
  nand_x1_sg U46197 ( .A(n30128), .B(n30129), .X(n41913) );
  nand_x1_sg U46198 ( .A(n30062), .B(n30063), .X(n41880) );
  nand_x1_sg U46199 ( .A(n30056), .B(n30057), .X(n41877) );
  nand_x1_sg U46200 ( .A(n29394), .B(n29395), .X(n41546) );
  nand_x1_sg U46201 ( .A(n29392), .B(n29393), .X(n41545) );
  nand_x1_sg U46202 ( .A(n30092), .B(n30093), .X(n41895) );
  nand_x1_sg U46203 ( .A(n30104), .B(n30105), .X(n41901) );
  nand_x1_sg U46204 ( .A(n30086), .B(n30087), .X(n41892) );
  nand_x1_sg U46205 ( .A(n30080), .B(n30081), .X(n41889) );
  nand_x1_sg U46206 ( .A(n29504), .B(n29505), .X(n41601) );
  nand_x1_sg U46207 ( .A(n29502), .B(n29503), .X(n41600) );
  nand_x1_sg U46208 ( .A(n29510), .B(n29511), .X(n41604) );
  nand_x1_sg U46209 ( .A(n29508), .B(n29509), .X(n41603) );
  nand_x1_sg U46210 ( .A(n29492), .B(n29493), .X(n41595) );
  nand_x1_sg U46211 ( .A(n29490), .B(n29491), .X(n41594) );
  nand_x1_sg U46212 ( .A(n29498), .B(n29499), .X(n41598) );
  nand_x1_sg U46213 ( .A(n29496), .B(n29497), .X(n41597) );
  nand_x1_sg U46214 ( .A(n29516), .B(n29517), .X(n41607) );
  nand_x1_sg U46215 ( .A(n29928), .B(n29929), .X(n41813) );
  nand_x1_sg U46216 ( .A(n29922), .B(n29923), .X(n41810) );
  nand_x1_sg U46217 ( .A(n29412), .B(n29413), .X(n41555) );
  nand_x1_sg U46218 ( .A(n29934), .B(n29935), .X(n41816) );
  nand_x1_sg U46219 ( .A(n29514), .B(n29515), .X(n41606) );
  nand_x1_sg U46220 ( .A(n29946), .B(n29947), .X(n41822) );
  nand_x1_sg U46221 ( .A(n29952), .B(n29953), .X(n41825) );
  nand_x1_sg U46222 ( .A(n29456), .B(n29457), .X(n41577) );
  nand_x1_sg U46223 ( .A(n29454), .B(n29455), .X(n41576) );
  nand_x1_sg U46224 ( .A(n29462), .B(n29463), .X(n41580) );
  nand_x1_sg U46225 ( .A(n29460), .B(n29461), .X(n41579) );
  nand_x1_sg U46226 ( .A(n29444), .B(n29445), .X(n41571) );
  nand_x1_sg U46227 ( .A(n29442), .B(n29443), .X(n41570) );
  nand_x1_sg U46228 ( .A(n29450), .B(n29451), .X(n41574) );
  nand_x1_sg U46229 ( .A(n29448), .B(n29449), .X(n41573) );
  nand_x1_sg U46230 ( .A(n29480), .B(n29481), .X(n41589) );
  nand_x1_sg U46231 ( .A(n29478), .B(n29479), .X(n41588) );
  nand_x1_sg U46232 ( .A(n29486), .B(n29487), .X(n41592) );
  nand_x1_sg U46233 ( .A(n29484), .B(n29485), .X(n41591) );
  nand_x1_sg U46234 ( .A(n29468), .B(n29469), .X(n41583) );
  nand_x1_sg U46235 ( .A(n29466), .B(n29467), .X(n41582) );
  nand_x1_sg U46236 ( .A(n29474), .B(n29475), .X(n41586) );
  nand_x1_sg U46237 ( .A(n29472), .B(n29473), .X(n41585) );
  nand_x1_sg U46238 ( .A(n29632), .B(n29633), .X(n41665) );
  nand_x1_sg U46239 ( .A(n29608), .B(n29609), .X(n41653) );
  nand_x1_sg U46240 ( .A(n29572), .B(n29573), .X(n41635) );
  nand_x1_sg U46241 ( .A(n29808), .B(n29809), .X(n41753) );
  nand_x1_sg U46242 ( .A(n29398), .B(n29399), .X(n41548) );
  nand_x1_sg U46243 ( .A(n29396), .B(n29397), .X(n41547) );
  nand_x1_sg U46244 ( .A(n29692), .B(n29693), .X(n41695) );
  nand_x1_sg U46245 ( .A(n29892), .B(n29893), .X(n41795) );
  nand_x1_sg U46246 ( .A(n29352), .B(n29353), .X(n41525) );
  nand_x1_sg U46247 ( .A(n30008), .B(n30009), .X(n41853) );
  nand_x1_sg U46248 ( .A(n29378), .B(n29379), .X(n41538) );
  nand_x1_sg U46249 ( .A(n29422), .B(n29423), .X(n41560) );
  nand_x1_sg U46250 ( .A(n29772), .B(n29773), .X(n41735) );
  nand_x1_sg U46251 ( .A(n29874), .B(n29875), .X(n41786) );
  nand_x1_sg U46252 ( .A(n29886), .B(n29887), .X(n41792) );
  nand_x1_sg U46253 ( .A(n29868), .B(n29869), .X(n41783) );
  nand_x1_sg U46254 ( .A(n29814), .B(n29815), .X(n41756) );
  nand_x1_sg U46255 ( .A(n29826), .B(n29827), .X(n41762) );
  nand_x1_sg U46256 ( .A(n29506), .B(n29507), .X(n41602) );
  nand_x1_sg U46257 ( .A(n29778), .B(n29779), .X(n41738) );
  nand_x1_sg U46258 ( .A(n29850), .B(n29851), .X(n41774) );
  nand_x1_sg U46259 ( .A(n29862), .B(n29863), .X(n41780) );
  nand_x1_sg U46260 ( .A(n29560), .B(n29561), .X(n41629) );
  nand_x1_sg U46261 ( .A(n29548), .B(n29549), .X(n41623) );
  nand_x1_sg U46262 ( .A(n29990), .B(n29991), .X(n41844) );
  nand_x1_sg U46263 ( .A(n29388), .B(n29389), .X(n41543) );
  nand_x1_sg U46264 ( .A(n29838), .B(n29839), .X(n41768) );
  nand_x1_sg U46265 ( .A(n29832), .B(n29833), .X(n41765) );
  nand_x1_sg U46266 ( .A(n29880), .B(n29881), .X(n41789) );
  nand_x1_sg U46267 ( .A(n29402), .B(n29403), .X(n41550) );
  nand_x1_sg U46268 ( .A(n30098), .B(n30099), .X(n41898) );
  nand_x1_sg U46269 ( .A(n29796), .B(n29797), .X(n41747) );
  nand_x1_sg U46270 ( .A(n29940), .B(n29941), .X(n41819) );
  nand_x1_sg U46271 ( .A(n29512), .B(n29513), .X(n41605) );
  nand_x1_sg U46272 ( .A(n29500), .B(n29501), .X(n41599) );
  nand_x1_sg U46273 ( .A(n29494), .B(n29495), .X(n41596) );
  nand_x1_sg U46274 ( .A(n29766), .B(n29767), .X(n41732) );
  nand_x1_sg U46275 ( .A(n30068), .B(n30069), .X(n41883) );
  nand_x1_sg U46276 ( .A(n29458), .B(n29459), .X(n41578) );
  nand_x1_sg U46277 ( .A(n29410), .B(n29411), .X(n41554) );
  nand_x1_sg U46278 ( .A(n29996), .B(n29997), .X(n41847) );
  nand_x1_sg U46279 ( .A(n29982), .B(n29983), .X(n41840) );
  nand_x1_sg U46280 ( .A(n29984), .B(n29985), .X(n41841) );
  nand_x1_sg U46281 ( .A(n29408), .B(n29409), .X(n41553) );
  nand_x1_sg U46282 ( .A(n29390), .B(n29391), .X(n41544) );
  nand_x1_sg U46283 ( .A(n29434), .B(n29435), .X(n41566) );
  nand_x1_sg U46284 ( .A(n30026), .B(n30027), .X(n41862) );
  nand_x1_sg U46285 ( .A(n30020), .B(n30021), .X(n41859) );
  nand_x1_sg U46286 ( .A(n29482), .B(n29483), .X(n41590) );
  nand_x1_sg U46287 ( .A(n29476), .B(n29477), .X(n41587) );
  nand_x1_sg U46288 ( .A(n30110), .B(n30111), .X(n41904) );
  nand_x1_sg U46289 ( .A(n30522), .B(n30523), .X(n42110) );
  nand_x1_sg U46290 ( .A(n29348), .B(n29349), .X(n41523) );
  nand_x1_sg U46291 ( .A(n29380), .B(n29381), .X(n41539) );
  nand_x1_sg U46292 ( .A(n30116), .B(n30117), .X(n41907) );
  nand_x1_sg U46293 ( .A(n29958), .B(n29959), .X(n41828) );
  nand_x1_sg U46294 ( .A(n29470), .B(n29471), .X(n41584) );
  nand_x1_sg U46295 ( .A(n29416), .B(n29417), .X(n41557) );
  nand_x1_sg U46296 ( .A(n29844), .B(n29845), .X(n41771) );
  nand_x1_sg U46297 ( .A(n29404), .B(n29405), .X(n41551) );
  nand_x1_sg U46298 ( .A(n29464), .B(n29465), .X(n41581) );
  nand_x1_sg U46299 ( .A(n29452), .B(n29453), .X(n41575) );
  nand_x1_sg U46300 ( .A(n29440), .B(n29441), .X(n41569) );
  nand_x1_sg U46301 ( .A(n29428), .B(n29429), .X(n41563) );
  nand_x1_sg U46302 ( .A(n30392), .B(n30393), .X(n42045) );
  nand_x1_sg U46303 ( .A(n30390), .B(n30391), .X(n42044) );
  nand_x1_sg U46304 ( .A(n30398), .B(n30399), .X(n42048) );
  nand_x1_sg U46305 ( .A(n30396), .B(n30397), .X(n42047) );
  nand_x1_sg U46306 ( .A(n30380), .B(n30381), .X(n42039) );
  nand_x1_sg U46307 ( .A(n30378), .B(n30379), .X(n42038) );
  nand_x1_sg U46308 ( .A(n30386), .B(n30387), .X(n42042) );
  nand_x1_sg U46309 ( .A(n30384), .B(n30385), .X(n42041) );
  nand_x1_sg U46310 ( .A(n30416), .B(n30417), .X(n42057) );
  nand_x1_sg U46311 ( .A(n30414), .B(n30415), .X(n42056) );
  nand_x1_sg U46312 ( .A(n30422), .B(n30423), .X(n42060) );
  nand_x1_sg U46313 ( .A(n30420), .B(n30421), .X(n42059) );
  nand_x1_sg U46314 ( .A(n30404), .B(n30405), .X(n42051) );
  nand_x1_sg U46315 ( .A(n30402), .B(n30403), .X(n42050) );
  nand_x1_sg U46316 ( .A(n30410), .B(n30411), .X(n42054) );
  nand_x1_sg U46317 ( .A(n30408), .B(n30409), .X(n42053) );
  nand_x1_sg U46318 ( .A(n30344), .B(n30345), .X(n42021) );
  nand_x1_sg U46319 ( .A(n30342), .B(n30343), .X(n42020) );
  nand_x1_sg U46320 ( .A(n30350), .B(n30351), .X(n42024) );
  nand_x1_sg U46321 ( .A(n30348), .B(n30349), .X(n42023) );
  nand_x1_sg U46322 ( .A(n30332), .B(n30333), .X(n42015) );
  nand_x1_sg U46323 ( .A(n30330), .B(n30331), .X(n42014) );
  nand_x1_sg U46324 ( .A(n30338), .B(n30339), .X(n42018) );
  nand_x1_sg U46325 ( .A(n30336), .B(n30337), .X(n42017) );
  nand_x1_sg U46326 ( .A(n30368), .B(n30369), .X(n42033) );
  nand_x1_sg U46327 ( .A(n30366), .B(n30367), .X(n42032) );
  nand_x1_sg U46328 ( .A(n30374), .B(n30375), .X(n42036) );
  nand_x1_sg U46329 ( .A(n30372), .B(n30373), .X(n42035) );
  nand_x1_sg U46330 ( .A(n30356), .B(n30357), .X(n42027) );
  nand_x1_sg U46331 ( .A(n30354), .B(n30355), .X(n42026) );
  nand_x1_sg U46332 ( .A(n30362), .B(n30363), .X(n42030) );
  nand_x1_sg U46333 ( .A(n30360), .B(n30361), .X(n42029) );
  nand_x1_sg U46334 ( .A(n30488), .B(n30489), .X(n42093) );
  nand_x1_sg U46335 ( .A(n30486), .B(n30487), .X(n42092) );
  nand_x1_sg U46336 ( .A(n30494), .B(n30495), .X(n42096) );
  nand_x1_sg U46337 ( .A(n30492), .B(n30493), .X(n42095) );
  nand_x1_sg U46338 ( .A(n30476), .B(n30477), .X(n42087) );
  nand_x1_sg U46339 ( .A(n30474), .B(n30475), .X(n42086) );
  nand_x1_sg U46340 ( .A(n30482), .B(n30483), .X(n42090) );
  nand_x1_sg U46341 ( .A(n30480), .B(n30481), .X(n42089) );
  nand_x1_sg U46342 ( .A(n30512), .B(n30513), .X(n42105) );
  nand_x1_sg U46343 ( .A(n30510), .B(n30511), .X(n42104) );
  nand_x1_sg U46344 ( .A(n30518), .B(n30519), .X(n42108) );
  nand_x1_sg U46345 ( .A(n30516), .B(n30517), .X(n42107) );
  nand_x1_sg U46346 ( .A(n30500), .B(n30501), .X(n42099) );
  nand_x1_sg U46347 ( .A(n30498), .B(n30499), .X(n42098) );
  nand_x1_sg U46348 ( .A(n30506), .B(n30507), .X(n42102) );
  nand_x1_sg U46349 ( .A(n30504), .B(n30505), .X(n42101) );
  nand_x1_sg U46350 ( .A(n30440), .B(n30441), .X(n42069) );
  nand_x1_sg U46351 ( .A(n30438), .B(n30439), .X(n42068) );
  nand_x1_sg U46352 ( .A(n30446), .B(n30447), .X(n42072) );
  nand_x1_sg U46353 ( .A(n30444), .B(n30445), .X(n42071) );
  nand_x1_sg U46354 ( .A(n30428), .B(n30429), .X(n42063) );
  nand_x1_sg U46355 ( .A(n30426), .B(n30427), .X(n42062) );
  nand_x1_sg U46356 ( .A(n30434), .B(n30435), .X(n42066) );
  nand_x1_sg U46357 ( .A(n30432), .B(n30433), .X(n42065) );
  nand_x1_sg U46358 ( .A(n30464), .B(n30465), .X(n42081) );
  nand_x1_sg U46359 ( .A(n30462), .B(n30463), .X(n42080) );
  nand_x1_sg U46360 ( .A(n30470), .B(n30471), .X(n42084) );
  nand_x1_sg U46361 ( .A(n30468), .B(n30469), .X(n42083) );
  nand_x1_sg U46362 ( .A(n30452), .B(n30453), .X(n42075) );
  nand_x1_sg U46363 ( .A(n30450), .B(n30451), .X(n42074) );
  nand_x1_sg U46364 ( .A(n30458), .B(n30459), .X(n42078) );
  nand_x1_sg U46365 ( .A(n30456), .B(n30457), .X(n42077) );
  nand_x1_sg U46366 ( .A(n30200), .B(n30201), .X(n41949) );
  nand_x1_sg U46367 ( .A(n30198), .B(n30199), .X(n41948) );
  nand_x1_sg U46368 ( .A(n30206), .B(n30207), .X(n41952) );
  nand_x1_sg U46369 ( .A(n30204), .B(n30205), .X(n41951) );
  nand_x1_sg U46370 ( .A(n30188), .B(n30189), .X(n41943) );
  nand_x1_sg U46371 ( .A(n30186), .B(n30187), .X(n41942) );
  nand_x1_sg U46372 ( .A(n30194), .B(n30195), .X(n41946) );
  nand_x1_sg U46373 ( .A(n30192), .B(n30193), .X(n41945) );
  nand_x1_sg U46374 ( .A(n30224), .B(n30225), .X(n41961) );
  nand_x1_sg U46375 ( .A(n30222), .B(n30223), .X(n41960) );
  nand_x1_sg U46376 ( .A(n30230), .B(n30231), .X(n41964) );
  nand_x1_sg U46377 ( .A(n30228), .B(n30229), .X(n41963) );
  nand_x1_sg U46378 ( .A(n30212), .B(n30213), .X(n41955) );
  nand_x1_sg U46379 ( .A(n30210), .B(n30211), .X(n41954) );
  nand_x1_sg U46380 ( .A(n30218), .B(n30219), .X(n41958) );
  nand_x1_sg U46381 ( .A(n30216), .B(n30217), .X(n41957) );
  nand_x1_sg U46382 ( .A(n30152), .B(n30153), .X(n41925) );
  nand_x1_sg U46383 ( .A(n30150), .B(n30151), .X(n41924) );
  nand_x1_sg U46384 ( .A(n30158), .B(n30159), .X(n41928) );
  nand_x1_sg U46385 ( .A(n30156), .B(n30157), .X(n41927) );
  nand_x1_sg U46386 ( .A(n30140), .B(n30141), .X(n41919) );
  nand_x1_sg U46387 ( .A(n30138), .B(n30139), .X(n41918) );
  nand_x1_sg U46388 ( .A(n30146), .B(n30147), .X(n41922) );
  nand_x1_sg U46389 ( .A(n30144), .B(n30145), .X(n41921) );
  nand_x1_sg U46390 ( .A(n30176), .B(n30177), .X(n41937) );
  nand_x1_sg U46391 ( .A(n30174), .B(n30175), .X(n41936) );
  nand_x1_sg U46392 ( .A(n30182), .B(n30183), .X(n41940) );
  nand_x1_sg U46393 ( .A(n30180), .B(n30181), .X(n41939) );
  nand_x1_sg U46394 ( .A(n30164), .B(n30165), .X(n41931) );
  nand_x1_sg U46395 ( .A(n30162), .B(n30163), .X(n41930) );
  nand_x1_sg U46396 ( .A(n30170), .B(n30171), .X(n41934) );
  nand_x1_sg U46397 ( .A(n30168), .B(n30169), .X(n41933) );
  nand_x1_sg U46398 ( .A(n30296), .B(n30297), .X(n41997) );
  nand_x1_sg U46399 ( .A(n30294), .B(n30295), .X(n41996) );
  nand_x1_sg U46400 ( .A(n30302), .B(n30303), .X(n42000) );
  nand_x1_sg U46401 ( .A(n30300), .B(n30301), .X(n41999) );
  nand_x1_sg U46402 ( .A(n30284), .B(n30285), .X(n41991) );
  nand_x1_sg U46403 ( .A(n30282), .B(n30283), .X(n41990) );
  nand_x1_sg U46404 ( .A(n30290), .B(n30291), .X(n41994) );
  nand_x1_sg U46405 ( .A(n30288), .B(n30289), .X(n41993) );
  nand_x1_sg U46406 ( .A(n30320), .B(n30321), .X(n42009) );
  nand_x1_sg U46407 ( .A(n30318), .B(n30319), .X(n42008) );
  nand_x1_sg U46408 ( .A(n30326), .B(n30327), .X(n42012) );
  nand_x1_sg U46409 ( .A(n30324), .B(n30325), .X(n42011) );
  nand_x1_sg U46410 ( .A(n30308), .B(n30309), .X(n42003) );
  nand_x1_sg U46411 ( .A(n30306), .B(n30307), .X(n42002) );
  nand_x1_sg U46412 ( .A(n30314), .B(n30315), .X(n42006) );
  nand_x1_sg U46413 ( .A(n30312), .B(n30313), .X(n42005) );
  nand_x1_sg U46414 ( .A(n30248), .B(n30249), .X(n41973) );
  nand_x1_sg U46415 ( .A(n30246), .B(n30247), .X(n41972) );
  nand_x1_sg U46416 ( .A(n30254), .B(n30255), .X(n41976) );
  nand_x1_sg U46417 ( .A(n30252), .B(n30253), .X(n41975) );
  nand_x1_sg U46418 ( .A(n30236), .B(n30237), .X(n41967) );
  nand_x1_sg U46419 ( .A(n30234), .B(n30235), .X(n41966) );
  nand_x1_sg U46420 ( .A(n30242), .B(n30243), .X(n41970) );
  nand_x1_sg U46421 ( .A(n30240), .B(n30241), .X(n41969) );
  nand_x1_sg U46422 ( .A(n30272), .B(n30273), .X(n41985) );
  nand_x1_sg U46423 ( .A(n30270), .B(n30271), .X(n41984) );
  nand_x1_sg U46424 ( .A(n30278), .B(n30279), .X(n41988) );
  nand_x1_sg U46425 ( .A(n30276), .B(n30277), .X(n41987) );
  nand_x1_sg U46426 ( .A(n30260), .B(n30261), .X(n41979) );
  nand_x1_sg U46427 ( .A(n30258), .B(n30259), .X(n41978) );
  nand_x1_sg U46428 ( .A(n30266), .B(n30267), .X(n41982) );
  nand_x1_sg U46429 ( .A(n30264), .B(n30265), .X(n41981) );
  nand_x1_sg U46430 ( .A(n30592), .B(n30593), .X(n42145) );
  nand_x1_sg U46431 ( .A(n30590), .B(n30591), .X(n42144) );
  nand_x1_sg U46432 ( .A(n30598), .B(n30599), .X(n42148) );
  nand_x1_sg U46433 ( .A(n30596), .B(n30597), .X(n42147) );
  nand_x1_sg U46434 ( .A(n30580), .B(n30581), .X(n42139) );
  nand_x1_sg U46435 ( .A(n30578), .B(n30579), .X(n42138) );
  nand_x1_sg U46436 ( .A(n30586), .B(n30587), .X(n42142) );
  nand_x1_sg U46437 ( .A(n30584), .B(n30585), .X(n42141) );
  nand_x1_sg U46438 ( .A(n30616), .B(n30617), .X(n42157) );
  nand_x1_sg U46439 ( .A(n30614), .B(n30615), .X(n42156) );
  nand_x1_sg U46440 ( .A(n30622), .B(n30623), .X(n42160) );
  nand_x1_sg U46441 ( .A(n30620), .B(n30621), .X(n42159) );
  nand_x1_sg U46442 ( .A(n30604), .B(n30605), .X(n42151) );
  nand_x1_sg U46443 ( .A(n30602), .B(n30603), .X(n42150) );
  nand_x1_sg U46444 ( .A(n30610), .B(n30611), .X(n42154) );
  nand_x1_sg U46445 ( .A(n30608), .B(n30609), .X(n42153) );
  nand_x1_sg U46446 ( .A(n30544), .B(n30545), .X(n42121) );
  nand_x1_sg U46447 ( .A(n30542), .B(n30543), .X(n42120) );
  nand_x1_sg U46448 ( .A(n30550), .B(n30551), .X(n42124) );
  nand_x1_sg U46449 ( .A(n30548), .B(n30549), .X(n42123) );
  nand_x1_sg U46450 ( .A(n30532), .B(n30533), .X(n42115) );
  nand_x1_sg U46451 ( .A(n30530), .B(n30531), .X(n42114) );
  nand_x1_sg U46452 ( .A(n30538), .B(n30539), .X(n42118) );
  nand_x1_sg U46453 ( .A(n30536), .B(n30537), .X(n42117) );
  nand_x1_sg U46454 ( .A(n30568), .B(n30569), .X(n42133) );
  nand_x1_sg U46455 ( .A(n30566), .B(n30567), .X(n42132) );
  nand_x1_sg U46456 ( .A(n30574), .B(n30575), .X(n42136) );
  nand_x1_sg U46457 ( .A(n30572), .B(n30573), .X(n42135) );
  nand_x1_sg U46458 ( .A(n30556), .B(n30557), .X(n42127) );
  nand_x1_sg U46459 ( .A(n30554), .B(n30555), .X(n42126) );
  nand_x1_sg U46460 ( .A(n30562), .B(n30563), .X(n42130) );
  nand_x1_sg U46461 ( .A(n30560), .B(n30561), .X(n42129) );
  nand_x1_sg U46462 ( .A(n30262), .B(n30263), .X(n41980) );
  nand_x1_sg U46463 ( .A(n30136), .B(n30137), .X(n41917) );
  nand_x1_sg U46464 ( .A(n30564), .B(n30565), .X(n42131) );
  nand_x1_sg U46465 ( .A(n30558), .B(n30559), .X(n42128) );
  nand_x1_sg U46466 ( .A(n30226), .B(n30227), .X(n41962) );
  nand_x1_sg U46467 ( .A(n29748), .B(n29749), .X(n41723) );
  nand_x1_sg U46468 ( .A(n30600), .B(n30601), .X(n42149) );
  nand_x1_sg U46469 ( .A(n30134), .B(n30135), .X(n41916) );
  nand_x1_sg U46470 ( .A(n30520), .B(n30521), .X(n42109) );
  nand_x1_sg U46471 ( .A(n30528), .B(n30529), .X(n42113) );
  nand_x1_sg U46472 ( .A(n30570), .B(n30571), .X(n42134) );
  nand_x1_sg U46473 ( .A(n30400), .B(n30401), .X(n42049) );
  nand_x1_sg U46474 ( .A(n57874), .B(n29326), .X(\shifter_0/n14056 ) );
  nand_x1_sg U46475 ( .A(n32434), .B(n32435), .X(n42814) );
  nand_x1_sg U46476 ( .A(n57302), .B(n32368), .X(n32435) );
  nand_x1_sg U46477 ( .A(n32379), .B(n32380), .X(n42812) );
  nand_x1_sg U46478 ( .A(n57304), .B(n32368), .X(n32380) );
  nand_x1_sg U46479 ( .A(n32366), .B(n32367), .X(n42811) );
  nand_x1_sg U46480 ( .A(n32389), .B(n32390), .X(n42813) );
  nand_x1_sg U46481 ( .A(n68264), .B(n32391), .X(n32390) );
  nand_x1_sg U46482 ( .A(n57306), .B(n32368), .X(n32389) );
  nand_x1_sg U46483 ( .A(n32392), .B(n32393), .X(n32391) );
  nand_x1_sg U46484 ( .A(n58759), .B(n58758), .X(n42355) );
  inv_x1_sg U46485 ( .A(n58757), .X(n58758) );
  inv_x1_sg U46486 ( .A(n58756), .X(n58759) );
  nand_x1_sg U46487 ( .A(n58754), .B(n58753), .X(n42354) );
  inv_x1_sg U46488 ( .A(n58752), .X(n58753) );
  inv_x1_sg U46489 ( .A(n58751), .X(n58754) );
  nand_x1_sg U46490 ( .A(n58749), .B(n58748), .X(n42358) );
  inv_x1_sg U46491 ( .A(n58747), .X(n58748) );
  inv_x1_sg U46492 ( .A(n58746), .X(n58749) );
  nand_x1_sg U46493 ( .A(n58744), .B(n58743), .X(n42357) );
  inv_x1_sg U46494 ( .A(n58742), .X(n58743) );
  inv_x1_sg U46495 ( .A(n58741), .X(n58744) );
  nand_x1_sg U46496 ( .A(n58739), .B(n58738), .X(n42349) );
  inv_x1_sg U46497 ( .A(n58737), .X(n58738) );
  inv_x1_sg U46498 ( .A(n58736), .X(n58739) );
  nand_x1_sg U46499 ( .A(n58734), .B(n58733), .X(n42348) );
  inv_x1_sg U46500 ( .A(n58732), .X(n58733) );
  inv_x1_sg U46501 ( .A(n58731), .X(n58734) );
  nand_x1_sg U46502 ( .A(n58729), .B(n58728), .X(n42352) );
  inv_x1_sg U46503 ( .A(n58727), .X(n58728) );
  inv_x1_sg U46504 ( .A(n58726), .X(n58729) );
  nand_x1_sg U46505 ( .A(n58724), .B(n58723), .X(n42351) );
  inv_x1_sg U46506 ( .A(n58722), .X(n58723) );
  inv_x1_sg U46507 ( .A(n58721), .X(n58724) );
  nand_x1_sg U46508 ( .A(n58719), .B(n58718), .X(n42367) );
  inv_x1_sg U46509 ( .A(n58717), .X(n58718) );
  inv_x1_sg U46510 ( .A(n58716), .X(n58719) );
  nand_x1_sg U46511 ( .A(n58714), .B(n58713), .X(n42366) );
  inv_x1_sg U46512 ( .A(n58712), .X(n58713) );
  inv_x1_sg U46513 ( .A(n58711), .X(n58714) );
  nand_x1_sg U46514 ( .A(n58709), .B(n58708), .X(n42370) );
  inv_x1_sg U46515 ( .A(n58707), .X(n58708) );
  inv_x1_sg U46516 ( .A(n58706), .X(n58709) );
  nand_x1_sg U46517 ( .A(n58704), .B(n58703), .X(n42369) );
  inv_x1_sg U46518 ( .A(n58702), .X(n58703) );
  inv_x1_sg U46519 ( .A(n58701), .X(n58704) );
  nand_x1_sg U46520 ( .A(n58699), .B(n58698), .X(n42361) );
  inv_x1_sg U46521 ( .A(n58697), .X(n58698) );
  inv_x1_sg U46522 ( .A(n58696), .X(n58699) );
  nand_x1_sg U46523 ( .A(n58694), .B(n58693), .X(n42360) );
  inv_x1_sg U46524 ( .A(n58692), .X(n58693) );
  inv_x1_sg U46525 ( .A(n58691), .X(n58694) );
  nand_x1_sg U46526 ( .A(n58689), .B(n58688), .X(n42364) );
  inv_x1_sg U46527 ( .A(n58687), .X(n58688) );
  inv_x1_sg U46528 ( .A(n58686), .X(n58689) );
  nand_x1_sg U46529 ( .A(n58684), .B(n58683), .X(n42363) );
  inv_x1_sg U46530 ( .A(n58682), .X(n58683) );
  inv_x1_sg U46531 ( .A(n58681), .X(n58684) );
  nand_x1_sg U46532 ( .A(n58679), .B(n58678), .X(n42331) );
  inv_x1_sg U46533 ( .A(n58677), .X(n58678) );
  inv_x1_sg U46534 ( .A(n58676), .X(n58679) );
  nand_x1_sg U46535 ( .A(n58674), .B(n58673), .X(n42330) );
  inv_x1_sg U46536 ( .A(n58672), .X(n58673) );
  inv_x1_sg U46537 ( .A(n58671), .X(n58674) );
  nand_x1_sg U46538 ( .A(n58669), .B(n58668), .X(n42334) );
  inv_x1_sg U46539 ( .A(n58667), .X(n58668) );
  inv_x1_sg U46540 ( .A(n58666), .X(n58669) );
  nand_x1_sg U46541 ( .A(n58664), .B(n58663), .X(n42333) );
  inv_x1_sg U46542 ( .A(n58662), .X(n58663) );
  inv_x1_sg U46543 ( .A(n58661), .X(n58664) );
  nand_x1_sg U46544 ( .A(n61861), .B(n61860), .X(n42769) );
  inv_x1_sg U46545 ( .A(n61859), .X(n61860) );
  inv_x1_sg U46546 ( .A(n61857), .X(n61861) );
  nand_x1_sg U46547 ( .A(n61854), .B(n61853), .X(n42766) );
  inv_x1_sg U46548 ( .A(n61852), .X(n61853) );
  inv_x1_sg U46549 ( .A(n61851), .X(n61854) );
  nand_x1_sg U46550 ( .A(n61849), .B(n61848), .X(n42230) );
  inv_x1_sg U46551 ( .A(n61847), .X(n61848) );
  inv_x1_sg U46552 ( .A(n61846), .X(n61849) );
  nand_x1_sg U46553 ( .A(n61844), .B(n61843), .X(n42229) );
  inv_x1_sg U46554 ( .A(n61842), .X(n61843) );
  inv_x1_sg U46555 ( .A(n61841), .X(n61844) );
  nand_x1_sg U46556 ( .A(n61839), .B(n61838), .X(n42343) );
  inv_x1_sg U46557 ( .A(n61837), .X(n61838) );
  inv_x1_sg U46558 ( .A(n61836), .X(n61839) );
  nand_x1_sg U46559 ( .A(n61834), .B(n61833), .X(n42342) );
  inv_x1_sg U46560 ( .A(n61832), .X(n61833) );
  inv_x1_sg U46561 ( .A(n61831), .X(n61834) );
  nand_x1_sg U46562 ( .A(n61829), .B(n61828), .X(n42346) );
  inv_x1_sg U46563 ( .A(n61827), .X(n61828) );
  inv_x1_sg U46564 ( .A(n61826), .X(n61829) );
  nand_x1_sg U46565 ( .A(n61824), .B(n61823), .X(n42345) );
  inv_x1_sg U46566 ( .A(n61822), .X(n61823) );
  inv_x1_sg U46567 ( .A(n61821), .X(n61824) );
  nand_x1_sg U46568 ( .A(n61819), .B(n61818), .X(n42337) );
  inv_x1_sg U46569 ( .A(n61817), .X(n61818) );
  inv_x1_sg U46570 ( .A(n61816), .X(n61819) );
  nand_x1_sg U46571 ( .A(n61814), .B(n61813), .X(n42336) );
  inv_x1_sg U46572 ( .A(n61812), .X(n61813) );
  inv_x1_sg U46573 ( .A(n61811), .X(n61814) );
  nand_x1_sg U46574 ( .A(n61809), .B(n61808), .X(n42340) );
  inv_x1_sg U46575 ( .A(n61807), .X(n61808) );
  inv_x1_sg U46576 ( .A(n61806), .X(n61809) );
  nand_x1_sg U46577 ( .A(n61804), .B(n61803), .X(n42339) );
  inv_x1_sg U46578 ( .A(n61802), .X(n61803) );
  inv_x1_sg U46579 ( .A(n61801), .X(n61804) );
  nand_x1_sg U46580 ( .A(n61799), .B(n61798), .X(n42403) );
  inv_x1_sg U46581 ( .A(n61797), .X(n61798) );
  inv_x1_sg U46582 ( .A(n61796), .X(n61799) );
  nand_x1_sg U46583 ( .A(n61794), .B(n61793), .X(n42402) );
  inv_x1_sg U46584 ( .A(n61792), .X(n61793) );
  inv_x1_sg U46585 ( .A(n61791), .X(n61794) );
  nand_x1_sg U46586 ( .A(n61789), .B(n61788), .X(n42406) );
  inv_x1_sg U46587 ( .A(n61787), .X(n61788) );
  inv_x1_sg U46588 ( .A(n61786), .X(n61789) );
  nand_x1_sg U46589 ( .A(n61784), .B(n61783), .X(n42405) );
  inv_x1_sg U46590 ( .A(n61782), .X(n61783) );
  inv_x1_sg U46591 ( .A(n61781), .X(n61784) );
  nand_x1_sg U46592 ( .A(n61779), .B(n61778), .X(n42397) );
  inv_x1_sg U46593 ( .A(n61777), .X(n61778) );
  inv_x1_sg U46594 ( .A(n61776), .X(n61779) );
  nand_x1_sg U46595 ( .A(n61774), .B(n61773), .X(n42396) );
  inv_x1_sg U46596 ( .A(n61772), .X(n61773) );
  inv_x1_sg U46597 ( .A(n61771), .X(n61774) );
  nand_x1_sg U46598 ( .A(n61769), .B(n61768), .X(n42400) );
  inv_x1_sg U46599 ( .A(n61767), .X(n61768) );
  inv_x1_sg U46600 ( .A(n61766), .X(n61769) );
  nand_x1_sg U46601 ( .A(n61764), .B(n61763), .X(n42399) );
  inv_x1_sg U46602 ( .A(n61762), .X(n61763) );
  inv_x1_sg U46603 ( .A(n61761), .X(n61764) );
  nand_x1_sg U46604 ( .A(n61759), .B(n61758), .X(n42784) );
  inv_x1_sg U46605 ( .A(n61757), .X(n61758) );
  inv_x1_sg U46606 ( .A(n61756), .X(n61759) );
  nand_x1_sg U46607 ( .A(n61754), .B(n61753), .X(n42781) );
  inv_x1_sg U46608 ( .A(n61752), .X(n61753) );
  inv_x1_sg U46609 ( .A(n61751), .X(n61754) );
  nand_x1_sg U46610 ( .A(n61749), .B(n61748), .X(n42778) );
  inv_x1_sg U46611 ( .A(n61747), .X(n61748) );
  inv_x1_sg U46612 ( .A(n61746), .X(n61749) );
  nand_x1_sg U46613 ( .A(n61744), .B(n61743), .X(n42775) );
  inv_x1_sg U46614 ( .A(n61742), .X(n61743) );
  inv_x1_sg U46615 ( .A(n61741), .X(n61744) );
  nand_x1_sg U46616 ( .A(n61739), .B(n61738), .X(n42410) );
  inv_x1_sg U46617 ( .A(n61737), .X(n61738) );
  inv_x1_sg U46618 ( .A(n61736), .X(n61739) );
  nand_x1_sg U46619 ( .A(n61734), .B(n61733), .X(n42409) );
  inv_x1_sg U46620 ( .A(n61732), .X(n61733) );
  inv_x1_sg U46621 ( .A(n61731), .X(n61734) );
  nand_x1_sg U46622 ( .A(n61729), .B(n61728), .X(n42413) );
  inv_x1_sg U46623 ( .A(n61727), .X(n61728) );
  inv_x1_sg U46624 ( .A(n61726), .X(n61729) );
  nand_x1_sg U46625 ( .A(n61724), .B(n61723), .X(n42412) );
  inv_x1_sg U46626 ( .A(n61722), .X(n61723) );
  inv_x1_sg U46627 ( .A(n61721), .X(n61724) );
  nand_x1_sg U46628 ( .A(n61719), .B(n61718), .X(n42379) );
  inv_x1_sg U46629 ( .A(n61717), .X(n61718) );
  inv_x1_sg U46630 ( .A(n61716), .X(n61719) );
  nand_x1_sg U46631 ( .A(n61714), .B(n61713), .X(n42378) );
  inv_x1_sg U46632 ( .A(n61712), .X(n61713) );
  inv_x1_sg U46633 ( .A(n61711), .X(n61714) );
  nand_x1_sg U46634 ( .A(n61709), .B(n61708), .X(n42382) );
  inv_x1_sg U46635 ( .A(n61707), .X(n61708) );
  inv_x1_sg U46636 ( .A(n61706), .X(n61709) );
  nand_x1_sg U46637 ( .A(n61704), .B(n61703), .X(n42381) );
  inv_x1_sg U46638 ( .A(n61702), .X(n61703) );
  inv_x1_sg U46639 ( .A(n61701), .X(n61704) );
  nand_x1_sg U46640 ( .A(n61699), .B(n61698), .X(n42373) );
  inv_x1_sg U46641 ( .A(n61697), .X(n61698) );
  inv_x1_sg U46642 ( .A(n61696), .X(n61699) );
  nand_x1_sg U46643 ( .A(n61694), .B(n61693), .X(n42372) );
  inv_x1_sg U46644 ( .A(n61692), .X(n61693) );
  inv_x1_sg U46645 ( .A(n61691), .X(n61694) );
  nand_x1_sg U46646 ( .A(n61689), .B(n61688), .X(n42376) );
  inv_x1_sg U46647 ( .A(n61687), .X(n61688) );
  inv_x1_sg U46648 ( .A(n61686), .X(n61689) );
  nand_x1_sg U46649 ( .A(n61684), .B(n61683), .X(n42375) );
  inv_x1_sg U46650 ( .A(n61682), .X(n61683) );
  inv_x1_sg U46651 ( .A(n61681), .X(n61684) );
  nand_x1_sg U46652 ( .A(n61679), .B(n61678), .X(n42391) );
  inv_x1_sg U46653 ( .A(n61677), .X(n61678) );
  inv_x1_sg U46654 ( .A(n61676), .X(n61679) );
  nand_x1_sg U46655 ( .A(n61674), .B(n61673), .X(n42390) );
  inv_x1_sg U46656 ( .A(n61672), .X(n61673) );
  inv_x1_sg U46657 ( .A(n61671), .X(n61674) );
  nand_x1_sg U46658 ( .A(n61669), .B(n61668), .X(n42394) );
  inv_x1_sg U46659 ( .A(n61667), .X(n61668) );
  inv_x1_sg U46660 ( .A(n61666), .X(n61669) );
  nand_x1_sg U46661 ( .A(n61664), .B(n61663), .X(n42393) );
  inv_x1_sg U46662 ( .A(n61662), .X(n61663) );
  inv_x1_sg U46663 ( .A(n61661), .X(n61664) );
  nand_x1_sg U46664 ( .A(n61659), .B(n61658), .X(n42385) );
  inv_x1_sg U46665 ( .A(n61657), .X(n61658) );
  inv_x1_sg U46666 ( .A(n61656), .X(n61659) );
  nand_x1_sg U46667 ( .A(n61654), .B(n61653), .X(n42384) );
  inv_x1_sg U46668 ( .A(n61652), .X(n61653) );
  inv_x1_sg U46669 ( .A(n61651), .X(n61654) );
  nand_x1_sg U46670 ( .A(n61649), .B(n61648), .X(n42388) );
  inv_x1_sg U46671 ( .A(n61647), .X(n61648) );
  inv_x1_sg U46672 ( .A(n61646), .X(n61649) );
  nand_x1_sg U46673 ( .A(n61644), .B(n61643), .X(n42387) );
  inv_x1_sg U46674 ( .A(n61642), .X(n61643) );
  inv_x1_sg U46675 ( .A(n61641), .X(n61644) );
  nand_x1_sg U46676 ( .A(n61639), .B(n61638), .X(n42292) );
  inv_x1_sg U46677 ( .A(n61637), .X(n61638) );
  inv_x1_sg U46678 ( .A(n61636), .X(n61639) );
  nand_x1_sg U46679 ( .A(n61634), .B(n61633), .X(n42291) );
  inv_x1_sg U46680 ( .A(n61632), .X(n61633) );
  inv_x1_sg U46681 ( .A(n61631), .X(n61634) );
  nand_x1_sg U46682 ( .A(n61629), .B(n61628), .X(n42295) );
  inv_x1_sg U46683 ( .A(n61627), .X(n61628) );
  inv_x1_sg U46684 ( .A(n61626), .X(n61629) );
  nand_x1_sg U46685 ( .A(n61624), .B(n61623), .X(n42294) );
  inv_x1_sg U46686 ( .A(n61622), .X(n61623) );
  inv_x1_sg U46687 ( .A(n61621), .X(n61624) );
  nand_x1_sg U46688 ( .A(n61619), .B(n61618), .X(n42286) );
  inv_x1_sg U46689 ( .A(n61617), .X(n61618) );
  inv_x1_sg U46690 ( .A(n61616), .X(n61619) );
  nand_x1_sg U46691 ( .A(n61614), .B(n61613), .X(n42285) );
  inv_x1_sg U46692 ( .A(n61612), .X(n61613) );
  inv_x1_sg U46693 ( .A(n61611), .X(n61614) );
  nand_x1_sg U46694 ( .A(n61609), .B(n61608), .X(n42289) );
  inv_x1_sg U46695 ( .A(n61607), .X(n61608) );
  inv_x1_sg U46696 ( .A(n61606), .X(n61609) );
  nand_x1_sg U46697 ( .A(n61604), .B(n61603), .X(n42288) );
  inv_x1_sg U46698 ( .A(n61602), .X(n61603) );
  inv_x1_sg U46699 ( .A(n61601), .X(n61604) );
  nand_x1_sg U46700 ( .A(n61599), .B(n61598), .X(n42304) );
  inv_x1_sg U46701 ( .A(n61597), .X(n61598) );
  inv_x1_sg U46702 ( .A(n61596), .X(n61599) );
  nand_x1_sg U46703 ( .A(n61594), .B(n61593), .X(n42303) );
  inv_x1_sg U46704 ( .A(n61592), .X(n61593) );
  inv_x1_sg U46705 ( .A(n61591), .X(n61594) );
  nand_x1_sg U46706 ( .A(n61589), .B(n61588), .X(n42307) );
  inv_x1_sg U46707 ( .A(n61587), .X(n61588) );
  inv_x1_sg U46708 ( .A(n61586), .X(n61589) );
  nand_x1_sg U46709 ( .A(n61584), .B(n61583), .X(n42306) );
  inv_x1_sg U46710 ( .A(n61582), .X(n61583) );
  inv_x1_sg U46711 ( .A(n61581), .X(n61584) );
  nand_x1_sg U46712 ( .A(n61579), .B(n61578), .X(n42298) );
  inv_x1_sg U46713 ( .A(n61577), .X(n61578) );
  inv_x1_sg U46714 ( .A(n61576), .X(n61579) );
  nand_x1_sg U46715 ( .A(n61574), .B(n61573), .X(n42297) );
  inv_x1_sg U46716 ( .A(n61572), .X(n61573) );
  inv_x1_sg U46717 ( .A(n61571), .X(n61574) );
  nand_x1_sg U46718 ( .A(n61569), .B(n61568), .X(n42301) );
  inv_x1_sg U46719 ( .A(n61567), .X(n61568) );
  inv_x1_sg U46720 ( .A(n61566), .X(n61569) );
  nand_x1_sg U46721 ( .A(n61564), .B(n61563), .X(n42300) );
  inv_x1_sg U46722 ( .A(n61562), .X(n61563) );
  inv_x1_sg U46723 ( .A(n61561), .X(n61564) );
  nand_x1_sg U46724 ( .A(n61559), .B(n61558), .X(n42268) );
  inv_x1_sg U46725 ( .A(n61557), .X(n61558) );
  inv_x1_sg U46726 ( .A(n61556), .X(n61559) );
  nand_x1_sg U46727 ( .A(n61554), .B(n61553), .X(n42267) );
  inv_x1_sg U46728 ( .A(n61552), .X(n61553) );
  inv_x1_sg U46729 ( .A(n61551), .X(n61554) );
  nand_x1_sg U46730 ( .A(n61549), .B(n61548), .X(n42271) );
  inv_x1_sg U46731 ( .A(n61547), .X(n61548) );
  inv_x1_sg U46732 ( .A(n61546), .X(n61549) );
  nand_x1_sg U46733 ( .A(n61544), .B(n61543), .X(n42270) );
  inv_x1_sg U46734 ( .A(n61542), .X(n61543) );
  inv_x1_sg U46735 ( .A(n61541), .X(n61544) );
  nand_x1_sg U46736 ( .A(n61539), .B(n61538), .X(n42262) );
  inv_x1_sg U46737 ( .A(n61537), .X(n61538) );
  inv_x1_sg U46738 ( .A(n61536), .X(n61539) );
  nand_x1_sg U46739 ( .A(n61534), .B(n61533), .X(n42261) );
  inv_x1_sg U46740 ( .A(n61532), .X(n61533) );
  inv_x1_sg U46741 ( .A(n61531), .X(n61534) );
  nand_x1_sg U46742 ( .A(n61529), .B(n61528), .X(n42265) );
  inv_x1_sg U46743 ( .A(n61527), .X(n61528) );
  inv_x1_sg U46744 ( .A(n61526), .X(n61529) );
  nand_x1_sg U46745 ( .A(n61524), .B(n61523), .X(n42264) );
  inv_x1_sg U46746 ( .A(n61522), .X(n61523) );
  inv_x1_sg U46747 ( .A(n61521), .X(n61524) );
  nand_x1_sg U46748 ( .A(n61519), .B(n61518), .X(n42280) );
  inv_x1_sg U46749 ( .A(n61517), .X(n61518) );
  inv_x1_sg U46750 ( .A(n61516), .X(n61519) );
  nand_x1_sg U46751 ( .A(n61514), .B(n61513), .X(n42279) );
  inv_x1_sg U46752 ( .A(n61512), .X(n61513) );
  inv_x1_sg U46753 ( .A(n61511), .X(n61514) );
  nand_x1_sg U46754 ( .A(n61509), .B(n61508), .X(n42283) );
  inv_x1_sg U46755 ( .A(n61507), .X(n61508) );
  inv_x1_sg U46756 ( .A(n61506), .X(n61509) );
  nand_x1_sg U46757 ( .A(n61504), .B(n61503), .X(n42282) );
  inv_x1_sg U46758 ( .A(n61502), .X(n61503) );
  inv_x1_sg U46759 ( .A(n61501), .X(n61504) );
  nand_x1_sg U46760 ( .A(n61499), .B(n61498), .X(n42274) );
  inv_x1_sg U46761 ( .A(n61497), .X(n61498) );
  inv_x1_sg U46762 ( .A(n61496), .X(n61499) );
  nand_x1_sg U46763 ( .A(n61494), .B(n61493), .X(n42273) );
  inv_x1_sg U46764 ( .A(n61492), .X(n61493) );
  inv_x1_sg U46765 ( .A(n61491), .X(n61494) );
  nand_x1_sg U46766 ( .A(n61489), .B(n61488), .X(n42277) );
  inv_x1_sg U46767 ( .A(n61487), .X(n61488) );
  inv_x1_sg U46768 ( .A(n61486), .X(n61489) );
  nand_x1_sg U46769 ( .A(n61484), .B(n61483), .X(n42276) );
  inv_x1_sg U46770 ( .A(n61482), .X(n61483) );
  inv_x1_sg U46771 ( .A(n61481), .X(n61484) );
  nand_x1_sg U46772 ( .A(n61479), .B(n61478), .X(n42317) );
  inv_x1_sg U46773 ( .A(n61477), .X(n61478) );
  inv_x1_sg U46774 ( .A(n61476), .X(n61479) );
  nand_x1_sg U46775 ( .A(n61474), .B(n61473), .X(n42316) );
  inv_x1_sg U46776 ( .A(n61472), .X(n61473) );
  inv_x1_sg U46777 ( .A(n61471), .X(n61474) );
  nand_x1_sg U46778 ( .A(n61469), .B(n61468), .X(n42320) );
  inv_x1_sg U46779 ( .A(n61467), .X(n61468) );
  inv_x1_sg U46780 ( .A(n61466), .X(n61469) );
  nand_x1_sg U46781 ( .A(n61464), .B(n61463), .X(n42319) );
  inv_x1_sg U46782 ( .A(n61462), .X(n61463) );
  inv_x1_sg U46783 ( .A(n61461), .X(n61464) );
  nand_x1_sg U46784 ( .A(n61459), .B(n61458), .X(n42311) );
  inv_x1_sg U46785 ( .A(n61457), .X(n61458) );
  inv_x1_sg U46786 ( .A(n61456), .X(n61459) );
  nand_x1_sg U46787 ( .A(n61454), .B(n61453), .X(n42310) );
  inv_x1_sg U46788 ( .A(n61452), .X(n61453) );
  inv_x1_sg U46789 ( .A(n61451), .X(n61454) );
  nand_x1_sg U46790 ( .A(n61449), .B(n61448), .X(n42314) );
  inv_x1_sg U46791 ( .A(n61447), .X(n61448) );
  inv_x1_sg U46792 ( .A(n61446), .X(n61449) );
  nand_x1_sg U46793 ( .A(n61444), .B(n61443), .X(n42313) );
  inv_x1_sg U46794 ( .A(n61442), .X(n61443) );
  inv_x1_sg U46795 ( .A(n61441), .X(n61444) );
  nand_x1_sg U46796 ( .A(n61439), .B(n61438), .X(n42324) );
  inv_x1_sg U46797 ( .A(n61437), .X(n61438) );
  inv_x1_sg U46798 ( .A(n61436), .X(n61439) );
  nand_x1_sg U46799 ( .A(n61434), .B(n61433), .X(n42323) );
  inv_x1_sg U46800 ( .A(n61432), .X(n61433) );
  inv_x1_sg U46801 ( .A(n61431), .X(n61434) );
  nand_x1_sg U46802 ( .A(n61429), .B(n61428), .X(n42327) );
  inv_x1_sg U46803 ( .A(n61427), .X(n61428) );
  inv_x1_sg U46804 ( .A(n61426), .X(n61429) );
  nand_x1_sg U46805 ( .A(n61424), .B(n61423), .X(n42326) );
  inv_x1_sg U46806 ( .A(n61422), .X(n61423) );
  inv_x1_sg U46807 ( .A(n61421), .X(n61424) );
  nand_x1_sg U46808 ( .A(n61419), .B(n61418), .X(n42475) );
  inv_x1_sg U46809 ( .A(n61417), .X(n61418) );
  inv_x1_sg U46810 ( .A(n61416), .X(n61419) );
  nand_x1_sg U46811 ( .A(n61414), .B(n61413), .X(n42321) );
  inv_x1_sg U46812 ( .A(n61412), .X(n61413) );
  inv_x1_sg U46813 ( .A(n61411), .X(n61414) );
  nand_x1_sg U46814 ( .A(n61409), .B(n61408), .X(n42472) );
  inv_x1_sg U46815 ( .A(n61407), .X(n61408) );
  inv_x1_sg U46816 ( .A(n61406), .X(n61409) );
  nand_x1_sg U46817 ( .A(n61404), .B(n61403), .X(n42469) );
  inv_x1_sg U46818 ( .A(n61402), .X(n61403) );
  inv_x1_sg U46819 ( .A(n61401), .X(n61404) );
  nand_x1_sg U46820 ( .A(n61399), .B(n61398), .X(n42463) );
  inv_x1_sg U46821 ( .A(n61397), .X(n61398) );
  inv_x1_sg U46822 ( .A(n61396), .X(n61399) );
  nand_x1_sg U46823 ( .A(n61394), .B(n61393), .X(n42308) );
  inv_x1_sg U46824 ( .A(n61392), .X(n61393) );
  inv_x1_sg U46825 ( .A(n61391), .X(n61394) );
  nand_x1_sg U46826 ( .A(n61389), .B(n61388), .X(n42460) );
  inv_x1_sg U46827 ( .A(n61387), .X(n61388) );
  inv_x1_sg U46828 ( .A(n61386), .X(n61389) );
  nand_x1_sg U46829 ( .A(n61384), .B(n61383), .X(n42457) );
  inv_x1_sg U46830 ( .A(n61382), .X(n61383) );
  inv_x1_sg U46831 ( .A(n61381), .X(n61384) );
  nand_x1_sg U46832 ( .A(n61379), .B(n61378), .X(n42454) );
  inv_x1_sg U46833 ( .A(n61377), .X(n61378) );
  inv_x1_sg U46834 ( .A(n61376), .X(n61379) );
  nand_x1_sg U46835 ( .A(n61374), .B(n61373), .X(n42466) );
  inv_x1_sg U46836 ( .A(n61372), .X(n61373) );
  inv_x1_sg U46837 ( .A(n61371), .X(n61374) );
  nand_x1_sg U46838 ( .A(n61369), .B(n61368), .X(n42451) );
  inv_x1_sg U46839 ( .A(n61367), .X(n61368) );
  inv_x1_sg U46840 ( .A(n61366), .X(n61369) );
  nand_x1_sg U46841 ( .A(n61364), .B(n61363), .X(n42448) );
  inv_x1_sg U46842 ( .A(n61362), .X(n61363) );
  inv_x1_sg U46843 ( .A(n61361), .X(n61364) );
  nand_x1_sg U46844 ( .A(n61359), .B(n61358), .X(n42442) );
  inv_x1_sg U46845 ( .A(n61357), .X(n61358) );
  inv_x1_sg U46846 ( .A(n61356), .X(n61359) );
  nand_x1_sg U46847 ( .A(n61354), .B(n61353), .X(n42439) );
  inv_x1_sg U46848 ( .A(n61352), .X(n61353) );
  inv_x1_sg U46849 ( .A(n61351), .X(n61354) );
  nand_x1_sg U46850 ( .A(n61349), .B(n61348), .X(n42436) );
  inv_x1_sg U46851 ( .A(n61347), .X(n61348) );
  inv_x1_sg U46852 ( .A(n61346), .X(n61349) );
  nand_x1_sg U46853 ( .A(n61344), .B(n61343), .X(n42787) );
  inv_x1_sg U46854 ( .A(n61342), .X(n61343) );
  inv_x1_sg U46855 ( .A(n61341), .X(n61344) );
  nand_x1_sg U46856 ( .A(n61339), .B(n61338), .X(n42433) );
  inv_x1_sg U46857 ( .A(n61337), .X(n61338) );
  inv_x1_sg U46858 ( .A(n61336), .X(n61339) );
  nand_x1_sg U46859 ( .A(n61334), .B(n61333), .X(n42445) );
  inv_x1_sg U46860 ( .A(n61332), .X(n61333) );
  inv_x1_sg U46861 ( .A(n61331), .X(n61334) );
  nand_x1_sg U46862 ( .A(n61329), .B(n61328), .X(n42427) );
  inv_x1_sg U46863 ( .A(n61327), .X(n61328) );
  inv_x1_sg U46864 ( .A(n61326), .X(n61329) );
  nand_x1_sg U46865 ( .A(n61324), .B(n61323), .X(n42424) );
  inv_x1_sg U46866 ( .A(n61322), .X(n61323) );
  inv_x1_sg U46867 ( .A(n61321), .X(n61324) );
  nand_x1_sg U46868 ( .A(n61319), .B(n61318), .X(n42613) );
  inv_x1_sg U46869 ( .A(n61317), .X(n61318) );
  inv_x1_sg U46870 ( .A(n61316), .X(n61319) );
  nand_x1_sg U46871 ( .A(n61314), .B(n61313), .X(n42610) );
  inv_x1_sg U46872 ( .A(n61312), .X(n61313) );
  inv_x1_sg U46873 ( .A(n61311), .X(n61314) );
  nand_x1_sg U46874 ( .A(n61309), .B(n61308), .X(n42571) );
  inv_x1_sg U46875 ( .A(n61307), .X(n61308) );
  inv_x1_sg U46876 ( .A(n61306), .X(n61309) );
  nand_x1_sg U46877 ( .A(n61304), .B(n61303), .X(n42649) );
  inv_x1_sg U46878 ( .A(n61302), .X(n61303) );
  inv_x1_sg U46879 ( .A(n61301), .X(n61304) );
  nand_x1_sg U46880 ( .A(n61299), .B(n61298), .X(n42259) );
  inv_x1_sg U46881 ( .A(n61297), .X(n61298) );
  inv_x1_sg U46882 ( .A(n61296), .X(n61299) );
  nand_x1_sg U46883 ( .A(n61294), .B(n61293), .X(n42417) );
  inv_x1_sg U46884 ( .A(n61292), .X(n61293) );
  inv_x1_sg U46885 ( .A(n61291), .X(n61294) );
  nand_x1_sg U46886 ( .A(n61289), .B(n61288), .X(n42258) );
  inv_x1_sg U46887 ( .A(n61287), .X(n61288) );
  inv_x1_sg U46888 ( .A(n61286), .X(n61289) );
  nand_x1_sg U46889 ( .A(n61284), .B(n61283), .X(n42421) );
  inv_x1_sg U46890 ( .A(n61282), .X(n61283) );
  inv_x1_sg U46891 ( .A(n61281), .X(n61284) );
  nand_x1_sg U46892 ( .A(n61279), .B(n61278), .X(n42589) );
  inv_x1_sg U46893 ( .A(n61277), .X(n61278) );
  inv_x1_sg U46894 ( .A(n61276), .X(n61279) );
  nand_x1_sg U46895 ( .A(n61274), .B(n61273), .X(n42586) );
  inv_x1_sg U46896 ( .A(n61272), .X(n61273) );
  inv_x1_sg U46897 ( .A(n61271), .X(n61274) );
  nand_x1_sg U46898 ( .A(n61269), .B(n61268), .X(n42580) );
  inv_x1_sg U46899 ( .A(n61267), .X(n61268) );
  inv_x1_sg U46900 ( .A(n61266), .X(n61269) );
  nand_x1_sg U46901 ( .A(n61264), .B(n61263), .X(n42577) );
  inv_x1_sg U46902 ( .A(n61262), .X(n61263) );
  inv_x1_sg U46903 ( .A(n61261), .X(n61264) );
  nand_x1_sg U46904 ( .A(n61259), .B(n61258), .X(n42607) );
  inv_x1_sg U46905 ( .A(n61257), .X(n61258) );
  inv_x1_sg U46906 ( .A(n61256), .X(n61259) );
  nand_x1_sg U46907 ( .A(n61254), .B(n61253), .X(n42604) );
  inv_x1_sg U46908 ( .A(n61252), .X(n61253) );
  inv_x1_sg U46909 ( .A(n61251), .X(n61254) );
  nand_x1_sg U46910 ( .A(n61249), .B(n61248), .X(n42598) );
  inv_x1_sg U46911 ( .A(n61247), .X(n61248) );
  inv_x1_sg U46912 ( .A(n61246), .X(n61249) );
  nand_x1_sg U46913 ( .A(n61244), .B(n61243), .X(n42595) );
  inv_x1_sg U46914 ( .A(n61242), .X(n61243) );
  inv_x1_sg U46915 ( .A(n61241), .X(n61244) );
  nand_x1_sg U46916 ( .A(n61239), .B(n61238), .X(n42592) );
  inv_x1_sg U46917 ( .A(n61237), .X(n61238) );
  inv_x1_sg U46918 ( .A(n61236), .X(n61239) );
  nand_x1_sg U46919 ( .A(n61234), .B(n61233), .X(n42601) );
  inv_x1_sg U46920 ( .A(n61232), .X(n61233) );
  inv_x1_sg U46921 ( .A(n61231), .X(n61234) );
  nand_x1_sg U46922 ( .A(n61229), .B(n61228), .X(n42658) );
  inv_x1_sg U46923 ( .A(n61227), .X(n61228) );
  inv_x1_sg U46924 ( .A(n61226), .X(n61229) );
  nand_x1_sg U46925 ( .A(n61224), .B(n61223), .X(n42250) );
  inv_x1_sg U46926 ( .A(n61222), .X(n61223) );
  inv_x1_sg U46927 ( .A(n61221), .X(n61224) );
  nand_x1_sg U46928 ( .A(n61219), .B(n61218), .X(n42643) );
  inv_x1_sg U46929 ( .A(n61217), .X(n61218) );
  inv_x1_sg U46930 ( .A(n61216), .X(n61219) );
  nand_x1_sg U46931 ( .A(n61214), .B(n61213), .X(n42631) );
  inv_x1_sg U46932 ( .A(n61212), .X(n61213) );
  inv_x1_sg U46933 ( .A(n61211), .X(n61214) );
  nand_x1_sg U46934 ( .A(n61209), .B(n61208), .X(n42574) );
  inv_x1_sg U46935 ( .A(n61207), .X(n61208) );
  inv_x1_sg U46936 ( .A(n61206), .X(n61209) );
  nand_x1_sg U46937 ( .A(n61204), .B(n61203), .X(n42583) );
  inv_x1_sg U46938 ( .A(n61202), .X(n61203) );
  inv_x1_sg U46939 ( .A(n61201), .X(n61204) );
  nand_x1_sg U46940 ( .A(n61199), .B(n61198), .X(n42251) );
  inv_x1_sg U46941 ( .A(n61197), .X(n61198) );
  inv_x1_sg U46942 ( .A(n61196), .X(n61199) );
  nand_x1_sg U46943 ( .A(n61194), .B(n61193), .X(n42682) );
  inv_x1_sg U46944 ( .A(n61192), .X(n61193) );
  inv_x1_sg U46945 ( .A(n61191), .X(n61194) );
  nand_x1_sg U46946 ( .A(n61189), .B(n61188), .X(n42667) );
  inv_x1_sg U46947 ( .A(n61187), .X(n61188) );
  inv_x1_sg U46948 ( .A(n61186), .X(n61189) );
  nand_x1_sg U46949 ( .A(n61184), .B(n61183), .X(n42189) );
  inv_x1_sg U46950 ( .A(n61182), .X(n61183) );
  inv_x1_sg U46951 ( .A(n61181), .X(n61184) );
  nand_x1_sg U46952 ( .A(n61179), .B(n61178), .X(n42257) );
  inv_x1_sg U46953 ( .A(n61177), .X(n61178) );
  inv_x1_sg U46954 ( .A(n61176), .X(n61179) );
  nand_x1_sg U46955 ( .A(n61174), .B(n61173), .X(n42616) );
  inv_x1_sg U46956 ( .A(n61172), .X(n61173) );
  inv_x1_sg U46957 ( .A(n61171), .X(n61174) );
  nand_x1_sg U46958 ( .A(n61169), .B(n61168), .X(n42243) );
  inv_x1_sg U46959 ( .A(n61167), .X(n61168) );
  inv_x1_sg U46960 ( .A(n61166), .X(n61169) );
  nand_x1_sg U46961 ( .A(n61164), .B(n61163), .X(n42414) );
  inv_x1_sg U46962 ( .A(n61162), .X(n61163) );
  inv_x1_sg U46963 ( .A(n61161), .X(n61164) );
  nand_x1_sg U46964 ( .A(n61159), .B(n61158), .X(n42688) );
  inv_x1_sg U46965 ( .A(n61157), .X(n61158) );
  inv_x1_sg U46966 ( .A(n61156), .X(n61159) );
  nand_x1_sg U46967 ( .A(n61154), .B(n61153), .X(n42685) );
  inv_x1_sg U46968 ( .A(n61152), .X(n61153) );
  inv_x1_sg U46969 ( .A(n61151), .X(n61154) );
  nand_x1_sg U46970 ( .A(n61149), .B(n61148), .X(n42177) );
  inv_x1_sg U46971 ( .A(n61147), .X(n61148) );
  inv_x1_sg U46972 ( .A(n61146), .X(n61149) );
  nand_x1_sg U46973 ( .A(n61144), .B(n61143), .X(n42174) );
  inv_x1_sg U46974 ( .A(n61142), .X(n61143) );
  inv_x1_sg U46975 ( .A(n61141), .X(n61144) );
  nand_x1_sg U46976 ( .A(n61139), .B(n61138), .X(n42679) );
  inv_x1_sg U46977 ( .A(n61137), .X(n61138) );
  inv_x1_sg U46978 ( .A(n61136), .X(n61139) );
  nand_x1_sg U46979 ( .A(n61134), .B(n61133), .X(n42676) );
  inv_x1_sg U46980 ( .A(n61132), .X(n61133) );
  inv_x1_sg U46981 ( .A(n61131), .X(n61134) );
  nand_x1_sg U46982 ( .A(n61129), .B(n61128), .X(n42673) );
  inv_x1_sg U46983 ( .A(n61127), .X(n61128) );
  inv_x1_sg U46984 ( .A(n61126), .X(n61129) );
  nand_x1_sg U46985 ( .A(n61124), .B(n61123), .X(n42670) );
  inv_x1_sg U46986 ( .A(n61122), .X(n61123) );
  inv_x1_sg U46987 ( .A(n61121), .X(n61124) );
  nand_x1_sg U46988 ( .A(n61119), .B(n61118), .X(n42328) );
  inv_x1_sg U46989 ( .A(n61117), .X(n61118) );
  inv_x1_sg U46990 ( .A(n61116), .X(n61119) );
  nand_x1_sg U46991 ( .A(n61114), .B(n61113), .X(n42411) );
  inv_x1_sg U46992 ( .A(n61112), .X(n61113) );
  inv_x1_sg U46993 ( .A(n61111), .X(n61114) );
  nand_x1_sg U46994 ( .A(n61109), .B(n61108), .X(n42386) );
  inv_x1_sg U46995 ( .A(n61107), .X(n61108) );
  inv_x1_sg U46996 ( .A(n61106), .X(n61109) );
  nand_x1_sg U46997 ( .A(n61104), .B(n61103), .X(n42541) );
  inv_x1_sg U46998 ( .A(n61102), .X(n61103) );
  inv_x1_sg U46999 ( .A(n61101), .X(n61104) );
  nand_x1_sg U47000 ( .A(n61099), .B(n61098), .X(n42715) );
  inv_x1_sg U47001 ( .A(n61097), .X(n61098) );
  inv_x1_sg U47002 ( .A(n61096), .X(n61099) );
  nand_x1_sg U47003 ( .A(n61094), .B(n61093), .X(n42165) );
  inv_x1_sg U47004 ( .A(n61092), .X(n61093) );
  inv_x1_sg U47005 ( .A(n61091), .X(n61094) );
  nand_x1_sg U47006 ( .A(n61089), .B(n61088), .X(n42419) );
  inv_x1_sg U47007 ( .A(n61087), .X(n61088) );
  inv_x1_sg U47008 ( .A(n61086), .X(n61089) );
  nand_x1_sg U47009 ( .A(n61084), .B(n61083), .X(n42724) );
  inv_x1_sg U47010 ( .A(n61082), .X(n61083) );
  inv_x1_sg U47011 ( .A(n61081), .X(n61084) );
  nand_x1_sg U47012 ( .A(n61079), .B(n61078), .X(n42628) );
  inv_x1_sg U47013 ( .A(n61077), .X(n61078) );
  inv_x1_sg U47014 ( .A(n61076), .X(n61079) );
  nand_x1_sg U47015 ( .A(n61074), .B(n61073), .X(n42625) );
  inv_x1_sg U47016 ( .A(n61072), .X(n61073) );
  inv_x1_sg U47017 ( .A(n61071), .X(n61074) );
  nand_x1_sg U47018 ( .A(n61069), .B(n61068), .X(n42622) );
  inv_x1_sg U47019 ( .A(n61067), .X(n61068) );
  inv_x1_sg U47020 ( .A(n61066), .X(n61069) );
  nand_x1_sg U47021 ( .A(n61064), .B(n61063), .X(n42619) );
  inv_x1_sg U47022 ( .A(n61062), .X(n61063) );
  inv_x1_sg U47023 ( .A(n61061), .X(n61064) );
  nand_x1_sg U47024 ( .A(n61059), .B(n61058), .X(n42640) );
  inv_x1_sg U47025 ( .A(n61057), .X(n61058) );
  inv_x1_sg U47026 ( .A(n61056), .X(n61059) );
  nand_x1_sg U47027 ( .A(n61054), .B(n61053), .X(n42646) );
  inv_x1_sg U47028 ( .A(n61052), .X(n61053) );
  inv_x1_sg U47029 ( .A(n61051), .X(n61054) );
  nand_x1_sg U47030 ( .A(n61049), .B(n61048), .X(n42634) );
  inv_x1_sg U47031 ( .A(n61047), .X(n61048) );
  inv_x1_sg U47032 ( .A(n61046), .X(n61049) );
  nand_x1_sg U47033 ( .A(n61044), .B(n61043), .X(n42637) );
  inv_x1_sg U47034 ( .A(n61042), .X(n61043) );
  inv_x1_sg U47035 ( .A(n61041), .X(n61044) );
  nand_x1_sg U47036 ( .A(n61039), .B(n61038), .X(n42664) );
  inv_x1_sg U47037 ( .A(n61037), .X(n61038) );
  inv_x1_sg U47038 ( .A(n61036), .X(n61039) );
  nand_x1_sg U47039 ( .A(n61034), .B(n61033), .X(n42661) );
  inv_x1_sg U47040 ( .A(n61032), .X(n61033) );
  inv_x1_sg U47041 ( .A(n61031), .X(n61034) );
  nand_x1_sg U47042 ( .A(n61029), .B(n61028), .X(n42655) );
  inv_x1_sg U47043 ( .A(n61027), .X(n61028) );
  inv_x1_sg U47044 ( .A(n61026), .X(n61029) );
  nand_x1_sg U47045 ( .A(n61024), .B(n61023), .X(n42652) );
  inv_x1_sg U47046 ( .A(n61022), .X(n61023) );
  inv_x1_sg U47047 ( .A(n61021), .X(n61024) );
  nand_x1_sg U47048 ( .A(n61019), .B(n61018), .X(n42192) );
  inv_x1_sg U47049 ( .A(n61017), .X(n61018) );
  inv_x1_sg U47050 ( .A(n61016), .X(n61019) );
  nand_x1_sg U47051 ( .A(n61014), .B(n61013), .X(n42423) );
  inv_x1_sg U47052 ( .A(n61012), .X(n61013) );
  inv_x1_sg U47053 ( .A(n61011), .X(n61014) );
  nand_x1_sg U47054 ( .A(n61009), .B(n61008), .X(n42219) );
  inv_x1_sg U47055 ( .A(n61007), .X(n61008) );
  inv_x1_sg U47056 ( .A(n61006), .X(n61009) );
  nand_x1_sg U47057 ( .A(n61004), .B(n61003), .X(n42742) );
  inv_x1_sg U47058 ( .A(n61002), .X(n61003) );
  inv_x1_sg U47059 ( .A(n61001), .X(n61004) );
  nand_x1_sg U47060 ( .A(n60999), .B(n60998), .X(n42290) );
  inv_x1_sg U47061 ( .A(n60997), .X(n60998) );
  inv_x1_sg U47062 ( .A(n60996), .X(n60999) );
  nand_x1_sg U47063 ( .A(n60994), .B(n60993), .X(n42287) );
  inv_x1_sg U47064 ( .A(n60992), .X(n60993) );
  inv_x1_sg U47065 ( .A(n60991), .X(n60994) );
  nand_x1_sg U47066 ( .A(n60989), .B(n60988), .X(n42284) );
  inv_x1_sg U47067 ( .A(n60987), .X(n60988) );
  inv_x1_sg U47068 ( .A(n60986), .X(n60989) );
  nand_x1_sg U47069 ( .A(n60984), .B(n60983), .X(n42281) );
  inv_x1_sg U47070 ( .A(n60982), .X(n60983) );
  inv_x1_sg U47071 ( .A(n60981), .X(n60984) );
  nand_x1_sg U47072 ( .A(n60979), .B(n60978), .X(n42293) );
  inv_x1_sg U47073 ( .A(n60977), .X(n60978) );
  inv_x1_sg U47074 ( .A(n60976), .X(n60979) );
  nand_x1_sg U47075 ( .A(n60974), .B(n60973), .X(n42249) );
  inv_x1_sg U47076 ( .A(n60972), .X(n60973) );
  inv_x1_sg U47077 ( .A(n60971), .X(n60974) );
  nand_x1_sg U47078 ( .A(n60969), .B(n60968), .X(n42299) );
  inv_x1_sg U47079 ( .A(n60967), .X(n60968) );
  inv_x1_sg U47080 ( .A(n60966), .X(n60969) );
  nand_x1_sg U47081 ( .A(n60964), .B(n60963), .X(n42296) );
  inv_x1_sg U47082 ( .A(n60962), .X(n60963) );
  inv_x1_sg U47083 ( .A(n60961), .X(n60964) );
  nand_x1_sg U47084 ( .A(n60959), .B(n60958), .X(n42772) );
  inv_x1_sg U47085 ( .A(n60957), .X(n60958) );
  inv_x1_sg U47086 ( .A(n60956), .X(n60959) );
  nand_x1_sg U47087 ( .A(n60954), .B(n60953), .X(n42305) );
  inv_x1_sg U47088 ( .A(n60952), .X(n60953) );
  inv_x1_sg U47089 ( .A(n60951), .X(n60954) );
  nand_x1_sg U47090 ( .A(n60949), .B(n60948), .X(n42341) );
  inv_x1_sg U47091 ( .A(n60947), .X(n60948) );
  inv_x1_sg U47092 ( .A(n60946), .X(n60949) );
  nand_x1_sg U47093 ( .A(n60944), .B(n60943), .X(n42228) );
  inv_x1_sg U47094 ( .A(n60942), .X(n60943) );
  inv_x1_sg U47095 ( .A(n60941), .X(n60944) );
  nand_x1_sg U47096 ( .A(n60939), .B(n60938), .X(n42344) );
  inv_x1_sg U47097 ( .A(n60937), .X(n60938) );
  inv_x1_sg U47098 ( .A(n60936), .X(n60939) );
  nand_x1_sg U47099 ( .A(n60934), .B(n60933), .X(n42335) );
  inv_x1_sg U47100 ( .A(n60932), .X(n60933) );
  inv_x1_sg U47101 ( .A(n60931), .X(n60934) );
  nand_x1_sg U47102 ( .A(n60929), .B(n60928), .X(n42332) );
  inv_x1_sg U47103 ( .A(n60927), .X(n60928) );
  inv_x1_sg U47104 ( .A(n60926), .X(n60929) );
  nand_x1_sg U47105 ( .A(n60924), .B(n60923), .X(n42329) );
  inv_x1_sg U47106 ( .A(n60922), .X(n60923) );
  inv_x1_sg U47107 ( .A(n60921), .X(n60924) );
  nand_x1_sg U47108 ( .A(n60919), .B(n60918), .X(n42266) );
  inv_x1_sg U47109 ( .A(n60917), .X(n60918) );
  inv_x1_sg U47110 ( .A(n60916), .X(n60919) );
  nand_x1_sg U47111 ( .A(n60914), .B(n60913), .X(n42263) );
  inv_x1_sg U47112 ( .A(n60912), .X(n60913) );
  inv_x1_sg U47113 ( .A(n60911), .X(n60914) );
  nand_x1_sg U47114 ( .A(n60909), .B(n60908), .X(n42318) );
  inv_x1_sg U47115 ( .A(n60907), .X(n60908) );
  inv_x1_sg U47116 ( .A(n60906), .X(n60909) );
  nand_x1_sg U47117 ( .A(n60904), .B(n60903), .X(n42315) );
  inv_x1_sg U47118 ( .A(n60902), .X(n60903) );
  inv_x1_sg U47119 ( .A(n60901), .X(n60904) );
  nand_x1_sg U47120 ( .A(n60899), .B(n60898), .X(n42312) );
  inv_x1_sg U47121 ( .A(n60897), .X(n60898) );
  inv_x1_sg U47122 ( .A(n60896), .X(n60899) );
  nand_x1_sg U47123 ( .A(n60894), .B(n60893), .X(n42309) );
  inv_x1_sg U47124 ( .A(n60892), .X(n60893) );
  inv_x1_sg U47125 ( .A(n60891), .X(n60894) );
  nand_x1_sg U47126 ( .A(n60889), .B(n60888), .X(n42275) );
  inv_x1_sg U47127 ( .A(n60887), .X(n60888) );
  inv_x1_sg U47128 ( .A(n60886), .X(n60889) );
  nand_x1_sg U47129 ( .A(n60884), .B(n60883), .X(n42278) );
  inv_x1_sg U47130 ( .A(n60882), .X(n60883) );
  inv_x1_sg U47131 ( .A(n60881), .X(n60884) );
  nand_x1_sg U47132 ( .A(n60879), .B(n60878), .X(n42260) );
  inv_x1_sg U47133 ( .A(n60877), .X(n60878) );
  inv_x1_sg U47134 ( .A(n60876), .X(n60879) );
  nand_x1_sg U47135 ( .A(n60874), .B(n60873), .X(n42269) );
  inv_x1_sg U47136 ( .A(n60872), .X(n60873) );
  inv_x1_sg U47137 ( .A(n60871), .X(n60874) );
  nand_x1_sg U47138 ( .A(n60869), .B(n60868), .X(n42302) );
  inv_x1_sg U47139 ( .A(n60867), .X(n60868) );
  inv_x1_sg U47140 ( .A(n60866), .X(n60869) );
  nand_x1_sg U47141 ( .A(n60864), .B(n60863), .X(n42248) );
  inv_x1_sg U47142 ( .A(n60862), .X(n60863) );
  inv_x1_sg U47143 ( .A(n60861), .X(n60864) );
  nand_x1_sg U47144 ( .A(n60859), .B(n60858), .X(n42325) );
  inv_x1_sg U47145 ( .A(n60857), .X(n60858) );
  inv_x1_sg U47146 ( .A(n60856), .X(n60859) );
  nand_x1_sg U47147 ( .A(n60854), .B(n60853), .X(n42247) );
  inv_x1_sg U47148 ( .A(n60852), .X(n60853) );
  inv_x1_sg U47149 ( .A(n60851), .X(n60854) );
  nand_x1_sg U47150 ( .A(n60849), .B(n60848), .X(n42322) );
  inv_x1_sg U47151 ( .A(n60847), .X(n60848) );
  inv_x1_sg U47152 ( .A(n60846), .X(n60849) );
  nand_x1_sg U47153 ( .A(n60844), .B(n60843), .X(n42272) );
  inv_x1_sg U47154 ( .A(n60842), .X(n60843) );
  inv_x1_sg U47155 ( .A(n60841), .X(n60844) );
  nand_x1_sg U47156 ( .A(n60839), .B(n60838), .X(n42508) );
  inv_x1_sg U47157 ( .A(n60837), .X(n60838) );
  inv_x1_sg U47158 ( .A(n60836), .X(n60839) );
  nand_x1_sg U47159 ( .A(n60834), .B(n60833), .X(n42505) );
  inv_x1_sg U47160 ( .A(n60832), .X(n60833) );
  inv_x1_sg U47161 ( .A(n60831), .X(n60834) );
  nand_x1_sg U47162 ( .A(n60829), .B(n60828), .X(n42502) );
  inv_x1_sg U47163 ( .A(n60827), .X(n60828) );
  inv_x1_sg U47164 ( .A(n60826), .X(n60829) );
  nand_x1_sg U47165 ( .A(n60824), .B(n60823), .X(n42499) );
  inv_x1_sg U47166 ( .A(n60822), .X(n60823) );
  inv_x1_sg U47167 ( .A(n60821), .X(n60824) );
  nand_x1_sg U47168 ( .A(n60819), .B(n60818), .X(n42517) );
  inv_x1_sg U47169 ( .A(n60817), .X(n60818) );
  inv_x1_sg U47170 ( .A(n60816), .X(n60819) );
  nand_x1_sg U47171 ( .A(n60814), .B(n60813), .X(n42514) );
  inv_x1_sg U47172 ( .A(n60812), .X(n60813) );
  inv_x1_sg U47173 ( .A(n60811), .X(n60814) );
  nand_x1_sg U47174 ( .A(n60809), .B(n60808), .X(n42520) );
  inv_x1_sg U47175 ( .A(n60807), .X(n60808) );
  inv_x1_sg U47176 ( .A(n60806), .X(n60809) );
  nand_x1_sg U47177 ( .A(n60804), .B(n60803), .X(n42511) );
  inv_x1_sg U47178 ( .A(n60802), .X(n60803) );
  inv_x1_sg U47179 ( .A(n60801), .X(n60804) );
  nand_x1_sg U47180 ( .A(n60799), .B(n60798), .X(n42565) );
  inv_x1_sg U47181 ( .A(n60797), .X(n60798) );
  inv_x1_sg U47182 ( .A(n60796), .X(n60799) );
  nand_x1_sg U47183 ( .A(n60794), .B(n60793), .X(n42246) );
  inv_x1_sg U47184 ( .A(n60792), .X(n60793) );
  inv_x1_sg U47185 ( .A(n60791), .X(n60794) );
  nand_x1_sg U47186 ( .A(n60789), .B(n60788), .X(n42556) );
  inv_x1_sg U47187 ( .A(n60787), .X(n60788) );
  inv_x1_sg U47188 ( .A(n60786), .X(n60789) );
  nand_x1_sg U47189 ( .A(n60784), .B(n60783), .X(n42550) );
  inv_x1_sg U47190 ( .A(n60782), .X(n60783) );
  inv_x1_sg U47191 ( .A(n60781), .X(n60784) );
  nand_x1_sg U47192 ( .A(n60779), .B(n60778), .X(n42562) );
  inv_x1_sg U47193 ( .A(n60777), .X(n60778) );
  inv_x1_sg U47194 ( .A(n60776), .X(n60779) );
  nand_x1_sg U47195 ( .A(n60774), .B(n60773), .X(n42568) );
  inv_x1_sg U47196 ( .A(n60772), .X(n60773) );
  inv_x1_sg U47197 ( .A(n60771), .X(n60774) );
  nand_x1_sg U47198 ( .A(n60769), .B(n60768), .X(n42553) );
  inv_x1_sg U47199 ( .A(n60767), .X(n60768) );
  inv_x1_sg U47200 ( .A(n60766), .X(n60769) );
  nand_x1_sg U47201 ( .A(n60764), .B(n60763), .X(n42559) );
  inv_x1_sg U47202 ( .A(n60762), .X(n60763) );
  inv_x1_sg U47203 ( .A(n60761), .X(n60764) );
  nand_x1_sg U47204 ( .A(n60759), .B(n60758), .X(n42493) );
  inv_x1_sg U47205 ( .A(n60757), .X(n60758) );
  inv_x1_sg U47206 ( .A(n60756), .X(n60759) );
  nand_x1_sg U47207 ( .A(n60754), .B(n60753), .X(n42496) );
  inv_x1_sg U47208 ( .A(n60752), .X(n60753) );
  inv_x1_sg U47209 ( .A(n60751), .X(n60754) );
  nand_x1_sg U47210 ( .A(n60749), .B(n60748), .X(n42523) );
  inv_x1_sg U47211 ( .A(n60747), .X(n60748) );
  inv_x1_sg U47212 ( .A(n60746), .X(n60749) );
  nand_x1_sg U47213 ( .A(n60744), .B(n60743), .X(n42535) );
  inv_x1_sg U47214 ( .A(n60742), .X(n60743) );
  inv_x1_sg U47215 ( .A(n60741), .X(n60744) );
  nand_x1_sg U47216 ( .A(n60739), .B(n60738), .X(n42254) );
  inv_x1_sg U47217 ( .A(n60737), .X(n60738) );
  inv_x1_sg U47218 ( .A(n60736), .X(n60739) );
  nand_x1_sg U47219 ( .A(n60734), .B(n60733), .X(n42255) );
  inv_x1_sg U47220 ( .A(n60732), .X(n60733) );
  inv_x1_sg U47221 ( .A(n60731), .X(n60734) );
  nand_x1_sg U47222 ( .A(n60729), .B(n60728), .X(n42490) );
  inv_x1_sg U47223 ( .A(n60727), .X(n60728) );
  inv_x1_sg U47224 ( .A(n60726), .X(n60729) );
  nand_x1_sg U47225 ( .A(n60724), .B(n60723), .X(n42256) );
  inv_x1_sg U47226 ( .A(n60722), .X(n60723) );
  inv_x1_sg U47227 ( .A(n60721), .X(n60724) );
  nand_x1_sg U47228 ( .A(n60719), .B(n60718), .X(n42547) );
  inv_x1_sg U47229 ( .A(n60717), .X(n60718) );
  inv_x1_sg U47230 ( .A(n60716), .X(n60719) );
  nand_x1_sg U47231 ( .A(n60714), .B(n60713), .X(n42544) );
  inv_x1_sg U47232 ( .A(n60712), .X(n60713) );
  inv_x1_sg U47233 ( .A(n60711), .X(n60714) );
  nand_x1_sg U47234 ( .A(n60709), .B(n60708), .X(n42526) );
  inv_x1_sg U47235 ( .A(n60707), .X(n60708) );
  inv_x1_sg U47236 ( .A(n60706), .X(n60709) );
  nand_x1_sg U47237 ( .A(n60704), .B(n60703), .X(n42529) );
  inv_x1_sg U47238 ( .A(n60702), .X(n60703) );
  inv_x1_sg U47239 ( .A(n60701), .X(n60704) );
  nand_x1_sg U47240 ( .A(n60699), .B(n60698), .X(n42487) );
  inv_x1_sg U47241 ( .A(n60697), .X(n60698) );
  inv_x1_sg U47242 ( .A(n60696), .X(n60699) );
  nand_x1_sg U47243 ( .A(n60694), .B(n60693), .X(n42484) );
  inv_x1_sg U47244 ( .A(n60692), .X(n60693) );
  inv_x1_sg U47245 ( .A(n60691), .X(n60694) );
  nand_x1_sg U47246 ( .A(n60689), .B(n60688), .X(n42478) );
  inv_x1_sg U47247 ( .A(n60687), .X(n60688) );
  inv_x1_sg U47248 ( .A(n60686), .X(n60689) );
  nand_x1_sg U47249 ( .A(n60684), .B(n60683), .X(n42481) );
  inv_x1_sg U47250 ( .A(n60682), .X(n60683) );
  inv_x1_sg U47251 ( .A(n60681), .X(n60684) );
  nand_x1_sg U47252 ( .A(n60679), .B(n60678), .X(n42188) );
  inv_x1_sg U47253 ( .A(n60677), .X(n60678) );
  inv_x1_sg U47254 ( .A(n60676), .X(n60679) );
  nand_x1_sg U47255 ( .A(n60674), .B(n60673), .X(n42187) );
  inv_x1_sg U47256 ( .A(n60672), .X(n60673) );
  inv_x1_sg U47257 ( .A(n60671), .X(n60674) );
  nand_x1_sg U47258 ( .A(n60669), .B(n60668), .X(n42191) );
  inv_x1_sg U47259 ( .A(n60667), .X(n60668) );
  inv_x1_sg U47260 ( .A(n60666), .X(n60669) );
  nand_x1_sg U47261 ( .A(n60664), .B(n60663), .X(n42190) );
  inv_x1_sg U47262 ( .A(n60662), .X(n60663) );
  inv_x1_sg U47263 ( .A(n60661), .X(n60664) );
  nand_x1_sg U47264 ( .A(n60659), .B(n60658), .X(n42182) );
  inv_x1_sg U47265 ( .A(n60657), .X(n60658) );
  inv_x1_sg U47266 ( .A(n60656), .X(n60659) );
  nand_x1_sg U47267 ( .A(n60654), .B(n60653), .X(n42181) );
  inv_x1_sg U47268 ( .A(n60652), .X(n60653) );
  inv_x1_sg U47269 ( .A(n60651), .X(n60654) );
  nand_x1_sg U47270 ( .A(n60649), .B(n60648), .X(n42185) );
  inv_x1_sg U47271 ( .A(n60647), .X(n60648) );
  inv_x1_sg U47272 ( .A(n60646), .X(n60649) );
  nand_x1_sg U47273 ( .A(n60644), .B(n60643), .X(n42184) );
  inv_x1_sg U47274 ( .A(n60642), .X(n60643) );
  inv_x1_sg U47275 ( .A(n60641), .X(n60644) );
  nand_x1_sg U47276 ( .A(n60639), .B(n60638), .X(n42200) );
  inv_x1_sg U47277 ( .A(n60637), .X(n60638) );
  inv_x1_sg U47278 ( .A(n60636), .X(n60639) );
  nand_x1_sg U47279 ( .A(n60634), .B(n60633), .X(n42199) );
  inv_x1_sg U47280 ( .A(n60632), .X(n60633) );
  inv_x1_sg U47281 ( .A(n60631), .X(n60634) );
  nand_x1_sg U47282 ( .A(n60629), .B(n60628), .X(n42203) );
  inv_x1_sg U47283 ( .A(n60627), .X(n60628) );
  inv_x1_sg U47284 ( .A(n60626), .X(n60629) );
  nand_x1_sg U47285 ( .A(n60624), .B(n60623), .X(n42202) );
  inv_x1_sg U47286 ( .A(n60622), .X(n60623) );
  inv_x1_sg U47287 ( .A(n60621), .X(n60624) );
  nand_x1_sg U47288 ( .A(n60619), .B(n60618), .X(n42194) );
  inv_x1_sg U47289 ( .A(n60617), .X(n60618) );
  inv_x1_sg U47290 ( .A(n60616), .X(n60619) );
  nand_x1_sg U47291 ( .A(n60614), .B(n60613), .X(n42193) );
  inv_x1_sg U47292 ( .A(n60612), .X(n60613) );
  inv_x1_sg U47293 ( .A(n60611), .X(n60614) );
  nand_x1_sg U47294 ( .A(n60609), .B(n60608), .X(n42197) );
  inv_x1_sg U47295 ( .A(n60607), .X(n60608) );
  inv_x1_sg U47296 ( .A(n60606), .X(n60609) );
  nand_x1_sg U47297 ( .A(n60604), .B(n60603), .X(n42196) );
  inv_x1_sg U47298 ( .A(n60602), .X(n60603) );
  inv_x1_sg U47299 ( .A(n60601), .X(n60604) );
  nand_x1_sg U47300 ( .A(n60599), .B(n60598), .X(n42164) );
  inv_x1_sg U47301 ( .A(n60597), .X(n60598) );
  inv_x1_sg U47302 ( .A(n60596), .X(n60599) );
  nand_x1_sg U47303 ( .A(n60594), .B(n60593), .X(n42163) );
  inv_x1_sg U47304 ( .A(n60592), .X(n60593) );
  inv_x1_sg U47305 ( .A(n60591), .X(n60594) );
  nand_x1_sg U47306 ( .A(n60589), .B(n60588), .X(n42253) );
  inv_x1_sg U47307 ( .A(n60587), .X(n60588) );
  inv_x1_sg U47308 ( .A(n60586), .X(n60589) );
  nand_x1_sg U47309 ( .A(n60584), .B(n60583), .X(n42252) );
  inv_x1_sg U47310 ( .A(n60582), .X(n60583) );
  inv_x1_sg U47311 ( .A(n60581), .X(n60584) );
  nand_x1_sg U47312 ( .A(n60579), .B(n60578), .X(n42721) );
  inv_x1_sg U47313 ( .A(n60577), .X(n60578) );
  inv_x1_sg U47314 ( .A(n60576), .X(n60579) );
  nand_x1_sg U47315 ( .A(n60574), .B(n60573), .X(n42718) );
  inv_x1_sg U47316 ( .A(n60572), .X(n60573) );
  inv_x1_sg U47317 ( .A(n60571), .X(n60574) );
  nand_x1_sg U47318 ( .A(n60569), .B(n60568), .X(n42167) );
  inv_x1_sg U47319 ( .A(n60567), .X(n60568) );
  inv_x1_sg U47320 ( .A(n60566), .X(n60569) );
  nand_x1_sg U47321 ( .A(n60564), .B(n60563), .X(n42166) );
  inv_x1_sg U47322 ( .A(n60562), .X(n60563) );
  inv_x1_sg U47323 ( .A(n60561), .X(n60564) );
  nand_x1_sg U47324 ( .A(n60559), .B(n60558), .X(n42176) );
  inv_x1_sg U47325 ( .A(n60557), .X(n60558) );
  inv_x1_sg U47326 ( .A(n60556), .X(n60559) );
  nand_x1_sg U47327 ( .A(n60554), .B(n60553), .X(n42175) );
  inv_x1_sg U47328 ( .A(n60552), .X(n60553) );
  inv_x1_sg U47329 ( .A(n60551), .X(n60554) );
  nand_x1_sg U47330 ( .A(n60549), .B(n60548), .X(n42179) );
  inv_x1_sg U47331 ( .A(n60547), .X(n60548) );
  inv_x1_sg U47332 ( .A(n60546), .X(n60549) );
  nand_x1_sg U47333 ( .A(n60544), .B(n60543), .X(n42178) );
  inv_x1_sg U47334 ( .A(n60542), .X(n60543) );
  inv_x1_sg U47335 ( .A(n60541), .X(n60544) );
  nand_x1_sg U47336 ( .A(n60539), .B(n60538), .X(n42170) );
  inv_x1_sg U47337 ( .A(n60537), .X(n60538) );
  inv_x1_sg U47338 ( .A(n60536), .X(n60539) );
  nand_x1_sg U47339 ( .A(n60534), .B(n60533), .X(n42169) );
  inv_x1_sg U47340 ( .A(n60532), .X(n60533) );
  inv_x1_sg U47341 ( .A(n60531), .X(n60534) );
  nand_x1_sg U47342 ( .A(n60529), .B(n60528), .X(n42173) );
  inv_x1_sg U47343 ( .A(n60527), .X(n60528) );
  inv_x1_sg U47344 ( .A(n60526), .X(n60529) );
  nand_x1_sg U47345 ( .A(n60524), .B(n60523), .X(n42172) );
  inv_x1_sg U47346 ( .A(n60522), .X(n60523) );
  inv_x1_sg U47347 ( .A(n60521), .X(n60524) );
  nand_x1_sg U47348 ( .A(n60519), .B(n60518), .X(n42239) );
  inv_x1_sg U47349 ( .A(n60517), .X(n60518) );
  inv_x1_sg U47350 ( .A(n60516), .X(n60519) );
  nand_x1_sg U47351 ( .A(n60514), .B(n60513), .X(n42238) );
  inv_x1_sg U47352 ( .A(n60512), .X(n60513) );
  inv_x1_sg U47353 ( .A(n60511), .X(n60514) );
  nand_x1_sg U47354 ( .A(n60509), .B(n60508), .X(n42242) );
  inv_x1_sg U47355 ( .A(n60507), .X(n60508) );
  inv_x1_sg U47356 ( .A(n60506), .X(n60509) );
  nand_x1_sg U47357 ( .A(n60504), .B(n60503), .X(n42241) );
  inv_x1_sg U47358 ( .A(n60502), .X(n60503) );
  inv_x1_sg U47359 ( .A(n60501), .X(n60504) );
  nand_x1_sg U47360 ( .A(n60499), .B(n60498), .X(n42233) );
  inv_x1_sg U47361 ( .A(n60497), .X(n60498) );
  inv_x1_sg U47362 ( .A(n60496), .X(n60499) );
  nand_x1_sg U47363 ( .A(n60494), .B(n60493), .X(n42232) );
  inv_x1_sg U47364 ( .A(n60492), .X(n60493) );
  inv_x1_sg U47365 ( .A(n60491), .X(n60494) );
  nand_x1_sg U47366 ( .A(n60489), .B(n60488), .X(n42236) );
  inv_x1_sg U47367 ( .A(n60487), .X(n60488) );
  inv_x1_sg U47368 ( .A(n60486), .X(n60489) );
  nand_x1_sg U47369 ( .A(n60484), .B(n60483), .X(n42235) );
  inv_x1_sg U47370 ( .A(n60482), .X(n60483) );
  inv_x1_sg U47371 ( .A(n60481), .X(n60484) );
  nand_x1_sg U47372 ( .A(n60479), .B(n60478), .X(n42739) );
  inv_x1_sg U47373 ( .A(n60477), .X(n60478) );
  inv_x1_sg U47374 ( .A(n60476), .X(n60479) );
  nand_x1_sg U47375 ( .A(n60474), .B(n60473), .X(n42757) );
  inv_x1_sg U47376 ( .A(n60472), .X(n60473) );
  inv_x1_sg U47377 ( .A(n60471), .X(n60474) );
  nand_x1_sg U47378 ( .A(n60469), .B(n60468), .X(n42736) );
  inv_x1_sg U47379 ( .A(n60467), .X(n60468) );
  inv_x1_sg U47380 ( .A(n60466), .X(n60469) );
  nand_x1_sg U47381 ( .A(n60464), .B(n60463), .X(n42733) );
  inv_x1_sg U47382 ( .A(n60462), .X(n60463) );
  inv_x1_sg U47383 ( .A(n60461), .X(n60464) );
  nand_x1_sg U47384 ( .A(n60459), .B(n60458), .X(n42763) );
  inv_x1_sg U47385 ( .A(n60457), .X(n60458) );
  inv_x1_sg U47386 ( .A(n60456), .X(n60459) );
  nand_x1_sg U47387 ( .A(n60454), .B(n60453), .X(n42760) );
  inv_x1_sg U47388 ( .A(n60452), .X(n60453) );
  inv_x1_sg U47389 ( .A(n60451), .X(n60454) );
  nand_x1_sg U47390 ( .A(n60449), .B(n60448), .X(n42751) );
  inv_x1_sg U47391 ( .A(n60447), .X(n60448) );
  inv_x1_sg U47392 ( .A(n60446), .X(n60449) );
  nand_x1_sg U47393 ( .A(n60444), .B(n60443), .X(n42748) );
  inv_x1_sg U47394 ( .A(n60442), .X(n60443) );
  inv_x1_sg U47395 ( .A(n60441), .X(n60444) );
  nand_x1_sg U47396 ( .A(n60439), .B(n60438), .X(n42212) );
  inv_x1_sg U47397 ( .A(n60437), .X(n60438) );
  inv_x1_sg U47398 ( .A(n60436), .X(n60439) );
  nand_x1_sg U47399 ( .A(n60434), .B(n60433), .X(n42211) );
  inv_x1_sg U47400 ( .A(n60432), .X(n60433) );
  inv_x1_sg U47401 ( .A(n60431), .X(n60434) );
  nand_x1_sg U47402 ( .A(n60429), .B(n60428), .X(n42215) );
  inv_x1_sg U47403 ( .A(n60427), .X(n60428) );
  inv_x1_sg U47404 ( .A(n60426), .X(n60429) );
  nand_x1_sg U47405 ( .A(n60424), .B(n60423), .X(n42214) );
  inv_x1_sg U47406 ( .A(n60422), .X(n60423) );
  inv_x1_sg U47407 ( .A(n60421), .X(n60424) );
  nand_x1_sg U47408 ( .A(n60419), .B(n60418), .X(n42206) );
  inv_x1_sg U47409 ( .A(n60417), .X(n60418) );
  inv_x1_sg U47410 ( .A(n60416), .X(n60419) );
  nand_x1_sg U47411 ( .A(n60414), .B(n60413), .X(n42205) );
  inv_x1_sg U47412 ( .A(n60412), .X(n60413) );
  inv_x1_sg U47413 ( .A(n60411), .X(n60414) );
  nand_x1_sg U47414 ( .A(n60409), .B(n60408), .X(n42209) );
  inv_x1_sg U47415 ( .A(n60407), .X(n60408) );
  inv_x1_sg U47416 ( .A(n60406), .X(n60409) );
  nand_x1_sg U47417 ( .A(n60404), .B(n60403), .X(n42208) );
  inv_x1_sg U47418 ( .A(n60402), .X(n60403) );
  inv_x1_sg U47419 ( .A(n60401), .X(n60404) );
  nand_x1_sg U47420 ( .A(n60399), .B(n60398), .X(n42224) );
  inv_x1_sg U47421 ( .A(n60397), .X(n60398) );
  inv_x1_sg U47422 ( .A(n60396), .X(n60399) );
  nand_x1_sg U47423 ( .A(n60394), .B(n60393), .X(n42223) );
  inv_x1_sg U47424 ( .A(n60392), .X(n60393) );
  inv_x1_sg U47425 ( .A(n60391), .X(n60394) );
  nand_x1_sg U47426 ( .A(n60389), .B(n60388), .X(n42227) );
  inv_x1_sg U47427 ( .A(n60387), .X(n60388) );
  inv_x1_sg U47428 ( .A(n60386), .X(n60389) );
  nand_x1_sg U47429 ( .A(n60384), .B(n60383), .X(n42226) );
  inv_x1_sg U47430 ( .A(n60382), .X(n60383) );
  inv_x1_sg U47431 ( .A(n60381), .X(n60384) );
  nand_x1_sg U47432 ( .A(n60379), .B(n60378), .X(n42218) );
  inv_x1_sg U47433 ( .A(n60377), .X(n60378) );
  inv_x1_sg U47434 ( .A(n60376), .X(n60379) );
  nand_x1_sg U47435 ( .A(n60374), .B(n60373), .X(n42217) );
  inv_x1_sg U47436 ( .A(n60372), .X(n60373) );
  inv_x1_sg U47437 ( .A(n60371), .X(n60374) );
  nand_x1_sg U47438 ( .A(n60369), .B(n60368), .X(n42221) );
  inv_x1_sg U47439 ( .A(n60367), .X(n60368) );
  inv_x1_sg U47440 ( .A(n60366), .X(n60369) );
  nand_x1_sg U47441 ( .A(n60364), .B(n60363), .X(n42220) );
  inv_x1_sg U47442 ( .A(n60362), .X(n60363) );
  inv_x1_sg U47443 ( .A(n60361), .X(n60364) );
  nand_x1_sg U47444 ( .A(n60359), .B(n60358), .X(n42216) );
  inv_x1_sg U47445 ( .A(n60357), .X(n60358) );
  inv_x1_sg U47446 ( .A(n60356), .X(n60359) );
  nand_x1_sg U47447 ( .A(n60354), .B(n60353), .X(n42245) );
  inv_x1_sg U47448 ( .A(n60352), .X(n60353) );
  inv_x1_sg U47449 ( .A(n60351), .X(n60354) );
  nand_x1_sg U47450 ( .A(n60349), .B(n60348), .X(n42198) );
  inv_x1_sg U47451 ( .A(n60347), .X(n60348) );
  inv_x1_sg U47452 ( .A(n60346), .X(n60349) );
  nand_x1_sg U47453 ( .A(n60344), .B(n60343), .X(n42195) );
  inv_x1_sg U47454 ( .A(n60342), .X(n60343) );
  inv_x1_sg U47455 ( .A(n60341), .X(n60344) );
  nand_x1_sg U47456 ( .A(n60339), .B(n60338), .X(n42162) );
  inv_x1_sg U47457 ( .A(n60337), .X(n60338) );
  inv_x1_sg U47458 ( .A(n60336), .X(n60339) );
  nand_x1_sg U47459 ( .A(n60334), .B(n60333), .X(n42244) );
  inv_x1_sg U47460 ( .A(n60332), .X(n60333) );
  inv_x1_sg U47461 ( .A(n60331), .X(n60334) );
  nand_x1_sg U47462 ( .A(n60329), .B(n60328), .X(n42416) );
  inv_x1_sg U47463 ( .A(n60327), .X(n60328) );
  inv_x1_sg U47464 ( .A(n60326), .X(n60329) );
  nand_x1_sg U47465 ( .A(n60324), .B(n60323), .X(n42359) );
  inv_x1_sg U47466 ( .A(n60322), .X(n60323) );
  inv_x1_sg U47467 ( .A(n60321), .X(n60324) );
  nand_x1_sg U47468 ( .A(n60319), .B(n60318), .X(n42371) );
  inv_x1_sg U47469 ( .A(n60317), .X(n60318) );
  inv_x1_sg U47470 ( .A(n60316), .X(n60319) );
  nand_x1_sg U47471 ( .A(n60314), .B(n60313), .X(n42415) );
  inv_x1_sg U47472 ( .A(n60312), .X(n60313) );
  inv_x1_sg U47473 ( .A(n60311), .X(n60314) );
  nand_x1_sg U47474 ( .A(n60309), .B(n60308), .X(n42368) );
  inv_x1_sg U47475 ( .A(n60307), .X(n60308) );
  inv_x1_sg U47476 ( .A(n60306), .X(n60309) );
  nand_x1_sg U47477 ( .A(n60304), .B(n60303), .X(n42362) );
  inv_x1_sg U47478 ( .A(n60302), .X(n60303) );
  inv_x1_sg U47479 ( .A(n60301), .X(n60304) );
  nand_x1_sg U47480 ( .A(n60299), .B(n60298), .X(n42240) );
  inv_x1_sg U47481 ( .A(n60297), .X(n60298) );
  inv_x1_sg U47482 ( .A(n60296), .X(n60299) );
  nand_x1_sg U47483 ( .A(n60294), .B(n60293), .X(n42234) );
  inv_x1_sg U47484 ( .A(n60292), .X(n60293) );
  inv_x1_sg U47485 ( .A(n60291), .X(n60294) );
  nand_x1_sg U47486 ( .A(n60289), .B(n60288), .X(n42231) );
  inv_x1_sg U47487 ( .A(n60287), .X(n60288) );
  inv_x1_sg U47488 ( .A(n60286), .X(n60289) );
  nand_x1_sg U47489 ( .A(n60284), .B(n60283), .X(n42225) );
  inv_x1_sg U47490 ( .A(n60282), .X(n60283) );
  inv_x1_sg U47491 ( .A(n60281), .X(n60284) );
  nand_x1_sg U47492 ( .A(n60279), .B(n60278), .X(n42694) );
  inv_x1_sg U47493 ( .A(n60277), .X(n60278) );
  inv_x1_sg U47494 ( .A(n60276), .X(n60279) );
  nand_x1_sg U47495 ( .A(n60274), .B(n60273), .X(n42691) );
  inv_x1_sg U47496 ( .A(n60272), .X(n60273) );
  inv_x1_sg U47497 ( .A(n60271), .X(n60274) );
  nand_x1_sg U47498 ( .A(n60269), .B(n60268), .X(n42186) );
  inv_x1_sg U47499 ( .A(n60267), .X(n60268) );
  inv_x1_sg U47500 ( .A(n60266), .X(n60269) );
  nand_x1_sg U47501 ( .A(n60264), .B(n60263), .X(n42183) );
  inv_x1_sg U47502 ( .A(n60262), .X(n60263) );
  inv_x1_sg U47503 ( .A(n60261), .X(n60264) );
  nand_x1_sg U47504 ( .A(n60259), .B(n60258), .X(n42703) );
  inv_x1_sg U47505 ( .A(n60257), .X(n60258) );
  inv_x1_sg U47506 ( .A(n60256), .X(n60259) );
  nand_x1_sg U47507 ( .A(n60254), .B(n60253), .X(n42180) );
  inv_x1_sg U47508 ( .A(n60252), .X(n60253) );
  inv_x1_sg U47509 ( .A(n60251), .X(n60254) );
  nand_x1_sg U47510 ( .A(n60249), .B(n60248), .X(n42700) );
  inv_x1_sg U47511 ( .A(n60247), .X(n60248) );
  inv_x1_sg U47512 ( .A(n60246), .X(n60249) );
  nand_x1_sg U47513 ( .A(n60244), .B(n60243), .X(n42697) );
  inv_x1_sg U47514 ( .A(n60242), .X(n60243) );
  inv_x1_sg U47515 ( .A(n60241), .X(n60244) );
  nand_x1_sg U47516 ( .A(n60239), .B(n60238), .X(n42213) );
  inv_x1_sg U47517 ( .A(n60237), .X(n60238) );
  inv_x1_sg U47518 ( .A(n60236), .X(n60239) );
  nand_x1_sg U47519 ( .A(n60234), .B(n60233), .X(n42210) );
  inv_x1_sg U47520 ( .A(n60232), .X(n60233) );
  inv_x1_sg U47521 ( .A(n60231), .X(n60234) );
  nand_x1_sg U47522 ( .A(n60229), .B(n60228), .X(n42207) );
  inv_x1_sg U47523 ( .A(n60227), .X(n60228) );
  inv_x1_sg U47524 ( .A(n60226), .X(n60229) );
  nand_x1_sg U47525 ( .A(n60224), .B(n60223), .X(n42204) );
  inv_x1_sg U47526 ( .A(n60222), .X(n60223) );
  inv_x1_sg U47527 ( .A(n60221), .X(n60224) );
  nand_x1_sg U47528 ( .A(n60219), .B(n60218), .X(n42161) );
  inv_x1_sg U47529 ( .A(n60217), .X(n60218) );
  inv_x1_sg U47530 ( .A(n60216), .X(n60219) );
  nand_x1_sg U47531 ( .A(n60214), .B(n60213), .X(n42745) );
  inv_x1_sg U47532 ( .A(n60212), .X(n60213) );
  inv_x1_sg U47533 ( .A(n60211), .X(n60214) );
  nand_x1_sg U47534 ( .A(n60209), .B(n60208), .X(n42754) );
  inv_x1_sg U47535 ( .A(n60207), .X(n60208) );
  inv_x1_sg U47536 ( .A(n60206), .X(n60209) );
  nand_x1_sg U47537 ( .A(n60204), .B(n60203), .X(n42222) );
  inv_x1_sg U47538 ( .A(n60202), .X(n60203) );
  inv_x1_sg U47539 ( .A(n60201), .X(n60204) );
  nand_x1_sg U47540 ( .A(n60199), .B(n60198), .X(n42353) );
  inv_x1_sg U47541 ( .A(n60197), .X(n60198) );
  inv_x1_sg U47542 ( .A(n60196), .X(n60199) );
  nand_x1_sg U47543 ( .A(n60194), .B(n60193), .X(n42347) );
  inv_x1_sg U47544 ( .A(n60192), .X(n60193) );
  inv_x1_sg U47545 ( .A(n60191), .X(n60194) );
  nand_x1_sg U47546 ( .A(n60189), .B(n60188), .X(n42338) );
  inv_x1_sg U47547 ( .A(n60187), .X(n60188) );
  inv_x1_sg U47548 ( .A(n60186), .X(n60189) );
  nand_x1_sg U47549 ( .A(n60184), .B(n60183), .X(n42401) );
  inv_x1_sg U47550 ( .A(n60182), .X(n60183) );
  inv_x1_sg U47551 ( .A(n60181), .X(n60184) );
  nand_x1_sg U47552 ( .A(n60179), .B(n60178), .X(n42356) );
  inv_x1_sg U47553 ( .A(n60177), .X(n60178) );
  inv_x1_sg U47554 ( .A(n60176), .X(n60179) );
  nand_x1_sg U47555 ( .A(n60174), .B(n60173), .X(n42420) );
  inv_x1_sg U47556 ( .A(n60172), .X(n60173) );
  inv_x1_sg U47557 ( .A(n60171), .X(n60174) );
  nand_x1_sg U47558 ( .A(n60169), .B(n60168), .X(n42350) );
  inv_x1_sg U47559 ( .A(n60167), .X(n60168) );
  inv_x1_sg U47560 ( .A(n60166), .X(n60169) );
  nand_x1_sg U47561 ( .A(n60164), .B(n60163), .X(n42404) );
  inv_x1_sg U47562 ( .A(n60162), .X(n60163) );
  inv_x1_sg U47563 ( .A(n60161), .X(n60164) );
  nand_x1_sg U47564 ( .A(n60159), .B(n60158), .X(n42712) );
  inv_x1_sg U47565 ( .A(n60157), .X(n60158) );
  inv_x1_sg U47566 ( .A(n60156), .X(n60159) );
  nand_x1_sg U47567 ( .A(n60154), .B(n60153), .X(n42418) );
  inv_x1_sg U47568 ( .A(n60152), .X(n60153) );
  inv_x1_sg U47569 ( .A(n60151), .X(n60154) );
  nand_x1_sg U47570 ( .A(n60149), .B(n60148), .X(n42709) );
  inv_x1_sg U47571 ( .A(n60147), .X(n60148) );
  inv_x1_sg U47572 ( .A(n60146), .X(n60149) );
  nand_x1_sg U47573 ( .A(n60144), .B(n60143), .X(n42706) );
  inv_x1_sg U47574 ( .A(n60142), .X(n60143) );
  inv_x1_sg U47575 ( .A(n60141), .X(n60144) );
  nand_x1_sg U47576 ( .A(n60139), .B(n60138), .X(n42422) );
  inv_x1_sg U47577 ( .A(n60137), .X(n60138) );
  inv_x1_sg U47578 ( .A(n60136), .X(n60139) );
  nand_x1_sg U47579 ( .A(n60134), .B(n60133), .X(n42407) );
  inv_x1_sg U47580 ( .A(n60132), .X(n60133) );
  inv_x1_sg U47581 ( .A(n60131), .X(n60134) );
  nand_x1_sg U47582 ( .A(n60129), .B(n60128), .X(n42730) );
  inv_x1_sg U47583 ( .A(n60127), .X(n60128) );
  inv_x1_sg U47584 ( .A(n60126), .X(n60129) );
  nand_x1_sg U47585 ( .A(n60124), .B(n60123), .X(n42727) );
  inv_x1_sg U47586 ( .A(n60122), .X(n60123) );
  inv_x1_sg U47587 ( .A(n60121), .X(n60124) );
  nand_x1_sg U47588 ( .A(n60119), .B(n60118), .X(n42398) );
  inv_x1_sg U47589 ( .A(n60117), .X(n60118) );
  inv_x1_sg U47590 ( .A(n60116), .X(n60119) );
  nand_x1_sg U47591 ( .A(n60114), .B(n60113), .X(n42395) );
  inv_x1_sg U47592 ( .A(n60112), .X(n60113) );
  inv_x1_sg U47593 ( .A(n60111), .X(n60114) );
  nand_x1_sg U47594 ( .A(n60109), .B(n60108), .X(n42365) );
  inv_x1_sg U47595 ( .A(n60107), .X(n60108) );
  inv_x1_sg U47596 ( .A(n60106), .X(n60109) );
  nand_x1_sg U47597 ( .A(n60104), .B(n60103), .X(n42538) );
  inv_x1_sg U47598 ( .A(n60102), .X(n60103) );
  inv_x1_sg U47599 ( .A(n60101), .X(n60104) );
  nand_x1_sg U47600 ( .A(n60099), .B(n60098), .X(n42237) );
  inv_x1_sg U47601 ( .A(n60097), .X(n60098) );
  inv_x1_sg U47602 ( .A(n60096), .X(n60099) );
  nand_x1_sg U47603 ( .A(n60094), .B(n60093), .X(n42201) );
  inv_x1_sg U47604 ( .A(n60092), .X(n60093) );
  inv_x1_sg U47605 ( .A(n60091), .X(n60094) );
  nand_x1_sg U47606 ( .A(n60089), .B(n60088), .X(n42171) );
  inv_x1_sg U47607 ( .A(n60087), .X(n60088) );
  inv_x1_sg U47608 ( .A(n60086), .X(n60089) );
  nand_x1_sg U47609 ( .A(n60084), .B(n60083), .X(n42168) );
  inv_x1_sg U47610 ( .A(n60082), .X(n60083) );
  inv_x1_sg U47611 ( .A(n60081), .X(n60084) );
  nand_x1_sg U47612 ( .A(n60079), .B(n60078), .X(n42383) );
  inv_x1_sg U47613 ( .A(n60077), .X(n60078) );
  inv_x1_sg U47614 ( .A(n60076), .X(n60079) );
  nand_x1_sg U47615 ( .A(n60074), .B(n60073), .X(n42380) );
  inv_x1_sg U47616 ( .A(n60072), .X(n60073) );
  inv_x1_sg U47617 ( .A(n60071), .X(n60074) );
  nand_x1_sg U47618 ( .A(n60069), .B(n60068), .X(n42377) );
  inv_x1_sg U47619 ( .A(n60067), .X(n60068) );
  inv_x1_sg U47620 ( .A(n60066), .X(n60069) );
  nand_x1_sg U47621 ( .A(n60064), .B(n60063), .X(n42374) );
  inv_x1_sg U47622 ( .A(n60062), .X(n60063) );
  inv_x1_sg U47623 ( .A(n60061), .X(n60064) );
  nand_x1_sg U47624 ( .A(n60059), .B(n60058), .X(n42408) );
  inv_x1_sg U47625 ( .A(n60057), .X(n60058) );
  inv_x1_sg U47626 ( .A(n60056), .X(n60059) );
  nand_x1_sg U47627 ( .A(n60054), .B(n60053), .X(n42532) );
  inv_x1_sg U47628 ( .A(n60052), .X(n60053) );
  inv_x1_sg U47629 ( .A(n60051), .X(n60054) );
  nand_x1_sg U47630 ( .A(n60049), .B(n60048), .X(n42392) );
  inv_x1_sg U47631 ( .A(n60047), .X(n60048) );
  inv_x1_sg U47632 ( .A(n60046), .X(n60049) );
  nand_x1_sg U47633 ( .A(n60044), .B(n60043), .X(n42389) );
  inv_x1_sg U47634 ( .A(n60042), .X(n60043) );
  inv_x1_sg U47635 ( .A(n60041), .X(n60044) );
  nand_x1_sg U47636 ( .A(n60039), .B(n60038), .X(n42552) );
  inv_x1_sg U47637 ( .A(n60037), .X(n60038) );
  inv_x1_sg U47638 ( .A(n60036), .X(n60039) );
  nand_x1_sg U47639 ( .A(n60034), .B(n60033), .X(n42551) );
  inv_x1_sg U47640 ( .A(n60032), .X(n60033) );
  inv_x1_sg U47641 ( .A(n60031), .X(n60034) );
  nand_x1_sg U47642 ( .A(n60029), .B(n60028), .X(n42555) );
  inv_x1_sg U47643 ( .A(n60027), .X(n60028) );
  inv_x1_sg U47644 ( .A(n60026), .X(n60029) );
  nand_x1_sg U47645 ( .A(n60024), .B(n60023), .X(n42554) );
  inv_x1_sg U47646 ( .A(n60022), .X(n60023) );
  inv_x1_sg U47647 ( .A(n60021), .X(n60024) );
  nand_x1_sg U47648 ( .A(n60019), .B(n60018), .X(n42546) );
  inv_x1_sg U47649 ( .A(n60017), .X(n60018) );
  inv_x1_sg U47650 ( .A(n60016), .X(n60019) );
  nand_x1_sg U47651 ( .A(n60014), .B(n60013), .X(n42545) );
  inv_x1_sg U47652 ( .A(n60012), .X(n60013) );
  inv_x1_sg U47653 ( .A(n60011), .X(n60014) );
  nand_x1_sg U47654 ( .A(n60009), .B(n60008), .X(n42549) );
  inv_x1_sg U47655 ( .A(n60007), .X(n60008) );
  inv_x1_sg U47656 ( .A(n60006), .X(n60009) );
  nand_x1_sg U47657 ( .A(n60004), .B(n60003), .X(n42548) );
  inv_x1_sg U47658 ( .A(n60002), .X(n60003) );
  inv_x1_sg U47659 ( .A(n60001), .X(n60004) );
  nand_x1_sg U47660 ( .A(n59999), .B(n59998), .X(n42564) );
  inv_x1_sg U47661 ( .A(n59997), .X(n59998) );
  inv_x1_sg U47662 ( .A(n59996), .X(n59999) );
  nand_x1_sg U47663 ( .A(n59994), .B(n59993), .X(n42563) );
  inv_x1_sg U47664 ( .A(n59992), .X(n59993) );
  inv_x1_sg U47665 ( .A(n59991), .X(n59994) );
  nand_x1_sg U47666 ( .A(n59989), .B(n59988), .X(n42567) );
  inv_x1_sg U47667 ( .A(n59987), .X(n59988) );
  inv_x1_sg U47668 ( .A(n59986), .X(n59989) );
  nand_x1_sg U47669 ( .A(n59984), .B(n59983), .X(n42566) );
  inv_x1_sg U47670 ( .A(n59982), .X(n59983) );
  inv_x1_sg U47671 ( .A(n59981), .X(n59984) );
  nand_x1_sg U47672 ( .A(n59979), .B(n59978), .X(n42558) );
  inv_x1_sg U47673 ( .A(n59977), .X(n59978) );
  inv_x1_sg U47674 ( .A(n59976), .X(n59979) );
  nand_x1_sg U47675 ( .A(n59974), .B(n59973), .X(n42557) );
  inv_x1_sg U47676 ( .A(n59972), .X(n59973) );
  inv_x1_sg U47677 ( .A(n59971), .X(n59974) );
  nand_x1_sg U47678 ( .A(n59969), .B(n59968), .X(n42561) );
  inv_x1_sg U47679 ( .A(n59967), .X(n59968) );
  inv_x1_sg U47680 ( .A(n59966), .X(n59969) );
  nand_x1_sg U47681 ( .A(n59964), .B(n59963), .X(n42560) );
  inv_x1_sg U47682 ( .A(n59962), .X(n59963) );
  inv_x1_sg U47683 ( .A(n59961), .X(n59964) );
  nand_x1_sg U47684 ( .A(n59959), .B(n59958), .X(n42528) );
  inv_x1_sg U47685 ( .A(n59957), .X(n59958) );
  inv_x1_sg U47686 ( .A(n59956), .X(n59959) );
  nand_x1_sg U47687 ( .A(n59954), .B(n59953), .X(n42527) );
  inv_x1_sg U47688 ( .A(n59952), .X(n59953) );
  inv_x1_sg U47689 ( .A(n59951), .X(n59954) );
  nand_x1_sg U47690 ( .A(n59949), .B(n59948), .X(n42531) );
  inv_x1_sg U47691 ( .A(n59947), .X(n59948) );
  inv_x1_sg U47692 ( .A(n59946), .X(n59949) );
  nand_x1_sg U47693 ( .A(n59944), .B(n59943), .X(n42530) );
  inv_x1_sg U47694 ( .A(n59942), .X(n59943) );
  inv_x1_sg U47695 ( .A(n59941), .X(n59944) );
  nand_x1_sg U47696 ( .A(n59939), .B(n59938), .X(n42522) );
  inv_x1_sg U47697 ( .A(n59937), .X(n59938) );
  inv_x1_sg U47698 ( .A(n59936), .X(n59939) );
  nand_x1_sg U47699 ( .A(n59934), .B(n59933), .X(n42521) );
  inv_x1_sg U47700 ( .A(n59932), .X(n59933) );
  inv_x1_sg U47701 ( .A(n59931), .X(n59934) );
  nand_x1_sg U47702 ( .A(n59929), .B(n59928), .X(n42525) );
  inv_x1_sg U47703 ( .A(n59927), .X(n59928) );
  inv_x1_sg U47704 ( .A(n59926), .X(n59929) );
  nand_x1_sg U47705 ( .A(n59924), .B(n59923), .X(n42524) );
  inv_x1_sg U47706 ( .A(n59922), .X(n59923) );
  inv_x1_sg U47707 ( .A(n59921), .X(n59924) );
  nand_x1_sg U47708 ( .A(n59919), .B(n59918), .X(n42540) );
  inv_x1_sg U47709 ( .A(n59917), .X(n59918) );
  inv_x1_sg U47710 ( .A(n59916), .X(n59919) );
  nand_x1_sg U47711 ( .A(n59914), .B(n59913), .X(n42539) );
  inv_x1_sg U47712 ( .A(n59912), .X(n59913) );
  inv_x1_sg U47713 ( .A(n59911), .X(n59914) );
  nand_x1_sg U47714 ( .A(n59909), .B(n59908), .X(n42543) );
  inv_x1_sg U47715 ( .A(n59907), .X(n59908) );
  inv_x1_sg U47716 ( .A(n59906), .X(n59909) );
  nand_x1_sg U47717 ( .A(n59904), .B(n59903), .X(n42542) );
  inv_x1_sg U47718 ( .A(n59902), .X(n59903) );
  inv_x1_sg U47719 ( .A(n59901), .X(n59904) );
  nand_x1_sg U47720 ( .A(n59899), .B(n59898), .X(n42534) );
  inv_x1_sg U47721 ( .A(n59897), .X(n59898) );
  inv_x1_sg U47722 ( .A(n59896), .X(n59899) );
  nand_x1_sg U47723 ( .A(n59894), .B(n59893), .X(n42533) );
  inv_x1_sg U47724 ( .A(n59892), .X(n59893) );
  inv_x1_sg U47725 ( .A(n59891), .X(n59894) );
  nand_x1_sg U47726 ( .A(n59889), .B(n59888), .X(n42537) );
  inv_x1_sg U47727 ( .A(n59887), .X(n59888) );
  inv_x1_sg U47728 ( .A(n59886), .X(n59889) );
  nand_x1_sg U47729 ( .A(n59884), .B(n59883), .X(n42536) );
  inv_x1_sg U47730 ( .A(n59882), .X(n59883) );
  inv_x1_sg U47731 ( .A(n59881), .X(n59884) );
  nand_x1_sg U47732 ( .A(n59879), .B(n59878), .X(n42600) );
  inv_x1_sg U47733 ( .A(n59877), .X(n59878) );
  inv_x1_sg U47734 ( .A(n59876), .X(n59879) );
  nand_x1_sg U47735 ( .A(n59874), .B(n59873), .X(n42599) );
  inv_x1_sg U47736 ( .A(n59872), .X(n59873) );
  inv_x1_sg U47737 ( .A(n59871), .X(n59874) );
  nand_x1_sg U47738 ( .A(n59869), .B(n59868), .X(n42603) );
  inv_x1_sg U47739 ( .A(n59867), .X(n59868) );
  inv_x1_sg U47740 ( .A(n59866), .X(n59869) );
  nand_x1_sg U47741 ( .A(n59864), .B(n59863), .X(n42602) );
  inv_x1_sg U47742 ( .A(n59862), .X(n59863) );
  inv_x1_sg U47743 ( .A(n59861), .X(n59864) );
  nand_x1_sg U47744 ( .A(n59859), .B(n59858), .X(n42594) );
  inv_x1_sg U47745 ( .A(n59857), .X(n59858) );
  inv_x1_sg U47746 ( .A(n59856), .X(n59859) );
  nand_x1_sg U47747 ( .A(n59854), .B(n59853), .X(n42593) );
  inv_x1_sg U47748 ( .A(n59852), .X(n59853) );
  inv_x1_sg U47749 ( .A(n59851), .X(n59854) );
  nand_x1_sg U47750 ( .A(n59849), .B(n59848), .X(n42597) );
  inv_x1_sg U47751 ( .A(n59847), .X(n59848) );
  inv_x1_sg U47752 ( .A(n59846), .X(n59849) );
  nand_x1_sg U47753 ( .A(n59844), .B(n59843), .X(n42596) );
  inv_x1_sg U47754 ( .A(n59842), .X(n59843) );
  inv_x1_sg U47755 ( .A(n59841), .X(n59844) );
  nand_x1_sg U47756 ( .A(n59839), .B(n59838), .X(n42612) );
  inv_x1_sg U47757 ( .A(n59837), .X(n59838) );
  inv_x1_sg U47758 ( .A(n59836), .X(n59839) );
  nand_x1_sg U47759 ( .A(n59834), .B(n59833), .X(n42611) );
  inv_x1_sg U47760 ( .A(n59832), .X(n59833) );
  inv_x1_sg U47761 ( .A(n59831), .X(n59834) );
  nand_x1_sg U47762 ( .A(n59829), .B(n59828), .X(n42615) );
  inv_x1_sg U47763 ( .A(n59827), .X(n59828) );
  inv_x1_sg U47764 ( .A(n59826), .X(n59829) );
  nand_x1_sg U47765 ( .A(n59824), .B(n59823), .X(n42614) );
  inv_x1_sg U47766 ( .A(n59822), .X(n59823) );
  inv_x1_sg U47767 ( .A(n59821), .X(n59824) );
  nand_x1_sg U47768 ( .A(n59819), .B(n59818), .X(n42606) );
  inv_x1_sg U47769 ( .A(n59817), .X(n59818) );
  inv_x1_sg U47770 ( .A(n59816), .X(n59819) );
  nand_x1_sg U47771 ( .A(n59814), .B(n59813), .X(n42605) );
  inv_x1_sg U47772 ( .A(n59812), .X(n59813) );
  inv_x1_sg U47773 ( .A(n59811), .X(n59814) );
  nand_x1_sg U47774 ( .A(n59809), .B(n59808), .X(n42609) );
  inv_x1_sg U47775 ( .A(n59807), .X(n59808) );
  inv_x1_sg U47776 ( .A(n59806), .X(n59809) );
  nand_x1_sg U47777 ( .A(n59804), .B(n59803), .X(n42608) );
  inv_x1_sg U47778 ( .A(n59802), .X(n59803) );
  inv_x1_sg U47779 ( .A(n59801), .X(n59804) );
  nand_x1_sg U47780 ( .A(n59799), .B(n59798), .X(n42576) );
  inv_x1_sg U47781 ( .A(n59797), .X(n59798) );
  inv_x1_sg U47782 ( .A(n59796), .X(n59799) );
  nand_x1_sg U47783 ( .A(n59794), .B(n59793), .X(n42575) );
  inv_x1_sg U47784 ( .A(n59792), .X(n59793) );
  inv_x1_sg U47785 ( .A(n59791), .X(n59794) );
  nand_x1_sg U47786 ( .A(n59789), .B(n59788), .X(n42579) );
  inv_x1_sg U47787 ( .A(n59787), .X(n59788) );
  inv_x1_sg U47788 ( .A(n59786), .X(n59789) );
  nand_x1_sg U47789 ( .A(n59784), .B(n59783), .X(n42578) );
  inv_x1_sg U47790 ( .A(n59782), .X(n59783) );
  inv_x1_sg U47791 ( .A(n59781), .X(n59784) );
  nand_x1_sg U47792 ( .A(n59779), .B(n59778), .X(n42570) );
  inv_x1_sg U47793 ( .A(n59777), .X(n59778) );
  inv_x1_sg U47794 ( .A(n59776), .X(n59779) );
  nand_x1_sg U47795 ( .A(n59774), .B(n59773), .X(n42569) );
  inv_x1_sg U47796 ( .A(n59772), .X(n59773) );
  inv_x1_sg U47797 ( .A(n59771), .X(n59774) );
  nand_x1_sg U47798 ( .A(n59769), .B(n59768), .X(n42573) );
  inv_x1_sg U47799 ( .A(n59767), .X(n59768) );
  inv_x1_sg U47800 ( .A(n59766), .X(n59769) );
  nand_x1_sg U47801 ( .A(n59764), .B(n59763), .X(n42572) );
  inv_x1_sg U47802 ( .A(n59762), .X(n59763) );
  inv_x1_sg U47803 ( .A(n59761), .X(n59764) );
  nand_x1_sg U47804 ( .A(n59759), .B(n59758), .X(n42588) );
  inv_x1_sg U47805 ( .A(n59757), .X(n59758) );
  inv_x1_sg U47806 ( .A(n59756), .X(n59759) );
  nand_x1_sg U47807 ( .A(n59754), .B(n59753), .X(n42587) );
  inv_x1_sg U47808 ( .A(n59752), .X(n59753) );
  inv_x1_sg U47809 ( .A(n59751), .X(n59754) );
  nand_x1_sg U47810 ( .A(n59749), .B(n59748), .X(n42591) );
  inv_x1_sg U47811 ( .A(n59747), .X(n59748) );
  inv_x1_sg U47812 ( .A(n59746), .X(n59749) );
  nand_x1_sg U47813 ( .A(n59744), .B(n59743), .X(n42590) );
  inv_x1_sg U47814 ( .A(n59742), .X(n59743) );
  inv_x1_sg U47815 ( .A(n59741), .X(n59744) );
  nand_x1_sg U47816 ( .A(n59739), .B(n59738), .X(n42582) );
  inv_x1_sg U47817 ( .A(n59737), .X(n59738) );
  inv_x1_sg U47818 ( .A(n59736), .X(n59739) );
  nand_x1_sg U47819 ( .A(n59734), .B(n59733), .X(n42581) );
  inv_x1_sg U47820 ( .A(n59732), .X(n59733) );
  inv_x1_sg U47821 ( .A(n59731), .X(n59734) );
  nand_x1_sg U47822 ( .A(n59729), .B(n59728), .X(n42585) );
  inv_x1_sg U47823 ( .A(n59727), .X(n59728) );
  inv_x1_sg U47824 ( .A(n59726), .X(n59729) );
  nand_x1_sg U47825 ( .A(n59724), .B(n59723), .X(n42584) );
  inv_x1_sg U47826 ( .A(n59722), .X(n59723) );
  inv_x1_sg U47827 ( .A(n59721), .X(n59724) );
  nand_x1_sg U47828 ( .A(n59719), .B(n59718), .X(n42456) );
  inv_x1_sg U47829 ( .A(n59717), .X(n59718) );
  inv_x1_sg U47830 ( .A(n59716), .X(n59719) );
  nand_x1_sg U47831 ( .A(n59714), .B(n59713), .X(n42455) );
  inv_x1_sg U47832 ( .A(n59712), .X(n59713) );
  inv_x1_sg U47833 ( .A(n59711), .X(n59714) );
  nand_x1_sg U47834 ( .A(n59709), .B(n59708), .X(n42459) );
  inv_x1_sg U47835 ( .A(n59707), .X(n59708) );
  inv_x1_sg U47836 ( .A(n59706), .X(n59709) );
  nand_x1_sg U47837 ( .A(n59704), .B(n59703), .X(n42458) );
  inv_x1_sg U47838 ( .A(n59702), .X(n59703) );
  inv_x1_sg U47839 ( .A(n59701), .X(n59704) );
  nand_x1_sg U47840 ( .A(n59699), .B(n59698), .X(n42450) );
  inv_x1_sg U47841 ( .A(n59697), .X(n59698) );
  inv_x1_sg U47842 ( .A(n59696), .X(n59699) );
  nand_x1_sg U47843 ( .A(n59694), .B(n59693), .X(n42449) );
  inv_x1_sg U47844 ( .A(n59692), .X(n59693) );
  inv_x1_sg U47845 ( .A(n59691), .X(n59694) );
  nand_x1_sg U47846 ( .A(n59689), .B(n59688), .X(n42453) );
  inv_x1_sg U47847 ( .A(n59687), .X(n59688) );
  inv_x1_sg U47848 ( .A(n59686), .X(n59689) );
  nand_x1_sg U47849 ( .A(n59684), .B(n59683), .X(n42452) );
  inv_x1_sg U47850 ( .A(n59682), .X(n59683) );
  inv_x1_sg U47851 ( .A(n59681), .X(n59684) );
  nand_x1_sg U47852 ( .A(n59679), .B(n59678), .X(n42468) );
  inv_x1_sg U47853 ( .A(n59677), .X(n59678) );
  inv_x1_sg U47854 ( .A(n59676), .X(n59679) );
  nand_x1_sg U47855 ( .A(n59674), .B(n59673), .X(n42467) );
  inv_x1_sg U47856 ( .A(n59672), .X(n59673) );
  inv_x1_sg U47857 ( .A(n59671), .X(n59674) );
  nand_x1_sg U47858 ( .A(n59669), .B(n59668), .X(n42471) );
  inv_x1_sg U47859 ( .A(n59667), .X(n59668) );
  inv_x1_sg U47860 ( .A(n59666), .X(n59669) );
  nand_x1_sg U47861 ( .A(n59664), .B(n59663), .X(n42470) );
  inv_x1_sg U47862 ( .A(n59662), .X(n59663) );
  inv_x1_sg U47863 ( .A(n59661), .X(n59664) );
  nand_x1_sg U47864 ( .A(n59659), .B(n59658), .X(n42462) );
  inv_x1_sg U47865 ( .A(n59657), .X(n59658) );
  inv_x1_sg U47866 ( .A(n59656), .X(n59659) );
  nand_x1_sg U47867 ( .A(n59654), .B(n59653), .X(n42461) );
  inv_x1_sg U47868 ( .A(n59652), .X(n59653) );
  inv_x1_sg U47869 ( .A(n59651), .X(n59654) );
  nand_x1_sg U47870 ( .A(n59649), .B(n59648), .X(n42465) );
  inv_x1_sg U47871 ( .A(n59647), .X(n59648) );
  inv_x1_sg U47872 ( .A(n59646), .X(n59649) );
  nand_x1_sg U47873 ( .A(n59644), .B(n59643), .X(n42464) );
  inv_x1_sg U47874 ( .A(n59642), .X(n59643) );
  inv_x1_sg U47875 ( .A(n59641), .X(n59644) );
  nand_x1_sg U47876 ( .A(n59639), .B(n59638), .X(n42435) );
  inv_x1_sg U47877 ( .A(n59637), .X(n59638) );
  inv_x1_sg U47878 ( .A(n59636), .X(n59639) );
  nand_x1_sg U47879 ( .A(n59634), .B(n59633), .X(n42434) );
  inv_x1_sg U47880 ( .A(n59632), .X(n59633) );
  inv_x1_sg U47881 ( .A(n59631), .X(n59634) );
  nand_x1_sg U47882 ( .A(n59629), .B(n59628), .X(n42795) );
  inv_x1_sg U47883 ( .A(n59627), .X(n59628) );
  inv_x1_sg U47884 ( .A(n59626), .X(n59629) );
  nand_x1_sg U47885 ( .A(n59624), .B(n59623), .X(n42430) );
  inv_x1_sg U47886 ( .A(n59622), .X(n59623) );
  inv_x1_sg U47887 ( .A(n59621), .X(n59624) );
  nand_x1_sg U47888 ( .A(n59619), .B(n59618), .X(n42426) );
  inv_x1_sg U47889 ( .A(n59617), .X(n59618) );
  inv_x1_sg U47890 ( .A(n59616), .X(n59619) );
  nand_x1_sg U47891 ( .A(n59614), .B(n59613), .X(n42425) );
  inv_x1_sg U47892 ( .A(n59612), .X(n59613) );
  inv_x1_sg U47893 ( .A(n59611), .X(n59614) );
  nand_x1_sg U47894 ( .A(n59609), .B(n59608), .X(n42429) );
  inv_x1_sg U47895 ( .A(n59607), .X(n59608) );
  inv_x1_sg U47896 ( .A(n59606), .X(n59609) );
  nand_x1_sg U47897 ( .A(n59604), .B(n59603), .X(n42428) );
  inv_x1_sg U47898 ( .A(n59602), .X(n59603) );
  inv_x1_sg U47899 ( .A(n59601), .X(n59604) );
  nand_x1_sg U47900 ( .A(n59599), .B(n59598), .X(n42444) );
  inv_x1_sg U47901 ( .A(n59597), .X(n59598) );
  inv_x1_sg U47902 ( .A(n59596), .X(n59599) );
  nand_x1_sg U47903 ( .A(n59594), .B(n59593), .X(n42443) );
  inv_x1_sg U47904 ( .A(n59592), .X(n59593) );
  inv_x1_sg U47905 ( .A(n59591), .X(n59594) );
  nand_x1_sg U47906 ( .A(n59589), .B(n59588), .X(n42447) );
  inv_x1_sg U47907 ( .A(n59587), .X(n59588) );
  inv_x1_sg U47908 ( .A(n59586), .X(n59589) );
  nand_x1_sg U47909 ( .A(n59584), .B(n59583), .X(n42446) );
  inv_x1_sg U47910 ( .A(n59582), .X(n59583) );
  inv_x1_sg U47911 ( .A(n59581), .X(n59584) );
  nand_x1_sg U47912 ( .A(n59579), .B(n59578), .X(n42438) );
  inv_x1_sg U47913 ( .A(n59577), .X(n59578) );
  inv_x1_sg U47914 ( .A(n59576), .X(n59579) );
  nand_x1_sg U47915 ( .A(n59574), .B(n59573), .X(n42437) );
  inv_x1_sg U47916 ( .A(n59572), .X(n59573) );
  inv_x1_sg U47917 ( .A(n59571), .X(n59574) );
  nand_x1_sg U47918 ( .A(n59569), .B(n59568), .X(n42441) );
  inv_x1_sg U47919 ( .A(n59567), .X(n59568) );
  inv_x1_sg U47920 ( .A(n59566), .X(n59569) );
  nand_x1_sg U47921 ( .A(n59564), .B(n59563), .X(n42440) );
  inv_x1_sg U47922 ( .A(n59562), .X(n59563) );
  inv_x1_sg U47923 ( .A(n59561), .X(n59564) );
  nand_x1_sg U47924 ( .A(n59559), .B(n59558), .X(n42504) );
  inv_x1_sg U47925 ( .A(n59557), .X(n59558) );
  inv_x1_sg U47926 ( .A(n59556), .X(n59559) );
  nand_x1_sg U47927 ( .A(n59554), .B(n59553), .X(n42503) );
  inv_x1_sg U47928 ( .A(n59552), .X(n59553) );
  inv_x1_sg U47929 ( .A(n59551), .X(n59554) );
  nand_x1_sg U47930 ( .A(n59549), .B(n59548), .X(n42507) );
  inv_x1_sg U47931 ( .A(n59547), .X(n59548) );
  inv_x1_sg U47932 ( .A(n59546), .X(n59549) );
  nand_x1_sg U47933 ( .A(n59544), .B(n59543), .X(n42506) );
  inv_x1_sg U47934 ( .A(n59542), .X(n59543) );
  inv_x1_sg U47935 ( .A(n59541), .X(n59544) );
  nand_x1_sg U47936 ( .A(n59539), .B(n59538), .X(n42498) );
  inv_x1_sg U47937 ( .A(n59537), .X(n59538) );
  inv_x1_sg U47938 ( .A(n59536), .X(n59539) );
  nand_x1_sg U47939 ( .A(n59534), .B(n59533), .X(n42497) );
  inv_x1_sg U47940 ( .A(n59532), .X(n59533) );
  inv_x1_sg U47941 ( .A(n59531), .X(n59534) );
  nand_x1_sg U47942 ( .A(n59529), .B(n59528), .X(n42501) );
  inv_x1_sg U47943 ( .A(n59527), .X(n59528) );
  inv_x1_sg U47944 ( .A(n59526), .X(n59529) );
  nand_x1_sg U47945 ( .A(n59524), .B(n59523), .X(n42500) );
  inv_x1_sg U47946 ( .A(n59522), .X(n59523) );
  inv_x1_sg U47947 ( .A(n59521), .X(n59524) );
  nand_x1_sg U47948 ( .A(n59519), .B(n59518), .X(n42516) );
  inv_x1_sg U47949 ( .A(n59517), .X(n59518) );
  inv_x1_sg U47950 ( .A(n59516), .X(n59519) );
  nand_x1_sg U47951 ( .A(n59514), .B(n59513), .X(n42515) );
  inv_x1_sg U47952 ( .A(n59512), .X(n59513) );
  inv_x1_sg U47953 ( .A(n59511), .X(n59514) );
  nand_x1_sg U47954 ( .A(n59509), .B(n59508), .X(n42519) );
  inv_x1_sg U47955 ( .A(n59507), .X(n59508) );
  inv_x1_sg U47956 ( .A(n59506), .X(n59509) );
  nand_x1_sg U47957 ( .A(n59504), .B(n59503), .X(n42518) );
  inv_x1_sg U47958 ( .A(n59502), .X(n59503) );
  inv_x1_sg U47959 ( .A(n59501), .X(n59504) );
  nand_x1_sg U47960 ( .A(n59499), .B(n59498), .X(n42510) );
  inv_x1_sg U47961 ( .A(n59497), .X(n59498) );
  inv_x1_sg U47962 ( .A(n59496), .X(n59499) );
  nand_x1_sg U47963 ( .A(n59494), .B(n59493), .X(n42509) );
  inv_x1_sg U47964 ( .A(n59492), .X(n59493) );
  inv_x1_sg U47965 ( .A(n59491), .X(n59494) );
  nand_x1_sg U47966 ( .A(n59489), .B(n59488), .X(n42513) );
  inv_x1_sg U47967 ( .A(n59487), .X(n59488) );
  inv_x1_sg U47968 ( .A(n59486), .X(n59489) );
  nand_x1_sg U47969 ( .A(n59484), .B(n59483), .X(n42512) );
  inv_x1_sg U47970 ( .A(n59482), .X(n59483) );
  inv_x1_sg U47971 ( .A(n59481), .X(n59484) );
  nand_x1_sg U47972 ( .A(n59479), .B(n59478), .X(n42480) );
  inv_x1_sg U47973 ( .A(n59477), .X(n59478) );
  inv_x1_sg U47974 ( .A(n59476), .X(n59479) );
  nand_x1_sg U47975 ( .A(n59474), .B(n59473), .X(n42479) );
  inv_x1_sg U47976 ( .A(n59472), .X(n59473) );
  inv_x1_sg U47977 ( .A(n59471), .X(n59474) );
  nand_x1_sg U47978 ( .A(n59469), .B(n59468), .X(n42483) );
  inv_x1_sg U47979 ( .A(n59467), .X(n59468) );
  inv_x1_sg U47980 ( .A(n59466), .X(n59469) );
  nand_x1_sg U47981 ( .A(n59464), .B(n59463), .X(n42482) );
  inv_x1_sg U47982 ( .A(n59462), .X(n59463) );
  inv_x1_sg U47983 ( .A(n59461), .X(n59464) );
  nand_x1_sg U47984 ( .A(n59459), .B(n59458), .X(n42474) );
  inv_x1_sg U47985 ( .A(n59457), .X(n59458) );
  inv_x1_sg U47986 ( .A(n59456), .X(n59459) );
  nand_x1_sg U47987 ( .A(n59454), .B(n59453), .X(n42473) );
  inv_x1_sg U47988 ( .A(n59452), .X(n59453) );
  inv_x1_sg U47989 ( .A(n59451), .X(n59454) );
  nand_x1_sg U47990 ( .A(n59449), .B(n59448), .X(n42477) );
  inv_x1_sg U47991 ( .A(n59447), .X(n59448) );
  inv_x1_sg U47992 ( .A(n59446), .X(n59449) );
  nand_x1_sg U47993 ( .A(n59444), .B(n59443), .X(n42476) );
  inv_x1_sg U47994 ( .A(n59442), .X(n59443) );
  inv_x1_sg U47995 ( .A(n59441), .X(n59444) );
  nand_x1_sg U47996 ( .A(n59439), .B(n59438), .X(n42492) );
  inv_x1_sg U47997 ( .A(n59437), .X(n59438) );
  inv_x1_sg U47998 ( .A(n59436), .X(n59439) );
  nand_x1_sg U47999 ( .A(n59434), .B(n59433), .X(n42491) );
  inv_x1_sg U48000 ( .A(n59432), .X(n59433) );
  inv_x1_sg U48001 ( .A(n59431), .X(n59434) );
  nand_x1_sg U48002 ( .A(n59429), .B(n59428), .X(n42495) );
  inv_x1_sg U48003 ( .A(n59427), .X(n59428) );
  inv_x1_sg U48004 ( .A(n59426), .X(n59429) );
  nand_x1_sg U48005 ( .A(n59424), .B(n59423), .X(n42494) );
  inv_x1_sg U48006 ( .A(n59422), .X(n59423) );
  inv_x1_sg U48007 ( .A(n59421), .X(n59424) );
  nand_x1_sg U48008 ( .A(n59419), .B(n59418), .X(n42486) );
  inv_x1_sg U48009 ( .A(n59417), .X(n59418) );
  inv_x1_sg U48010 ( .A(n59416), .X(n59419) );
  nand_x1_sg U48011 ( .A(n59414), .B(n59413), .X(n42485) );
  inv_x1_sg U48012 ( .A(n59412), .X(n59413) );
  inv_x1_sg U48013 ( .A(n59411), .X(n59414) );
  nand_x1_sg U48014 ( .A(n59409), .B(n59408), .X(n42489) );
  inv_x1_sg U48015 ( .A(n59407), .X(n59408) );
  inv_x1_sg U48016 ( .A(n59406), .X(n59409) );
  nand_x1_sg U48017 ( .A(n59404), .B(n59403), .X(n42488) );
  inv_x1_sg U48018 ( .A(n59402), .X(n59403) );
  inv_x1_sg U48019 ( .A(n59401), .X(n59404) );
  nand_x1_sg U48020 ( .A(n59399), .B(n59398), .X(n42744) );
  inv_x1_sg U48021 ( .A(n59397), .X(n59398) );
  inv_x1_sg U48022 ( .A(n59396), .X(n59399) );
  nand_x1_sg U48023 ( .A(n59394), .B(n59393), .X(n42743) );
  inv_x1_sg U48024 ( .A(n59392), .X(n59393) );
  inv_x1_sg U48025 ( .A(n59391), .X(n59394) );
  nand_x1_sg U48026 ( .A(n59389), .B(n59388), .X(n42747) );
  inv_x1_sg U48027 ( .A(n59387), .X(n59388) );
  inv_x1_sg U48028 ( .A(n59386), .X(n59389) );
  nand_x1_sg U48029 ( .A(n59384), .B(n59383), .X(n42746) );
  inv_x1_sg U48030 ( .A(n59382), .X(n59383) );
  inv_x1_sg U48031 ( .A(n59381), .X(n59384) );
  nand_x1_sg U48032 ( .A(n59379), .B(n59378), .X(n42738) );
  inv_x1_sg U48033 ( .A(n59377), .X(n59378) );
  inv_x1_sg U48034 ( .A(n59376), .X(n59379) );
  nand_x1_sg U48035 ( .A(n59374), .B(n59373), .X(n42737) );
  inv_x1_sg U48036 ( .A(n59372), .X(n59373) );
  inv_x1_sg U48037 ( .A(n59371), .X(n59374) );
  nand_x1_sg U48038 ( .A(n59369), .B(n59368), .X(n42741) );
  inv_x1_sg U48039 ( .A(n59367), .X(n59368) );
  inv_x1_sg U48040 ( .A(n59366), .X(n59369) );
  nand_x1_sg U48041 ( .A(n59364), .B(n59363), .X(n42740) );
  inv_x1_sg U48042 ( .A(n59362), .X(n59363) );
  inv_x1_sg U48043 ( .A(n59361), .X(n59364) );
  nand_x1_sg U48044 ( .A(n59359), .B(n59358), .X(n42756) );
  inv_x1_sg U48045 ( .A(n59357), .X(n59358) );
  inv_x1_sg U48046 ( .A(n59356), .X(n59359) );
  nand_x1_sg U48047 ( .A(n59354), .B(n59353), .X(n42755) );
  inv_x1_sg U48048 ( .A(n59352), .X(n59353) );
  inv_x1_sg U48049 ( .A(n59351), .X(n59354) );
  nand_x1_sg U48050 ( .A(n59349), .B(n59348), .X(n42759) );
  inv_x1_sg U48051 ( .A(n59347), .X(n59348) );
  inv_x1_sg U48052 ( .A(n59346), .X(n59349) );
  nand_x1_sg U48053 ( .A(n59344), .B(n59343), .X(n42758) );
  inv_x1_sg U48054 ( .A(n59342), .X(n59343) );
  inv_x1_sg U48055 ( .A(n59341), .X(n59344) );
  nand_x1_sg U48056 ( .A(n59339), .B(n59338), .X(n42750) );
  inv_x1_sg U48057 ( .A(n59337), .X(n59338) );
  inv_x1_sg U48058 ( .A(n59336), .X(n59339) );
  nand_x1_sg U48059 ( .A(n59334), .B(n59333), .X(n42749) );
  inv_x1_sg U48060 ( .A(n59332), .X(n59333) );
  inv_x1_sg U48061 ( .A(n59331), .X(n59334) );
  nand_x1_sg U48062 ( .A(n59329), .B(n59328), .X(n42753) );
  inv_x1_sg U48063 ( .A(n59327), .X(n59328) );
  inv_x1_sg U48064 ( .A(n59326), .X(n59329) );
  nand_x1_sg U48065 ( .A(n59324), .B(n59323), .X(n42752) );
  inv_x1_sg U48066 ( .A(n59322), .X(n59323) );
  inv_x1_sg U48067 ( .A(n59321), .X(n59324) );
  nand_x1_sg U48068 ( .A(n59319), .B(n59318), .X(n42720) );
  inv_x1_sg U48069 ( .A(n59317), .X(n59318) );
  inv_x1_sg U48070 ( .A(n59316), .X(n59319) );
  nand_x1_sg U48071 ( .A(n59314), .B(n59313), .X(n42719) );
  inv_x1_sg U48072 ( .A(n59312), .X(n59313) );
  inv_x1_sg U48073 ( .A(n59311), .X(n59314) );
  nand_x1_sg U48074 ( .A(n59309), .B(n59308), .X(n42723) );
  inv_x1_sg U48075 ( .A(n59307), .X(n59308) );
  inv_x1_sg U48076 ( .A(n59306), .X(n59309) );
  nand_x1_sg U48077 ( .A(n59304), .B(n59303), .X(n42722) );
  inv_x1_sg U48078 ( .A(n59302), .X(n59303) );
  inv_x1_sg U48079 ( .A(n59301), .X(n59304) );
  nand_x1_sg U48080 ( .A(n59299), .B(n59298), .X(n42714) );
  inv_x1_sg U48081 ( .A(n59297), .X(n59298) );
  inv_x1_sg U48082 ( .A(n59296), .X(n59299) );
  nand_x1_sg U48083 ( .A(n59294), .B(n59293), .X(n42713) );
  inv_x1_sg U48084 ( .A(n59292), .X(n59293) );
  inv_x1_sg U48085 ( .A(n59291), .X(n59294) );
  nand_x1_sg U48086 ( .A(n59289), .B(n59288), .X(n42717) );
  inv_x1_sg U48087 ( .A(n59287), .X(n59288) );
  inv_x1_sg U48088 ( .A(n59286), .X(n59289) );
  nand_x1_sg U48089 ( .A(n59284), .B(n59283), .X(n42716) );
  inv_x1_sg U48090 ( .A(n59282), .X(n59283) );
  inv_x1_sg U48091 ( .A(n59281), .X(n59284) );
  nand_x1_sg U48092 ( .A(n59279), .B(n59278), .X(n42732) );
  inv_x1_sg U48093 ( .A(n59277), .X(n59278) );
  inv_x1_sg U48094 ( .A(n59276), .X(n59279) );
  nand_x1_sg U48095 ( .A(n59274), .B(n59273), .X(n42731) );
  inv_x1_sg U48096 ( .A(n59272), .X(n59273) );
  inv_x1_sg U48097 ( .A(n59271), .X(n59274) );
  nand_x1_sg U48098 ( .A(n59269), .B(n59268), .X(n42735) );
  inv_x1_sg U48099 ( .A(n59267), .X(n59268) );
  inv_x1_sg U48100 ( .A(n59266), .X(n59269) );
  nand_x1_sg U48101 ( .A(n59264), .B(n59263), .X(n42734) );
  inv_x1_sg U48102 ( .A(n59262), .X(n59263) );
  inv_x1_sg U48103 ( .A(n59261), .X(n59264) );
  nand_x1_sg U48104 ( .A(n59259), .B(n59258), .X(n42726) );
  inv_x1_sg U48105 ( .A(n59257), .X(n59258) );
  inv_x1_sg U48106 ( .A(n59256), .X(n59259) );
  nand_x1_sg U48107 ( .A(n59254), .B(n59253), .X(n42725) );
  inv_x1_sg U48108 ( .A(n59252), .X(n59253) );
  inv_x1_sg U48109 ( .A(n59251), .X(n59254) );
  nand_x1_sg U48110 ( .A(n59249), .B(n59248), .X(n42729) );
  inv_x1_sg U48111 ( .A(n59247), .X(n59248) );
  inv_x1_sg U48112 ( .A(n59246), .X(n59249) );
  nand_x1_sg U48113 ( .A(n59244), .B(n59243), .X(n42728) );
  inv_x1_sg U48114 ( .A(n59242), .X(n59243) );
  inv_x1_sg U48115 ( .A(n59241), .X(n59244) );
  nand_x1_sg U48116 ( .A(n59239), .B(n59238), .X(n42432) );
  inv_x1_sg U48117 ( .A(n59237), .X(n59238) );
  inv_x1_sg U48118 ( .A(n59236), .X(n59239) );
  nand_x1_sg U48119 ( .A(n59234), .B(n59233), .X(n42431) );
  inv_x1_sg U48120 ( .A(n59232), .X(n59233) );
  inv_x1_sg U48121 ( .A(n59231), .X(n59234) );
  nand_x1_sg U48122 ( .A(n59229), .B(n59228), .X(n42797) );
  inv_x1_sg U48123 ( .A(n59227), .X(n59228) );
  inv_x1_sg U48124 ( .A(n59226), .X(n59229) );
  nand_x1_sg U48125 ( .A(n59224), .B(n59223), .X(n42796) );
  inv_x1_sg U48126 ( .A(n59222), .X(n59223) );
  inv_x1_sg U48127 ( .A(n59221), .X(n59224) );
  nand_x1_sg U48128 ( .A(n59219), .B(n59218), .X(n42786) );
  inv_x1_sg U48129 ( .A(n59217), .X(n59218) );
  inv_x1_sg U48130 ( .A(n59216), .X(n59219) );
  nand_x1_sg U48131 ( .A(n59214), .B(n59213), .X(n42785) );
  inv_x1_sg U48132 ( .A(n59212), .X(n59213) );
  inv_x1_sg U48133 ( .A(n59211), .X(n59214) );
  nand_x1_sg U48134 ( .A(n59209), .B(n59208), .X(n42789) );
  inv_x1_sg U48135 ( .A(n59207), .X(n59208) );
  inv_x1_sg U48136 ( .A(n59206), .X(n59209) );
  nand_x1_sg U48137 ( .A(n59204), .B(n59203), .X(n42788) );
  inv_x1_sg U48138 ( .A(n59202), .X(n59203) );
  inv_x1_sg U48139 ( .A(n59201), .X(n59204) );
  nand_x1_sg U48140 ( .A(n59199), .B(n59198), .X(n42790) );
  inv_x1_sg U48141 ( .A(n59197), .X(n59198) );
  inv_x1_sg U48142 ( .A(n59196), .X(n59199) );
  nand_x1_sg U48143 ( .A(n59194), .B(n59193), .X(n42798) );
  inv_x1_sg U48144 ( .A(n59192), .X(n59193) );
  inv_x1_sg U48145 ( .A(n59191), .X(n59194) );
  nand_x1_sg U48146 ( .A(n59189), .B(n59188), .X(n42800) );
  inv_x1_sg U48147 ( .A(n59187), .X(n59188) );
  inv_x1_sg U48148 ( .A(n59186), .X(n59189) );
  nand_x1_sg U48149 ( .A(n59184), .B(n59183), .X(n42799) );
  inv_x1_sg U48150 ( .A(n59182), .X(n59183) );
  inv_x1_sg U48151 ( .A(n59181), .X(n59184) );
  nand_x1_sg U48152 ( .A(n59179), .B(n59178), .X(n42792) );
  inv_x1_sg U48153 ( .A(n59177), .X(n59178) );
  inv_x1_sg U48154 ( .A(n59176), .X(n59179) );
  nand_x1_sg U48155 ( .A(n59174), .B(n59173), .X(n42791) );
  inv_x1_sg U48156 ( .A(n59172), .X(n59173) );
  inv_x1_sg U48157 ( .A(n59171), .X(n59174) );
  nand_x1_sg U48158 ( .A(n59169), .B(n59168), .X(n42794) );
  inv_x1_sg U48159 ( .A(n59167), .X(n59168) );
  inv_x1_sg U48160 ( .A(n59166), .X(n59169) );
  nand_x1_sg U48161 ( .A(n59164), .B(n59163), .X(n42793) );
  inv_x1_sg U48162 ( .A(n59162), .X(n59163) );
  inv_x1_sg U48163 ( .A(n59161), .X(n59164) );
  nand_x1_sg U48164 ( .A(n59159), .B(n59158), .X(n42768) );
  inv_x1_sg U48165 ( .A(n59157), .X(n59158) );
  inv_x1_sg U48166 ( .A(n59156), .X(n59159) );
  nand_x1_sg U48167 ( .A(n59154), .B(n59153), .X(n42767) );
  inv_x1_sg U48168 ( .A(n59152), .X(n59153) );
  inv_x1_sg U48169 ( .A(n59151), .X(n59154) );
  nand_x1_sg U48170 ( .A(n59149), .B(n59148), .X(n42771) );
  inv_x1_sg U48171 ( .A(n59147), .X(n59148) );
  inv_x1_sg U48172 ( .A(n59146), .X(n59149) );
  nand_x1_sg U48173 ( .A(n59144), .B(n59143), .X(n42770) );
  inv_x1_sg U48174 ( .A(n59142), .X(n59143) );
  inv_x1_sg U48175 ( .A(n59141), .X(n59144) );
  nand_x1_sg U48176 ( .A(n59139), .B(n59138), .X(n42762) );
  inv_x1_sg U48177 ( .A(n59137), .X(n59138) );
  inv_x1_sg U48178 ( .A(n59136), .X(n59139) );
  nand_x1_sg U48179 ( .A(n59134), .B(n59133), .X(n42761) );
  inv_x1_sg U48180 ( .A(n59132), .X(n59133) );
  inv_x1_sg U48181 ( .A(n59131), .X(n59134) );
  nand_x1_sg U48182 ( .A(n59129), .B(n59128), .X(n42765) );
  inv_x1_sg U48183 ( .A(n59127), .X(n59128) );
  inv_x1_sg U48184 ( .A(n59126), .X(n59129) );
  nand_x1_sg U48185 ( .A(n59124), .B(n59123), .X(n42764) );
  inv_x1_sg U48186 ( .A(n59122), .X(n59123) );
  inv_x1_sg U48187 ( .A(n59121), .X(n59124) );
  nand_x1_sg U48188 ( .A(n59119), .B(n59118), .X(n42780) );
  inv_x1_sg U48189 ( .A(n59117), .X(n59118) );
  inv_x1_sg U48190 ( .A(n59116), .X(n59119) );
  nand_x1_sg U48191 ( .A(n59114), .B(n59113), .X(n42779) );
  inv_x1_sg U48192 ( .A(n59112), .X(n59113) );
  inv_x1_sg U48193 ( .A(n59111), .X(n59114) );
  nand_x1_sg U48194 ( .A(n59109), .B(n59108), .X(n42783) );
  inv_x1_sg U48195 ( .A(n59107), .X(n59108) );
  inv_x1_sg U48196 ( .A(n59106), .X(n59109) );
  nand_x1_sg U48197 ( .A(n59104), .B(n59103), .X(n42782) );
  inv_x1_sg U48198 ( .A(n59102), .X(n59103) );
  inv_x1_sg U48199 ( .A(n59101), .X(n59104) );
  nand_x1_sg U48200 ( .A(n59099), .B(n59098), .X(n42774) );
  inv_x1_sg U48201 ( .A(n59097), .X(n59098) );
  inv_x1_sg U48202 ( .A(n59096), .X(n59099) );
  nand_x1_sg U48203 ( .A(n59094), .B(n59093), .X(n42773) );
  inv_x1_sg U48204 ( .A(n59092), .X(n59093) );
  inv_x1_sg U48205 ( .A(n59091), .X(n59094) );
  nand_x1_sg U48206 ( .A(n59089), .B(n59088), .X(n42777) );
  inv_x1_sg U48207 ( .A(n59087), .X(n59088) );
  inv_x1_sg U48208 ( .A(n59086), .X(n59089) );
  nand_x1_sg U48209 ( .A(n59084), .B(n59083), .X(n42776) );
  inv_x1_sg U48210 ( .A(n59082), .X(n59083) );
  inv_x1_sg U48211 ( .A(n59081), .X(n59084) );
  nand_x1_sg U48212 ( .A(n59079), .B(n59078), .X(n42648) );
  inv_x1_sg U48213 ( .A(n59077), .X(n59078) );
  inv_x1_sg U48214 ( .A(n59076), .X(n59079) );
  nand_x1_sg U48215 ( .A(n59074), .B(n59073), .X(n42647) );
  inv_x1_sg U48216 ( .A(n59072), .X(n59073) );
  inv_x1_sg U48217 ( .A(n59071), .X(n59074) );
  nand_x1_sg U48218 ( .A(n59069), .B(n59068), .X(n42651) );
  inv_x1_sg U48219 ( .A(n59067), .X(n59068) );
  inv_x1_sg U48220 ( .A(n59066), .X(n59069) );
  nand_x1_sg U48221 ( .A(n59064), .B(n59063), .X(n42650) );
  inv_x1_sg U48222 ( .A(n59062), .X(n59063) );
  inv_x1_sg U48223 ( .A(n59061), .X(n59064) );
  nand_x1_sg U48224 ( .A(n59059), .B(n59058), .X(n42642) );
  inv_x1_sg U48225 ( .A(n59057), .X(n59058) );
  inv_x1_sg U48226 ( .A(n59056), .X(n59059) );
  nand_x1_sg U48227 ( .A(n59054), .B(n59053), .X(n42641) );
  inv_x1_sg U48228 ( .A(n59052), .X(n59053) );
  inv_x1_sg U48229 ( .A(n59051), .X(n59054) );
  nand_x1_sg U48230 ( .A(n59049), .B(n59048), .X(n42645) );
  inv_x1_sg U48231 ( .A(n59047), .X(n59048) );
  inv_x1_sg U48232 ( .A(n59046), .X(n59049) );
  nand_x1_sg U48233 ( .A(n59044), .B(n59043), .X(n42644) );
  inv_x1_sg U48234 ( .A(n59042), .X(n59043) );
  inv_x1_sg U48235 ( .A(n59041), .X(n59044) );
  nand_x1_sg U48236 ( .A(n59039), .B(n59038), .X(n42660) );
  inv_x1_sg U48237 ( .A(n59037), .X(n59038) );
  inv_x1_sg U48238 ( .A(n59036), .X(n59039) );
  nand_x1_sg U48239 ( .A(n59034), .B(n59033), .X(n42659) );
  inv_x1_sg U48240 ( .A(n59032), .X(n59033) );
  inv_x1_sg U48241 ( .A(n59031), .X(n59034) );
  nand_x1_sg U48242 ( .A(n59029), .B(n59028), .X(n42663) );
  inv_x1_sg U48243 ( .A(n59027), .X(n59028) );
  inv_x1_sg U48244 ( .A(n59026), .X(n59029) );
  nand_x1_sg U48245 ( .A(n59024), .B(n59023), .X(n42662) );
  inv_x1_sg U48246 ( .A(n59022), .X(n59023) );
  inv_x1_sg U48247 ( .A(n59021), .X(n59024) );
  nand_x1_sg U48248 ( .A(n59019), .B(n59018), .X(n42654) );
  inv_x1_sg U48249 ( .A(n59017), .X(n59018) );
  inv_x1_sg U48250 ( .A(n59016), .X(n59019) );
  nand_x1_sg U48251 ( .A(n59014), .B(n59013), .X(n42653) );
  inv_x1_sg U48252 ( .A(n59012), .X(n59013) );
  inv_x1_sg U48253 ( .A(n59011), .X(n59014) );
  nand_x1_sg U48254 ( .A(n59009), .B(n59008), .X(n42657) );
  inv_x1_sg U48255 ( .A(n59007), .X(n59008) );
  inv_x1_sg U48256 ( .A(n59006), .X(n59009) );
  nand_x1_sg U48257 ( .A(n59004), .B(n59003), .X(n42656) );
  inv_x1_sg U48258 ( .A(n59002), .X(n59003) );
  inv_x1_sg U48259 ( .A(n59001), .X(n59004) );
  nand_x1_sg U48260 ( .A(n58999), .B(n58998), .X(n42624) );
  inv_x1_sg U48261 ( .A(n58997), .X(n58998) );
  inv_x1_sg U48262 ( .A(n58996), .X(n58999) );
  nand_x1_sg U48263 ( .A(n58994), .B(n58993), .X(n42623) );
  inv_x1_sg U48264 ( .A(n58992), .X(n58993) );
  inv_x1_sg U48265 ( .A(n58991), .X(n58994) );
  nand_x1_sg U48266 ( .A(n58989), .B(n58988), .X(n42627) );
  inv_x1_sg U48267 ( .A(n58987), .X(n58988) );
  inv_x1_sg U48268 ( .A(n58986), .X(n58989) );
  nand_x1_sg U48269 ( .A(n58984), .B(n58983), .X(n42626) );
  inv_x1_sg U48270 ( .A(n58982), .X(n58983) );
  inv_x1_sg U48271 ( .A(n58981), .X(n58984) );
  nand_x1_sg U48272 ( .A(n58979), .B(n58978), .X(n42618) );
  inv_x1_sg U48273 ( .A(n58977), .X(n58978) );
  inv_x1_sg U48274 ( .A(n58976), .X(n58979) );
  nand_x1_sg U48275 ( .A(n58974), .B(n58973), .X(n42617) );
  inv_x1_sg U48276 ( .A(n58972), .X(n58973) );
  inv_x1_sg U48277 ( .A(n58971), .X(n58974) );
  nand_x1_sg U48278 ( .A(n58969), .B(n58968), .X(n42621) );
  inv_x1_sg U48279 ( .A(n58967), .X(n58968) );
  inv_x1_sg U48280 ( .A(n58966), .X(n58969) );
  nand_x1_sg U48281 ( .A(n58964), .B(n58963), .X(n42620) );
  inv_x1_sg U48282 ( .A(n58962), .X(n58963) );
  inv_x1_sg U48283 ( .A(n58961), .X(n58964) );
  nand_x1_sg U48284 ( .A(n58959), .B(n58958), .X(n42636) );
  inv_x1_sg U48285 ( .A(n58957), .X(n58958) );
  inv_x1_sg U48286 ( .A(n58956), .X(n58959) );
  nand_x1_sg U48287 ( .A(n58954), .B(n58953), .X(n42635) );
  inv_x1_sg U48288 ( .A(n58952), .X(n58953) );
  inv_x1_sg U48289 ( .A(n58951), .X(n58954) );
  nand_x1_sg U48290 ( .A(n58949), .B(n58948), .X(n42639) );
  inv_x1_sg U48291 ( .A(n58947), .X(n58948) );
  inv_x1_sg U48292 ( .A(n58946), .X(n58949) );
  nand_x1_sg U48293 ( .A(n58944), .B(n58943), .X(n42638) );
  inv_x1_sg U48294 ( .A(n58942), .X(n58943) );
  inv_x1_sg U48295 ( .A(n58941), .X(n58944) );
  nand_x1_sg U48296 ( .A(n58939), .B(n58938), .X(n42630) );
  inv_x1_sg U48297 ( .A(n58937), .X(n58938) );
  inv_x1_sg U48298 ( .A(n58936), .X(n58939) );
  nand_x1_sg U48299 ( .A(n58934), .B(n58933), .X(n42629) );
  inv_x1_sg U48300 ( .A(n58932), .X(n58933) );
  inv_x1_sg U48301 ( .A(n58931), .X(n58934) );
  nand_x1_sg U48302 ( .A(n58929), .B(n58928), .X(n42633) );
  inv_x1_sg U48303 ( .A(n58927), .X(n58928) );
  inv_x1_sg U48304 ( .A(n58926), .X(n58929) );
  nand_x1_sg U48305 ( .A(n58924), .B(n58923), .X(n42632) );
  inv_x1_sg U48306 ( .A(n58922), .X(n58923) );
  inv_x1_sg U48307 ( .A(n58921), .X(n58924) );
  nand_x1_sg U48308 ( .A(n58919), .B(n58918), .X(n42696) );
  inv_x1_sg U48309 ( .A(n58917), .X(n58918) );
  inv_x1_sg U48310 ( .A(n58916), .X(n58919) );
  nand_x1_sg U48311 ( .A(n58914), .B(n58913), .X(n42695) );
  inv_x1_sg U48312 ( .A(n58912), .X(n58913) );
  inv_x1_sg U48313 ( .A(n58911), .X(n58914) );
  nand_x1_sg U48314 ( .A(n58909), .B(n58908), .X(n42699) );
  inv_x1_sg U48315 ( .A(n58907), .X(n58908) );
  inv_x1_sg U48316 ( .A(n58906), .X(n58909) );
  nand_x1_sg U48317 ( .A(n58904), .B(n58903), .X(n42698) );
  inv_x1_sg U48318 ( .A(n58902), .X(n58903) );
  inv_x1_sg U48319 ( .A(n58901), .X(n58904) );
  nand_x1_sg U48320 ( .A(n58899), .B(n58898), .X(n42690) );
  inv_x1_sg U48321 ( .A(n58897), .X(n58898) );
  inv_x1_sg U48322 ( .A(n58896), .X(n58899) );
  nand_x1_sg U48323 ( .A(n58894), .B(n58893), .X(n42689) );
  inv_x1_sg U48324 ( .A(n58892), .X(n58893) );
  inv_x1_sg U48325 ( .A(n58891), .X(n58894) );
  nand_x1_sg U48326 ( .A(n58889), .B(n58888), .X(n42693) );
  inv_x1_sg U48327 ( .A(n58887), .X(n58888) );
  inv_x1_sg U48328 ( .A(n58886), .X(n58889) );
  nand_x1_sg U48329 ( .A(n58884), .B(n58883), .X(n42692) );
  inv_x1_sg U48330 ( .A(n58882), .X(n58883) );
  inv_x1_sg U48331 ( .A(n58881), .X(n58884) );
  nand_x1_sg U48332 ( .A(n58879), .B(n58878), .X(n42708) );
  inv_x1_sg U48333 ( .A(n58877), .X(n58878) );
  inv_x1_sg U48334 ( .A(n58876), .X(n58879) );
  nand_x1_sg U48335 ( .A(n58874), .B(n58873), .X(n42707) );
  inv_x1_sg U48336 ( .A(n58872), .X(n58873) );
  inv_x1_sg U48337 ( .A(n58871), .X(n58874) );
  nand_x1_sg U48338 ( .A(n58869), .B(n58868), .X(n42711) );
  inv_x1_sg U48339 ( .A(n58867), .X(n58868) );
  inv_x1_sg U48340 ( .A(n58866), .X(n58869) );
  nand_x1_sg U48341 ( .A(n58864), .B(n58863), .X(n42710) );
  inv_x1_sg U48342 ( .A(n58862), .X(n58863) );
  inv_x1_sg U48343 ( .A(n58861), .X(n58864) );
  nand_x1_sg U48344 ( .A(n58859), .B(n58858), .X(n42702) );
  inv_x1_sg U48345 ( .A(n58857), .X(n58858) );
  inv_x1_sg U48346 ( .A(n58856), .X(n58859) );
  nand_x1_sg U48347 ( .A(n58854), .B(n58853), .X(n42701) );
  inv_x1_sg U48348 ( .A(n58852), .X(n58853) );
  inv_x1_sg U48349 ( .A(n58851), .X(n58854) );
  nand_x1_sg U48350 ( .A(n58849), .B(n58848), .X(n42705) );
  inv_x1_sg U48351 ( .A(n58847), .X(n58848) );
  inv_x1_sg U48352 ( .A(n58846), .X(n58849) );
  nand_x1_sg U48353 ( .A(n58844), .B(n58843), .X(n42704) );
  inv_x1_sg U48354 ( .A(n58842), .X(n58843) );
  inv_x1_sg U48355 ( .A(n58841), .X(n58844) );
  nand_x1_sg U48356 ( .A(n58839), .B(n58838), .X(n42672) );
  inv_x1_sg U48357 ( .A(n58837), .X(n58838) );
  inv_x1_sg U48358 ( .A(n58836), .X(n58839) );
  nand_x1_sg U48359 ( .A(n58834), .B(n58833), .X(n42671) );
  inv_x1_sg U48360 ( .A(n58832), .X(n58833) );
  inv_x1_sg U48361 ( .A(n58831), .X(n58834) );
  nand_x1_sg U48362 ( .A(n58829), .B(n58828), .X(n42675) );
  inv_x1_sg U48363 ( .A(n58827), .X(n58828) );
  inv_x1_sg U48364 ( .A(n58826), .X(n58829) );
  nand_x1_sg U48365 ( .A(n58824), .B(n58823), .X(n42674) );
  inv_x1_sg U48366 ( .A(n58822), .X(n58823) );
  inv_x1_sg U48367 ( .A(n58821), .X(n58824) );
  nand_x1_sg U48368 ( .A(n58819), .B(n58818), .X(n42666) );
  inv_x1_sg U48369 ( .A(n58817), .X(n58818) );
  inv_x1_sg U48370 ( .A(n58816), .X(n58819) );
  nand_x1_sg U48371 ( .A(n58814), .B(n58813), .X(n42665) );
  inv_x1_sg U48372 ( .A(n58812), .X(n58813) );
  inv_x1_sg U48373 ( .A(n58811), .X(n58814) );
  nand_x1_sg U48374 ( .A(n58809), .B(n58808), .X(n42669) );
  inv_x1_sg U48375 ( .A(n58807), .X(n58808) );
  inv_x1_sg U48376 ( .A(n58806), .X(n58809) );
  nand_x1_sg U48377 ( .A(n58804), .B(n58803), .X(n42668) );
  inv_x1_sg U48378 ( .A(n58802), .X(n58803) );
  inv_x1_sg U48379 ( .A(n58801), .X(n58804) );
  nand_x1_sg U48380 ( .A(n58799), .B(n58798), .X(n42684) );
  inv_x1_sg U48381 ( .A(n58797), .X(n58798) );
  inv_x1_sg U48382 ( .A(n58796), .X(n58799) );
  nand_x1_sg U48383 ( .A(n58794), .B(n58793), .X(n42683) );
  inv_x1_sg U48384 ( .A(n58792), .X(n58793) );
  inv_x1_sg U48385 ( .A(n58791), .X(n58794) );
  nand_x1_sg U48386 ( .A(n58789), .B(n58788), .X(n42687) );
  inv_x1_sg U48387 ( .A(n58787), .X(n58788) );
  inv_x1_sg U48388 ( .A(n58786), .X(n58789) );
  nand_x1_sg U48389 ( .A(n58784), .B(n58783), .X(n42686) );
  inv_x1_sg U48390 ( .A(n58782), .X(n58783) );
  inv_x1_sg U48391 ( .A(n58781), .X(n58784) );
  nand_x1_sg U48392 ( .A(n58779), .B(n58778), .X(n42678) );
  inv_x1_sg U48393 ( .A(n58777), .X(n58778) );
  inv_x1_sg U48394 ( .A(n58776), .X(n58779) );
  nand_x1_sg U48395 ( .A(n58774), .B(n58773), .X(n42677) );
  inv_x1_sg U48396 ( .A(n58772), .X(n58773) );
  inv_x1_sg U48397 ( .A(n58771), .X(n58774) );
  nand_x1_sg U48398 ( .A(n58769), .B(n58768), .X(n42681) );
  inv_x1_sg U48399 ( .A(n58767), .X(n58768) );
  inv_x1_sg U48400 ( .A(n58766), .X(n58769) );
  nand_x1_sg U48401 ( .A(n58764), .B(n58763), .X(n42680) );
  inv_x1_sg U48402 ( .A(n58762), .X(n58763) );
  inv_x1_sg U48403 ( .A(n58761), .X(n58764) );
  nand_x1_sg U48404 ( .A(n32818), .B(n32819), .X(n42823) );
  nand_x1_sg U48405 ( .A(n34224), .B(n34225), .X(n43469) );
  nand_x1_sg U48406 ( .A(n34226), .B(n57167), .X(n34225) );
  nand_x1_sg U48407 ( .A(n32812), .B(n32813), .X(n42820) );
  nand_x1_sg U48408 ( .A(n40871), .B(n32803), .X(n32812) );
  nand_x1_sg U48409 ( .A(n32814), .B(n32815), .X(n42821) );
  nand_x1_sg U48410 ( .A(n40870), .B(n57170), .X(n32814) );
  nand_x1_sg U48411 ( .A(n32823), .B(n32824), .X(n42825) );
  nand_x1_sg U48412 ( .A(n40869), .B(n57170), .X(n32823) );
  nand_x1_sg U48413 ( .A(n32804), .B(n32805), .X(n42816) );
  nand_x1_sg U48414 ( .A(n40868), .B(n57170), .X(n32804) );
  nand_x1_sg U48415 ( .A(n32825), .B(n32826), .X(n42826) );
  nand_x1_sg U48416 ( .A(n40875), .B(n57170), .X(n32825) );
  nand_x1_sg U48417 ( .A(n32816), .B(n32817), .X(n42822) );
  nand_x1_sg U48418 ( .A(n40874), .B(n57170), .X(n32816) );
  nand_x1_sg U48419 ( .A(n32821), .B(n32822), .X(n42824) );
  nand_x1_sg U48420 ( .A(n40873), .B(n57170), .X(n32821) );
  nand_x1_sg U48421 ( .A(n32829), .B(n32830), .X(n42828) );
  nand_x1_sg U48422 ( .A(n40872), .B(n57170), .X(n32829) );
  nand_x1_sg U48423 ( .A(n32827), .B(n32828), .X(n42827) );
  nand_x1_sg U48424 ( .A(n40880), .B(n57170), .X(n32827) );
  nand_x1_sg U48425 ( .A(n32808), .B(n32809), .X(n42818) );
  nand_x1_sg U48426 ( .A(n40879), .B(n57170), .X(n32808) );
  nand_x1_sg U48427 ( .A(n51057), .B(n57294), .X(n32809) );
  nand_x1_sg U48428 ( .A(n32810), .B(n32811), .X(n42819) );
  nand_x1_sg U48429 ( .A(n40878), .B(n57170), .X(n32810) );
  nand_x1_sg U48430 ( .A(n32806), .B(n32807), .X(n42817) );
  nand_x1_sg U48431 ( .A(n40877), .B(n57170), .X(n32806) );
  nand_x1_sg U48432 ( .A(n57310), .B(n57294), .X(n32807) );
  nand_x1_sg U48433 ( .A(n32800), .B(n32801), .X(n42815) );
  nand_x1_sg U48434 ( .A(n40876), .B(n57170), .X(n32800) );
  nand_x1_sg U48435 ( .A(n40220), .B(n40221), .X(\filter_0/n11501 ) );
  nand_x1_sg U48436 ( .A(n57536), .B(n40222), .X(n40220) );
  nand_x1_sg U48437 ( .A(n68336), .B(n40223), .X(n40222) );
  nand_x1_sg U48438 ( .A(n40215), .B(n40216), .X(\filter_0/n11502 ) );
  nand_x1_sg U48439 ( .A(n57558), .B(n40217), .X(n40216) );
  nand_x1_sg U48440 ( .A(n68335), .B(n40218), .X(n40217) );
  nand_x1_sg U48441 ( .A(n40210), .B(n40211), .X(\filter_0/n11503 ) );
  nand_x1_sg U48442 ( .A(n57534), .B(n40212), .X(n40211) );
  nand_x1_sg U48443 ( .A(n68334), .B(n40213), .X(n40212) );
  nand_x1_sg U48444 ( .A(n40205), .B(n40206), .X(\filter_0/n11504 ) );
  nand_x1_sg U48445 ( .A(n57551), .B(n40207), .X(n40206) );
  nand_x1_sg U48446 ( .A(n68333), .B(n40208), .X(n40207) );
  nand_x1_sg U48447 ( .A(n40200), .B(n40201), .X(\filter_0/n11505 ) );
  nand_x1_sg U48448 ( .A(n57558), .B(n40202), .X(n40201) );
  nand_x1_sg U48449 ( .A(n68332), .B(n40203), .X(n40202) );
  nand_x1_sg U48450 ( .A(n40195), .B(n40196), .X(\filter_0/n11506 ) );
  nand_x1_sg U48451 ( .A(n57554), .B(n40197), .X(n40196) );
  nand_x1_sg U48452 ( .A(n68331), .B(n40198), .X(n40197) );
  nand_x1_sg U48453 ( .A(n40190), .B(n40191), .X(\filter_0/n11507 ) );
  nand_x1_sg U48454 ( .A(n57537), .B(n40192), .X(n40191) );
  nand_x1_sg U48455 ( .A(n68330), .B(n40193), .X(n40192) );
  nand_x1_sg U48456 ( .A(n40185), .B(n40186), .X(\filter_0/n11508 ) );
  nand_x1_sg U48457 ( .A(n57558), .B(n40187), .X(n40186) );
  nand_x1_sg U48458 ( .A(n68329), .B(n40188), .X(n40187) );
  nand_x1_sg U48459 ( .A(n40180), .B(n40181), .X(\filter_0/n11509 ) );
  nand_x1_sg U48460 ( .A(n57558), .B(n40182), .X(n40181) );
  nand_x1_sg U48461 ( .A(n68328), .B(n40183), .X(n40182) );
  nand_x1_sg U48462 ( .A(n40175), .B(n40176), .X(\filter_0/n11510 ) );
  nand_x1_sg U48463 ( .A(n57537), .B(n40177), .X(n40176) );
  nand_x1_sg U48464 ( .A(n68327), .B(n40178), .X(n40177) );
  nand_x1_sg U48465 ( .A(n40170), .B(n40171), .X(\filter_0/n11511 ) );
  nand_x1_sg U48466 ( .A(n57552), .B(n40172), .X(n40171) );
  nand_x1_sg U48467 ( .A(n68326), .B(n40173), .X(n40172) );
  nand_x1_sg U48468 ( .A(n40165), .B(n40166), .X(\filter_0/n11512 ) );
  nand_x1_sg U48469 ( .A(n57554), .B(n40167), .X(n40166) );
  nand_x1_sg U48470 ( .A(n68325), .B(n40168), .X(n40167) );
  nand_x1_sg U48471 ( .A(n40160), .B(n40161), .X(\filter_0/n11513 ) );
  nand_x1_sg U48472 ( .A(n57550), .B(n40162), .X(n40161) );
  nand_x1_sg U48473 ( .A(n68324), .B(n40163), .X(n40162) );
  nand_x1_sg U48474 ( .A(n40155), .B(n40156), .X(\filter_0/n11514 ) );
  nand_x1_sg U48475 ( .A(n57558), .B(n40157), .X(n40156) );
  nand_x1_sg U48476 ( .A(n68323), .B(n40158), .X(n40157) );
  nand_x1_sg U48477 ( .A(n40150), .B(n40151), .X(\filter_0/n11515 ) );
  nand_x1_sg U48478 ( .A(n57533), .B(n40152), .X(n40151) );
  nand_x1_sg U48479 ( .A(n68322), .B(n40153), .X(n40152) );
  nand_x1_sg U48480 ( .A(n40145), .B(n40146), .X(\filter_0/n11516 ) );
  nand_x1_sg U48481 ( .A(n57552), .B(n40147), .X(n40146) );
  nand_x1_sg U48482 ( .A(n68321), .B(n40148), .X(n40147) );
  nand_x1_sg U48483 ( .A(n40140), .B(n40141), .X(\filter_0/n11517 ) );
  nand_x1_sg U48484 ( .A(n57550), .B(n40142), .X(n40141) );
  nand_x1_sg U48485 ( .A(n68320), .B(n40143), .X(n40142) );
  nand_x1_sg U48486 ( .A(n40135), .B(n40136), .X(\filter_0/n11518 ) );
  nand_x1_sg U48487 ( .A(n57554), .B(n40137), .X(n40136) );
  nand_x1_sg U48488 ( .A(n68319), .B(n40138), .X(n40137) );
  nand_x1_sg U48489 ( .A(n40130), .B(n40131), .X(\filter_0/n11519 ) );
  nand_x1_sg U48490 ( .A(n57551), .B(n40132), .X(n40131) );
  nand_x1_sg U48491 ( .A(n68318), .B(n40133), .X(n40132) );
  nand_x1_sg U48492 ( .A(n40125), .B(n40126), .X(\filter_0/n11520 ) );
  nand_x1_sg U48493 ( .A(n57533), .B(n40127), .X(n40126) );
  nand_x1_sg U48494 ( .A(n68317), .B(n40128), .X(n40127) );
  nand_x1_sg U48495 ( .A(n40120), .B(n40121), .X(\filter_0/n11521 ) );
  nand_x1_sg U48496 ( .A(n57552), .B(n40122), .X(n40121) );
  nand_x1_sg U48497 ( .A(n68316), .B(n40123), .X(n40122) );
  nand_x1_sg U48498 ( .A(n40115), .B(n40116), .X(\filter_0/n11522 ) );
  nand_x1_sg U48499 ( .A(n57534), .B(n40117), .X(n40116) );
  nand_x1_sg U48500 ( .A(n68315), .B(n40118), .X(n40117) );
  nand_x1_sg U48501 ( .A(n40110), .B(n40111), .X(\filter_0/n11523 ) );
  nand_x1_sg U48502 ( .A(n57557), .B(n40112), .X(n40111) );
  nand_x1_sg U48503 ( .A(n68314), .B(n40113), .X(n40112) );
  nand_x1_sg U48504 ( .A(n40105), .B(n40106), .X(\filter_0/n11524 ) );
  nand_x1_sg U48505 ( .A(n57551), .B(n40107), .X(n40106) );
  nand_x1_sg U48506 ( .A(n68313), .B(n40108), .X(n40107) );
  nand_x1_sg U48507 ( .A(n40100), .B(n40101), .X(\filter_0/n11525 ) );
  nand_x1_sg U48508 ( .A(n57534), .B(n40102), .X(n40101) );
  nand_x1_sg U48509 ( .A(n68312), .B(n40103), .X(n40102) );
  nand_x1_sg U48510 ( .A(n40095), .B(n40096), .X(\filter_0/n11526 ) );
  nand_x1_sg U48511 ( .A(n57535), .B(n40097), .X(n40096) );
  nand_x1_sg U48512 ( .A(n68311), .B(n40098), .X(n40097) );
  nand_x1_sg U48513 ( .A(n40090), .B(n40091), .X(\filter_0/n11527 ) );
  nand_x1_sg U48514 ( .A(n57538), .B(n40092), .X(n40091) );
  nand_x1_sg U48515 ( .A(n68310), .B(n40093), .X(n40092) );
  nand_x1_sg U48516 ( .A(n40085), .B(n40086), .X(\filter_0/n11528 ) );
  nand_x1_sg U48517 ( .A(n57550), .B(n40087), .X(n40086) );
  nand_x1_sg U48518 ( .A(n68309), .B(n40088), .X(n40087) );
  nand_x1_sg U48519 ( .A(n40080), .B(n40081), .X(\filter_0/n11529 ) );
  nand_x1_sg U48520 ( .A(n57554), .B(n40082), .X(n40081) );
  nand_x1_sg U48521 ( .A(n68308), .B(n40083), .X(n40082) );
  nand_x1_sg U48522 ( .A(n40075), .B(n40076), .X(\filter_0/n11530 ) );
  nand_x1_sg U48523 ( .A(n57551), .B(n40077), .X(n40076) );
  nand_x1_sg U48524 ( .A(n68307), .B(n40078), .X(n40077) );
  nand_x1_sg U48525 ( .A(n40070), .B(n40071), .X(\filter_0/n11531 ) );
  nand_x1_sg U48526 ( .A(n57536), .B(n40072), .X(n40071) );
  nand_x1_sg U48527 ( .A(n68306), .B(n40073), .X(n40072) );
  nand_x1_sg U48528 ( .A(n40065), .B(n40066), .X(\filter_0/n11532 ) );
  nand_x1_sg U48529 ( .A(n57551), .B(n40067), .X(n40066) );
  nand_x1_sg U48530 ( .A(n68305), .B(n40068), .X(n40067) );
  nand_x1_sg U48531 ( .A(n40060), .B(n40061), .X(\filter_0/n11533 ) );
  nand_x1_sg U48532 ( .A(n57533), .B(n40062), .X(n40061) );
  nand_x1_sg U48533 ( .A(n68304), .B(n40063), .X(n40062) );
  nand_x1_sg U48534 ( .A(n40055), .B(n40056), .X(\filter_0/n11534 ) );
  nand_x1_sg U48535 ( .A(n57550), .B(n40057), .X(n40056) );
  nand_x1_sg U48536 ( .A(n68303), .B(n40058), .X(n40057) );
  nand_x1_sg U48537 ( .A(n40050), .B(n40051), .X(\filter_0/n11535 ) );
  nand_x1_sg U48538 ( .A(n57534), .B(n40052), .X(n40051) );
  nand_x1_sg U48539 ( .A(n68302), .B(n40053), .X(n40052) );
  nand_x1_sg U48540 ( .A(n40045), .B(n40046), .X(\filter_0/n11536 ) );
  nand_x1_sg U48541 ( .A(n57550), .B(n40047), .X(n40046) );
  nand_x1_sg U48542 ( .A(n68301), .B(n40048), .X(n40047) );
  nand_x1_sg U48543 ( .A(n40040), .B(n40041), .X(\filter_0/n11537 ) );
  nand_x1_sg U48544 ( .A(n57551), .B(n40042), .X(n40041) );
  nand_x1_sg U48545 ( .A(n68300), .B(n40043), .X(n40042) );
  nand_x1_sg U48546 ( .A(n40035), .B(n40036), .X(\filter_0/n11538 ) );
  nand_x1_sg U48547 ( .A(n57551), .B(n40037), .X(n40036) );
  nand_x1_sg U48548 ( .A(n68299), .B(n40038), .X(n40037) );
  nand_x1_sg U48549 ( .A(n40030), .B(n40031), .X(\filter_0/n11539 ) );
  nand_x1_sg U48550 ( .A(n57554), .B(n40032), .X(n40031) );
  nand_x1_sg U48551 ( .A(n68298), .B(n40033), .X(n40032) );
  nand_x1_sg U48552 ( .A(n40025), .B(n40026), .X(\filter_0/n11540 ) );
  nand_x1_sg U48553 ( .A(n57550), .B(n40027), .X(n40026) );
  nand_x1_sg U48554 ( .A(n68297), .B(n40028), .X(n40027) );
  nand_x1_sg U48555 ( .A(n40020), .B(n40021), .X(\filter_0/n11541 ) );
  nand_x1_sg U48556 ( .A(n57533), .B(n40022), .X(n40021) );
  nand_x1_sg U48557 ( .A(n68296), .B(n40023), .X(n40022) );
  nand_x1_sg U48558 ( .A(n40015), .B(n40016), .X(\filter_0/n11542 ) );
  nand_x1_sg U48559 ( .A(n57535), .B(n40017), .X(n40016) );
  nand_x1_sg U48560 ( .A(n68295), .B(n40018), .X(n40017) );
  nand_x1_sg U48561 ( .A(n40010), .B(n40011), .X(\filter_0/n11543 ) );
  nand_x1_sg U48562 ( .A(n57533), .B(n40012), .X(n40011) );
  nand_x1_sg U48563 ( .A(n68294), .B(n40013), .X(n40012) );
  nand_x1_sg U48564 ( .A(n40005), .B(n40006), .X(\filter_0/n11544 ) );
  nand_x1_sg U48565 ( .A(n57550), .B(n40007), .X(n40006) );
  nand_x1_sg U48566 ( .A(n68293), .B(n40008), .X(n40007) );
  nand_x1_sg U48567 ( .A(n40000), .B(n40001), .X(\filter_0/n11545 ) );
  nand_x1_sg U48568 ( .A(n57535), .B(n40002), .X(n40001) );
  nand_x1_sg U48569 ( .A(n68292), .B(n40003), .X(n40002) );
  nand_x1_sg U48570 ( .A(n39995), .B(n39996), .X(\filter_0/n11546 ) );
  nand_x1_sg U48571 ( .A(n57536), .B(n39997), .X(n39996) );
  nand_x1_sg U48572 ( .A(n68291), .B(n39998), .X(n39997) );
  nand_x1_sg U48573 ( .A(n39990), .B(n39991), .X(\filter_0/n11547 ) );
  nand_x1_sg U48574 ( .A(n57533), .B(n39992), .X(n39991) );
  nand_x1_sg U48575 ( .A(n68290), .B(n39993), .X(n39992) );
  nand_x1_sg U48576 ( .A(n39985), .B(n39986), .X(\filter_0/n11548 ) );
  nand_x1_sg U48577 ( .A(n57554), .B(n39987), .X(n39986) );
  nand_x1_sg U48578 ( .A(n68289), .B(n39988), .X(n39987) );
  nand_x1_sg U48579 ( .A(n39980), .B(n39981), .X(\filter_0/n11549 ) );
  nand_x1_sg U48580 ( .A(n57534), .B(n39982), .X(n39981) );
  nand_x1_sg U48581 ( .A(n68288), .B(n39983), .X(n39982) );
  nand_x1_sg U48582 ( .A(n39975), .B(n39976), .X(\filter_0/n11550 ) );
  nand_x1_sg U48583 ( .A(n57534), .B(n39977), .X(n39976) );
  nand_x1_sg U48584 ( .A(n68287), .B(n39978), .X(n39977) );
  nand_x1_sg U48585 ( .A(n39970), .B(n39971), .X(\filter_0/n11551 ) );
  nand_x1_sg U48586 ( .A(n57534), .B(n39972), .X(n39971) );
  nand_x1_sg U48587 ( .A(n68286), .B(n39973), .X(n39972) );
  nand_x1_sg U48588 ( .A(n39965), .B(n39966), .X(\filter_0/n11552 ) );
  nand_x1_sg U48589 ( .A(n57534), .B(n39967), .X(n39966) );
  nand_x1_sg U48590 ( .A(n68285), .B(n39968), .X(n39967) );
  nand_x1_sg U48591 ( .A(n39960), .B(n39961), .X(\filter_0/n11553 ) );
  nand_x1_sg U48592 ( .A(n57558), .B(n39962), .X(n39961) );
  nand_x1_sg U48593 ( .A(n68284), .B(n39963), .X(n39962) );
  nand_x1_sg U48594 ( .A(n39955), .B(n39956), .X(\filter_0/n11554 ) );
  nand_x1_sg U48595 ( .A(n57554), .B(n39957), .X(n39956) );
  nand_x1_sg U48596 ( .A(n68283), .B(n39958), .X(n39957) );
  nand_x1_sg U48597 ( .A(n39950), .B(n39951), .X(\filter_0/n11555 ) );
  nand_x1_sg U48598 ( .A(n57533), .B(n39952), .X(n39951) );
  nand_x1_sg U48599 ( .A(n68282), .B(n39953), .X(n39952) );
  nand_x1_sg U48600 ( .A(n39945), .B(n39946), .X(\filter_0/n11556 ) );
  nand_x1_sg U48601 ( .A(n57551), .B(n39947), .X(n39946) );
  nand_x1_sg U48602 ( .A(n68281), .B(n39948), .X(n39947) );
  nand_x1_sg U48603 ( .A(n39940), .B(n39941), .X(\filter_0/n11557 ) );
  nand_x1_sg U48604 ( .A(n57550), .B(n39942), .X(n39941) );
  nand_x1_sg U48605 ( .A(n68280), .B(n39943), .X(n39942) );
  nand_x1_sg U48606 ( .A(n39935), .B(n39936), .X(\filter_0/n11558 ) );
  nand_x1_sg U48607 ( .A(n57533), .B(n39937), .X(n39936) );
  nand_x1_sg U48608 ( .A(n68279), .B(n39938), .X(n39937) );
  nand_x1_sg U48609 ( .A(n39930), .B(n39931), .X(\filter_0/n11559 ) );
  nand_x1_sg U48610 ( .A(n57558), .B(n39932), .X(n39931) );
  nand_x1_sg U48611 ( .A(n68278), .B(n39933), .X(n39932) );
  nand_x1_sg U48612 ( .A(n39925), .B(n39926), .X(\filter_0/n11560 ) );
  nand_x1_sg U48613 ( .A(n57558), .B(n39927), .X(n39926) );
  nand_x1_sg U48614 ( .A(n68277), .B(n39928), .X(n39927) );
  nand_x1_sg U48615 ( .A(n39920), .B(n39921), .X(\filter_0/n11561 ) );
  nand_x1_sg U48616 ( .A(n57538), .B(n39922), .X(n39921) );
  nand_x1_sg U48617 ( .A(n68276), .B(n39923), .X(n39922) );
  nand_x1_sg U48618 ( .A(n39915), .B(n39916), .X(\filter_0/n11562 ) );
  nand_x1_sg U48619 ( .A(n57553), .B(n39917), .X(n39916) );
  nand_x1_sg U48620 ( .A(n68275), .B(n39918), .X(n39917) );
  nand_x1_sg U48621 ( .A(n39910), .B(n39911), .X(\filter_0/n11563 ) );
  nand_x1_sg U48622 ( .A(n57550), .B(n39912), .X(n39911) );
  nand_x1_sg U48623 ( .A(n68274), .B(n39913), .X(n39912) );
  nand_x1_sg U48624 ( .A(n39905), .B(n39906), .X(\filter_0/n11564 ) );
  nand_x1_sg U48625 ( .A(n57558), .B(n39907), .X(n39906) );
  nand_x1_sg U48626 ( .A(n68273), .B(n39908), .X(n39907) );
  nand_x1_sg U48627 ( .A(n39903), .B(n39904), .X(\filter_0/n11565 ) );
  nand_x1_sg U48628 ( .A(n39901), .B(n39902), .X(\filter_0/n11566 ) );
  nand_x1_sg U48629 ( .A(n39899), .B(n39900), .X(\filter_0/n11567 ) );
  nand_x1_sg U48630 ( .A(n39897), .B(n39898), .X(\filter_0/n11568 ) );
  nand_x1_sg U48631 ( .A(n39895), .B(n39896), .X(\filter_0/n11569 ) );
  nand_x1_sg U48632 ( .A(n39893), .B(n39894), .X(\filter_0/n11570 ) );
  nand_x1_sg U48633 ( .A(n39891), .B(n39892), .X(\filter_0/n11571 ) );
  nand_x1_sg U48634 ( .A(n39889), .B(n39890), .X(\filter_0/n11572 ) );
  nand_x1_sg U48635 ( .A(n39887), .B(n39888), .X(\filter_0/n11573 ) );
  nand_x1_sg U48636 ( .A(n39885), .B(n39886), .X(\filter_0/n11574 ) );
  nand_x1_sg U48637 ( .A(n39883), .B(n39884), .X(\filter_0/n11575 ) );
  nand_x1_sg U48638 ( .A(n39881), .B(n39882), .X(\filter_0/n11576 ) );
  nand_x1_sg U48639 ( .A(n39879), .B(n39880), .X(\filter_0/n11577 ) );
  nand_x1_sg U48640 ( .A(n39877), .B(n39878), .X(\filter_0/n11578 ) );
  nand_x1_sg U48641 ( .A(n39875), .B(n39876), .X(\filter_0/n11579 ) );
  nand_x1_sg U48642 ( .A(n39873), .B(n39874), .X(\filter_0/n11580 ) );
  nand_x1_sg U48643 ( .A(n39871), .B(n39872), .X(\filter_0/n11581 ) );
  nand_x1_sg U48644 ( .A(n39869), .B(n39870), .X(\filter_0/n11582 ) );
  nand_x1_sg U48645 ( .A(n39867), .B(n39868), .X(\filter_0/n11583 ) );
  nand_x1_sg U48646 ( .A(n39865), .B(n39866), .X(\filter_0/n11584 ) );
  nand_x1_sg U48647 ( .A(n39863), .B(n39864), .X(\filter_0/n11585 ) );
  nand_x1_sg U48648 ( .A(n39861), .B(n39862), .X(\filter_0/n11586 ) );
  nand_x1_sg U48649 ( .A(n39859), .B(n39860), .X(\filter_0/n11587 ) );
  nand_x1_sg U48650 ( .A(n39857), .B(n39858), .X(\filter_0/n11588 ) );
  nand_x1_sg U48651 ( .A(n39855), .B(n39856), .X(\filter_0/n11589 ) );
  nand_x1_sg U48652 ( .A(n39853), .B(n39854), .X(\filter_0/n11590 ) );
  nand_x1_sg U48653 ( .A(n39851), .B(n39852), .X(\filter_0/n11591 ) );
  nand_x1_sg U48654 ( .A(n39849), .B(n39850), .X(\filter_0/n11592 ) );
  nand_x1_sg U48655 ( .A(n39847), .B(n39848), .X(\filter_0/n11593 ) );
  nand_x1_sg U48656 ( .A(n39845), .B(n39846), .X(\filter_0/n11594 ) );
  nand_x1_sg U48657 ( .A(n39843), .B(n39844), .X(\filter_0/n11595 ) );
  nand_x1_sg U48658 ( .A(n39841), .B(n39842), .X(\filter_0/n11596 ) );
  nand_x1_sg U48659 ( .A(n35387), .B(n35388), .X(n44048) );
  nand_x1_sg U48660 ( .A(n35381), .B(n35382), .X(n44045) );
  nand_x1_sg U48661 ( .A(n35371), .B(n35372), .X(n44040) );
  nand_x1_sg U48662 ( .A(n35365), .B(n35366), .X(n44037) );
  nand_x1_sg U48663 ( .A(n35323), .B(n35324), .X(n44016) );
  nand_x1_sg U48664 ( .A(n34391), .B(n34392), .X(n43550) );
  nand_x1_sg U48665 ( .A(n35317), .B(n35318), .X(n44013) );
  nand_x1_sg U48666 ( .A(n35311), .B(n35312), .X(n44010) );
  nand_x1_sg U48667 ( .A(n35359), .B(n35360), .X(n44034) );
  nand_x1_sg U48668 ( .A(n35353), .B(n35354), .X(n44031) );
  nand_x1_sg U48669 ( .A(n35337), .B(n35338), .X(n44023) );
  nand_x1_sg U48670 ( .A(n35333), .B(n35334), .X(n44021) );
  nand_x1_sg U48671 ( .A(n35209), .B(n35210), .X(n43959) );
  nand_x1_sg U48672 ( .A(n35197), .B(n35198), .X(n43953) );
  nand_x1_sg U48673 ( .A(n35399), .B(n35400), .X(n44054) );
  nand_x1_sg U48674 ( .A(n35393), .B(n35394), .X(n44051) );
  nand_x1_sg U48675 ( .A(n35283), .B(n35284), .X(n43996) );
  nand_x1_sg U48676 ( .A(n35295), .B(n35296), .X(n44002) );
  nand_x1_sg U48677 ( .A(n35281), .B(n35282), .X(n43995) );
  nand_x1_sg U48678 ( .A(n35275), .B(n35276), .X(n43992) );
  nand_x1_sg U48679 ( .A(n34917), .B(n34918), .X(n43813) );
  nand_x1_sg U48680 ( .A(n34911), .B(n34912), .X(n43810) );
  nand_x1_sg U48681 ( .A(n34905), .B(n34906), .X(n43807) );
  nand_x1_sg U48682 ( .A(n34899), .B(n34900), .X(n43804) );
  nand_x1_sg U48683 ( .A(n34941), .B(n34942), .X(n43825) );
  nand_x1_sg U48684 ( .A(n34953), .B(n34954), .X(n43831) );
  nand_x1_sg U48685 ( .A(n34935), .B(n34936), .X(n43822) );
  nand_x1_sg U48686 ( .A(n34929), .B(n34930), .X(n43819) );
  nand_x1_sg U48687 ( .A(n34985), .B(n34986), .X(n43847) );
  nand_x1_sg U48688 ( .A(n34979), .B(n34980), .X(n43844) );
  nand_x1_sg U48689 ( .A(n34973), .B(n34974), .X(n43841) );
  nand_x1_sg U48690 ( .A(n34969), .B(n34970), .X(n43839) );
  nand_x1_sg U48691 ( .A(n34881), .B(n34882), .X(n43795) );
  nand_x1_sg U48692 ( .A(n34875), .B(n34876), .X(n43792) );
  nand_x1_sg U48693 ( .A(n35021), .B(n35022), .X(n43865) );
  nand_x1_sg U48694 ( .A(n34337), .B(n34338), .X(n43523) );
  nand_x1_sg U48695 ( .A(n34355), .B(n34356), .X(n43532) );
  nand_x1_sg U48696 ( .A(n34353), .B(n34354), .X(n43531) );
  nand_x1_sg U48697 ( .A(n34863), .B(n34864), .X(n43786) );
  nand_x1_sg U48698 ( .A(n34857), .B(n34858), .X(n43783) );
  nand_x1_sg U48699 ( .A(n34821), .B(n34822), .X(n43765) );
  nand_x1_sg U48700 ( .A(n34815), .B(n34816), .X(n43762) );
  nand_x1_sg U48701 ( .A(n34809), .B(n34810), .X(n43759) );
  nand_x1_sg U48702 ( .A(n34803), .B(n34804), .X(n43756) );
  nand_x1_sg U48703 ( .A(n35027), .B(n35028), .X(n43868) );
  nand_x1_sg U48704 ( .A(n34357), .B(n34358), .X(n43533) );
  nand_x1_sg U48705 ( .A(n34335), .B(n34336), .X(n43522) );
  nand_x1_sg U48706 ( .A(n34349), .B(n34350), .X(n43529) );
  nand_x1_sg U48707 ( .A(n34827), .B(n34828), .X(n43768) );
  nand_x1_sg U48708 ( .A(n34839), .B(n34840), .X(n43774) );
  nand_x1_sg U48709 ( .A(n34575), .B(n34576), .X(n43642) );
  nand_x1_sg U48710 ( .A(n34393), .B(n34394), .X(n43551) );
  nand_x1_sg U48711 ( .A(n35139), .B(n35140), .X(n43924) );
  nand_x1_sg U48712 ( .A(n35133), .B(n35134), .X(n43921) );
  nand_x1_sg U48713 ( .A(n35127), .B(n35128), .X(n43918) );
  nand_x1_sg U48714 ( .A(n35121), .B(n35122), .X(n43915) );
  nand_x1_sg U48715 ( .A(n35163), .B(n35164), .X(n43936) );
  nand_x1_sg U48716 ( .A(n35175), .B(n35176), .X(n43942) );
  nand_x1_sg U48717 ( .A(n35157), .B(n35158), .X(n43933) );
  nand_x1_sg U48718 ( .A(n35151), .B(n35152), .X(n43930) );
  nand_x1_sg U48719 ( .A(n35233), .B(n35234), .X(n43971) );
  nand_x1_sg U48720 ( .A(n34379), .B(n34380), .X(n43544) );
  nand_x1_sg U48721 ( .A(n35229), .B(n35230), .X(n43969) );
  nand_x1_sg U48722 ( .A(n35225), .B(n35226), .X(n43967) );
  nand_x1_sg U48723 ( .A(n35269), .B(n35270), .X(n43989) );
  nand_x1_sg U48724 ( .A(n35257), .B(n35258), .X(n43983) );
  nand_x1_sg U48725 ( .A(n35219), .B(n35220), .X(n43964) );
  nand_x1_sg U48726 ( .A(n35203), .B(n35204), .X(n43956) );
  nand_x1_sg U48727 ( .A(n35115), .B(n35116), .X(n43912) );
  nand_x1_sg U48728 ( .A(n34367), .B(n34368), .X(n43538) );
  nand_x1_sg U48729 ( .A(n35109), .B(n35110), .X(n43909) );
  nand_x1_sg U48730 ( .A(n35103), .B(n35104), .X(n43906) );
  nand_x1_sg U48731 ( .A(n35015), .B(n35016), .X(n43862) );
  nand_x1_sg U48732 ( .A(n35009), .B(n35010), .X(n43859) );
  nand_x1_sg U48733 ( .A(n34997), .B(n34998), .X(n43853) );
  nand_x1_sg U48734 ( .A(n34991), .B(n34992), .X(n43850) );
  nand_x1_sg U48735 ( .A(n35049), .B(n35050), .X(n43879) );
  nand_x1_sg U48736 ( .A(n35045), .B(n35046), .X(n43877) );
  nand_x1_sg U48737 ( .A(n35039), .B(n35040), .X(n43874) );
  nand_x1_sg U48738 ( .A(n35033), .B(n35034), .X(n43871) );
  nand_x1_sg U48739 ( .A(n35073), .B(n35074), .X(n43891) );
  nand_x1_sg U48740 ( .A(n35085), .B(n35086), .X(n43897) );
  nand_x1_sg U48741 ( .A(n35067), .B(n35068), .X(n43888) );
  nand_x1_sg U48742 ( .A(n35061), .B(n35062), .X(n43885) );
  nand_x1_sg U48743 ( .A(n34579), .B(n34580), .X(n43644) );
  nand_x1_sg U48744 ( .A(n34577), .B(n34578), .X(n43643) );
  nand_x1_sg U48745 ( .A(n34585), .B(n34586), .X(n43647) );
  nand_x1_sg U48746 ( .A(n34583), .B(n34584), .X(n43646) );
  nand_x1_sg U48747 ( .A(n34567), .B(n34568), .X(n43638) );
  nand_x1_sg U48748 ( .A(n34565), .B(n34566), .X(n43637) );
  nand_x1_sg U48749 ( .A(n34573), .B(n34574), .X(n43641) );
  nand_x1_sg U48750 ( .A(n34571), .B(n34572), .X(n43640) );
  nand_x1_sg U48751 ( .A(n34603), .B(n34604), .X(n43656) );
  nand_x1_sg U48752 ( .A(n34601), .B(n34602), .X(n43655) );
  nand_x1_sg U48753 ( .A(n34609), .B(n34610), .X(n43659) );
  nand_x1_sg U48754 ( .A(n34607), .B(n34608), .X(n43658) );
  nand_x1_sg U48755 ( .A(n34591), .B(n34592), .X(n43650) );
  nand_x1_sg U48756 ( .A(n34589), .B(n34590), .X(n43649) );
  nand_x1_sg U48757 ( .A(n34597), .B(n34598), .X(n43653) );
  nand_x1_sg U48758 ( .A(n34595), .B(n34596), .X(n43652) );
  nand_x1_sg U48759 ( .A(n34531), .B(n34532), .X(n43620) );
  nand_x1_sg U48760 ( .A(n34529), .B(n34530), .X(n43619) );
  nand_x1_sg U48761 ( .A(n34537), .B(n34538), .X(n43623) );
  nand_x1_sg U48762 ( .A(n34535), .B(n34536), .X(n43622) );
  nand_x1_sg U48763 ( .A(n34519), .B(n34520), .X(n43614) );
  nand_x1_sg U48764 ( .A(n34517), .B(n34518), .X(n43613) );
  nand_x1_sg U48765 ( .A(n34525), .B(n34526), .X(n43617) );
  nand_x1_sg U48766 ( .A(n34523), .B(n34524), .X(n43616) );
  nand_x1_sg U48767 ( .A(n34555), .B(n34556), .X(n43632) );
  nand_x1_sg U48768 ( .A(n34553), .B(n34554), .X(n43631) );
  nand_x1_sg U48769 ( .A(n34561), .B(n34562), .X(n43635) );
  nand_x1_sg U48770 ( .A(n34559), .B(n34560), .X(n43634) );
  nand_x1_sg U48771 ( .A(n34543), .B(n34544), .X(n43626) );
  nand_x1_sg U48772 ( .A(n34541), .B(n34542), .X(n43625) );
  nand_x1_sg U48773 ( .A(n34549), .B(n34550), .X(n43629) );
  nand_x1_sg U48774 ( .A(n34547), .B(n34548), .X(n43628) );
  nand_x1_sg U48775 ( .A(n34671), .B(n34672), .X(n43690) );
  nand_x1_sg U48776 ( .A(n34669), .B(n34670), .X(n43689) );
  nand_x1_sg U48777 ( .A(n34677), .B(n34678), .X(n43693) );
  nand_x1_sg U48778 ( .A(n34675), .B(n34676), .X(n43692) );
  nand_x1_sg U48779 ( .A(n34659), .B(n34660), .X(n43684) );
  nand_x1_sg U48780 ( .A(n34657), .B(n34658), .X(n43683) );
  nand_x1_sg U48781 ( .A(n34665), .B(n34666), .X(n43687) );
  nand_x1_sg U48782 ( .A(n34663), .B(n34664), .X(n43686) );
  nand_x1_sg U48783 ( .A(n34693), .B(n34694), .X(n43701) );
  nand_x1_sg U48784 ( .A(n34691), .B(n34692), .X(n43700) );
  nand_x1_sg U48785 ( .A(n34699), .B(n34700), .X(n43704) );
  nand_x1_sg U48786 ( .A(n34697), .B(n34698), .X(n43703) );
  nand_x1_sg U48787 ( .A(n34683), .B(n34684), .X(n43696) );
  nand_x1_sg U48788 ( .A(n34681), .B(n34682), .X(n43695) );
  nand_x1_sg U48789 ( .A(n34689), .B(n34690), .X(n43699) );
  nand_x1_sg U48790 ( .A(n34687), .B(n34688), .X(n43698) );
  nand_x1_sg U48791 ( .A(n34625), .B(n34626), .X(n43667) );
  nand_x1_sg U48792 ( .A(n34623), .B(n34624), .X(n43666) );
  nand_x1_sg U48793 ( .A(n34631), .B(n34632), .X(n43670) );
  nand_x1_sg U48794 ( .A(n34629), .B(n34630), .X(n43669) );
  nand_x1_sg U48795 ( .A(n34613), .B(n34614), .X(n43661) );
  nand_x1_sg U48796 ( .A(n34611), .B(n34612), .X(n43660) );
  nand_x1_sg U48797 ( .A(n34619), .B(n34620), .X(n43664) );
  nand_x1_sg U48798 ( .A(n34617), .B(n34618), .X(n43663) );
  nand_x1_sg U48799 ( .A(n34649), .B(n34650), .X(n43679) );
  nand_x1_sg U48800 ( .A(n34647), .B(n34648), .X(n43678) );
  nand_x1_sg U48801 ( .A(n34655), .B(n34656), .X(n43682) );
  nand_x1_sg U48802 ( .A(n34653), .B(n34654), .X(n43681) );
  nand_x1_sg U48803 ( .A(n34637), .B(n34638), .X(n43673) );
  nand_x1_sg U48804 ( .A(n34635), .B(n34636), .X(n43672) );
  nand_x1_sg U48805 ( .A(n34643), .B(n34644), .X(n43676) );
  nand_x1_sg U48806 ( .A(n34641), .B(n34642), .X(n43675) );
  nand_x1_sg U48807 ( .A(n34303), .B(n34304), .X(n43506) );
  nand_x1_sg U48808 ( .A(n34301), .B(n34302), .X(n43505) );
  nand_x1_sg U48809 ( .A(n34309), .B(n34310), .X(n43509) );
  nand_x1_sg U48810 ( .A(n34307), .B(n34308), .X(n43508) );
  nand_x1_sg U48811 ( .A(n34291), .B(n34292), .X(n43500) );
  nand_x1_sg U48812 ( .A(n34289), .B(n34290), .X(n43499) );
  nand_x1_sg U48813 ( .A(n34297), .B(n34298), .X(n43503) );
  nand_x1_sg U48814 ( .A(n34295), .B(n34296), .X(n43502) );
  nand_x1_sg U48815 ( .A(n34333), .B(n34334), .X(n43521) );
  nand_x1_sg U48816 ( .A(n34331), .B(n34332), .X(n43520) );
  nand_x1_sg U48817 ( .A(n35487), .B(n35488), .X(n44098) );
  nand_x1_sg U48818 ( .A(n35485), .B(n35486), .X(n44097) );
  nand_x1_sg U48819 ( .A(n34387), .B(n34388), .X(n43548) );
  nand_x1_sg U48820 ( .A(n34385), .B(n34386), .X(n43547) );
  nand_x1_sg U48821 ( .A(n35499), .B(n35500), .X(n44104) );
  nand_x1_sg U48822 ( .A(n35497), .B(n35498), .X(n44103) );
  nand_x1_sg U48823 ( .A(n35505), .B(n35506), .X(n44107) );
  nand_x1_sg U48824 ( .A(n35503), .B(n35504), .X(n44106) );
  nand_x1_sg U48825 ( .A(n34401), .B(n34402), .X(n43555) );
  nand_x1_sg U48826 ( .A(n34399), .B(n34400), .X(n43554) );
  nand_x1_sg U48827 ( .A(n35247), .B(n35248), .X(n43978) );
  nand_x1_sg U48828 ( .A(n35237), .B(n35238), .X(n43973) );
  nand_x1_sg U48829 ( .A(n35213), .B(n35214), .X(n43961) );
  nand_x1_sg U48830 ( .A(n35417), .B(n35418), .X(n44063) );
  nand_x1_sg U48831 ( .A(n34375), .B(n34376), .X(n43542) );
  nand_x1_sg U48832 ( .A(n34373), .B(n34374), .X(n43541) );
  nand_x1_sg U48833 ( .A(n35263), .B(n35264), .X(n43986) );
  nand_x1_sg U48834 ( .A(n34397), .B(n34398), .X(n43553) );
  nand_x1_sg U48835 ( .A(n34411), .B(n34412), .X(n43560) );
  nand_x1_sg U48836 ( .A(n34409), .B(n34410), .X(n43559) );
  nand_x1_sg U48837 ( .A(n34417), .B(n34418), .X(n43563) );
  nand_x1_sg U48838 ( .A(n34415), .B(n34416), .X(n43562) );
  nand_x1_sg U48839 ( .A(n34483), .B(n34484), .X(n43596) );
  nand_x1_sg U48840 ( .A(n34481), .B(n34482), .X(n43595) );
  nand_x1_sg U48841 ( .A(n34489), .B(n34490), .X(n43599) );
  nand_x1_sg U48842 ( .A(n34487), .B(n34488), .X(n43598) );
  nand_x1_sg U48843 ( .A(n34471), .B(n34472), .X(n43590) );
  nand_x1_sg U48844 ( .A(n34469), .B(n34470), .X(n43589) );
  nand_x1_sg U48845 ( .A(n34477), .B(n34478), .X(n43593) );
  nand_x1_sg U48846 ( .A(n34475), .B(n34476), .X(n43592) );
  nand_x1_sg U48847 ( .A(n34507), .B(n34508), .X(n43608) );
  nand_x1_sg U48848 ( .A(n34505), .B(n34506), .X(n43607) );
  nand_x1_sg U48849 ( .A(n34513), .B(n34514), .X(n43611) );
  nand_x1_sg U48850 ( .A(n34511), .B(n34512), .X(n43610) );
  nand_x1_sg U48851 ( .A(n34495), .B(n34496), .X(n43602) );
  nand_x1_sg U48852 ( .A(n34493), .B(n34494), .X(n43601) );
  nand_x1_sg U48853 ( .A(n34501), .B(n34502), .X(n43605) );
  nand_x1_sg U48854 ( .A(n34499), .B(n34500), .X(n43604) );
  nand_x1_sg U48855 ( .A(n34435), .B(n34436), .X(n43572) );
  nand_x1_sg U48856 ( .A(n34433), .B(n34434), .X(n43571) );
  nand_x1_sg U48857 ( .A(n34441), .B(n34442), .X(n43575) );
  nand_x1_sg U48858 ( .A(n34439), .B(n34440), .X(n43574) );
  nand_x1_sg U48859 ( .A(n34423), .B(n34424), .X(n43566) );
  nand_x1_sg U48860 ( .A(n34421), .B(n34422), .X(n43565) );
  nand_x1_sg U48861 ( .A(n34429), .B(n34430), .X(n43569) );
  nand_x1_sg U48862 ( .A(n34427), .B(n34428), .X(n43568) );
  nand_x1_sg U48863 ( .A(n34459), .B(n34460), .X(n43584) );
  nand_x1_sg U48864 ( .A(n34457), .B(n34458), .X(n43583) );
  nand_x1_sg U48865 ( .A(n34465), .B(n34466), .X(n43587) );
  nand_x1_sg U48866 ( .A(n34463), .B(n34464), .X(n43586) );
  nand_x1_sg U48867 ( .A(n34447), .B(n34448), .X(n43578) );
  nand_x1_sg U48868 ( .A(n34445), .B(n34446), .X(n43577) );
  nand_x1_sg U48869 ( .A(n34453), .B(n34454), .X(n43581) );
  nand_x1_sg U48870 ( .A(n34451), .B(n34452), .X(n43580) );
  nand_x1_sg U48871 ( .A(n35047), .B(n35048), .X(n43878) );
  nand_x1_sg U48872 ( .A(n34233), .B(n34234), .X(n43471) );
  nand_x1_sg U48873 ( .A(n35053), .B(n35054), .X(n43881) );
  nand_x1_sg U48874 ( .A(n35051), .B(n35052), .X(n43880) );
  nand_x1_sg U48875 ( .A(n35037), .B(n35038), .X(n43873) );
  nand_x1_sg U48876 ( .A(n35035), .B(n35036), .X(n43872) );
  nand_x1_sg U48877 ( .A(n35043), .B(n35044), .X(n43876) );
  nand_x1_sg U48878 ( .A(n35041), .B(n35042), .X(n43875) );
  nand_x1_sg U48879 ( .A(n35071), .B(n35072), .X(n43890) );
  nand_x1_sg U48880 ( .A(n35069), .B(n35070), .X(n43889) );
  nand_x1_sg U48881 ( .A(n35077), .B(n35078), .X(n43893) );
  nand_x1_sg U48882 ( .A(n35075), .B(n35076), .X(n43892) );
  nand_x1_sg U48883 ( .A(n35059), .B(n35060), .X(n43884) );
  nand_x1_sg U48884 ( .A(n35057), .B(n35058), .X(n43883) );
  nand_x1_sg U48885 ( .A(n35065), .B(n35066), .X(n43887) );
  nand_x1_sg U48886 ( .A(n35063), .B(n35064), .X(n43886) );
  nand_x1_sg U48887 ( .A(n35001), .B(n35002), .X(n43855) );
  nand_x1_sg U48888 ( .A(n34999), .B(n35000), .X(n43854) );
  nand_x1_sg U48889 ( .A(n35007), .B(n35008), .X(n43858) );
  nand_x1_sg U48890 ( .A(n35005), .B(n35006), .X(n43857) );
  nand_x1_sg U48891 ( .A(n34989), .B(n34990), .X(n43849) );
  nand_x1_sg U48892 ( .A(n34987), .B(n34988), .X(n43848) );
  nand_x1_sg U48893 ( .A(n34995), .B(n34996), .X(n43852) );
  nand_x1_sg U48894 ( .A(n34993), .B(n34994), .X(n43851) );
  nand_x1_sg U48895 ( .A(n35025), .B(n35026), .X(n43867) );
  nand_x1_sg U48896 ( .A(n35023), .B(n35024), .X(n43866) );
  nand_x1_sg U48897 ( .A(n35031), .B(n35032), .X(n43870) );
  nand_x1_sg U48898 ( .A(n35029), .B(n35030), .X(n43869) );
  nand_x1_sg U48899 ( .A(n35013), .B(n35014), .X(n43861) );
  nand_x1_sg U48900 ( .A(n35011), .B(n35012), .X(n43860) );
  nand_x1_sg U48901 ( .A(n35019), .B(n35020), .X(n43864) );
  nand_x1_sg U48902 ( .A(n35017), .B(n35018), .X(n43863) );
  nand_x1_sg U48903 ( .A(n35143), .B(n35144), .X(n43926) );
  nand_x1_sg U48904 ( .A(n35141), .B(n35142), .X(n43925) );
  nand_x1_sg U48905 ( .A(n35149), .B(n35150), .X(n43929) );
  nand_x1_sg U48906 ( .A(n35147), .B(n35148), .X(n43928) );
  nand_x1_sg U48907 ( .A(n35131), .B(n35132), .X(n43920) );
  nand_x1_sg U48908 ( .A(n35129), .B(n35130), .X(n43919) );
  nand_x1_sg U48909 ( .A(n35137), .B(n35138), .X(n43923) );
  nand_x1_sg U48910 ( .A(n35135), .B(n35136), .X(n43922) );
  nand_x1_sg U48911 ( .A(n35167), .B(n35168), .X(n43938) );
  nand_x1_sg U48912 ( .A(n35165), .B(n35166), .X(n43937) );
  nand_x1_sg U48913 ( .A(n35173), .B(n35174), .X(n43941) );
  nand_x1_sg U48914 ( .A(n35171), .B(n35172), .X(n43940) );
  nand_x1_sg U48915 ( .A(n35155), .B(n35156), .X(n43932) );
  nand_x1_sg U48916 ( .A(n35153), .B(n35154), .X(n43931) );
  nand_x1_sg U48917 ( .A(n35161), .B(n35162), .X(n43935) );
  nand_x1_sg U48918 ( .A(n35159), .B(n35160), .X(n43934) );
  nand_x1_sg U48919 ( .A(n35095), .B(n35096), .X(n43902) );
  nand_x1_sg U48920 ( .A(n35093), .B(n35094), .X(n43901) );
  nand_x1_sg U48921 ( .A(n35101), .B(n35102), .X(n43905) );
  nand_x1_sg U48922 ( .A(n35099), .B(n35100), .X(n43904) );
  nand_x1_sg U48923 ( .A(n35083), .B(n35084), .X(n43896) );
  nand_x1_sg U48924 ( .A(n35081), .B(n35082), .X(n43895) );
  nand_x1_sg U48925 ( .A(n35089), .B(n35090), .X(n43899) );
  nand_x1_sg U48926 ( .A(n35087), .B(n35088), .X(n43898) );
  nand_x1_sg U48927 ( .A(n35119), .B(n35120), .X(n43914) );
  nand_x1_sg U48928 ( .A(n35117), .B(n35118), .X(n43913) );
  nand_x1_sg U48929 ( .A(n35125), .B(n35126), .X(n43917) );
  nand_x1_sg U48930 ( .A(n35123), .B(n35124), .X(n43916) );
  nand_x1_sg U48931 ( .A(n35107), .B(n35108), .X(n43908) );
  nand_x1_sg U48932 ( .A(n35105), .B(n35106), .X(n43907) );
  nand_x1_sg U48933 ( .A(n35113), .B(n35114), .X(n43911) );
  nand_x1_sg U48934 ( .A(n35111), .B(n35112), .X(n43910) );
  nand_x1_sg U48935 ( .A(n34861), .B(n34862), .X(n43785) );
  nand_x1_sg U48936 ( .A(n34859), .B(n34860), .X(n43784) );
  nand_x1_sg U48937 ( .A(n34867), .B(n34868), .X(n43788) );
  nand_x1_sg U48938 ( .A(n34865), .B(n34866), .X(n43787) );
  nand_x1_sg U48939 ( .A(n34849), .B(n34850), .X(n43779) );
  nand_x1_sg U48940 ( .A(n34847), .B(n34848), .X(n43778) );
  nand_x1_sg U48941 ( .A(n34855), .B(n34856), .X(n43782) );
  nand_x1_sg U48942 ( .A(n34853), .B(n34854), .X(n43781) );
  nand_x1_sg U48943 ( .A(n34885), .B(n34886), .X(n43797) );
  nand_x1_sg U48944 ( .A(n34883), .B(n34884), .X(n43796) );
  nand_x1_sg U48945 ( .A(n34891), .B(n34892), .X(n43800) );
  nand_x1_sg U48946 ( .A(n34889), .B(n34890), .X(n43799) );
  nand_x1_sg U48947 ( .A(n34873), .B(n34874), .X(n43791) );
  nand_x1_sg U48948 ( .A(n34871), .B(n34872), .X(n43790) );
  nand_x1_sg U48949 ( .A(n34879), .B(n34880), .X(n43794) );
  nand_x1_sg U48950 ( .A(n34877), .B(n34878), .X(n43793) );
  nand_x1_sg U48951 ( .A(n34813), .B(n34814), .X(n43761) );
  nand_x1_sg U48952 ( .A(n34811), .B(n34812), .X(n43760) );
  nand_x1_sg U48953 ( .A(n34819), .B(n34820), .X(n43764) );
  nand_x1_sg U48954 ( .A(n34817), .B(n34818), .X(n43763) );
  nand_x1_sg U48955 ( .A(n34801), .B(n34802), .X(n43755) );
  nand_x1_sg U48956 ( .A(n34799), .B(n34800), .X(n43754) );
  nand_x1_sg U48957 ( .A(n34807), .B(n34808), .X(n43758) );
  nand_x1_sg U48958 ( .A(n34805), .B(n34806), .X(n43757) );
  nand_x1_sg U48959 ( .A(n34837), .B(n34838), .X(n43773) );
  nand_x1_sg U48960 ( .A(n34835), .B(n34836), .X(n43772) );
  nand_x1_sg U48961 ( .A(n34843), .B(n34844), .X(n43776) );
  nand_x1_sg U48962 ( .A(n34841), .B(n34842), .X(n43775) );
  nand_x1_sg U48963 ( .A(n34825), .B(n34826), .X(n43767) );
  nand_x1_sg U48964 ( .A(n34823), .B(n34824), .X(n43766) );
  nand_x1_sg U48965 ( .A(n34831), .B(n34832), .X(n43770) );
  nand_x1_sg U48966 ( .A(n34829), .B(n34830), .X(n43769) );
  nand_x1_sg U48967 ( .A(n34957), .B(n34958), .X(n43833) );
  nand_x1_sg U48968 ( .A(n34955), .B(n34956), .X(n43832) );
  nand_x1_sg U48969 ( .A(n34963), .B(n34964), .X(n43836) );
  nand_x1_sg U48970 ( .A(n34961), .B(n34962), .X(n43835) );
  nand_x1_sg U48971 ( .A(n34945), .B(n34946), .X(n43827) );
  nand_x1_sg U48972 ( .A(n34943), .B(n34944), .X(n43826) );
  nand_x1_sg U48973 ( .A(n34951), .B(n34952), .X(n43830) );
  nand_x1_sg U48974 ( .A(n34949), .B(n34950), .X(n43829) );
  nand_x1_sg U48975 ( .A(n34977), .B(n34978), .X(n43843) );
  nand_x1_sg U48976 ( .A(n34975), .B(n34976), .X(n43842) );
  nand_x1_sg U48977 ( .A(n34983), .B(n34984), .X(n43846) );
  nand_x1_sg U48978 ( .A(n34981), .B(n34982), .X(n43845) );
  nand_x1_sg U48979 ( .A(n34967), .B(n34968), .X(n43838) );
  nand_x1_sg U48980 ( .A(n34237), .B(n34238), .X(n43473) );
  nand_x1_sg U48981 ( .A(n34971), .B(n34972), .X(n43840) );
  nand_x1_sg U48982 ( .A(n34241), .B(n34242), .X(n43475) );
  nand_x1_sg U48983 ( .A(n34909), .B(n34910), .X(n43809) );
  nand_x1_sg U48984 ( .A(n34907), .B(n34908), .X(n43808) );
  nand_x1_sg U48985 ( .A(n34915), .B(n34916), .X(n43812) );
  nand_x1_sg U48986 ( .A(n34913), .B(n34914), .X(n43811) );
  nand_x1_sg U48987 ( .A(n34897), .B(n34898), .X(n43803) );
  nand_x1_sg U48988 ( .A(n34895), .B(n34896), .X(n43802) );
  nand_x1_sg U48989 ( .A(n34903), .B(n34904), .X(n43806) );
  nand_x1_sg U48990 ( .A(n34901), .B(n34902), .X(n43805) );
  nand_x1_sg U48991 ( .A(n34933), .B(n34934), .X(n43821) );
  nand_x1_sg U48992 ( .A(n34931), .B(n34932), .X(n43820) );
  nand_x1_sg U48993 ( .A(n34939), .B(n34940), .X(n43824) );
  nand_x1_sg U48994 ( .A(n34937), .B(n34938), .X(n43823) );
  nand_x1_sg U48995 ( .A(n34921), .B(n34922), .X(n43815) );
  nand_x1_sg U48996 ( .A(n34919), .B(n34920), .X(n43814) );
  nand_x1_sg U48997 ( .A(n34927), .B(n34928), .X(n43818) );
  nand_x1_sg U48998 ( .A(n34925), .B(n34926), .X(n43817) );
  nand_x1_sg U48999 ( .A(n35403), .B(n35404), .X(n44056) );
  nand_x1_sg U49000 ( .A(n35401), .B(n35402), .X(n44055) );
  nand_x1_sg U49001 ( .A(n35409), .B(n35410), .X(n44059) );
  nand_x1_sg U49002 ( .A(n35407), .B(n35408), .X(n44058) );
  nand_x1_sg U49003 ( .A(n35391), .B(n35392), .X(n44050) );
  nand_x1_sg U49004 ( .A(n35389), .B(n35390), .X(n44049) );
  nand_x1_sg U49005 ( .A(n35397), .B(n35398), .X(n44053) );
  nand_x1_sg U49006 ( .A(n35395), .B(n35396), .X(n44052) );
  nand_x1_sg U49007 ( .A(n35427), .B(n35428), .X(n44068) );
  nand_x1_sg U49008 ( .A(n35425), .B(n35426), .X(n44067) );
  nand_x1_sg U49009 ( .A(n35433), .B(n35434), .X(n44071) );
  nand_x1_sg U49010 ( .A(n35431), .B(n35432), .X(n44070) );
  nand_x1_sg U49011 ( .A(n35415), .B(n35416), .X(n44062) );
  nand_x1_sg U49012 ( .A(n35413), .B(n35414), .X(n44061) );
  nand_x1_sg U49013 ( .A(n35421), .B(n35422), .X(n44065) );
  nand_x1_sg U49014 ( .A(n35419), .B(n35420), .X(n44064) );
  nand_x1_sg U49015 ( .A(n35357), .B(n35358), .X(n44033) );
  nand_x1_sg U49016 ( .A(n35355), .B(n35356), .X(n44032) );
  nand_x1_sg U49017 ( .A(n35363), .B(n35364), .X(n44036) );
  nand_x1_sg U49018 ( .A(n35361), .B(n35362), .X(n44035) );
  nand_x1_sg U49019 ( .A(n35345), .B(n35346), .X(n44027) );
  nand_x1_sg U49020 ( .A(n35343), .B(n35344), .X(n44026) );
  nand_x1_sg U49021 ( .A(n35351), .B(n35352), .X(n44030) );
  nand_x1_sg U49022 ( .A(n35349), .B(n35350), .X(n44029) );
  nand_x1_sg U49023 ( .A(n35379), .B(n35380), .X(n44044) );
  nand_x1_sg U49024 ( .A(n35377), .B(n35378), .X(n44043) );
  nand_x1_sg U49025 ( .A(n35385), .B(n35386), .X(n44047) );
  nand_x1_sg U49026 ( .A(n35383), .B(n35384), .X(n44046) );
  nand_x1_sg U49027 ( .A(n35369), .B(n35370), .X(n44039) );
  nand_x1_sg U49028 ( .A(n35367), .B(n35368), .X(n44038) );
  nand_x1_sg U49029 ( .A(n35375), .B(n35376), .X(n44042) );
  nand_x1_sg U49030 ( .A(n35373), .B(n35374), .X(n44041) );
  nand_x1_sg U49031 ( .A(n35461), .B(n35462), .X(n44085) );
  nand_x1_sg U49032 ( .A(n35459), .B(n35460), .X(n44084) );
  nand_x1_sg U49033 ( .A(n35439), .B(n35440), .X(n44074) );
  nand_x1_sg U49034 ( .A(n35467), .B(n35468), .X(n44088) );
  nand_x1_sg U49035 ( .A(n35465), .B(n35466), .X(n44087) );
  nand_x1_sg U49036 ( .A(n35463), .B(n35464), .X(n44086) );
  nand_x1_sg U49037 ( .A(n35471), .B(n35472), .X(n44090) );
  nand_x1_sg U49038 ( .A(n35469), .B(n35470), .X(n44089) );
  nand_x1_sg U49039 ( .A(n35493), .B(n35494), .X(n44101) );
  nand_x1_sg U49040 ( .A(n35491), .B(n35492), .X(n44100) );
  nand_x1_sg U49041 ( .A(n35473), .B(n35474), .X(n44091) );
  nand_x1_sg U49042 ( .A(n35489), .B(n35490), .X(n44099) );
  nand_x1_sg U49043 ( .A(n35477), .B(n35478), .X(n44093) );
  nand_x1_sg U49044 ( .A(n35475), .B(n35476), .X(n44092) );
  nand_x1_sg U49045 ( .A(n35481), .B(n35482), .X(n44095) );
  nand_x1_sg U49046 ( .A(n35479), .B(n35480), .X(n44094) );
  nand_x1_sg U49047 ( .A(n35429), .B(n35430), .X(n44069) );
  nand_x1_sg U49048 ( .A(n35437), .B(n35438), .X(n44073) );
  nand_x1_sg U49049 ( .A(n35445), .B(n35446), .X(n44077) );
  nand_x1_sg U49050 ( .A(n35443), .B(n35444), .X(n44076) );
  nand_x1_sg U49051 ( .A(n35423), .B(n35424), .X(n44066) );
  nand_x1_sg U49052 ( .A(n34363), .B(n34364), .X(n43536) );
  nand_x1_sg U49053 ( .A(n34361), .B(n34362), .X(n43535) );
  nand_x1_sg U49054 ( .A(n34359), .B(n34360), .X(n43534) );
  nand_x1_sg U49055 ( .A(n35435), .B(n35436), .X(n44072) );
  nand_x1_sg U49056 ( .A(n35453), .B(n35454), .X(n44081) );
  nand_x1_sg U49057 ( .A(n35457), .B(n35458), .X(n44083) );
  nand_x1_sg U49058 ( .A(n35455), .B(n35456), .X(n44082) );
  nand_x1_sg U49059 ( .A(n35451), .B(n35452), .X(n44080) );
  nand_x1_sg U49060 ( .A(n35449), .B(n35450), .X(n44079) );
  nand_x1_sg U49061 ( .A(n35441), .B(n35442), .X(n44075) );
  nand_x1_sg U49062 ( .A(n35447), .B(n35448), .X(n44078) );
  nand_x1_sg U49063 ( .A(n35231), .B(n35232), .X(n43970) );
  nand_x1_sg U49064 ( .A(n34245), .B(n34246), .X(n43477) );
  nand_x1_sg U49065 ( .A(n34230), .B(n34231), .X(n43470) );
  nand_x1_sg U49066 ( .A(n35235), .B(n35236), .X(n43972) );
  nand_x1_sg U49067 ( .A(n35223), .B(n35224), .X(n43966) );
  nand_x1_sg U49068 ( .A(n35221), .B(n35222), .X(n43965) );
  nand_x1_sg U49069 ( .A(n35227), .B(n35228), .X(n43968) );
  nand_x1_sg U49070 ( .A(n34259), .B(n34260), .X(n43484) );
  nand_x1_sg U49071 ( .A(n35249), .B(n35250), .X(n43979) );
  nand_x1_sg U49072 ( .A(n34255), .B(n34256), .X(n43482) );
  nand_x1_sg U49073 ( .A(n35255), .B(n35256), .X(n43982) );
  nand_x1_sg U49074 ( .A(n35253), .B(n35254), .X(n43981) );
  nand_x1_sg U49075 ( .A(n35239), .B(n35240), .X(n43974) );
  nand_x1_sg U49076 ( .A(n34257), .B(n34258), .X(n43483) );
  nand_x1_sg U49077 ( .A(n35245), .B(n35246), .X(n43977) );
  nand_x1_sg U49078 ( .A(n35243), .B(n35244), .X(n43976) );
  nand_x1_sg U49079 ( .A(n35189), .B(n35190), .X(n43949) );
  nand_x1_sg U49080 ( .A(n34251), .B(n34252), .X(n43480) );
  nand_x1_sg U49081 ( .A(n35195), .B(n35196), .X(n43952) );
  nand_x1_sg U49082 ( .A(n35193), .B(n35194), .X(n43951) );
  nand_x1_sg U49083 ( .A(n35179), .B(n35180), .X(n43944) );
  nand_x1_sg U49084 ( .A(n35177), .B(n35178), .X(n43943) );
  nand_x1_sg U49085 ( .A(n35185), .B(n35186), .X(n43947) );
  nand_x1_sg U49086 ( .A(n35183), .B(n35184), .X(n43946) );
  nand_x1_sg U49087 ( .A(n34235), .B(n34236), .X(n43472) );
  nand_x1_sg U49088 ( .A(n35211), .B(n35212), .X(n43960) );
  nand_x1_sg U49089 ( .A(n35217), .B(n35218), .X(n43963) );
  nand_x1_sg U49090 ( .A(n35215), .B(n35216), .X(n43962) );
  nand_x1_sg U49091 ( .A(n35201), .B(n35202), .X(n43955) );
  nand_x1_sg U49092 ( .A(n35199), .B(n35200), .X(n43954) );
  nand_x1_sg U49093 ( .A(n35207), .B(n35208), .X(n43958) );
  nand_x1_sg U49094 ( .A(n35205), .B(n35206), .X(n43957) );
  nand_x1_sg U49095 ( .A(n35315), .B(n35316), .X(n44012) );
  nand_x1_sg U49096 ( .A(n35313), .B(n35314), .X(n44011) );
  nand_x1_sg U49097 ( .A(n35321), .B(n35322), .X(n44015) );
  nand_x1_sg U49098 ( .A(n35319), .B(n35320), .X(n44014) );
  nand_x1_sg U49099 ( .A(n35305), .B(n35306), .X(n44007) );
  nand_x1_sg U49100 ( .A(n35303), .B(n35304), .X(n44006) );
  nand_x1_sg U49101 ( .A(n35309), .B(n35310), .X(n44009) );
  nand_x1_sg U49102 ( .A(n34249), .B(n34250), .X(n43479) );
  nand_x1_sg U49103 ( .A(n35335), .B(n35336), .X(n44022) );
  nand_x1_sg U49104 ( .A(n34253), .B(n34254), .X(n43481) );
  nand_x1_sg U49105 ( .A(n35339), .B(n35340), .X(n44024) );
  nand_x1_sg U49106 ( .A(n34243), .B(n34244), .X(n43476) );
  nand_x1_sg U49107 ( .A(n35325), .B(n35326), .X(n44017) );
  nand_x1_sg U49108 ( .A(n34247), .B(n34248), .X(n43478) );
  nand_x1_sg U49109 ( .A(n35331), .B(n35332), .X(n44020) );
  nand_x1_sg U49110 ( .A(n35329), .B(n35330), .X(n44019) );
  nand_x1_sg U49111 ( .A(n35273), .B(n35274), .X(n43991) );
  nand_x1_sg U49112 ( .A(n35271), .B(n35272), .X(n43990) );
  nand_x1_sg U49113 ( .A(n35279), .B(n35280), .X(n43994) );
  nand_x1_sg U49114 ( .A(n35277), .B(n35278), .X(n43993) );
  nand_x1_sg U49115 ( .A(n35261), .B(n35262), .X(n43985) );
  nand_x1_sg U49116 ( .A(n35259), .B(n35260), .X(n43984) );
  nand_x1_sg U49117 ( .A(n35267), .B(n35268), .X(n43988) );
  nand_x1_sg U49118 ( .A(n35265), .B(n35266), .X(n43987) );
  nand_x1_sg U49119 ( .A(n35293), .B(n35294), .X(n44001) );
  nand_x1_sg U49120 ( .A(n35291), .B(n35292), .X(n44000) );
  nand_x1_sg U49121 ( .A(n35299), .B(n35300), .X(n44004) );
  nand_x1_sg U49122 ( .A(n35297), .B(n35298), .X(n44003) );
  nand_x1_sg U49123 ( .A(n34269), .B(n34270), .X(n43489) );
  nand_x1_sg U49124 ( .A(n34267), .B(n34268), .X(n43488) );
  nand_x1_sg U49125 ( .A(n35287), .B(n35288), .X(n43998) );
  nand_x1_sg U49126 ( .A(n35285), .B(n35286), .X(n43997) );
  nand_x1_sg U49127 ( .A(n34707), .B(n34708), .X(n43708) );
  nand_x1_sg U49128 ( .A(n34701), .B(n34702), .X(n43705) );
  nand_x1_sg U49129 ( .A(n34271), .B(n34272), .X(n43490) );
  nand_x1_sg U49130 ( .A(n34713), .B(n34714), .X(n43711) );
  nand_x1_sg U49131 ( .A(n34725), .B(n34726), .X(n43717) );
  nand_x1_sg U49132 ( .A(n34719), .B(n34720), .X(n43714) );
  nand_x1_sg U49133 ( .A(n34581), .B(n34582), .X(n43645) );
  nand_x1_sg U49134 ( .A(n34605), .B(n34606), .X(n43657) );
  nand_x1_sg U49135 ( .A(n34569), .B(n34570), .X(n43639) );
  nand_x1_sg U49136 ( .A(n34563), .B(n34564), .X(n43636) );
  nand_x1_sg U49137 ( .A(n34557), .B(n34558), .X(n43633) );
  nand_x1_sg U49138 ( .A(n34551), .B(n34552), .X(n43630) );
  nand_x1_sg U49139 ( .A(n34599), .B(n34600), .X(n43654) );
  nand_x1_sg U49140 ( .A(n34615), .B(n34616), .X(n43662) );
  nand_x1_sg U49141 ( .A(n34593), .B(n34594), .X(n43651) );
  nand_x1_sg U49142 ( .A(n34587), .B(n34588), .X(n43648) );
  nand_x1_sg U49143 ( .A(n34341), .B(n34342), .X(n43525) );
  nand_x1_sg U49144 ( .A(n34343), .B(n34344), .X(n43526) );
  nand_x1_sg U49145 ( .A(n34533), .B(n34534), .X(n43621) );
  nand_x1_sg U49146 ( .A(n34527), .B(n34528), .X(n43618) );
  nand_x1_sg U49147 ( .A(n34479), .B(n34480), .X(n43594) );
  nand_x1_sg U49148 ( .A(n34345), .B(n34346), .X(n43527) );
  nand_x1_sg U49149 ( .A(n34485), .B(n34486), .X(n43597) );
  nand_x1_sg U49150 ( .A(n34461), .B(n34462), .X(n43585) );
  nand_x1_sg U49151 ( .A(n34497), .B(n34498), .X(n43603) );
  nand_x1_sg U49152 ( .A(n34515), .B(n34516), .X(n43612) );
  nand_x1_sg U49153 ( .A(n34545), .B(n34546), .X(n43627) );
  nand_x1_sg U49154 ( .A(n34521), .B(n34522), .X(n43615) );
  nand_x1_sg U49155 ( .A(n34503), .B(n34504), .X(n43606) );
  nand_x1_sg U49156 ( .A(n34509), .B(n34510), .X(n43609) );
  nand_x1_sg U49157 ( .A(n34539), .B(n34540), .X(n43624) );
  nand_x1_sg U49158 ( .A(n34491), .B(n34492), .X(n43600) );
  nand_x1_sg U49159 ( .A(n35509), .B(n35510), .X(n44109) );
  nand_x1_sg U49160 ( .A(n34887), .B(n34888), .X(n43798) );
  nand_x1_sg U49161 ( .A(n34869), .B(n34870), .X(n43789) );
  nand_x1_sg U49162 ( .A(n35405), .B(n35406), .X(n44057) );
  nand_x1_sg U49163 ( .A(n35341), .B(n35342), .X(n44025) );
  nand_x1_sg U49164 ( .A(n35507), .B(n35508), .X(n44108) );
  nand_x1_sg U49165 ( .A(n34673), .B(n34674), .X(n43691) );
  nand_x1_sg U49166 ( .A(n34695), .B(n34696), .X(n43702) );
  nand_x1_sg U49167 ( .A(n35181), .B(n35182), .X(n43945) );
  nand_x1_sg U49168 ( .A(n34389), .B(n34390), .X(n43549) );
  nand_x1_sg U49169 ( .A(n35307), .B(n35308), .X(n44008) );
  nand_x1_sg U49170 ( .A(n35097), .B(n35098), .X(n43903) );
  nand_x1_sg U49171 ( .A(n35301), .B(n35302), .X(n44005) );
  nand_x1_sg U49172 ( .A(n35289), .B(n35290), .X(n43999) );
  nand_x1_sg U49173 ( .A(n35327), .B(n35328), .X(n44018) );
  nand_x1_sg U49174 ( .A(n35347), .B(n35348), .X(n44028) );
  nand_x1_sg U49175 ( .A(n34621), .B(n34622), .X(n43665) );
  nand_x1_sg U49176 ( .A(n34667), .B(n34668), .X(n43688) );
  nand_x1_sg U49177 ( .A(n34645), .B(n34646), .X(n43677) );
  nand_x1_sg U49178 ( .A(n34627), .B(n34628), .X(n43668) );
  nand_x1_sg U49179 ( .A(n34661), .B(n34662), .X(n43685) );
  nand_x1_sg U49180 ( .A(n34239), .B(n34240), .X(n43474) );
  nand_x1_sg U49181 ( .A(n34639), .B(n34640), .X(n43674) );
  nand_x1_sg U49182 ( .A(n34633), .B(n34634), .X(n43671) );
  nand_x1_sg U49183 ( .A(n34263), .B(n34264), .X(n43486) );
  nand_x1_sg U49184 ( .A(n34261), .B(n34262), .X(n43485) );
  nand_x1_sg U49185 ( .A(n34685), .B(n34686), .X(n43697) );
  nand_x1_sg U49186 ( .A(n34679), .B(n34680), .X(n43694) );
  nand_x1_sg U49187 ( .A(n34651), .B(n34652), .X(n43680) );
  nand_x1_sg U49188 ( .A(n34265), .B(n34266), .X(n43487) );
  nand_x1_sg U49189 ( .A(n35003), .B(n35004), .X(n43856) );
  nand_x1_sg U49190 ( .A(n34369), .B(n34370), .X(n43539) );
  nand_x1_sg U49191 ( .A(n35169), .B(n35170), .X(n43939) );
  nand_x1_sg U49192 ( .A(n35091), .B(n35092), .X(n43900) );
  nand_x1_sg U49193 ( .A(n35055), .B(n35056), .X(n43882) );
  nand_x1_sg U49194 ( .A(n35079), .B(n35080), .X(n43894) );
  nand_x1_sg U49195 ( .A(n35191), .B(n35192), .X(n43950) );
  nand_x1_sg U49196 ( .A(n34277), .B(n34278), .X(n43493) );
  nand_x1_sg U49197 ( .A(n34381), .B(n34382), .X(n43545) );
  nand_x1_sg U49198 ( .A(n35187), .B(n35188), .X(n43948) );
  nand_x1_sg U49199 ( .A(n34413), .B(n34414), .X(n43561) );
  nand_x1_sg U49200 ( .A(n34283), .B(n34284), .X(n43496) );
  nand_x1_sg U49201 ( .A(n34407), .B(n34408), .X(n43558) );
  nand_x1_sg U49202 ( .A(n35251), .B(n35252), .X(n43980) );
  nand_x1_sg U49203 ( .A(n34285), .B(n34286), .X(n43497) );
  nand_x1_sg U49204 ( .A(n35501), .B(n35502), .X(n44105) );
  nand_x1_sg U49205 ( .A(n34281), .B(n34282), .X(n43495) );
  nand_x1_sg U49206 ( .A(n34965), .B(n34966), .X(n43837) );
  nand_x1_sg U49207 ( .A(n34755), .B(n34756), .X(n43732) );
  nand_x1_sg U49208 ( .A(n34749), .B(n34750), .X(n43729) );
  nand_x1_sg U49209 ( .A(n34743), .B(n34744), .X(n43726) );
  nand_x1_sg U49210 ( .A(n34737), .B(n34738), .X(n43723) );
  nand_x1_sg U49211 ( .A(n34779), .B(n34780), .X(n43744) );
  nand_x1_sg U49212 ( .A(n34791), .B(n34792), .X(n43750) );
  nand_x1_sg U49213 ( .A(n34773), .B(n34774), .X(n43741) );
  nand_x1_sg U49214 ( .A(n34767), .B(n34768), .X(n43738) );
  nand_x1_sg U49215 ( .A(n34845), .B(n34846), .X(n43777) );
  nand_x1_sg U49216 ( .A(n35241), .B(n35242), .X(n43975) );
  nand_x1_sg U49217 ( .A(n34833), .B(n34834), .X(n43771) );
  nand_x1_sg U49218 ( .A(n34851), .B(n34852), .X(n43780) );
  nand_x1_sg U49219 ( .A(n34959), .B(n34960), .X(n43834) );
  nand_x1_sg U49220 ( .A(n34893), .B(n34894), .X(n43801) );
  nand_x1_sg U49221 ( .A(n34923), .B(n34924), .X(n43816) );
  nand_x1_sg U49222 ( .A(n34947), .B(n34948), .X(n43828) );
  nand_x1_sg U49223 ( .A(n34425), .B(n34426), .X(n43567) );
  nand_x1_sg U49224 ( .A(n34321), .B(n34322), .X(n43515) );
  nand_x1_sg U49225 ( .A(n34419), .B(n34420), .X(n43564) );
  nand_x1_sg U49226 ( .A(n35483), .B(n35484), .X(n44096) );
  nand_x1_sg U49227 ( .A(n34317), .B(n34318), .X(n43513) );
  nand_x1_sg U49228 ( .A(n34319), .B(n34320), .X(n43514) );
  nand_x1_sg U49229 ( .A(n34443), .B(n34444), .X(n43576) );
  nand_x1_sg U49230 ( .A(n34437), .B(n34438), .X(n43573) );
  nand_x1_sg U49231 ( .A(n34323), .B(n34324), .X(n43516) );
  nand_x1_sg U49232 ( .A(n34325), .B(n34326), .X(n43517) );
  nand_x1_sg U49233 ( .A(n34473), .B(n34474), .X(n43591) );
  nand_x1_sg U49234 ( .A(n34467), .B(n34468), .X(n43588) );
  nand_x1_sg U49235 ( .A(n34449), .B(n34450), .X(n43579) );
  nand_x1_sg U49236 ( .A(n34327), .B(n34328), .X(n43518) );
  nand_x1_sg U49237 ( .A(n34455), .B(n34456), .X(n43582) );
  nand_x1_sg U49238 ( .A(n34431), .B(n34432), .X(n43570) );
  nand_x1_sg U49239 ( .A(n35411), .B(n35412), .X(n44060) );
  nand_x1_sg U49240 ( .A(n34311), .B(n34312), .X(n43510) );
  nand_x1_sg U49241 ( .A(n34329), .B(n34330), .X(n43519) );
  nand_x1_sg U49242 ( .A(n34313), .B(n34314), .X(n43511) );
  nand_x1_sg U49243 ( .A(n34403), .B(n34404), .X(n43556) );
  nand_x1_sg U49244 ( .A(n34315), .B(n34316), .X(n43512) );
  nand_x1_sg U49245 ( .A(n34395), .B(n34396), .X(n43552) );
  nand_x1_sg U49246 ( .A(n34377), .B(n34378), .X(n43543) );
  nand_x1_sg U49247 ( .A(n35495), .B(n35496), .X(n44102) );
  nand_x1_sg U49248 ( .A(n34293), .B(n34294), .X(n43501) );
  nand_x1_sg U49249 ( .A(n34299), .B(n34300), .X(n43504) );
  nand_x1_sg U49250 ( .A(n34371), .B(n34372), .X(n43540) );
  nand_x1_sg U49251 ( .A(n34383), .B(n34384), .X(n43546) );
  nand_x1_sg U49252 ( .A(n34305), .B(n34306), .X(n43507) );
  nand_x1_sg U49253 ( .A(n34287), .B(n34288), .X(n43498) );
  nand_x1_sg U49254 ( .A(n34405), .B(n34406), .X(n43557) );
  nand_x1_sg U49255 ( .A(n34765), .B(n34766), .X(n43737) );
  nand_x1_sg U49256 ( .A(n34763), .B(n34764), .X(n43736) );
  nand_x1_sg U49257 ( .A(n34771), .B(n34772), .X(n43740) );
  nand_x1_sg U49258 ( .A(n34769), .B(n34770), .X(n43739) );
  nand_x1_sg U49259 ( .A(n34753), .B(n34754), .X(n43731) );
  nand_x1_sg U49260 ( .A(n34751), .B(n34752), .X(n43730) );
  nand_x1_sg U49261 ( .A(n34759), .B(n34760), .X(n43734) );
  nand_x1_sg U49262 ( .A(n34757), .B(n34758), .X(n43733) );
  nand_x1_sg U49263 ( .A(n34789), .B(n34790), .X(n43749) );
  nand_x1_sg U49264 ( .A(n34787), .B(n34788), .X(n43748) );
  nand_x1_sg U49265 ( .A(n34795), .B(n34796), .X(n43752) );
  nand_x1_sg U49266 ( .A(n34793), .B(n34794), .X(n43751) );
  nand_x1_sg U49267 ( .A(n34777), .B(n34778), .X(n43743) );
  nand_x1_sg U49268 ( .A(n34775), .B(n34776), .X(n43742) );
  nand_x1_sg U49269 ( .A(n34783), .B(n34784), .X(n43746) );
  nand_x1_sg U49270 ( .A(n34781), .B(n34782), .X(n43745) );
  nand_x1_sg U49271 ( .A(n34717), .B(n34718), .X(n43713) );
  nand_x1_sg U49272 ( .A(n34715), .B(n34716), .X(n43712) );
  nand_x1_sg U49273 ( .A(n34723), .B(n34724), .X(n43716) );
  nand_x1_sg U49274 ( .A(n34721), .B(n34722), .X(n43715) );
  nand_x1_sg U49275 ( .A(n34705), .B(n34706), .X(n43707) );
  nand_x1_sg U49276 ( .A(n34703), .B(n34704), .X(n43706) );
  nand_x1_sg U49277 ( .A(n34711), .B(n34712), .X(n43710) );
  nand_x1_sg U49278 ( .A(n34709), .B(n34710), .X(n43709) );
  nand_x1_sg U49279 ( .A(n34741), .B(n34742), .X(n43725) );
  nand_x1_sg U49280 ( .A(n34739), .B(n34740), .X(n43724) );
  nand_x1_sg U49281 ( .A(n34747), .B(n34748), .X(n43728) );
  nand_x1_sg U49282 ( .A(n34745), .B(n34746), .X(n43727) );
  nand_x1_sg U49283 ( .A(n34729), .B(n34730), .X(n43719) );
  nand_x1_sg U49284 ( .A(n34727), .B(n34728), .X(n43718) );
  nand_x1_sg U49285 ( .A(n34735), .B(n34736), .X(n43722) );
  nand_x1_sg U49286 ( .A(n34733), .B(n34734), .X(n43721) );
  nand_x1_sg U49287 ( .A(n34347), .B(n34348), .X(n43528) );
  nand_x1_sg U49288 ( .A(n34273), .B(n34274), .X(n43491) );
  nand_x1_sg U49289 ( .A(n34797), .B(n34798), .X(n43753) );
  nand_x1_sg U49290 ( .A(n34339), .B(n34340), .X(n43524) );
  nand_x1_sg U49291 ( .A(n35145), .B(n35146), .X(n43927) );
  nand_x1_sg U49292 ( .A(n34275), .B(n34276), .X(n43492) );
  nand_x1_sg U49293 ( .A(n34365), .B(n34366), .X(n43537) );
  nand_x1_sg U49294 ( .A(n34279), .B(n34280), .X(n43494) );
  nand_x1_sg U49295 ( .A(n34761), .B(n34762), .X(n43735) );
  nand_x1_sg U49296 ( .A(n34785), .B(n34786), .X(n43747) );
  nand_x1_sg U49297 ( .A(n34731), .B(n34732), .X(n43720) );
  nand_x1_sg U49298 ( .A(n34351), .B(n34352), .X(n43530) );
  nand_x1_sg U49299 ( .A(n39839), .B(n39840), .X(\filter_0/n12237 ) );
  nand_x1_sg U49300 ( .A(n34140), .B(n34141), .X(n43432) );
  nand_x1_sg U49301 ( .A(n40518), .B(n57178), .X(n34141) );
  nand_x1_sg U49302 ( .A(n34156), .B(n34157), .X(n43440) );
  nand_x1_sg U49303 ( .A(n40517), .B(n57178), .X(n34157) );
  nand_x1_sg U49304 ( .A(n34136), .B(n34137), .X(n43430) );
  nand_x1_sg U49305 ( .A(n40516), .B(n57178), .X(n34137) );
  nand_x1_sg U49306 ( .A(n34146), .B(n34147), .X(n43435) );
  nand_x1_sg U49307 ( .A(n40515), .B(n57178), .X(n34147) );
  nand_x1_sg U49308 ( .A(n34160), .B(n34161), .X(n43442) );
  nand_x1_sg U49309 ( .A(n40514), .B(n57178), .X(n34161) );
  nand_x1_sg U49310 ( .A(n34144), .B(n34145), .X(n43434) );
  nand_x1_sg U49311 ( .A(n40513), .B(n57178), .X(n34145) );
  nand_x1_sg U49312 ( .A(n34150), .B(n34151), .X(n43437) );
  nand_x1_sg U49313 ( .A(n40512), .B(n34134), .X(n34151) );
  nand_x1_sg U49314 ( .A(n34154), .B(n34155), .X(n43439) );
  nand_x1_sg U49315 ( .A(n40511), .B(n57178), .X(n34155) );
  nand_x1_sg U49316 ( .A(n34162), .B(n34163), .X(n43443) );
  nand_x1_sg U49317 ( .A(n40510), .B(n57178), .X(n34163) );
  nand_x1_sg U49318 ( .A(n34164), .B(n34165), .X(n43444) );
  nand_x1_sg U49319 ( .A(n40506), .B(n57178), .X(n34165) );
  nand_x1_sg U49320 ( .A(n34166), .B(n34167), .X(n43445) );
  nand_x1_sg U49321 ( .A(n40474), .B(n57178), .X(n34167) );
  nand_x1_sg U49322 ( .A(n34168), .B(n34169), .X(n43446) );
  nand_x1_sg U49323 ( .A(n40442), .B(n57178), .X(n34169) );
  nand_x1_sg U49324 ( .A(n34132), .B(n34133), .X(n43429) );
  nand_x1_sg U49325 ( .A(n40411), .B(n57178), .X(n34133) );
  nand_x1_sg U49326 ( .A(n34152), .B(n34153), .X(n43438) );
  nand_x1_sg U49327 ( .A(n40509), .B(n57178), .X(n34153) );
  nand_x1_sg U49328 ( .A(n34170), .B(n34171), .X(n43447) );
  nand_x1_sg U49329 ( .A(n40379), .B(n57178), .X(n34171) );
  nand_x1_sg U49330 ( .A(n34142), .B(n34143), .X(n43433) );
  nand_x1_sg U49331 ( .A(n40345), .B(n57178), .X(n34143) );
  nand_x1_sg U49332 ( .A(n34158), .B(n34159), .X(n43441) );
  nand_x1_sg U49333 ( .A(n40508), .B(n57178), .X(n34159) );
  nand_x1_sg U49334 ( .A(n34138), .B(n34139), .X(n43431) );
  nand_x1_sg U49335 ( .A(n40507), .B(n57178), .X(n34139) );
  nand_x1_sg U49336 ( .A(n34172), .B(n34173), .X(n43448) );
  nand_x1_sg U49337 ( .A(n40311), .B(n57178), .X(n34173) );
  nand_x1_sg U49338 ( .A(n34148), .B(n34149), .X(n43436) );
  nand_x1_sg U49339 ( .A(n40277), .B(n57178), .X(n34149) );
  nand_x1_sg U49340 ( .A(n33103), .B(n33104), .X(n42952) );
  nand_x1_sg U49341 ( .A(n40530), .B(n57268), .X(n33104) );
  nand_x1_sg U49342 ( .A(n33111), .B(n33112), .X(n42956) );
  nand_x1_sg U49343 ( .A(n40529), .B(n57268), .X(n33112) );
  nand_x1_sg U49344 ( .A(n33095), .B(n33096), .X(n42949) );
  nand_x1_sg U49345 ( .A(n40528), .B(n57268), .X(n33096) );
  nand_x1_sg U49346 ( .A(n33115), .B(n33116), .X(n42958) );
  nand_x1_sg U49347 ( .A(n40527), .B(n57268), .X(n33116) );
  nand_x1_sg U49348 ( .A(n33117), .B(n33118), .X(n42959) );
  nand_x1_sg U49349 ( .A(n40526), .B(n57268), .X(n33118) );
  nand_x1_sg U49350 ( .A(n33109), .B(n33110), .X(n42955) );
  nand_x1_sg U49351 ( .A(n40525), .B(n57268), .X(n33110) );
  nand_x1_sg U49352 ( .A(n33107), .B(n33108), .X(n42954) );
  nand_x1_sg U49353 ( .A(n40524), .B(n57268), .X(n33108) );
  nand_x1_sg U49354 ( .A(n33101), .B(n33102), .X(n42951) );
  nand_x1_sg U49355 ( .A(n40523), .B(n57268), .X(n33102) );
  nand_x1_sg U49356 ( .A(n33119), .B(n33120), .X(n42960) );
  nand_x1_sg U49357 ( .A(n40522), .B(n57268), .X(n33120) );
  nand_x1_sg U49358 ( .A(n33121), .B(n33122), .X(n42961) );
  nand_x1_sg U49359 ( .A(n40505), .B(n57268), .X(n33122) );
  nand_x1_sg U49360 ( .A(n33123), .B(n33124), .X(n42962) );
  nand_x1_sg U49361 ( .A(n40473), .B(n57268), .X(n33124) );
  nand_x1_sg U49362 ( .A(n33125), .B(n33126), .X(n42963) );
  nand_x1_sg U49363 ( .A(n40441), .B(n57268), .X(n33126) );
  nand_x1_sg U49364 ( .A(n33127), .B(n33128), .X(n42964) );
  nand_x1_sg U49365 ( .A(n40410), .B(n57268), .X(n33128) );
  nand_x1_sg U49366 ( .A(n33099), .B(n33100), .X(n42950) );
  nand_x1_sg U49367 ( .A(n40521), .B(n57268), .X(n33100) );
  nand_x1_sg U49368 ( .A(n33129), .B(n33130), .X(n42965) );
  nand_x1_sg U49369 ( .A(n40378), .B(n57268), .X(n33130) );
  nand_x1_sg U49370 ( .A(n33131), .B(n33132), .X(n42966) );
  nand_x1_sg U49371 ( .A(n40344), .B(n33097), .X(n33132) );
  nand_x1_sg U49372 ( .A(n33113), .B(n33114), .X(n42957) );
  nand_x1_sg U49373 ( .A(n40520), .B(n57268), .X(n33114) );
  nand_x1_sg U49374 ( .A(n33105), .B(n33106), .X(n42953) );
  nand_x1_sg U49375 ( .A(n40519), .B(n57268), .X(n33106) );
  nand_x1_sg U49376 ( .A(n33133), .B(n33134), .X(n42967) );
  nand_x1_sg U49377 ( .A(n40310), .B(n57268), .X(n33134) );
  nand_x1_sg U49378 ( .A(n33135), .B(n33136), .X(n42968) );
  nand_x1_sg U49379 ( .A(n40276), .B(n57268), .X(n33136) );
  nand_x1_sg U49380 ( .A(n32943), .B(n32944), .X(n42878) );
  nand_x1_sg U49381 ( .A(n40542), .B(n57284), .X(n32944) );
  nand_x1_sg U49382 ( .A(n32939), .B(n32940), .X(n42876) );
  nand_x1_sg U49383 ( .A(n40541), .B(n57284), .X(n32940) );
  nand_x1_sg U49384 ( .A(n32931), .B(n32932), .X(n42872) );
  nand_x1_sg U49385 ( .A(n40540), .B(n57284), .X(n32932) );
  nand_x1_sg U49386 ( .A(n32927), .B(n32928), .X(n42870) );
  nand_x1_sg U49387 ( .A(n40539), .B(n57284), .X(n32928) );
  nand_x1_sg U49388 ( .A(n32945), .B(n32946), .X(n42879) );
  nand_x1_sg U49389 ( .A(n40538), .B(n57284), .X(n32946) );
  nand_x1_sg U49390 ( .A(n32937), .B(n32938), .X(n42875) );
  nand_x1_sg U49391 ( .A(n40537), .B(n57284), .X(n32938) );
  nand_x1_sg U49392 ( .A(n32929), .B(n32930), .X(n42871) );
  nand_x1_sg U49393 ( .A(n40536), .B(n57284), .X(n32930) );
  nand_x1_sg U49394 ( .A(n32947), .B(n32948), .X(n42880) );
  nand_x1_sg U49395 ( .A(n40535), .B(n57284), .X(n32948) );
  nand_x1_sg U49396 ( .A(n32923), .B(n32924), .X(n42869) );
  nand_x1_sg U49397 ( .A(n40534), .B(n57284), .X(n32924) );
  nand_x1_sg U49398 ( .A(n32949), .B(n32950), .X(n42881) );
  nand_x1_sg U49399 ( .A(n40504), .B(n57284), .X(n32950) );
  nand_x1_sg U49400 ( .A(n32951), .B(n32952), .X(n42882) );
  nand_x1_sg U49401 ( .A(n40472), .B(n57284), .X(n32952) );
  nand_x1_sg U49402 ( .A(n32953), .B(n32954), .X(n42883) );
  nand_x1_sg U49403 ( .A(n40440), .B(n57284), .X(n32954) );
  nand_x1_sg U49404 ( .A(n32955), .B(n32956), .X(n42884) );
  nand_x1_sg U49405 ( .A(n40409), .B(n57284), .X(n32956) );
  nand_x1_sg U49406 ( .A(n32957), .B(n32958), .X(n42885) );
  nand_x1_sg U49407 ( .A(n40377), .B(n57284), .X(n32958) );
  nand_x1_sg U49408 ( .A(n32933), .B(n32934), .X(n42873) );
  nand_x1_sg U49409 ( .A(n40533), .B(n57284), .X(n32934) );
  nand_x1_sg U49410 ( .A(n32959), .B(n32960), .X(n42886) );
  nand_x1_sg U49411 ( .A(n40343), .B(n32925), .X(n32960) );
  nand_x1_sg U49412 ( .A(n32941), .B(n32942), .X(n42877) );
  nand_x1_sg U49413 ( .A(n40532), .B(n57284), .X(n32942) );
  nand_x1_sg U49414 ( .A(n32961), .B(n32962), .X(n42887) );
  nand_x1_sg U49415 ( .A(n40309), .B(n57284), .X(n32962) );
  nand_x1_sg U49416 ( .A(n32935), .B(n32936), .X(n42874) );
  nand_x1_sg U49417 ( .A(n40531), .B(n57284), .X(n32936) );
  nand_x1_sg U49418 ( .A(n32963), .B(n32964), .X(n42888) );
  nand_x1_sg U49419 ( .A(n40275), .B(n57284), .X(n32964) );
  nand_x1_sg U49420 ( .A(n33662), .B(n33663), .X(n43212) );
  nand_x1_sg U49421 ( .A(n40554), .B(n57219), .X(n33663) );
  nand_x1_sg U49422 ( .A(n33670), .B(n33671), .X(n43216) );
  nand_x1_sg U49423 ( .A(n40553), .B(n57219), .X(n33671) );
  nand_x1_sg U49424 ( .A(n33654), .B(n33655), .X(n43209) );
  nand_x1_sg U49425 ( .A(n40552), .B(n57219), .X(n33655) );
  nand_x1_sg U49426 ( .A(n33674), .B(n33675), .X(n43218) );
  nand_x1_sg U49427 ( .A(n40551), .B(n57219), .X(n33675) );
  nand_x1_sg U49428 ( .A(n33676), .B(n33677), .X(n43219) );
  nand_x1_sg U49429 ( .A(n40550), .B(n57219), .X(n33677) );
  nand_x1_sg U49430 ( .A(n33668), .B(n33669), .X(n43215) );
  nand_x1_sg U49431 ( .A(n40549), .B(n57219), .X(n33669) );
  nand_x1_sg U49432 ( .A(n33666), .B(n33667), .X(n43214) );
  nand_x1_sg U49433 ( .A(n40548), .B(n57219), .X(n33667) );
  nand_x1_sg U49434 ( .A(n33660), .B(n33661), .X(n43211) );
  nand_x1_sg U49435 ( .A(n40547), .B(n57219), .X(n33661) );
  nand_x1_sg U49436 ( .A(n33678), .B(n33679), .X(n43220) );
  nand_x1_sg U49437 ( .A(n40546), .B(n57219), .X(n33679) );
  nand_x1_sg U49438 ( .A(n33680), .B(n33681), .X(n43221) );
  nand_x1_sg U49439 ( .A(n40503), .B(n57219), .X(n33681) );
  nand_x1_sg U49440 ( .A(n33682), .B(n33683), .X(n43222) );
  nand_x1_sg U49441 ( .A(n40471), .B(n57219), .X(n33683) );
  nand_x1_sg U49442 ( .A(n33684), .B(n33685), .X(n43223) );
  nand_x1_sg U49443 ( .A(n40439), .B(n57219), .X(n33685) );
  nand_x1_sg U49444 ( .A(n33686), .B(n33687), .X(n43224) );
  nand_x1_sg U49445 ( .A(n40408), .B(n57219), .X(n33687) );
  nand_x1_sg U49446 ( .A(n33658), .B(n33659), .X(n43210) );
  nand_x1_sg U49447 ( .A(n40545), .B(n57219), .X(n33659) );
  nand_x1_sg U49448 ( .A(n33688), .B(n33689), .X(n43225) );
  nand_x1_sg U49449 ( .A(n40376), .B(n57219), .X(n33689) );
  nand_x1_sg U49450 ( .A(n33690), .B(n33691), .X(n43226) );
  nand_x1_sg U49451 ( .A(n40342), .B(n33656), .X(n33691) );
  nand_x1_sg U49452 ( .A(n33672), .B(n33673), .X(n43217) );
  nand_x1_sg U49453 ( .A(n40544), .B(n57219), .X(n33673) );
  nand_x1_sg U49454 ( .A(n33664), .B(n33665), .X(n43213) );
  nand_x1_sg U49455 ( .A(n40543), .B(n57219), .X(n33665) );
  nand_x1_sg U49456 ( .A(n33692), .B(n33693), .X(n43227) );
  nand_x1_sg U49457 ( .A(n40308), .B(n57219), .X(n33693) );
  nand_x1_sg U49458 ( .A(n33694), .B(n33695), .X(n43228) );
  nand_x1_sg U49459 ( .A(n40248), .B(n57219), .X(n33695) );
  nand_x1_sg U49460 ( .A(n33704), .B(n33705), .X(n43232) );
  nand_x1_sg U49461 ( .A(n40566), .B(n57215), .X(n33705) );
  nand_x1_sg U49462 ( .A(n33712), .B(n33713), .X(n43236) );
  nand_x1_sg U49463 ( .A(n40565), .B(n57215), .X(n33713) );
  nand_x1_sg U49464 ( .A(n33696), .B(n33697), .X(n43229) );
  nand_x1_sg U49465 ( .A(n40564), .B(n57215), .X(n33697) );
  nand_x1_sg U49466 ( .A(n33716), .B(n33717), .X(n43238) );
  nand_x1_sg U49467 ( .A(n40563), .B(n57215), .X(n33717) );
  nand_x1_sg U49468 ( .A(n33718), .B(n33719), .X(n43239) );
  nand_x1_sg U49469 ( .A(n40562), .B(n57215), .X(n33719) );
  nand_x1_sg U49470 ( .A(n33710), .B(n33711), .X(n43235) );
  nand_x1_sg U49471 ( .A(n40561), .B(n57215), .X(n33711) );
  nand_x1_sg U49472 ( .A(n33708), .B(n33709), .X(n43234) );
  nand_x1_sg U49473 ( .A(n40560), .B(n57215), .X(n33709) );
  nand_x1_sg U49474 ( .A(n33702), .B(n33703), .X(n43231) );
  nand_x1_sg U49475 ( .A(n40559), .B(n57215), .X(n33703) );
  nand_x1_sg U49476 ( .A(n33720), .B(n33721), .X(n43240) );
  nand_x1_sg U49477 ( .A(n40558), .B(n57215), .X(n33721) );
  nand_x1_sg U49478 ( .A(n33722), .B(n33723), .X(n43241) );
  nand_x1_sg U49479 ( .A(n40502), .B(n57215), .X(n33723) );
  nand_x1_sg U49480 ( .A(n33724), .B(n33725), .X(n43242) );
  nand_x1_sg U49481 ( .A(n40470), .B(n57215), .X(n33725) );
  nand_x1_sg U49482 ( .A(n33726), .B(n33727), .X(n43243) );
  nand_x1_sg U49483 ( .A(n40438), .B(n57215), .X(n33727) );
  nand_x1_sg U49484 ( .A(n33728), .B(n33729), .X(n43244) );
  nand_x1_sg U49485 ( .A(n40407), .B(n57215), .X(n33729) );
  nand_x1_sg U49486 ( .A(n33700), .B(n33701), .X(n43230) );
  nand_x1_sg U49487 ( .A(n40557), .B(n57215), .X(n33701) );
  nand_x1_sg U49488 ( .A(n33730), .B(n33731), .X(n43245) );
  nand_x1_sg U49489 ( .A(n40375), .B(n57215), .X(n33731) );
  nand_x1_sg U49490 ( .A(n33732), .B(n33733), .X(n43246) );
  nand_x1_sg U49491 ( .A(n40341), .B(n33698), .X(n33733) );
  nand_x1_sg U49492 ( .A(n33714), .B(n33715), .X(n43237) );
  nand_x1_sg U49493 ( .A(n40556), .B(n57215), .X(n33715) );
  nand_x1_sg U49494 ( .A(n33706), .B(n33707), .X(n43233) );
  nand_x1_sg U49495 ( .A(n40555), .B(n57215), .X(n33707) );
  nand_x1_sg U49496 ( .A(n33734), .B(n33735), .X(n43247) );
  nand_x1_sg U49497 ( .A(n40307), .B(n57215), .X(n33735) );
  nand_x1_sg U49498 ( .A(n33736), .B(n33737), .X(n43248) );
  nand_x1_sg U49499 ( .A(n40274), .B(n57215), .X(n33737) );
  nand_x1_sg U49500 ( .A(n33575), .B(n33576), .X(n43172) );
  nand_x1_sg U49501 ( .A(n40578), .B(n57226), .X(n33576) );
  nand_x1_sg U49502 ( .A(n33583), .B(n33584), .X(n43176) );
  nand_x1_sg U49503 ( .A(n40577), .B(n33569), .X(n33584) );
  nand_x1_sg U49504 ( .A(n33577), .B(n33578), .X(n43173) );
  nand_x1_sg U49505 ( .A(n40576), .B(n57226), .X(n33578) );
  nand_x1_sg U49506 ( .A(n33587), .B(n33588), .X(n43178) );
  nand_x1_sg U49507 ( .A(n40575), .B(n57226), .X(n33588) );
  nand_x1_sg U49508 ( .A(n33589), .B(n33590), .X(n43179) );
  nand_x1_sg U49509 ( .A(n40574), .B(n57226), .X(n33590) );
  nand_x1_sg U49510 ( .A(n33581), .B(n33582), .X(n43175) );
  nand_x1_sg U49511 ( .A(n40573), .B(n57226), .X(n33582) );
  nand_x1_sg U49512 ( .A(n33567), .B(n33568), .X(n43169) );
  nand_x1_sg U49513 ( .A(n40572), .B(n57226), .X(n33568) );
  nand_x1_sg U49514 ( .A(n33571), .B(n33572), .X(n43170) );
  nand_x1_sg U49515 ( .A(n40571), .B(n57226), .X(n33572) );
  nand_x1_sg U49516 ( .A(n33591), .B(n33592), .X(n43180) );
  nand_x1_sg U49517 ( .A(n40570), .B(n57226), .X(n33592) );
  nand_x1_sg U49518 ( .A(n33593), .B(n33594), .X(n43181) );
  nand_x1_sg U49519 ( .A(n40501), .B(n57226), .X(n33594) );
  nand_x1_sg U49520 ( .A(n33595), .B(n33596), .X(n43182) );
  nand_x1_sg U49521 ( .A(n40469), .B(n57226), .X(n33596) );
  nand_x1_sg U49522 ( .A(n33573), .B(n33574), .X(n43171) );
  nand_x1_sg U49523 ( .A(n40569), .B(n57226), .X(n33574) );
  nand_x1_sg U49524 ( .A(n33597), .B(n33598), .X(n43183) );
  nand_x1_sg U49525 ( .A(n40437), .B(n57226), .X(n33598) );
  nand_x1_sg U49526 ( .A(n33579), .B(n33580), .X(n43174) );
  nand_x1_sg U49527 ( .A(n40568), .B(n57226), .X(n33580) );
  nand_x1_sg U49528 ( .A(n33599), .B(n33600), .X(n43184) );
  nand_x1_sg U49529 ( .A(n40406), .B(n57226), .X(n33600) );
  nand_x1_sg U49530 ( .A(n33601), .B(n33602), .X(n43185) );
  nand_x1_sg U49531 ( .A(n40374), .B(n57226), .X(n33602) );
  nand_x1_sg U49532 ( .A(n33585), .B(n33586), .X(n43177) );
  nand_x1_sg U49533 ( .A(n40567), .B(n57226), .X(n33586) );
  nand_x1_sg U49534 ( .A(n33603), .B(n33604), .X(n43186) );
  nand_x1_sg U49535 ( .A(n40340), .B(n57226), .X(n33604) );
  nand_x1_sg U49536 ( .A(n33605), .B(n33606), .X(n43187) );
  nand_x1_sg U49537 ( .A(n40306), .B(n57226), .X(n33606) );
  nand_x1_sg U49538 ( .A(n33607), .B(n33608), .X(n43188) );
  nand_x1_sg U49539 ( .A(n40273), .B(n57226), .X(n33608) );
  nand_x1_sg U49540 ( .A(n33630), .B(n33631), .X(n43198) );
  nand_x1_sg U49541 ( .A(n40589), .B(n57223), .X(n33631) );
  nand_x1_sg U49542 ( .A(n33626), .B(n33627), .X(n43196) );
  nand_x1_sg U49543 ( .A(n40588), .B(n57223), .X(n33627) );
  nand_x1_sg U49544 ( .A(n33632), .B(n33633), .X(n43199) );
  nand_x1_sg U49545 ( .A(n40587), .B(n57223), .X(n33633) );
  nand_x1_sg U49546 ( .A(n33634), .B(n33635), .X(n43200) );
  nand_x1_sg U49547 ( .A(n40500), .B(n57223), .X(n33635) );
  nand_x1_sg U49548 ( .A(n33618), .B(n33619), .X(n43192) );
  nand_x1_sg U49549 ( .A(n40586), .B(n57223), .X(n33619) );
  nand_x1_sg U49550 ( .A(n33624), .B(n33625), .X(n43195) );
  nand_x1_sg U49551 ( .A(n40585), .B(n57223), .X(n33625) );
  nand_x1_sg U49552 ( .A(n33636), .B(n33637), .X(n43201) );
  nand_x1_sg U49553 ( .A(n40468), .B(n57223), .X(n33637) );
  nand_x1_sg U49554 ( .A(n33638), .B(n33639), .X(n43202) );
  nand_x1_sg U49555 ( .A(n40436), .B(n57223), .X(n33639) );
  nand_x1_sg U49556 ( .A(n33614), .B(n33615), .X(n43190) );
  nand_x1_sg U49557 ( .A(n40584), .B(n57223), .X(n33615) );
  nand_x1_sg U49558 ( .A(n33640), .B(n33641), .X(n43203) );
  nand_x1_sg U49559 ( .A(n40405), .B(n57223), .X(n33641) );
  nand_x1_sg U49560 ( .A(n33622), .B(n33623), .X(n43194) );
  nand_x1_sg U49561 ( .A(n40583), .B(n57223), .X(n33623) );
  nand_x1_sg U49562 ( .A(n33642), .B(n33643), .X(n43204) );
  nand_x1_sg U49563 ( .A(n40373), .B(n57223), .X(n33643) );
  nand_x1_sg U49564 ( .A(n33616), .B(n33617), .X(n43191) );
  nand_x1_sg U49565 ( .A(n40582), .B(n57223), .X(n33617) );
  nand_x1_sg U49566 ( .A(n33644), .B(n33645), .X(n43205) );
  nand_x1_sg U49567 ( .A(n40339), .B(n57223), .X(n33645) );
  nand_x1_sg U49568 ( .A(n33620), .B(n33621), .X(n43193) );
  nand_x1_sg U49569 ( .A(n40581), .B(n57223), .X(n33621) );
  nand_x1_sg U49570 ( .A(n33646), .B(n33647), .X(n43206) );
  nand_x1_sg U49571 ( .A(n40305), .B(n33612), .X(n33647) );
  nand_x1_sg U49572 ( .A(n33628), .B(n33629), .X(n43197) );
  nand_x1_sg U49573 ( .A(n40580), .B(n57223), .X(n33629) );
  nand_x1_sg U49574 ( .A(n33648), .B(n33649), .X(n43207) );
  nand_x1_sg U49575 ( .A(n40272), .B(n57223), .X(n33649) );
  nand_x1_sg U49576 ( .A(n33610), .B(n33611), .X(n43189) );
  nand_x1_sg U49577 ( .A(n40579), .B(n57223), .X(n33611) );
  nand_x1_sg U49578 ( .A(n33650), .B(n33651), .X(n43208) );
  nand_x1_sg U49579 ( .A(n40247), .B(n57223), .X(n33651) );
  nand_x1_sg U49580 ( .A(n32878), .B(n32879), .X(n42849) );
  nand_x1_sg U49581 ( .A(n40592), .B(n57288), .X(n32879) );
  nand_x1_sg U49582 ( .A(n32882), .B(n32883), .X(n42850) );
  nand_x1_sg U49583 ( .A(n40591), .B(n57288), .X(n32883) );
  nand_x1_sg U49584 ( .A(n32884), .B(n32885), .X(n42851) );
  nand_x1_sg U49585 ( .A(n40590), .B(n57288), .X(n32885) );
  nand_x1_sg U49586 ( .A(n32886), .B(n32887), .X(n42852) );
  nand_x1_sg U49587 ( .A(n40499), .B(n57288), .X(n32887) );
  nand_x1_sg U49588 ( .A(n32890), .B(n32891), .X(n42854) );
  nand_x1_sg U49589 ( .A(n40404), .B(n57288), .X(n32891) );
  nand_x1_sg U49590 ( .A(n32888), .B(n32889), .X(n42853) );
  nand_x1_sg U49591 ( .A(n40467), .B(n57288), .X(n32889) );
  nand_x1_sg U49592 ( .A(n32892), .B(n32893), .X(n42855) );
  nand_x1_sg U49593 ( .A(n40372), .B(n57288), .X(n32893) );
  nand_x1_sg U49594 ( .A(n32906), .B(n32907), .X(n42862) );
  nand_x1_sg U49595 ( .A(n40403), .B(n57288), .X(n32907) );
  nand_x1_sg U49596 ( .A(n32894), .B(n32895), .X(n42856) );
  nand_x1_sg U49597 ( .A(n40338), .B(n57288), .X(n32895) );
  nand_x1_sg U49598 ( .A(n32908), .B(n32909), .X(n42863) );
  nand_x1_sg U49599 ( .A(n40371), .B(n57288), .X(n32909) );
  nand_x1_sg U49600 ( .A(n32896), .B(n32897), .X(n42857) );
  nand_x1_sg U49601 ( .A(n40304), .B(n57288), .X(n32897) );
  nand_x1_sg U49602 ( .A(n32910), .B(n32911), .X(n42864) );
  nand_x1_sg U49603 ( .A(n40337), .B(n57288), .X(n32911) );
  nand_x1_sg U49604 ( .A(n32898), .B(n32899), .X(n42858) );
  nand_x1_sg U49605 ( .A(n40271), .B(n57288), .X(n32899) );
  nand_x1_sg U49606 ( .A(n32912), .B(n32913), .X(n42865) );
  nand_x1_sg U49607 ( .A(n40303), .B(n57288), .X(n32913) );
  nand_x1_sg U49608 ( .A(n32900), .B(n32901), .X(n42859) );
  nand_x1_sg U49609 ( .A(n40246), .B(n57288), .X(n32901) );
  nand_x1_sg U49610 ( .A(n32914), .B(n32915), .X(n42866) );
  nand_x1_sg U49611 ( .A(n40270), .B(n32880), .X(n32915) );
  nand_x1_sg U49612 ( .A(n32902), .B(n32903), .X(n42860) );
  nand_x1_sg U49613 ( .A(n40233), .B(n57288), .X(n32903) );
  nand_x1_sg U49614 ( .A(n32916), .B(n32917), .X(n42867) );
  nand_x1_sg U49615 ( .A(n40245), .B(n57288), .X(n32917) );
  nand_x1_sg U49616 ( .A(n32904), .B(n32905), .X(n42861) );
  nand_x1_sg U49617 ( .A(n40231), .B(n57288), .X(n32905) );
  nand_x1_sg U49618 ( .A(n32918), .B(n32919), .X(n42868) );
  nand_x1_sg U49619 ( .A(n40230), .B(n57288), .X(n32919) );
  nand_x1_sg U49620 ( .A(n33145), .B(n33146), .X(n42972) );
  nand_x1_sg U49621 ( .A(n40603), .B(n57264), .X(n33146) );
  nand_x1_sg U49622 ( .A(n33153), .B(n33154), .X(n42976) );
  nand_x1_sg U49623 ( .A(n40602), .B(n57264), .X(n33154) );
  nand_x1_sg U49624 ( .A(n33137), .B(n33138), .X(n42969) );
  nand_x1_sg U49625 ( .A(n40601), .B(n57264), .X(n33138) );
  nand_x1_sg U49626 ( .A(n33157), .B(n33158), .X(n42978) );
  nand_x1_sg U49627 ( .A(n40600), .B(n57264), .X(n33158) );
  nand_x1_sg U49628 ( .A(n33159), .B(n33160), .X(n42979) );
  nand_x1_sg U49629 ( .A(n40599), .B(n57264), .X(n33160) );
  nand_x1_sg U49630 ( .A(n33151), .B(n33152), .X(n42975) );
  nand_x1_sg U49631 ( .A(n40598), .B(n57264), .X(n33152) );
  nand_x1_sg U49632 ( .A(n33149), .B(n33150), .X(n42974) );
  nand_x1_sg U49633 ( .A(n40597), .B(n57264), .X(n33150) );
  nand_x1_sg U49634 ( .A(n33143), .B(n33144), .X(n42971) );
  nand_x1_sg U49635 ( .A(n40596), .B(n57264), .X(n33144) );
  nand_x1_sg U49636 ( .A(n33161), .B(n33162), .X(n42980) );
  nand_x1_sg U49637 ( .A(n40498), .B(n57264), .X(n33162) );
  nand_x1_sg U49638 ( .A(n33163), .B(n33164), .X(n42981) );
  nand_x1_sg U49639 ( .A(n40466), .B(n57264), .X(n33164) );
  nand_x1_sg U49640 ( .A(n33165), .B(n33166), .X(n42982) );
  nand_x1_sg U49641 ( .A(n40435), .B(n57264), .X(n33166) );
  nand_x1_sg U49642 ( .A(n33167), .B(n33168), .X(n42983) );
  nand_x1_sg U49643 ( .A(n40402), .B(n57264), .X(n33168) );
  nand_x1_sg U49644 ( .A(n33169), .B(n33170), .X(n42984) );
  nand_x1_sg U49645 ( .A(n40370), .B(n57264), .X(n33170) );
  nand_x1_sg U49646 ( .A(n33141), .B(n33142), .X(n42970) );
  nand_x1_sg U49647 ( .A(n40595), .B(n57264), .X(n33142) );
  nand_x1_sg U49648 ( .A(n33171), .B(n33172), .X(n42985) );
  nand_x1_sg U49649 ( .A(n40336), .B(n57264), .X(n33172) );
  nand_x1_sg U49650 ( .A(n33173), .B(n33174), .X(n42986) );
  nand_x1_sg U49651 ( .A(n40302), .B(n33139), .X(n33174) );
  nand_x1_sg U49652 ( .A(n33155), .B(n33156), .X(n42977) );
  nand_x1_sg U49653 ( .A(n40594), .B(n57264), .X(n33156) );
  nand_x1_sg U49654 ( .A(n33147), .B(n33148), .X(n42973) );
  nand_x1_sg U49655 ( .A(n40593), .B(n57264), .X(n33148) );
  nand_x1_sg U49656 ( .A(n33175), .B(n33176), .X(n42987) );
  nand_x1_sg U49657 ( .A(n40269), .B(n57264), .X(n33176) );
  nand_x1_sg U49658 ( .A(n33177), .B(n33178), .X(n42988) );
  nand_x1_sg U49659 ( .A(n40244), .B(n57264), .X(n33178) );
  nand_x1_sg U49660 ( .A(n33188), .B(n33189), .X(n42992) );
  nand_x1_sg U49661 ( .A(n40614), .B(n57260), .X(n33189) );
  nand_x1_sg U49662 ( .A(n33196), .B(n33197), .X(n42996) );
  nand_x1_sg U49663 ( .A(n40613), .B(n57260), .X(n33197) );
  nand_x1_sg U49664 ( .A(n33190), .B(n33191), .X(n42993) );
  nand_x1_sg U49665 ( .A(n40612), .B(n57260), .X(n33191) );
  nand_x1_sg U49666 ( .A(n33200), .B(n33201), .X(n42998) );
  nand_x1_sg U49667 ( .A(n40611), .B(n57260), .X(n33201) );
  nand_x1_sg U49668 ( .A(n33202), .B(n33203), .X(n42999) );
  nand_x1_sg U49669 ( .A(n40610), .B(n57260), .X(n33203) );
  nand_x1_sg U49670 ( .A(n33194), .B(n33195), .X(n42995) );
  nand_x1_sg U49671 ( .A(n40609), .B(n57260), .X(n33195) );
  nand_x1_sg U49672 ( .A(n33180), .B(n33181), .X(n42989) );
  nand_x1_sg U49673 ( .A(n40608), .B(n57260), .X(n33181) );
  nand_x1_sg U49674 ( .A(n33184), .B(n33185), .X(n42990) );
  nand_x1_sg U49675 ( .A(n40607), .B(n57260), .X(n33185) );
  nand_x1_sg U49676 ( .A(n33204), .B(n33205), .X(n43000) );
  nand_x1_sg U49677 ( .A(n40497), .B(n57260), .X(n33205) );
  nand_x1_sg U49678 ( .A(n33206), .B(n33207), .X(n43001) );
  nand_x1_sg U49679 ( .A(n40465), .B(n57260), .X(n33207) );
  nand_x1_sg U49680 ( .A(n33208), .B(n33209), .X(n43002) );
  nand_x1_sg U49681 ( .A(n40434), .B(n57260), .X(n33209) );
  nand_x1_sg U49682 ( .A(n33186), .B(n33187), .X(n42991) );
  nand_x1_sg U49683 ( .A(n40606), .B(n57260), .X(n33187) );
  nand_x1_sg U49684 ( .A(n33210), .B(n33211), .X(n43003) );
  nand_x1_sg U49685 ( .A(n40401), .B(n57260), .X(n33211) );
  nand_x1_sg U49686 ( .A(n33192), .B(n33193), .X(n42994) );
  nand_x1_sg U49687 ( .A(n40605), .B(n57260), .X(n33193) );
  nand_x1_sg U49688 ( .A(n33212), .B(n33213), .X(n43004) );
  nand_x1_sg U49689 ( .A(n40369), .B(n57260), .X(n33213) );
  nand_x1_sg U49690 ( .A(n33214), .B(n33215), .X(n43005) );
  nand_x1_sg U49691 ( .A(n40335), .B(n57260), .X(n33215) );
  nand_x1_sg U49692 ( .A(n33198), .B(n33199), .X(n42997) );
  nand_x1_sg U49693 ( .A(n40604), .B(n33182), .X(n33199) );
  nand_x1_sg U49694 ( .A(n33216), .B(n33217), .X(n43006) );
  nand_x1_sg U49695 ( .A(n40301), .B(n57260), .X(n33217) );
  nand_x1_sg U49696 ( .A(n33218), .B(n33219), .X(n43007) );
  nand_x1_sg U49697 ( .A(n40268), .B(n57260), .X(n33219) );
  nand_x1_sg U49698 ( .A(n33220), .B(n33221), .X(n43008) );
  nand_x1_sg U49699 ( .A(n40243), .B(n57260), .X(n33221) );
  nand_x1_sg U49700 ( .A(n33231), .B(n33232), .X(n43012) );
  nand_x1_sg U49701 ( .A(n40625), .B(n57256), .X(n33232) );
  nand_x1_sg U49702 ( .A(n33239), .B(n33240), .X(n43016) );
  nand_x1_sg U49703 ( .A(n40624), .B(n57256), .X(n33240) );
  nand_x1_sg U49704 ( .A(n33223), .B(n33224), .X(n43009) );
  nand_x1_sg U49705 ( .A(n40623), .B(n57256), .X(n33224) );
  nand_x1_sg U49706 ( .A(n33243), .B(n33244), .X(n43018) );
  nand_x1_sg U49707 ( .A(n40622), .B(n57256), .X(n33244) );
  nand_x1_sg U49708 ( .A(n33245), .B(n33246), .X(n43019) );
  nand_x1_sg U49709 ( .A(n40621), .B(n57256), .X(n33246) );
  nand_x1_sg U49710 ( .A(n33237), .B(n33238), .X(n43015) );
  nand_x1_sg U49711 ( .A(n40620), .B(n57256), .X(n33238) );
  nand_x1_sg U49712 ( .A(n33235), .B(n33236), .X(n43014) );
  nand_x1_sg U49713 ( .A(n40619), .B(n57256), .X(n33236) );
  nand_x1_sg U49714 ( .A(n33229), .B(n33230), .X(n43011) );
  nand_x1_sg U49715 ( .A(n40618), .B(n57256), .X(n33230) );
  nand_x1_sg U49716 ( .A(n33247), .B(n33248), .X(n43020) );
  nand_x1_sg U49717 ( .A(n40496), .B(n57256), .X(n33248) );
  nand_x1_sg U49718 ( .A(n33249), .B(n33250), .X(n43021) );
  nand_x1_sg U49719 ( .A(n40464), .B(n57256), .X(n33250) );
  nand_x1_sg U49720 ( .A(n33251), .B(n33252), .X(n43022) );
  nand_x1_sg U49721 ( .A(n40433), .B(n57256), .X(n33252) );
  nand_x1_sg U49722 ( .A(n33253), .B(n33254), .X(n43023) );
  nand_x1_sg U49723 ( .A(n40400), .B(n57256), .X(n33254) );
  nand_x1_sg U49724 ( .A(n33255), .B(n33256), .X(n43024) );
  nand_x1_sg U49725 ( .A(n40368), .B(n57256), .X(n33256) );
  nand_x1_sg U49726 ( .A(n33227), .B(n33228), .X(n43010) );
  nand_x1_sg U49727 ( .A(n40617), .B(n57256), .X(n33228) );
  nand_x1_sg U49728 ( .A(n33257), .B(n33258), .X(n43025) );
  nand_x1_sg U49729 ( .A(n40334), .B(n57256), .X(n33258) );
  nand_x1_sg U49730 ( .A(n33259), .B(n33260), .X(n43026) );
  nand_x1_sg U49731 ( .A(n40300), .B(n33225), .X(n33260) );
  nand_x1_sg U49732 ( .A(n33241), .B(n33242), .X(n43017) );
  nand_x1_sg U49733 ( .A(n40616), .B(n57256), .X(n33242) );
  nand_x1_sg U49734 ( .A(n33233), .B(n33234), .X(n43013) );
  nand_x1_sg U49735 ( .A(n40615), .B(n57256), .X(n33234) );
  nand_x1_sg U49736 ( .A(n33261), .B(n33262), .X(n43027) );
  nand_x1_sg U49737 ( .A(n40267), .B(n57256), .X(n33262) );
  nand_x1_sg U49738 ( .A(n33263), .B(n33264), .X(n43028) );
  nand_x1_sg U49739 ( .A(n40242), .B(n57256), .X(n33264) );
  nand_x1_sg U49740 ( .A(n32994), .B(n32995), .X(n42902) );
  nand_x1_sg U49741 ( .A(n40637), .B(n57280), .X(n32995) );
  nand_x1_sg U49742 ( .A(n32984), .B(n32985), .X(n42897) );
  nand_x1_sg U49743 ( .A(n40636), .B(n32968), .X(n32985) );
  nand_x1_sg U49744 ( .A(n32974), .B(n32975), .X(n42892) );
  nand_x1_sg U49745 ( .A(n40635), .B(n57280), .X(n32975) );
  nand_x1_sg U49746 ( .A(n32992), .B(n32993), .X(n42901) );
  nand_x1_sg U49747 ( .A(n40634), .B(n57280), .X(n32993) );
  nand_x1_sg U49748 ( .A(n33004), .B(n33005), .X(n42907) );
  nand_x1_sg U49749 ( .A(n40633), .B(n57280), .X(n33005) );
  nand_x1_sg U49750 ( .A(n33002), .B(n33003), .X(n42906) );
  nand_x1_sg U49751 ( .A(n40632), .B(n57280), .X(n33003) );
  nand_x1_sg U49752 ( .A(n32970), .B(n32971), .X(n42890) );
  nand_x1_sg U49753 ( .A(n40495), .B(n57280), .X(n32971) );
  nand_x1_sg U49754 ( .A(n32998), .B(n32999), .X(n42904) );
  nand_x1_sg U49755 ( .A(n40463), .B(n57280), .X(n32999) );
  nand_x1_sg U49756 ( .A(n32978), .B(n32979), .X(n42894) );
  nand_x1_sg U49757 ( .A(n40631), .B(n57280), .X(n32979) );
  nand_x1_sg U49758 ( .A(n33000), .B(n33001), .X(n42905) );
  nand_x1_sg U49759 ( .A(n40432), .B(n57280), .X(n33001) );
  nand_x1_sg U49760 ( .A(n32966), .B(n32967), .X(n42889) );
  nand_x1_sg U49761 ( .A(n40630), .B(n57280), .X(n32967) );
  nand_x1_sg U49762 ( .A(n32982), .B(n32983), .X(n42896) );
  nand_x1_sg U49763 ( .A(n40399), .B(n57280), .X(n32983) );
  nand_x1_sg U49764 ( .A(n32976), .B(n32977), .X(n42893) );
  nand_x1_sg U49765 ( .A(n40629), .B(n57280), .X(n32977) );
  nand_x1_sg U49766 ( .A(n33006), .B(n33007), .X(n42908) );
  nand_x1_sg U49767 ( .A(n40367), .B(n57280), .X(n33007) );
  nand_x1_sg U49768 ( .A(n32988), .B(n32989), .X(n42899) );
  nand_x1_sg U49769 ( .A(n40628), .B(n57280), .X(n32989) );
  nand_x1_sg U49770 ( .A(n32996), .B(n32997), .X(n42903) );
  nand_x1_sg U49771 ( .A(n40333), .B(n57280), .X(n32997) );
  nand_x1_sg U49772 ( .A(n32980), .B(n32981), .X(n42895) );
  nand_x1_sg U49773 ( .A(n40627), .B(n57280), .X(n32981) );
  nand_x1_sg U49774 ( .A(n32972), .B(n32973), .X(n42891) );
  nand_x1_sg U49775 ( .A(n40299), .B(n57280), .X(n32973) );
  nand_x1_sg U49776 ( .A(n32990), .B(n32991), .X(n42900) );
  nand_x1_sg U49777 ( .A(n40626), .B(n57280), .X(n32991) );
  nand_x1_sg U49778 ( .A(n32986), .B(n32987), .X(n42898) );
  nand_x1_sg U49779 ( .A(n40266), .B(n57280), .X(n32987) );
  nand_x1_sg U49780 ( .A(n33747), .B(n33748), .X(n43252) );
  nand_x1_sg U49781 ( .A(n40649), .B(n57211), .X(n33748) );
  nand_x1_sg U49782 ( .A(n33755), .B(n33756), .X(n43256) );
  nand_x1_sg U49783 ( .A(n40648), .B(n57211), .X(n33756) );
  nand_x1_sg U49784 ( .A(n33739), .B(n33740), .X(n43249) );
  nand_x1_sg U49785 ( .A(n40647), .B(n57211), .X(n33740) );
  nand_x1_sg U49786 ( .A(n33759), .B(n33760), .X(n43258) );
  nand_x1_sg U49787 ( .A(n40646), .B(n57211), .X(n33760) );
  nand_x1_sg U49788 ( .A(n33761), .B(n33762), .X(n43259) );
  nand_x1_sg U49789 ( .A(n40645), .B(n57211), .X(n33762) );
  nand_x1_sg U49790 ( .A(n33753), .B(n33754), .X(n43255) );
  nand_x1_sg U49791 ( .A(n40644), .B(n57211), .X(n33754) );
  nand_x1_sg U49792 ( .A(n33751), .B(n33752), .X(n43254) );
  nand_x1_sg U49793 ( .A(n40643), .B(n57211), .X(n33752) );
  nand_x1_sg U49794 ( .A(n33745), .B(n33746), .X(n43251) );
  nand_x1_sg U49795 ( .A(n40642), .B(n57211), .X(n33746) );
  nand_x1_sg U49796 ( .A(n33763), .B(n33764), .X(n43260) );
  nand_x1_sg U49797 ( .A(n40641), .B(n57211), .X(n33764) );
  nand_x1_sg U49798 ( .A(n33765), .B(n33766), .X(n43261) );
  nand_x1_sg U49799 ( .A(n40494), .B(n57211), .X(n33766) );
  nand_x1_sg U49800 ( .A(n33767), .B(n33768), .X(n43262) );
  nand_x1_sg U49801 ( .A(n40462), .B(n57211), .X(n33768) );
  nand_x1_sg U49802 ( .A(n33769), .B(n33770), .X(n43263) );
  nand_x1_sg U49803 ( .A(n40431), .B(n57211), .X(n33770) );
  nand_x1_sg U49804 ( .A(n33771), .B(n33772), .X(n43264) );
  nand_x1_sg U49805 ( .A(n40398), .B(n57211), .X(n33772) );
  nand_x1_sg U49806 ( .A(n33743), .B(n33744), .X(n43250) );
  nand_x1_sg U49807 ( .A(n40640), .B(n57211), .X(n33744) );
  nand_x1_sg U49808 ( .A(n33773), .B(n33774), .X(n43265) );
  nand_x1_sg U49809 ( .A(n40366), .B(n57211), .X(n33774) );
  nand_x1_sg U49810 ( .A(n33775), .B(n33776), .X(n43266) );
  nand_x1_sg U49811 ( .A(n40332), .B(n33741), .X(n33776) );
  nand_x1_sg U49812 ( .A(n33757), .B(n33758), .X(n43257) );
  nand_x1_sg U49813 ( .A(n40639), .B(n57211), .X(n33758) );
  nand_x1_sg U49814 ( .A(n33749), .B(n33750), .X(n43253) );
  nand_x1_sg U49815 ( .A(n40638), .B(n57211), .X(n33750) );
  nand_x1_sg U49816 ( .A(n33777), .B(n33778), .X(n43267) );
  nand_x1_sg U49817 ( .A(n40298), .B(n57211), .X(n33778) );
  nand_x1_sg U49818 ( .A(n33779), .B(n33780), .X(n43268) );
  nand_x1_sg U49819 ( .A(n40265), .B(n57211), .X(n33780) );
  nand_x1_sg U49820 ( .A(n33792), .B(n33793), .X(n43272) );
  nand_x1_sg U49821 ( .A(n40661), .B(n57207), .X(n33793) );
  nand_x1_sg U49822 ( .A(n33800), .B(n33801), .X(n43276) );
  nand_x1_sg U49823 ( .A(n40660), .B(n33786), .X(n33801) );
  nand_x1_sg U49824 ( .A(n33784), .B(n33785), .X(n43269) );
  nand_x1_sg U49825 ( .A(n40659), .B(n57207), .X(n33785) );
  nand_x1_sg U49826 ( .A(n33804), .B(n33805), .X(n43278) );
  nand_x1_sg U49827 ( .A(n40658), .B(n57207), .X(n33805) );
  nand_x1_sg U49828 ( .A(n33806), .B(n33807), .X(n43279) );
  nand_x1_sg U49829 ( .A(n40657), .B(n57207), .X(n33807) );
  nand_x1_sg U49830 ( .A(n33798), .B(n33799), .X(n43275) );
  nand_x1_sg U49831 ( .A(n40656), .B(n57207), .X(n33799) );
  nand_x1_sg U49832 ( .A(n33796), .B(n33797), .X(n43274) );
  nand_x1_sg U49833 ( .A(n40655), .B(n57207), .X(n33797) );
  nand_x1_sg U49834 ( .A(n33790), .B(n33791), .X(n43271) );
  nand_x1_sg U49835 ( .A(n40654), .B(n57207), .X(n33791) );
  nand_x1_sg U49836 ( .A(n33808), .B(n33809), .X(n43280) );
  nand_x1_sg U49837 ( .A(n40653), .B(n57207), .X(n33809) );
  nand_x1_sg U49838 ( .A(n33810), .B(n33811), .X(n43281) );
  nand_x1_sg U49839 ( .A(n40493), .B(n57207), .X(n33811) );
  nand_x1_sg U49840 ( .A(n33812), .B(n33813), .X(n43282) );
  nand_x1_sg U49841 ( .A(n40461), .B(n57207), .X(n33813) );
  nand_x1_sg U49842 ( .A(n33814), .B(n33815), .X(n43283) );
  nand_x1_sg U49843 ( .A(n40430), .B(n57207), .X(n33815) );
  nand_x1_sg U49844 ( .A(n33816), .B(n33817), .X(n43284) );
  nand_x1_sg U49845 ( .A(n40397), .B(n57207), .X(n33817) );
  nand_x1_sg U49846 ( .A(n33788), .B(n33789), .X(n43270) );
  nand_x1_sg U49847 ( .A(n40652), .B(n57207), .X(n33789) );
  nand_x1_sg U49848 ( .A(n33818), .B(n33819), .X(n43285) );
  nand_x1_sg U49849 ( .A(n40365), .B(n57207), .X(n33819) );
  nand_x1_sg U49850 ( .A(n33820), .B(n33821), .X(n43286) );
  nand_x1_sg U49851 ( .A(n40331), .B(n57207), .X(n33821) );
  nand_x1_sg U49852 ( .A(n33802), .B(n33803), .X(n43277) );
  nand_x1_sg U49853 ( .A(n40651), .B(n57207), .X(n33803) );
  nand_x1_sg U49854 ( .A(n33794), .B(n33795), .X(n43273) );
  nand_x1_sg U49855 ( .A(n40650), .B(n57207), .X(n33795) );
  nand_x1_sg U49856 ( .A(n33822), .B(n33823), .X(n43287) );
  nand_x1_sg U49857 ( .A(n40297), .B(n57207), .X(n33823) );
  nand_x1_sg U49858 ( .A(n33824), .B(n33825), .X(n43288) );
  nand_x1_sg U49859 ( .A(n40264), .B(n57207), .X(n33825) );
  nand_x1_sg U49860 ( .A(n33834), .B(n33835), .X(n43292) );
  nand_x1_sg U49861 ( .A(n40673), .B(n57204), .X(n33835) );
  nand_x1_sg U49862 ( .A(n33842), .B(n33843), .X(n43296) );
  nand_x1_sg U49863 ( .A(n40672), .B(n33828), .X(n33843) );
  nand_x1_sg U49864 ( .A(n33836), .B(n33837), .X(n43293) );
  nand_x1_sg U49865 ( .A(n40671), .B(n57204), .X(n33837) );
  nand_x1_sg U49866 ( .A(n33846), .B(n33847), .X(n43298) );
  nand_x1_sg U49867 ( .A(n40670), .B(n57204), .X(n33847) );
  nand_x1_sg U49868 ( .A(n33848), .B(n33849), .X(n43299) );
  nand_x1_sg U49869 ( .A(n40669), .B(n57204), .X(n33849) );
  nand_x1_sg U49870 ( .A(n33840), .B(n33841), .X(n43295) );
  nand_x1_sg U49871 ( .A(n40668), .B(n57204), .X(n33841) );
  nand_x1_sg U49872 ( .A(n33826), .B(n33827), .X(n43289) );
  nand_x1_sg U49873 ( .A(n40667), .B(n57204), .X(n33827) );
  nand_x1_sg U49874 ( .A(n33830), .B(n33831), .X(n43290) );
  nand_x1_sg U49875 ( .A(n40666), .B(n57204), .X(n33831) );
  nand_x1_sg U49876 ( .A(n33850), .B(n33851), .X(n43300) );
  nand_x1_sg U49877 ( .A(n40665), .B(n57204), .X(n33851) );
  nand_x1_sg U49878 ( .A(n33852), .B(n33853), .X(n43301) );
  nand_x1_sg U49879 ( .A(n40492), .B(n57204), .X(n33853) );
  nand_x1_sg U49880 ( .A(n33854), .B(n33855), .X(n43302) );
  nand_x1_sg U49881 ( .A(n40460), .B(n57204), .X(n33855) );
  nand_x1_sg U49882 ( .A(n33832), .B(n33833), .X(n43291) );
  nand_x1_sg U49883 ( .A(n40664), .B(n57204), .X(n33833) );
  nand_x1_sg U49884 ( .A(n33856), .B(n33857), .X(n43303) );
  nand_x1_sg U49885 ( .A(n40429), .B(n57204), .X(n33857) );
  nand_x1_sg U49886 ( .A(n33838), .B(n33839), .X(n43294) );
  nand_x1_sg U49887 ( .A(n40663), .B(n57204), .X(n33839) );
  nand_x1_sg U49888 ( .A(n33858), .B(n33859), .X(n43304) );
  nand_x1_sg U49889 ( .A(n40396), .B(n57204), .X(n33859) );
  nand_x1_sg U49890 ( .A(n33860), .B(n33861), .X(n43305) );
  nand_x1_sg U49891 ( .A(n40364), .B(n57204), .X(n33861) );
  nand_x1_sg U49892 ( .A(n33844), .B(n33845), .X(n43297) );
  nand_x1_sg U49893 ( .A(n40662), .B(n57204), .X(n33845) );
  nand_x1_sg U49894 ( .A(n33862), .B(n33863), .X(n43306) );
  nand_x1_sg U49895 ( .A(n40330), .B(n57204), .X(n33863) );
  nand_x1_sg U49896 ( .A(n33864), .B(n33865), .X(n43307) );
  nand_x1_sg U49897 ( .A(n40296), .B(n57204), .X(n33865) );
  nand_x1_sg U49898 ( .A(n33866), .B(n33867), .X(n43308) );
  nand_x1_sg U49899 ( .A(n40241), .B(n57204), .X(n33867) );
  nand_x1_sg U49900 ( .A(n33877), .B(n33878), .X(n43312) );
  nand_x1_sg U49901 ( .A(n40686), .B(n57201), .X(n33878) );
  nand_x1_sg U49902 ( .A(n33885), .B(n33886), .X(n43316) );
  nand_x1_sg U49903 ( .A(n40685), .B(n57201), .X(n33886) );
  nand_x1_sg U49904 ( .A(n33879), .B(n33880), .X(n43313) );
  nand_x1_sg U49905 ( .A(n40684), .B(n57201), .X(n33880) );
  nand_x1_sg U49906 ( .A(n33889), .B(n33890), .X(n43318) );
  nand_x1_sg U49907 ( .A(n40683), .B(n57201), .X(n33890) );
  nand_x1_sg U49908 ( .A(n33891), .B(n33892), .X(n43319) );
  nand_x1_sg U49909 ( .A(n40682), .B(n57201), .X(n33892) );
  nand_x1_sg U49910 ( .A(n33883), .B(n33884), .X(n43315) );
  nand_x1_sg U49911 ( .A(n40681), .B(n57201), .X(n33884) );
  nand_x1_sg U49912 ( .A(n33869), .B(n33870), .X(n43309) );
  nand_x1_sg U49913 ( .A(n40680), .B(n57201), .X(n33870) );
  nand_x1_sg U49914 ( .A(n33873), .B(n33874), .X(n43310) );
  nand_x1_sg U49915 ( .A(n40679), .B(n57201), .X(n33874) );
  nand_x1_sg U49916 ( .A(n33893), .B(n33894), .X(n43320) );
  nand_x1_sg U49917 ( .A(n40678), .B(n57201), .X(n33894) );
  nand_x1_sg U49918 ( .A(n33895), .B(n33896), .X(n43321) );
  nand_x1_sg U49919 ( .A(n40677), .B(n57201), .X(n33896) );
  nand_x1_sg U49920 ( .A(n33897), .B(n33898), .X(n43322) );
  nand_x1_sg U49921 ( .A(n40491), .B(n57201), .X(n33898) );
  nand_x1_sg U49922 ( .A(n33875), .B(n33876), .X(n43311) );
  nand_x1_sg U49923 ( .A(n40676), .B(n57201), .X(n33876) );
  nand_x1_sg U49924 ( .A(n33899), .B(n33900), .X(n43323) );
  nand_x1_sg U49925 ( .A(n40459), .B(n57201), .X(n33900) );
  nand_x1_sg U49926 ( .A(n33881), .B(n33882), .X(n43314) );
  nand_x1_sg U49927 ( .A(n40675), .B(n57201), .X(n33882) );
  nand_x1_sg U49928 ( .A(n33901), .B(n33902), .X(n43324) );
  nand_x1_sg U49929 ( .A(n40428), .B(n57201), .X(n33902) );
  nand_x1_sg U49930 ( .A(n33903), .B(n33904), .X(n43325) );
  nand_x1_sg U49931 ( .A(n40395), .B(n57201), .X(n33904) );
  nand_x1_sg U49932 ( .A(n33887), .B(n33888), .X(n43317) );
  nand_x1_sg U49933 ( .A(n40674), .B(n33871), .X(n33888) );
  nand_x1_sg U49934 ( .A(n33905), .B(n33906), .X(n43326) );
  nand_x1_sg U49935 ( .A(n40363), .B(n57201), .X(n33906) );
  nand_x1_sg U49936 ( .A(n33907), .B(n33908), .X(n43327) );
  nand_x1_sg U49937 ( .A(n40329), .B(n57201), .X(n33908) );
  nand_x1_sg U49938 ( .A(n33909), .B(n33910), .X(n43328) );
  nand_x1_sg U49939 ( .A(n40295), .B(n57201), .X(n33910) );
  nand_x1_sg U49940 ( .A(n33406), .B(n33407), .X(n43092) );
  nand_x1_sg U49941 ( .A(n40698), .B(n57240), .X(n33407) );
  nand_x1_sg U49942 ( .A(n33414), .B(n33415), .X(n43096) );
  nand_x1_sg U49943 ( .A(n40697), .B(n57240), .X(n33415) );
  nand_x1_sg U49944 ( .A(n33398), .B(n33399), .X(n43089) );
  nand_x1_sg U49945 ( .A(n40696), .B(n57240), .X(n33399) );
  nand_x1_sg U49946 ( .A(n33418), .B(n33419), .X(n43098) );
  nand_x1_sg U49947 ( .A(n40695), .B(n57240), .X(n33419) );
  nand_x1_sg U49948 ( .A(n33420), .B(n33421), .X(n43099) );
  nand_x1_sg U49949 ( .A(n40694), .B(n57240), .X(n33421) );
  nand_x1_sg U49950 ( .A(n33412), .B(n33413), .X(n43095) );
  nand_x1_sg U49951 ( .A(n40693), .B(n57240), .X(n33413) );
  nand_x1_sg U49952 ( .A(n33410), .B(n33411), .X(n43094) );
  nand_x1_sg U49953 ( .A(n40692), .B(n57240), .X(n33411) );
  nand_x1_sg U49954 ( .A(n33404), .B(n33405), .X(n43091) );
  nand_x1_sg U49955 ( .A(n40691), .B(n57240), .X(n33405) );
  nand_x1_sg U49956 ( .A(n33422), .B(n33423), .X(n43100) );
  nand_x1_sg U49957 ( .A(n40690), .B(n57240), .X(n33423) );
  nand_x1_sg U49958 ( .A(n33424), .B(n33425), .X(n43101) );
  nand_x1_sg U49959 ( .A(n40490), .B(n57240), .X(n33425) );
  nand_x1_sg U49960 ( .A(n33426), .B(n33427), .X(n43102) );
  nand_x1_sg U49961 ( .A(n40458), .B(n57240), .X(n33427) );
  nand_x1_sg U49962 ( .A(n33428), .B(n33429), .X(n43103) );
  nand_x1_sg U49963 ( .A(n40427), .B(n57240), .X(n33429) );
  nand_x1_sg U49964 ( .A(n33430), .B(n33431), .X(n43104) );
  nand_x1_sg U49965 ( .A(n40394), .B(n57240), .X(n33431) );
  nand_x1_sg U49966 ( .A(n33402), .B(n33403), .X(n43090) );
  nand_x1_sg U49967 ( .A(n40689), .B(n57240), .X(n33403) );
  nand_x1_sg U49968 ( .A(n33432), .B(n33433), .X(n43105) );
  nand_x1_sg U49969 ( .A(n40362), .B(n57240), .X(n33433) );
  nand_x1_sg U49970 ( .A(n33434), .B(n33435), .X(n43106) );
  nand_x1_sg U49971 ( .A(n40328), .B(n33400), .X(n33435) );
  nand_x1_sg U49972 ( .A(n33416), .B(n33417), .X(n43097) );
  nand_x1_sg U49973 ( .A(n40688), .B(n57240), .X(n33417) );
  nand_x1_sg U49974 ( .A(n33408), .B(n33409), .X(n43093) );
  nand_x1_sg U49975 ( .A(n40687), .B(n57240), .X(n33409) );
  nand_x1_sg U49976 ( .A(n33436), .B(n33437), .X(n43107) );
  nand_x1_sg U49977 ( .A(n40294), .B(n57240), .X(n33437) );
  nand_x1_sg U49978 ( .A(n33438), .B(n33439), .X(n43108) );
  nand_x1_sg U49979 ( .A(n40263), .B(n57240), .X(n33439) );
  nand_x1_sg U49980 ( .A(n33448), .B(n33449), .X(n43112) );
  nand_x1_sg U49981 ( .A(n40710), .B(n57236), .X(n33449) );
  nand_x1_sg U49982 ( .A(n33456), .B(n33457), .X(n43116) );
  nand_x1_sg U49983 ( .A(n40709), .B(n57236), .X(n33457) );
  nand_x1_sg U49984 ( .A(n33440), .B(n33441), .X(n43109) );
  nand_x1_sg U49985 ( .A(n40708), .B(n57236), .X(n33441) );
  nand_x1_sg U49986 ( .A(n33460), .B(n33461), .X(n43118) );
  nand_x1_sg U49987 ( .A(n40707), .B(n57236), .X(n33461) );
  nand_x1_sg U49988 ( .A(n33462), .B(n33463), .X(n43119) );
  nand_x1_sg U49989 ( .A(n40706), .B(n57236), .X(n33463) );
  nand_x1_sg U49990 ( .A(n33454), .B(n33455), .X(n43115) );
  nand_x1_sg U49991 ( .A(n40705), .B(n57236), .X(n33455) );
  nand_x1_sg U49992 ( .A(n33452), .B(n33453), .X(n43114) );
  nand_x1_sg U49993 ( .A(n40704), .B(n57236), .X(n33453) );
  nand_x1_sg U49994 ( .A(n33446), .B(n33447), .X(n43111) );
  nand_x1_sg U49995 ( .A(n40703), .B(n57236), .X(n33447) );
  nand_x1_sg U49996 ( .A(n33464), .B(n33465), .X(n43120) );
  nand_x1_sg U49997 ( .A(n40702), .B(n57236), .X(n33465) );
  nand_x1_sg U49998 ( .A(n33466), .B(n33467), .X(n43121) );
  nand_x1_sg U49999 ( .A(n40489), .B(n57236), .X(n33467) );
  nand_x1_sg U50000 ( .A(n33468), .B(n33469), .X(n43122) );
  nand_x1_sg U50001 ( .A(n40457), .B(n57236), .X(n33469) );
  nand_x1_sg U50002 ( .A(n33470), .B(n33471), .X(n43123) );
  nand_x1_sg U50003 ( .A(n40426), .B(n57236), .X(n33471) );
  nand_x1_sg U50004 ( .A(n33472), .B(n33473), .X(n43124) );
  nand_x1_sg U50005 ( .A(n40393), .B(n57236), .X(n33473) );
  nand_x1_sg U50006 ( .A(n33444), .B(n33445), .X(n43110) );
  nand_x1_sg U50007 ( .A(n40701), .B(n57236), .X(n33445) );
  nand_x1_sg U50008 ( .A(n33474), .B(n33475), .X(n43125) );
  nand_x1_sg U50009 ( .A(n40361), .B(n57236), .X(n33475) );
  nand_x1_sg U50010 ( .A(n33476), .B(n33477), .X(n43126) );
  nand_x1_sg U50011 ( .A(n40327), .B(n33442), .X(n33477) );
  nand_x1_sg U50012 ( .A(n33458), .B(n33459), .X(n43117) );
  nand_x1_sg U50013 ( .A(n40700), .B(n57236), .X(n33459) );
  nand_x1_sg U50014 ( .A(n33450), .B(n33451), .X(n43113) );
  nand_x1_sg U50015 ( .A(n40699), .B(n57236), .X(n33451) );
  nand_x1_sg U50016 ( .A(n33478), .B(n33479), .X(n43127) );
  nand_x1_sg U50017 ( .A(n40293), .B(n57236), .X(n33479) );
  nand_x1_sg U50018 ( .A(n33480), .B(n33481), .X(n43128) );
  nand_x1_sg U50019 ( .A(n40262), .B(n57236), .X(n33481) );
  nand_x1_sg U50020 ( .A(n33047), .B(n33048), .X(n42927) );
  nand_x1_sg U50021 ( .A(n40722), .B(n57276), .X(n33048) );
  nand_x1_sg U50022 ( .A(n33027), .B(n33028), .X(n42917) );
  nand_x1_sg U50023 ( .A(n40721), .B(n33011), .X(n33028) );
  nand_x1_sg U50024 ( .A(n33017), .B(n33018), .X(n42912) );
  nand_x1_sg U50025 ( .A(n40720), .B(n57276), .X(n33018) );
  nand_x1_sg U50026 ( .A(n33019), .B(n33020), .X(n42913) );
  nand_x1_sg U50027 ( .A(n40719), .B(n57276), .X(n33020) );
  nand_x1_sg U50028 ( .A(n33035), .B(n33036), .X(n42921) );
  nand_x1_sg U50029 ( .A(n40718), .B(n57276), .X(n33036) );
  nand_x1_sg U50030 ( .A(n33045), .B(n33046), .X(n42926) );
  nand_x1_sg U50031 ( .A(n40717), .B(n57276), .X(n33046) );
  nand_x1_sg U50032 ( .A(n33041), .B(n33042), .X(n42924) );
  nand_x1_sg U50033 ( .A(n40716), .B(n57276), .X(n33042) );
  nand_x1_sg U50034 ( .A(n33013), .B(n33014), .X(n42910) );
  nand_x1_sg U50035 ( .A(n40715), .B(n57276), .X(n33014) );
  nand_x1_sg U50036 ( .A(n33025), .B(n33026), .X(n42916) );
  nand_x1_sg U50037 ( .A(n40714), .B(n57276), .X(n33026) );
  nand_x1_sg U50038 ( .A(n33009), .B(n33010), .X(n42909) );
  nand_x1_sg U50039 ( .A(n40488), .B(n57276), .X(n33010) );
  nand_x1_sg U50040 ( .A(n33037), .B(n33038), .X(n42922) );
  nand_x1_sg U50041 ( .A(n40456), .B(n57276), .X(n33038) );
  nand_x1_sg U50042 ( .A(n33029), .B(n33030), .X(n42918) );
  nand_x1_sg U50043 ( .A(n40425), .B(n57276), .X(n33030) );
  nand_x1_sg U50044 ( .A(n33049), .B(n33050), .X(n42928) );
  nand_x1_sg U50045 ( .A(n40392), .B(n57276), .X(n33050) );
  nand_x1_sg U50046 ( .A(n33023), .B(n33024), .X(n42915) );
  nand_x1_sg U50047 ( .A(n40360), .B(n57276), .X(n33024) );
  nand_x1_sg U50048 ( .A(n33031), .B(n33032), .X(n42919) );
  nand_x1_sg U50049 ( .A(n40713), .B(n57276), .X(n33032) );
  nand_x1_sg U50050 ( .A(n33039), .B(n33040), .X(n42923) );
  nand_x1_sg U50051 ( .A(n40326), .B(n57276), .X(n33040) );
  nand_x1_sg U50052 ( .A(n33043), .B(n33044), .X(n42925) );
  nand_x1_sg U50053 ( .A(n40712), .B(n57276), .X(n33044) );
  nand_x1_sg U50054 ( .A(n33015), .B(n33016), .X(n42911) );
  nand_x1_sg U50055 ( .A(n40292), .B(n57276), .X(n33016) );
  nand_x1_sg U50056 ( .A(n33021), .B(n33022), .X(n42914) );
  nand_x1_sg U50057 ( .A(n40711), .B(n57276), .X(n33022) );
  nand_x1_sg U50058 ( .A(n33033), .B(n33034), .X(n42920) );
  nand_x1_sg U50059 ( .A(n40261), .B(n57276), .X(n33034) );
  nand_x1_sg U50060 ( .A(n34185), .B(n34186), .X(n43452) );
  nand_x1_sg U50061 ( .A(n40735), .B(n57174), .X(n34186) );
  nand_x1_sg U50062 ( .A(n34201), .B(n34202), .X(n43460) );
  nand_x1_sg U50063 ( .A(n40734), .B(n57174), .X(n34202) );
  nand_x1_sg U50064 ( .A(n34181), .B(n34182), .X(n43450) );
  nand_x1_sg U50065 ( .A(n40733), .B(n57174), .X(n34182) );
  nand_x1_sg U50066 ( .A(n34205), .B(n34206), .X(n43462) );
  nand_x1_sg U50067 ( .A(n40732), .B(n57174), .X(n34206) );
  nand_x1_sg U50068 ( .A(n34207), .B(n34208), .X(n43463) );
  nand_x1_sg U50069 ( .A(n40731), .B(n57174), .X(n34208) );
  nand_x1_sg U50070 ( .A(n34189), .B(n34190), .X(n43454) );
  nand_x1_sg U50071 ( .A(n40730), .B(n57174), .X(n34190) );
  nand_x1_sg U50072 ( .A(n34199), .B(n34200), .X(n43459) );
  nand_x1_sg U50073 ( .A(n40729), .B(n57174), .X(n34200) );
  nand_x1_sg U50074 ( .A(n34191), .B(n34192), .X(n43455) );
  nand_x1_sg U50075 ( .A(n40728), .B(n57174), .X(n34192) );
  nand_x1_sg U50076 ( .A(n34209), .B(n34210), .X(n43464) );
  nand_x1_sg U50077 ( .A(n40727), .B(n57174), .X(n34210) );
  nand_x1_sg U50078 ( .A(n34195), .B(n34196), .X(n43457) );
  nand_x1_sg U50079 ( .A(n40726), .B(n34179), .X(n34196) );
  nand_x1_sg U50080 ( .A(n34211), .B(n34212), .X(n43465) );
  nand_x1_sg U50081 ( .A(n40487), .B(n57174), .X(n34212) );
  nand_x1_sg U50082 ( .A(n34193), .B(n34194), .X(n43456) );
  nand_x1_sg U50083 ( .A(n40455), .B(n57174), .X(n34194) );
  nand_x1_sg U50084 ( .A(n34177), .B(n34178), .X(n43449) );
  nand_x1_sg U50085 ( .A(n40424), .B(n57174), .X(n34178) );
  nand_x1_sg U50086 ( .A(n34197), .B(n34198), .X(n43458) );
  nand_x1_sg U50087 ( .A(n40725), .B(n57174), .X(n34198) );
  nand_x1_sg U50088 ( .A(n34213), .B(n34214), .X(n43466) );
  nand_x1_sg U50089 ( .A(n40391), .B(n57174), .X(n34214) );
  nand_x1_sg U50090 ( .A(n34187), .B(n34188), .X(n43453) );
  nand_x1_sg U50091 ( .A(n40359), .B(n57174), .X(n34188) );
  nand_x1_sg U50092 ( .A(n34203), .B(n34204), .X(n43461) );
  nand_x1_sg U50093 ( .A(n40724), .B(n57174), .X(n34204) );
  nand_x1_sg U50094 ( .A(n34183), .B(n34184), .X(n43451) );
  nand_x1_sg U50095 ( .A(n40723), .B(n57174), .X(n34184) );
  nand_x1_sg U50096 ( .A(n34215), .B(n34216), .X(n43467) );
  nand_x1_sg U50097 ( .A(n40325), .B(n57174), .X(n34216) );
  nand_x1_sg U50098 ( .A(n34217), .B(n34218), .X(n43468) );
  nand_x1_sg U50099 ( .A(n40291), .B(n57174), .X(n34218) );
  nand_x1_sg U50100 ( .A(n33275), .B(n33276), .X(n43032) );
  nand_x1_sg U50101 ( .A(n40747), .B(n57252), .X(n33276) );
  nand_x1_sg U50102 ( .A(n33283), .B(n33284), .X(n43036) );
  nand_x1_sg U50103 ( .A(n40746), .B(n57252), .X(n33284) );
  nand_x1_sg U50104 ( .A(n33267), .B(n33268), .X(n43029) );
  nand_x1_sg U50105 ( .A(n40745), .B(n57252), .X(n33268) );
  nand_x1_sg U50106 ( .A(n33287), .B(n33288), .X(n43038) );
  nand_x1_sg U50107 ( .A(n40744), .B(n57252), .X(n33288) );
  nand_x1_sg U50108 ( .A(n33289), .B(n33290), .X(n43039) );
  nand_x1_sg U50109 ( .A(n40743), .B(n57252), .X(n33290) );
  nand_x1_sg U50110 ( .A(n33281), .B(n33282), .X(n43035) );
  nand_x1_sg U50111 ( .A(n40742), .B(n57252), .X(n33282) );
  nand_x1_sg U50112 ( .A(n33279), .B(n33280), .X(n43034) );
  nand_x1_sg U50113 ( .A(n40741), .B(n57252), .X(n33280) );
  nand_x1_sg U50114 ( .A(n33273), .B(n33274), .X(n43031) );
  nand_x1_sg U50115 ( .A(n40740), .B(n57252), .X(n33274) );
  nand_x1_sg U50116 ( .A(n33291), .B(n33292), .X(n43040) );
  nand_x1_sg U50117 ( .A(n40739), .B(n57252), .X(n33292) );
  nand_x1_sg U50118 ( .A(n33293), .B(n33294), .X(n43041) );
  nand_x1_sg U50119 ( .A(n40486), .B(n57252), .X(n33294) );
  nand_x1_sg U50120 ( .A(n33295), .B(n33296), .X(n43042) );
  nand_x1_sg U50121 ( .A(n40454), .B(n57252), .X(n33296) );
  nand_x1_sg U50122 ( .A(n33297), .B(n33298), .X(n43043) );
  nand_x1_sg U50123 ( .A(n40423), .B(n57252), .X(n33298) );
  nand_x1_sg U50124 ( .A(n33299), .B(n33300), .X(n43044) );
  nand_x1_sg U50125 ( .A(n40390), .B(n57252), .X(n33300) );
  nand_x1_sg U50126 ( .A(n33271), .B(n33272), .X(n43030) );
  nand_x1_sg U50127 ( .A(n40738), .B(n57252), .X(n33272) );
  nand_x1_sg U50128 ( .A(n33301), .B(n33302), .X(n43045) );
  nand_x1_sg U50129 ( .A(n40358), .B(n57252), .X(n33302) );
  nand_x1_sg U50130 ( .A(n33303), .B(n33304), .X(n43046) );
  nand_x1_sg U50131 ( .A(n40324), .B(n33269), .X(n33304) );
  nand_x1_sg U50132 ( .A(n33285), .B(n33286), .X(n43037) );
  nand_x1_sg U50133 ( .A(n40737), .B(n57252), .X(n33286) );
  nand_x1_sg U50134 ( .A(n33277), .B(n33278), .X(n43033) );
  nand_x1_sg U50135 ( .A(n40736), .B(n57252), .X(n33278) );
  nand_x1_sg U50136 ( .A(n33305), .B(n33306), .X(n43047) );
  nand_x1_sg U50137 ( .A(n40290), .B(n57252), .X(n33306) );
  nand_x1_sg U50138 ( .A(n33307), .B(n33308), .X(n43048) );
  nand_x1_sg U50139 ( .A(n40260), .B(n57252), .X(n33308) );
  nand_x1_sg U50140 ( .A(n33319), .B(n33320), .X(n43052) );
  nand_x1_sg U50141 ( .A(n40759), .B(n57248), .X(n33320) );
  nand_x1_sg U50142 ( .A(n33327), .B(n33328), .X(n43056) );
  nand_x1_sg U50143 ( .A(n40758), .B(n57248), .X(n33328) );
  nand_x1_sg U50144 ( .A(n33321), .B(n33322), .X(n43053) );
  nand_x1_sg U50145 ( .A(n40757), .B(n57248), .X(n33322) );
  nand_x1_sg U50146 ( .A(n33331), .B(n33332), .X(n43058) );
  nand_x1_sg U50147 ( .A(n40756), .B(n57248), .X(n33332) );
  nand_x1_sg U50148 ( .A(n33333), .B(n33334), .X(n43059) );
  nand_x1_sg U50149 ( .A(n40755), .B(n57248), .X(n33334) );
  nand_x1_sg U50150 ( .A(n33325), .B(n33326), .X(n43055) );
  nand_x1_sg U50151 ( .A(n40754), .B(n57248), .X(n33326) );
  nand_x1_sg U50152 ( .A(n33311), .B(n33312), .X(n43049) );
  nand_x1_sg U50153 ( .A(n40753), .B(n57248), .X(n33312) );
  nand_x1_sg U50154 ( .A(n33315), .B(n33316), .X(n43050) );
  nand_x1_sg U50155 ( .A(n40752), .B(n57248), .X(n33316) );
  nand_x1_sg U50156 ( .A(n33335), .B(n33336), .X(n43060) );
  nand_x1_sg U50157 ( .A(n40751), .B(n57248), .X(n33336) );
  nand_x1_sg U50158 ( .A(n33337), .B(n33338), .X(n43061) );
  nand_x1_sg U50159 ( .A(n40485), .B(n57248), .X(n33338) );
  nand_x1_sg U50160 ( .A(n33339), .B(n33340), .X(n43062) );
  nand_x1_sg U50161 ( .A(n40453), .B(n57248), .X(n33340) );
  nand_x1_sg U50162 ( .A(n33317), .B(n33318), .X(n43051) );
  nand_x1_sg U50163 ( .A(n40750), .B(n57248), .X(n33318) );
  nand_x1_sg U50164 ( .A(n33341), .B(n33342), .X(n43063) );
  nand_x1_sg U50165 ( .A(n40422), .B(n57248), .X(n33342) );
  nand_x1_sg U50166 ( .A(n33323), .B(n33324), .X(n43054) );
  nand_x1_sg U50167 ( .A(n40749), .B(n57248), .X(n33324) );
  nand_x1_sg U50168 ( .A(n33343), .B(n33344), .X(n43064) );
  nand_x1_sg U50169 ( .A(n40389), .B(n57248), .X(n33344) );
  nand_x1_sg U50170 ( .A(n33345), .B(n33346), .X(n43065) );
  nand_x1_sg U50171 ( .A(n40357), .B(n57248), .X(n33346) );
  nand_x1_sg U50172 ( .A(n33329), .B(n33330), .X(n43057) );
  nand_x1_sg U50173 ( .A(n40748), .B(n33313), .X(n33330) );
  nand_x1_sg U50174 ( .A(n33347), .B(n33348), .X(n43066) );
  nand_x1_sg U50175 ( .A(n40323), .B(n57248), .X(n33348) );
  nand_x1_sg U50176 ( .A(n33349), .B(n33350), .X(n43067) );
  nand_x1_sg U50177 ( .A(n40289), .B(n57248), .X(n33350) );
  nand_x1_sg U50178 ( .A(n33351), .B(n33352), .X(n43068) );
  nand_x1_sg U50179 ( .A(n40259), .B(n57248), .X(n33352) );
  nand_x1_sg U50180 ( .A(n33373), .B(n33374), .X(n43078) );
  nand_x1_sg U50181 ( .A(n40770), .B(n57244), .X(n33374) );
  nand_x1_sg U50182 ( .A(n33369), .B(n33370), .X(n43076) );
  nand_x1_sg U50183 ( .A(n40769), .B(n57244), .X(n33370) );
  nand_x1_sg U50184 ( .A(n33375), .B(n33376), .X(n43079) );
  nand_x1_sg U50185 ( .A(n40768), .B(n57244), .X(n33376) );
  nand_x1_sg U50186 ( .A(n33377), .B(n33378), .X(n43080) );
  nand_x1_sg U50187 ( .A(n40484), .B(n57244), .X(n33378) );
  nand_x1_sg U50188 ( .A(n33361), .B(n33362), .X(n43072) );
  nand_x1_sg U50189 ( .A(n40767), .B(n57244), .X(n33362) );
  nand_x1_sg U50190 ( .A(n33367), .B(n33368), .X(n43075) );
  nand_x1_sg U50191 ( .A(n40766), .B(n57244), .X(n33368) );
  nand_x1_sg U50192 ( .A(n33379), .B(n33380), .X(n43081) );
  nand_x1_sg U50193 ( .A(n40452), .B(n57244), .X(n33380) );
  nand_x1_sg U50194 ( .A(n33381), .B(n33382), .X(n43082) );
  nand_x1_sg U50195 ( .A(n40421), .B(n57244), .X(n33382) );
  nand_x1_sg U50196 ( .A(n33357), .B(n33358), .X(n43070) );
  nand_x1_sg U50197 ( .A(n40765), .B(n57244), .X(n33358) );
  nand_x1_sg U50198 ( .A(n33383), .B(n33384), .X(n43083) );
  nand_x1_sg U50199 ( .A(n40388), .B(n57244), .X(n33384) );
  nand_x1_sg U50200 ( .A(n33365), .B(n33366), .X(n43074) );
  nand_x1_sg U50201 ( .A(n40764), .B(n57244), .X(n33366) );
  nand_x1_sg U50202 ( .A(n33385), .B(n33386), .X(n43084) );
  nand_x1_sg U50203 ( .A(n40356), .B(n57244), .X(n33386) );
  nand_x1_sg U50204 ( .A(n33359), .B(n33360), .X(n43071) );
  nand_x1_sg U50205 ( .A(n40763), .B(n57244), .X(n33360) );
  nand_x1_sg U50206 ( .A(n33387), .B(n33388), .X(n43085) );
  nand_x1_sg U50207 ( .A(n40322), .B(n57244), .X(n33388) );
  nand_x1_sg U50208 ( .A(n33363), .B(n33364), .X(n43073) );
  nand_x1_sg U50209 ( .A(n40762), .B(n57244), .X(n33364) );
  nand_x1_sg U50210 ( .A(n33389), .B(n33390), .X(n43086) );
  nand_x1_sg U50211 ( .A(n40288), .B(n33355), .X(n33390) );
  nand_x1_sg U50212 ( .A(n33371), .B(n33372), .X(n43077) );
  nand_x1_sg U50213 ( .A(n40761), .B(n57244), .X(n33372) );
  nand_x1_sg U50214 ( .A(n33391), .B(n33392), .X(n43087) );
  nand_x1_sg U50215 ( .A(n40258), .B(n57244), .X(n33392) );
  nand_x1_sg U50216 ( .A(n33353), .B(n33354), .X(n43069) );
  nand_x1_sg U50217 ( .A(n40760), .B(n57244), .X(n33354) );
  nand_x1_sg U50218 ( .A(n33393), .B(n33394), .X(n43088) );
  nand_x1_sg U50219 ( .A(n40240), .B(n57244), .X(n33394) );
  nand_x1_sg U50220 ( .A(n32836), .B(n32837), .X(n42830) );
  nand_x1_sg U50221 ( .A(n40774), .B(n57292), .X(n32837) );
  nand_x1_sg U50222 ( .A(n32838), .B(n32839), .X(n42831) );
  nand_x1_sg U50223 ( .A(n40773), .B(n57292), .X(n32839) );
  nand_x1_sg U50224 ( .A(n32840), .B(n32841), .X(n42832) );
  nand_x1_sg U50225 ( .A(n40772), .B(n57292), .X(n32841) );
  nand_x1_sg U50226 ( .A(n32842), .B(n32843), .X(n42833) );
  nand_x1_sg U50227 ( .A(n40771), .B(n57292), .X(n32843) );
  nand_x1_sg U50228 ( .A(n32844), .B(n32845), .X(n42834) );
  nand_x1_sg U50229 ( .A(n40483), .B(n57292), .X(n32845) );
  nand_x1_sg U50230 ( .A(n32846), .B(n32847), .X(n42835) );
  nand_x1_sg U50231 ( .A(n40451), .B(n57292), .X(n32847) );
  nand_x1_sg U50232 ( .A(n32850), .B(n32851), .X(n42837) );
  nand_x1_sg U50233 ( .A(n40355), .B(n57292), .X(n32851) );
  nand_x1_sg U50234 ( .A(n32848), .B(n32849), .X(n42836) );
  nand_x1_sg U50235 ( .A(n40420), .B(n57292), .X(n32849) );
  nand_x1_sg U50236 ( .A(n32852), .B(n32853), .X(n42838) );
  nand_x1_sg U50237 ( .A(n40321), .B(n57292), .X(n32853) );
  nand_x1_sg U50238 ( .A(n32862), .B(n32863), .X(n42843) );
  nand_x1_sg U50239 ( .A(n40354), .B(n57292), .X(n32863) );
  nand_x1_sg U50240 ( .A(n32854), .B(n32855), .X(n42839) );
  nand_x1_sg U50241 ( .A(n40287), .B(n57292), .X(n32855) );
  nand_x1_sg U50242 ( .A(n32864), .B(n32865), .X(n42844) );
  nand_x1_sg U50243 ( .A(n40320), .B(n57292), .X(n32865) );
  nand_x1_sg U50244 ( .A(n32856), .B(n32857), .X(n42840) );
  nand_x1_sg U50245 ( .A(n40257), .B(n57292), .X(n32857) );
  nand_x1_sg U50246 ( .A(n32866), .B(n32867), .X(n42845) );
  nand_x1_sg U50247 ( .A(n40286), .B(n57292), .X(n32867) );
  nand_x1_sg U50248 ( .A(n32858), .B(n32859), .X(n42841) );
  nand_x1_sg U50249 ( .A(n40239), .B(n32834), .X(n32859) );
  nand_x1_sg U50250 ( .A(n32868), .B(n32869), .X(n42846) );
  nand_x1_sg U50251 ( .A(n40256), .B(n57292), .X(n32869) );
  nand_x1_sg U50252 ( .A(n32832), .B(n32833), .X(n42829) );
  nand_x1_sg U50253 ( .A(n40232), .B(n57292), .X(n32833) );
  nand_x1_sg U50254 ( .A(n32870), .B(n32871), .X(n42847) );
  nand_x1_sg U50255 ( .A(n40238), .B(n57292), .X(n32871) );
  nand_x1_sg U50256 ( .A(n32860), .B(n32861), .X(n42842) );
  nand_x1_sg U50257 ( .A(n40229), .B(n57292), .X(n32861) );
  nand_x1_sg U50258 ( .A(n32872), .B(n32873), .X(n42848) );
  nand_x1_sg U50259 ( .A(n40228), .B(n57292), .X(n32873) );
  nand_x1_sg U50260 ( .A(n33490), .B(n33491), .X(n43132) );
  nand_x1_sg U50261 ( .A(n40785), .B(n57232), .X(n33491) );
  nand_x1_sg U50262 ( .A(n33498), .B(n33499), .X(n43136) );
  nand_x1_sg U50263 ( .A(n40784), .B(n33484), .X(n33499) );
  nand_x1_sg U50264 ( .A(n33482), .B(n33483), .X(n43129) );
  nand_x1_sg U50265 ( .A(n40783), .B(n57232), .X(n33483) );
  nand_x1_sg U50266 ( .A(n33502), .B(n33503), .X(n43138) );
  nand_x1_sg U50267 ( .A(n40782), .B(n57232), .X(n33503) );
  nand_x1_sg U50268 ( .A(n33504), .B(n33505), .X(n43139) );
  nand_x1_sg U50269 ( .A(n40781), .B(n57232), .X(n33505) );
  nand_x1_sg U50270 ( .A(n33496), .B(n33497), .X(n43135) );
  nand_x1_sg U50271 ( .A(n40780), .B(n57232), .X(n33497) );
  nand_x1_sg U50272 ( .A(n33494), .B(n33495), .X(n43134) );
  nand_x1_sg U50273 ( .A(n40779), .B(n57232), .X(n33495) );
  nand_x1_sg U50274 ( .A(n33488), .B(n33489), .X(n43131) );
  nand_x1_sg U50275 ( .A(n40778), .B(n57232), .X(n33489) );
  nand_x1_sg U50276 ( .A(n33506), .B(n33507), .X(n43140) );
  nand_x1_sg U50277 ( .A(n40482), .B(n57232), .X(n33507) );
  nand_x1_sg U50278 ( .A(n33508), .B(n33509), .X(n43141) );
  nand_x1_sg U50279 ( .A(n40450), .B(n57232), .X(n33509) );
  nand_x1_sg U50280 ( .A(n33510), .B(n33511), .X(n43142) );
  nand_x1_sg U50281 ( .A(n40419), .B(n57232), .X(n33511) );
  nand_x1_sg U50282 ( .A(n33512), .B(n33513), .X(n43143) );
  nand_x1_sg U50283 ( .A(n40387), .B(n57232), .X(n33513) );
  nand_x1_sg U50284 ( .A(n33514), .B(n33515), .X(n43144) );
  nand_x1_sg U50285 ( .A(n40353), .B(n57232), .X(n33515) );
  nand_x1_sg U50286 ( .A(n33486), .B(n33487), .X(n43130) );
  nand_x1_sg U50287 ( .A(n40777), .B(n57232), .X(n33487) );
  nand_x1_sg U50288 ( .A(n33516), .B(n33517), .X(n43145) );
  nand_x1_sg U50289 ( .A(n40319), .B(n57232), .X(n33517) );
  nand_x1_sg U50290 ( .A(n33518), .B(n33519), .X(n43146) );
  nand_x1_sg U50291 ( .A(n40285), .B(n57232), .X(n33519) );
  nand_x1_sg U50292 ( .A(n33500), .B(n33501), .X(n43137) );
  nand_x1_sg U50293 ( .A(n40776), .B(n57232), .X(n33501) );
  nand_x1_sg U50294 ( .A(n33492), .B(n33493), .X(n43133) );
  nand_x1_sg U50295 ( .A(n40775), .B(n57232), .X(n33493) );
  nand_x1_sg U50296 ( .A(n33520), .B(n33521), .X(n43147) );
  nand_x1_sg U50297 ( .A(n40255), .B(n57232), .X(n33521) );
  nand_x1_sg U50298 ( .A(n33522), .B(n33523), .X(n43148) );
  nand_x1_sg U50299 ( .A(n40237), .B(n57232), .X(n33523) );
  nand_x1_sg U50300 ( .A(n33533), .B(n33534), .X(n43152) );
  nand_x1_sg U50301 ( .A(n40796), .B(n57229), .X(n33534) );
  nand_x1_sg U50302 ( .A(n33541), .B(n33542), .X(n43156) );
  nand_x1_sg U50303 ( .A(n40795), .B(n33527), .X(n33542) );
  nand_x1_sg U50304 ( .A(n33535), .B(n33536), .X(n43153) );
  nand_x1_sg U50305 ( .A(n40794), .B(n57229), .X(n33536) );
  nand_x1_sg U50306 ( .A(n33545), .B(n33546), .X(n43158) );
  nand_x1_sg U50307 ( .A(n40793), .B(n57229), .X(n33546) );
  nand_x1_sg U50308 ( .A(n33547), .B(n33548), .X(n43159) );
  nand_x1_sg U50309 ( .A(n40792), .B(n57229), .X(n33548) );
  nand_x1_sg U50310 ( .A(n33539), .B(n33540), .X(n43155) );
  nand_x1_sg U50311 ( .A(n40791), .B(n57229), .X(n33540) );
  nand_x1_sg U50312 ( .A(n33525), .B(n33526), .X(n43149) );
  nand_x1_sg U50313 ( .A(n40790), .B(n57229), .X(n33526) );
  nand_x1_sg U50314 ( .A(n33529), .B(n33530), .X(n43150) );
  nand_x1_sg U50315 ( .A(n40789), .B(n57229), .X(n33530) );
  nand_x1_sg U50316 ( .A(n33549), .B(n33550), .X(n43160) );
  nand_x1_sg U50317 ( .A(n40481), .B(n57229), .X(n33550) );
  nand_x1_sg U50318 ( .A(n33551), .B(n33552), .X(n43161) );
  nand_x1_sg U50319 ( .A(n40449), .B(n57229), .X(n33552) );
  nand_x1_sg U50320 ( .A(n33553), .B(n33554), .X(n43162) );
  nand_x1_sg U50321 ( .A(n40418), .B(n57229), .X(n33554) );
  nand_x1_sg U50322 ( .A(n33531), .B(n33532), .X(n43151) );
  nand_x1_sg U50323 ( .A(n40788), .B(n57229), .X(n33532) );
  nand_x1_sg U50324 ( .A(n33555), .B(n33556), .X(n43163) );
  nand_x1_sg U50325 ( .A(n40386), .B(n57229), .X(n33556) );
  nand_x1_sg U50326 ( .A(n33537), .B(n33538), .X(n43154) );
  nand_x1_sg U50327 ( .A(n40787), .B(n57229), .X(n33538) );
  nand_x1_sg U50328 ( .A(n33557), .B(n33558), .X(n43164) );
  nand_x1_sg U50329 ( .A(n40352), .B(n57229), .X(n33558) );
  nand_x1_sg U50330 ( .A(n33559), .B(n33560), .X(n43165) );
  nand_x1_sg U50331 ( .A(n40318), .B(n57229), .X(n33560) );
  nand_x1_sg U50332 ( .A(n33543), .B(n33544), .X(n43157) );
  nand_x1_sg U50333 ( .A(n40786), .B(n57229), .X(n33544) );
  nand_x1_sg U50334 ( .A(n33561), .B(n33562), .X(n43166) );
  nand_x1_sg U50335 ( .A(n40284), .B(n57229), .X(n33562) );
  nand_x1_sg U50336 ( .A(n33563), .B(n33564), .X(n43167) );
  nand_x1_sg U50337 ( .A(n40254), .B(n57229), .X(n33564) );
  nand_x1_sg U50338 ( .A(n33565), .B(n33566), .X(n43168) );
  nand_x1_sg U50339 ( .A(n40236), .B(n57229), .X(n33566) );
  nand_x1_sg U50340 ( .A(n34097), .B(n34098), .X(n43412) );
  nand_x1_sg U50341 ( .A(n40808), .B(n57181), .X(n34098) );
  nand_x1_sg U50342 ( .A(n34105), .B(n34106), .X(n43416) );
  nand_x1_sg U50343 ( .A(n40807), .B(n34091), .X(n34106) );
  nand_x1_sg U50344 ( .A(n34089), .B(n34090), .X(n43409) );
  nand_x1_sg U50345 ( .A(n40806), .B(n57181), .X(n34090) );
  nand_x1_sg U50346 ( .A(n34109), .B(n34110), .X(n43418) );
  nand_x1_sg U50347 ( .A(n40805), .B(n57181), .X(n34110) );
  nand_x1_sg U50348 ( .A(n34111), .B(n34112), .X(n43419) );
  nand_x1_sg U50349 ( .A(n40804), .B(n57181), .X(n34112) );
  nand_x1_sg U50350 ( .A(n34103), .B(n34104), .X(n43415) );
  nand_x1_sg U50351 ( .A(n40803), .B(n57181), .X(n34104) );
  nand_x1_sg U50352 ( .A(n34101), .B(n34102), .X(n43414) );
  nand_x1_sg U50353 ( .A(n40802), .B(n57181), .X(n34102) );
  nand_x1_sg U50354 ( .A(n34095), .B(n34096), .X(n43411) );
  nand_x1_sg U50355 ( .A(n40801), .B(n57181), .X(n34096) );
  nand_x1_sg U50356 ( .A(n34113), .B(n34114), .X(n43420) );
  nand_x1_sg U50357 ( .A(n40800), .B(n57181), .X(n34114) );
  nand_x1_sg U50358 ( .A(n34115), .B(n34116), .X(n43421) );
  nand_x1_sg U50359 ( .A(n40480), .B(n57181), .X(n34116) );
  nand_x1_sg U50360 ( .A(n34117), .B(n34118), .X(n43422) );
  nand_x1_sg U50361 ( .A(n40448), .B(n57181), .X(n34118) );
  nand_x1_sg U50362 ( .A(n34119), .B(n34120), .X(n43423) );
  nand_x1_sg U50363 ( .A(n40417), .B(n57181), .X(n34120) );
  nand_x1_sg U50364 ( .A(n34121), .B(n34122), .X(n43424) );
  nand_x1_sg U50365 ( .A(n40385), .B(n57181), .X(n34122) );
  nand_x1_sg U50366 ( .A(n34093), .B(n34094), .X(n43410) );
  nand_x1_sg U50367 ( .A(n40799), .B(n57181), .X(n34094) );
  nand_x1_sg U50368 ( .A(n34123), .B(n34124), .X(n43425) );
  nand_x1_sg U50369 ( .A(n40351), .B(n57181), .X(n34124) );
  nand_x1_sg U50370 ( .A(n34125), .B(n34126), .X(n43426) );
  nand_x1_sg U50371 ( .A(n40317), .B(n57181), .X(n34126) );
  nand_x1_sg U50372 ( .A(n34107), .B(n34108), .X(n43417) );
  nand_x1_sg U50373 ( .A(n40798), .B(n57181), .X(n34108) );
  nand_x1_sg U50374 ( .A(n34099), .B(n34100), .X(n43413) );
  nand_x1_sg U50375 ( .A(n40797), .B(n57181), .X(n34100) );
  nand_x1_sg U50376 ( .A(n34127), .B(n34128), .X(n43427) );
  nand_x1_sg U50377 ( .A(n40283), .B(n57181), .X(n34128) );
  nand_x1_sg U50378 ( .A(n34129), .B(n34130), .X(n43428) );
  nand_x1_sg U50379 ( .A(n40253), .B(n57181), .X(n34130) );
  nand_x1_sg U50380 ( .A(n33080), .B(n33081), .X(n42942) );
  nand_x1_sg U50381 ( .A(n40820), .B(n57272), .X(n33081) );
  nand_x1_sg U50382 ( .A(n33070), .B(n33071), .X(n42937) );
  nand_x1_sg U50383 ( .A(n40819), .B(n33054), .X(n33071) );
  nand_x1_sg U50384 ( .A(n33060), .B(n33061), .X(n42932) );
  nand_x1_sg U50385 ( .A(n40818), .B(n57272), .X(n33061) );
  nand_x1_sg U50386 ( .A(n33078), .B(n33079), .X(n42941) );
  nand_x1_sg U50387 ( .A(n40817), .B(n57272), .X(n33079) );
  nand_x1_sg U50388 ( .A(n33090), .B(n33091), .X(n42947) );
  nand_x1_sg U50389 ( .A(n40816), .B(n57272), .X(n33091) );
  nand_x1_sg U50390 ( .A(n33088), .B(n33089), .X(n42946) );
  nand_x1_sg U50391 ( .A(n40815), .B(n57272), .X(n33089) );
  nand_x1_sg U50392 ( .A(n33056), .B(n33057), .X(n42930) );
  nand_x1_sg U50393 ( .A(n40479), .B(n57272), .X(n33057) );
  nand_x1_sg U50394 ( .A(n33084), .B(n33085), .X(n42944) );
  nand_x1_sg U50395 ( .A(n40447), .B(n57272), .X(n33085) );
  nand_x1_sg U50396 ( .A(n33064), .B(n33065), .X(n42934) );
  nand_x1_sg U50397 ( .A(n40814), .B(n57272), .X(n33065) );
  nand_x1_sg U50398 ( .A(n33086), .B(n33087), .X(n42945) );
  nand_x1_sg U50399 ( .A(n40416), .B(n57272), .X(n33087) );
  nand_x1_sg U50400 ( .A(n33052), .B(n33053), .X(n42929) );
  nand_x1_sg U50401 ( .A(n40813), .B(n57272), .X(n33053) );
  nand_x1_sg U50402 ( .A(n33068), .B(n33069), .X(n42936) );
  nand_x1_sg U50403 ( .A(n40384), .B(n57272), .X(n33069) );
  nand_x1_sg U50404 ( .A(n33062), .B(n33063), .X(n42933) );
  nand_x1_sg U50405 ( .A(n40812), .B(n57272), .X(n33063) );
  nand_x1_sg U50406 ( .A(n33092), .B(n33093), .X(n42948) );
  nand_x1_sg U50407 ( .A(n40350), .B(n57272), .X(n33093) );
  nand_x1_sg U50408 ( .A(n33074), .B(n33075), .X(n42939) );
  nand_x1_sg U50409 ( .A(n40811), .B(n57272), .X(n33075) );
  nand_x1_sg U50410 ( .A(n33082), .B(n33083), .X(n42943) );
  nand_x1_sg U50411 ( .A(n40316), .B(n57272), .X(n33083) );
  nand_x1_sg U50412 ( .A(n33066), .B(n33067), .X(n42935) );
  nand_x1_sg U50413 ( .A(n40810), .B(n57272), .X(n33067) );
  nand_x1_sg U50414 ( .A(n33058), .B(n33059), .X(n42931) );
  nand_x1_sg U50415 ( .A(n40282), .B(n57272), .X(n33059) );
  nand_x1_sg U50416 ( .A(n33076), .B(n33077), .X(n42940) );
  nand_x1_sg U50417 ( .A(n40809), .B(n57272), .X(n33077) );
  nand_x1_sg U50418 ( .A(n33072), .B(n33073), .X(n42938) );
  nand_x1_sg U50419 ( .A(n40252), .B(n57272), .X(n33073) );
  nand_x1_sg U50420 ( .A(n34007), .B(n34008), .X(n43372) );
  nand_x1_sg U50421 ( .A(n40831), .B(n57189), .X(n34008) );
  nand_x1_sg U50422 ( .A(n34015), .B(n34016), .X(n43376) );
  nand_x1_sg U50423 ( .A(n40830), .B(n57189), .X(n34016) );
  nand_x1_sg U50424 ( .A(n33999), .B(n34000), .X(n43369) );
  nand_x1_sg U50425 ( .A(n40829), .B(n57189), .X(n34000) );
  nand_x1_sg U50426 ( .A(n34019), .B(n34020), .X(n43378) );
  nand_x1_sg U50427 ( .A(n40828), .B(n57189), .X(n34020) );
  nand_x1_sg U50428 ( .A(n34021), .B(n34022), .X(n43379) );
  nand_x1_sg U50429 ( .A(n40827), .B(n57189), .X(n34022) );
  nand_x1_sg U50430 ( .A(n34013), .B(n34014), .X(n43375) );
  nand_x1_sg U50431 ( .A(n40826), .B(n57189), .X(n34014) );
  nand_x1_sg U50432 ( .A(n34011), .B(n34012), .X(n43374) );
  nand_x1_sg U50433 ( .A(n40825), .B(n57189), .X(n34012) );
  nand_x1_sg U50434 ( .A(n34005), .B(n34006), .X(n43371) );
  nand_x1_sg U50435 ( .A(n40824), .B(n57189), .X(n34006) );
  nand_x1_sg U50436 ( .A(n34023), .B(n34024), .X(n43380) );
  nand_x1_sg U50437 ( .A(n40478), .B(n57189), .X(n34024) );
  nand_x1_sg U50438 ( .A(n34025), .B(n34026), .X(n43381) );
  nand_x1_sg U50439 ( .A(n40446), .B(n57189), .X(n34026) );
  nand_x1_sg U50440 ( .A(n34027), .B(n34028), .X(n43382) );
  nand_x1_sg U50441 ( .A(n40415), .B(n57189), .X(n34028) );
  nand_x1_sg U50442 ( .A(n34029), .B(n34030), .X(n43383) );
  nand_x1_sg U50443 ( .A(n40383), .B(n57189), .X(n34030) );
  nand_x1_sg U50444 ( .A(n34031), .B(n34032), .X(n43384) );
  nand_x1_sg U50445 ( .A(n40349), .B(n57189), .X(n34032) );
  nand_x1_sg U50446 ( .A(n34003), .B(n34004), .X(n43370) );
  nand_x1_sg U50447 ( .A(n40823), .B(n57189), .X(n34004) );
  nand_x1_sg U50448 ( .A(n34033), .B(n34034), .X(n43385) );
  nand_x1_sg U50449 ( .A(n40315), .B(n57189), .X(n34034) );
  nand_x1_sg U50450 ( .A(n34035), .B(n34036), .X(n43386) );
  nand_x1_sg U50451 ( .A(n40281), .B(n34001), .X(n34036) );
  nand_x1_sg U50452 ( .A(n34017), .B(n34018), .X(n43377) );
  nand_x1_sg U50453 ( .A(n40822), .B(n57189), .X(n34018) );
  nand_x1_sg U50454 ( .A(n34009), .B(n34010), .X(n43373) );
  nand_x1_sg U50455 ( .A(n40821), .B(n57189), .X(n34010) );
  nand_x1_sg U50456 ( .A(n34037), .B(n34038), .X(n43387) );
  nand_x1_sg U50457 ( .A(n40251), .B(n57189), .X(n34038) );
  nand_x1_sg U50458 ( .A(n34039), .B(n34040), .X(n43388) );
  nand_x1_sg U50459 ( .A(n40235), .B(n57189), .X(n34040) );
  nand_x1_sg U50460 ( .A(n34052), .B(n34053), .X(n43392) );
  nand_x1_sg U50461 ( .A(n40842), .B(n57185), .X(n34053) );
  nand_x1_sg U50462 ( .A(n34060), .B(n34061), .X(n43396) );
  nand_x1_sg U50463 ( .A(n40841), .B(n57185), .X(n34061) );
  nand_x1_sg U50464 ( .A(n34044), .B(n34045), .X(n43389) );
  nand_x1_sg U50465 ( .A(n40840), .B(n57185), .X(n34045) );
  nand_x1_sg U50466 ( .A(n34064), .B(n34065), .X(n43398) );
  nand_x1_sg U50467 ( .A(n40839), .B(n57185), .X(n34065) );
  nand_x1_sg U50468 ( .A(n34066), .B(n34067), .X(n43399) );
  nand_x1_sg U50469 ( .A(n40838), .B(n57185), .X(n34067) );
  nand_x1_sg U50470 ( .A(n34058), .B(n34059), .X(n43395) );
  nand_x1_sg U50471 ( .A(n40837), .B(n57185), .X(n34059) );
  nand_x1_sg U50472 ( .A(n34056), .B(n34057), .X(n43394) );
  nand_x1_sg U50473 ( .A(n40836), .B(n57185), .X(n34057) );
  nand_x1_sg U50474 ( .A(n34050), .B(n34051), .X(n43391) );
  nand_x1_sg U50475 ( .A(n40835), .B(n57185), .X(n34051) );
  nand_x1_sg U50476 ( .A(n34068), .B(n34069), .X(n43400) );
  nand_x1_sg U50477 ( .A(n40477), .B(n57185), .X(n34069) );
  nand_x1_sg U50478 ( .A(n34070), .B(n34071), .X(n43401) );
  nand_x1_sg U50479 ( .A(n40445), .B(n57185), .X(n34071) );
  nand_x1_sg U50480 ( .A(n34072), .B(n34073), .X(n43402) );
  nand_x1_sg U50481 ( .A(n40414), .B(n57185), .X(n34073) );
  nand_x1_sg U50482 ( .A(n34074), .B(n34075), .X(n43403) );
  nand_x1_sg U50483 ( .A(n40382), .B(n57185), .X(n34075) );
  nand_x1_sg U50484 ( .A(n34076), .B(n34077), .X(n43404) );
  nand_x1_sg U50485 ( .A(n40348), .B(n57185), .X(n34077) );
  nand_x1_sg U50486 ( .A(n34048), .B(n34049), .X(n43390) );
  nand_x1_sg U50487 ( .A(n40834), .B(n57185), .X(n34049) );
  nand_x1_sg U50488 ( .A(n34078), .B(n34079), .X(n43405) );
  nand_x1_sg U50489 ( .A(n40314), .B(n57185), .X(n34079) );
  nand_x1_sg U50490 ( .A(n34080), .B(n34081), .X(n43406) );
  nand_x1_sg U50491 ( .A(n40280), .B(n34046), .X(n34081) );
  nand_x1_sg U50492 ( .A(n34062), .B(n34063), .X(n43397) );
  nand_x1_sg U50493 ( .A(n40833), .B(n57185), .X(n34063) );
  nand_x1_sg U50494 ( .A(n34054), .B(n34055), .X(n43393) );
  nand_x1_sg U50495 ( .A(n40832), .B(n57185), .X(n34055) );
  nand_x1_sg U50496 ( .A(n34082), .B(n34083), .X(n43407) );
  nand_x1_sg U50497 ( .A(n40250), .B(n57185), .X(n34083) );
  nand_x1_sg U50498 ( .A(n34084), .B(n34085), .X(n43408) );
  nand_x1_sg U50499 ( .A(n40234), .B(n57185), .X(n34085) );
  nand_x1_sg U50500 ( .A(n33921), .B(n33922), .X(n43332) );
  nand_x1_sg U50501 ( .A(n40854), .B(n57197), .X(n33922) );
  nand_x1_sg U50502 ( .A(n33929), .B(n33930), .X(n43336) );
  nand_x1_sg U50503 ( .A(n40853), .B(n57197), .X(n33930) );
  nand_x1_sg U50504 ( .A(n33923), .B(n33924), .X(n43333) );
  nand_x1_sg U50505 ( .A(n40852), .B(n57197), .X(n33924) );
  nand_x1_sg U50506 ( .A(n33933), .B(n33934), .X(n43338) );
  nand_x1_sg U50507 ( .A(n40851), .B(n57197), .X(n33934) );
  nand_x1_sg U50508 ( .A(n33935), .B(n33936), .X(n43339) );
  nand_x1_sg U50509 ( .A(n40850), .B(n57197), .X(n33936) );
  nand_x1_sg U50510 ( .A(n33927), .B(n33928), .X(n43335) );
  nand_x1_sg U50511 ( .A(n40849), .B(n57197), .X(n33928) );
  nand_x1_sg U50512 ( .A(n33913), .B(n33914), .X(n43329) );
  nand_x1_sg U50513 ( .A(n40848), .B(n57197), .X(n33914) );
  nand_x1_sg U50514 ( .A(n33917), .B(n33918), .X(n43330) );
  nand_x1_sg U50515 ( .A(n40847), .B(n57197), .X(n33918) );
  nand_x1_sg U50516 ( .A(n33937), .B(n33938), .X(n43340) );
  nand_x1_sg U50517 ( .A(n40846), .B(n57197), .X(n33938) );
  nand_x1_sg U50518 ( .A(n33939), .B(n33940), .X(n43341) );
  nand_x1_sg U50519 ( .A(n40476), .B(n57197), .X(n33940) );
  nand_x1_sg U50520 ( .A(n33941), .B(n33942), .X(n43342) );
  nand_x1_sg U50521 ( .A(n40444), .B(n57197), .X(n33942) );
  nand_x1_sg U50522 ( .A(n33919), .B(n33920), .X(n43331) );
  nand_x1_sg U50523 ( .A(n40845), .B(n57197), .X(n33920) );
  nand_x1_sg U50524 ( .A(n33943), .B(n33944), .X(n43343) );
  nand_x1_sg U50525 ( .A(n40413), .B(n57197), .X(n33944) );
  nand_x1_sg U50526 ( .A(n33925), .B(n33926), .X(n43334) );
  nand_x1_sg U50527 ( .A(n40844), .B(n57197), .X(n33926) );
  nand_x1_sg U50528 ( .A(n33945), .B(n33946), .X(n43344) );
  nand_x1_sg U50529 ( .A(n40381), .B(n57197), .X(n33946) );
  nand_x1_sg U50530 ( .A(n33947), .B(n33948), .X(n43345) );
  nand_x1_sg U50531 ( .A(n40347), .B(n57197), .X(n33948) );
  nand_x1_sg U50532 ( .A(n33931), .B(n33932), .X(n43337) );
  nand_x1_sg U50533 ( .A(n40843), .B(n33915), .X(n33932) );
  nand_x1_sg U50534 ( .A(n33949), .B(n33950), .X(n43346) );
  nand_x1_sg U50535 ( .A(n40313), .B(n57197), .X(n33950) );
  nand_x1_sg U50536 ( .A(n33951), .B(n33952), .X(n43347) );
  nand_x1_sg U50537 ( .A(n40279), .B(n57197), .X(n33952) );
  nand_x1_sg U50538 ( .A(n33953), .B(n33954), .X(n43348) );
  nand_x1_sg U50539 ( .A(n40249), .B(n57197), .X(n33954) );
  nand_x1_sg U50540 ( .A(n33964), .B(n33965), .X(n43352) );
  nand_x1_sg U50541 ( .A(n40867), .B(n57193), .X(n33965) );
  nand_x1_sg U50542 ( .A(n33972), .B(n33973), .X(n43356) );
  nand_x1_sg U50543 ( .A(n40866), .B(n57193), .X(n33973) );
  nand_x1_sg U50544 ( .A(n33966), .B(n33967), .X(n43353) );
  nand_x1_sg U50545 ( .A(n40865), .B(n57193), .X(n33967) );
  nand_x1_sg U50546 ( .A(n33976), .B(n33977), .X(n43358) );
  nand_x1_sg U50547 ( .A(n40864), .B(n57193), .X(n33977) );
  nand_x1_sg U50548 ( .A(n33978), .B(n33979), .X(n43359) );
  nand_x1_sg U50549 ( .A(n40863), .B(n57193), .X(n33979) );
  nand_x1_sg U50550 ( .A(n33970), .B(n33971), .X(n43355) );
  nand_x1_sg U50551 ( .A(n40862), .B(n57193), .X(n33971) );
  nand_x1_sg U50552 ( .A(n33956), .B(n33957), .X(n43349) );
  nand_x1_sg U50553 ( .A(n40861), .B(n57193), .X(n33957) );
  nand_x1_sg U50554 ( .A(n33960), .B(n33961), .X(n43350) );
  nand_x1_sg U50555 ( .A(n40860), .B(n57193), .X(n33961) );
  nand_x1_sg U50556 ( .A(n33980), .B(n33981), .X(n43360) );
  nand_x1_sg U50557 ( .A(n40859), .B(n57193), .X(n33981) );
  nand_x1_sg U50558 ( .A(n33982), .B(n33983), .X(n43361) );
  nand_x1_sg U50559 ( .A(n40858), .B(n57193), .X(n33983) );
  nand_x1_sg U50560 ( .A(n33984), .B(n33985), .X(n43362) );
  nand_x1_sg U50561 ( .A(n40475), .B(n57193), .X(n33985) );
  nand_x1_sg U50562 ( .A(n33962), .B(n33963), .X(n43351) );
  nand_x1_sg U50563 ( .A(n40857), .B(n57193), .X(n33963) );
  nand_x1_sg U50564 ( .A(n33986), .B(n33987), .X(n43363) );
  nand_x1_sg U50565 ( .A(n40443), .B(n57193), .X(n33987) );
  nand_x1_sg U50566 ( .A(n33968), .B(n33969), .X(n43354) );
  nand_x1_sg U50567 ( .A(n40856), .B(n57193), .X(n33969) );
  nand_x1_sg U50568 ( .A(n33988), .B(n33989), .X(n43364) );
  nand_x1_sg U50569 ( .A(n40412), .B(n57193), .X(n33989) );
  nand_x1_sg U50570 ( .A(n33990), .B(n33991), .X(n43365) );
  nand_x1_sg U50571 ( .A(n40380), .B(n57193), .X(n33991) );
  nand_x1_sg U50572 ( .A(n33974), .B(n33975), .X(n43357) );
  nand_x1_sg U50573 ( .A(n40855), .B(n33958), .X(n33975) );
  nand_x1_sg U50574 ( .A(n33992), .B(n33993), .X(n43366) );
  nand_x1_sg U50575 ( .A(n40346), .B(n57193), .X(n33993) );
  nand_x1_sg U50576 ( .A(n33994), .B(n33995), .X(n43367) );
  nand_x1_sg U50577 ( .A(n40312), .B(n57193), .X(n33995) );
  nand_x1_sg U50578 ( .A(n33996), .B(n33997), .X(n43368) );
  nand_x1_sg U50579 ( .A(n40278), .B(n57193), .X(n33997) );
  nand_x1_sg U50580 ( .A(n39701), .B(n39703), .X(n46195) );
  nand_x1_sg U50581 ( .A(n39697), .B(n39698), .X(n46194) );
  nand_x1_sg U50582 ( .A(n35796), .B(n35797), .X(n44250) );
  nand_x1_sg U50583 ( .A(n35810), .B(n35811), .X(n44257) );
  nand_x1_sg U50584 ( .A(n35802), .B(n35803), .X(n44253) );
  nand_x1_sg U50585 ( .A(n35794), .B(n35795), .X(n44249) );
  nand_x1_sg U50586 ( .A(n35804), .B(n35805), .X(n44254) );
  nand_x1_sg U50587 ( .A(n35806), .B(n35807), .X(n44255) );
  nand_x1_sg U50588 ( .A(n35798), .B(n35799), .X(n44251) );
  nand_x1_sg U50589 ( .A(n35800), .B(n35801), .X(n44252) );
  nand_x1_sg U50590 ( .A(n35782), .B(n35783), .X(n44243) );
  nand_x1_sg U50591 ( .A(n35816), .B(n35817), .X(n44260) );
  nand_x1_sg U50592 ( .A(n35788), .B(n35789), .X(n44246) );
  nand_x1_sg U50593 ( .A(n35780), .B(n35781), .X(n44242) );
  nand_x1_sg U50594 ( .A(n35790), .B(n35791), .X(n44247) );
  nand_x1_sg U50595 ( .A(n35792), .B(n35793), .X(n44248) );
  nand_x1_sg U50596 ( .A(n35784), .B(n35785), .X(n44244) );
  nand_x1_sg U50597 ( .A(n35786), .B(n35787), .X(n44245) );
  nand_x1_sg U50598 ( .A(n35824), .B(n35825), .X(n44264) );
  nand_x1_sg U50599 ( .A(n35808), .B(n35809), .X(n44256) );
  nand_x1_sg U50600 ( .A(n35830), .B(n35831), .X(n44267) );
  nand_x1_sg U50601 ( .A(n35822), .B(n35823), .X(n44263) );
  nand_x1_sg U50602 ( .A(n35832), .B(n35833), .X(n44268) );
  nand_x1_sg U50603 ( .A(n35834), .B(n35835), .X(n44269) );
  nand_x1_sg U50604 ( .A(n35826), .B(n35827), .X(n44265) );
  nand_x1_sg U50605 ( .A(n35828), .B(n35829), .X(n44266) );
  nand_x1_sg U50606 ( .A(n35818), .B(n35819), .X(n44261) );
  nand_x1_sg U50607 ( .A(n35820), .B(n35821), .X(n44262) );
  nand_x1_sg U50608 ( .A(n35812), .B(n35813), .X(n44258) );
  nand_x1_sg U50609 ( .A(n35814), .B(n35815), .X(n44259) );
  nand_x1_sg U50610 ( .A(n35710), .B(n35711), .X(n44207) );
  nand_x1_sg U50611 ( .A(n35716), .B(n35717), .X(n44210) );
  nand_x1_sg U50612 ( .A(n35722), .B(n35723), .X(n44213) );
  nand_x1_sg U50613 ( .A(n35728), .B(n35729), .X(n44216) );
  nand_x1_sg U50614 ( .A(n35736), .B(n35737), .X(n44220) );
  nand_x1_sg U50615 ( .A(n35768), .B(n35769), .X(n44236) );
  nand_x1_sg U50616 ( .A(n35742), .B(n35743), .X(n44223) );
  nand_x1_sg U50617 ( .A(n35734), .B(n35735), .X(n44219) );
  nand_x1_sg U50618 ( .A(n35744), .B(n35745), .X(n44224) );
  nand_x1_sg U50619 ( .A(n35746), .B(n35747), .X(n44225) );
  nand_x1_sg U50620 ( .A(n35738), .B(n35739), .X(n44221) );
  nand_x1_sg U50621 ( .A(n35740), .B(n35741), .X(n44222) );
  nand_x1_sg U50622 ( .A(n35718), .B(n35719), .X(n44211) );
  nand_x1_sg U50623 ( .A(n35720), .B(n35721), .X(n44212) );
  nand_x1_sg U50624 ( .A(n35712), .B(n35713), .X(n44208) );
  nand_x1_sg U50625 ( .A(n35714), .B(n35715), .X(n44209) );
  nand_x1_sg U50626 ( .A(n35730), .B(n35731), .X(n44217) );
  nand_x1_sg U50627 ( .A(n35732), .B(n35733), .X(n44218) );
  nand_x1_sg U50628 ( .A(n35724), .B(n35725), .X(n44214) );
  nand_x1_sg U50629 ( .A(n35726), .B(n35727), .X(n44215) );
  nand_x1_sg U50630 ( .A(n35748), .B(n35749), .X(n44226) );
  nand_x1_sg U50631 ( .A(n35754), .B(n35755), .X(n44229) );
  nand_x1_sg U50632 ( .A(n35774), .B(n35775), .X(n44239) );
  nand_x1_sg U50633 ( .A(n35766), .B(n35767), .X(n44235) );
  nand_x1_sg U50634 ( .A(n35776), .B(n35777), .X(n44240) );
  nand_x1_sg U50635 ( .A(n35778), .B(n35779), .X(n44241) );
  nand_x1_sg U50636 ( .A(n35770), .B(n35771), .X(n44237) );
  nand_x1_sg U50637 ( .A(n35772), .B(n35773), .X(n44238) );
  nand_x1_sg U50638 ( .A(n35756), .B(n35757), .X(n44230) );
  nand_x1_sg U50639 ( .A(n35758), .B(n35759), .X(n44231) );
  nand_x1_sg U50640 ( .A(n35750), .B(n35751), .X(n44227) );
  nand_x1_sg U50641 ( .A(n35752), .B(n35753), .X(n44228) );
  nand_x1_sg U50642 ( .A(n35706), .B(n35707), .X(n44206) );
  nand_x1_sg U50643 ( .A(n35760), .B(n35761), .X(n44232) );
  nand_x1_sg U50644 ( .A(n35762), .B(n35763), .X(n44233) );
  nand_x1_sg U50645 ( .A(n35764), .B(n35765), .X(n44234) );
  nand_x1_sg U50646 ( .A(n35533), .B(n35534), .X(n44119) );
  nand_x1_sg U50647 ( .A(n35526), .B(n35527), .X(n44116) );
  nand_x1_sg U50648 ( .A(n35519), .B(n35520), .X(n44113) );
  nand_x1_sg U50649 ( .A(n35511), .B(n35512), .X(n44110) );
  nand_x1_sg U50650 ( .A(n35699), .B(n35700), .X(n44203) );
  nand_x1_sg U50651 ( .A(n35693), .B(n35694), .X(n44200) );
  nand_x1_sg U50652 ( .A(n35641), .B(n35642), .X(n44170) );
  nand_x1_sg U50653 ( .A(n35635), .B(n35636), .X(n44167) );
  nand_x1_sg U50654 ( .A(n35678), .B(n35679), .X(n44191) );
  nand_x1_sg U50655 ( .A(n35674), .B(n35675), .X(n44188) );
  inv_x1_sg U50656 ( .A(n35607), .X(n68242) );
  nand_x1_sg U50657 ( .A(n35658), .B(n35659), .X(n44179) );
  nand_x1_sg U50658 ( .A(n35652), .B(n35653), .X(n44176) );
  nand_x1_sg U50659 ( .A(n35662), .B(n35663), .X(n44182) );
  nand_x1_sg U50660 ( .A(n35668), .B(n35669), .X(n44185) );
  inv_x1_sg U50661 ( .A(n35595), .X(n68243) );
  nand_x1_sg U50662 ( .A(n35586), .B(n35587), .X(n44143) );
  nand_x1_sg U50663 ( .A(n35682), .B(n35683), .X(n44194) );
  nand_x1_sg U50664 ( .A(n35647), .B(n35648), .X(n44173) );
  nand_x1_sg U50665 ( .A(n35623), .B(n35624), .X(n44161) );
  nand_x1_sg U50666 ( .A(n35599), .B(n35600), .X(n44149) );
  nand_x1_sg U50667 ( .A(n35593), .B(n35594), .X(n44146) );
  nand_x1_sg U50668 ( .A(n35605), .B(n35606), .X(n44152) );
  nand_x1_sg U50669 ( .A(n35611), .B(n35612), .X(n44155) );
  nand_x1_sg U50670 ( .A(n35629), .B(n35630), .X(n44164) );
  nand_x1_sg U50671 ( .A(n35617), .B(n35618), .X(n44158) );
  nand_x1_sg U50672 ( .A(n35580), .B(n35581), .X(n44140) );
  nand_x1_sg U50673 ( .A(n35574), .B(n35575), .X(n44137) );
  nand_x1_sg U50674 ( .A(n35555), .B(n35556), .X(n44128) );
  nand_x1_sg U50675 ( .A(n35547), .B(n35548), .X(n44125) );
  nand_x1_sg U50676 ( .A(n35562), .B(n35563), .X(n44131) );
  nand_x1_sg U50677 ( .A(n35568), .B(n35569), .X(n44134) );
  nand_x1_sg U50678 ( .A(n35688), .B(n35689), .X(n44197) );
  nand_x1_sg U50679 ( .A(n35540), .B(n35541), .X(n44122) );
  nand_x1_sg U50680 ( .A(n35584), .B(n35585), .X(n44142) );
  nand_x1_sg U50681 ( .A(n35582), .B(n35583), .X(n44141) );
  nand_x1_sg U50682 ( .A(n35591), .B(n35592), .X(n44145) );
  nand_x1_sg U50683 ( .A(n35589), .B(n35590), .X(n44144) );
  nand_x1_sg U50684 ( .A(n35603), .B(n35604), .X(n44151) );
  nand_x1_sg U50685 ( .A(n35566), .B(n35567), .X(n44133) );
  nand_x1_sg U50686 ( .A(n35564), .B(n35565), .X(n44132) );
  nand_x1_sg U50687 ( .A(n35550), .B(n35551), .X(n44126) );
  nand_x1_sg U50688 ( .A(n35666), .B(n35667), .X(n44184) );
  nand_x1_sg U50689 ( .A(n35664), .B(n35665), .X(n44183) );
  nand_x1_sg U50690 ( .A(n35672), .B(n35673), .X(n44187) );
  nand_x1_sg U50691 ( .A(n35670), .B(n35671), .X(n44186) );
  nand_x1_sg U50692 ( .A(n35697), .B(n35698), .X(n44202) );
  nand_x1_sg U50693 ( .A(n35695), .B(n35696), .X(n44201) );
  nand_x1_sg U50694 ( .A(n35703), .B(n35704), .X(n44205) );
  nand_x1_sg U50695 ( .A(n35701), .B(n35702), .X(n44204) );
  nand_x1_sg U50696 ( .A(n35686), .B(n35687), .X(n44196) );
  nand_x1_sg U50697 ( .A(n35684), .B(n35685), .X(n44195) );
  nand_x1_sg U50698 ( .A(n35690), .B(n35691), .X(n44198) );
  nand_x1_sg U50699 ( .A(n35633), .B(n35634), .X(n44166) );
  nand_x1_sg U50700 ( .A(n35631), .B(n35632), .X(n44165) );
  nand_x1_sg U50701 ( .A(n35639), .B(n35640), .X(n44169) );
  nand_x1_sg U50702 ( .A(n35637), .B(n35638), .X(n44168) );
  nand_x1_sg U50703 ( .A(n35621), .B(n35622), .X(n44160) );
  nand_x1_sg U50704 ( .A(n35619), .B(n35620), .X(n44159) );
  nand_x1_sg U50705 ( .A(n35627), .B(n35628), .X(n44163) );
  nand_x1_sg U50706 ( .A(n35625), .B(n35626), .X(n44162) );
  nand_x1_sg U50707 ( .A(n35656), .B(n35657), .X(n44178) );
  nand_x1_sg U50708 ( .A(n35654), .B(n35655), .X(n44177) );
  nand_x1_sg U50709 ( .A(n35645), .B(n35646), .X(n44172) );
  nand_x1_sg U50710 ( .A(n35643), .B(n35644), .X(n44171) );
  nand_x1_sg U50711 ( .A(n35650), .B(n35651), .X(n44175) );
  nand_x1_sg U50712 ( .A(n36381), .B(n36382), .X(n44539) );
  nand_x1_sg U50713 ( .A(n38329), .B(n38330), .X(n45513) );
  nand_x1_sg U50714 ( .A(n36389), .B(n36390), .X(n44543) );
  nand_x1_sg U50715 ( .A(n38327), .B(n38328), .X(n45512) );
  nand_x1_sg U50716 ( .A(n36391), .B(n36392), .X(n44544) );
  nand_x1_sg U50717 ( .A(n38319), .B(n38320), .X(n45508) );
  nand_x1_sg U50718 ( .A(n36433), .B(n36434), .X(n44565) );
  nand_x1_sg U50719 ( .A(n38325), .B(n38326), .X(n45511) );
  nand_x1_sg U50720 ( .A(n36435), .B(n36436), .X(n44566) );
  nand_x1_sg U50721 ( .A(n37595), .B(n37596), .X(n45146) );
  nand_x1_sg U50722 ( .A(n36427), .B(n36428), .X(n44562) );
  nand_x1_sg U50723 ( .A(n37597), .B(n37598), .X(n45147) );
  nand_x1_sg U50724 ( .A(n37567), .B(n37568), .X(n45132) );
  nand_x1_sg U50725 ( .A(n38323), .B(n38324), .X(n45510) );
  nand_x1_sg U50726 ( .A(n37549), .B(n37550), .X(n45123) );
  nand_x1_sg U50727 ( .A(n38321), .B(n38322), .X(n45509) );
  nand_x1_sg U50728 ( .A(n37569), .B(n37570), .X(n45133) );
  nand_x1_sg U50729 ( .A(n38331), .B(n38332), .X(n45514) );
  nand_x1_sg U50730 ( .A(n37575), .B(n37576), .X(n45136) );
  nand_x1_sg U50731 ( .A(n37593), .B(n37594), .X(n45145) );
  nand_x1_sg U50732 ( .A(n37577), .B(n37578), .X(n45137) );
  nand_x1_sg U50733 ( .A(n37539), .B(n37540), .X(n45118) );
  nand_x1_sg U50734 ( .A(n37579), .B(n37580), .X(n45138) );
  nand_x1_sg U50735 ( .A(n37541), .B(n37542), .X(n45119) );
  nand_x1_sg U50736 ( .A(n37571), .B(n37572), .X(n45134) );
  nand_x1_sg U50737 ( .A(n37533), .B(n37534), .X(n45115) );
  nand_x1_sg U50738 ( .A(n37573), .B(n37574), .X(n45135) );
  nand_x1_sg U50739 ( .A(n37535), .B(n37536), .X(n45116) );
  nand_x1_sg U50740 ( .A(n37551), .B(n37552), .X(n45124) );
  nand_x1_sg U50741 ( .A(n37529), .B(n37530), .X(n45113) );
  nand_x1_sg U50742 ( .A(n37553), .B(n37554), .X(n45125) );
  nand_x1_sg U50743 ( .A(n37543), .B(n37544), .X(n45120) );
  nand_x1_sg U50744 ( .A(n37545), .B(n37546), .X(n45121) );
  nand_x1_sg U50745 ( .A(n37555), .B(n37556), .X(n45126) );
  nand_x1_sg U50746 ( .A(n37547), .B(n37548), .X(n45122) );
  nand_x1_sg U50747 ( .A(n37561), .B(n37562), .X(n45129) );
  nand_x1_sg U50748 ( .A(n37563), .B(n37564), .X(n45130) );
  nand_x1_sg U50749 ( .A(n37513), .B(n37514), .X(n45105) );
  nand_x1_sg U50750 ( .A(n37565), .B(n37566), .X(n45131) );
  nand_x1_sg U50751 ( .A(n37515), .B(n37516), .X(n45106) );
  nand_x1_sg U50752 ( .A(n37557), .B(n37558), .X(n45127) );
  nand_x1_sg U50753 ( .A(n37507), .B(n37508), .X(n45102) );
  nand_x1_sg U50754 ( .A(n37559), .B(n37560), .X(n45128) );
  nand_x1_sg U50755 ( .A(n37509), .B(n37510), .X(n45103) );
  nand_x1_sg U50756 ( .A(n36637), .B(n36638), .X(n44667) );
  nand_x1_sg U50757 ( .A(n37525), .B(n37526), .X(n45111) );
  nand_x1_sg U50758 ( .A(n36639), .B(n36640), .X(n44668) );
  nand_x1_sg U50759 ( .A(n37527), .B(n37528), .X(n45112) );
  nand_x1_sg U50760 ( .A(n36631), .B(n36632), .X(n44664) );
  nand_x1_sg U50761 ( .A(n37519), .B(n37520), .X(n45108) );
  nand_x1_sg U50762 ( .A(n36633), .B(n36634), .X(n44665) );
  nand_x1_sg U50763 ( .A(n37521), .B(n37522), .X(n45109) );
  nand_x1_sg U50764 ( .A(n36661), .B(n36662), .X(n44679) );
  nand_x1_sg U50765 ( .A(n36649), .B(n36650), .X(n44673) );
  nand_x1_sg U50766 ( .A(n36663), .B(n36664), .X(n44680) );
  nand_x1_sg U50767 ( .A(n36651), .B(n36652), .X(n44674) );
  nand_x1_sg U50768 ( .A(n36655), .B(n36656), .X(n44676) );
  nand_x1_sg U50769 ( .A(n36643), .B(n36644), .X(n44670) );
  nand_x1_sg U50770 ( .A(n36657), .B(n36658), .X(n44677) );
  nand_x1_sg U50771 ( .A(n36645), .B(n36646), .X(n44671) );
  nand_x1_sg U50772 ( .A(n36673), .B(n36674), .X(n44685) );
  nand_x1_sg U50773 ( .A(n36613), .B(n36614), .X(n44655) );
  nand_x1_sg U50774 ( .A(n36675), .B(n36676), .X(n44686) );
  nand_x1_sg U50775 ( .A(n36615), .B(n36616), .X(n44656) );
  nand_x1_sg U50776 ( .A(n36667), .B(n36668), .X(n44682) );
  nand_x1_sg U50777 ( .A(n36607), .B(n36608), .X(n44652) );
  nand_x1_sg U50778 ( .A(n36669), .B(n36670), .X(n44683) );
  nand_x1_sg U50779 ( .A(n36609), .B(n36610), .X(n44653) );
  nand_x1_sg U50780 ( .A(n36589), .B(n36590), .X(n44643) );
  nand_x1_sg U50781 ( .A(n36625), .B(n36626), .X(n44661) );
  nand_x1_sg U50782 ( .A(n36591), .B(n36592), .X(n44644) );
  nand_x1_sg U50783 ( .A(n36627), .B(n36628), .X(n44662) );
  nand_x1_sg U50784 ( .A(n36583), .B(n36584), .X(n44640) );
  nand_x1_sg U50785 ( .A(n36619), .B(n36620), .X(n44658) );
  nand_x1_sg U50786 ( .A(n36585), .B(n36586), .X(n44641) );
  nand_x1_sg U50787 ( .A(n36621), .B(n36622), .X(n44659) );
  nand_x1_sg U50788 ( .A(n36601), .B(n36602), .X(n44649) );
  nand_x1_sg U50789 ( .A(n36685), .B(n36686), .X(n44691) );
  nand_x1_sg U50790 ( .A(n36603), .B(n36604), .X(n44650) );
  nand_x1_sg U50791 ( .A(n36687), .B(n36688), .X(n44692) );
  nand_x1_sg U50792 ( .A(n36595), .B(n36596), .X(n44646) );
  nand_x1_sg U50793 ( .A(n36679), .B(n36680), .X(n44688) );
  nand_x1_sg U50794 ( .A(n36597), .B(n36598), .X(n44647) );
  nand_x1_sg U50795 ( .A(n36681), .B(n36682), .X(n44689) );
  nand_x1_sg U50796 ( .A(n36577), .B(n36578), .X(n44637) );
  nand_x1_sg U50797 ( .A(n36697), .B(n36698), .X(n44697) );
  nand_x1_sg U50798 ( .A(n36579), .B(n36580), .X(n44638) );
  nand_x1_sg U50799 ( .A(n36699), .B(n36700), .X(n44698) );
  nand_x1_sg U50800 ( .A(n36571), .B(n36572), .X(n44634) );
  nand_x1_sg U50801 ( .A(n36691), .B(n36692), .X(n44694) );
  nand_x1_sg U50802 ( .A(n36573), .B(n36574), .X(n44635) );
  nand_x1_sg U50803 ( .A(n36693), .B(n36694), .X(n44695) );
  nand_x1_sg U50804 ( .A(n38147), .B(n38148), .X(n45422) );
  nand_x1_sg U50805 ( .A(n36039), .B(n36040), .X(n44368) );
  nand_x1_sg U50806 ( .A(n37683), .B(n37684), .X(n45190) );
  nand_x1_sg U50807 ( .A(n36041), .B(n36042), .X(n44369) );
  nand_x1_sg U50808 ( .A(n37681), .B(n37682), .X(n45189) );
  nand_x1_sg U50809 ( .A(n38315), .B(n38316), .X(n45506) );
  nand_x1_sg U50810 ( .A(n37673), .B(n37674), .X(n45185) );
  nand_x1_sg U50811 ( .A(n38313), .B(n38314), .X(n45505) );
  nand_x1_sg U50812 ( .A(n37679), .B(n37680), .X(n45188) );
  nand_x1_sg U50813 ( .A(n36565), .B(n36566), .X(n44631) );
  nand_x1_sg U50814 ( .A(n36843), .B(n36844), .X(n44770) );
  nand_x1_sg U50815 ( .A(n36567), .B(n36568), .X(n44632) );
  nand_x1_sg U50816 ( .A(n36835), .B(n36836), .X(n44766) );
  nand_x1_sg U50817 ( .A(n36559), .B(n36560), .X(n44628) );
  nand_x1_sg U50818 ( .A(n36837), .B(n36838), .X(n44767) );
  nand_x1_sg U50819 ( .A(n36561), .B(n36562), .X(n44629) );
  nand_x1_sg U50820 ( .A(n36805), .B(n36806), .X(n44751) );
  nand_x1_sg U50821 ( .A(n36553), .B(n36554), .X(n44625) );
  nand_x1_sg U50822 ( .A(n36807), .B(n36808), .X(n44752) );
  nand_x1_sg U50823 ( .A(n36555), .B(n36556), .X(n44626) );
  nand_x1_sg U50824 ( .A(n36799), .B(n36800), .X(n44748) );
  nand_x1_sg U50825 ( .A(n36547), .B(n36548), .X(n44622) );
  nand_x1_sg U50826 ( .A(n36801), .B(n36802), .X(n44749) );
  nand_x1_sg U50827 ( .A(n36549), .B(n36550), .X(n44623) );
  nand_x1_sg U50828 ( .A(n36817), .B(n36818), .X(n44757) );
  nand_x1_sg U50829 ( .A(n36445), .B(n36446), .X(n44571) );
  nand_x1_sg U50830 ( .A(n36819), .B(n36820), .X(n44758) );
  nand_x1_sg U50831 ( .A(n36447), .B(n36448), .X(n44572) );
  nand_x1_sg U50832 ( .A(n36811), .B(n36812), .X(n44754) );
  nand_x1_sg U50833 ( .A(n36439), .B(n36440), .X(n44568) );
  nand_x1_sg U50834 ( .A(n36813), .B(n36814), .X(n44755) );
  nand_x1_sg U50835 ( .A(n36441), .B(n36442), .X(n44569) );
  nand_x1_sg U50836 ( .A(n36877), .B(n36878), .X(n44787) );
  nand_x1_sg U50837 ( .A(n36457), .B(n36458), .X(n44577) );
  nand_x1_sg U50838 ( .A(n36879), .B(n36880), .X(n44788) );
  nand_x1_sg U50839 ( .A(n36459), .B(n36460), .X(n44578) );
  nand_x1_sg U50840 ( .A(n36871), .B(n36872), .X(n44784) );
  nand_x1_sg U50841 ( .A(n36451), .B(n36452), .X(n44574) );
  nand_x1_sg U50842 ( .A(n36873), .B(n36874), .X(n44785) );
  nand_x1_sg U50843 ( .A(n36453), .B(n36454), .X(n44575) );
  nand_x1_sg U50844 ( .A(n36889), .B(n36890), .X(n44793) );
  nand_x1_sg U50845 ( .A(n36829), .B(n36830), .X(n44763) );
  nand_x1_sg U50846 ( .A(n36891), .B(n36892), .X(n44794) );
  nand_x1_sg U50847 ( .A(n36831), .B(n36832), .X(n44764) );
  nand_x1_sg U50848 ( .A(n36883), .B(n36884), .X(n44790) );
  nand_x1_sg U50849 ( .A(n36823), .B(n36824), .X(n44760) );
  nand_x1_sg U50850 ( .A(n36885), .B(n36886), .X(n44791) );
  nand_x1_sg U50851 ( .A(n36825), .B(n36826), .X(n44761) );
  nand_x1_sg U50852 ( .A(n36853), .B(n36854), .X(n44775) );
  nand_x1_sg U50853 ( .A(n36841), .B(n36842), .X(n44769) );
  nand_x1_sg U50854 ( .A(n36723), .B(n36724), .X(n44710) );
  nand_x1_sg U50855 ( .A(n36855), .B(n36856), .X(n44776) );
  nand_x1_sg U50856 ( .A(n36715), .B(n36716), .X(n44706) );
  nand_x1_sg U50857 ( .A(n36847), .B(n36848), .X(n44772) );
  nand_x1_sg U50858 ( .A(n36717), .B(n36718), .X(n44707) );
  nand_x1_sg U50859 ( .A(n36849), .B(n36850), .X(n44773) );
  nand_x1_sg U50860 ( .A(n36781), .B(n36782), .X(n44739) );
  nand_x1_sg U50861 ( .A(n36865), .B(n36866), .X(n44781) );
  nand_x1_sg U50862 ( .A(n36783), .B(n36784), .X(n44740) );
  nand_x1_sg U50863 ( .A(n36867), .B(n36868), .X(n44782) );
  nand_x1_sg U50864 ( .A(n36775), .B(n36776), .X(n44736) );
  nand_x1_sg U50865 ( .A(n36859), .B(n36860), .X(n44778) );
  nand_x1_sg U50866 ( .A(n36777), .B(n36778), .X(n44737) );
  nand_x1_sg U50867 ( .A(n36861), .B(n36862), .X(n44779) );
  nand_x1_sg U50868 ( .A(n36793), .B(n36794), .X(n44745) );
  nand_x1_sg U50869 ( .A(n36733), .B(n36734), .X(n44715) );
  nand_x1_sg U50870 ( .A(n36795), .B(n36796), .X(n44746) );
  nand_x1_sg U50871 ( .A(n36735), .B(n36736), .X(n44716) );
  nand_x1_sg U50872 ( .A(n36787), .B(n36788), .X(n44742) );
  nand_x1_sg U50873 ( .A(n36727), .B(n36728), .X(n44712) );
  nand_x1_sg U50874 ( .A(n36789), .B(n36790), .X(n44743) );
  nand_x1_sg U50875 ( .A(n36729), .B(n36730), .X(n44713) );
  nand_x1_sg U50876 ( .A(n36757), .B(n36758), .X(n44727) );
  nand_x1_sg U50877 ( .A(n36745), .B(n36746), .X(n44721) );
  nand_x1_sg U50878 ( .A(n36759), .B(n36760), .X(n44728) );
  nand_x1_sg U50879 ( .A(n36747), .B(n36748), .X(n44722) );
  nand_x1_sg U50880 ( .A(n36751), .B(n36752), .X(n44724) );
  nand_x1_sg U50881 ( .A(n36739), .B(n36740), .X(n44718) );
  nand_x1_sg U50882 ( .A(n36753), .B(n36754), .X(n44725) );
  nand_x1_sg U50883 ( .A(n36741), .B(n36742), .X(n44719) );
  nand_x1_sg U50884 ( .A(n36769), .B(n36770), .X(n44733) );
  nand_x1_sg U50885 ( .A(n36709), .B(n36710), .X(n44703) );
  nand_x1_sg U50886 ( .A(n36771), .B(n36772), .X(n44734) );
  nand_x1_sg U50887 ( .A(n36711), .B(n36712), .X(n44704) );
  nand_x1_sg U50888 ( .A(n36763), .B(n36764), .X(n44730) );
  nand_x1_sg U50889 ( .A(n36703), .B(n36704), .X(n44700) );
  nand_x1_sg U50890 ( .A(n36765), .B(n36766), .X(n44731) );
  nand_x1_sg U50891 ( .A(n36705), .B(n36706), .X(n44701) );
  nand_x1_sg U50892 ( .A(n36241), .B(n36242), .X(n44469) );
  nand_x1_sg U50893 ( .A(n36721), .B(n36722), .X(n44709) );
  nand_x1_sg U50894 ( .A(n36349), .B(n36350), .X(n44523) );
  nand_x1_sg U50895 ( .A(n36223), .B(n36224), .X(n44460) );
  nand_x1_sg U50896 ( .A(n36369), .B(n36370), .X(n44533) );
  nand_x1_sg U50897 ( .A(n36243), .B(n36244), .X(n44470) );
  nand_x1_sg U50898 ( .A(n36371), .B(n36372), .X(n44534) );
  nand_x1_sg U50899 ( .A(n36249), .B(n36250), .X(n44473) );
  nand_x1_sg U50900 ( .A(n36263), .B(n36264), .X(n44480) );
  nand_x1_sg U50901 ( .A(n36251), .B(n36252), .X(n44474) );
  nand_x1_sg U50902 ( .A(n36265), .B(n36266), .X(n44481) );
  nand_x1_sg U50903 ( .A(n36253), .B(n36254), .X(n44475) );
  nand_x1_sg U50904 ( .A(n36229), .B(n36230), .X(n44463) );
  nand_x1_sg U50905 ( .A(n36245), .B(n36246), .X(n44471) );
  nand_x1_sg U50906 ( .A(n36235), .B(n36236), .X(n44466) );
  nand_x1_sg U50907 ( .A(n36247), .B(n36248), .X(n44472) );
  nand_x1_sg U50908 ( .A(n36343), .B(n36344), .X(n44520) );
  nand_x1_sg U50909 ( .A(n36225), .B(n36226), .X(n44461) );
  nand_x1_sg U50910 ( .A(n36261), .B(n36262), .X(n44479) );
  nand_x1_sg U50911 ( .A(n36227), .B(n36228), .X(n44462) );
  nand_x1_sg U50912 ( .A(n36345), .B(n36346), .X(n44521) );
  nand_x1_sg U50913 ( .A(n36219), .B(n36220), .X(n44458) );
  nand_x1_sg U50914 ( .A(n36347), .B(n36348), .X(n44522) );
  nand_x1_sg U50915 ( .A(n36221), .B(n36222), .X(n44459) );
  nand_x1_sg U50916 ( .A(n36167), .B(n36168), .X(n44432) );
  nand_x1_sg U50917 ( .A(n36237), .B(n36238), .X(n44467) );
  nand_x1_sg U50918 ( .A(n36173), .B(n36174), .X(n44435) );
  nand_x1_sg U50919 ( .A(n36239), .B(n36240), .X(n44468) );
  nand_x1_sg U50920 ( .A(n36157), .B(n36158), .X(n44427) );
  nand_x1_sg U50921 ( .A(n36231), .B(n36232), .X(n44464) );
  nand_x1_sg U50922 ( .A(n36159), .B(n36160), .X(n44428) );
  nand_x1_sg U50923 ( .A(n36233), .B(n36234), .X(n44465) );
  nand_x1_sg U50924 ( .A(n36151), .B(n36152), .X(n44424) );
  nand_x1_sg U50925 ( .A(n36357), .B(n36358), .X(n44527) );
  nand_x1_sg U50926 ( .A(n36153), .B(n36154), .X(n44425) );
  nand_x1_sg U50927 ( .A(n36359), .B(n36360), .X(n44528) );
  nand_x1_sg U50928 ( .A(n36149), .B(n36150), .X(n44423) );
  nand_x1_sg U50929 ( .A(n36351), .B(n36352), .X(n44524) );
  nand_x1_sg U50930 ( .A(n36155), .B(n36156), .X(n44426) );
  nand_x1_sg U50931 ( .A(n36353), .B(n36354), .X(n44525) );
  nand_x1_sg U50932 ( .A(n36163), .B(n36164), .X(n44430) );
  nand_x1_sg U50933 ( .A(n36367), .B(n36368), .X(n44532) );
  nand_x1_sg U50934 ( .A(n36179), .B(n36180), .X(n44438) );
  nand_x1_sg U50935 ( .A(n36165), .B(n36166), .X(n44431) );
  nand_x1_sg U50936 ( .A(n36199), .B(n36200), .X(n44448) );
  nand_x1_sg U50937 ( .A(n36161), .B(n36162), .X(n44429) );
  nand_x1_sg U50938 ( .A(n36201), .B(n36202), .X(n44449) );
  nand_x1_sg U50939 ( .A(n36117), .B(n36118), .X(n44407) );
  nand_x1_sg U50940 ( .A(n36489), .B(n36490), .X(n44593) );
  nand_x1_sg U50941 ( .A(n36175), .B(n36176), .X(n44436) );
  nand_x1_sg U50942 ( .A(n36491), .B(n36492), .X(n44594) );
  nand_x1_sg U50943 ( .A(n36177), .B(n36178), .X(n44437) );
  nand_x1_sg U50944 ( .A(n36483), .B(n36484), .X(n44590) );
  nand_x1_sg U50945 ( .A(n36169), .B(n36170), .X(n44433) );
  nand_x1_sg U50946 ( .A(n36485), .B(n36486), .X(n44591) );
  nand_x1_sg U50947 ( .A(n36171), .B(n36172), .X(n44434) );
  nand_x1_sg U50948 ( .A(n36501), .B(n36502), .X(n44599) );
  nand_x1_sg U50949 ( .A(n36213), .B(n36214), .X(n44455) );
  nand_x1_sg U50950 ( .A(n36503), .B(n36504), .X(n44600) );
  nand_x1_sg U50951 ( .A(n36215), .B(n36216), .X(n44456) );
  nand_x1_sg U50952 ( .A(n36495), .B(n36496), .X(n44596) );
  nand_x1_sg U50953 ( .A(n36207), .B(n36208), .X(n44452) );
  nand_x1_sg U50954 ( .A(n36497), .B(n36498), .X(n44597) );
  nand_x1_sg U50955 ( .A(n36209), .B(n36210), .X(n44453) );
  nand_x1_sg U50956 ( .A(n36477), .B(n36478), .X(n44587) );
  nand_x1_sg U50957 ( .A(n36211), .B(n36212), .X(n44454) );
  nand_x1_sg U50958 ( .A(n36479), .B(n36480), .X(n44588) );
  nand_x1_sg U50959 ( .A(n36217), .B(n36218), .X(n44457) );
  nand_x1_sg U50960 ( .A(n36471), .B(n36472), .X(n44584) );
  nand_x1_sg U50961 ( .A(n36203), .B(n36204), .X(n44450) );
  nand_x1_sg U50962 ( .A(n36473), .B(n36474), .X(n44585) );
  nand_x1_sg U50963 ( .A(n36205), .B(n36206), .X(n44451) );
  nand_x1_sg U50964 ( .A(n36481), .B(n36482), .X(n44589) );
  nand_x1_sg U50965 ( .A(n36187), .B(n36188), .X(n44442) );
  nand_x1_sg U50966 ( .A(n36469), .B(n36470), .X(n44583) );
  nand_x1_sg U50967 ( .A(n36189), .B(n36190), .X(n44443) );
  nand_x1_sg U50968 ( .A(n36475), .B(n36476), .X(n44586) );
  nand_x1_sg U50969 ( .A(n36181), .B(n36182), .X(n44439) );
  nand_x1_sg U50970 ( .A(n36467), .B(n36468), .X(n44582) );
  nand_x1_sg U50971 ( .A(n36183), .B(n36184), .X(n44440) );
  nand_x1_sg U50972 ( .A(n36529), .B(n36530), .X(n44613) );
  nand_x1_sg U50973 ( .A(n36197), .B(n36198), .X(n44447) );
  nand_x1_sg U50974 ( .A(n36511), .B(n36512), .X(n44604) );
  nand_x1_sg U50975 ( .A(n36531), .B(n36532), .X(n44614) );
  nand_x1_sg U50976 ( .A(n36395), .B(n36396), .X(n44546) );
  nand_x1_sg U50977 ( .A(n36523), .B(n36524), .X(n44610) );
  nand_x1_sg U50978 ( .A(n36397), .B(n36398), .X(n44547) );
  nand_x1_sg U50979 ( .A(n36525), .B(n36526), .X(n44611) );
  nand_x1_sg U50980 ( .A(n36393), .B(n36394), .X(n44545) );
  nand_x1_sg U50981 ( .A(n36527), .B(n36528), .X(n44612) );
  nand_x1_sg U50982 ( .A(n36375), .B(n36376), .X(n44536) );
  nand_x1_sg U50983 ( .A(n36507), .B(n36508), .X(n44602) );
  nand_x1_sg U50984 ( .A(n36407), .B(n36408), .X(n44552) );
  nand_x1_sg U50985 ( .A(n36519), .B(n36520), .X(n44608) );
  nand_x1_sg U50986 ( .A(n36409), .B(n36410), .X(n44553) );
  nand_x1_sg U50987 ( .A(n36521), .B(n36522), .X(n44609) );
  nand_x1_sg U50988 ( .A(n36401), .B(n36402), .X(n44549) );
  nand_x1_sg U50989 ( .A(n36499), .B(n36500), .X(n44598) );
  nand_x1_sg U50990 ( .A(n36403), .B(n36404), .X(n44550) );
  nand_x1_sg U50991 ( .A(n36487), .B(n36488), .X(n44592) );
  nand_x1_sg U50992 ( .A(n36383), .B(n36384), .X(n44540) );
  nand_x1_sg U50993 ( .A(n36505), .B(n36506), .X(n44601) );
  nand_x1_sg U50994 ( .A(n36385), .B(n36386), .X(n44541) );
  nand_x1_sg U50995 ( .A(n36493), .B(n36494), .X(n44595) );
  nand_x1_sg U50996 ( .A(n36377), .B(n36378), .X(n44537) );
  nand_x1_sg U50997 ( .A(n36515), .B(n36516), .X(n44606) );
  nand_x1_sg U50998 ( .A(n36379), .B(n36380), .X(n44538) );
  nand_x1_sg U50999 ( .A(n36517), .B(n36518), .X(n44607) );
  nand_x1_sg U51000 ( .A(n36387), .B(n36388), .X(n44542) );
  nand_x1_sg U51001 ( .A(n36509), .B(n36510), .X(n44603) );
  nand_x1_sg U51002 ( .A(n37043), .B(n37044), .X(n44870) );
  nand_x1_sg U51003 ( .A(n36429), .B(n36430), .X(n44563) );
  nand_x1_sg U51004 ( .A(n37055), .B(n37056), .X(n44876) );
  nand_x1_sg U51005 ( .A(n36461), .B(n36462), .X(n44579) );
  nand_x1_sg U51006 ( .A(n37061), .B(n37062), .X(n44879) );
  nand_x1_sg U51007 ( .A(n36425), .B(n36426), .X(n44561) );
  nand_x1_sg U51008 ( .A(n37403), .B(n37404), .X(n45050) );
  nand_x1_sg U51009 ( .A(n36463), .B(n36464), .X(n44580) );
  nand_x1_sg U51010 ( .A(n35965), .B(n35966), .X(n44331) );
  nand_x1_sg U51011 ( .A(n36465), .B(n36466), .X(n44581) );
  nand_x1_sg U51012 ( .A(n35973), .B(n35974), .X(n44335) );
  nand_x1_sg U51013 ( .A(n36399), .B(n36400), .X(n44548) );
  nand_x1_sg U51014 ( .A(n35961), .B(n35962), .X(n44329) );
  nand_x1_sg U51015 ( .A(n36413), .B(n36414), .X(n44555) );
  nand_x1_sg U51016 ( .A(n35967), .B(n35968), .X(n44332) );
  nand_x1_sg U51017 ( .A(n36419), .B(n36420), .X(n44558) );
  nand_x1_sg U51018 ( .A(n35959), .B(n35960), .X(n44328) );
  nand_x1_sg U51019 ( .A(n36411), .B(n36412), .X(n44554) );
  nand_x1_sg U51020 ( .A(n36021), .B(n36022), .X(n44359) );
  nand_x1_sg U51021 ( .A(n36421), .B(n36422), .X(n44559) );
  nand_x1_sg U51022 ( .A(n36023), .B(n36024), .X(n44360) );
  nand_x1_sg U51023 ( .A(n36423), .B(n36424), .X(n44560) );
  nand_x1_sg U51024 ( .A(n36015), .B(n36016), .X(n44356) );
  nand_x1_sg U51025 ( .A(n36415), .B(n36416), .X(n44556) );
  nand_x1_sg U51026 ( .A(n36017), .B(n36018), .X(n44357) );
  nand_x1_sg U51027 ( .A(n36417), .B(n36418), .X(n44557) );
  nand_x1_sg U51028 ( .A(n36013), .B(n36014), .X(n44355) );
  nand_x1_sg U51029 ( .A(n35981), .B(n35982), .X(n44339) );
  nand_x1_sg U51030 ( .A(n36005), .B(n36006), .X(n44351) );
  nand_x1_sg U51031 ( .A(n35983), .B(n35984), .X(n44340) );
  nand_x1_sg U51032 ( .A(n36011), .B(n36012), .X(n44354) );
  nand_x1_sg U51033 ( .A(n35975), .B(n35976), .X(n44336) );
  nand_x1_sg U51034 ( .A(n35999), .B(n36000), .X(n44348) );
  nand_x1_sg U51035 ( .A(n35977), .B(n35978), .X(n44337) );
  nand_x1_sg U51036 ( .A(n35991), .B(n35992), .X(n44344) );
  nand_x1_sg U51037 ( .A(n35993), .B(n35994), .X(n44345) );
  nand_x1_sg U51038 ( .A(n35979), .B(n35980), .X(n44338) );
  nand_x1_sg U51039 ( .A(n35995), .B(n35996), .X(n44346) );
  nand_x1_sg U51040 ( .A(n35997), .B(n35998), .X(n44347) );
  nand_x1_sg U51041 ( .A(n35987), .B(n35988), .X(n44342) );
  nand_x1_sg U51042 ( .A(n35985), .B(n35986), .X(n44341) );
  nand_x1_sg U51043 ( .A(n35989), .B(n35990), .X(n44343) );
  nand_x1_sg U51044 ( .A(n36007), .B(n36008), .X(n44352) );
  nand_x1_sg U51045 ( .A(n35969), .B(n35970), .X(n44333) );
  nand_x1_sg U51046 ( .A(n36009), .B(n36010), .X(n44353) );
  nand_x1_sg U51047 ( .A(n35971), .B(n35972), .X(n44334) );
  nand_x1_sg U51048 ( .A(n36001), .B(n36002), .X(n44349) );
  nand_x1_sg U51049 ( .A(n35963), .B(n35964), .X(n44330) );
  nand_x1_sg U51050 ( .A(n35939), .B(n35940), .X(n44318) );
  nand_x1_sg U51051 ( .A(n36003), .B(n36004), .X(n44350) );
  nand_x1_sg U51052 ( .A(n35953), .B(n35954), .X(n44325) );
  nand_x1_sg U51053 ( .A(n35905), .B(n35906), .X(n44301) );
  nand_x1_sg U51054 ( .A(n35935), .B(n35936), .X(n44316) );
  nand_x1_sg U51055 ( .A(n35907), .B(n35908), .X(n44302) );
  nand_x1_sg U51056 ( .A(n35955), .B(n35956), .X(n44326) );
  nand_x1_sg U51057 ( .A(n35903), .B(n35904), .X(n44300) );
  nand_x1_sg U51058 ( .A(n35957), .B(n35958), .X(n44327) );
  nand_x1_sg U51059 ( .A(n35891), .B(n35892), .X(n44294) );
  nand_x1_sg U51060 ( .A(n35909), .B(n35910), .X(n44303) );
  nand_x1_sg U51061 ( .A(n35917), .B(n35918), .X(n44307) );
  nand_x1_sg U51062 ( .A(n35923), .B(n35924), .X(n44310) );
  nand_x1_sg U51063 ( .A(n35919), .B(n35920), .X(n44308) );
  nand_x1_sg U51064 ( .A(n35929), .B(n35930), .X(n44313) );
  nand_x1_sg U51065 ( .A(n35911), .B(n35912), .X(n44304) );
  nand_x1_sg U51066 ( .A(n35921), .B(n35922), .X(n44309) );
  nand_x1_sg U51067 ( .A(n35913), .B(n35914), .X(n44305) );
  nand_x1_sg U51068 ( .A(n35931), .B(n35932), .X(n44314) );
  nand_x1_sg U51069 ( .A(n35893), .B(n35894), .X(n44295) );
  nand_x1_sg U51070 ( .A(n35933), .B(n35934), .X(n44315) );
  nand_x1_sg U51071 ( .A(n35895), .B(n35896), .X(n44296) );
  nand_x1_sg U51072 ( .A(n35925), .B(n35926), .X(n44311) );
  nand_x1_sg U51073 ( .A(n35887), .B(n35888), .X(n44292) );
  nand_x1_sg U51074 ( .A(n35927), .B(n35928), .X(n44312) );
  nand_x1_sg U51075 ( .A(n35889), .B(n35890), .X(n44293) );
  nand_x1_sg U51076 ( .A(n36145), .B(n36146), .X(n44421) );
  nand_x1_sg U51077 ( .A(n35897), .B(n35898), .X(n44297) );
  nand_x1_sg U51078 ( .A(n36147), .B(n36148), .X(n44422) );
  nand_x1_sg U51079 ( .A(n35885), .B(n35886), .X(n44291) );
  nand_x1_sg U51080 ( .A(n36139), .B(n36140), .X(n44418) );
  nand_x1_sg U51081 ( .A(n35899), .B(n35900), .X(n44298) );
  nand_x1_sg U51082 ( .A(n36141), .B(n36142), .X(n44419) );
  nand_x1_sg U51083 ( .A(n35901), .B(n35902), .X(n44299) );
  nand_x1_sg U51084 ( .A(n36101), .B(n36102), .X(n44399) );
  nand_x1_sg U51085 ( .A(n35943), .B(n35944), .X(n44320) );
  nand_x1_sg U51086 ( .A(n36137), .B(n36138), .X(n44417) );
  nand_x1_sg U51087 ( .A(n35945), .B(n35946), .X(n44321) );
  nand_x1_sg U51088 ( .A(n36143), .B(n36144), .X(n44420) );
  nand_x1_sg U51089 ( .A(n35937), .B(n35938), .X(n44317) );
  nand_x1_sg U51090 ( .A(n37343), .B(n37344), .X(n45020) );
  nand_x1_sg U51091 ( .A(n36135), .B(n36136), .X(n44416) );
  nand_x1_sg U51092 ( .A(n37355), .B(n37356), .X(n45026) );
  nand_x1_sg U51093 ( .A(n36111), .B(n36112), .X(n44404) );
  nand_x1_sg U51094 ( .A(n37357), .B(n37358), .X(n45027) );
  nand_x1_sg U51095 ( .A(n36113), .B(n36114), .X(n44405) );
  nand_x1_sg U51096 ( .A(n37351), .B(n37352), .X(n45024) );
  nand_x1_sg U51097 ( .A(n36105), .B(n36106), .X(n44401) );
  nand_x1_sg U51098 ( .A(n37353), .B(n37354), .X(n45025) );
  nand_x1_sg U51099 ( .A(n36107), .B(n36108), .X(n44402) );
  nand_x1_sg U51100 ( .A(n36059), .B(n36060), .X(n44378) );
  nand_x1_sg U51101 ( .A(n36131), .B(n36132), .X(n44414) );
  nand_x1_sg U51102 ( .A(n36061), .B(n36062), .X(n44379) );
  nand_x1_sg U51103 ( .A(n36133), .B(n36134), .X(n44415) );
  nand_x1_sg U51104 ( .A(n36053), .B(n36054), .X(n44375) );
  nand_x1_sg U51105 ( .A(n36129), .B(n36130), .X(n44413) );
  nand_x1_sg U51106 ( .A(n36055), .B(n36056), .X(n44376) );
  nand_x1_sg U51107 ( .A(n36103), .B(n36104), .X(n44400) );
  nand_x1_sg U51108 ( .A(n36063), .B(n36064), .X(n44380) );
  nand_x1_sg U51109 ( .A(n35883), .B(n35884), .X(n44290) );
  nand_x1_sg U51110 ( .A(n36051), .B(n36052), .X(n44374) );
  nand_x1_sg U51111 ( .A(n37345), .B(n37346), .X(n45021) );
  nand_x1_sg U51112 ( .A(n36057), .B(n36058), .X(n44377) );
  nand_x1_sg U51113 ( .A(n36115), .B(n36116), .X(n44406) );
  nand_x1_sg U51114 ( .A(n36049), .B(n36050), .X(n44373) );
  nand_x1_sg U51115 ( .A(n37339), .B(n37340), .X(n45018) );
  nand_x1_sg U51116 ( .A(n36033), .B(n36034), .X(n44365) );
  nand_x1_sg U51117 ( .A(n36125), .B(n36126), .X(n44411) );
  nand_x1_sg U51118 ( .A(n36035), .B(n36036), .X(n44366) );
  nand_x1_sg U51119 ( .A(n36127), .B(n36128), .X(n44412) );
  nand_x1_sg U51120 ( .A(n36027), .B(n36028), .X(n44362) );
  nand_x1_sg U51121 ( .A(n36119), .B(n36120), .X(n44408) );
  nand_x1_sg U51122 ( .A(n36029), .B(n36030), .X(n44363) );
  nand_x1_sg U51123 ( .A(n36121), .B(n36122), .X(n44409) );
  nand_x1_sg U51124 ( .A(n36043), .B(n36044), .X(n44370) );
  nand_x1_sg U51125 ( .A(n37347), .B(n37348), .X(n45022) );
  nand_x1_sg U51126 ( .A(n36025), .B(n36026), .X(n44361) );
  nand_x1_sg U51127 ( .A(n37349), .B(n37350), .X(n45023) );
  nand_x1_sg U51128 ( .A(n36045), .B(n36046), .X(n44371) );
  nand_x1_sg U51129 ( .A(n37341), .B(n37342), .X(n45019) );
  nand_x1_sg U51130 ( .A(n37999), .B(n38000), .X(n45348) );
  nand_x1_sg U51131 ( .A(n36047), .B(n36048), .X(n44372) );
  nand_x1_sg U51132 ( .A(n38077), .B(n38078), .X(n45387) );
  nand_x1_sg U51133 ( .A(n36087), .B(n36088), .X(n44392) );
  nand_x1_sg U51134 ( .A(n38075), .B(n38076), .X(n45386) );
  nand_x1_sg U51135 ( .A(n36069), .B(n36070), .X(n44383) );
  nand_x1_sg U51136 ( .A(n37711), .B(n37712), .X(n45204) );
  nand_x1_sg U51137 ( .A(n36089), .B(n36090), .X(n44393) );
  nand_x1_sg U51138 ( .A(n37709), .B(n37710), .X(n45203) );
  nand_x1_sg U51139 ( .A(n36095), .B(n36096), .X(n44396) );
  nand_x1_sg U51140 ( .A(n37715), .B(n37716), .X(n45206) );
  nand_x1_sg U51141 ( .A(n36097), .B(n36098), .X(n44397) );
  nand_x1_sg U51142 ( .A(n37713), .B(n37714), .X(n45205) );
  nand_x1_sg U51143 ( .A(n36099), .B(n36100), .X(n44398) );
  nand_x1_sg U51144 ( .A(n37701), .B(n37702), .X(n45199) );
  nand_x1_sg U51145 ( .A(n36091), .B(n36092), .X(n44394) );
  nand_x1_sg U51146 ( .A(n37699), .B(n37700), .X(n45198) );
  nand_x1_sg U51147 ( .A(n36093), .B(n36094), .X(n44395) );
  nand_x1_sg U51148 ( .A(n37707), .B(n37708), .X(n45202) );
  nand_x1_sg U51149 ( .A(n36071), .B(n36072), .X(n44384) );
  nand_x1_sg U51150 ( .A(n37705), .B(n37706), .X(n45201) );
  nand_x1_sg U51151 ( .A(n36073), .B(n36074), .X(n44385) );
  nand_x1_sg U51152 ( .A(n37723), .B(n37724), .X(n45210) );
  nand_x1_sg U51153 ( .A(n36065), .B(n36066), .X(n44381) );
  nand_x1_sg U51154 ( .A(n37721), .B(n37722), .X(n45209) );
  nand_x1_sg U51155 ( .A(n36067), .B(n36068), .X(n44382) );
  nand_x1_sg U51156 ( .A(n37729), .B(n37730), .X(n45213) );
  nand_x1_sg U51157 ( .A(n36083), .B(n36084), .X(n44390) );
  nand_x1_sg U51158 ( .A(n37727), .B(n37728), .X(n45212) );
  nand_x1_sg U51159 ( .A(n36085), .B(n36086), .X(n44391) );
  nand_x1_sg U51160 ( .A(n37725), .B(n37726), .X(n45211) );
  nand_x1_sg U51161 ( .A(n36077), .B(n36078), .X(n44387) );
  nand_x1_sg U51162 ( .A(n37719), .B(n37720), .X(n45208) );
  nand_x1_sg U51163 ( .A(n36079), .B(n36080), .X(n44388) );
  nand_x1_sg U51164 ( .A(n37703), .B(n37704), .X(n45200) );
  nand_x1_sg U51165 ( .A(n37997), .B(n37998), .X(n45347) );
  nand_x1_sg U51166 ( .A(n37717), .B(n37718), .X(n45207) );
  nand_x1_sg U51167 ( .A(n38073), .B(n38074), .X(n45385) );
  nand_x1_sg U51168 ( .A(n37627), .B(n37628), .X(n45162) );
  nand_x1_sg U51169 ( .A(n38001), .B(n38002), .X(n45349) );
  nand_x1_sg U51170 ( .A(n38129), .B(n38130), .X(n45413) );
  nand_x1_sg U51171 ( .A(n37657), .B(n37658), .X(n45177) );
  nand_x1_sg U51172 ( .A(n37647), .B(n37648), .X(n45172) );
  nand_x1_sg U51173 ( .A(n37613), .B(n37614), .X(n45155) );
  nand_x1_sg U51174 ( .A(n37645), .B(n37646), .X(n45171) );
  nand_x1_sg U51175 ( .A(n37881), .B(n37882), .X(n45289) );
  nand_x1_sg U51176 ( .A(n37649), .B(n37650), .X(n45173) );
  nand_x1_sg U51177 ( .A(n37653), .B(n37654), .X(n45175) );
  nand_x1_sg U51178 ( .A(n38133), .B(n38134), .X(n45415) );
  nand_x1_sg U51179 ( .A(n37655), .B(n37656), .X(n45176) );
  nand_x1_sg U51180 ( .A(n37651), .B(n37652), .X(n45174) );
  nand_x1_sg U51181 ( .A(n38363), .B(n38364), .X(n45530) );
  nand_x1_sg U51182 ( .A(n38131), .B(n38132), .X(n45414) );
  nand_x1_sg U51183 ( .A(n38357), .B(n38358), .X(n45527) );
  nand_x1_sg U51184 ( .A(n38139), .B(n38140), .X(n45418) );
  nand_x1_sg U51185 ( .A(n37659), .B(n37660), .X(n45178) );
  nand_x1_sg U51186 ( .A(n38299), .B(n38300), .X(n45498) );
  nand_x1_sg U51187 ( .A(n37661), .B(n37662), .X(n45179) );
  nand_x1_sg U51188 ( .A(n38281), .B(n38282), .X(n45489) );
  nand_x1_sg U51189 ( .A(n37891), .B(n37892), .X(n45294) );
  nand_x1_sg U51190 ( .A(n38015), .B(n38016), .X(n45356) );
  nand_x1_sg U51191 ( .A(n38401), .B(n38402), .X(n45549) );
  nand_x1_sg U51192 ( .A(n38145), .B(n38146), .X(n45421) );
  nand_x1_sg U51193 ( .A(n38369), .B(n38370), .X(n45533) );
  nand_x1_sg U51194 ( .A(n38303), .B(n38304), .X(n45500) );
  nand_x1_sg U51195 ( .A(n37663), .B(n37664), .X(n45180) );
  nand_x1_sg U51196 ( .A(n38317), .B(n38318), .X(n45507) );
  nand_x1_sg U51197 ( .A(n38383), .B(n38384), .X(n45540) );
  nand_x1_sg U51198 ( .A(n38149), .B(n38150), .X(n45423) );
  nand_x1_sg U51199 ( .A(n37633), .B(n37634), .X(n45165) );
  nand_x1_sg U51200 ( .A(n37227), .B(n37228), .X(n44962) );
  nand_x1_sg U51201 ( .A(n37671), .B(n37672), .X(n45184) );
  nand_x1_sg U51202 ( .A(n37219), .B(n37220), .X(n44958) );
  nand_x1_sg U51203 ( .A(n37669), .B(n37670), .X(n45183) );
  nand_x1_sg U51204 ( .A(n37221), .B(n37222), .X(n44959) );
  nand_x1_sg U51205 ( .A(n37677), .B(n37678), .X(n45187) );
  nand_x1_sg U51206 ( .A(n38345), .B(n38346), .X(n45521) );
  nand_x1_sg U51207 ( .A(n37675), .B(n37676), .X(n45186) );
  nand_x1_sg U51208 ( .A(n38125), .B(n38126), .X(n45411) );
  nand_x1_sg U51209 ( .A(n37693), .B(n37694), .X(n45195) );
  nand_x1_sg U51210 ( .A(n38115), .B(n38116), .X(n45406) );
  nand_x1_sg U51211 ( .A(n37691), .B(n37692), .X(n45194) );
  nand_x1_sg U51212 ( .A(n37825), .B(n37826), .X(n45261) );
  nand_x1_sg U51213 ( .A(n37697), .B(n37698), .X(n45197) );
  nand_x1_sg U51214 ( .A(n38337), .B(n38338), .X(n45517) );
  nand_x1_sg U51215 ( .A(n37695), .B(n37696), .X(n45196) );
  nand_x1_sg U51216 ( .A(n38225), .B(n38226), .X(n45461) );
  nand_x1_sg U51217 ( .A(n37667), .B(n37668), .X(n45182) );
  nand_x1_sg U51218 ( .A(n38223), .B(n38224), .X(n45460) );
  nand_x1_sg U51219 ( .A(n37685), .B(n37686), .X(n45191) );
  nand_x1_sg U51220 ( .A(n38229), .B(n38230), .X(n45463) );
  nand_x1_sg U51221 ( .A(n37689), .B(n37690), .X(n45193) );
  nand_x1_sg U51222 ( .A(n38227), .B(n38228), .X(n45462) );
  nand_x1_sg U51223 ( .A(n37687), .B(n37688), .X(n45192) );
  nand_x1_sg U51224 ( .A(n38217), .B(n38218), .X(n45457) );
  nand_x1_sg U51225 ( .A(n38393), .B(n38394), .X(n45545) );
  nand_x1_sg U51226 ( .A(n38215), .B(n38216), .X(n45456) );
  nand_x1_sg U51227 ( .A(n38107), .B(n38108), .X(n45402) );
  nand_x1_sg U51228 ( .A(n38221), .B(n38222), .X(n45459) );
  nand_x1_sg U51229 ( .A(n37777), .B(n37778), .X(n45237) );
  nand_x1_sg U51230 ( .A(n38219), .B(n38220), .X(n45458) );
  nand_x1_sg U51231 ( .A(n37665), .B(n37666), .X(n45181) );
  nand_x1_sg U51232 ( .A(n38241), .B(n38242), .X(n45469) );
  nand_x1_sg U51233 ( .A(n38143), .B(n38144), .X(n45420) );
  nand_x1_sg U51234 ( .A(n38239), .B(n38240), .X(n45468) );
  nand_x1_sg U51235 ( .A(n38141), .B(n38142), .X(n45419) );
  nand_x1_sg U51236 ( .A(n38245), .B(n38246), .X(n45471) );
  nand_x1_sg U51237 ( .A(n37601), .B(n37602), .X(n45149) );
  nand_x1_sg U51238 ( .A(n38243), .B(n38244), .X(n45470) );
  nand_x1_sg U51239 ( .A(n38105), .B(n38106), .X(n45401) );
  nand_x1_sg U51240 ( .A(n38233), .B(n38234), .X(n45465) );
  nand_x1_sg U51241 ( .A(n38127), .B(n38128), .X(n45412) );
  nand_x1_sg U51242 ( .A(n38231), .B(n38232), .X(n45464) );
  nand_x1_sg U51243 ( .A(n38123), .B(n38124), .X(n45410) );
  nand_x1_sg U51244 ( .A(n38237), .B(n38238), .X(n45467) );
  nand_x1_sg U51245 ( .A(n38343), .B(n38344), .X(n45520) );
  nand_x1_sg U51246 ( .A(n38269), .B(n38270), .X(n45483) );
  nand_x1_sg U51247 ( .A(n38235), .B(n38236), .X(n45466) );
  nand_x1_sg U51248 ( .A(n38259), .B(n38260), .X(n45478) );
  nand_x1_sg U51249 ( .A(n38193), .B(n38194), .X(n45445) );
  nand_x1_sg U51250 ( .A(n38257), .B(n38258), .X(n45477) );
  nand_x1_sg U51251 ( .A(n38191), .B(n38192), .X(n45444) );
  nand_x1_sg U51252 ( .A(n38263), .B(n38264), .X(n45480) );
  nand_x1_sg U51253 ( .A(n38197), .B(n38198), .X(n45447) );
  nand_x1_sg U51254 ( .A(n38261), .B(n38262), .X(n45479) );
  nand_x1_sg U51255 ( .A(n38195), .B(n38196), .X(n45446) );
  nand_x1_sg U51256 ( .A(n38279), .B(n38280), .X(n45488) );
  nand_x1_sg U51257 ( .A(n38185), .B(n38186), .X(n45441) );
  nand_x1_sg U51258 ( .A(n38277), .B(n38278), .X(n45487) );
  nand_x1_sg U51259 ( .A(n38183), .B(n38184), .X(n45440) );
  nand_x1_sg U51260 ( .A(n36755), .B(n36756), .X(n44726) );
  nand_x1_sg U51261 ( .A(n38189), .B(n38190), .X(n45443) );
  nand_x1_sg U51262 ( .A(n36761), .B(n36762), .X(n44729) );
  nand_x1_sg U51263 ( .A(n38187), .B(n38188), .X(n45442) );
  nand_x1_sg U51264 ( .A(n36779), .B(n36780), .X(n44738) );
  nand_x1_sg U51265 ( .A(n38209), .B(n38210), .X(n45453) );
  nand_x1_sg U51266 ( .A(n36767), .B(n36768), .X(n44732) );
  nand_x1_sg U51267 ( .A(n38207), .B(n38208), .X(n45452) );
  nand_x1_sg U51268 ( .A(n36581), .B(n36582), .X(n44639) );
  nand_x1_sg U51269 ( .A(n38213), .B(n38214), .X(n45455) );
  nand_x1_sg U51270 ( .A(n36665), .B(n36666), .X(n44681) );
  nand_x1_sg U51271 ( .A(n38211), .B(n38212), .X(n45454) );
  nand_x1_sg U51272 ( .A(n36671), .B(n36672), .X(n44684) );
  nand_x1_sg U51273 ( .A(n38201), .B(n38202), .X(n45449) );
  nand_x1_sg U51274 ( .A(n36713), .B(n36714), .X(n44705) );
  nand_x1_sg U51275 ( .A(n38199), .B(n38200), .X(n45448) );
  nand_x1_sg U51276 ( .A(n38251), .B(n38252), .X(n45474) );
  nand_x1_sg U51277 ( .A(n38205), .B(n38206), .X(n45451) );
  nand_x1_sg U51278 ( .A(n36851), .B(n36852), .X(n44774) );
  nand_x1_sg U51279 ( .A(n38203), .B(n38204), .X(n45450) );
  nand_x1_sg U51280 ( .A(n36863), .B(n36864), .X(n44780) );
  nand_x1_sg U51281 ( .A(n38267), .B(n38268), .X(n45482) );
  nand_x1_sg U51282 ( .A(n36575), .B(n36576), .X(n44636) );
  nand_x1_sg U51283 ( .A(n38265), .B(n38266), .X(n45481) );
  nand_x1_sg U51284 ( .A(n36791), .B(n36792), .X(n44744) );
  nand_x1_sg U51285 ( .A(n38271), .B(n38272), .X(n45484) );
  nand_x1_sg U51286 ( .A(n36551), .B(n36552), .X(n44624) );
  nand_x1_sg U51287 ( .A(n36797), .B(n36798), .X(n44747) );
  nand_x1_sg U51288 ( .A(n36617), .B(n36618), .X(n44657) );
  nand_x1_sg U51289 ( .A(n38255), .B(n38256), .X(n45476) );
  nand_x1_sg U51290 ( .A(n36605), .B(n36606), .X(n44651) );
  nand_x1_sg U51291 ( .A(n38253), .B(n38254), .X(n45475) );
  nand_x1_sg U51292 ( .A(n36443), .B(n36444), .X(n44570) );
  nand_x1_sg U51293 ( .A(n37139), .B(n37140), .X(n44918) );
  nand_x1_sg U51294 ( .A(n36449), .B(n36450), .X(n44573) );
  nand_x1_sg U51295 ( .A(n37145), .B(n37146), .X(n44921) );
  nand_x1_sg U51296 ( .A(n36455), .B(n36456), .X(n44576) );
  nand_x1_sg U51297 ( .A(n37157), .B(n37158), .X(n44927) );
  nand_x1_sg U51298 ( .A(n36557), .B(n36558), .X(n44627) );
  nand_x1_sg U51299 ( .A(n37163), .B(n37164), .X(n44930) );
  nand_x1_sg U51300 ( .A(n38121), .B(n38122), .X(n45409) );
  nand_x1_sg U51301 ( .A(n35859), .B(n35860), .X(n44278) );
  nand_x1_sg U51302 ( .A(n38119), .B(n38120), .X(n45408) );
  nand_x1_sg U51303 ( .A(n35861), .B(n35862), .X(n44279) );
  nand_x1_sg U51304 ( .A(n36569), .B(n36570), .X(n44633) );
  nand_x1_sg U51305 ( .A(n38137), .B(n38138), .X(n45417) );
  nand_x1_sg U51306 ( .A(n38111), .B(n38112), .X(n45404) );
  nand_x1_sg U51307 ( .A(n38135), .B(n38136), .X(n45416) );
  nand_x1_sg U51308 ( .A(n38113), .B(n38114), .X(n45405) );
  nand_x1_sg U51309 ( .A(n36887), .B(n36888), .X(n44792) );
  nand_x1_sg U51310 ( .A(n36037), .B(n36038), .X(n44367) );
  nand_x1_sg U51311 ( .A(n37007), .B(n37008), .X(n44852) );
  nand_x1_sg U51312 ( .A(n36647), .B(n36648), .X(n44672) );
  nand_x1_sg U51313 ( .A(n37025), .B(n37026), .X(n44861) );
  nand_x1_sg U51314 ( .A(n36677), .B(n36678), .X(n44687) );
  nand_x1_sg U51315 ( .A(n37013), .B(n37014), .X(n44855) );
  nand_x1_sg U51316 ( .A(n36653), .B(n36654), .X(n44675) );
  nand_x1_sg U51317 ( .A(n36815), .B(n36816), .X(n44756) );
  nand_x1_sg U51318 ( .A(n36659), .B(n36660), .X(n44678) );
  nand_x1_sg U51319 ( .A(n36833), .B(n36834), .X(n44765) );
  nand_x1_sg U51320 ( .A(n36689), .B(n36690), .X(n44693) );
  nand_x1_sg U51321 ( .A(n36869), .B(n36870), .X(n44783) );
  nand_x1_sg U51322 ( .A(n36695), .B(n36696), .X(n44696) );
  nand_x1_sg U51323 ( .A(n36875), .B(n36876), .X(n44786) );
  nand_x1_sg U51324 ( .A(n36587), .B(n36588), .X(n44642) );
  nand_x1_sg U51325 ( .A(n36545), .B(n36546), .X(n44621) );
  nand_x1_sg U51326 ( .A(n38155), .B(n38156), .X(n45426) );
  nand_x1_sg U51327 ( .A(n36593), .B(n36594), .X(n44645) );
  nand_x1_sg U51328 ( .A(n38153), .B(n38154), .X(n45425) );
  nand_x1_sg U51329 ( .A(n35873), .B(n35874), .X(n44285) );
  nand_x1_sg U51330 ( .A(n38151), .B(n38152), .X(n45424) );
  nand_x1_sg U51331 ( .A(n36629), .B(n36630), .X(n44663) );
  nand_x1_sg U51332 ( .A(n37315), .B(n37316), .X(n45006) );
  nand_x1_sg U51333 ( .A(n36737), .B(n36738), .X(n44717) );
  nand_x1_sg U51334 ( .A(n37321), .B(n37322), .X(n45009) );
  nand_x1_sg U51335 ( .A(n36743), .B(n36744), .X(n44720) );
  nand_x1_sg U51336 ( .A(n38169), .B(n38170), .X(n45433) );
  nand_x1_sg U51337 ( .A(n36839), .B(n36840), .X(n44768) );
  nand_x1_sg U51338 ( .A(n38167), .B(n38168), .X(n45432) );
  nand_x1_sg U51339 ( .A(n36821), .B(n36822), .X(n44759) );
  nand_x1_sg U51340 ( .A(n38173), .B(n38174), .X(n45435) );
  nand_x1_sg U51341 ( .A(n36701), .B(n36702), .X(n44699) );
  nand_x1_sg U51342 ( .A(n38171), .B(n38172), .X(n45434) );
  nand_x1_sg U51343 ( .A(n36707), .B(n36708), .X(n44702) );
  nand_x1_sg U51344 ( .A(n38161), .B(n38162), .X(n45429) );
  nand_x1_sg U51345 ( .A(n36719), .B(n36720), .X(n44708) );
  nand_x1_sg U51346 ( .A(n38159), .B(n38160), .X(n45428) );
  nand_x1_sg U51347 ( .A(n36725), .B(n36726), .X(n44711) );
  nand_x1_sg U51348 ( .A(n38165), .B(n38166), .X(n45431) );
  nand_x1_sg U51349 ( .A(n36405), .B(n36406), .X(n44551) );
  nand_x1_sg U51350 ( .A(n38163), .B(n38164), .X(n45430) );
  nand_x1_sg U51351 ( .A(n36431), .B(n36432), .X(n44564) );
  nand_x1_sg U51352 ( .A(n38297), .B(n38298), .X(n45497) );
  nand_x1_sg U51353 ( .A(n38179), .B(n38180), .X(n45438) );
  nand_x1_sg U51354 ( .A(n38295), .B(n38296), .X(n45496) );
  nand_x1_sg U51355 ( .A(n38177), .B(n38178), .X(n45437) );
  nand_x1_sg U51356 ( .A(n35855), .B(n35856), .X(n44276) );
  nand_x1_sg U51357 ( .A(n38181), .B(n38182), .X(n45439) );
  nand_x1_sg U51358 ( .A(n35857), .B(n35858), .X(n44277) );
  nand_x1_sg U51359 ( .A(n36267), .B(n36268), .X(n44482) );
  nand_x1_sg U51360 ( .A(n35849), .B(n35850), .X(n44273) );
  nand_x1_sg U51361 ( .A(n35867), .B(n35868), .X(n44282) );
  nand_x1_sg U51362 ( .A(n35851), .B(n35852), .X(n44274) );
  nand_x1_sg U51363 ( .A(n35869), .B(n35870), .X(n44283) );
  nand_x1_sg U51364 ( .A(n37589), .B(n37590), .X(n45143) );
  nand_x1_sg U51365 ( .A(n38157), .B(n38158), .X(n45427) );
  nand_x1_sg U51366 ( .A(n37265), .B(n37266), .X(n44981) );
  nand_x1_sg U51367 ( .A(n37591), .B(n37592), .X(n45144) );
  nand_x1_sg U51368 ( .A(n38293), .B(n38294), .X(n45495) );
  nand_x1_sg U51369 ( .A(n37583), .B(n37584), .X(n45140) );
  nand_x1_sg U51370 ( .A(n37271), .B(n37272), .X(n44984) );
  nand_x1_sg U51371 ( .A(n37585), .B(n37586), .X(n45141) );
  nand_x1_sg U51372 ( .A(n37303), .B(n37304), .X(n45000) );
  nand_x1_sg U51373 ( .A(n37193), .B(n37194), .X(n44945) );
  nand_x1_sg U51374 ( .A(n37309), .B(n37310), .X(n45003) );
  nand_x1_sg U51375 ( .A(n37199), .B(n37200), .X(n44948) );
  nand_x1_sg U51376 ( .A(n36535), .B(n36536), .X(n44616) );
  nand_x1_sg U51377 ( .A(n37235), .B(n37236), .X(n44966) );
  nand_x1_sg U51378 ( .A(n36537), .B(n36538), .X(n44617) );
  nand_x1_sg U51379 ( .A(n37247), .B(n37248), .X(n44972) );
  nand_x1_sg U51380 ( .A(n37211), .B(n37212), .X(n44954) );
  nand_x1_sg U51381 ( .A(n37109), .B(n37110), .X(n44903) );
  nand_x1_sg U51382 ( .A(n37217), .B(n37218), .X(n44957) );
  nand_x1_sg U51383 ( .A(n37115), .B(n37116), .X(n44906) );
  nand_x1_sg U51384 ( .A(n37223), .B(n37224), .X(n44960) );
  nand_x1_sg U51385 ( .A(n37127), .B(n37128), .X(n44912) );
  nand_x1_sg U51386 ( .A(n37241), .B(n37242), .X(n44969) );
  nand_x1_sg U51387 ( .A(n37205), .B(n37206), .X(n44951) );
  nand_x1_sg U51388 ( .A(n37073), .B(n37074), .X(n44885) );
  nand_x1_sg U51389 ( .A(n37175), .B(n37176), .X(n44936) );
  nand_x1_sg U51390 ( .A(n37079), .B(n37080), .X(n44888) );
  nand_x1_sg U51391 ( .A(n37181), .B(n37182), .X(n44939) );
  nand_x1_sg U51392 ( .A(n37091), .B(n37092), .X(n44894) );
  nand_x1_sg U51393 ( .A(n37291), .B(n37292), .X(n44994) );
  nand_x1_sg U51394 ( .A(n37097), .B(n37098), .X(n44897) );
  nand_x1_sg U51395 ( .A(n37297), .B(n37298), .X(n44997) );
  nand_x1_sg U51396 ( .A(n37037), .B(n37038), .X(n44867) );
  nand_x1_sg U51397 ( .A(n37259), .B(n37260), .X(n44978) );
  nand_x1_sg U51398 ( .A(n37031), .B(n37032), .X(n44864) );
  nand_x1_sg U51399 ( .A(n37385), .B(n37386), .X(n45041) );
  nand_x1_sg U51400 ( .A(n36361), .B(n36362), .X(n44529) );
  nand_x1_sg U51401 ( .A(n37405), .B(n37406), .X(n45051) );
  nand_x1_sg U51402 ( .A(n37277), .B(n37278), .X(n44987) );
  nand_x1_sg U51403 ( .A(n37411), .B(n37412), .X(n45054) );
  nand_x1_sg U51404 ( .A(n37421), .B(n37422), .X(n45059) );
  nand_x1_sg U51405 ( .A(n37413), .B(n37414), .X(n45055) );
  nand_x1_sg U51406 ( .A(n37423), .B(n37424), .X(n45060) );
  nand_x1_sg U51407 ( .A(n37415), .B(n37416), .X(n45056) );
  nand_x1_sg U51408 ( .A(n37391), .B(n37392), .X(n45044) );
  nand_x1_sg U51409 ( .A(n37407), .B(n37408), .X(n45052) );
  nand_x1_sg U51410 ( .A(n37397), .B(n37398), .X(n45047) );
  nand_x1_sg U51411 ( .A(n37409), .B(n37410), .X(n45053) );
  nand_x1_sg U51412 ( .A(n37425), .B(n37426), .X(n45061) );
  nand_x1_sg U51413 ( .A(n37387), .B(n37388), .X(n45042) );
  nand_x1_sg U51414 ( .A(n37419), .B(n37420), .X(n45058) );
  nand_x1_sg U51415 ( .A(n37389), .B(n37390), .X(n45043) );
  nand_x1_sg U51416 ( .A(n37427), .B(n37428), .X(n45062) );
  nand_x1_sg U51417 ( .A(n37381), .B(n37382), .X(n45039) );
  nand_x1_sg U51418 ( .A(n37429), .B(n37430), .X(n45063) );
  nand_x1_sg U51419 ( .A(n37383), .B(n37384), .X(n45040) );
  nand_x1_sg U51420 ( .A(n37311), .B(n37312), .X(n45004) );
  nand_x1_sg U51421 ( .A(n37399), .B(n37400), .X(n45048) );
  nand_x1_sg U51422 ( .A(n37313), .B(n37314), .X(n45005) );
  nand_x1_sg U51423 ( .A(n37401), .B(n37402), .X(n45049) );
  nand_x1_sg U51424 ( .A(n37305), .B(n37306), .X(n45001) );
  nand_x1_sg U51425 ( .A(n37393), .B(n37394), .X(n45045) );
  nand_x1_sg U51426 ( .A(n37307), .B(n37308), .X(n45002) );
  nand_x1_sg U51427 ( .A(n37395), .B(n37396), .X(n45046) );
  nand_x1_sg U51428 ( .A(n37323), .B(n37324), .X(n45010) );
  nand_x1_sg U51429 ( .A(n37439), .B(n37440), .X(n45068) );
  nand_x1_sg U51430 ( .A(n37325), .B(n37326), .X(n45011) );
  nand_x1_sg U51431 ( .A(n37441), .B(n37442), .X(n45069) );
  nand_x1_sg U51432 ( .A(n37317), .B(n37318), .X(n45007) );
  nand_x1_sg U51433 ( .A(n37433), .B(n37434), .X(n45065) );
  nand_x1_sg U51434 ( .A(n37319), .B(n37320), .X(n45008) );
  nand_x1_sg U51435 ( .A(n37435), .B(n37436), .X(n45066) );
  nand_x1_sg U51436 ( .A(n37287), .B(n37288), .X(n44992) );
  nand_x1_sg U51437 ( .A(n37417), .B(n37418), .X(n45057) );
  nand_x1_sg U51438 ( .A(n37289), .B(n37290), .X(n44993) );
  nand_x1_sg U51439 ( .A(n37431), .B(n37432), .X(n45064) );
  nand_x1_sg U51440 ( .A(n37281), .B(n37282), .X(n44989) );
  nand_x1_sg U51441 ( .A(n37437), .B(n37438), .X(n45067) );
  nand_x1_sg U51442 ( .A(n37363), .B(n37364), .X(n45030) );
  nand_x1_sg U51443 ( .A(n37283), .B(n37284), .X(n44990) );
  nand_x1_sg U51444 ( .A(n37463), .B(n37464), .X(n45080) );
  nand_x1_sg U51445 ( .A(n37299), .B(n37300), .X(n44998) );
  nand_x1_sg U51446 ( .A(n37465), .B(n37466), .X(n45081) );
  nand_x1_sg U51447 ( .A(n37301), .B(n37302), .X(n44999) );
  nand_x1_sg U51448 ( .A(n37457), .B(n37458), .X(n45077) );
  nand_x1_sg U51449 ( .A(n37293), .B(n37294), .X(n44995) );
  nand_x1_sg U51450 ( .A(n37459), .B(n37460), .X(n45078) );
  nand_x1_sg U51451 ( .A(n37295), .B(n37296), .X(n44996) );
  nand_x1_sg U51452 ( .A(n37475), .B(n37476), .X(n45086) );
  nand_x1_sg U51453 ( .A(n37375), .B(n37376), .X(n45036) );
  nand_x1_sg U51454 ( .A(n37477), .B(n37478), .X(n45087) );
  nand_x1_sg U51455 ( .A(n37377), .B(n37378), .X(n45037) );
  nand_x1_sg U51456 ( .A(n37469), .B(n37470), .X(n45083) );
  nand_x1_sg U51457 ( .A(n37369), .B(n37370), .X(n45033) );
  nand_x1_sg U51458 ( .A(n37471), .B(n37472), .X(n45084) );
  nand_x1_sg U51459 ( .A(n37371), .B(n37372), .X(n45034) );
  nand_x1_sg U51460 ( .A(n37445), .B(n37446), .X(n45071) );
  nand_x1_sg U51461 ( .A(n37373), .B(n37374), .X(n45035) );
  nand_x1_sg U51462 ( .A(n37447), .B(n37448), .X(n45072) );
  nand_x1_sg U51463 ( .A(n37379), .B(n37380), .X(n45038) );
  nand_x1_sg U51464 ( .A(n36333), .B(n36334), .X(n44515) );
  nand_x1_sg U51465 ( .A(n37365), .B(n37366), .X(n45031) );
  nand_x1_sg U51466 ( .A(n36335), .B(n36336), .X(n44516) );
  nand_x1_sg U51467 ( .A(n37367), .B(n37368), .X(n45032) );
  nand_x1_sg U51468 ( .A(n37455), .B(n37456), .X(n45076) );
  nand_x1_sg U51469 ( .A(n37335), .B(n37336), .X(n45016) );
  nand_x1_sg U51470 ( .A(n36331), .B(n36332), .X(n44514) );
  nand_x1_sg U51471 ( .A(n37337), .B(n37338), .X(n45017) );
  nand_x1_sg U51472 ( .A(n37443), .B(n37444), .X(n45070) );
  nand_x1_sg U51473 ( .A(n37329), .B(n37330), .X(n45013) );
  nand_x1_sg U51474 ( .A(n36325), .B(n36326), .X(n44511) );
  nand_x1_sg U51475 ( .A(n37331), .B(n37332), .X(n45014) );
  nand_x1_sg U51476 ( .A(n37501), .B(n37502), .X(n45099) );
  nand_x1_sg U51477 ( .A(n37359), .B(n37360), .X(n45028) );
  nand_x1_sg U51478 ( .A(n37503), .B(n37504), .X(n45100) );
  nand_x1_sg U51479 ( .A(n37333), .B(n37334), .X(n45015) );
  nand_x1_sg U51480 ( .A(n37497), .B(n37498), .X(n45097) );
  nand_x1_sg U51481 ( .A(n37361), .B(n37362), .X(n45029) );
  nand_x1_sg U51482 ( .A(n36297), .B(n36298), .X(n44497) );
  nand_x1_sg U51483 ( .A(n37499), .B(n37500), .X(n45098) );
  nand_x1_sg U51484 ( .A(n36277), .B(n36278), .X(n44487) );
  nand_x1_sg U51485 ( .A(n37487), .B(n37488), .X(n45092) );
  nand_x1_sg U51486 ( .A(n36279), .B(n36280), .X(n44488) );
  nand_x1_sg U51487 ( .A(n37481), .B(n37482), .X(n45089) );
  nand_x1_sg U51488 ( .A(n36271), .B(n36272), .X(n44484) );
  nand_x1_sg U51489 ( .A(n37493), .B(n37494), .X(n45095) );
  nand_x1_sg U51490 ( .A(n36273), .B(n36274), .X(n44485) );
  nand_x1_sg U51491 ( .A(n37495), .B(n37496), .X(n45096) );
  nand_x1_sg U51492 ( .A(n36281), .B(n36282), .X(n44489) );
  nand_x1_sg U51493 ( .A(n37473), .B(n37474), .X(n45085) );
  nand_x1_sg U51494 ( .A(n36275), .B(n36276), .X(n44486) );
  nand_x1_sg U51495 ( .A(n37461), .B(n37462), .X(n45079) );
  nand_x1_sg U51496 ( .A(n36283), .B(n36284), .X(n44490) );
  nand_x1_sg U51497 ( .A(n37479), .B(n37480), .X(n45088) );
  nand_x1_sg U51498 ( .A(n36285), .B(n36286), .X(n44491) );
  nand_x1_sg U51499 ( .A(n37467), .B(n37468), .X(n45082) );
  nand_x1_sg U51500 ( .A(n36327), .B(n36328), .X(n44512) );
  nand_x1_sg U51501 ( .A(n37489), .B(n37490), .X(n45093) );
  nand_x1_sg U51502 ( .A(n36329), .B(n36330), .X(n44513) );
  nand_x1_sg U51503 ( .A(n37491), .B(n37492), .X(n45094) );
  nand_x1_sg U51504 ( .A(n36321), .B(n36322), .X(n44509) );
  nand_x1_sg U51505 ( .A(n37483), .B(n37484), .X(n45090) );
  nand_x1_sg U51506 ( .A(n36323), .B(n36324), .X(n44510) );
  nand_x1_sg U51507 ( .A(n37485), .B(n37486), .X(n45091) );
  nand_x1_sg U51508 ( .A(n36337), .B(n36338), .X(n44517) );
  nand_x1_sg U51509 ( .A(n36289), .B(n36290), .X(n44493) );
  nand_x1_sg U51510 ( .A(n36319), .B(n36320), .X(n44508) );
  nand_x1_sg U51511 ( .A(n36291), .B(n36292), .X(n44494) );
  nand_x1_sg U51512 ( .A(n36339), .B(n36340), .X(n44518) );
  nand_x1_sg U51513 ( .A(n36287), .B(n36288), .X(n44492) );
  nand_x1_sg U51514 ( .A(n36341), .B(n36342), .X(n44519) );
  nand_x1_sg U51515 ( .A(n36269), .B(n36270), .X(n44483) );
  nand_x1_sg U51516 ( .A(n36305), .B(n36306), .X(n44501) );
  nand_x1_sg U51517 ( .A(n36301), .B(n36302), .X(n44499) );
  nand_x1_sg U51518 ( .A(n36293), .B(n36294), .X(n44495) );
  nand_x1_sg U51519 ( .A(n36303), .B(n36304), .X(n44500) );
  nand_x1_sg U51520 ( .A(n36307), .B(n36308), .X(n44502) );
  nand_x1_sg U51521 ( .A(n36295), .B(n36296), .X(n44496) );
  nand_x1_sg U51522 ( .A(n37005), .B(n37006), .X(n44851) );
  nand_x1_sg U51523 ( .A(n36313), .B(n36314), .X(n44505) );
  nand_x1_sg U51524 ( .A(n37069), .B(n37070), .X(n44883) );
  nand_x1_sg U51525 ( .A(n36315), .B(n36316), .X(n44506) );
  nand_x1_sg U51526 ( .A(n37071), .B(n37072), .X(n44884) );
  nand_x1_sg U51527 ( .A(n36317), .B(n36318), .X(n44507) );
  nand_x1_sg U51528 ( .A(n37063), .B(n37064), .X(n44880) );
  nand_x1_sg U51529 ( .A(n36309), .B(n36310), .X(n44503) );
  nand_x1_sg U51530 ( .A(n37065), .B(n37066), .X(n44881) );
  nand_x1_sg U51531 ( .A(n36311), .B(n36312), .X(n44504) );
  nand_x1_sg U51532 ( .A(n37081), .B(n37082), .X(n44889) );
  nand_x1_sg U51533 ( .A(n37021), .B(n37022), .X(n44859) );
  nand_x1_sg U51534 ( .A(n37083), .B(n37084), .X(n44890) );
  nand_x1_sg U51535 ( .A(n37023), .B(n37024), .X(n44860) );
  nand_x1_sg U51536 ( .A(n37075), .B(n37076), .X(n44886) );
  nand_x1_sg U51537 ( .A(n37015), .B(n37016), .X(n44856) );
  nand_x1_sg U51538 ( .A(n37077), .B(n37078), .X(n44887) );
  nand_x1_sg U51539 ( .A(n37017), .B(n37018), .X(n44857) );
  nand_x1_sg U51540 ( .A(n37045), .B(n37046), .X(n44871) );
  nand_x1_sg U51541 ( .A(n37033), .B(n37034), .X(n44865) );
  nand_x1_sg U51542 ( .A(n37047), .B(n37048), .X(n44872) );
  nand_x1_sg U51543 ( .A(n37035), .B(n37036), .X(n44866) );
  nand_x1_sg U51544 ( .A(n37039), .B(n37040), .X(n44868) );
  nand_x1_sg U51545 ( .A(n37027), .B(n37028), .X(n44862) );
  nand_x1_sg U51546 ( .A(n37041), .B(n37042), .X(n44869) );
  nand_x1_sg U51547 ( .A(n37029), .B(n37030), .X(n44863) );
  nand_x1_sg U51548 ( .A(n37057), .B(n37058), .X(n44877) );
  nand_x1_sg U51549 ( .A(n36997), .B(n36998), .X(n44847) );
  nand_x1_sg U51550 ( .A(n37059), .B(n37060), .X(n44878) );
  nand_x1_sg U51551 ( .A(n36999), .B(n37000), .X(n44848) );
  nand_x1_sg U51552 ( .A(n37051), .B(n37052), .X(n44874) );
  nand_x1_sg U51553 ( .A(n36991), .B(n36992), .X(n44844) );
  nand_x1_sg U51554 ( .A(n37053), .B(n37054), .X(n44875) );
  nand_x1_sg U51555 ( .A(n36993), .B(n36994), .X(n44845) );
  nand_x1_sg U51556 ( .A(n36925), .B(n36926), .X(n44811) );
  nand_x1_sg U51557 ( .A(n37009), .B(n37010), .X(n44853) );
  nand_x1_sg U51558 ( .A(n36927), .B(n36928), .X(n44812) );
  nand_x1_sg U51559 ( .A(n37011), .B(n37012), .X(n44854) );
  nand_x1_sg U51560 ( .A(n36919), .B(n36920), .X(n44808) );
  nand_x1_sg U51561 ( .A(n37003), .B(n37004), .X(n44850) );
  nand_x1_sg U51562 ( .A(n36985), .B(n36986), .X(n44841) );
  nand_x1_sg U51563 ( .A(n36921), .B(n36922), .X(n44809) );
  nand_x1_sg U51564 ( .A(n36987), .B(n36988), .X(n44842) );
  nand_x1_sg U51565 ( .A(n36937), .B(n36938), .X(n44817) );
  nand_x1_sg U51566 ( .A(n36979), .B(n36980), .X(n44838) );
  nand_x1_sg U51567 ( .A(n36939), .B(n36940), .X(n44818) );
  nand_x1_sg U51568 ( .A(n36981), .B(n36982), .X(n44839) );
  nand_x1_sg U51569 ( .A(n36931), .B(n36932), .X(n44814) );
  nand_x1_sg U51570 ( .A(n36949), .B(n36950), .X(n44823) );
  nand_x1_sg U51571 ( .A(n36933), .B(n36934), .X(n44815) );
  nand_x1_sg U51572 ( .A(n36951), .B(n36952), .X(n44824) );
  nand_x1_sg U51573 ( .A(n36901), .B(n36902), .X(n44799) );
  nand_x1_sg U51574 ( .A(n36943), .B(n36944), .X(n44820) );
  nand_x1_sg U51575 ( .A(n36903), .B(n36904), .X(n44800) );
  nand_x1_sg U51576 ( .A(n36945), .B(n36946), .X(n44821) );
  nand_x1_sg U51577 ( .A(n36895), .B(n36896), .X(n44796) );
  nand_x1_sg U51578 ( .A(n36961), .B(n36962), .X(n44829) );
  nand_x1_sg U51579 ( .A(n36897), .B(n36898), .X(n44797) );
  nand_x1_sg U51580 ( .A(n36963), .B(n36964), .X(n44830) );
  nand_x1_sg U51581 ( .A(n36913), .B(n36914), .X(n44805) );
  nand_x1_sg U51582 ( .A(n36955), .B(n36956), .X(n44826) );
  nand_x1_sg U51583 ( .A(n36915), .B(n36916), .X(n44806) );
  nand_x1_sg U51584 ( .A(n36957), .B(n36958), .X(n44827) );
  nand_x1_sg U51585 ( .A(n36907), .B(n36908), .X(n44802) );
  nand_x1_sg U51586 ( .A(n37213), .B(n37214), .X(n44955) );
  nand_x1_sg U51587 ( .A(n36909), .B(n36910), .X(n44803) );
  nand_x1_sg U51588 ( .A(n37215), .B(n37216), .X(n44956) );
  nand_x1_sg U51589 ( .A(n36973), .B(n36974), .X(n44835) );
  nand_x1_sg U51590 ( .A(n37207), .B(n37208), .X(n44952) );
  nand_x1_sg U51591 ( .A(n36975), .B(n36976), .X(n44836) );
  nand_x1_sg U51592 ( .A(n37209), .B(n37210), .X(n44953) );
  nand_x1_sg U51593 ( .A(n36967), .B(n36968), .X(n44832) );
  nand_x1_sg U51594 ( .A(n37225), .B(n37226), .X(n44961) );
  nand_x1_sg U51595 ( .A(n36969), .B(n36970), .X(n44833) );
  nand_x1_sg U51596 ( .A(n37607), .B(n37608), .X(n45152) );
  nand_x1_sg U51597 ( .A(n37189), .B(n37190), .X(n44943) );
  nand_x1_sg U51598 ( .A(n37251), .B(n37252), .X(n44974) );
  nand_x1_sg U51599 ( .A(n37191), .B(n37192), .X(n44944) );
  nand_x1_sg U51600 ( .A(n37243), .B(n37244), .X(n44970) );
  nand_x1_sg U51601 ( .A(n37183), .B(n37184), .X(n44940) );
  nand_x1_sg U51602 ( .A(n37245), .B(n37246), .X(n44971) );
  nand_x1_sg U51603 ( .A(n37185), .B(n37186), .X(n44941) );
  nand_x1_sg U51604 ( .A(n37117), .B(n37118), .X(n44907) );
  nand_x1_sg U51605 ( .A(n37201), .B(n37202), .X(n44949) );
  nand_x1_sg U51606 ( .A(n37119), .B(n37120), .X(n44908) );
  nand_x1_sg U51607 ( .A(n37203), .B(n37204), .X(n44950) );
  nand_x1_sg U51608 ( .A(n37111), .B(n37112), .X(n44904) );
  nand_x1_sg U51609 ( .A(n37195), .B(n37196), .X(n44946) );
  nand_x1_sg U51610 ( .A(n37113), .B(n37114), .X(n44905) );
  nand_x1_sg U51611 ( .A(n37197), .B(n37198), .X(n44947) );
  nand_x1_sg U51612 ( .A(n37129), .B(n37130), .X(n44913) );
  nand_x1_sg U51613 ( .A(n37261), .B(n37262), .X(n44979) );
  nand_x1_sg U51614 ( .A(n37131), .B(n37132), .X(n44914) );
  nand_x1_sg U51615 ( .A(n37263), .B(n37264), .X(n44980) );
  nand_x1_sg U51616 ( .A(n37123), .B(n37124), .X(n44910) );
  nand_x1_sg U51617 ( .A(n37255), .B(n37256), .X(n44976) );
  nand_x1_sg U51618 ( .A(n37125), .B(n37126), .X(n44911) );
  nand_x1_sg U51619 ( .A(n37257), .B(n37258), .X(n44977) );
  nand_x1_sg U51620 ( .A(n37093), .B(n37094), .X(n44895) );
  nand_x1_sg U51621 ( .A(n37273), .B(n37274), .X(n44985) );
  nand_x1_sg U51622 ( .A(n37095), .B(n37096), .X(n44896) );
  nand_x1_sg U51623 ( .A(n37275), .B(n37276), .X(n44986) );
  nand_x1_sg U51624 ( .A(n37087), .B(n37088), .X(n44892) );
  nand_x1_sg U51625 ( .A(n37267), .B(n37268), .X(n44982) );
  nand_x1_sg U51626 ( .A(n37089), .B(n37090), .X(n44893) );
  nand_x1_sg U51627 ( .A(n37269), .B(n37270), .X(n44983) );
  nand_x1_sg U51628 ( .A(n37105), .B(n37106), .X(n44901) );
  nand_x1_sg U51629 ( .A(n37237), .B(n37238), .X(n44967) );
  nand_x1_sg U51630 ( .A(n37107), .B(n37108), .X(n44902) );
  nand_x1_sg U51631 ( .A(n37239), .B(n37240), .X(n44968) );
  nand_x1_sg U51632 ( .A(n37099), .B(n37100), .X(n44898) );
  nand_x1_sg U51633 ( .A(n37231), .B(n37232), .X(n44964) );
  nand_x1_sg U51634 ( .A(n37101), .B(n37102), .X(n44899) );
  nand_x1_sg U51635 ( .A(n37233), .B(n37234), .X(n44965) );
  nand_x1_sg U51636 ( .A(n37165), .B(n37166), .X(n44931) );
  nand_x1_sg U51637 ( .A(n37249), .B(n37250), .X(n44973) );
  nand_x1_sg U51638 ( .A(n36959), .B(n36960), .X(n44828) );
  nand_x1_sg U51639 ( .A(n37167), .B(n37168), .X(n44932) );
  nand_x1_sg U51640 ( .A(n38373), .B(n38374), .X(n45535) );
  nand_x1_sg U51641 ( .A(n37159), .B(n37160), .X(n44928) );
  nand_x1_sg U51642 ( .A(n38371), .B(n38372), .X(n45534) );
  nand_x1_sg U51643 ( .A(n37161), .B(n37162), .X(n44929) );
  nand_x1_sg U51644 ( .A(n38375), .B(n38376), .X(n45536) );
  nand_x1_sg U51645 ( .A(n37177), .B(n37178), .X(n44937) );
  nand_x1_sg U51646 ( .A(n36953), .B(n36954), .X(n44825) );
  nand_x1_sg U51647 ( .A(n37179), .B(n37180), .X(n44938) );
  nand_x1_sg U51648 ( .A(n38361), .B(n38362), .X(n45529) );
  nand_x1_sg U51649 ( .A(n37171), .B(n37172), .X(n44934) );
  nand_x1_sg U51650 ( .A(n38359), .B(n38360), .X(n45528) );
  nand_x1_sg U51651 ( .A(n37173), .B(n37174), .X(n44935) );
  nand_x1_sg U51652 ( .A(n38367), .B(n38368), .X(n45532) );
  nand_x1_sg U51653 ( .A(n37141), .B(n37142), .X(n44919) );
  nand_x1_sg U51654 ( .A(n38365), .B(n38366), .X(n45531) );
  nand_x1_sg U51655 ( .A(n37143), .B(n37144), .X(n44920) );
  nand_x1_sg U51656 ( .A(n38387), .B(n38388), .X(n45542) );
  nand_x1_sg U51657 ( .A(n37135), .B(n37136), .X(n44916) );
  nand_x1_sg U51658 ( .A(n38385), .B(n38386), .X(n45541) );
  nand_x1_sg U51659 ( .A(n37137), .B(n37138), .X(n44917) );
  nand_x1_sg U51660 ( .A(n38391), .B(n38392), .X(n45544) );
  nand_x1_sg U51661 ( .A(n37153), .B(n37154), .X(n44925) );
  nand_x1_sg U51662 ( .A(n38389), .B(n38390), .X(n45543) );
  nand_x1_sg U51663 ( .A(n37155), .B(n37156), .X(n44926) );
  nand_x1_sg U51664 ( .A(n38377), .B(n38378), .X(n45537) );
  nand_x1_sg U51665 ( .A(n37147), .B(n37148), .X(n44922) );
  nand_x1_sg U51666 ( .A(n36977), .B(n36978), .X(n44837) );
  nand_x1_sg U51667 ( .A(n37149), .B(n37150), .X(n44923) );
  nand_x1_sg U51668 ( .A(n38381), .B(n38382), .X(n45539) );
  nand_x1_sg U51669 ( .A(n38405), .B(n38406), .X(n45551) );
  nand_x1_sg U51670 ( .A(n38379), .B(n38380), .X(n45538) );
  nand_x1_sg U51671 ( .A(n38403), .B(n38404), .X(n45550) );
  nand_x1_sg U51672 ( .A(n37931), .B(n37932), .X(n45314) );
  nand_x1_sg U51673 ( .A(n38397), .B(n38398), .X(n45547) );
  nand_x1_sg U51674 ( .A(n37919), .B(n37920), .X(n45308) );
  nand_x1_sg U51675 ( .A(n38395), .B(n38396), .X(n45546) );
  nand_x1_sg U51676 ( .A(n37897), .B(n37898), .X(n45297) );
  nand_x1_sg U51677 ( .A(n38399), .B(n38400), .X(n45548) );
  nand_x1_sg U51678 ( .A(n38309), .B(n38310), .X(n45503) );
  nand_x1_sg U51679 ( .A(n37885), .B(n37886), .X(n45291) );
  nand_x1_sg U51680 ( .A(n35941), .B(n35942), .X(n44319) );
  nand_x1_sg U51681 ( .A(n37925), .B(n37926), .X(n45311) );
  nand_x1_sg U51682 ( .A(n37799), .B(n37800), .X(n45248) );
  nand_x1_sg U51683 ( .A(n38347), .B(n38348), .X(n45522) );
  nand_x1_sg U51684 ( .A(n38287), .B(n38288), .X(n45492) );
  nand_x1_sg U51685 ( .A(n37941), .B(n37942), .X(n45319) );
  nand_x1_sg U51686 ( .A(n36923), .B(n36924), .X(n44810) );
  nand_x1_sg U51687 ( .A(n37947), .B(n37948), .X(n45322) );
  nand_x1_sg U51688 ( .A(n35915), .B(n35916), .X(n44306) );
  nand_x1_sg U51689 ( .A(n38275), .B(n38276), .X(n45486) );
  nand_x1_sg U51690 ( .A(n38311), .B(n38312), .X(n45504) );
  nand_x1_sg U51691 ( .A(n38273), .B(n38274), .X(n45485) );
  nand_x1_sg U51692 ( .A(n36941), .B(n36942), .X(n44819) );
  nand_x1_sg U51693 ( .A(n38249), .B(n38250), .X(n45473) );
  nand_x1_sg U51694 ( .A(n36947), .B(n36948), .X(n44822) );
  nand_x1_sg U51695 ( .A(n38247), .B(n38248), .X(n45472) );
  nand_x1_sg U51696 ( .A(n36019), .B(n36020), .X(n44358) );
  nand_x1_sg U51697 ( .A(n38301), .B(n38302), .X(n45499) );
  nand_x1_sg U51698 ( .A(n36109), .B(n36110), .X(n44403) );
  nand_x1_sg U51699 ( .A(n38289), .B(n38290), .X(n45493) );
  nand_x1_sg U51700 ( .A(n38341), .B(n38342), .X(n45519) );
  nand_x1_sg U51701 ( .A(n38283), .B(n38284), .X(n45490) );
  nand_x1_sg U51702 ( .A(n38339), .B(n38340), .X(n45518) );
  nand_x1_sg U51703 ( .A(n38291), .B(n38292), .X(n45494) );
  nand_x1_sg U51704 ( .A(n36075), .B(n36076), .X(n44386) );
  nand_x1_sg U51705 ( .A(n37871), .B(n37872), .X(n45284) );
  nand_x1_sg U51706 ( .A(n37623), .B(n37624), .X(n45160) );
  nand_x1_sg U51707 ( .A(n37603), .B(n37604), .X(n45150) );
  nand_x1_sg U51708 ( .A(n37957), .B(n37958), .X(n45327) );
  nand_x1_sg U51709 ( .A(n37847), .B(n37848), .X(n45272) );
  nand_x1_sg U51710 ( .A(n37625), .B(n37626), .X(n45161) );
  nand_x1_sg U51711 ( .A(n37813), .B(n37814), .X(n45255) );
  nand_x1_sg U51712 ( .A(n36081), .B(n36082), .X(n44389) );
  nand_x1_sg U51713 ( .A(n36123), .B(n36124), .X(n44410) );
  nand_x1_sg U51714 ( .A(n37639), .B(n37640), .X(n45168) );
  nand_x1_sg U51715 ( .A(n37605), .B(n37606), .X(n45151) );
  nand_x1_sg U51716 ( .A(n37643), .B(n37644), .X(n45170) );
  nand_x1_sg U51717 ( .A(n36031), .B(n36032), .X(n44364) );
  nand_x1_sg U51718 ( .A(n38349), .B(n38350), .X(n45523) );
  nand_x1_sg U51719 ( .A(n37641), .B(n37642), .X(n45169) );
  nand_x1_sg U51720 ( .A(n37829), .B(n37830), .X(n45263) );
  nand_x1_sg U51721 ( .A(n37631), .B(n37632), .X(n45164) );
  nand_x1_sg U51722 ( .A(n37827), .B(n37828), .X(n45262) );
  nand_x1_sg U51723 ( .A(n37629), .B(n37630), .X(n45163) );
  nand_x1_sg U51724 ( .A(n37833), .B(n37834), .X(n45265) );
  nand_x1_sg U51725 ( .A(n37637), .B(n37638), .X(n45167) );
  nand_x1_sg U51726 ( .A(n37831), .B(n37832), .X(n45264) );
  nand_x1_sg U51727 ( .A(n37635), .B(n37636), .X(n45166) );
  nand_x1_sg U51728 ( .A(n37821), .B(n37822), .X(n45259) );
  nand_x1_sg U51729 ( .A(n37617), .B(n37618), .X(n45157) );
  nand_x1_sg U51730 ( .A(n37819), .B(n37820), .X(n45258) );
  nand_x1_sg U51731 ( .A(n37615), .B(n37616), .X(n45156) );
  nand_x1_sg U51732 ( .A(n36513), .B(n36514), .X(n44605) );
  nand_x1_sg U51733 ( .A(n37621), .B(n37622), .X(n45159) );
  nand_x1_sg U51734 ( .A(n37823), .B(n37824), .X(n45260) );
  nand_x1_sg U51735 ( .A(n37619), .B(n37620), .X(n45158) );
  nand_x1_sg U51736 ( .A(n36355), .B(n36356), .X(n44526) );
  nand_x1_sg U51737 ( .A(n37753), .B(n37754), .X(n45225) );
  nand_x1_sg U51738 ( .A(n36185), .B(n36186), .X(n44441) );
  nand_x1_sg U51739 ( .A(n38285), .B(n38286), .X(n45491) );
  nand_x1_sg U51740 ( .A(n37845), .B(n37846), .X(n45271) );
  nand_x1_sg U51741 ( .A(n38355), .B(n38356), .X(n45526) );
  nand_x1_sg U51742 ( .A(n37843), .B(n37844), .X(n45270) );
  nand_x1_sg U51743 ( .A(n38353), .B(n38354), .X(n45525) );
  nand_x1_sg U51744 ( .A(n37837), .B(n37838), .X(n45267) );
  nand_x1_sg U51745 ( .A(n37985), .B(n37986), .X(n45341) );
  nand_x1_sg U51746 ( .A(n37835), .B(n37836), .X(n45266) );
  nand_x1_sg U51747 ( .A(n37983), .B(n37984), .X(n45340) );
  nand_x1_sg U51748 ( .A(n37841), .B(n37842), .X(n45269) );
  nand_x1_sg U51749 ( .A(n38335), .B(n38336), .X(n45516) );
  nand_x1_sg U51750 ( .A(n37839), .B(n37840), .X(n45268) );
  nand_x1_sg U51751 ( .A(n38333), .B(n38334), .X(n45515) );
  nand_x1_sg U51752 ( .A(n37793), .B(n37794), .X(n45245) );
  nand_x1_sg U51753 ( .A(n37611), .B(n37612), .X(n45154) );
  nand_x1_sg U51754 ( .A(n37791), .B(n37792), .X(n45244) );
  nand_x1_sg U51755 ( .A(n37609), .B(n37610), .X(n45153) );
  nand_x1_sg U51756 ( .A(n37797), .B(n37798), .X(n45247) );
  nand_x1_sg U51757 ( .A(n38351), .B(n38352), .X(n45524) );
  nand_x1_sg U51758 ( .A(n37863), .B(n37864), .X(n45280) );
  nand_x1_sg U51759 ( .A(n37795), .B(n37796), .X(n45246) );
  nand_x1_sg U51760 ( .A(n37869), .B(n37870), .X(n45283) );
  nand_x1_sg U51761 ( .A(n37785), .B(n37786), .X(n45241) );
  nand_x1_sg U51762 ( .A(n37867), .B(n37868), .X(n45282) );
  nand_x1_sg U51763 ( .A(n37783), .B(n37784), .X(n45240) );
  nand_x1_sg U51764 ( .A(n37889), .B(n37890), .X(n45293) );
  nand_x1_sg U51765 ( .A(n37789), .B(n37790), .X(n45243) );
  nand_x1_sg U51766 ( .A(n37887), .B(n37888), .X(n45292) );
  nand_x1_sg U51767 ( .A(n37787), .B(n37788), .X(n45242) );
  nand_x1_sg U51768 ( .A(n36195), .B(n36196), .X(n44446) );
  nand_x1_sg U51769 ( .A(n37811), .B(n37812), .X(n45254) );
  nand_x1_sg U51770 ( .A(n35863), .B(n35864), .X(n44280) );
  nand_x1_sg U51771 ( .A(n37809), .B(n37810), .X(n45253) );
  nand_x1_sg U51772 ( .A(n36191), .B(n36192), .X(n44444) );
  nand_x1_sg U51773 ( .A(n37817), .B(n37818), .X(n45257) );
  nand_x1_sg U51774 ( .A(n37883), .B(n37884), .X(n45290) );
  nand_x1_sg U51775 ( .A(n37815), .B(n37816), .X(n45256) );
  nand_x1_sg U51776 ( .A(n36373), .B(n36374), .X(n44535) );
  nand_x1_sg U51777 ( .A(n37803), .B(n37804), .X(n45250) );
  nand_x1_sg U51778 ( .A(n37581), .B(n37582), .X(n45139) );
  nand_x1_sg U51779 ( .A(n37801), .B(n37802), .X(n45249) );
  nand_x1_sg U51780 ( .A(n36193), .B(n36194), .X(n44445) );
  nand_x1_sg U51781 ( .A(n37807), .B(n37808), .X(n45252) );
  nand_x1_sg U51782 ( .A(n37587), .B(n37588), .X(n45142) );
  nand_x1_sg U51783 ( .A(n37805), .B(n37806), .X(n45251) );
  nand_x1_sg U51784 ( .A(n37133), .B(n37134), .X(n44915) );
  nand_x1_sg U51785 ( .A(n37875), .B(n37876), .X(n45286) );
  nand_x1_sg U51786 ( .A(n37849), .B(n37850), .X(n45273) );
  nand_x1_sg U51787 ( .A(n37873), .B(n37874), .X(n45285) );
  nand_x1_sg U51788 ( .A(n37169), .B(n37170), .X(n44933) );
  nand_x1_sg U51789 ( .A(n37879), .B(n37880), .X(n45288) );
  nand_x1_sg U51790 ( .A(n37253), .B(n37254), .X(n44975) );
  nand_x1_sg U51791 ( .A(n37877), .B(n37878), .X(n45287) );
  nand_x1_sg U51792 ( .A(n37151), .B(n37152), .X(n44924) );
  nand_x1_sg U51793 ( .A(n37865), .B(n37866), .X(n45281) );
  nand_x1_sg U51794 ( .A(n36541), .B(n36542), .X(n44619) );
  nand_x1_sg U51795 ( .A(n36363), .B(n36364), .X(n44530) );
  nand_x1_sg U51796 ( .A(n36809), .B(n36810), .X(n44753) );
  nand_x1_sg U51797 ( .A(n37861), .B(n37862), .X(n45279) );
  nand_x1_sg U51798 ( .A(n36803), .B(n36804), .X(n44750) );
  nand_x1_sg U51799 ( .A(n37859), .B(n37860), .X(n45278) );
  nand_x1_sg U51800 ( .A(n36543), .B(n36544), .X(n44620) );
  nand_x1_sg U51801 ( .A(n37853), .B(n37854), .X(n45275) );
  nand_x1_sg U51802 ( .A(n37735), .B(n37736), .X(n45216) );
  nand_x1_sg U51803 ( .A(n37851), .B(n37852), .X(n45274) );
  nand_x1_sg U51804 ( .A(n36899), .B(n36900), .X(n44798) );
  nand_x1_sg U51805 ( .A(n37857), .B(n37858), .X(n45277) );
  nand_x1_sg U51806 ( .A(n36911), .B(n36912), .X(n44804) );
  nand_x1_sg U51807 ( .A(n37855), .B(n37856), .X(n45276) );
  nand_x1_sg U51808 ( .A(n36893), .B(n36894), .X(n44795) );
  nand_x1_sg U51809 ( .A(n37749), .B(n37750), .X(n45223) );
  nand_x1_sg U51810 ( .A(n37085), .B(n37086), .X(n44891) );
  nand_x1_sg U51811 ( .A(n37747), .B(n37748), .X(n45222) );
  nand_x1_sg U51812 ( .A(n37733), .B(n37734), .X(n45215) );
  nand_x1_sg U51813 ( .A(n37187), .B(n37188), .X(n44942) );
  nand_x1_sg U51814 ( .A(n37731), .B(n37732), .X(n45214) );
  nand_x1_sg U51815 ( .A(n37121), .B(n37122), .X(n44909) );
  nand_x1_sg U51816 ( .A(n36539), .B(n36540), .X(n44618) );
  nand_x1_sg U51817 ( .A(n37743), .B(n37744), .X(n45220) );
  nand_x1_sg U51818 ( .A(n37739), .B(n37740), .X(n45218) );
  nand_x1_sg U51819 ( .A(n37741), .B(n37742), .X(n45219) );
  nand_x1_sg U51820 ( .A(n35951), .B(n35952), .X(n44324) );
  nand_x1_sg U51821 ( .A(n37229), .B(n37230), .X(n44963) );
  nand_x1_sg U51822 ( .A(n36365), .B(n36366), .X(n44531) );
  nand_x1_sg U51823 ( .A(n37745), .B(n37746), .X(n45221) );
  nand_x1_sg U51824 ( .A(n35949), .B(n35950), .X(n44323) );
  nand_x1_sg U51825 ( .A(n37103), .B(n37104), .X(n44900) );
  nand_x1_sg U51826 ( .A(n35947), .B(n35948), .X(n44322) );
  nand_x1_sg U51827 ( .A(n35865), .B(n35866), .X(n44281) );
  nand_x1_sg U51828 ( .A(n37737), .B(n37738), .X(n45217) );
  nand_x1_sg U51829 ( .A(n37751), .B(n37752), .X(n45224) );
  nand_x1_sg U51830 ( .A(n37279), .B(n37280), .X(n44988) );
  nand_x1_sg U51831 ( .A(n36599), .B(n36600), .X(n44648) );
  nand_x1_sg U51832 ( .A(n36881), .B(n36882), .X(n44789) );
  nand_x1_sg U51833 ( .A(n37067), .B(n37068), .X(n44882) );
  nand_x1_sg U51834 ( .A(n37755), .B(n37756), .X(n45226) );
  nand_x1_sg U51835 ( .A(n37019), .B(n37020), .X(n44858) );
  nand_x1_sg U51836 ( .A(n35877), .B(n35878), .X(n44287) );
  nand_x1_sg U51837 ( .A(n36929), .B(n36930), .X(n44813) );
  nand_x1_sg U51838 ( .A(n37285), .B(n37286), .X(n44991) );
  nand_x1_sg U51839 ( .A(n36965), .B(n36966), .X(n44831) );
  nand_x1_sg U51840 ( .A(n36533), .B(n36534), .X(n44615) );
  nand_x1_sg U51841 ( .A(n36845), .B(n36846), .X(n44771) );
  nand_x1_sg U51842 ( .A(n37769), .B(n37770), .X(n45233) );
  nand_x1_sg U51843 ( .A(n35875), .B(n35876), .X(n44286) );
  nand_x1_sg U51844 ( .A(n37773), .B(n37774), .X(n45235) );
  nand_x1_sg U51845 ( .A(n36827), .B(n36828), .X(n44762) );
  nand_x1_sg U51846 ( .A(n37771), .B(n37772), .X(n45234) );
  nand_x1_sg U51847 ( .A(n36563), .B(n36564), .X(n44630) );
  nand_x1_sg U51848 ( .A(n37763), .B(n37764), .X(n45230) );
  nand_x1_sg U51849 ( .A(n35871), .B(n35872), .X(n44284) );
  nand_x1_sg U51850 ( .A(n37761), .B(n37762), .X(n45229) );
  nand_x1_sg U51851 ( .A(n36731), .B(n36732), .X(n44714) );
  nand_x1_sg U51852 ( .A(n37767), .B(n37768), .X(n45232) );
  nand_x1_sg U51853 ( .A(n37781), .B(n37782), .X(n45239) );
  nand_x1_sg U51854 ( .A(n37765), .B(n37766), .X(n45231) );
  nand_x1_sg U51855 ( .A(n37779), .B(n37780), .X(n45238) );
  nand_x1_sg U51856 ( .A(n38037), .B(n38038), .X(n45367) );
  nand_x1_sg U51857 ( .A(n35879), .B(n35880), .X(n44288) );
  nand_x1_sg U51858 ( .A(n38035), .B(n38036), .X(n45366) );
  nand_x1_sg U51859 ( .A(n37775), .B(n37776), .X(n45236) );
  nand_x1_sg U51860 ( .A(n35845), .B(n35846), .X(n44272) );
  nand_x1_sg U51861 ( .A(n36995), .B(n36996), .X(n44846) );
  nand_x1_sg U51862 ( .A(n38041), .B(n38042), .X(n45369) );
  nand_x1_sg U51863 ( .A(n37001), .B(n37002), .X(n44849) );
  nand_x1_sg U51864 ( .A(n38025), .B(n38026), .X(n45361) );
  nand_x1_sg U51865 ( .A(n35881), .B(n35882), .X(n44289) );
  nand_x1_sg U51866 ( .A(n38023), .B(n38024), .X(n45360) );
  nand_x1_sg U51867 ( .A(n37759), .B(n37760), .X(n45228) );
  nand_x1_sg U51868 ( .A(n38031), .B(n38032), .X(n45364) );
  nand_x1_sg U51869 ( .A(n35853), .B(n35854), .X(n44275) );
  nand_x1_sg U51870 ( .A(n38029), .B(n38030), .X(n45363) );
  nand_x1_sg U51871 ( .A(n37327), .B(n37328), .X(n45012) );
  nand_x1_sg U51872 ( .A(n38047), .B(n38048), .X(n45372) );
  nand_x1_sg U51873 ( .A(n37757), .B(n37758), .X(n45227) );
  nand_x1_sg U51874 ( .A(n36917), .B(n36918), .X(n44807) );
  nand_x1_sg U51875 ( .A(n38045), .B(n38046), .X(n45371) );
  nand_x1_sg U51876 ( .A(n38013), .B(n38014), .X(n45355) );
  nand_x1_sg U51877 ( .A(n38053), .B(n38054), .X(n45375) );
  nand_x1_sg U51878 ( .A(n38011), .B(n38012), .X(n45354) );
  nand_x1_sg U51879 ( .A(n38051), .B(n38052), .X(n45374) );
  nand_x1_sg U51880 ( .A(n38095), .B(n38096), .X(n45396) );
  nand_x1_sg U51881 ( .A(n38043), .B(n38044), .X(n45370) );
  nand_x1_sg U51882 ( .A(n36935), .B(n36936), .X(n44816) );
  nand_x1_sg U51883 ( .A(n38033), .B(n38034), .X(n45365) );
  nand_x1_sg U51884 ( .A(n38089), .B(n38090), .X(n45393) );
  nand_x1_sg U51885 ( .A(n38027), .B(n38028), .X(n45362) );
  nand_x1_sg U51886 ( .A(n38093), .B(n38094), .X(n45395) );
  nand_x1_sg U51887 ( .A(n38039), .B(n38040), .X(n45368) );
  nand_x1_sg U51888 ( .A(n38087), .B(n38088), .X(n45392) );
  nand_x1_sg U51889 ( .A(n38007), .B(n38008), .X(n45352) );
  nand_x1_sg U51890 ( .A(n36971), .B(n36972), .X(n44834) );
  nand_x1_sg U51891 ( .A(n38005), .B(n38006), .X(n45351) );
  nand_x1_sg U51892 ( .A(n36989), .B(n36990), .X(n44843) );
  nand_x1_sg U51893 ( .A(n38003), .B(n38004), .X(n45350) );
  nand_x1_sg U51894 ( .A(n38091), .B(n38092), .X(n45394) );
  nand_x1_sg U51895 ( .A(n37599), .B(n37600), .X(n45148) );
  nand_x1_sg U51896 ( .A(n36983), .B(n36984), .X(n44840) );
  nand_x1_sg U51897 ( .A(n37991), .B(n37992), .X(n45344) );
  nand_x1_sg U51898 ( .A(n37049), .B(n37050), .X(n44873) );
  nand_x1_sg U51899 ( .A(n37989), .B(n37990), .X(n45343) );
  nand_x1_sg U51900 ( .A(n38103), .B(n38104), .X(n45400) );
  nand_x1_sg U51901 ( .A(n37995), .B(n37996), .X(n45346) );
  nand_x1_sg U51902 ( .A(n38101), .B(n38102), .X(n45399) );
  nand_x1_sg U51903 ( .A(n37993), .B(n37994), .X(n45345) );
  nand_x1_sg U51904 ( .A(n38085), .B(n38086), .X(n45391) );
  nand_x1_sg U51905 ( .A(n38021), .B(n38022), .X(n45359) );
  nand_x1_sg U51906 ( .A(n38099), .B(n38100), .X(n45398) );
  nand_x1_sg U51907 ( .A(n38019), .B(n38020), .X(n45358) );
  nand_x1_sg U51908 ( .A(n38097), .B(n38098), .X(n45397) );
  nand_x1_sg U51909 ( .A(n38009), .B(n38010), .X(n45353) );
  nand_x1_sg U51910 ( .A(n38083), .B(n38084), .X(n45390) );
  nand_x1_sg U51911 ( .A(n38017), .B(n38018), .X(n45357) );
  nand_x1_sg U51912 ( .A(n38061), .B(n38062), .X(n45379) );
  nand_x1_sg U51913 ( .A(n36905), .B(n36906), .X(n44801) );
  nand_x1_sg U51914 ( .A(n37921), .B(n37922), .X(n45309) );
  nand_x1_sg U51915 ( .A(n38059), .B(n38060), .X(n45378) );
  nand_x1_sg U51916 ( .A(n37929), .B(n37930), .X(n45313) );
  nand_x1_sg U51917 ( .A(n38067), .B(n38068), .X(n45382) );
  nand_x1_sg U51918 ( .A(n37927), .B(n37928), .X(n45312) );
  nand_x1_sg U51919 ( .A(n38065), .B(n38066), .X(n45381) );
  nand_x1_sg U51920 ( .A(n37951), .B(n37952), .X(n45324) );
  nand_x1_sg U51921 ( .A(n38057), .B(n38058), .X(n45377) );
  nand_x1_sg U51922 ( .A(n37949), .B(n37950), .X(n45323) );
  nand_x1_sg U51923 ( .A(n38063), .B(n38064), .X(n45380) );
  nand_x1_sg U51924 ( .A(n36299), .B(n36300), .X(n44498) );
  nand_x1_sg U51925 ( .A(n38049), .B(n38050), .X(n45373) );
  nand_x1_sg U51926 ( .A(n37953), .B(n37954), .X(n45325) );
  nand_x1_sg U51927 ( .A(n38055), .B(n38056), .X(n45376) );
  nand_x1_sg U51928 ( .A(n37939), .B(n37940), .X(n45318) );
  nand_x1_sg U51929 ( .A(n38081), .B(n38082), .X(n45389) );
  nand_x1_sg U51930 ( .A(n37937), .B(n37938), .X(n45317) );
  nand_x1_sg U51931 ( .A(n38079), .B(n38080), .X(n45388) );
  nand_x1_sg U51932 ( .A(n37945), .B(n37946), .X(n45321) );
  nand_x1_sg U51933 ( .A(n37523), .B(n37524), .X(n45110) );
  nand_x1_sg U51934 ( .A(n37943), .B(n37944), .X(n45320) );
  nand_x1_sg U51935 ( .A(n37537), .B(n37538), .X(n45117) );
  nand_x1_sg U51936 ( .A(n37901), .B(n37902), .X(n45299) );
  nand_x1_sg U51937 ( .A(n38069), .B(n38070), .X(n45383) );
  nand_x1_sg U51938 ( .A(n37899), .B(n37900), .X(n45298) );
  nand_x1_sg U51939 ( .A(n37531), .B(n37532), .X(n45114) );
  nand_x1_sg U51940 ( .A(n37451), .B(n37452), .X(n45074) );
  nand_x1_sg U51941 ( .A(n38071), .B(n38072), .X(n45384) );
  nand_x1_sg U51942 ( .A(n37453), .B(n37454), .X(n45075) );
  nand_x1_sg U51943 ( .A(n37505), .B(n37506), .X(n45101) );
  nand_x1_sg U51944 ( .A(n36257), .B(n36258), .X(n44477) );
  nand_x1_sg U51945 ( .A(n37511), .B(n37512), .X(n45104) );
  nand_x1_sg U51946 ( .A(n36259), .B(n36260), .X(n44478) );
  nand_x1_sg U51947 ( .A(n37517), .B(n37518), .X(n45107) );
  nand_x1_sg U51948 ( .A(n37895), .B(n37896), .X(n45296) );
  nand_x1_sg U51949 ( .A(n37935), .B(n37936), .X(n45316) );
  nand_x1_sg U51950 ( .A(n37893), .B(n37894), .X(n45295) );
  nand_x1_sg U51951 ( .A(n37933), .B(n37934), .X(n45315) );
  nand_x1_sg U51952 ( .A(n37913), .B(n37914), .X(n45305) );
  nand_x1_sg U51953 ( .A(n37923), .B(n37924), .X(n45310) );
  nand_x1_sg U51954 ( .A(n37977), .B(n37978), .X(n45337) );
  nand_x1_sg U51955 ( .A(n37911), .B(n37912), .X(n45304) );
  nand_x1_sg U51956 ( .A(n37449), .B(n37450), .X(n45073) );
  nand_x1_sg U51957 ( .A(n37917), .B(n37918), .X(n45307) );
  nand_x1_sg U51958 ( .A(n37981), .B(n37982), .X(n45339) );
  nand_x1_sg U51959 ( .A(n37915), .B(n37916), .X(n45306) );
  nand_x1_sg U51960 ( .A(n37979), .B(n37980), .X(n45338) );
  nand_x1_sg U51961 ( .A(n37905), .B(n37906), .X(n45301) );
  nand_x1_sg U51962 ( .A(n36749), .B(n36750), .X(n44723) );
  nand_x1_sg U51963 ( .A(n37903), .B(n37904), .X(n45300) );
  nand_x1_sg U51964 ( .A(n36785), .B(n36786), .X(n44741) );
  nand_x1_sg U51965 ( .A(n37909), .B(n37910), .X(n45303) );
  nand_x1_sg U51966 ( .A(n37959), .B(n37960), .X(n45328) );
  nand_x1_sg U51967 ( .A(n37907), .B(n37908), .X(n45302) );
  nand_x1_sg U51968 ( .A(n36773), .B(n36774), .X(n44735) );
  nand_x1_sg U51969 ( .A(n37971), .B(n37972), .X(n45334) );
  nand_x1_sg U51970 ( .A(n37955), .B(n37956), .X(n45326) );
  nand_x1_sg U51971 ( .A(n37969), .B(n37970), .X(n45333) );
  nand_x1_sg U51972 ( .A(n36857), .B(n36858), .X(n44777) );
  nand_x1_sg U51973 ( .A(n37975), .B(n37976), .X(n45336) );
  nand_x1_sg U51974 ( .A(n36683), .B(n36684), .X(n44690) );
  nand_x1_sg U51975 ( .A(n37973), .B(n37974), .X(n45335) );
  nand_x1_sg U51976 ( .A(n36635), .B(n36636), .X(n44666) );
  nand_x1_sg U51977 ( .A(n37963), .B(n37964), .X(n45330) );
  nand_x1_sg U51978 ( .A(n38117), .B(n38118), .X(n45407) );
  nand_x1_sg U51979 ( .A(n37961), .B(n37962), .X(n45329) );
  nand_x1_sg U51980 ( .A(n36437), .B(n36438), .X(n44567) );
  nand_x1_sg U51981 ( .A(n37967), .B(n37968), .X(n45332) );
  nand_x1_sg U51982 ( .A(n36611), .B(n36612), .X(n44654) );
  nand_x1_sg U51983 ( .A(n37965), .B(n37966), .X(n45331) );
  nand_x1_sg U51984 ( .A(n36623), .B(n36624), .X(n44660) );
  nand_x1_sg U51985 ( .A(n38307), .B(n38308), .X(n45502) );
  nand_x1_sg U51986 ( .A(n38109), .B(n38110), .X(n45403) );
  nand_x1_sg U51987 ( .A(n38305), .B(n38306), .X(n45501) );
  nand_x1_sg U51988 ( .A(n36641), .B(n36642), .X(n44669) );
  nand_x1_sg U51989 ( .A(n37987), .B(n37988), .X(n45342) );
  nand_x1_sg U51990 ( .A(n38175), .B(n38176), .X(n45436) );
  nand_x1_sg U51991 ( .A(n36255), .B(n36256), .X(n44476) );
  nand_x1_sg U51992 ( .A(n57607), .B(n39834), .X(n10398) );
  nand_x1_sg U51993 ( .A(n38647), .B(n38648), .X(n45669) );
  nand_x1_sg U51994 ( .A(w_15[19]), .B(n57569), .X(n38648) );
  nand_x1_sg U51995 ( .A(n39631), .B(n39632), .X(n46161) );
  nand_x1_sg U51996 ( .A(w_15[18]), .B(n57604), .X(n39632) );
  nand_x1_sg U51997 ( .A(n39559), .B(n39560), .X(n46125) );
  nand_x1_sg U51998 ( .A(w_15[17]), .B(n57601), .X(n39560) );
  nand_x1_sg U51999 ( .A(n39529), .B(n39530), .X(n46110) );
  nand_x1_sg U52000 ( .A(w_15[16]), .B(n57563), .X(n39530) );
  nand_x1_sg U52001 ( .A(n39271), .B(n39272), .X(n45981) );
  nand_x1_sg U52002 ( .A(w_15[15]), .B(n57621), .X(n39272) );
  nand_x1_sg U52003 ( .A(n38641), .B(n38642), .X(n45666) );
  nand_x1_sg U52004 ( .A(w_15[14]), .B(n57569), .X(n38642) );
  nand_x1_sg U52005 ( .A(n39385), .B(n39386), .X(n46038) );
  nand_x1_sg U52006 ( .A(w_15[13]), .B(n57630), .X(n39386) );
  nand_x1_sg U52007 ( .A(n39391), .B(n39392), .X(n46041) );
  nand_x1_sg U52008 ( .A(w_15[12]), .B(n57569), .X(n39392) );
  nand_x1_sg U52009 ( .A(n38743), .B(n38744), .X(n45717) );
  nand_x1_sg U52010 ( .A(w_15[11]), .B(n57573), .X(n38744) );
  nand_x1_sg U52011 ( .A(n39397), .B(n39398), .X(n46044) );
  nand_x1_sg U52012 ( .A(w_15[10]), .B(n57615), .X(n39398) );
  nand_x1_sg U52013 ( .A(n39403), .B(n39404), .X(n46047) );
  nand_x1_sg U52014 ( .A(w_15[9]), .B(n57624), .X(n39404) );
  nand_x1_sg U52015 ( .A(n38735), .B(n38736), .X(n45713) );
  nand_x1_sg U52016 ( .A(w_15[8]), .B(n57572), .X(n38736) );
  nand_x1_sg U52017 ( .A(n39193), .B(n39194), .X(n45942) );
  nand_x1_sg U52018 ( .A(w_15[7]), .B(n57596), .X(n39194) );
  nand_x1_sg U52019 ( .A(n38737), .B(n38738), .X(n45714) );
  nand_x1_sg U52020 ( .A(w_15[6]), .B(n57572), .X(n38738) );
  nand_x1_sg U52021 ( .A(n39199), .B(n39200), .X(n45945) );
  nand_x1_sg U52022 ( .A(w_15[5]), .B(n57596), .X(n39200) );
  nand_x1_sg U52023 ( .A(n39205), .B(n39206), .X(n45948) );
  nand_x1_sg U52024 ( .A(w_15[4]), .B(n57596), .X(n39206) );
  nand_x1_sg U52025 ( .A(n39211), .B(n39212), .X(n45951) );
  nand_x1_sg U52026 ( .A(w_15[3]), .B(n57597), .X(n39212) );
  nand_x1_sg U52027 ( .A(n39265), .B(n39266), .X(n45978) );
  nand_x1_sg U52028 ( .A(w_15[2]), .B(n57600), .X(n39266) );
  nand_x1_sg U52029 ( .A(n38745), .B(n38746), .X(n45718) );
  nand_x1_sg U52030 ( .A(w_15[1]), .B(n57573), .X(n38746) );
  nand_x1_sg U52031 ( .A(n38747), .B(n38748), .X(n45719) );
  nand_x1_sg U52032 ( .A(w_15[0]), .B(n57573), .X(n38748) );
  nand_x1_sg U52033 ( .A(n38739), .B(n38740), .X(n45715) );
  nand_x1_sg U52034 ( .A(w_14[19]), .B(n57573), .X(n38740) );
  nand_x1_sg U52035 ( .A(n38741), .B(n38742), .X(n45716) );
  nand_x1_sg U52036 ( .A(w_14[18]), .B(n57573), .X(n38742) );
  nand_x1_sg U52037 ( .A(n39393), .B(n39394), .X(n46042) );
  nand_x1_sg U52038 ( .A(w_14[17]), .B(n57625), .X(n39394) );
  nand_x1_sg U52039 ( .A(n39395), .B(n39396), .X(n46043) );
  nand_x1_sg U52040 ( .A(w_14[16]), .B(n57629), .X(n39396) );
  nand_x1_sg U52041 ( .A(n39387), .B(n39388), .X(n46039) );
  nand_x1_sg U52042 ( .A(w_14[15]), .B(n57630), .X(n39388) );
  nand_x1_sg U52043 ( .A(n39389), .B(n39390), .X(n46040) );
  nand_x1_sg U52044 ( .A(w_14[14]), .B(n57568), .X(n39390) );
  nand_x1_sg U52045 ( .A(n39405), .B(n39406), .X(n46048) );
  nand_x1_sg U52046 ( .A(w_14[13]), .B(n57617), .X(n39406) );
  nand_x1_sg U52047 ( .A(n39407), .B(n39408), .X(n46049) );
  nand_x1_sg U52048 ( .A(w_14[12]), .B(n57622), .X(n39408) );
  nand_x1_sg U52049 ( .A(n39399), .B(n39400), .X(n46045) );
  nand_x1_sg U52050 ( .A(w_14[11]), .B(n57569), .X(n39400) );
  nand_x1_sg U52051 ( .A(n39401), .B(n39402), .X(n46046) );
  nand_x1_sg U52052 ( .A(w_14[10]), .B(n57564), .X(n39402) );
  nand_x1_sg U52053 ( .A(n39441), .B(n39442), .X(n46066) );
  nand_x1_sg U52054 ( .A(w_14[9]), .B(n57600), .X(n39442) );
  nand_x1_sg U52055 ( .A(n39443), .B(n39444), .X(n46067) );
  nand_x1_sg U52056 ( .A(w_14[8]), .B(n57625), .X(n39444) );
  nand_x1_sg U52057 ( .A(n39435), .B(n39436), .X(n46063) );
  nand_x1_sg U52058 ( .A(w_14[7]), .B(n57600), .X(n39436) );
  nand_x1_sg U52059 ( .A(n39437), .B(n39438), .X(n46064) );
  nand_x1_sg U52060 ( .A(w_14[6]), .B(n57600), .X(n39438) );
  nand_x1_sg U52061 ( .A(n39453), .B(n39454), .X(n46072) );
  nand_x1_sg U52062 ( .A(w_14[5]), .B(n57600), .X(n39454) );
  nand_x1_sg U52063 ( .A(n39455), .B(n39456), .X(n46073) );
  nand_x1_sg U52064 ( .A(w_14[4]), .B(n57629), .X(n39456) );
  nand_x1_sg U52065 ( .A(n39447), .B(n39448), .X(n46069) );
  nand_x1_sg U52066 ( .A(w_14[3]), .B(n57622), .X(n39448) );
  nand_x1_sg U52067 ( .A(n39449), .B(n39450), .X(n46070) );
  nand_x1_sg U52068 ( .A(w_14[2]), .B(n57623), .X(n39450) );
  nand_x1_sg U52069 ( .A(n39417), .B(n39418), .X(n46054) );
  nand_x1_sg U52070 ( .A(w_14[1]), .B(n57600), .X(n39418) );
  nand_x1_sg U52071 ( .A(n39419), .B(n39420), .X(n46055) );
  nand_x1_sg U52072 ( .A(w_14[0]), .B(n57618), .X(n39420) );
  nand_x1_sg U52073 ( .A(n39411), .B(n39412), .X(n46051) );
  nand_x1_sg U52074 ( .A(w_13[19]), .B(n57623), .X(n39412) );
  nand_x1_sg U52075 ( .A(n39413), .B(n39414), .X(n46052) );
  nand_x1_sg U52076 ( .A(w_13[18]), .B(n57620), .X(n39414) );
  nand_x1_sg U52077 ( .A(n39429), .B(n39430), .X(n46060) );
  nand_x1_sg U52078 ( .A(w_13[17]), .B(n57600), .X(n39430) );
  nand_x1_sg U52079 ( .A(n39431), .B(n39432), .X(n46061) );
  nand_x1_sg U52080 ( .A(w_13[16]), .B(n57600), .X(n39432) );
  nand_x1_sg U52081 ( .A(n39423), .B(n39424), .X(n46057) );
  nand_x1_sg U52082 ( .A(w_13[15]), .B(n57600), .X(n39424) );
  nand_x1_sg U52083 ( .A(n39425), .B(n39426), .X(n46058) );
  nand_x1_sg U52084 ( .A(w_13[14]), .B(n57600), .X(n39426) );
  nand_x1_sg U52085 ( .A(n39489), .B(n39490), .X(n46090) );
  nand_x1_sg U52086 ( .A(w_13[13]), .B(n57625), .X(n39490) );
  nand_x1_sg U52087 ( .A(n39491), .B(n39492), .X(n46091) );
  nand_x1_sg U52088 ( .A(w_13[12]), .B(n57624), .X(n39492) );
  nand_x1_sg U52089 ( .A(n39483), .B(n39484), .X(n46087) );
  nand_x1_sg U52090 ( .A(w_13[11]), .B(n57624), .X(n39484) );
  nand_x1_sg U52091 ( .A(n39485), .B(n39486), .X(n46088) );
  nand_x1_sg U52092 ( .A(w_13[10]), .B(n57624), .X(n39486) );
  nand_x1_sg U52093 ( .A(n39501), .B(n39502), .X(n46096) );
  nand_x1_sg U52094 ( .A(w_13[9]), .B(n57562), .X(n39502) );
  nand_x1_sg U52095 ( .A(n39503), .B(n39504), .X(n46097) );
  nand_x1_sg U52096 ( .A(w_13[8]), .B(n57618), .X(n39504) );
  nand_x1_sg U52097 ( .A(n39495), .B(n39496), .X(n46093) );
  nand_x1_sg U52098 ( .A(w_13[7]), .B(n57615), .X(n39496) );
  nand_x1_sg U52099 ( .A(n39497), .B(n39498), .X(n46094) );
  nand_x1_sg U52100 ( .A(w_13[6]), .B(n57562), .X(n39498) );
  nand_x1_sg U52101 ( .A(n39465), .B(n39466), .X(n46078) );
  nand_x1_sg U52102 ( .A(w_13[5]), .B(n57632), .X(n39466) );
  nand_x1_sg U52103 ( .A(n39467), .B(n39468), .X(n46079) );
  nand_x1_sg U52104 ( .A(w_13[4]), .B(n57568), .X(n39468) );
  nand_x1_sg U52105 ( .A(n39459), .B(n39460), .X(n46075) );
  nand_x1_sg U52106 ( .A(w_13[3]), .B(n57569), .X(n39460) );
  nand_x1_sg U52107 ( .A(n39461), .B(n39462), .X(n46076) );
  nand_x1_sg U52108 ( .A(w_13[2]), .B(n57566), .X(n39462) );
  nand_x1_sg U52109 ( .A(n39477), .B(n39478), .X(n46084) );
  nand_x1_sg U52110 ( .A(w_13[1]), .B(n57624), .X(n39478) );
  nand_x1_sg U52111 ( .A(n39479), .B(n39480), .X(n46085) );
  nand_x1_sg U52112 ( .A(w_13[0]), .B(n57624), .X(n39480) );
  nand_x1_sg U52113 ( .A(n39471), .B(n39472), .X(n46081) );
  nand_x1_sg U52114 ( .A(w_12[19]), .B(n57615), .X(n39472) );
  nand_x1_sg U52115 ( .A(n39473), .B(n39474), .X(n46082) );
  nand_x1_sg U52116 ( .A(w_12[18]), .B(n57618), .X(n39474) );
  nand_x1_sg U52117 ( .A(n39633), .B(n39634), .X(n46162) );
  nand_x1_sg U52118 ( .A(w_12[17]), .B(n57604), .X(n39634) );
  nand_x1_sg U52119 ( .A(n39635), .B(n39636), .X(n46163) );
  nand_x1_sg U52120 ( .A(w_12[16]), .B(n57604), .X(n39636) );
  nand_x1_sg U52121 ( .A(n39627), .B(n39628), .X(n46159) );
  nand_x1_sg U52122 ( .A(w_12[15]), .B(n57604), .X(n39628) );
  nand_x1_sg U52123 ( .A(n39629), .B(n39630), .X(n46160) );
  nand_x1_sg U52124 ( .A(w_12[14]), .B(n57604), .X(n39630) );
  nand_x1_sg U52125 ( .A(n39645), .B(n39646), .X(n46168) );
  nand_x1_sg U52126 ( .A(w_12[13]), .B(n57605), .X(n39646) );
  nand_x1_sg U52127 ( .A(n39647), .B(n39648), .X(n46169) );
  nand_x1_sg U52128 ( .A(w_12[12]), .B(n57605), .X(n39648) );
  nand_x1_sg U52129 ( .A(n39639), .B(n39640), .X(n46165) );
  nand_x1_sg U52130 ( .A(w_12[11]), .B(n57605), .X(n39640) );
  nand_x1_sg U52131 ( .A(n39641), .B(n39642), .X(n46166) );
  nand_x1_sg U52132 ( .A(w_12[10]), .B(n57605), .X(n39642) );
  nand_x1_sg U52133 ( .A(n39609), .B(n39610), .X(n46150) );
  nand_x1_sg U52134 ( .A(w_12[9]), .B(n57603), .X(n39610) );
  nand_x1_sg U52135 ( .A(n39611), .B(n39612), .X(n46151) );
  nand_x1_sg U52136 ( .A(w_12[8]), .B(n57603), .X(n39612) );
  nand_x1_sg U52137 ( .A(n39603), .B(n39604), .X(n46147) );
  nand_x1_sg U52138 ( .A(w_12[7]), .B(n57603), .X(n39604) );
  nand_x1_sg U52139 ( .A(n39605), .B(n39606), .X(n46148) );
  nand_x1_sg U52140 ( .A(w_12[6]), .B(n57603), .X(n39606) );
  nand_x1_sg U52141 ( .A(n39621), .B(n39622), .X(n46156) );
  nand_x1_sg U52142 ( .A(w_12[5]), .B(n57604), .X(n39622) );
  nand_x1_sg U52143 ( .A(n39623), .B(n39624), .X(n46157) );
  nand_x1_sg U52144 ( .A(w_12[4]), .B(n57604), .X(n39624) );
  nand_x1_sg U52145 ( .A(n39615), .B(n39616), .X(n46153) );
  nand_x1_sg U52146 ( .A(w_12[3]), .B(n57603), .X(n39616) );
  nand_x1_sg U52147 ( .A(n39617), .B(n39618), .X(n46154) );
  nand_x1_sg U52148 ( .A(w_12[2]), .B(n57603), .X(n39618) );
  nand_x1_sg U52149 ( .A(n39681), .B(n39682), .X(n46186) );
  nand_x1_sg U52150 ( .A(w_12[1]), .B(n57606), .X(n39682) );
  nand_x1_sg U52151 ( .A(n39683), .B(n39684), .X(n46187) );
  nand_x1_sg U52152 ( .A(w_12[0]), .B(n57606), .X(n39684) );
  nand_x1_sg U52153 ( .A(n39675), .B(n39676), .X(n46183) );
  nand_x1_sg U52154 ( .A(w_11[19]), .B(n57606), .X(n39676) );
  nand_x1_sg U52155 ( .A(n39677), .B(n39678), .X(n46184) );
  nand_x1_sg U52156 ( .A(w_11[18]), .B(n57606), .X(n39678) );
  nand_x1_sg U52157 ( .A(n39693), .B(n39694), .X(n46192) );
  nand_x1_sg U52158 ( .A(w_11[17]), .B(n57628), .X(n39694) );
  nand_x1_sg U52159 ( .A(n39695), .B(n39696), .X(n46193) );
  nand_x1_sg U52160 ( .A(w_11[16]), .B(n57625), .X(n39696) );
  nand_x1_sg U52161 ( .A(n39687), .B(n39688), .X(n46189) );
  nand_x1_sg U52162 ( .A(w_11[15]), .B(n57606), .X(n39688) );
  nand_x1_sg U52163 ( .A(n39689), .B(n39690), .X(n46190) );
  nand_x1_sg U52164 ( .A(w_11[14]), .B(n57606), .X(n39690) );
  nand_x1_sg U52165 ( .A(n39657), .B(n39658), .X(n46174) );
  nand_x1_sg U52166 ( .A(w_11[13]), .B(n57622), .X(n39658) );
  nand_x1_sg U52167 ( .A(n39659), .B(n39660), .X(n46175) );
  nand_x1_sg U52168 ( .A(w_11[12]), .B(n57622), .X(n39660) );
  nand_x1_sg U52169 ( .A(n39651), .B(n39652), .X(n46171) );
  nand_x1_sg U52170 ( .A(w_11[11]), .B(n57605), .X(n39652) );
  nand_x1_sg U52171 ( .A(n39653), .B(n39654), .X(n46172) );
  nand_x1_sg U52172 ( .A(w_11[10]), .B(n57605), .X(n39654) );
  nand_x1_sg U52173 ( .A(n39669), .B(n39670), .X(n46180) );
  nand_x1_sg U52174 ( .A(w_11[9]), .B(n57622), .X(n39670) );
  nand_x1_sg U52175 ( .A(n39671), .B(n39672), .X(n46181) );
  nand_x1_sg U52176 ( .A(w_11[8]), .B(n57622), .X(n39672) );
  nand_x1_sg U52177 ( .A(n39663), .B(n39664), .X(n46177) );
  nand_x1_sg U52178 ( .A(w_11[7]), .B(n57622), .X(n39664) );
  nand_x1_sg U52179 ( .A(n39665), .B(n39666), .X(n46178) );
  nand_x1_sg U52180 ( .A(w_11[6]), .B(n57622), .X(n39666) );
  nand_x1_sg U52181 ( .A(n39537), .B(n39538), .X(n46114) );
  nand_x1_sg U52182 ( .A(w_11[5]), .B(n57568), .X(n39538) );
  nand_x1_sg U52183 ( .A(n39539), .B(n39540), .X(n46115) );
  nand_x1_sg U52184 ( .A(w_11[4]), .B(n57568), .X(n39540) );
  nand_x1_sg U52185 ( .A(n39531), .B(n39532), .X(n46111) );
  nand_x1_sg U52186 ( .A(w_11[3]), .B(n57569), .X(n39532) );
  nand_x1_sg U52187 ( .A(n39533), .B(n39534), .X(n46112) );
  nand_x1_sg U52188 ( .A(w_11[2]), .B(n57566), .X(n39534) );
  nand_x1_sg U52189 ( .A(n39549), .B(n39550), .X(n46120) );
  nand_x1_sg U52190 ( .A(w_11[1]), .B(n57601), .X(n39550) );
  nand_x1_sg U52191 ( .A(n39551), .B(n39552), .X(n46121) );
  nand_x1_sg U52192 ( .A(w_11[0]), .B(n57601), .X(n39552) );
  nand_x1_sg U52193 ( .A(n39543), .B(n39544), .X(n46117) );
  nand_x1_sg U52194 ( .A(w_10[19]), .B(n57564), .X(n39544) );
  nand_x1_sg U52195 ( .A(n39545), .B(n39546), .X(n46118) );
  nand_x1_sg U52196 ( .A(w_10[18]), .B(n57624), .X(n39546) );
  nand_x1_sg U52197 ( .A(n39513), .B(n39514), .X(n46102) );
  nand_x1_sg U52198 ( .A(w_10[17]), .B(n57619), .X(n39514) );
  nand_x1_sg U52199 ( .A(n39515), .B(n39516), .X(n46103) );
  nand_x1_sg U52200 ( .A(w_10[16]), .B(n57567), .X(n39516) );
  nand_x1_sg U52201 ( .A(n39507), .B(n39508), .X(n46099) );
  nand_x1_sg U52202 ( .A(w_10[15]), .B(n57616), .X(n39508) );
  nand_x1_sg U52203 ( .A(n39509), .B(n39510), .X(n46100) );
  nand_x1_sg U52204 ( .A(w_10[14]), .B(n57615), .X(n39510) );
  nand_x1_sg U52205 ( .A(n39525), .B(n39526), .X(n46108) );
  nand_x1_sg U52206 ( .A(w_10[13]), .B(n57564), .X(n39526) );
  nand_x1_sg U52207 ( .A(n39527), .B(n39528), .X(n46109) );
  nand_x1_sg U52208 ( .A(w_10[12]), .B(n57565), .X(n39528) );
  nand_x1_sg U52209 ( .A(n39519), .B(n39520), .X(n46105) );
  nand_x1_sg U52210 ( .A(w_10[11]), .B(n57568), .X(n39520) );
  nand_x1_sg U52211 ( .A(n39521), .B(n39522), .X(n46106) );
  nand_x1_sg U52212 ( .A(w_10[10]), .B(n57619), .X(n39522) );
  nand_x1_sg U52213 ( .A(n39585), .B(n39586), .X(n46138) );
  nand_x1_sg U52214 ( .A(w_10[9]), .B(n57601), .X(n39586) );
  nand_x1_sg U52215 ( .A(n39587), .B(n39588), .X(n46139) );
  nand_x1_sg U52216 ( .A(w_10[8]), .B(n57566), .X(n39588) );
  nand_x1_sg U52217 ( .A(n39579), .B(n39580), .X(n46135) );
  nand_x1_sg U52218 ( .A(w_10[7]), .B(n57602), .X(n39580) );
  nand_x1_sg U52219 ( .A(n39581), .B(n39582), .X(n46136) );
  nand_x1_sg U52220 ( .A(w_10[6]), .B(n57602), .X(n39582) );
  nand_x1_sg U52221 ( .A(n39597), .B(n39598), .X(n46144) );
  nand_x1_sg U52222 ( .A(w_10[5]), .B(n57603), .X(n39598) );
  nand_x1_sg U52223 ( .A(n39599), .B(n39600), .X(n46145) );
  nand_x1_sg U52224 ( .A(w_10[4]), .B(n57602), .X(n39600) );
  nand_x1_sg U52225 ( .A(n39591), .B(n39592), .X(n46141) );
  nand_x1_sg U52226 ( .A(w_10[3]), .B(n57567), .X(n39592) );
  nand_x1_sg U52227 ( .A(n39593), .B(n39594), .X(n46142) );
  nand_x1_sg U52228 ( .A(w_10[2]), .B(n57606), .X(n39594) );
  nand_x1_sg U52229 ( .A(n39561), .B(n39562), .X(n46126) );
  nand_x1_sg U52230 ( .A(w_10[1]), .B(n57601), .X(n39562) );
  nand_x1_sg U52231 ( .A(n39563), .B(n39564), .X(n46127) );
  nand_x1_sg U52232 ( .A(w_10[0]), .B(n57601), .X(n39564) );
  nand_x1_sg U52233 ( .A(n39555), .B(n39556), .X(n46123) );
  nand_x1_sg U52234 ( .A(w_9[19]), .B(n57601), .X(n39556) );
  nand_x1_sg U52235 ( .A(n39557), .B(n39558), .X(n46124) );
  nand_x1_sg U52236 ( .A(w_9[18]), .B(n57601), .X(n39558) );
  nand_x1_sg U52237 ( .A(n39573), .B(n39574), .X(n46132) );
  nand_x1_sg U52238 ( .A(w_9[17]), .B(n57602), .X(n39574) );
  nand_x1_sg U52239 ( .A(n39575), .B(n39576), .X(n46133) );
  nand_x1_sg U52240 ( .A(w_9[16]), .B(n57602), .X(n39576) );
  nand_x1_sg U52241 ( .A(n39567), .B(n39568), .X(n46129) );
  nand_x1_sg U52242 ( .A(w_9[15]), .B(n57602), .X(n39568) );
  nand_x1_sg U52243 ( .A(n39569), .B(n39570), .X(n46130) );
  nand_x1_sg U52244 ( .A(w_9[14]), .B(n57602), .X(n39570) );
  nand_x1_sg U52245 ( .A(n39129), .B(n39130), .X(n45910) );
  nand_x1_sg U52246 ( .A(w_9[13]), .B(n57592), .X(n39130) );
  nand_x1_sg U52247 ( .A(n39131), .B(n39132), .X(n45911) );
  nand_x1_sg U52248 ( .A(w_9[12]), .B(n57592), .X(n39132) );
  nand_x1_sg U52249 ( .A(n39123), .B(n39124), .X(n45907) );
  nand_x1_sg U52250 ( .A(w_9[11]), .B(n57592), .X(n39124) );
  nand_x1_sg U52251 ( .A(n39125), .B(n39126), .X(n45908) );
  nand_x1_sg U52252 ( .A(w_9[10]), .B(n57592), .X(n39126) );
  nand_x1_sg U52253 ( .A(n39141), .B(n39142), .X(n45916) );
  nand_x1_sg U52254 ( .A(w_9[9]), .B(n57593), .X(n39142) );
  nand_x1_sg U52255 ( .A(n39143), .B(n39144), .X(n45917) );
  nand_x1_sg U52256 ( .A(w_9[8]), .B(n57593), .X(n39144) );
  nand_x1_sg U52257 ( .A(n39135), .B(n39136), .X(n45913) );
  nand_x1_sg U52258 ( .A(w_9[7]), .B(n57593), .X(n39136) );
  nand_x1_sg U52259 ( .A(n39137), .B(n39138), .X(n45914) );
  nand_x1_sg U52260 ( .A(w_9[6]), .B(n57593), .X(n39138) );
  nand_x1_sg U52261 ( .A(n39105), .B(n39106), .X(n45898) );
  nand_x1_sg U52262 ( .A(w_9[5]), .B(n57591), .X(n39106) );
  nand_x1_sg U52263 ( .A(n39107), .B(n39108), .X(n45899) );
  nand_x1_sg U52264 ( .A(w_9[4]), .B(n57591), .X(n39108) );
  nand_x1_sg U52265 ( .A(n39099), .B(n39100), .X(n45895) );
  nand_x1_sg U52266 ( .A(w_9[3]), .B(n57591), .X(n39100) );
  nand_x1_sg U52267 ( .A(n39101), .B(n39102), .X(n45896) );
  nand_x1_sg U52268 ( .A(w_9[2]), .B(n57591), .X(n39102) );
  nand_x1_sg U52269 ( .A(n39117), .B(n39118), .X(n45904) );
  nand_x1_sg U52270 ( .A(w_9[1]), .B(n57592), .X(n39118) );
  nand_x1_sg U52271 ( .A(n39119), .B(n39120), .X(n45905) );
  nand_x1_sg U52272 ( .A(w_9[0]), .B(n57592), .X(n39120) );
  nand_x1_sg U52273 ( .A(n39111), .B(n39112), .X(n45901) );
  nand_x1_sg U52274 ( .A(w_8[19]), .B(n57591), .X(n39112) );
  nand_x1_sg U52275 ( .A(n39113), .B(n39114), .X(n45902) );
  nand_x1_sg U52276 ( .A(w_8[18]), .B(n57591), .X(n39114) );
  nand_x1_sg U52277 ( .A(n39177), .B(n39178), .X(n45934) );
  nand_x1_sg U52278 ( .A(w_8[17]), .B(n57595), .X(n39178) );
  nand_x1_sg U52279 ( .A(n39179), .B(n39180), .X(n45935) );
  nand_x1_sg U52280 ( .A(w_8[16]), .B(n57595), .X(n39180) );
  nand_x1_sg U52281 ( .A(n39171), .B(n39172), .X(n45931) );
  nand_x1_sg U52282 ( .A(w_8[15]), .B(n57595), .X(n39172) );
  nand_x1_sg U52283 ( .A(n39173), .B(n39174), .X(n45932) );
  nand_x1_sg U52284 ( .A(w_8[14]), .B(n57595), .X(n39174) );
  nand_x1_sg U52285 ( .A(n39189), .B(n39190), .X(n45940) );
  nand_x1_sg U52286 ( .A(w_8[13]), .B(n57596), .X(n39190) );
  nand_x1_sg U52287 ( .A(n39191), .B(n39192), .X(n45941) );
  nand_x1_sg U52288 ( .A(w_8[12]), .B(n57596), .X(n39192) );
  nand_x1_sg U52289 ( .A(n39183), .B(n39184), .X(n45937) );
  nand_x1_sg U52290 ( .A(w_8[11]), .B(n57595), .X(n39184) );
  nand_x1_sg U52291 ( .A(n39185), .B(n39186), .X(n45938) );
  nand_x1_sg U52292 ( .A(w_8[10]), .B(n57595), .X(n39186) );
  nand_x1_sg U52293 ( .A(n39153), .B(n39154), .X(n45922) );
  nand_x1_sg U52294 ( .A(w_8[9]), .B(n57594), .X(n39154) );
  nand_x1_sg U52295 ( .A(n39155), .B(n39156), .X(n45923) );
  nand_x1_sg U52296 ( .A(w_8[8]), .B(n57594), .X(n39156) );
  nand_x1_sg U52297 ( .A(n39147), .B(n39148), .X(n45919) );
  nand_x1_sg U52298 ( .A(w_8[7]), .B(n57593), .X(n39148) );
  nand_x1_sg U52299 ( .A(n39149), .B(n39150), .X(n45920) );
  nand_x1_sg U52300 ( .A(w_8[6]), .B(n57593), .X(n39150) );
  nand_x1_sg U52301 ( .A(n39165), .B(n39166), .X(n45928) );
  nand_x1_sg U52302 ( .A(w_8[5]), .B(n57594), .X(n39166) );
  nand_x1_sg U52303 ( .A(n39167), .B(n39168), .X(n45929) );
  nand_x1_sg U52304 ( .A(w_8[4]), .B(n57594), .X(n39168) );
  nand_x1_sg U52305 ( .A(n39159), .B(n39160), .X(n45925) );
  nand_x1_sg U52306 ( .A(w_8[3]), .B(n57594), .X(n39160) );
  nand_x1_sg U52307 ( .A(n39161), .B(n39162), .X(n45926) );
  nand_x1_sg U52308 ( .A(w_8[2]), .B(n57594), .X(n39162) );
  nand_x1_sg U52309 ( .A(n38943), .B(n38944), .X(n45817) );
  nand_x1_sg U52310 ( .A(w_8[1]), .B(n57582), .X(n38944) );
  nand_x1_sg U52311 ( .A(n38945), .B(n38946), .X(n45818) );
  nand_x1_sg U52312 ( .A(w_8[0]), .B(n57582), .X(n38946) );
  nand_x1_sg U52313 ( .A(n38937), .B(n38938), .X(n45814) );
  nand_x1_sg U52314 ( .A(w_7[19]), .B(n57582), .X(n38938) );
  nand_x1_sg U52315 ( .A(n38939), .B(n38940), .X(n45815) );
  nand_x1_sg U52316 ( .A(w_7[18]), .B(n57582), .X(n38940) );
  nand_x1_sg U52317 ( .A(n39035), .B(n39036), .X(n45863) );
  nand_x1_sg U52318 ( .A(w_7[17]), .B(n57587), .X(n39036) );
  nand_x1_sg U52319 ( .A(n38891), .B(n38892), .X(n45791) );
  nand_x1_sg U52320 ( .A(w_7[16]), .B(n57579), .X(n38892) );
  nand_x1_sg U52321 ( .A(n38635), .B(n38636), .X(n45663) );
  nand_x1_sg U52322 ( .A(w_7[15]), .B(n57569), .X(n38636) );
  nand_x1_sg U52323 ( .A(n38689), .B(n38690), .X(n45690) );
  nand_x1_sg U52324 ( .A(w_7[14]), .B(n57570), .X(n38690) );
  nand_x1_sg U52325 ( .A(n38649), .B(n38650), .X(n45670) );
  nand_x1_sg U52326 ( .A(w_7[13]), .B(n57565), .X(n38650) );
  nand_x1_sg U52327 ( .A(n38651), .B(n38652), .X(n45671) );
  nand_x1_sg U52328 ( .A(w_7[12]), .B(n57564), .X(n38652) );
  nand_x1_sg U52329 ( .A(n38643), .B(n38644), .X(n45667) );
  nand_x1_sg U52330 ( .A(w_7[11]), .B(n57569), .X(n38644) );
  nand_x1_sg U52331 ( .A(n38645), .B(n38646), .X(n45668) );
  nand_x1_sg U52332 ( .A(w_7[10]), .B(n57569), .X(n38646) );
  nand_x1_sg U52333 ( .A(n38661), .B(n38662), .X(n45676) );
  nand_x1_sg U52334 ( .A(w_7[9]), .B(n57615), .X(n38662) );
  nand_x1_sg U52335 ( .A(n38663), .B(n38664), .X(n45677) );
  nand_x1_sg U52336 ( .A(w_7[8]), .B(n57567), .X(n38664) );
  nand_x1_sg U52337 ( .A(n38655), .B(n38656), .X(n45673) );
  nand_x1_sg U52338 ( .A(w_7[7]), .B(n57566), .X(n38656) );
  nand_x1_sg U52339 ( .A(n38657), .B(n38658), .X(n45674) );
  nand_x1_sg U52340 ( .A(w_7[6]), .B(n57565), .X(n38658) );
  nand_x1_sg U52341 ( .A(n39081), .B(n39082), .X(n45886) );
  nand_x1_sg U52342 ( .A(w_7[5]), .B(n57590), .X(n39082) );
  nand_x1_sg U52343 ( .A(n39083), .B(n39084), .X(n45887) );
  nand_x1_sg U52344 ( .A(w_7[4]), .B(n57590), .X(n39084) );
  nand_x1_sg U52345 ( .A(n39075), .B(n39076), .X(n45883) );
  nand_x1_sg U52346 ( .A(w_7[3]), .B(n57589), .X(n39076) );
  nand_x1_sg U52347 ( .A(n39077), .B(n39078), .X(n45884) );
  nand_x1_sg U52348 ( .A(w_7[2]), .B(n57589), .X(n39078) );
  nand_x1_sg U52349 ( .A(n39093), .B(n39094), .X(n45892) );
  nand_x1_sg U52350 ( .A(w_7[1]), .B(n57590), .X(n39094) );
  nand_x1_sg U52351 ( .A(n39095), .B(n39096), .X(n45893) );
  nand_x1_sg U52352 ( .A(w_7[0]), .B(n57590), .X(n39096) );
  nand_x1_sg U52353 ( .A(n39087), .B(n39088), .X(n45889) );
  nand_x1_sg U52354 ( .A(w_6[19]), .B(n57590), .X(n39088) );
  nand_x1_sg U52355 ( .A(n39089), .B(n39090), .X(n45890) );
  nand_x1_sg U52356 ( .A(w_6[18]), .B(n57590), .X(n39090) );
  nand_x1_sg U52357 ( .A(n38917), .B(n38918), .X(n45804) );
  nand_x1_sg U52358 ( .A(w_6[17]), .B(n57580), .X(n38918) );
  nand_x1_sg U52359 ( .A(n38979), .B(n38980), .X(n45835) );
  nand_x1_sg U52360 ( .A(w_6[16]), .B(n57584), .X(n38980) );
  nand_x1_sg U52361 ( .A(n39053), .B(n39054), .X(n45872) );
  nand_x1_sg U52362 ( .A(w_6[15]), .B(n57588), .X(n39054) );
  nand_x1_sg U52363 ( .A(n38985), .B(n38986), .X(n45838) );
  nand_x1_sg U52364 ( .A(w_6[14]), .B(n57584), .X(n38986) );
  nand_x1_sg U52365 ( .A(n38931), .B(n38932), .X(n45811) );
  nand_x1_sg U52366 ( .A(w_6[13]), .B(n57581), .X(n38932) );
  nand_x1_sg U52367 ( .A(n38933), .B(n38934), .X(n45812) );
  nand_x1_sg U52368 ( .A(w_6[12]), .B(n57581), .X(n38934) );
  nand_x1_sg U52369 ( .A(n38925), .B(n38926), .X(n45808) );
  nand_x1_sg U52370 ( .A(w_6[11]), .B(n57581), .X(n38926) );
  nand_x1_sg U52371 ( .A(n38927), .B(n38928), .X(n45809) );
  nand_x1_sg U52372 ( .A(w_6[10]), .B(n57581), .X(n38928) );
  nand_x1_sg U52373 ( .A(n39321), .B(n39322), .X(n46006) );
  nand_x1_sg U52374 ( .A(w_6[9]), .B(n57622), .X(n39322) );
  nand_x1_sg U52375 ( .A(n39323), .B(n39324), .X(n46007) );
  nand_x1_sg U52376 ( .A(w_6[8]), .B(n57622), .X(n39324) );
  nand_x1_sg U52377 ( .A(n39315), .B(n39316), .X(n46003) );
  nand_x1_sg U52378 ( .A(w_6[7]), .B(n57624), .X(n39316) );
  nand_x1_sg U52379 ( .A(n39317), .B(n39318), .X(n46004) );
  nand_x1_sg U52380 ( .A(w_6[6]), .B(n57623), .X(n39318) );
  nand_x1_sg U52381 ( .A(n39333), .B(n39334), .X(n46012) );
  nand_x1_sg U52382 ( .A(w_6[5]), .B(n57623), .X(n39334) );
  nand_x1_sg U52383 ( .A(n39335), .B(n39336), .X(n46013) );
  nand_x1_sg U52384 ( .A(w_6[4]), .B(n57620), .X(n39336) );
  nand_x1_sg U52385 ( .A(n39327), .B(n39328), .X(n46009) );
  nand_x1_sg U52386 ( .A(w_6[3]), .B(n57623), .X(n39328) );
  nand_x1_sg U52387 ( .A(n39329), .B(n39330), .X(n46010) );
  nand_x1_sg U52388 ( .A(w_6[2]), .B(n57620), .X(n39330) );
  nand_x1_sg U52389 ( .A(n39297), .B(n39298), .X(n45994) );
  nand_x1_sg U52390 ( .A(w_6[1]), .B(n57622), .X(n39298) );
  nand_x1_sg U52391 ( .A(n39299), .B(n39300), .X(n45995) );
  nand_x1_sg U52392 ( .A(w_6[0]), .B(n57622), .X(n39300) );
  nand_x1_sg U52393 ( .A(n39291), .B(n39292), .X(n45991) );
  nand_x1_sg U52394 ( .A(w_5[19]), .B(n57617), .X(n39292) );
  nand_x1_sg U52395 ( .A(n39293), .B(n39294), .X(n45992) );
  nand_x1_sg U52396 ( .A(w_5[18]), .B(n57600), .X(n39294) );
  nand_x1_sg U52397 ( .A(n39309), .B(n39310), .X(n46000) );
  nand_x1_sg U52398 ( .A(w_5[17]), .B(n57600), .X(n39310) );
  nand_x1_sg U52399 ( .A(n39311), .B(n39312), .X(n46001) );
  nand_x1_sg U52400 ( .A(w_5[16]), .B(n57624), .X(n39312) );
  nand_x1_sg U52401 ( .A(n39303), .B(n39304), .X(n45997) );
  nand_x1_sg U52402 ( .A(w_5[15]), .B(n57617), .X(n39304) );
  nand_x1_sg U52403 ( .A(n39305), .B(n39306), .X(n45998) );
  nand_x1_sg U52404 ( .A(w_5[14]), .B(n57622), .X(n39306) );
  nand_x1_sg U52405 ( .A(n39369), .B(n39370), .X(n46030) );
  nand_x1_sg U52406 ( .A(w_5[13]), .B(n57564), .X(n39370) );
  nand_x1_sg U52407 ( .A(n39371), .B(n39372), .X(n46031) );
  nand_x1_sg U52408 ( .A(w_5[12]), .B(n57632), .X(n39372) );
  nand_x1_sg U52409 ( .A(n39363), .B(n39364), .X(n46027) );
  nand_x1_sg U52410 ( .A(w_5[11]), .B(n57568), .X(n39364) );
  nand_x1_sg U52411 ( .A(n39365), .B(n39366), .X(n46028) );
  nand_x1_sg U52412 ( .A(w_5[10]), .B(n57569), .X(n39366) );
  nand_x1_sg U52413 ( .A(n39381), .B(n39382), .X(n46036) );
  nand_x1_sg U52414 ( .A(w_5[9]), .B(n57632), .X(n39382) );
  nand_x1_sg U52415 ( .A(n39383), .B(n39384), .X(n46037) );
  nand_x1_sg U52416 ( .A(w_5[8]), .B(n57632), .X(n39384) );
  nand_x1_sg U52417 ( .A(n39375), .B(n39376), .X(n46033) );
  nand_x1_sg U52418 ( .A(w_5[7]), .B(n57632), .X(n39376) );
  nand_x1_sg U52419 ( .A(n39377), .B(n39378), .X(n46034) );
  nand_x1_sg U52420 ( .A(w_5[6]), .B(n38414), .X(n39378) );
  nand_x1_sg U52421 ( .A(n39345), .B(n39346), .X(n46018) );
  nand_x1_sg U52422 ( .A(w_5[5]), .B(n57615), .X(n39346) );
  nand_x1_sg U52423 ( .A(n39347), .B(n39348), .X(n46019) );
  nand_x1_sg U52424 ( .A(w_5[4]), .B(n57616), .X(n39348) );
  nand_x1_sg U52425 ( .A(n39339), .B(n39340), .X(n46015) );
  nand_x1_sg U52426 ( .A(w_5[3]), .B(n57621), .X(n39340) );
  nand_x1_sg U52427 ( .A(n39341), .B(n39342), .X(n46016) );
  nand_x1_sg U52428 ( .A(w_5[2]), .B(n57630), .X(n39342) );
  nand_x1_sg U52429 ( .A(n39357), .B(n39358), .X(n46024) );
  nand_x1_sg U52430 ( .A(w_5[1]), .B(n57565), .X(n39358) );
  nand_x1_sg U52431 ( .A(n39359), .B(n39360), .X(n46025) );
  nand_x1_sg U52432 ( .A(w_5[0]), .B(n57567), .X(n39360) );
  nand_x1_sg U52433 ( .A(n39351), .B(n39352), .X(n46021) );
  nand_x1_sg U52434 ( .A(w_4[19]), .B(n57621), .X(n39352) );
  nand_x1_sg U52435 ( .A(n39353), .B(n39354), .X(n46022) );
  nand_x1_sg U52436 ( .A(w_4[18]), .B(n57625), .X(n39354) );
  nand_x1_sg U52437 ( .A(n39225), .B(n39226), .X(n45958) );
  nand_x1_sg U52438 ( .A(w_4[17]), .B(n57598), .X(n39226) );
  nand_x1_sg U52439 ( .A(n39227), .B(n39228), .X(n45959) );
  nand_x1_sg U52440 ( .A(w_4[16]), .B(n57598), .X(n39228) );
  nand_x1_sg U52441 ( .A(n39219), .B(n39220), .X(n45955) );
  nand_x1_sg U52442 ( .A(w_4[15]), .B(n57597), .X(n39220) );
  nand_x1_sg U52443 ( .A(n39221), .B(n39222), .X(n45956) );
  nand_x1_sg U52444 ( .A(w_4[14]), .B(n57597), .X(n39222) );
  nand_x1_sg U52445 ( .A(n39237), .B(n39238), .X(n45964) );
  nand_x1_sg U52446 ( .A(w_4[13]), .B(n57598), .X(n39238) );
  nand_x1_sg U52447 ( .A(n39239), .B(n39240), .X(n45965) );
  nand_x1_sg U52448 ( .A(w_4[12]), .B(n57598), .X(n39240) );
  nand_x1_sg U52449 ( .A(n39231), .B(n39232), .X(n45961) );
  nand_x1_sg U52450 ( .A(w_4[11]), .B(n57598), .X(n39232) );
  nand_x1_sg U52451 ( .A(n39233), .B(n39234), .X(n45962) );
  nand_x1_sg U52452 ( .A(w_4[10]), .B(n57598), .X(n39234) );
  nand_x1_sg U52453 ( .A(n39201), .B(n39202), .X(n45946) );
  nand_x1_sg U52454 ( .A(w_4[9]), .B(n57596), .X(n39202) );
  nand_x1_sg U52455 ( .A(n39203), .B(n39204), .X(n45947) );
  nand_x1_sg U52456 ( .A(w_4[8]), .B(n57596), .X(n39204) );
  nand_x1_sg U52457 ( .A(n39195), .B(n39196), .X(n45943) );
  nand_x1_sg U52458 ( .A(w_4[7]), .B(n57596), .X(n39196) );
  nand_x1_sg U52459 ( .A(n39197), .B(n39198), .X(n45944) );
  nand_x1_sg U52460 ( .A(w_4[6]), .B(n57596), .X(n39198) );
  nand_x1_sg U52461 ( .A(n39213), .B(n39214), .X(n45952) );
  nand_x1_sg U52462 ( .A(w_4[5]), .B(n57597), .X(n39214) );
  nand_x1_sg U52463 ( .A(n39215), .B(n39216), .X(n45953) );
  nand_x1_sg U52464 ( .A(w_4[4]), .B(n57597), .X(n39216) );
  nand_x1_sg U52465 ( .A(n39207), .B(n39208), .X(n45949) );
  nand_x1_sg U52466 ( .A(w_4[3]), .B(n57597), .X(n39208) );
  nand_x1_sg U52467 ( .A(n39209), .B(n39210), .X(n45950) );
  nand_x1_sg U52468 ( .A(w_4[2]), .B(n57597), .X(n39210) );
  nand_x1_sg U52469 ( .A(n39273), .B(n39274), .X(n45982) );
  nand_x1_sg U52470 ( .A(w_4[1]), .B(n57618), .X(n39274) );
  nand_x1_sg U52471 ( .A(n39275), .B(n39276), .X(n45983) );
  nand_x1_sg U52472 ( .A(w_4[0]), .B(n57619), .X(n39276) );
  nand_x1_sg U52473 ( .A(n39267), .B(n39268), .X(n45979) );
  nand_x1_sg U52474 ( .A(w_3[19]), .B(n57624), .X(n39268) );
  nand_x1_sg U52475 ( .A(n39269), .B(n39270), .X(n45980) );
  nand_x1_sg U52476 ( .A(w_3[18]), .B(n57621), .X(n39270) );
  nand_x1_sg U52477 ( .A(n39285), .B(n39286), .X(n45988) );
  nand_x1_sg U52478 ( .A(w_3[17]), .B(n57624), .X(n39286) );
  nand_x1_sg U52479 ( .A(n39287), .B(n39288), .X(n45989) );
  nand_x1_sg U52480 ( .A(w_3[16]), .B(n57567), .X(n39288) );
  nand_x1_sg U52481 ( .A(n39279), .B(n39280), .X(n45985) );
  nand_x1_sg U52482 ( .A(w_3[15]), .B(n57629), .X(n39280) );
  nand_x1_sg U52483 ( .A(n39281), .B(n39282), .X(n45986) );
  nand_x1_sg U52484 ( .A(w_3[14]), .B(n57618), .X(n39282) );
  nand_x1_sg U52485 ( .A(n39249), .B(n39250), .X(n45970) );
  nand_x1_sg U52486 ( .A(w_3[13]), .B(n57599), .X(n39250) );
  nand_x1_sg U52487 ( .A(n39251), .B(n39252), .X(n45971) );
  nand_x1_sg U52488 ( .A(w_3[12]), .B(n57599), .X(n39252) );
  nand_x1_sg U52489 ( .A(n39243), .B(n39244), .X(n45967) );
  nand_x1_sg U52490 ( .A(w_3[11]), .B(n57599), .X(n39244) );
  nand_x1_sg U52491 ( .A(n39245), .B(n39246), .X(n45968) );
  nand_x1_sg U52492 ( .A(w_3[10]), .B(n57599), .X(n39246) );
  nand_x1_sg U52493 ( .A(n39261), .B(n39262), .X(n45976) );
  nand_x1_sg U52494 ( .A(w_3[9]), .B(n57616), .X(n39262) );
  nand_x1_sg U52495 ( .A(n39263), .B(n39264), .X(n45977) );
  nand_x1_sg U52496 ( .A(w_3[8]), .B(n57621), .X(n39264) );
  nand_x1_sg U52497 ( .A(n39255), .B(n39256), .X(n45973) );
  nand_x1_sg U52498 ( .A(w_3[7]), .B(n57599), .X(n39256) );
  nand_x1_sg U52499 ( .A(n39257), .B(n39258), .X(n45974) );
  nand_x1_sg U52500 ( .A(w_3[6]), .B(n57599), .X(n39258) );
  nand_x1_sg U52501 ( .A(n38541), .B(n38542), .X(n45616) );
  nand_x1_sg U52502 ( .A(w_3[5]), .B(n57564), .X(n38542) );
  nand_x1_sg U52503 ( .A(n38543), .B(n38544), .X(n45617) );
  nand_x1_sg U52504 ( .A(w_3[4]), .B(n57564), .X(n38544) );
  nand_x1_sg U52505 ( .A(n38535), .B(n38536), .X(n45613) );
  nand_x1_sg U52506 ( .A(w_3[3]), .B(n57615), .X(n38536) );
  nand_x1_sg U52507 ( .A(n38537), .B(n38538), .X(n45614) );
  nand_x1_sg U52508 ( .A(w_3[2]), .B(n57568), .X(n38538) );
  nand_x1_sg U52509 ( .A(n38539), .B(n38540), .X(n45615) );
  nand_x1_sg U52510 ( .A(w_3[1]), .B(n57569), .X(n38540) );
  nand_x1_sg U52511 ( .A(n38519), .B(n38520), .X(n45605) );
  nand_x1_sg U52512 ( .A(w_3[0]), .B(n57620), .X(n38520) );
  nand_x1_sg U52513 ( .A(n38531), .B(n38532), .X(n45611) );
  nand_x1_sg U52514 ( .A(w_2[19]), .B(n57566), .X(n38532) );
  nand_x1_sg U52515 ( .A(n38533), .B(n38534), .X(n45612) );
  nand_x1_sg U52516 ( .A(w_2[18]), .B(n57566), .X(n38534) );
  nand_x1_sg U52517 ( .A(n38505), .B(n38506), .X(n45598) );
  nand_x1_sg U52518 ( .A(w_2[17]), .B(n57621), .X(n38506) );
  nand_x1_sg U52519 ( .A(n38511), .B(n38512), .X(n45601) );
  nand_x1_sg U52520 ( .A(w_2[16]), .B(n57562), .X(n38512) );
  nand_x1_sg U52521 ( .A(n38517), .B(n38518), .X(n45604) );
  nand_x1_sg U52522 ( .A(w_2[15]), .B(n57568), .X(n38518) );
  nand_x1_sg U52523 ( .A(n38503), .B(n38504), .X(n45597) );
  nand_x1_sg U52524 ( .A(w_2[14]), .B(n57615), .X(n38504) );
  nand_x1_sg U52525 ( .A(n38527), .B(n38528), .X(n45609) );
  nand_x1_sg U52526 ( .A(w_2[13]), .B(n57615), .X(n38528) );
  nand_x1_sg U52527 ( .A(n38529), .B(n38530), .X(n45610) );
  nand_x1_sg U52528 ( .A(w_2[12]), .B(n57563), .X(n38530) );
  nand_x1_sg U52529 ( .A(n38521), .B(n38522), .X(n45606) );
  nand_x1_sg U52530 ( .A(w_2[11]), .B(n57569), .X(n38522) );
  nand_x1_sg U52531 ( .A(n38523), .B(n38524), .X(n45607) );
  nand_x1_sg U52532 ( .A(w_2[10]), .B(n57620), .X(n38524) );
  nand_x1_sg U52533 ( .A(n38569), .B(n38570), .X(n45630) );
  nand_x1_sg U52534 ( .A(w_2[9]), .B(n57565), .X(n38570) );
  nand_x1_sg U52535 ( .A(n38571), .B(n38572), .X(n45631) );
  nand_x1_sg U52536 ( .A(w_2[8]), .B(n57565), .X(n38572) );
  nand_x1_sg U52537 ( .A(n38563), .B(n38564), .X(n45627) );
  nand_x1_sg U52538 ( .A(w_2[7]), .B(n57565), .X(n38564) );
  nand_x1_sg U52539 ( .A(n38565), .B(n38566), .X(n45628) );
  nand_x1_sg U52540 ( .A(w_2[6]), .B(n57565), .X(n38566) );
  nand_x1_sg U52541 ( .A(n38579), .B(n38580), .X(n45635) );
  nand_x1_sg U52542 ( .A(w_2[5]), .B(n57566), .X(n38580) );
  nand_x1_sg U52543 ( .A(n38573), .B(n38574), .X(n45632) );
  nand_x1_sg U52544 ( .A(w_2[4]), .B(n57565), .X(n38574) );
  nand_x1_sg U52545 ( .A(n38561), .B(n38562), .X(n45626) );
  nand_x1_sg U52546 ( .A(w_2[3]), .B(n57565), .X(n38562) );
  nand_x1_sg U52547 ( .A(n38559), .B(n38560), .X(n45625) );
  nand_x1_sg U52548 ( .A(w_2[2]), .B(n57565), .X(n38560) );
  nand_x1_sg U52549 ( .A(n38555), .B(n38556), .X(n45623) );
  nand_x1_sg U52550 ( .A(w_2[1]), .B(n57564), .X(n38556) );
  nand_x1_sg U52551 ( .A(n38557), .B(n38558), .X(n45624) );
  nand_x1_sg U52552 ( .A(w_2[0]), .B(n57564), .X(n38558) );
  nand_x1_sg U52553 ( .A(n38549), .B(n38550), .X(n45620) );
  nand_x1_sg U52554 ( .A(w_1[19]), .B(n57564), .X(n38550) );
  nand_x1_sg U52555 ( .A(n38551), .B(n38552), .X(n45621) );
  nand_x1_sg U52556 ( .A(w_1[18]), .B(n57564), .X(n38552) );
  nand_x1_sg U52557 ( .A(n38567), .B(n38568), .X(n45629) );
  nand_x1_sg U52558 ( .A(w_1[17]), .B(n57565), .X(n38568) );
  nand_x1_sg U52559 ( .A(n38547), .B(n38548), .X(n45619) );
  nand_x1_sg U52560 ( .A(w_1[16]), .B(n57564), .X(n38548) );
  nand_x1_sg U52561 ( .A(n38553), .B(n38554), .X(n45622) );
  nand_x1_sg U52562 ( .A(w_1[15]), .B(n57564), .X(n38554) );
  nand_x1_sg U52563 ( .A(n38545), .B(n38546), .X(n45618) );
  nand_x1_sg U52564 ( .A(w_1[14]), .B(n57564), .X(n38546) );
  nand_x1_sg U52565 ( .A(n39673), .B(n39674), .X(n46182) );
  nand_x1_sg U52566 ( .A(w_1[13]), .B(n57564), .X(n39674) );
  nand_x1_sg U52567 ( .A(n39679), .B(n39680), .X(n46185) );
  nand_x1_sg U52568 ( .A(w_1[12]), .B(n57606), .X(n39680) );
  nand_x1_sg U52569 ( .A(n39241), .B(n39242), .X(n45966) );
  nand_x1_sg U52570 ( .A(w_1[11]), .B(n57598), .X(n39242) );
  nand_x1_sg U52571 ( .A(n39259), .B(n39260), .X(n45975) );
  nand_x1_sg U52572 ( .A(w_1[10]), .B(n57599), .X(n39260) );
  nand_x1_sg U52573 ( .A(n39601), .B(n39602), .X(n46146) );
  nand_x1_sg U52574 ( .A(w_1[9]), .B(n57604), .X(n39602) );
  nand_x1_sg U52575 ( .A(n39691), .B(n39692), .X(n46191) );
  nand_x1_sg U52576 ( .A(w_1[8]), .B(n57606), .X(n39692) );
  nand_x1_sg U52577 ( .A(n39685), .B(n39686), .X(n46188) );
  nand_x1_sg U52578 ( .A(w_1[7]), .B(n57606), .X(n39686) );
  nand_x1_sg U52579 ( .A(n39325), .B(n39326), .X(n46008) );
  nand_x1_sg U52580 ( .A(w_1[6]), .B(n57623), .X(n39326) );
  nand_x1_sg U52581 ( .A(n38483), .B(n38484), .X(n45587) );
  nand_x1_sg U52582 ( .A(w_1[5]), .B(n57563), .X(n38484) );
  nand_x1_sg U52583 ( .A(n38467), .B(n38468), .X(n45579) );
  nand_x1_sg U52584 ( .A(w_1[4]), .B(n57562), .X(n38468) );
  nand_x1_sg U52585 ( .A(n39577), .B(n39578), .X(n46134) );
  nand_x1_sg U52586 ( .A(w_1[3]), .B(n57602), .X(n39578) );
  nand_x1_sg U52587 ( .A(n38461), .B(n38462), .X(n45576) );
  nand_x1_sg U52588 ( .A(w_1[2]), .B(n57562), .X(n38462) );
  nand_x1_sg U52589 ( .A(n38469), .B(n38470), .X(n45580) );
  nand_x1_sg U52590 ( .A(w_1[1]), .B(n57563), .X(n38470) );
  nand_x1_sg U52591 ( .A(n39331), .B(n39332), .X(n46011) );
  nand_x1_sg U52592 ( .A(w_1[0]), .B(n57620), .X(n39332) );
  nand_x1_sg U52593 ( .A(n38463), .B(n38464), .X(n45577) );
  nand_x1_sg U52594 ( .A(w_0[19]), .B(n57562), .X(n38464) );
  nand_x1_sg U52595 ( .A(n38465), .B(n38466), .X(n45578) );
  nand_x1_sg U52596 ( .A(w_0[18]), .B(n57562), .X(n38466) );
  nand_x1_sg U52597 ( .A(n38475), .B(n38476), .X(n45583) );
  nand_x1_sg U52598 ( .A(w_0[17]), .B(n57563), .X(n38476) );
  nand_x1_sg U52599 ( .A(n38477), .B(n38478), .X(n45584) );
  nand_x1_sg U52600 ( .A(w_0[16]), .B(n57563), .X(n38478) );
  nand_x1_sg U52601 ( .A(n38473), .B(n38474), .X(n45582) );
  nand_x1_sg U52602 ( .A(w_0[15]), .B(n57563), .X(n38474) );
  nand_x1_sg U52603 ( .A(n38485), .B(n38486), .X(n45588) );
  nand_x1_sg U52604 ( .A(w_0[14]), .B(n57563), .X(n38486) );
  nand_x1_sg U52605 ( .A(n38513), .B(n38514), .X(n45602) );
  nand_x1_sg U52606 ( .A(w_0[13]), .B(n57567), .X(n38514) );
  nand_x1_sg U52607 ( .A(n38515), .B(n38516), .X(n45603) );
  nand_x1_sg U52608 ( .A(w_0[12]), .B(n57615), .X(n38516) );
  nand_x1_sg U52609 ( .A(n38507), .B(n38508), .X(n45599) );
  nand_x1_sg U52610 ( .A(w_0[11]), .B(n57628), .X(n38508) );
  nand_x1_sg U52611 ( .A(n38509), .B(n38510), .X(n45600) );
  nand_x1_sg U52612 ( .A(w_0[10]), .B(n57563), .X(n38510) );
  nand_x1_sg U52613 ( .A(n38493), .B(n38494), .X(n45592) );
  nand_x1_sg U52614 ( .A(w_0[9]), .B(n57622), .X(n38494) );
  nand_x1_sg U52615 ( .A(n38495), .B(n38496), .X(n45593) );
  nand_x1_sg U52616 ( .A(w_0[8]), .B(n57623), .X(n38496) );
  nand_x1_sg U52617 ( .A(n38487), .B(n38488), .X(n45589) );
  nand_x1_sg U52618 ( .A(w_0[7]), .B(n57630), .X(n38488) );
  nand_x1_sg U52619 ( .A(n38489), .B(n38490), .X(n45590) );
  nand_x1_sg U52620 ( .A(w_0[6]), .B(n57600), .X(n38490) );
  nand_x1_sg U52621 ( .A(n38497), .B(n38498), .X(n45594) );
  nand_x1_sg U52622 ( .A(w_0[5]), .B(n57618), .X(n38498) );
  nand_x1_sg U52623 ( .A(n39355), .B(n39356), .X(n46023) );
  nand_x1_sg U52624 ( .A(w_0[4]), .B(n57617), .X(n39356) );
  nand_x1_sg U52625 ( .A(n38499), .B(n38500), .X(n45595) );
  nand_x1_sg U52626 ( .A(w_0[3]), .B(n57616), .X(n38500) );
  nand_x1_sg U52627 ( .A(n38501), .B(n38502), .X(n45596) );
  nand_x1_sg U52628 ( .A(w_0[2]), .B(n57617), .X(n38502) );
  nand_x1_sg U52629 ( .A(n38695), .B(n38696), .X(n45693) );
  nand_x1_sg U52630 ( .A(w_0[1]), .B(n57570), .X(n38696) );
  nand_x1_sg U52631 ( .A(n38671), .B(n38672), .X(n45681) );
  nand_x1_sg U52632 ( .A(w_0[0]), .B(n57567), .X(n38672) );
  nand_x1_sg U52633 ( .A(n38677), .B(n38678), .X(n45684) );
  nand_x1_sg U52634 ( .A(i_15[19]), .B(n57566), .X(n38678) );
  nand_x1_sg U52635 ( .A(n38683), .B(n38684), .X(n45687) );
  nand_x1_sg U52636 ( .A(i_15[18]), .B(n57615), .X(n38684) );
  nand_x1_sg U52637 ( .A(n38705), .B(n38706), .X(n45698) );
  nand_x1_sg U52638 ( .A(i_15[17]), .B(n57571), .X(n38706) );
  nand_x1_sg U52639 ( .A(n38707), .B(n38708), .X(n45699) );
  nand_x1_sg U52640 ( .A(i_15[16]), .B(n57571), .X(n38708) );
  nand_x1_sg U52641 ( .A(n38699), .B(n38700), .X(n45695) );
  nand_x1_sg U52642 ( .A(i_15[15]), .B(n57570), .X(n38700) );
  nand_x1_sg U52643 ( .A(n38701), .B(n38702), .X(n45696) );
  nand_x1_sg U52644 ( .A(i_15[14]), .B(n57570), .X(n38702) );
  nand_x1_sg U52645 ( .A(n38679), .B(n38680), .X(n45685) );
  nand_x1_sg U52646 ( .A(i_15[13]), .B(n57564), .X(n38680) );
  nand_x1_sg U52647 ( .A(n38681), .B(n38682), .X(n45686) );
  nand_x1_sg U52648 ( .A(i_15[12]), .B(n57567), .X(n38682) );
  nand_x1_sg U52649 ( .A(n38673), .B(n38674), .X(n45682) );
  nand_x1_sg U52650 ( .A(i_15[11]), .B(n57566), .X(n38674) );
  nand_x1_sg U52651 ( .A(n38675), .B(n38676), .X(n45683) );
  nand_x1_sg U52652 ( .A(i_15[10]), .B(n57615), .X(n38676) );
  nand_x1_sg U52653 ( .A(n38691), .B(n38692), .X(n45691) );
  nand_x1_sg U52654 ( .A(i_15[9]), .B(n57570), .X(n38692) );
  nand_x1_sg U52655 ( .A(n38693), .B(n38694), .X(n45692) );
  nand_x1_sg U52656 ( .A(i_15[8]), .B(n57570), .X(n38694) );
  nand_x1_sg U52657 ( .A(n38685), .B(n38686), .X(n45688) );
  nand_x1_sg U52658 ( .A(i_15[7]), .B(n57570), .X(n38686) );
  nand_x1_sg U52659 ( .A(n38687), .B(n38688), .X(n45689) );
  nand_x1_sg U52660 ( .A(i_15[6]), .B(n57570), .X(n38688) );
  nand_x1_sg U52661 ( .A(n38525), .B(n38526), .X(n45608) );
  nand_x1_sg U52662 ( .A(i_15[5]), .B(n57562), .X(n38526) );
  nand_x1_sg U52663 ( .A(n38491), .B(n38492), .X(n45591) );
  nand_x1_sg U52664 ( .A(i_15[4]), .B(n57625), .X(n38492) );
  nand_x1_sg U52665 ( .A(n38449), .B(n38450), .X(n45570) );
  nand_x1_sg U52666 ( .A(i_15[3]), .B(n57562), .X(n38450) );
  nand_x1_sg U52667 ( .A(n38451), .B(n38452), .X(n45571) );
  nand_x1_sg U52668 ( .A(i_15[2]), .B(n57562), .X(n38452) );
  nand_x1_sg U52669 ( .A(n38591), .B(n38592), .X(n45641) );
  nand_x1_sg U52670 ( .A(i_15[1]), .B(n57566), .X(n38592) );
  nand_x1_sg U52671 ( .A(n38709), .B(n38710), .X(n45700) );
  nand_x1_sg U52672 ( .A(i_15[0]), .B(n57571), .X(n38710) );
  nand_x1_sg U52673 ( .A(n38727), .B(n38728), .X(n45709) );
  nand_x1_sg U52674 ( .A(i_14[19]), .B(n57572), .X(n38728) );
  nand_x1_sg U52675 ( .A(n38447), .B(n38448), .X(n45569) );
  nand_x1_sg U52676 ( .A(i_14[18]), .B(n57563), .X(n38448) );
  nand_x1_sg U52677 ( .A(n38717), .B(n38718), .X(n45704) );
  nand_x1_sg U52678 ( .A(i_14[17]), .B(n57571), .X(n38718) );
  nand_x1_sg U52679 ( .A(n38703), .B(n38704), .X(n45697) );
  nand_x1_sg U52680 ( .A(i_14[16]), .B(n57571), .X(n38704) );
  nand_x1_sg U52681 ( .A(n38719), .B(n38720), .X(n45705) );
  nand_x1_sg U52682 ( .A(i_14[15]), .B(n57571), .X(n38720) );
  nand_x1_sg U52683 ( .A(n38721), .B(n38722), .X(n45706) );
  nand_x1_sg U52684 ( .A(i_14[14]), .B(n57572), .X(n38722) );
  nand_x1_sg U52685 ( .A(n38713), .B(n38714), .X(n45702) );
  nand_x1_sg U52686 ( .A(i_14[13]), .B(n57571), .X(n38714) );
  nand_x1_sg U52687 ( .A(n38715), .B(n38716), .X(n45703) );
  nand_x1_sg U52688 ( .A(i_14[12]), .B(n57571), .X(n38716) );
  nand_x1_sg U52689 ( .A(n38711), .B(n38712), .X(n45701) );
  nand_x1_sg U52690 ( .A(i_14[11]), .B(n57571), .X(n38712) );
  nand_x1_sg U52691 ( .A(n38697), .B(n38698), .X(n45694) );
  nand_x1_sg U52692 ( .A(i_14[10]), .B(n57570), .X(n38698) );
  nand_x1_sg U52693 ( .A(n38597), .B(n38598), .X(n45644) );
  nand_x1_sg U52694 ( .A(i_14[9]), .B(n57567), .X(n38598) );
  nand_x1_sg U52695 ( .A(n38585), .B(n38586), .X(n45638) );
  nand_x1_sg U52696 ( .A(i_14[8]), .B(n57566), .X(n38586) );
  nand_x1_sg U52697 ( .A(n38599), .B(n38600), .X(n45645) );
  nand_x1_sg U52698 ( .A(i_14[7]), .B(n57567), .X(n38600) );
  nand_x1_sg U52699 ( .A(n38605), .B(n38606), .X(n45648) );
  nand_x1_sg U52700 ( .A(i_14[6]), .B(n57567), .X(n38606) );
  nand_x1_sg U52701 ( .A(n38607), .B(n38608), .X(n45649) );
  nand_x1_sg U52702 ( .A(i_14[5]), .B(n57567), .X(n38608) );
  nand_x1_sg U52703 ( .A(n38609), .B(n38610), .X(n45650) );
  nand_x1_sg U52704 ( .A(i_14[4]), .B(n57567), .X(n38610) );
  nand_x1_sg U52705 ( .A(n38601), .B(n38602), .X(n45646) );
  nand_x1_sg U52706 ( .A(i_14[3]), .B(n57567), .X(n38602) );
  nand_x1_sg U52707 ( .A(n38603), .B(n38604), .X(n45647) );
  nand_x1_sg U52708 ( .A(i_14[2]), .B(n57567), .X(n38604) );
  nand_x1_sg U52709 ( .A(n38581), .B(n38582), .X(n45636) );
  nand_x1_sg U52710 ( .A(i_14[1]), .B(n57566), .X(n38582) );
  nand_x1_sg U52711 ( .A(n38583), .B(n38584), .X(n45637) );
  nand_x1_sg U52712 ( .A(i_14[0]), .B(n57566), .X(n38584) );
  nand_x1_sg U52713 ( .A(n38575), .B(n38576), .X(n45633) );
  nand_x1_sg U52714 ( .A(i_13[19]), .B(n57565), .X(n38576) );
  nand_x1_sg U52715 ( .A(n38577), .B(n38578), .X(n45634) );
  nand_x1_sg U52716 ( .A(i_13[18]), .B(n57566), .X(n38578) );
  nand_x1_sg U52717 ( .A(n38593), .B(n38594), .X(n45642) );
  nand_x1_sg U52718 ( .A(i_13[17]), .B(n57566), .X(n38594) );
  nand_x1_sg U52719 ( .A(n38595), .B(n38596), .X(n45643) );
  nand_x1_sg U52720 ( .A(i_13[16]), .B(n57567), .X(n38596) );
  nand_x1_sg U52721 ( .A(n38587), .B(n38588), .X(n45639) );
  nand_x1_sg U52722 ( .A(i_13[15]), .B(n57566), .X(n38588) );
  nand_x1_sg U52723 ( .A(n38589), .B(n38590), .X(n45640) );
  nand_x1_sg U52724 ( .A(i_13[14]), .B(n57566), .X(n38590) );
  nand_x1_sg U52725 ( .A(n38637), .B(n38638), .X(n45664) );
  nand_x1_sg U52726 ( .A(i_13[13]), .B(n57569), .X(n38638) );
  nand_x1_sg U52727 ( .A(n38639), .B(n38640), .X(n45665) );
  nand_x1_sg U52728 ( .A(i_13[12]), .B(n57569), .X(n38640) );
  nand_x1_sg U52729 ( .A(n38631), .B(n38632), .X(n45661) );
  nand_x1_sg U52730 ( .A(i_13[11]), .B(n57569), .X(n38632) );
  nand_x1_sg U52731 ( .A(n38633), .B(n38634), .X(n45662) );
  nand_x1_sg U52732 ( .A(i_13[10]), .B(n57569), .X(n38634) );
  nand_x1_sg U52733 ( .A(n38665), .B(n38666), .X(n45678) );
  nand_x1_sg U52734 ( .A(i_13[9]), .B(n57564), .X(n38666) );
  nand_x1_sg U52735 ( .A(n38629), .B(n38630), .X(n45660) );
  nand_x1_sg U52736 ( .A(i_13[8]), .B(n57568), .X(n38630) );
  nand_x1_sg U52737 ( .A(n38667), .B(n38668), .X(n45679) );
  nand_x1_sg U52738 ( .A(i_13[7]), .B(n57565), .X(n38668) );
  nand_x1_sg U52739 ( .A(n38669), .B(n38670), .X(n45680) );
  nand_x1_sg U52740 ( .A(i_13[6]), .B(n57564), .X(n38670) );
  nand_x1_sg U52741 ( .A(n38619), .B(n38620), .X(n45655) );
  nand_x1_sg U52742 ( .A(i_13[5]), .B(n57568), .X(n38620) );
  nand_x1_sg U52743 ( .A(n38621), .B(n38622), .X(n45656) );
  nand_x1_sg U52744 ( .A(i_13[4]), .B(n57568), .X(n38622) );
  nand_x1_sg U52745 ( .A(n38613), .B(n38614), .X(n45652) );
  nand_x1_sg U52746 ( .A(i_13[3]), .B(n57568), .X(n38614) );
  nand_x1_sg U52747 ( .A(n38615), .B(n38616), .X(n45653) );
  nand_x1_sg U52748 ( .A(i_13[2]), .B(n57568), .X(n38616) );
  nand_x1_sg U52749 ( .A(n38623), .B(n38624), .X(n45657) );
  nand_x1_sg U52750 ( .A(i_13[1]), .B(n57568), .X(n38624) );
  nand_x1_sg U52751 ( .A(n38611), .B(n38612), .X(n45651) );
  nand_x1_sg U52752 ( .A(i_13[0]), .B(n57567), .X(n38612) );
  nand_x1_sg U52753 ( .A(n38625), .B(n38626), .X(n45658) );
  nand_x1_sg U52754 ( .A(i_12[19]), .B(n57568), .X(n38626) );
  nand_x1_sg U52755 ( .A(n38627), .B(n38628), .X(n45659) );
  nand_x1_sg U52756 ( .A(i_12[18]), .B(n57568), .X(n38628) );
  nand_x1_sg U52757 ( .A(n39187), .B(n39188), .X(n45939) );
  nand_x1_sg U52758 ( .A(i_12[17]), .B(n57595), .X(n39188) );
  nand_x1_sg U52759 ( .A(n39319), .B(n39320), .X(n46005) );
  nand_x1_sg U52760 ( .A(i_12[16]), .B(n57620), .X(n39320) );
  nand_x1_sg U52761 ( .A(n38443), .B(n38444), .X(n45567) );
  nand_x1_sg U52762 ( .A(i_12[15]), .B(n57623), .X(n38444) );
  nand_x1_sg U52763 ( .A(n39313), .B(n39314), .X(n46002) );
  nand_x1_sg U52764 ( .A(i_12[14]), .B(n57600), .X(n39314) );
  nand_x1_sg U52765 ( .A(n39373), .B(n39374), .X(n46032) );
  nand_x1_sg U52766 ( .A(i_12[13]), .B(n38414), .X(n39374) );
  nand_x1_sg U52767 ( .A(n39409), .B(n39410), .X(n46050) );
  nand_x1_sg U52768 ( .A(i_12[12]), .B(n57621), .X(n39410) );
  nand_x1_sg U52769 ( .A(n38441), .B(n38442), .X(n45566) );
  nand_x1_sg U52770 ( .A(i_12[11]), .B(n57615), .X(n38442) );
  nand_x1_sg U52771 ( .A(n38439), .B(n38440), .X(n45565) );
  nand_x1_sg U52772 ( .A(i_12[10]), .B(n57563), .X(n38440) );
  nand_x1_sg U52773 ( .A(n39301), .B(n39302), .X(n45996) );
  nand_x1_sg U52774 ( .A(i_12[9]), .B(n57624), .X(n39302) );
  nand_x1_sg U52775 ( .A(n39307), .B(n39308), .X(n45999) );
  nand_x1_sg U52776 ( .A(i_12[8]), .B(n57600), .X(n39308) );
  nand_x1_sg U52777 ( .A(n38435), .B(n38436), .X(n45563) );
  nand_x1_sg U52778 ( .A(i_12[7]), .B(n57625), .X(n38436) );
  nand_x1_sg U52779 ( .A(n38433), .B(n38434), .X(n45562) );
  nand_x1_sg U52780 ( .A(i_12[6]), .B(n57618), .X(n38434) );
  nand_x1_sg U52781 ( .A(n39295), .B(n39296), .X(n45993) );
  nand_x1_sg U52782 ( .A(i_12[5]), .B(n57619), .X(n39296) );
  nand_x1_sg U52783 ( .A(n39253), .B(n39254), .X(n45972) );
  nand_x1_sg U52784 ( .A(i_12[4]), .B(n57599), .X(n39254) );
  nand_x1_sg U52785 ( .A(n38437), .B(n38438), .X(n45564) );
  nand_x1_sg U52786 ( .A(i_12[3]), .B(n57619), .X(n38438) );
  nand_x1_sg U52787 ( .A(n39289), .B(n39290), .X(n45990) );
  nand_x1_sg U52788 ( .A(i_12[2]), .B(n57616), .X(n39290) );
  nand_x1_sg U52789 ( .A(n39439), .B(n39440), .X(n46065) );
  nand_x1_sg U52790 ( .A(i_12[1]), .B(n57600), .X(n39440) );
  nand_x1_sg U52791 ( .A(n39445), .B(n39446), .X(n46068) );
  nand_x1_sg U52792 ( .A(i_12[0]), .B(n57620), .X(n39446) );
  nand_x1_sg U52793 ( .A(n39493), .B(n39494), .X(n46092) );
  nand_x1_sg U52794 ( .A(i_11[19]), .B(n57569), .X(n39494) );
  nand_x1_sg U52795 ( .A(n39499), .B(n39500), .X(n46095) );
  nand_x1_sg U52796 ( .A(i_11[18]), .B(n57562), .X(n39500) );
  nand_x1_sg U52797 ( .A(n39451), .B(n39452), .X(n46071) );
  nand_x1_sg U52798 ( .A(i_11[17]), .B(n57621), .X(n39452) );
  nand_x1_sg U52799 ( .A(n39433), .B(n39434), .X(n46062) );
  nand_x1_sg U52800 ( .A(i_11[16]), .B(n57600), .X(n39434) );
  nand_x1_sg U52801 ( .A(n39505), .B(n39506), .X(n46098) );
  nand_x1_sg U52802 ( .A(i_11[15]), .B(n57617), .X(n39506) );
  nand_x1_sg U52803 ( .A(n39481), .B(n39482), .X(n46086) );
  nand_x1_sg U52804 ( .A(i_11[14]), .B(n57624), .X(n39482) );
  nand_x1_sg U52805 ( .A(n39343), .B(n39344), .X(n46017) );
  nand_x1_sg U52806 ( .A(i_11[13]), .B(n57617), .X(n39344) );
  nand_x1_sg U52807 ( .A(n39415), .B(n39416), .X(n46053) );
  nand_x1_sg U52808 ( .A(i_11[12]), .B(n57619), .X(n39416) );
  nand_x1_sg U52809 ( .A(n38459), .B(n38460), .X(n45575) );
  nand_x1_sg U52810 ( .A(i_11[11]), .B(n57562), .X(n38460) );
  nand_x1_sg U52811 ( .A(n39337), .B(n39338), .X(n46014) );
  nand_x1_sg U52812 ( .A(i_11[10]), .B(n57624), .X(n39338) );
  nand_x1_sg U52813 ( .A(n39517), .B(n39518), .X(n46104) );
  nand_x1_sg U52814 ( .A(i_11[9]), .B(n57617), .X(n39518) );
  nand_x1_sg U52815 ( .A(n39523), .B(n39524), .X(n46107) );
  nand_x1_sg U52816 ( .A(i_11[8]), .B(n57562), .X(n39524) );
  nand_x1_sg U52817 ( .A(n39511), .B(n39512), .X(n46101) );
  nand_x1_sg U52818 ( .A(i_11[7]), .B(n57628), .X(n39512) );
  nand_x1_sg U52819 ( .A(n39421), .B(n39422), .X(n46056) );
  nand_x1_sg U52820 ( .A(i_11[6]), .B(n57616), .X(n39422) );
  nand_x1_sg U52821 ( .A(n38431), .B(n38432), .X(n45561) );
  nand_x1_sg U52822 ( .A(i_11[5]), .B(n57563), .X(n38432) );
  nand_x1_sg U52823 ( .A(n38935), .B(n38936), .X(n45813) );
  nand_x1_sg U52824 ( .A(i_11[4]), .B(n57581), .X(n38936) );
  nand_x1_sg U52825 ( .A(n38427), .B(n38428), .X(n45559) );
  nand_x1_sg U52826 ( .A(i_11[3]), .B(n57624), .X(n38428) );
  nand_x1_sg U52827 ( .A(n39109), .B(n39110), .X(n45900) );
  nand_x1_sg U52828 ( .A(i_11[2]), .B(n57591), .X(n39110) );
  nand_x1_sg U52829 ( .A(n39115), .B(n39116), .X(n45903) );
  nand_x1_sg U52830 ( .A(i_11[1]), .B(n57591), .X(n39116) );
  nand_x1_sg U52831 ( .A(n39133), .B(n39134), .X(n45912) );
  nand_x1_sg U52832 ( .A(i_11[0]), .B(n57592), .X(n39134) );
  nand_x1_sg U52833 ( .A(n38429), .B(n38430), .X(n45560) );
  nand_x1_sg U52834 ( .A(i_10[19]), .B(n57624), .X(n38430) );
  nand_x1_sg U52835 ( .A(n39139), .B(n39140), .X(n45915) );
  nand_x1_sg U52836 ( .A(i_10[18]), .B(n57593), .X(n39140) );
  nand_x1_sg U52837 ( .A(n39643), .B(n39644), .X(n46167) );
  nand_x1_sg U52838 ( .A(i_10[17]), .B(n57605), .X(n39644) );
  nand_x1_sg U52839 ( .A(n38653), .B(n38654), .X(n45672) );
  nand_x1_sg U52840 ( .A(i_10[16]), .B(n57615), .X(n38654) );
  nand_x1_sg U52841 ( .A(n38423), .B(n38424), .X(n45557) );
  nand_x1_sg U52842 ( .A(i_10[15]), .B(n57600), .X(n38424) );
  nand_x1_sg U52843 ( .A(n38421), .B(n38422), .X(n45556) );
  nand_x1_sg U52844 ( .A(i_10[14]), .B(n57615), .X(n38422) );
  nand_x1_sg U52845 ( .A(n39637), .B(n39638), .X(n46164) );
  nand_x1_sg U52846 ( .A(i_10[13]), .B(n57604), .X(n39638) );
  nand_x1_sg U52847 ( .A(n38659), .B(n38660), .X(n45675) );
  nand_x1_sg U52848 ( .A(i_10[12]), .B(n57568), .X(n38660) );
  nand_x1_sg U52849 ( .A(n38425), .B(n38426), .X(n45558) );
  nand_x1_sg U52850 ( .A(i_10[11]), .B(n57624), .X(n38426) );
  nand_x1_sg U52851 ( .A(n39625), .B(n39626), .X(n46158) );
  nand_x1_sg U52852 ( .A(i_10[10]), .B(n57604), .X(n39626) );
  nand_x1_sg U52853 ( .A(n39151), .B(n39152), .X(n45921) );
  nand_x1_sg U52854 ( .A(i_10[9]), .B(n57593), .X(n39152) );
  nand_x1_sg U52855 ( .A(n39157), .B(n39158), .X(n45924) );
  nand_x1_sg U52856 ( .A(i_10[8]), .B(n57594), .X(n39158) );
  nand_x1_sg U52857 ( .A(n38419), .B(n38420), .X(n45555) );
  nand_x1_sg U52858 ( .A(i_10[7]), .B(n57618), .X(n38420) );
  nand_x1_sg U52859 ( .A(n39175), .B(n39176), .X(n45933) );
  nand_x1_sg U52860 ( .A(i_10[6]), .B(n57595), .X(n39176) );
  nand_x1_sg U52861 ( .A(n39145), .B(n39146), .X(n45918) );
  nand_x1_sg U52862 ( .A(i_10[5]), .B(n57593), .X(n39146) );
  nand_x1_sg U52863 ( .A(n39169), .B(n39170), .X(n45930) );
  nand_x1_sg U52864 ( .A(i_10[4]), .B(n57594), .X(n39170) );
  nand_x1_sg U52865 ( .A(n39163), .B(n39164), .X(n45927) );
  nand_x1_sg U52866 ( .A(i_10[3]), .B(n57594), .X(n39164) );
  nand_x1_sg U52867 ( .A(n39181), .B(n39182), .X(n45936) );
  nand_x1_sg U52868 ( .A(i_10[2]), .B(n57595), .X(n39182) );
  nand_x1_sg U52869 ( .A(n38617), .B(n38618), .X(n45654) );
  nand_x1_sg U52870 ( .A(i_10[1]), .B(n57568), .X(n38618) );
  nand_x1_sg U52871 ( .A(n39071), .B(n39072), .X(n45881) );
  nand_x1_sg U52872 ( .A(i_10[0]), .B(n57589), .X(n39072) );
  nand_x1_sg U52873 ( .A(n39085), .B(n39086), .X(n45888) );
  nand_x1_sg U52874 ( .A(i_9[19]), .B(n57590), .X(n39086) );
  nand_x1_sg U52875 ( .A(n39091), .B(n39092), .X(n45891) );
  nand_x1_sg U52876 ( .A(i_9[18]), .B(n57590), .X(n39092) );
  nand_x1_sg U52877 ( .A(n39073), .B(n39074), .X(n45882) );
  nand_x1_sg U52878 ( .A(i_9[17]), .B(n57589), .X(n39074) );
  nand_x1_sg U52879 ( .A(n38941), .B(n38942), .X(n45816) );
  nand_x1_sg U52880 ( .A(i_9[16]), .B(n57582), .X(n38942) );
  nand_x1_sg U52881 ( .A(n39103), .B(n39104), .X(n45897) );
  nand_x1_sg U52882 ( .A(i_9[15]), .B(n57591), .X(n39104) );
  nand_x1_sg U52883 ( .A(n39079), .B(n39080), .X(n45885) );
  nand_x1_sg U52884 ( .A(i_9[14]), .B(n57589), .X(n39080) );
  nand_x1_sg U52885 ( .A(n39127), .B(n39128), .X(n45909) );
  nand_x1_sg U52886 ( .A(i_9[13]), .B(n57592), .X(n39128) );
  nand_x1_sg U52887 ( .A(n39217), .B(n39218), .X(n45954) );
  nand_x1_sg U52888 ( .A(i_9[12]), .B(n57597), .X(n39218) );
  nand_x1_sg U52889 ( .A(n39223), .B(n39224), .X(n45957) );
  nand_x1_sg U52890 ( .A(i_9[11]), .B(n57597), .X(n39224) );
  nand_x1_sg U52891 ( .A(n39229), .B(n39230), .X(n45960) );
  nand_x1_sg U52892 ( .A(i_9[10]), .B(n57598), .X(n39230) );
  nand_x1_sg U52893 ( .A(n38471), .B(n38472), .X(n45581) );
  nand_x1_sg U52894 ( .A(i_9[9]), .B(n57563), .X(n38472) );
  nand_x1_sg U52895 ( .A(n38839), .B(n38840), .X(n45765) );
  nand_x1_sg U52896 ( .A(i_9[8]), .B(n57577), .X(n38840) );
  nand_x1_sg U52897 ( .A(n38929), .B(n38930), .X(n45810) );
  nand_x1_sg U52898 ( .A(i_9[7]), .B(n57581), .X(n38930) );
  nand_x1_sg U52899 ( .A(n39097), .B(n39098), .X(n45894) );
  nand_x1_sg U52900 ( .A(i_9[6]), .B(n57590), .X(n39098) );
  nand_x1_sg U52901 ( .A(n38827), .B(n38828), .X(n45759) );
  nand_x1_sg U52902 ( .A(i_9[5]), .B(n57576), .X(n38828) );
  nand_x1_sg U52903 ( .A(n38833), .B(n38834), .X(n45762) );
  nand_x1_sg U52904 ( .A(i_9[4]), .B(n57577), .X(n38834) );
  nand_x1_sg U52905 ( .A(n39059), .B(n39060), .X(n45875) );
  nand_x1_sg U52906 ( .A(i_9[3]), .B(n57588), .X(n39060) );
  nand_x1_sg U52907 ( .A(n38877), .B(n38878), .X(n45784) );
  nand_x1_sg U52908 ( .A(i_9[2]), .B(n57578), .X(n38878) );
  nand_x1_sg U52909 ( .A(n38803), .B(n38804), .X(n45747) );
  nand_x1_sg U52910 ( .A(i_9[1]), .B(n57575), .X(n38804) );
  nand_x1_sg U52911 ( .A(n38809), .B(n38810), .X(n45750) );
  nand_x1_sg U52912 ( .A(i_9[0]), .B(n57575), .X(n38810) );
  nand_x1_sg U52913 ( .A(n38815), .B(n38816), .X(n45753) );
  nand_x1_sg U52914 ( .A(i_8[19]), .B(n57576), .X(n38816) );
  nand_x1_sg U52915 ( .A(n38821), .B(n38822), .X(n45756) );
  nand_x1_sg U52916 ( .A(i_8[18]), .B(n57576), .X(n38822) );
  nand_x1_sg U52917 ( .A(n39361), .B(n39362), .X(n46026) );
  nand_x1_sg U52918 ( .A(i_8[17]), .B(n57625), .X(n39362) );
  nand_x1_sg U52919 ( .A(n39367), .B(n39368), .X(n46029) );
  nand_x1_sg U52920 ( .A(i_8[16]), .B(n57618), .X(n39368) );
  nand_x1_sg U52921 ( .A(n39379), .B(n39380), .X(n46035) );
  nand_x1_sg U52922 ( .A(i_8[15]), .B(n57562), .X(n39380) );
  nand_x1_sg U52923 ( .A(n39457), .B(n39458), .X(n46074) );
  nand_x1_sg U52924 ( .A(i_8[14]), .B(n57632), .X(n39458) );
  nand_x1_sg U52925 ( .A(n38479), .B(n38480), .X(n45585) );
  nand_x1_sg U52926 ( .A(i_8[13]), .B(n57563), .X(n38480) );
  nand_x1_sg U52927 ( .A(n38481), .B(n38482), .X(n45586) );
  nand_x1_sg U52928 ( .A(i_8[12]), .B(n57563), .X(n38482) );
  nand_x1_sg U52929 ( .A(n39235), .B(n39236), .X(n45963) );
  nand_x1_sg U52930 ( .A(i_8[11]), .B(n57598), .X(n39236) );
  nand_x1_sg U52931 ( .A(n39349), .B(n39350), .X(n46020) );
  nand_x1_sg U52932 ( .A(i_8[10]), .B(n57622), .X(n39350) );
  nand_x1_sg U52933 ( .A(n38417), .B(n38418), .X(n45554) );
  nand_x1_sg U52934 ( .A(i_8[9]), .B(n57600), .X(n38418) );
  nand_x1_sg U52935 ( .A(n39547), .B(n39548), .X(n46119) );
  nand_x1_sg U52936 ( .A(i_8[8]), .B(n57600), .X(n39548) );
  nand_x1_sg U52937 ( .A(n39121), .B(n39122), .X(n45906) );
  nand_x1_sg U52938 ( .A(i_8[7]), .B(n57592), .X(n39122) );
  nand_x1_sg U52939 ( .A(n38923), .B(n38924), .X(n45807) );
  nand_x1_sg U52940 ( .A(i_8[6]), .B(n57581), .X(n38924) );
  nand_x1_sg U52941 ( .A(n39463), .B(n39464), .X(n46077) );
  nand_x1_sg U52942 ( .A(i_8[5]), .B(n57619), .X(n39464) );
  nand_x1_sg U52943 ( .A(n39469), .B(n39470), .X(n46080) );
  nand_x1_sg U52944 ( .A(i_8[4]), .B(n57616), .X(n39470) );
  nand_x1_sg U52945 ( .A(n39475), .B(n39476), .X(n46083) );
  nand_x1_sg U52946 ( .A(i_8[3]), .B(n57617), .X(n39476) );
  nand_x1_sg U52947 ( .A(n39541), .B(n39542), .X(n46116) );
  nand_x1_sg U52948 ( .A(i_8[2]), .B(n57622), .X(n39542) );
  nand_x1_sg U52949 ( .A(n39649), .B(n39650), .X(n46170) );
  nand_x1_sg U52950 ( .A(i_8[1]), .B(n57605), .X(n39650) );
  nand_x1_sg U52951 ( .A(n39655), .B(n39656), .X(n46173) );
  nand_x1_sg U52952 ( .A(i_8[0]), .B(n57605), .X(n39656) );
  nand_x1_sg U52953 ( .A(n39661), .B(n39662), .X(n46176) );
  nand_x1_sg U52954 ( .A(i_7[19]), .B(n57565), .X(n39662) );
  nand_x1_sg U52955 ( .A(n39667), .B(n39668), .X(n46179) );
  nand_x1_sg U52956 ( .A(i_7[18]), .B(n57562), .X(n39668) );
  nand_x1_sg U52957 ( .A(n39583), .B(n39584), .X(n46137) );
  nand_x1_sg U52958 ( .A(i_7[17]), .B(n57602), .X(n39584) );
  nand_x1_sg U52959 ( .A(n39589), .B(n39590), .X(n46140) );
  nand_x1_sg U52960 ( .A(i_7[16]), .B(n57624), .X(n39590) );
  nand_x1_sg U52961 ( .A(n39607), .B(n39608), .X(n46149) );
  nand_x1_sg U52962 ( .A(i_7[15]), .B(n57603), .X(n39608) );
  nand_x1_sg U52963 ( .A(n39613), .B(n39614), .X(n46152) );
  nand_x1_sg U52964 ( .A(i_7[14]), .B(n57603), .X(n39614) );
  nand_x1_sg U52965 ( .A(n39535), .B(n39536), .X(n46113) );
  nand_x1_sg U52966 ( .A(i_7[13]), .B(n57566), .X(n39536) );
  nand_x1_sg U52967 ( .A(n39553), .B(n39554), .X(n46122) );
  nand_x1_sg U52968 ( .A(i_7[12]), .B(n57601), .X(n39554) );
  nand_x1_sg U52969 ( .A(n39565), .B(n39566), .X(n46128) );
  nand_x1_sg U52970 ( .A(i_7[11]), .B(n57601), .X(n39566) );
  nand_x1_sg U52971 ( .A(n39571), .B(n39572), .X(n46131) );
  nand_x1_sg U52972 ( .A(i_7[10]), .B(n57602), .X(n39572) );
  nand_x1_sg U52973 ( .A(n39247), .B(n39248), .X(n45969) );
  nand_x1_sg U52974 ( .A(i_7[9]), .B(n57599), .X(n39248) );
  nand_x1_sg U52975 ( .A(n39277), .B(n39278), .X(n45984) );
  nand_x1_sg U52976 ( .A(i_7[8]), .B(n57616), .X(n39278) );
  nand_x1_sg U52977 ( .A(n39427), .B(n39428), .X(n46059) );
  nand_x1_sg U52978 ( .A(i_7[7]), .B(n57600), .X(n39428) );
  nand_x1_sg U52979 ( .A(n39487), .B(n39488), .X(n46089) );
  nand_x1_sg U52980 ( .A(i_7[6]), .B(n57624), .X(n39488) );
  nand_x1_sg U52981 ( .A(n38779), .B(n38780), .X(n45735) );
  nand_x1_sg U52982 ( .A(i_7[5]), .B(n57598), .X(n38780) );
  nand_x1_sg U52983 ( .A(n38785), .B(n38786), .X(n45738) );
  nand_x1_sg U52984 ( .A(i_7[4]), .B(n57598), .X(n38786) );
  nand_x1_sg U52985 ( .A(n38457), .B(n38458), .X(n45574) );
  nand_x1_sg U52986 ( .A(i_7[3]), .B(n57562), .X(n38458) );
  nand_x1_sg U52987 ( .A(n38445), .B(n38446), .X(n45568) );
  nand_x1_sg U52988 ( .A(i_7[2]), .B(n57616), .X(n38446) );
  nand_x1_sg U52989 ( .A(n38755), .B(n38756), .X(n45723) );
  nand_x1_sg U52990 ( .A(i_7[1]), .B(n57573), .X(n38756) );
  nand_x1_sg U52991 ( .A(n38761), .B(n38762), .X(n45726) );
  nand_x1_sg U52992 ( .A(i_7[0]), .B(n57574), .X(n38762) );
  nand_x1_sg U52993 ( .A(n38767), .B(n38768), .X(n45729) );
  nand_x1_sg U52994 ( .A(i_6[19]), .B(n57574), .X(n38768) );
  nand_x1_sg U52995 ( .A(n38773), .B(n38774), .X(n45732) );
  nand_x1_sg U52996 ( .A(i_6[18]), .B(n57574), .X(n38774) );
  nand_x1_sg U52997 ( .A(n39619), .B(n39620), .X(n46155) );
  nand_x1_sg U52998 ( .A(i_6[17]), .B(n57603), .X(n39620) );
  nand_x1_sg U52999 ( .A(n39595), .B(n39596), .X(n46143) );
  nand_x1_sg U53000 ( .A(i_6[16]), .B(n57569), .X(n39596) );
  nand_x1_sg U53001 ( .A(n38749), .B(n38750), .X(n45720) );
  nand_x1_sg U53002 ( .A(i_6[15]), .B(n57573), .X(n38750) );
  nand_x1_sg U53003 ( .A(n39283), .B(n39284), .X(n45987) );
  nand_x1_sg U53004 ( .A(i_6[14]), .B(n57617), .X(n39284) );
  nand_x1_sg U53005 ( .A(n38791), .B(n38792), .X(n45741) );
  nand_x1_sg U53006 ( .A(i_6[13]), .B(n57598), .X(n38792) );
  nand_x1_sg U53007 ( .A(n38797), .B(n38798), .X(n45744) );
  nand_x1_sg U53008 ( .A(i_6[12]), .B(n57575), .X(n38798) );
  nand_x1_sg U53009 ( .A(n38453), .B(n38454), .X(n45572) );
  nand_x1_sg U53010 ( .A(i_6[11]), .B(n57562), .X(n38454) );
  nand_x1_sg U53011 ( .A(n38455), .B(n38456), .X(n45573) );
  nand_x1_sg U53012 ( .A(i_6[10]), .B(n57562), .X(n38456) );
  nand_x1_sg U53013 ( .A(n38867), .B(n38868), .X(n45779) );
  nand_x1_sg U53014 ( .A(i_6[9]), .B(n57578), .X(n38868) );
  nand_x1_sg U53015 ( .A(n38869), .B(n38870), .X(n45780) );
  nand_x1_sg U53016 ( .A(i_6[8]), .B(n57578), .X(n38870) );
  nand_x1_sg U53017 ( .A(n38861), .B(n38862), .X(n45776) );
  nand_x1_sg U53018 ( .A(i_6[7]), .B(n57600), .X(n38862) );
  nand_x1_sg U53019 ( .A(n38863), .B(n38864), .X(n45777) );
  nand_x1_sg U53020 ( .A(i_6[6]), .B(n57605), .X(n38864) );
  nand_x1_sg U53021 ( .A(n38879), .B(n38880), .X(n45785) );
  nand_x1_sg U53022 ( .A(i_6[5]), .B(n57578), .X(n38880) );
  nand_x1_sg U53023 ( .A(n38881), .B(n38882), .X(n45786) );
  nand_x1_sg U53024 ( .A(i_6[4]), .B(n57578), .X(n38882) );
  nand_x1_sg U53025 ( .A(n38873), .B(n38874), .X(n45782) );
  nand_x1_sg U53026 ( .A(i_6[3]), .B(n57578), .X(n38874) );
  nand_x1_sg U53027 ( .A(n38875), .B(n38876), .X(n45783) );
  nand_x1_sg U53028 ( .A(i_6[2]), .B(n57578), .X(n38876) );
  nand_x1_sg U53029 ( .A(n38855), .B(n38856), .X(n45773) );
  nand_x1_sg U53030 ( .A(i_6[1]), .B(n57620), .X(n38856) );
  nand_x1_sg U53031 ( .A(n38857), .B(n38858), .X(n45774) );
  nand_x1_sg U53032 ( .A(i_6[0]), .B(n57565), .X(n38858) );
  nand_x1_sg U53033 ( .A(n38849), .B(n38850), .X(n45770) );
  nand_x1_sg U53034 ( .A(i_5[19]), .B(n57563), .X(n38850) );
  nand_x1_sg U53035 ( .A(n38851), .B(n38852), .X(n45771) );
  nand_x1_sg U53036 ( .A(i_5[18]), .B(n57616), .X(n38852) );
  nand_x1_sg U53037 ( .A(n38729), .B(n38730), .X(n45710) );
  nand_x1_sg U53038 ( .A(i_5[17]), .B(n57572), .X(n38730) );
  nand_x1_sg U53039 ( .A(n38853), .B(n38854), .X(n45772) );
  nand_x1_sg U53040 ( .A(i_5[16]), .B(n57617), .X(n38854) );
  nand_x1_sg U53041 ( .A(n38845), .B(n38846), .X(n45768) );
  nand_x1_sg U53042 ( .A(i_5[15]), .B(n57577), .X(n38846) );
  nand_x1_sg U53043 ( .A(n38847), .B(n38848), .X(n45769) );
  nand_x1_sg U53044 ( .A(i_5[14]), .B(n57623), .X(n38848) );
  nand_x1_sg U53045 ( .A(n38907), .B(n38908), .X(n45799) );
  nand_x1_sg U53046 ( .A(i_5[13]), .B(n57580), .X(n38908) );
  nand_x1_sg U53047 ( .A(n38909), .B(n38910), .X(n45800) );
  nand_x1_sg U53048 ( .A(i_5[12]), .B(n57580), .X(n38910) );
  nand_x1_sg U53049 ( .A(n38901), .B(n38902), .X(n45796) );
  nand_x1_sg U53050 ( .A(i_5[11]), .B(n57580), .X(n38902) );
  nand_x1_sg U53051 ( .A(n38903), .B(n38904), .X(n45797) );
  nand_x1_sg U53052 ( .A(i_5[10]), .B(n57580), .X(n38904) );
  nand_x1_sg U53053 ( .A(n38905), .B(n38906), .X(n45798) );
  nand_x1_sg U53054 ( .A(i_5[9]), .B(n57580), .X(n38906) );
  nand_x1_sg U53055 ( .A(n38885), .B(n38886), .X(n45788) );
  nand_x1_sg U53056 ( .A(i_5[8]), .B(n57579), .X(n38886) );
  nand_x1_sg U53057 ( .A(n38897), .B(n38898), .X(n45794) );
  nand_x1_sg U53058 ( .A(i_5[7]), .B(n57579), .X(n38898) );
  nand_x1_sg U53059 ( .A(n38899), .B(n38900), .X(n45795) );
  nand_x1_sg U53060 ( .A(i_5[6]), .B(n57579), .X(n38900) );
  nand_x1_sg U53061 ( .A(n38871), .B(n38872), .X(n45781) );
  nand_x1_sg U53062 ( .A(i_5[5]), .B(n57578), .X(n38872) );
  nand_x1_sg U53063 ( .A(n38859), .B(n38860), .X(n45775) );
  nand_x1_sg U53064 ( .A(i_5[4]), .B(n57618), .X(n38860) );
  nand_x1_sg U53065 ( .A(n38883), .B(n38884), .X(n45787) );
  nand_x1_sg U53066 ( .A(i_5[3]), .B(n57579), .X(n38884) );
  nand_x1_sg U53067 ( .A(n38865), .B(n38866), .X(n45778) );
  nand_x1_sg U53068 ( .A(i_5[2]), .B(n57578), .X(n38866) );
  nand_x1_sg U53069 ( .A(n38893), .B(n38894), .X(n45792) );
  nand_x1_sg U53070 ( .A(i_5[1]), .B(n57579), .X(n38894) );
  nand_x1_sg U53071 ( .A(n38895), .B(n38896), .X(n45793) );
  nand_x1_sg U53072 ( .A(i_5[0]), .B(n57579), .X(n38896) );
  nand_x1_sg U53073 ( .A(n38887), .B(n38888), .X(n45789) );
  nand_x1_sg U53074 ( .A(i_4[19]), .B(n57579), .X(n38888) );
  nand_x1_sg U53075 ( .A(n38889), .B(n38890), .X(n45790) );
  nand_x1_sg U53076 ( .A(i_4[18]), .B(n57579), .X(n38890) );
  nand_x1_sg U53077 ( .A(n38781), .B(n38782), .X(n45736) );
  nand_x1_sg U53078 ( .A(i_4[17]), .B(n57598), .X(n38782) );
  nand_x1_sg U53079 ( .A(n38783), .B(n38784), .X(n45737) );
  nand_x1_sg U53080 ( .A(i_4[16]), .B(n57623), .X(n38784) );
  nand_x1_sg U53081 ( .A(n38775), .B(n38776), .X(n45733) );
  nand_x1_sg U53082 ( .A(i_4[15]), .B(n57598), .X(n38776) );
  nand_x1_sg U53083 ( .A(n38777), .B(n38778), .X(n45734) );
  nand_x1_sg U53084 ( .A(i_4[14]), .B(n57598), .X(n38778) );
  nand_x1_sg U53085 ( .A(n38793), .B(n38794), .X(n45742) );
  nand_x1_sg U53086 ( .A(i_4[13]), .B(n57575), .X(n38794) );
  nand_x1_sg U53087 ( .A(n38795), .B(n38796), .X(n45743) );
  nand_x1_sg U53088 ( .A(i_4[12]), .B(n57575), .X(n38796) );
  nand_x1_sg U53089 ( .A(n38787), .B(n38788), .X(n45739) );
  nand_x1_sg U53090 ( .A(i_4[11]), .B(n57598), .X(n38788) );
  nand_x1_sg U53091 ( .A(n38789), .B(n38790), .X(n45740) );
  nand_x1_sg U53092 ( .A(i_4[10]), .B(n57623), .X(n38790) );
  nand_x1_sg U53093 ( .A(n38757), .B(n38758), .X(n45724) );
  nand_x1_sg U53094 ( .A(i_4[9]), .B(n57574), .X(n38758) );
  nand_x1_sg U53095 ( .A(n38759), .B(n38760), .X(n45725) );
  nand_x1_sg U53096 ( .A(i_4[8]), .B(n57574), .X(n38760) );
  nand_x1_sg U53097 ( .A(n38751), .B(n38752), .X(n45721) );
  nand_x1_sg U53098 ( .A(i_4[7]), .B(n57573), .X(n38752) );
  nand_x1_sg U53099 ( .A(n38753), .B(n38754), .X(n45722) );
  nand_x1_sg U53100 ( .A(i_4[6]), .B(n57573), .X(n38754) );
  nand_x1_sg U53101 ( .A(n38769), .B(n38770), .X(n45730) );
  nand_x1_sg U53102 ( .A(i_4[5]), .B(n57574), .X(n38770) );
  nand_x1_sg U53103 ( .A(n38771), .B(n38772), .X(n45731) );
  nand_x1_sg U53104 ( .A(i_4[4]), .B(n57574), .X(n38772) );
  nand_x1_sg U53105 ( .A(n38763), .B(n38764), .X(n45727) );
  nand_x1_sg U53106 ( .A(i_4[3]), .B(n57574), .X(n38764) );
  nand_x1_sg U53107 ( .A(n38765), .B(n38766), .X(n45728) );
  nand_x1_sg U53108 ( .A(i_4[2]), .B(n57574), .X(n38766) );
  nand_x1_sg U53109 ( .A(n38829), .B(n38830), .X(n45760) );
  nand_x1_sg U53110 ( .A(i_4[1]), .B(n57577), .X(n38830) );
  nand_x1_sg U53111 ( .A(n38831), .B(n38832), .X(n45761) );
  nand_x1_sg U53112 ( .A(i_4[0]), .B(n57577), .X(n38832) );
  nand_x1_sg U53113 ( .A(n38823), .B(n38824), .X(n45757) );
  nand_x1_sg U53114 ( .A(i_3[19]), .B(n57576), .X(n38824) );
  nand_x1_sg U53115 ( .A(n38825), .B(n38826), .X(n45758) );
  nand_x1_sg U53116 ( .A(i_3[18]), .B(n57576), .X(n38826) );
  nand_x1_sg U53117 ( .A(n38841), .B(n38842), .X(n45766) );
  nand_x1_sg U53118 ( .A(i_3[17]), .B(n57577), .X(n38842) );
  nand_x1_sg U53119 ( .A(n38843), .B(n38844), .X(n45767) );
  nand_x1_sg U53120 ( .A(i_3[16]), .B(n57577), .X(n38844) );
  nand_x1_sg U53121 ( .A(n38835), .B(n38836), .X(n45763) );
  nand_x1_sg U53122 ( .A(i_3[15]), .B(n57577), .X(n38836) );
  nand_x1_sg U53123 ( .A(n38837), .B(n38838), .X(n45764) );
  nand_x1_sg U53124 ( .A(i_3[14]), .B(n57577), .X(n38838) );
  nand_x1_sg U53125 ( .A(n38805), .B(n38806), .X(n45748) );
  nand_x1_sg U53126 ( .A(i_3[13]), .B(n57575), .X(n38806) );
  nand_x1_sg U53127 ( .A(n38807), .B(n38808), .X(n45749) );
  nand_x1_sg U53128 ( .A(i_3[12]), .B(n57575), .X(n38808) );
  nand_x1_sg U53129 ( .A(n38799), .B(n38800), .X(n45745) );
  nand_x1_sg U53130 ( .A(i_3[11]), .B(n57575), .X(n38800) );
  nand_x1_sg U53131 ( .A(n38801), .B(n38802), .X(n45746) );
  nand_x1_sg U53132 ( .A(i_3[10]), .B(n57575), .X(n38802) );
  nand_x1_sg U53133 ( .A(n38817), .B(n38818), .X(n45754) );
  nand_x1_sg U53134 ( .A(i_3[9]), .B(n57576), .X(n38818) );
  nand_x1_sg U53135 ( .A(n38819), .B(n38820), .X(n45755) );
  nand_x1_sg U53136 ( .A(i_3[8]), .B(n57576), .X(n38820) );
  nand_x1_sg U53137 ( .A(n38811), .B(n38812), .X(n45751) );
  nand_x1_sg U53138 ( .A(i_3[7]), .B(n57576), .X(n38812) );
  nand_x1_sg U53139 ( .A(n38813), .B(n38814), .X(n45752) );
  nand_x1_sg U53140 ( .A(i_3[6]), .B(n57576), .X(n38814) );
  nand_x1_sg U53141 ( .A(n39037), .B(n39038), .X(n45864) );
  nand_x1_sg U53142 ( .A(i_3[5]), .B(n57587), .X(n39038) );
  nand_x1_sg U53143 ( .A(n39039), .B(n39040), .X(n45865) );
  nand_x1_sg U53144 ( .A(i_3[4]), .B(n57587), .X(n39040) );
  nand_x1_sg U53145 ( .A(n39031), .B(n39032), .X(n45861) );
  nand_x1_sg U53146 ( .A(i_3[3]), .B(n57587), .X(n39032) );
  nand_x1_sg U53147 ( .A(n39033), .B(n39034), .X(n45862) );
  nand_x1_sg U53148 ( .A(i_3[2]), .B(n57587), .X(n39034) );
  nand_x1_sg U53149 ( .A(n39015), .B(n39016), .X(n45853) );
  nand_x1_sg U53150 ( .A(i_3[1]), .B(n57586), .X(n39016) );
  nand_x1_sg U53151 ( .A(n39029), .B(n39030), .X(n45860) );
  nand_x1_sg U53152 ( .A(i_3[0]), .B(n57587), .X(n39030) );
  nand_x1_sg U53153 ( .A(n39017), .B(n39018), .X(n45854) );
  nand_x1_sg U53154 ( .A(i_2[19]), .B(n57586), .X(n39018) );
  nand_x1_sg U53155 ( .A(n39019), .B(n39020), .X(n45855) );
  nand_x1_sg U53156 ( .A(i_2[18]), .B(n57586), .X(n39020) );
  nand_x1_sg U53157 ( .A(n39011), .B(n39012), .X(n45851) );
  nand_x1_sg U53158 ( .A(i_2[17]), .B(n57586), .X(n39012) );
  nand_x1_sg U53159 ( .A(n39013), .B(n39014), .X(n45852) );
  nand_x1_sg U53160 ( .A(i_2[16]), .B(n57586), .X(n39014) );
  nand_x1_sg U53161 ( .A(n39007), .B(n39008), .X(n45849) );
  nand_x1_sg U53162 ( .A(i_2[15]), .B(n57585), .X(n39008) );
  nand_x1_sg U53163 ( .A(n39009), .B(n39010), .X(n45850) );
  nand_x1_sg U53164 ( .A(i_2[14]), .B(n57586), .X(n39010) );
  nand_x1_sg U53165 ( .A(n39023), .B(n39024), .X(n45857) );
  nand_x1_sg U53166 ( .A(i_2[13]), .B(n57586), .X(n39024) );
  nand_x1_sg U53167 ( .A(n39025), .B(n39026), .X(n45858) );
  nand_x1_sg U53168 ( .A(i_2[12]), .B(n57586), .X(n39026) );
  nand_x1_sg U53169 ( .A(n39005), .B(n39006), .X(n45848) );
  nand_x1_sg U53170 ( .A(i_2[11]), .B(n57585), .X(n39006) );
  nand_x1_sg U53171 ( .A(n39021), .B(n39022), .X(n45856) );
  nand_x1_sg U53172 ( .A(i_2[10]), .B(n57586), .X(n39022) );
  nand_x1_sg U53173 ( .A(n39069), .B(n39070), .X(n45880) );
  nand_x1_sg U53174 ( .A(i_2[9]), .B(n57589), .X(n39070) );
  nand_x1_sg U53175 ( .A(n39027), .B(n39028), .X(n45859) );
  nand_x1_sg U53176 ( .A(i_2[8]), .B(n57587), .X(n39028) );
  nand_x1_sg U53177 ( .A(n39041), .B(n39042), .X(n45866) );
  nand_x1_sg U53178 ( .A(i_2[7]), .B(n57587), .X(n39042) );
  nand_x1_sg U53179 ( .A(n39047), .B(n39048), .X(n45869) );
  nand_x1_sg U53180 ( .A(i_2[6]), .B(n57588), .X(n39048) );
  nand_x1_sg U53181 ( .A(n38723), .B(n38724), .X(n45707) );
  nand_x1_sg U53182 ( .A(i_2[5]), .B(n57572), .X(n38724) );
  nand_x1_sg U53183 ( .A(n38725), .B(n38726), .X(n45708) );
  nand_x1_sg U53184 ( .A(i_2[4]), .B(n57572), .X(n38726) );
  nand_x1_sg U53185 ( .A(n39065), .B(n39066), .X(n45878) );
  nand_x1_sg U53186 ( .A(i_2[3]), .B(n57589), .X(n39066) );
  nand_x1_sg U53187 ( .A(n39067), .B(n39068), .X(n45879) );
  nand_x1_sg U53188 ( .A(i_2[2]), .B(n57589), .X(n39068) );
  nand_x1_sg U53189 ( .A(n39049), .B(n39050), .X(n45870) );
  nand_x1_sg U53190 ( .A(i_2[1]), .B(n57588), .X(n39050) );
  nand_x1_sg U53191 ( .A(n39051), .B(n39052), .X(n45871) );
  nand_x1_sg U53192 ( .A(i_2[0]), .B(n57588), .X(n39052) );
  nand_x1_sg U53193 ( .A(n39043), .B(n39044), .X(n45867) );
  nand_x1_sg U53194 ( .A(i_1[19]), .B(n57587), .X(n39044) );
  nand_x1_sg U53195 ( .A(n39045), .B(n39046), .X(n45868) );
  nand_x1_sg U53196 ( .A(i_1[18]), .B(n57588), .X(n39046) );
  nand_x1_sg U53197 ( .A(n39061), .B(n39062), .X(n45876) );
  nand_x1_sg U53198 ( .A(i_1[17]), .B(n57588), .X(n39062) );
  nand_x1_sg U53199 ( .A(n39063), .B(n39064), .X(n45877) );
  nand_x1_sg U53200 ( .A(i_1[16]), .B(n57589), .X(n39064) );
  nand_x1_sg U53201 ( .A(n39055), .B(n39056), .X(n45873) );
  nand_x1_sg U53202 ( .A(i_1[15]), .B(n57588), .X(n39056) );
  nand_x1_sg U53203 ( .A(n39057), .B(n39058), .X(n45874) );
  nand_x1_sg U53204 ( .A(i_1[14]), .B(n57588), .X(n39058) );
  nand_x1_sg U53205 ( .A(n38963), .B(n38964), .X(n45827) );
  nand_x1_sg U53206 ( .A(i_1[13]), .B(n57583), .X(n38964) );
  nand_x1_sg U53207 ( .A(n38965), .B(n38966), .X(n45828) );
  nand_x1_sg U53208 ( .A(i_1[12]), .B(n57583), .X(n38966) );
  nand_x1_sg U53209 ( .A(n38957), .B(n38958), .X(n45824) );
  nand_x1_sg U53210 ( .A(i_1[11]), .B(n57583), .X(n38958) );
  nand_x1_sg U53211 ( .A(n38959), .B(n38960), .X(n45825) );
  nand_x1_sg U53212 ( .A(i_1[10]), .B(n57583), .X(n38960) );
  nand_x1_sg U53213 ( .A(n38967), .B(n38968), .X(n45829) );
  nand_x1_sg U53214 ( .A(i_1[9]), .B(n57583), .X(n38968) );
  nand_x1_sg U53215 ( .A(n38955), .B(n38956), .X(n45823) );
  nand_x1_sg U53216 ( .A(i_1[8]), .B(n57583), .X(n38956) );
  nand_x1_sg U53217 ( .A(n38961), .B(n38962), .X(n45826) );
  nand_x1_sg U53218 ( .A(i_1[7]), .B(n57583), .X(n38962) );
  nand_x1_sg U53219 ( .A(n38953), .B(n38954), .X(n45822) );
  nand_x1_sg U53220 ( .A(i_1[6]), .B(n57582), .X(n38954) );
  nand_x1_sg U53221 ( .A(n38919), .B(n38920), .X(n45805) );
  nand_x1_sg U53222 ( .A(i_1[5]), .B(n57581), .X(n38920) );
  nand_x1_sg U53223 ( .A(n38921), .B(n38922), .X(n45806) );
  nand_x1_sg U53224 ( .A(i_1[4]), .B(n57581), .X(n38922) );
  nand_x1_sg U53225 ( .A(n38913), .B(n38914), .X(n45802) );
  nand_x1_sg U53226 ( .A(i_1[3]), .B(n57580), .X(n38914) );
  nand_x1_sg U53227 ( .A(n38915), .B(n38916), .X(n45803) );
  nand_x1_sg U53228 ( .A(i_1[2]), .B(n57580), .X(n38916) );
  nand_x1_sg U53229 ( .A(n38947), .B(n38948), .X(n45819) );
  nand_x1_sg U53230 ( .A(i_1[1]), .B(n57582), .X(n38948) );
  nand_x1_sg U53231 ( .A(n38911), .B(n38912), .X(n45801) );
  nand_x1_sg U53232 ( .A(i_1[0]), .B(n57580), .X(n38912) );
  nand_x1_sg U53233 ( .A(n38949), .B(n38950), .X(n45820) );
  nand_x1_sg U53234 ( .A(i_0[19]), .B(n57582), .X(n38950) );
  nand_x1_sg U53235 ( .A(n38951), .B(n38952), .X(n45821) );
  nand_x1_sg U53236 ( .A(i_0[18]), .B(n57582), .X(n38952) );
  nand_x1_sg U53237 ( .A(n38973), .B(n38974), .X(n45832) );
  nand_x1_sg U53238 ( .A(i_0[17]), .B(n57584), .X(n38974) );
  nand_x1_sg U53239 ( .A(n38991), .B(n38992), .X(n45841) );
  nand_x1_sg U53240 ( .A(i_0[16]), .B(n57585), .X(n38992) );
  nand_x1_sg U53241 ( .A(n38993), .B(n38994), .X(n45842) );
  nand_x1_sg U53242 ( .A(i_0[15]), .B(n57585), .X(n38994) );
  nand_x1_sg U53243 ( .A(n38999), .B(n39000), .X(n45845) );
  nand_x1_sg U53244 ( .A(i_0[14]), .B(n57585), .X(n39000) );
  nand_x1_sg U53245 ( .A(n39001), .B(n39002), .X(n45846) );
  nand_x1_sg U53246 ( .A(i_0[13]), .B(n57585), .X(n39002) );
  nand_x1_sg U53247 ( .A(n39003), .B(n39004), .X(n45847) );
  nand_x1_sg U53248 ( .A(i_0[12]), .B(n57585), .X(n39004) );
  nand_x1_sg U53249 ( .A(n38995), .B(n38996), .X(n45843) );
  nand_x1_sg U53250 ( .A(i_0[11]), .B(n57585), .X(n38996) );
  nand_x1_sg U53251 ( .A(n38997), .B(n38998), .X(n45844) );
  nand_x1_sg U53252 ( .A(i_0[10]), .B(n57585), .X(n38998) );
  nand_x1_sg U53253 ( .A(n38975), .B(n38976), .X(n45833) );
  nand_x1_sg U53254 ( .A(i_0[9]), .B(n57584), .X(n38976) );
  nand_x1_sg U53255 ( .A(n38977), .B(n38978), .X(n45834) );
  nand_x1_sg U53256 ( .A(i_0[8]), .B(n57584), .X(n38978) );
  nand_x1_sg U53257 ( .A(n38969), .B(n38970), .X(n45830) );
  nand_x1_sg U53258 ( .A(i_0[7]), .B(n57583), .X(n38970) );
  nand_x1_sg U53259 ( .A(n38971), .B(n38972), .X(n45831) );
  nand_x1_sg U53260 ( .A(i_0[6]), .B(n57583), .X(n38972) );
  nand_x1_sg U53261 ( .A(n38987), .B(n38988), .X(n45839) );
  nand_x1_sg U53262 ( .A(i_0[5]), .B(n57584), .X(n38988) );
  nand_x1_sg U53263 ( .A(n38989), .B(n38990), .X(n45840) );
  nand_x1_sg U53264 ( .A(i_0[4]), .B(n57584), .X(n38990) );
  nand_x1_sg U53265 ( .A(n38981), .B(n38982), .X(n45836) );
  nand_x1_sg U53266 ( .A(i_0[3]), .B(n57584), .X(n38982) );
  nand_x1_sg U53267 ( .A(n38983), .B(n38984), .X(n45837) );
  nand_x1_sg U53268 ( .A(i_0[2]), .B(n57584), .X(n38984) );
  nand_x1_sg U53269 ( .A(n38731), .B(n38732), .X(n45711) );
  nand_x1_sg U53270 ( .A(i_0[1]), .B(n57572), .X(n38732) );
  nand_x1_sg U53271 ( .A(n38733), .B(n38734), .X(n45712) );
  nand_x1_sg U53272 ( .A(i_0[0]), .B(n57572), .X(n38734) );
  nand_x1_sg U53273 ( .A(n39706), .B(n39707), .X(n10462) );
  nand_x1_sg U53274 ( .A(i_mask[0]), .B(n57619), .X(n39707) );
  nand_x1_sg U53275 ( .A(n39708), .B(n39709), .X(n10461) );
  nand_x1_sg U53276 ( .A(i_mask[1]), .B(n57628), .X(n39709) );
  nand_x1_sg U53277 ( .A(n39710), .B(n39711), .X(n10460) );
  nand_x1_sg U53278 ( .A(i_mask[2]), .B(n57629), .X(n39711) );
  nand_x1_sg U53279 ( .A(n39712), .B(n39713), .X(n10459) );
  nand_x1_sg U53280 ( .A(i_mask[3]), .B(n57630), .X(n39713) );
  nand_x1_sg U53281 ( .A(n39714), .B(n39715), .X(n10458) );
  nand_x1_sg U53282 ( .A(i_mask[4]), .B(n57632), .X(n39715) );
  nand_x1_sg U53283 ( .A(n39716), .B(n39717), .X(n10457) );
  nand_x1_sg U53284 ( .A(i_mask[5]), .B(n57615), .X(n39717) );
  nand_x1_sg U53285 ( .A(n39718), .B(n39719), .X(n10456) );
  nand_x1_sg U53286 ( .A(i_mask[6]), .B(n57618), .X(n39719) );
  nand_x1_sg U53287 ( .A(n39720), .B(n39721), .X(n10455) );
  nand_x1_sg U53288 ( .A(i_mask[7]), .B(n57629), .X(n39721) );
  nand_x1_sg U53289 ( .A(n39722), .B(n39723), .X(n10454) );
  nand_x1_sg U53290 ( .A(i_mask[8]), .B(n57625), .X(n39723) );
  nand_x1_sg U53291 ( .A(n39724), .B(n39725), .X(n10453) );
  nand_x1_sg U53292 ( .A(i_mask[9]), .B(n57632), .X(n39725) );
  nand_x1_sg U53293 ( .A(n39726), .B(n39727), .X(n10452) );
  nand_x1_sg U53294 ( .A(i_mask[10]), .B(n57615), .X(n39727) );
  nand_x1_sg U53295 ( .A(n39728), .B(n39729), .X(n10451) );
  nand_x1_sg U53296 ( .A(i_mask[11]), .B(n57629), .X(n39729) );
  nand_x1_sg U53297 ( .A(n39730), .B(n39731), .X(n10450) );
  nand_x1_sg U53298 ( .A(i_mask[12]), .B(n57629), .X(n39731) );
  nand_x1_sg U53299 ( .A(n39732), .B(n39733), .X(n10449) );
  nand_x1_sg U53300 ( .A(i_mask[13]), .B(n57630), .X(n39733) );
  nand_x1_sg U53301 ( .A(n39734), .B(n39735), .X(n10448) );
  nand_x1_sg U53302 ( .A(i_mask[14]), .B(n57625), .X(n39735) );
  nand_x1_sg U53303 ( .A(n39736), .B(n39737), .X(n10447) );
  nand_x1_sg U53304 ( .A(i_mask[15]), .B(n57625), .X(n39737) );
  nand_x1_sg U53305 ( .A(n39738), .B(n39739), .X(n10446) );
  nand_x1_sg U53306 ( .A(i_mask[16]), .B(n57600), .X(n39739) );
  nand_x1_sg U53307 ( .A(n39740), .B(n39741), .X(n10445) );
  nand_x1_sg U53308 ( .A(i_mask[17]), .B(n57624), .X(n39741) );
  nand_x1_sg U53309 ( .A(n39742), .B(n39743), .X(n10444) );
  nand_x1_sg U53310 ( .A(i_mask[18]), .B(n57623), .X(n39743) );
  nand_x1_sg U53311 ( .A(n39744), .B(n39745), .X(n10443) );
  nand_x1_sg U53312 ( .A(i_mask[19]), .B(n57625), .X(n39745) );
  nand_x1_sg U53313 ( .A(n39746), .B(n39747), .X(n10442) );
  nand_x1_sg U53314 ( .A(i_mask[20]), .B(n57623), .X(n39747) );
  nand_x1_sg U53315 ( .A(n39748), .B(n39749), .X(n10441) );
  nand_x1_sg U53316 ( .A(i_mask[21]), .B(n57618), .X(n39749) );
  nand_x1_sg U53317 ( .A(n39750), .B(n39751), .X(n10440) );
  nand_x1_sg U53318 ( .A(i_mask[22]), .B(n57619), .X(n39751) );
  nand_x1_sg U53319 ( .A(n39752), .B(n39753), .X(n10439) );
  nand_x1_sg U53320 ( .A(i_mask[23]), .B(n57616), .X(n39753) );
  nand_x1_sg U53321 ( .A(n39754), .B(n39755), .X(n10438) );
  nand_x1_sg U53322 ( .A(i_mask[24]), .B(n57617), .X(n39755) );
  nand_x1_sg U53323 ( .A(n39756), .B(n39757), .X(n10437) );
  nand_x1_sg U53324 ( .A(i_mask[25]), .B(n57628), .X(n39757) );
  nand_x1_sg U53325 ( .A(n39758), .B(n39759), .X(n10436) );
  nand_x1_sg U53326 ( .A(i_mask[26]), .B(n57628), .X(n39759) );
  nand_x1_sg U53327 ( .A(n39760), .B(n39761), .X(n10435) );
  nand_x1_sg U53328 ( .A(i_mask[27]), .B(n57618), .X(n39761) );
  nand_x1_sg U53329 ( .A(n39762), .B(n39763), .X(n10434) );
  nand_x1_sg U53330 ( .A(i_mask[28]), .B(n57628), .X(n39763) );
  nand_x1_sg U53331 ( .A(n39764), .B(n39765), .X(n10433) );
  nand_x1_sg U53332 ( .A(i_mask[29]), .B(n57628), .X(n39765) );
  nand_x1_sg U53333 ( .A(n39766), .B(n39767), .X(n10432) );
  nand_x1_sg U53334 ( .A(i_mask[30]), .B(n57619), .X(n39767) );
  nand_x1_sg U53335 ( .A(n39768), .B(n39769), .X(n10431) );
  nand_x1_sg U53336 ( .A(i_mask[31]), .B(n57616), .X(n39769) );
  nand_x1_sg U53337 ( .A(n39770), .B(n39771), .X(n10430) );
  nand_x1_sg U53338 ( .A(w_mask[0]), .B(n57617), .X(n39771) );
  nand_x1_sg U53339 ( .A(n39772), .B(n39773), .X(n10429) );
  nand_x1_sg U53340 ( .A(w_mask[1]), .B(n57628), .X(n39773) );
  nand_x1_sg U53341 ( .A(n39774), .B(n39775), .X(n10428) );
  nand_x1_sg U53342 ( .A(w_mask[2]), .B(n57625), .X(n39775) );
  nand_x1_sg U53343 ( .A(n39776), .B(n39777), .X(n10427) );
  nand_x1_sg U53344 ( .A(w_mask[3]), .B(n57629), .X(n39777) );
  nand_x1_sg U53345 ( .A(n39778), .B(n39779), .X(n10426) );
  nand_x1_sg U53346 ( .A(w_mask[4]), .B(n57630), .X(n39779) );
  nand_x1_sg U53347 ( .A(n39780), .B(n39781), .X(n10425) );
  nand_x1_sg U53348 ( .A(w_mask[5]), .B(n57621), .X(n39781) );
  nand_x1_sg U53349 ( .A(n39782), .B(n39783), .X(n10424) );
  nand_x1_sg U53350 ( .A(w_mask[6]), .B(n57625), .X(n39783) );
  nand_x1_sg U53351 ( .A(n39784), .B(n39785), .X(n10423) );
  nand_x1_sg U53352 ( .A(w_mask[7]), .B(n57629), .X(n39785) );
  nand_x1_sg U53353 ( .A(n39786), .B(n39787), .X(n10422) );
  nand_x1_sg U53354 ( .A(w_mask[8]), .B(n57630), .X(n39787) );
  nand_x1_sg U53355 ( .A(n39788), .B(n39789), .X(n10421) );
  nand_x1_sg U53356 ( .A(w_mask[9]), .B(n57620), .X(n39789) );
  nand_x1_sg U53357 ( .A(n39790), .B(n39791), .X(n10420) );
  nand_x1_sg U53358 ( .A(w_mask[10]), .B(n57625), .X(n39791) );
  nand_x1_sg U53359 ( .A(n39792), .B(n39793), .X(n10419) );
  nand_x1_sg U53360 ( .A(w_mask[11]), .B(n57615), .X(n39793) );
  nand_x1_sg U53361 ( .A(n39794), .B(n39795), .X(n10418) );
  nand_x1_sg U53362 ( .A(w_mask[12]), .B(n57600), .X(n39795) );
  nand_x1_sg U53363 ( .A(n39796), .B(n39797), .X(n10417) );
  nand_x1_sg U53364 ( .A(w_mask[13]), .B(n57620), .X(n39797) );
  nand_x1_sg U53365 ( .A(n39798), .B(n39799), .X(n10416) );
  nand_x1_sg U53366 ( .A(w_mask[14]), .B(n57615), .X(n39799) );
  nand_x1_sg U53367 ( .A(n39800), .B(n39801), .X(n10415) );
  nand_x1_sg U53368 ( .A(w_mask[15]), .B(n57630), .X(n39801) );
  nand_x1_sg U53369 ( .A(n39802), .B(n39803), .X(n10414) );
  nand_x1_sg U53370 ( .A(w_mask[16]), .B(n57621), .X(n39803) );
  nand_x1_sg U53371 ( .A(n39804), .B(n39805), .X(n10413) );
  nand_x1_sg U53372 ( .A(w_mask[17]), .B(n57615), .X(n39805) );
  nand_x1_sg U53373 ( .A(n39806), .B(n39807), .X(n10412) );
  nand_x1_sg U53374 ( .A(w_mask[18]), .B(n57616), .X(n39807) );
  nand_x1_sg U53375 ( .A(n39808), .B(n39809), .X(n10411) );
  nand_x1_sg U53376 ( .A(w_mask[19]), .B(n57624), .X(n39809) );
  nand_x1_sg U53377 ( .A(n39810), .B(n39811), .X(n10410) );
  nand_x1_sg U53378 ( .A(w_mask[20]), .B(n57630), .X(n39811) );
  nand_x1_sg U53379 ( .A(n39812), .B(n39813), .X(n10409) );
  nand_x1_sg U53380 ( .A(w_mask[21]), .B(n57615), .X(n39813) );
  nand_x1_sg U53381 ( .A(n39814), .B(n39815), .X(n10408) );
  nand_x1_sg U53382 ( .A(w_mask[22]), .B(n57624), .X(n39815) );
  nand_x1_sg U53383 ( .A(n39816), .B(n39817), .X(n10407) );
  nand_x1_sg U53384 ( .A(w_mask[23]), .B(n57630), .X(n39817) );
  nand_x1_sg U53385 ( .A(n39818), .B(n39819), .X(n10406) );
  nand_x1_sg U53386 ( .A(w_mask[24]), .B(n57625), .X(n39819) );
  nand_x1_sg U53387 ( .A(n39820), .B(n39821), .X(n10405) );
  nand_x1_sg U53388 ( .A(w_mask[25]), .B(n57624), .X(n39821) );
  nand_x1_sg U53389 ( .A(n39822), .B(n39823), .X(n10404) );
  nand_x1_sg U53390 ( .A(w_mask[26]), .B(n57624), .X(n39823) );
  nand_x1_sg U53391 ( .A(n39824), .B(n39825), .X(n10403) );
  nand_x1_sg U53392 ( .A(w_mask[27]), .B(n57615), .X(n39825) );
  nand_x1_sg U53393 ( .A(n39826), .B(n39827), .X(n10402) );
  nand_x1_sg U53394 ( .A(w_mask[28]), .B(n57567), .X(n39827) );
  nand_x1_sg U53395 ( .A(n39828), .B(n39829), .X(n10401) );
  nand_x1_sg U53396 ( .A(w_mask[29]), .B(n57615), .X(n39829) );
  nand_x1_sg U53397 ( .A(n39830), .B(n39831), .X(n10400) );
  nand_x1_sg U53398 ( .A(w_mask[30]), .B(n57619), .X(n39831) );
  nand_x1_sg U53399 ( .A(n39832), .B(n39833), .X(n10399) );
  nand_x1_sg U53400 ( .A(w_mask[31]), .B(n57615), .X(n39833) );
  nand_x1_sg U53401 ( .A(n38408), .B(n38409), .X(n45552) );
  inv_x1_sg U53402 ( .A(n35549), .X(n68246) );
  inv_x1_sg U53403 ( .A(n35522), .X(n68255) );
  inv_x1_sg U53404 ( .A(n35609), .X(n68239) );
  nand_x4_sg U53405 ( .A(n25964), .B(n25965), .X(n24146) );
  nand_x4_sg U53406 ( .A(n25784), .B(n25785), .X(n24116) );
  nand_x4_sg U53407 ( .A(n25544), .B(n25545), .X(n24076) );
  nand_x4_sg U53408 ( .A(n25212), .B(n25213), .X(n24011) );
  nand_x4_sg U53409 ( .A(n25062), .B(n25063), .X(n23986) );
  nand_x2_sg U53410 ( .A(n47377), .B(n57862), .X(n23168) );
  nand_x2_sg U53411 ( .A(n47381), .B(n57862), .X(n23069) );
  nand_x2_sg U53412 ( .A(n47383), .B(n57862), .X(n22992) );
  nand_x2_sg U53413 ( .A(n47385), .B(n57862), .X(n22886) );
  nand_x2_sg U53414 ( .A(n47387), .B(n57862), .X(n22798) );
  inv_x2_sg U53415 ( .A(n47446), .X(n47447) );
  inv_x2_sg U53416 ( .A(n47448), .X(n47449) );
  inv_x2_sg U53417 ( .A(n47450), .X(n47451) );
  inv_x2_sg U53418 ( .A(n47452), .X(n47453) );
  nor_x2_sg U53419 ( .A(n57023), .B(n22988), .X(n23164) );
  nor_x2_sg U53420 ( .A(n51501), .B(n57152), .X(n23153) );
  nor_x2_sg U53421 ( .A(n57027), .B(n22761), .X(n22937) );
  nor_x2_sg U53422 ( .A(n51505), .B(n57158), .X(n22926) );
  inv_x4_sg U53423 ( .A(n25870), .X(n67459) );
  inv_x4_sg U53424 ( .A(n25720), .X(n67464) );
  inv_x4_sg U53425 ( .A(n25480), .X(n67472) );
  inv_x4_sg U53426 ( .A(n25148), .X(n67270) );
  inv_x4_sg U53427 ( .A(n25028), .X(n67274) );
  nor_x4_sg U53428 ( .A(n24487), .B(n67096), .X(n24479) );
  nor_x2_sg U53429 ( .A(n47775), .B(n67096), .X(n24485) );
  inv_x1_sg U53430 ( .A(n35553), .X(n68235) );
  inv_x1_sg U53431 ( .A(n35543), .X(n68262) );
  inv_x1_sg U53432 ( .A(n35557), .X(n68245) );
  inv_x1_sg U53433 ( .A(n35515), .X(n68256) );
  inv_x1_sg U53434 ( .A(n35513), .X(n68238) );
  nand_x4_sg U53435 ( .A(n25694), .B(n25695), .X(n24101) );
  nand_x4_sg U53436 ( .A(n25514), .B(n25515), .X(n24071) );
  nand_x4_sg U53437 ( .A(n25182), .B(n25183), .X(n24006) );
  nand_x4_sg U53438 ( .A(n24942), .B(n24943), .X(n23966) );
  nand_x2_sg U53439 ( .A(n47379), .B(n57862), .X(n23157) );
  nand_x2_sg U53440 ( .A(n47451), .B(n57862), .X(n23036) );
  nand_x2_sg U53441 ( .A(n47449), .B(n57862), .X(n22979) );
  nand_x2_sg U53442 ( .A(n47453), .B(n57862), .X(n22875) );
  nand_x2_sg U53443 ( .A(n47389), .B(n57862), .X(n22765) );
  nand_x2_sg U53444 ( .A(n68430), .B(n68431), .X(n32613) );
  nor_x2_sg U53445 ( .A(n68430), .B(n58638), .X(n58172) );
  inv_x4_sg U53446 ( .A(n55007), .X(n68430) );
  nand_x2_sg U53447 ( .A(n68428), .B(n68429), .X(n32608) );
  nor_x2_sg U53448 ( .A(n68428), .B(n57104), .X(n58192) );
  inv_x4_sg U53449 ( .A(n55003), .X(n68428) );
  nand_x2_sg U53450 ( .A(n68426), .B(n68427), .X(n32605) );
  nor_x2_sg U53451 ( .A(n68426), .B(n57103), .X(n58217) );
  inv_x4_sg U53452 ( .A(n54999), .X(n68426) );
  nand_x2_sg U53453 ( .A(n68520), .B(n68521), .X(n32168) );
  nor_x2_sg U53454 ( .A(n68520), .B(n57104), .X(n58272) );
  inv_x4_sg U53455 ( .A(n55019), .X(n68520) );
  nand_x2_sg U53456 ( .A(n68518), .B(n68519), .X(n32163) );
  nor_x2_sg U53457 ( .A(n68518), .B(n57103), .X(n58292) );
  inv_x4_sg U53458 ( .A(n55015), .X(n68518) );
  nand_x2_sg U53459 ( .A(n68516), .B(n68517), .X(n32160) );
  nor_x2_sg U53460 ( .A(n68516), .B(n58638), .X(n58317) );
  inv_x4_sg U53461 ( .A(n55011), .X(n68516) );
  inv_x2_sg U53462 ( .A(n47454), .X(n47455) );
  inv_x2_sg U53463 ( .A(n47456), .X(n47457) );
  inv_x2_sg U53464 ( .A(n47458), .X(n47459) );
  inv_x2_sg U53465 ( .A(n47460), .X(n47461) );
  inv_x2_sg U53466 ( .A(n47462), .X(n47463) );
  inv_x2_sg U53467 ( .A(n47464), .X(n47465) );
  inv_x2_sg U53468 ( .A(n47466), .X(n47467) );
  nor_x2_sg U53469 ( .A(n47755), .B(n57153), .X(n23142) );
  nor_x2_sg U53470 ( .A(n57035), .B(n22988), .X(n23131) );
  nor_x2_sg U53471 ( .A(n47757), .B(n57159), .X(n22915) );
  nor_x2_sg U53472 ( .A(n57041), .B(n22761), .X(n22904) );
  inv_x4_sg U53473 ( .A(n25630), .X(n67467) );
  inv_x4_sg U53474 ( .A(n25450), .X(n67473) );
  inv_x4_sg U53475 ( .A(n25118), .X(n67271) );
  inv_x4_sg U53476 ( .A(n24998), .X(n67275) );
  inv_x4_sg U53477 ( .A(n25960), .X(n67456) );
  inv_x1_sg U53478 ( .A(n35542), .X(n68249) );
  inv_x1_sg U53479 ( .A(n35545), .X(n68263) );
  inv_x1_sg U53480 ( .A(n35524), .X(n68253) );
  inv_x1_sg U53481 ( .A(n35517), .X(n68257) );
  inv_x1_sg U53482 ( .A(n35601), .X(n68236) );
  inv_x1_sg U53483 ( .A(n35597), .X(n68244) );
  inv_x1_sg U53484 ( .A(n35521), .X(n68237) );
  nand_x4_sg U53485 ( .A(n25934), .B(n25935), .X(n24141) );
  nand_x4_sg U53486 ( .A(n25664), .B(n25665), .X(n24096) );
  nand_x4_sg U53487 ( .A(n25332), .B(n25333), .X(n24031) );
  nand_x4_sg U53488 ( .A(n25092), .B(n25093), .X(n23991) );
  nand_x4_sg U53489 ( .A(n24912), .B(n24913), .X(n23961) );
  nand_x2_sg U53490 ( .A(n47461), .B(n57862), .X(n23146) );
  nand_x2_sg U53491 ( .A(n47459), .B(n57862), .X(n23058) );
  nand_x2_sg U53492 ( .A(n47457), .B(n57862), .X(n23003) );
  nand_x2_sg U53493 ( .A(n47467), .B(n57862), .X(n22853) );
  nand_x2_sg U53494 ( .A(n47447), .B(n57862), .X(n22776) );
  nand_x2_sg U53495 ( .A(n56969), .B(n57166), .X(n34176) );
  nor_x2_sg U53496 ( .A(n68431), .B(n57104), .X(n58167) );
  inv_x4_sg U53497 ( .A(n55009), .X(n68431) );
  nor_x2_sg U53498 ( .A(n68429), .B(n57103), .X(n58187) );
  inv_x4_sg U53499 ( .A(n55005), .X(n68429) );
  nor_x2_sg U53500 ( .A(n68427), .B(n58638), .X(n58212) );
  inv_x4_sg U53501 ( .A(n55001), .X(n68427) );
  nor_x2_sg U53502 ( .A(n68521), .B(n57103), .X(n58267) );
  inv_x4_sg U53503 ( .A(n55021), .X(n68521) );
  nor_x2_sg U53504 ( .A(n68519), .B(n58638), .X(n58287) );
  inv_x4_sg U53505 ( .A(n55017), .X(n68519) );
  nor_x2_sg U53506 ( .A(n68517), .B(n57104), .X(n58312) );
  inv_x4_sg U53507 ( .A(n55013), .X(n68517) );
  inv_x2_sg U53508 ( .A(n47468), .X(n47469) );
  inv_x2_sg U53509 ( .A(n47470), .X(n47471) );
  inv_x2_sg U53510 ( .A(n47472), .X(n47473) );
  inv_x2_sg U53511 ( .A(n47474), .X(n47475) );
  inv_x2_sg U53512 ( .A(\shifter_0/reg_w_9 [0]), .X(n47520) );
  inv_x2_sg U53513 ( .A(\shifter_0/reg_w_9 [1]), .X(n47522) );
  inv_x2_sg U53514 ( .A(\shifter_0/reg_w_9 [5]), .X(n47524) );
  inv_x2_sg U53515 ( .A(\shifter_0/reg_w_14 [0]), .X(n47532) );
  inv_x2_sg U53516 ( .A(\shifter_0/reg_w_14 [5]), .X(n47534) );
  inv_x2_sg U53517 ( .A(\shifter_0/reg_i_9 [0]), .X(n47536) );
  inv_x2_sg U53518 ( .A(\shifter_0/reg_i_9 [1]), .X(n47538) );
  inv_x2_sg U53519 ( .A(\shifter_0/reg_i_9 [5]), .X(n47540) );
  inv_x2_sg U53520 ( .A(\shifter_0/reg_i_10 [1]), .X(n47544) );
  inv_x2_sg U53521 ( .A(\shifter_0/reg_i_14 [0]), .X(n47548) );
  inv_x2_sg U53522 ( .A(\shifter_0/reg_i_14 [5]), .X(n47550) );
  inv_x2_sg U53523 ( .A(\shifter_0/reg_i_9 [17]), .X(n47552) );
  inv_x2_sg U53524 ( .A(\shifter_0/reg_w_11 [17]), .X(n47704) );
  inv_x2_sg U53525 ( .A(\shifter_0/pointer [3]), .X(n47504) );
  inv_x2_sg U53526 ( .A(\shifter_0/reg_w_2 [2]), .X(n55232) );
  inv_x2_sg U53527 ( .A(\shifter_0/reg_i_2 [17]), .X(n55248) );
  inv_x2_sg U53528 ( .A(\shifter_0/reg_i_6 [16]), .X(n47568) );
  inv_x2_sg U53529 ( .A(\shifter_0/reg_w_6 [16]), .X(n47570) );
  nor_x2_sg U53530 ( .A(n51511), .B(n57152), .X(n23120) );
  nor_x2_sg U53531 ( .A(n57019), .B(n57153), .X(n23109) );
  nor_x2_sg U53532 ( .A(n51517), .B(n57158), .X(n22893) );
  nor_x2_sg U53533 ( .A(n57021), .B(n57159), .X(n22882) );
  inv_x4_sg U53534 ( .A(n25840), .X(n67460) );
  inv_x4_sg U53535 ( .A(n25600), .X(n67468) );
  inv_x4_sg U53536 ( .A(n25389), .X(n67262) );
  inv_x4_sg U53537 ( .A(n24968), .X(n67276) );
  inv_x4_sg U53538 ( .A(n25208), .X(n67268) );
  inv_x1_sg U53539 ( .A(n35558), .X(n68261) );
  inv_x1_sg U53540 ( .A(n35536), .X(n68259) );
  inv_x1_sg U53541 ( .A(n35529), .X(n68254) );
  inv_x1_sg U53542 ( .A(n35531), .X(n68250) );
  inv_x1_sg U53543 ( .A(n35588), .X(n68234) );
  inv_x1_sg U53544 ( .A(n35613), .X(n68248) );
  inv_x1_sg U53545 ( .A(n35528), .X(n68241) );
  nand_x4_sg U53546 ( .A(n25814), .B(n25815), .X(n24121) );
  nand_x4_sg U53547 ( .A(n25362), .B(n25363), .X(n24036) );
  nand_x2_sg U53548 ( .A(n47471), .B(n57862), .X(n23124) );
  nand_x2_sg U53549 ( .A(n47469), .B(n57862), .X(n23025) );
  nand_x2_sg U53550 ( .A(n47465), .B(n57862), .X(n22963) );
  nand_x2_sg U53551 ( .A(n47463), .B(n57862), .X(n22864) );
  nand_x2_sg U53552 ( .A(n47475), .B(n57862), .X(n22751) );
  nand_x4_sg U53553 ( .A(n25754), .B(n25755), .X(n24111) );
  nand_x4_sg U53554 ( .A(n25242), .B(n25243), .X(n24016) );
  nand_x4_sg U53555 ( .A(n25002), .B(n25003), .X(n23976) );
  nand_x2_sg U53556 ( .A(n56971), .B(n57166), .X(n34221) );
  nand_x2_sg U53557 ( .A(n68477), .B(n68478), .X(n32491) );
  inv_x4_sg U53558 ( .A(n56987), .X(n68477) );
  nand_x2_sg U53559 ( .A(n68577), .B(n68578), .X(n32048) );
  inv_x4_sg U53560 ( .A(n56983), .X(n68577) );
  inv_x2_sg U53561 ( .A(n47476), .X(n47477) );
  inv_x2_sg U53562 ( .A(n47478), .X(n47479) );
  inv_x2_sg U53563 ( .A(n47480), .X(n47481) );
  inv_x2_sg U53564 ( .A(\shifter_0/reg_i_4 [0]), .X(n47600) );
  inv_x2_sg U53565 ( .A(\shifter_0/reg_i_4 [1]), .X(n47602) );
  inv_x2_sg U53566 ( .A(\shifter_0/reg_i_4 [5]), .X(n47604) );
  inv_x2_sg U53567 ( .A(\shifter_0/reg_i_12 [0]), .X(n47616) );
  inv_x2_sg U53568 ( .A(\shifter_0/reg_i_12 [1]), .X(n47618) );
  inv_x2_sg U53569 ( .A(\shifter_0/reg_i_12 [5]), .X(n47620) );
  inv_x2_sg U53570 ( .A(\shifter_0/reg_i_13 [0]), .X(n47622) );
  inv_x2_sg U53571 ( .A(\shifter_0/reg_i_13 [1]), .X(n47624) );
  inv_x2_sg U53572 ( .A(\shifter_0/reg_i_13 [5]), .X(n47626) );
  inv_x2_sg U53573 ( .A(\shifter_0/reg_i_14 [19]), .X(n56672) );
  inv_x2_sg U53574 ( .A(\shifter_0/reg_w_4 [0]), .X(n47606) );
  inv_x2_sg U53575 ( .A(\shifter_0/reg_w_4 [1]), .X(n47608) );
  inv_x2_sg U53576 ( .A(\shifter_0/reg_w_4 [5]), .X(n47610) );
  inv_x2_sg U53577 ( .A(\shifter_0/reg_w_10 [0]), .X(n47526) );
  inv_x2_sg U53578 ( .A(\shifter_0/reg_w_10 [1]), .X(n47528) );
  inv_x2_sg U53579 ( .A(\shifter_0/reg_w_10 [5]), .X(n47530) );
  inv_x2_sg U53580 ( .A(\shifter_0/reg_w_11 [0]), .X(n47630) );
  inv_x2_sg U53581 ( .A(\shifter_0/reg_w_11 [1]), .X(n47632) );
  inv_x2_sg U53582 ( .A(\shifter_0/reg_w_11 [5]), .X(n47634) );
  inv_x2_sg U53583 ( .A(\shifter_0/reg_w_12 [0]), .X(n47636) );
  inv_x2_sg U53584 ( .A(\shifter_0/reg_w_12 [1]), .X(n47638) );
  inv_x2_sg U53585 ( .A(\shifter_0/reg_w_12 [5]), .X(n47640) );
  inv_x2_sg U53586 ( .A(\shifter_0/reg_w_13 [0]), .X(n47642) );
  inv_x2_sg U53587 ( .A(\shifter_0/reg_w_13 [1]), .X(n47644) );
  inv_x2_sg U53588 ( .A(\shifter_0/reg_w_13 [5]), .X(n47646) );
  inv_x2_sg U53589 ( .A(\shifter_0/reg_w_14 [1]), .X(n56696) );
  inv_x2_sg U53590 ( .A(\shifter_0/reg_w_14 [6]), .X(n47650) );
  inv_x2_sg U53591 ( .A(\shifter_0/reg_i_9 [2]), .X(n56740) );
  inv_x2_sg U53592 ( .A(\shifter_0/reg_i_10 [0]), .X(n47542) );
  inv_x2_sg U53593 ( .A(\shifter_0/reg_i_10 [2]), .X(n56748) );
  inv_x2_sg U53594 ( .A(\shifter_0/reg_i_10 [5]), .X(n47546) );
  inv_x2_sg U53595 ( .A(\shifter_0/reg_i_11 [0]), .X(n47652) );
  inv_x2_sg U53596 ( .A(\shifter_0/reg_i_11 [1]), .X(n47654) );
  inv_x2_sg U53597 ( .A(\shifter_0/reg_i_11 [5]), .X(n47656) );
  inv_x2_sg U53598 ( .A(\shifter_0/reg_i_14 [6]), .X(n47660) );
  inv_x2_sg U53599 ( .A(\shifter_0/reg_i_14 [10]), .X(n47662) );
  inv_x2_sg U53600 ( .A(\shifter_0/reg_w_14 [10]), .X(n47664) );
  inv_x2_sg U53601 ( .A(\shifter_0/reg_i_5 [0]), .X(n47672) );
  inv_x2_sg U53602 ( .A(\shifter_0/reg_i_5 [1]), .X(n47674) );
  inv_x2_sg U53603 ( .A(\shifter_0/reg_i_5 [5]), .X(n47676) );
  inv_x2_sg U53604 ( .A(\shifter_0/reg_i_12 [16]), .X(n47678) );
  inv_x2_sg U53605 ( .A(\shifter_0/reg_i_13 [16]), .X(n47680) );
  inv_x2_sg U53606 ( .A(\shifter_0/reg_i_14 [16]), .X(n47682) );
  inv_x2_sg U53607 ( .A(\shifter_0/reg_w_5 [0]), .X(n47684) );
  inv_x2_sg U53608 ( .A(\shifter_0/reg_w_5 [1]), .X(n47686) );
  inv_x2_sg U53609 ( .A(\shifter_0/reg_w_5 [5]), .X(n47688) );
  inv_x2_sg U53610 ( .A(\shifter_0/reg_w_12 [16]), .X(n47690) );
  inv_x2_sg U53611 ( .A(\shifter_0/reg_w_13 [16]), .X(n47692) );
  inv_x2_sg U53612 ( .A(\shifter_0/reg_i_5 [17]), .X(n47694) );
  inv_x2_sg U53613 ( .A(\shifter_0/reg_w_5 [17]), .X(n47696) );
  inv_x2_sg U53614 ( .A(\shifter_0/reg_i_10 [17]), .X(n56852) );
  inv_x2_sg U53615 ( .A(\shifter_0/reg_i_11 [17]), .X(n47700) );
  inv_x2_sg U53616 ( .A(\shifter_0/reg_w_9 [17]), .X(n47554) );
  inv_x2_sg U53617 ( .A(\shifter_0/reg_w_10 [17]), .X(n56856) );
  inv_x2_sg U53618 ( .A(\shifter_0/reg_w_11 [18]), .X(n51412) );
  inv_x2_sg U53619 ( .A(\shifter_0/reg_w_14 [17]), .X(n47706) );
  nor_x2_sg U53620 ( .A(n57168), .B(n51523), .X(n34175) );
  inv_x2_sg U53621 ( .A(\shifter_0/reg_i_2 [6]), .X(n55224) );
  inv_x2_sg U53622 ( .A(\shifter_0/reg_i_2 [10]), .X(n55228) );
  inv_x2_sg U53623 ( .A(\shifter_0/reg_i_6 [0]), .X(n47556) );
  inv_x2_sg U53624 ( .A(\shifter_0/reg_i_6 [1]), .X(n47558) );
  inv_x2_sg U53625 ( .A(\shifter_0/reg_i_6 [5]), .X(n47560) );
  inv_x2_sg U53626 ( .A(\shifter_0/reg_w_2 [6]), .X(n55236) );
  inv_x2_sg U53627 ( .A(\shifter_0/reg_w_2 [10]), .X(n55240) );
  inv_x2_sg U53628 ( .A(\shifter_0/reg_w_6 [0]), .X(n47562) );
  inv_x2_sg U53629 ( .A(\shifter_0/reg_w_6 [1]), .X(n47564) );
  inv_x2_sg U53630 ( .A(\shifter_0/reg_w_6 [5]), .X(n47566) );
  inv_x2_sg U53631 ( .A(\shifter_0/reg_i_3 [0]), .X(n47720) );
  inv_x2_sg U53632 ( .A(\shifter_0/reg_i_3 [1]), .X(n47722) );
  inv_x2_sg U53633 ( .A(\shifter_0/reg_i_3 [5]), .X(n47724) );
  inv_x2_sg U53634 ( .A(\shifter_0/reg_w_3 [1]), .X(n47728) );
  inv_x2_sg U53635 ( .A(\shifter_0/reg_w_3 [5]), .X(n47730) );
  inv_x2_sg U53636 ( .A(\shifter_0/reg_i_6 [17]), .X(n47732) );
  inv_x2_sg U53637 ( .A(\shifter_0/reg_w_3 [0]), .X(n47726) );
  inv_x2_sg U53638 ( .A(\shifter_0/reg_w_2 [17]), .X(n55250) );
  inv_x2_sg U53639 ( .A(\shifter_0/reg_w_6 [17]), .X(n47734) );
  inv_x2_sg U53640 ( .A(\shifter_0/reg_i_3 [16]), .X(n47736) );
  inv_x2_sg U53641 ( .A(\shifter_0/reg_w_3 [16]), .X(n47738) );
  nor_x2_sg U53642 ( .A(n57033), .B(n57152), .X(n23087) );
  nor_x2_sg U53643 ( .A(n57017), .B(n22988), .X(n23065) );
  nor_x2_sg U53644 ( .A(n47753), .B(n57153), .X(n23043) );
  nor_x2_sg U53645 ( .A(n57039), .B(n57158), .X(n22860) );
  nor_x2_sg U53646 ( .A(n57013), .B(n22761), .X(n22838) );
  nor_x2_sg U53647 ( .A(n47747), .B(n57159), .X(n22816) );
  inv_x4_sg U53648 ( .A(n24878), .X(n67279) );
  inv_x4_sg U53649 ( .A(n25930), .X(n67457) );
  inv_x4_sg U53650 ( .A(n25690), .X(n67465) );
  inv_x4_sg U53651 ( .A(n25510), .X(n67471) );
  inv_x4_sg U53652 ( .A(n25178), .X(n67269) );
  nor_x2_sg U53653 ( .A(n68388), .B(n32372), .X(n32382) );
  inv_x4_sg U53654 ( .A(n32386), .X(n68388) );
  nand_x2_sg U53655 ( .A(n68494), .B(n68495), .X(n32038) );
  inv_x4_sg U53656 ( .A(n55057), .X(n68495) );
  inv_x2_sg U53657 ( .A(n57085), .X(n58493) );
  inv_x2_sg U53658 ( .A(n57081), .X(n58532) );
  inv_x2_sg U53659 ( .A(n57089), .X(n58542) );
  nor_x2_sg U53660 ( .A(n31951), .B(n68572), .X(n31950) );
  nor_x2_sg U53661 ( .A(n23546), .B(n58384), .X(n58385) );
  nor_x2_sg U53662 ( .A(n57097), .B(n47775), .X(n23546) );
  inv_x1_sg U53663 ( .A(n35560), .X(n68260) );
  inv_x1_sg U53664 ( .A(n35538), .X(n68258) );
  inv_x1_sg U53665 ( .A(n35615), .X(n68247) );
  inv_x1_sg U53666 ( .A(n35576), .X(n68252) );
  inv_x1_sg U53667 ( .A(n35578), .X(n68251) );
  inv_x1_sg U53668 ( .A(n35570), .X(n68233) );
  inv_x1_sg U53669 ( .A(n35572), .X(n68232) );
  inv_x1_sg U53670 ( .A(n35535), .X(n68240) );
  nand_x2_sg U53671 ( .A(n47481), .B(n57862), .X(n23113) );
  nand_x2_sg U53672 ( .A(n47479), .B(n57862), .X(n23014) );
  nand_x2_sg U53673 ( .A(n47473), .B(n57862), .X(n22930) );
  nand_x2_sg U53674 ( .A(n47455), .B(n57862), .X(n22831) );
  nand_x2_sg U53675 ( .A(n47477), .B(n57862), .X(n22787) );
  nand_x4_sg U53676 ( .A(n25634), .B(n25635), .X(n24091) );
  nand_x4_sg U53677 ( .A(n25454), .B(n25455), .X(n24061) );
  nand_x4_sg U53678 ( .A(n25032), .B(n25033), .X(n23981) );
  nand_x4_sg U53679 ( .A(n24821), .B(n24822), .X(n23945) );
  nand_x4_sg U53680 ( .A(n25904), .B(n25905), .X(n24136) );
  nand_x4_sg U53681 ( .A(n25302), .B(n25303), .X(n24026) );
  nand_x2_sg U53682 ( .A(n68405), .B(n68406), .X(n32480) );
  nor_x2_sg U53683 ( .A(n24829), .B(n68406), .X(n25970) );
  inv_x4_sg U53684 ( .A(n55037), .X(n68406) );
  nand_x2_sg U53685 ( .A(n68408), .B(n68409), .X(n32644) );
  nor_x2_sg U53686 ( .A(n68409), .B(n57102), .X(n25551) );
  inv_x4_sg U53687 ( .A(n55287), .X(n68409) );
  nand_x2_sg U53688 ( .A(n68399), .B(n68400), .X(n32469) );
  nor_x2_sg U53689 ( .A(n24829), .B(n68400), .X(n25550) );
  inv_x4_sg U53690 ( .A(n55025), .X(n68400) );
  inv_x2_sg U53691 ( .A(\shifter_0/reg_i_4 [2]), .X(n51134) );
  inv_x2_sg U53692 ( .A(\shifter_0/reg_i_4 [6]), .X(n51136) );
  inv_x2_sg U53693 ( .A(\shifter_0/reg_i_4 [10]), .X(n51138) );
  inv_x2_sg U53694 ( .A(\shifter_0/reg_i_12 [2]), .X(n51200) );
  inv_x2_sg U53695 ( .A(\shifter_0/reg_i_12 [6]), .X(n51202) );
  inv_x2_sg U53696 ( .A(\shifter_0/reg_i_12 [10]), .X(n51204) );
  inv_x2_sg U53697 ( .A(\shifter_0/reg_i_13 [2]), .X(n51206) );
  inv_x2_sg U53698 ( .A(\shifter_0/reg_i_13 [6]), .X(n51208) );
  inv_x2_sg U53699 ( .A(\shifter_0/reg_i_13 [10]), .X(n51210) );
  inv_x2_sg U53700 ( .A(\shifter_0/reg_i_14 [14]), .X(n47628) );
  inv_x2_sg U53701 ( .A(\shifter_0/reg_w_4 [2]), .X(n51140) );
  inv_x2_sg U53702 ( .A(\shifter_0/reg_w_4 [6]), .X(n51142) );
  inv_x2_sg U53703 ( .A(\shifter_0/reg_w_4 [10]), .X(n51144) );
  inv_x2_sg U53704 ( .A(\shifter_0/reg_w_9 [2]), .X(n56674) );
  inv_x2_sg U53705 ( .A(n47482), .X(n47483) );
  inv_x2_sg U53706 ( .A(\shifter_0/reg_w_9 [6]), .X(n56676) );
  inv_x2_sg U53707 ( .A(\shifter_0/reg_w_10 [2]), .X(n56678) );
  inv_x2_sg U53708 ( .A(\shifter_0/reg_w_10 [6]), .X(n56680) );
  inv_x2_sg U53709 ( .A(\shifter_0/reg_w_11 [7]), .X(n56682) );
  inv_x2_sg U53710 ( .A(\shifter_0/reg_w_12 [2]), .X(n51222) );
  inv_x2_sg U53711 ( .A(\shifter_0/reg_w_12 [6]), .X(n51224) );
  inv_x2_sg U53712 ( .A(\shifter_0/reg_w_12 [10]), .X(n51226) );
  inv_x2_sg U53713 ( .A(\shifter_0/reg_w_13 [2]), .X(n51228) );
  inv_x2_sg U53714 ( .A(\shifter_0/reg_w_13 [6]), .X(n51230) );
  inv_x2_sg U53715 ( .A(\shifter_0/reg_w_13 [10]), .X(n51232) );
  inv_x2_sg U53716 ( .A(\shifter_0/reg_w_14 [2]), .X(n47648) );
  inv_x2_sg U53717 ( .A(\shifter_0/reg_w_14 [7]), .X(n51234) );
  inv_x2_sg U53718 ( .A(\shifter_0/reg_i_12 [14]), .X(n51236) );
  inv_x2_sg U53719 ( .A(\shifter_0/reg_i_13 [14]), .X(n51238) );
  inv_x2_sg U53720 ( .A(\shifter_0/reg_w_12 [14]), .X(n51240) );
  inv_x2_sg U53721 ( .A(\shifter_0/reg_w_13 [14]), .X(n51242) );
  inv_x2_sg U53722 ( .A(\shifter_0/reg_i_12 [3]), .X(n51244) );
  inv_x2_sg U53723 ( .A(\shifter_0/reg_i_12 [8]), .X(n51246) );
  inv_x2_sg U53724 ( .A(\shifter_0/reg_i_12 [12]), .X(n51248) );
  inv_x2_sg U53725 ( .A(\shifter_0/reg_i_13 [3]), .X(n51250) );
  inv_x2_sg U53726 ( .A(\shifter_0/reg_i_13 [8]), .X(n51252) );
  inv_x2_sg U53727 ( .A(\shifter_0/reg_i_13 [12]), .X(n51254) );
  inv_x2_sg U53728 ( .A(\shifter_0/reg_w_10 [3]), .X(n56722) );
  inv_x2_sg U53729 ( .A(\shifter_0/reg_w_11 [3]), .X(n51262) );
  inv_x2_sg U53730 ( .A(\shifter_0/reg_w_12 [3]), .X(n51264) );
  inv_x2_sg U53731 ( .A(\shifter_0/reg_w_12 [8]), .X(n51266) );
  inv_x2_sg U53732 ( .A(\shifter_0/reg_w_12 [12]), .X(n51268) );
  inv_x2_sg U53733 ( .A(\shifter_0/reg_w_13 [3]), .X(n51270) );
  inv_x2_sg U53734 ( .A(\shifter_0/reg_w_13 [8]), .X(n51272) );
  inv_x2_sg U53735 ( .A(\shifter_0/reg_w_13 [12]), .X(n51274) );
  inv_x2_sg U53736 ( .A(n47484), .X(n47485) );
  inv_x2_sg U53737 ( .A(\shifter_0/reg_i_9 [6]), .X(n56742) );
  inv_x2_sg U53738 ( .A(\shifter_0/reg_i_9 [10]), .X(n56744) );
  inv_x2_sg U53739 ( .A(\shifter_0/reg_i_9 [15]), .X(n51282) );
  inv_x2_sg U53740 ( .A(\shifter_0/reg_i_10 [6]), .X(n56750) );
  inv_x2_sg U53741 ( .A(\shifter_0/reg_i_10 [10]), .X(n56752) );
  inv_x2_sg U53742 ( .A(\shifter_0/reg_i_10 [14]), .X(n51288) );
  inv_x2_sg U53743 ( .A(\shifter_0/reg_i_11 [2]), .X(n51290) );
  inv_x2_sg U53744 ( .A(\shifter_0/reg_i_11 [7]), .X(n56756) );
  inv_x2_sg U53745 ( .A(\shifter_0/reg_i_11 [11]), .X(n56758) );
  inv_x2_sg U53746 ( .A(\shifter_0/reg_i_14 [1]), .X(n47658) );
  inv_x2_sg U53747 ( .A(\shifter_0/reg_i_14 [7]), .X(n51300) );
  inv_x2_sg U53748 ( .A(\shifter_0/reg_i_14 [11]), .X(n51302) );
  inv_x2_sg U53749 ( .A(\shifter_0/reg_w_9 [10]), .X(n56762) );
  inv_x2_sg U53750 ( .A(\shifter_0/reg_w_9 [15]), .X(n51306) );
  inv_x2_sg U53751 ( .A(\shifter_0/reg_w_10 [10]), .X(n56766) );
  inv_x2_sg U53752 ( .A(\shifter_0/reg_w_10 [14]), .X(n51310) );
  inv_x2_sg U53753 ( .A(\shifter_0/reg_w_11 [11]), .X(n56770) );
  inv_x2_sg U53754 ( .A(\shifter_0/reg_w_14 [11]), .X(n51316) );
  inv_x2_sg U53755 ( .A(\shifter_0/reg_w_14 [14]), .X(n47666) );
  inv_x2_sg U53756 ( .A(\shifter_0/reg_i_10 [19]), .X(n51322) );
  inv_x2_sg U53757 ( .A(\shifter_0/reg_w_11 [19]), .X(n56776) );
  inv_x2_sg U53758 ( .A(\shifter_0/reg_i_9 [8]), .X(n56792) );
  inv_x2_sg U53759 ( .A(\shifter_0/reg_i_10 [3]), .X(n56796) );
  inv_x2_sg U53760 ( .A(\shifter_0/reg_i_10 [12]), .X(n56800) );
  inv_x2_sg U53761 ( .A(\shifter_0/reg_i_11 [3]), .X(n51354) );
  inv_x2_sg U53762 ( .A(\shifter_0/reg_i_11 [9]), .X(n56804) );
  inv_x2_sg U53763 ( .A(\shifter_0/reg_i_11 [12]), .X(n51358) );
  inv_x2_sg U53764 ( .A(\shifter_0/reg_i_14 [8]), .X(n47668) );
  inv_x2_sg U53765 ( .A(n47486), .X(n47487) );
  inv_x2_sg U53766 ( .A(\shifter_0/reg_w_9 [8]), .X(n56810) );
  inv_x2_sg U53767 ( .A(\shifter_0/reg_w_10 [12]), .X(n56816) );
  inv_x2_sg U53768 ( .A(\shifter_0/reg_w_11 [9]), .X(n56818) );
  inv_x2_sg U53769 ( .A(\shifter_0/reg_w_11 [12]), .X(n51374) );
  inv_x2_sg U53770 ( .A(\shifter_0/reg_w_14 [8]), .X(n47670) );
  inv_x2_sg U53771 ( .A(\shifter_0/reg_i_5 [2]), .X(n51380) );
  inv_x2_sg U53772 ( .A(\shifter_0/reg_i_5 [6]), .X(n51382) );
  inv_x2_sg U53773 ( .A(\shifter_0/reg_i_5 [10]), .X(n51384) );
  inv_x2_sg U53774 ( .A(\shifter_0/reg_i_12 [17]), .X(n51388) );
  inv_x2_sg U53775 ( .A(\shifter_0/reg_i_13 [17]), .X(n51390) );
  inv_x2_sg U53776 ( .A(\shifter_0/reg_i_14 [18]), .X(n56834) );
  inv_x2_sg U53777 ( .A(\shifter_0/reg_w_5 [2]), .X(n51394) );
  inv_x2_sg U53778 ( .A(\shifter_0/reg_w_5 [6]), .X(n51396) );
  inv_x2_sg U53779 ( .A(\shifter_0/reg_w_5 [10]), .X(n51398) );
  inv_x2_sg U53780 ( .A(\shifter_0/reg_w_12 [18]), .X(n56842) );
  inv_x2_sg U53781 ( .A(\shifter_0/reg_w_13 [17]), .X(n51404) );
  inv_x2_sg U53782 ( .A(\shifter_0/reg_i_5 [18]), .X(n51406) );
  inv_x2_sg U53783 ( .A(\shifter_0/reg_w_5 [18]), .X(n51408) );
  inv_x2_sg U53784 ( .A(\shifter_0/reg_i_9 [18]), .X(n56850) );
  inv_x2_sg U53785 ( .A(\shifter_0/reg_i_10 [18]), .X(n47698) );
  inv_x2_sg U53786 ( .A(n47488), .X(n47489) );
  inv_x2_sg U53787 ( .A(\shifter_0/reg_w_9 [18]), .X(n56854) );
  inv_x2_sg U53788 ( .A(\shifter_0/reg_w_10 [18]), .X(n47702) );
  inv_x2_sg U53789 ( .A(\shifter_0/reg_w_14 [18]), .X(n56858) );
  inv_x2_sg U53790 ( .A(\shifter_0/reg_i_11 [16]), .X(n56860) );
  inv_x2_sg U53791 ( .A(\shifter_0/reg_w_11 [16]), .X(n56862) );
  nor_x2_sg U53792 ( .A(n57168), .B(n51525), .X(n34088) );
  inv_x2_sg U53793 ( .A(\shifter_0/pointer [2]), .X(n53714) );
  inv_x2_sg U53794 ( .A(\shifter_0/reg_i_2 [0]), .X(n47506) );
  inv_x2_sg U53795 ( .A(\shifter_0/reg_i_2 [1]), .X(n51150) );
  inv_x2_sg U53796 ( .A(\shifter_0/reg_i_2 [4]), .X(n51152) );
  inv_x2_sg U53797 ( .A(\shifter_0/reg_i_2 [5]), .X(n47508) );
  inv_x2_sg U53798 ( .A(\shifter_0/reg_i_6 [2]), .X(n56868) );
  inv_x2_sg U53799 ( .A(\shifter_0/reg_i_6 [6]), .X(n56870) );
  inv_x2_sg U53800 ( .A(\shifter_0/reg_i_6 [10]), .X(n56872) );
  inv_x2_sg U53801 ( .A(\shifter_0/reg_w_2 [0]), .X(n47510) );
  inv_x2_sg U53802 ( .A(\shifter_0/reg_w_2 [1]), .X(n47512) );
  inv_x2_sg U53803 ( .A(\shifter_0/reg_w_2 [5]), .X(n47514) );
  inv_x2_sg U53804 ( .A(\shifter_0/reg_w_6 [2]), .X(n56876) );
  inv_x2_sg U53805 ( .A(\shifter_0/reg_w_6 [6]), .X(n56878) );
  inv_x2_sg U53806 ( .A(\shifter_0/reg_w_6 [10]), .X(n56880) );
  inv_x2_sg U53807 ( .A(\shifter_0/reg_i_6 [3]), .X(n47708) );
  inv_x2_sg U53808 ( .A(\shifter_0/reg_i_6 [8]), .X(n47710) );
  inv_x2_sg U53809 ( .A(\shifter_0/reg_i_6 [12]), .X(n47712) );
  inv_x2_sg U53810 ( .A(\shifter_0/reg_w_6 [3]), .X(n47714) );
  inv_x2_sg U53811 ( .A(\shifter_0/reg_w_6 [8]), .X(n47716) );
  inv_x2_sg U53812 ( .A(\shifter_0/reg_w_6 [12]), .X(n47718) );
  inv_x2_sg U53813 ( .A(\shifter_0/reg_i_3 [2]), .X(n51452) );
  inv_x2_sg U53814 ( .A(\shifter_0/reg_i_3 [6]), .X(n51454) );
  inv_x2_sg U53815 ( .A(\shifter_0/reg_i_3 [10]), .X(n51456) );
  inv_x2_sg U53816 ( .A(\shifter_0/reg_w_3 [2]), .X(n51458) );
  inv_x2_sg U53817 ( .A(\shifter_0/reg_w_3 [6]), .X(n51460) );
  inv_x2_sg U53818 ( .A(\shifter_0/reg_w_3 [10]), .X(n51462) );
  inv_x2_sg U53819 ( .A(\shifter_0/reg_i_2 [16]), .X(n47516) );
  inv_x2_sg U53820 ( .A(\shifter_0/reg_i_3 [12]), .X(n51468) );
  inv_x2_sg U53821 ( .A(\shifter_0/reg_i_6 [18]), .X(n51472) );
  inv_x2_sg U53822 ( .A(\shifter_0/reg_w_2 [16]), .X(n47518) );
  inv_x2_sg U53823 ( .A(\shifter_0/reg_w_3 [3]), .X(n51474) );
  inv_x2_sg U53824 ( .A(\shifter_0/reg_w_3 [8]), .X(n51476) );
  inv_x2_sg U53825 ( .A(\shifter_0/reg_w_6 [18]), .X(n51482) );
  inv_x2_sg U53826 ( .A(\shifter_0/reg_i_3 [17]), .X(n51484) );
  inv_x2_sg U53827 ( .A(\shifter_0/reg_w_3 [17]), .X(n51486) );
  inv_x2_sg U53828 ( .A(\filter_0/N13 ), .X(n51056) );
  nor_x2_sg U53829 ( .A(n51513), .B(n57153), .X(n23175) );
  nor_x2_sg U53830 ( .A(n47751), .B(n22988), .X(n22999) );
  nor_x2_sg U53831 ( .A(n47749), .B(n57152), .X(n22986) );
  nor_x2_sg U53832 ( .A(n51519), .B(n57159), .X(n22948) );
  nor_x2_sg U53833 ( .A(n47745), .B(n22761), .X(n22772) );
  nor_x2_sg U53834 ( .A(n47743), .B(n57158), .X(n22759) );
  inv_x4_sg U53835 ( .A(n25810), .X(n67461) );
  inv_x4_sg U53836 ( .A(n25660), .X(n67466) );
  inv_x4_sg U53837 ( .A(n25358), .X(n67263) );
  inv_x4_sg U53838 ( .A(n25088), .X(n67272) );
  inv_x4_sg U53839 ( .A(n24938), .X(n67277) );
  nor_x4_sg U53840 ( .A(n57113), .B(n57168), .X(n32803) );
  nand_x4_sg U53841 ( .A(n33396), .B(n34042), .X(n34041) );
  inv_x4_sg U53842 ( .A(n22548), .X(n67160) );
  inv_x4_sg U53843 ( .A(n24692), .X(n67101) );
  nor_x2_sg U53844 ( .A(n24692), .B(n57099), .X(n58121) );
  nand_x4_sg U53845 ( .A(n23308), .B(n22471), .X(n24692) );
  inv_x4_sg U53846 ( .A(n32482), .X(n68265) );
  nand_x4_sg U53847 ( .A(n68265), .B(n32436), .X(n32368) );
  inv_x4_sg U53848 ( .A(n47490), .X(n47491) );
  nand_x4_sg U53849 ( .A(n47491), .B(n31993), .X(n31968) );
  inv_x2_sg U53850 ( .A(n51551), .X(n58499) );
  inv_x2_sg U53851 ( .A(n57075), .X(n58513) );
  inv_x2_sg U53852 ( .A(n51547), .X(n58520) );
  inv_x2_sg U53853 ( .A(n51553), .X(n58548) );
  inv_x2_sg U53854 ( .A(n57071), .X(n58562) );
  inv_x2_sg U53855 ( .A(n51545), .X(n58569) );
  inv_x2_sg U53856 ( .A(n47773), .X(n58576) );
  nor_x2_sg U53857 ( .A(n57097), .B(n29336), .X(n23309) );
  nor_x8_sg U53858 ( .A(n68574), .B(n68572), .X(n29336) );
  nand_x4_sg U53859 ( .A(n26178), .B(n67574), .X(n26177) );
  inv_x4_sg U53860 ( .A(n34222), .X(n67574) );
  nor_x2_sg U53861 ( .A(n32083), .B(n32084), .X(n32072) );
  nor_x2_sg U53862 ( .A(n32074), .B(n68556), .X(n32073) );
  nand_x4_sg U53863 ( .A(n57958), .B(n57957), .X(n57962) );
  nand_x4_sg U53864 ( .A(n25874), .B(n25875), .X(n24131) );
  nand_x4_sg U53865 ( .A(n25724), .B(n25725), .X(n24106) );
  nand_x4_sg U53866 ( .A(n25424), .B(n25425), .X(n24055) );
  nand_x4_sg U53867 ( .A(n25272), .B(n25273), .X(n24021) );
  nand_x4_sg U53868 ( .A(n24852), .B(n24853), .X(n23951) );
  nand_x2_sg U53869 ( .A(n68412), .B(n68413), .X(n32652) );
  nor_x2_sg U53870 ( .A(n68413), .B(n57102), .X(n25821) );
  inv_x4_sg U53871 ( .A(n55295), .X(n68413) );
  nand_x2_sg U53872 ( .A(n68403), .B(n68404), .X(n32477) );
  nor_x2_sg U53873 ( .A(n24829), .B(n68404), .X(n25820) );
  inv_x4_sg U53874 ( .A(n55033), .X(n68404) );
  nand_x2_sg U53875 ( .A(n68410), .B(n68411), .X(n32647) );
  nor_x2_sg U53876 ( .A(n68411), .B(n57102), .X(n25701) );
  inv_x4_sg U53877 ( .A(n55291), .X(n68411) );
  nand_x2_sg U53878 ( .A(n68401), .B(n68402), .X(n32472) );
  nor_x2_sg U53879 ( .A(n24829), .B(n68402), .X(n25700) );
  inv_x4_sg U53880 ( .A(n55029), .X(n68402) );
  nand_x2_sg U53881 ( .A(n68501), .B(n68502), .X(n32207) );
  nor_x2_sg U53882 ( .A(n68502), .B(n57102), .X(n25219) );
  inv_x4_sg U53883 ( .A(n55307), .X(n68502) );
  nand_x2_sg U53884 ( .A(n68492), .B(n68493), .X(n32035) );
  nor_x2_sg U53885 ( .A(n24829), .B(n68493), .X(n25218) );
  inv_x4_sg U53886 ( .A(n55053), .X(n68493) );
  nand_x2_sg U53887 ( .A(n68499), .B(n68500), .X(n32202) );
  nor_x2_sg U53888 ( .A(n68500), .B(n57102), .X(n25099) );
  inv_x4_sg U53889 ( .A(n55303), .X(n68500) );
  nand_x2_sg U53890 ( .A(n68490), .B(n68491), .X(n32030) );
  nor_x2_sg U53891 ( .A(n24829), .B(n68491), .X(n25098) );
  inv_x4_sg U53892 ( .A(n55049), .X(n68491) );
  nand_x2_sg U53893 ( .A(n68497), .B(n68498), .X(n32199) );
  nor_x2_sg U53894 ( .A(n68498), .B(n57102), .X(n24949) );
  inv_x4_sg U53895 ( .A(n55299), .X(n68498) );
  nand_x2_sg U53896 ( .A(n68488), .B(n68489), .X(n32027) );
  nor_x2_sg U53897 ( .A(n24829), .B(n68489), .X(n24948) );
  inv_x4_sg U53898 ( .A(n55045), .X(n68489) );
  nand_x2_sg U53899 ( .A(n68479), .B(n68480), .X(n32495) );
  inv_x4_sg U53900 ( .A(n56991), .X(n68479) );
  inv_x4_sg U53901 ( .A(n56989), .X(n68478) );
  nand_x2_sg U53902 ( .A(n68414), .B(n68415), .X(n32655) );
  nor_x2_sg U53903 ( .A(n68415), .B(n57102), .X(n25971) );
  inv_x4_sg U53904 ( .A(n55311), .X(n68415) );
  nand_x2_sg U53905 ( .A(n68503), .B(n68504), .X(n32210) );
  nor_x2_sg U53906 ( .A(n68504), .B(n57102), .X(n25369) );
  inv_x4_sg U53907 ( .A(n55315), .X(n68504) );
  nand_x2_sg U53908 ( .A(n68579), .B(n68580), .X(n32052) );
  inv_x4_sg U53909 ( .A(n56979), .X(n68579) );
  nand_x2_sg U53910 ( .A(n68432), .B(n68433), .X(n32616) );
  nor_x2_sg U53911 ( .A(n68432), .B(n57103), .X(n58147) );
  inv_x4_sg U53912 ( .A(n55039), .X(n68432) );
  nand_x2_sg U53913 ( .A(n68522), .B(n68523), .X(n32171) );
  nor_x2_sg U53914 ( .A(n68522), .B(n58638), .X(n58247) );
  inv_x4_sg U53915 ( .A(n55059), .X(n68522) );
  inv_x4_sg U53916 ( .A(n56985), .X(n68578) );
  inv_x2_sg U53917 ( .A(\mask_0/reg_i_mask [1]), .X(n51070) );
  inv_x2_sg U53918 ( .A(\mask_0/reg_i_mask [2]), .X(n51072) );
  inv_x2_sg U53919 ( .A(\mask_0/reg_i_mask [3]), .X(n51074) );
  inv_x2_sg U53920 ( .A(\mask_0/reg_i_mask [6]), .X(n51076) );
  inv_x2_sg U53921 ( .A(\mask_0/reg_i_mask [7]), .X(n51078) );
  inv_x2_sg U53922 ( .A(\mask_0/reg_i_mask [8]), .X(n51080) );
  inv_x2_sg U53923 ( .A(\mask_0/reg_i_mask [9]), .X(n51082) );
  inv_x2_sg U53924 ( .A(\mask_0/reg_i_mask [10]), .X(n51084) );
  inv_x2_sg U53925 ( .A(\mask_0/reg_i_mask [11]), .X(n51086) );
  inv_x2_sg U53926 ( .A(\mask_0/reg_i_mask [12]), .X(n51088) );
  inv_x2_sg U53927 ( .A(\mask_0/reg_i_mask [13]), .X(n51090) );
  inv_x2_sg U53928 ( .A(\mask_0/reg_i_mask [14]), .X(n51092) );
  inv_x2_sg U53929 ( .A(\mask_0/reg_i_mask [15]), .X(n51094) );
  inv_x2_sg U53930 ( .A(\mask_0/reg_i_mask [16]), .X(n51096) );
  inv_x2_sg U53931 ( .A(\mask_0/reg_i_mask [18]), .X(n51098) );
  inv_x2_sg U53932 ( .A(\mask_0/reg_i_mask [19]), .X(n51100) );
  inv_x2_sg U53933 ( .A(\mask_0/reg_i_mask [20]), .X(n51102) );
  inv_x2_sg U53934 ( .A(\mask_0/reg_i_mask [21]), .X(n51104) );
  inv_x2_sg U53935 ( .A(\mask_0/reg_i_mask [22]), .X(n51106) );
  inv_x2_sg U53936 ( .A(\mask_0/reg_i_mask [23]), .X(n51108) );
  inv_x2_sg U53937 ( .A(\mask_0/reg_i_mask [24]), .X(n51110) );
  inv_x2_sg U53938 ( .A(\mask_0/reg_i_mask [25]), .X(n51112) );
  inv_x2_sg U53939 ( .A(\mask_0/reg_i_mask [26]), .X(n51114) );
  inv_x2_sg U53940 ( .A(\mask_0/reg_i_mask [27]), .X(n51116) );
  inv_x2_sg U53941 ( .A(\mask_0/reg_w_mask [0]), .X(n51118) );
  inv_x2_sg U53942 ( .A(\mask_0/reg_w_mask [4]), .X(n51120) );
  inv_x2_sg U53943 ( .A(\mask_0/reg_w_mask [5]), .X(n51122) );
  inv_x2_sg U53944 ( .A(\mask_0/reg_w_mask [17]), .X(n51124) );
  inv_x2_sg U53945 ( .A(\mask_0/reg_w_mask [28]), .X(n51126) );
  inv_x2_sg U53946 ( .A(\mask_0/reg_w_mask [29]), .X(n51128) );
  inv_x2_sg U53947 ( .A(\mask_0/reg_w_mask [30]), .X(n51130) );
  inv_x2_sg U53948 ( .A(\mask_0/reg_w_mask [31]), .X(n51132) );
  inv_x2_sg U53949 ( .A(\filter_0/reg_i_11 [13]), .X(n55782) );
  inv_x2_sg U53950 ( .A(\shifter_0/reg_i_4 [7]), .X(n55072) );
  inv_x2_sg U53951 ( .A(\shifter_0/reg_i_4 [11]), .X(n55074) );
  inv_x2_sg U53952 ( .A(\shifter_0/reg_i_4 [19]), .X(n55076) );
  inv_x2_sg U53953 ( .A(\shifter_0/reg_i_12 [7]), .X(n56660) );
  inv_x2_sg U53954 ( .A(\shifter_0/reg_i_12 [11]), .X(n56662) );
  inv_x2_sg U53955 ( .A(\shifter_0/reg_i_12 [19]), .X(n56664) );
  inv_x2_sg U53956 ( .A(\shifter_0/reg_i_13 [7]), .X(n56666) );
  inv_x2_sg U53957 ( .A(\shifter_0/reg_i_13 [11]), .X(n56668) );
  inv_x2_sg U53958 ( .A(\shifter_0/reg_i_13 [19]), .X(n56670) );
  inv_x2_sg U53959 ( .A(\shifter_0/reg_i_14 [15]), .X(n51212) );
  inv_x2_sg U53960 ( .A(\shifter_0/reg_w_4 [7]), .X(n55078) );
  inv_x2_sg U53961 ( .A(\shifter_0/reg_w_4 [11]), .X(n55080) );
  inv_x2_sg U53962 ( .A(\shifter_0/reg_w_4 [19]), .X(n55082) );
  inv_x2_sg U53963 ( .A(\shifter_0/reg_w_11 [2]), .X(n51218) );
  inv_x2_sg U53964 ( .A(\shifter_0/reg_w_11 [6]), .X(n51220) );
  inv_x2_sg U53965 ( .A(\shifter_0/reg_w_12 [7]), .X(n56684) );
  inv_x2_sg U53966 ( .A(\shifter_0/reg_w_12 [11]), .X(n56686) );
  inv_x2_sg U53967 ( .A(\shifter_0/reg_w_12 [19]), .X(n56688) );
  inv_x2_sg U53968 ( .A(\shifter_0/reg_w_13 [7]), .X(n56690) );
  inv_x2_sg U53969 ( .A(\shifter_0/reg_w_13 [11]), .X(n56692) );
  inv_x2_sg U53970 ( .A(\shifter_0/reg_w_13 [19]), .X(n56694) );
  inv_x2_sg U53971 ( .A(\shifter_0/reg_i_12 [15]), .X(n56698) );
  inv_x2_sg U53972 ( .A(\shifter_0/reg_i_13 [15]), .X(n56700) );
  inv_x2_sg U53973 ( .A(\shifter_0/reg_w_12 [15]), .X(n56702) );
  inv_x2_sg U53974 ( .A(\shifter_0/reg_w_13 [15]), .X(n56704) );
  inv_x2_sg U53975 ( .A(\shifter_0/reg_i_4 [14]), .X(n51146) );
  inv_x2_sg U53976 ( .A(\shifter_0/reg_w_4 [14]), .X(n51148) );
  inv_x2_sg U53977 ( .A(\shifter_0/reg_i_0 [0]), .X(n51182) );
  inv_x2_sg U53978 ( .A(\shifter_0/reg_i_0 [1]), .X(n51184) );
  inv_x2_sg U53979 ( .A(\shifter_0/reg_w_0 [0]), .X(n51186) );
  inv_x2_sg U53980 ( .A(\shifter_0/reg_w_0 [1]), .X(n51188) );
  inv_x2_sg U53981 ( .A(\shifter_0/reg_i_12 [4]), .X(n56706) );
  inv_x2_sg U53982 ( .A(\shifter_0/reg_i_12 [9]), .X(n56708) );
  inv_x2_sg U53983 ( .A(\shifter_0/reg_i_12 [13]), .X(n56710) );
  inv_x2_sg U53984 ( .A(\shifter_0/reg_i_13 [4]), .X(n56712) );
  inv_x2_sg U53985 ( .A(\shifter_0/reg_i_13 [9]), .X(n56714) );
  inv_x2_sg U53986 ( .A(\shifter_0/reg_i_13 [13]), .X(n56716) );
  inv_x2_sg U53987 ( .A(\shifter_0/reg_i_14 [12]), .X(n51256) );
  inv_x2_sg U53988 ( .A(\shifter_0/reg_w_9 [3]), .X(n56720) );
  inv_x2_sg U53989 ( .A(\shifter_0/reg_w_10 [4]), .X(n51260) );
  inv_x2_sg U53990 ( .A(\shifter_0/reg_w_11 [4]), .X(n56724) );
  inv_x2_sg U53991 ( .A(\shifter_0/reg_w_12 [4]), .X(n56726) );
  inv_x2_sg U53992 ( .A(\shifter_0/reg_w_12 [9]), .X(n56728) );
  inv_x2_sg U53993 ( .A(\shifter_0/reg_w_12 [13]), .X(n56730) );
  inv_x2_sg U53994 ( .A(\shifter_0/reg_w_13 [4]), .X(n56732) );
  inv_x2_sg U53995 ( .A(\shifter_0/reg_w_13 [9]), .X(n56734) );
  inv_x2_sg U53996 ( .A(\shifter_0/reg_w_13 [13]), .X(n56736) );
  inv_x2_sg U53997 ( .A(\shifter_0/reg_w_14 [3]), .X(n51276) );
  inv_x2_sg U53998 ( .A(n47492), .X(n47493) );
  inv_x2_sg U53999 ( .A(\shifter_0/reg_i_9 [14]), .X(n56746) );
  inv_x2_sg U54000 ( .A(\shifter_0/reg_i_10 [15]), .X(n56754) );
  inv_x2_sg U54001 ( .A(\shifter_0/reg_i_11 [6]), .X(n51292) );
  inv_x2_sg U54002 ( .A(\shifter_0/reg_i_11 [10]), .X(n51294) );
  inv_x2_sg U54003 ( .A(\shifter_0/reg_i_11 [15]), .X(n56760) );
  inv_x2_sg U54004 ( .A(\shifter_0/reg_i_14 [2]), .X(n51298) );
  inv_x2_sg U54005 ( .A(n47494), .X(n47495) );
  inv_x2_sg U54006 ( .A(\shifter_0/reg_w_9 [14]), .X(n56764) );
  inv_x2_sg U54007 ( .A(\shifter_0/reg_w_10 [15]), .X(n56768) );
  inv_x2_sg U54008 ( .A(\shifter_0/reg_w_11 [10]), .X(n51312) );
  inv_x2_sg U54009 ( .A(\shifter_0/reg_w_11 [15]), .X(n56772) );
  inv_x2_sg U54010 ( .A(\shifter_0/reg_w_14 [15]), .X(n51318) );
  inv_x2_sg U54011 ( .A(\shifter_0/reg_i_11 [19]), .X(n56774) );
  inv_x2_sg U54012 ( .A(\shifter_0/reg_w_14 [19]), .X(n51328) );
  inv_x2_sg U54013 ( .A(\shifter_0/reg_i_5 [3]), .X(n51330) );
  inv_x2_sg U54014 ( .A(\shifter_0/reg_i_5 [8]), .X(n51332) );
  inv_x2_sg U54015 ( .A(\shifter_0/reg_i_5 [12]), .X(n51334) );
  inv_x2_sg U54016 ( .A(\shifter_0/reg_w_5 [3]), .X(n51336) );
  inv_x2_sg U54017 ( .A(\shifter_0/reg_w_5 [8]), .X(n51338) );
  inv_x2_sg U54018 ( .A(\shifter_0/reg_w_5 [12]), .X(n51340) );
  inv_x2_sg U54019 ( .A(\shifter_0/reg_i_9 [3]), .X(n56790) );
  inv_x2_sg U54020 ( .A(\shifter_0/reg_i_9 [12]), .X(n56794) );
  inv_x2_sg U54021 ( .A(\shifter_0/reg_i_10 [4]), .X(n51348) );
  inv_x2_sg U54022 ( .A(\shifter_0/reg_i_10 [8]), .X(n56798) );
  inv_x2_sg U54023 ( .A(\shifter_0/reg_i_10 [13]), .X(n51352) );
  inv_x2_sg U54024 ( .A(\shifter_0/reg_i_11 [4]), .X(n56802) );
  inv_x2_sg U54025 ( .A(\shifter_0/reg_i_11 [8]), .X(n51356) );
  inv_x2_sg U54026 ( .A(\shifter_0/reg_i_11 [13]), .X(n56806) );
  inv_x2_sg U54027 ( .A(\shifter_0/reg_i_14 [3]), .X(n51360) );
  inv_x2_sg U54028 ( .A(\shifter_0/reg_i_14 [9]), .X(n51362) );
  inv_x2_sg U54029 ( .A(\shifter_0/reg_w_9 [12]), .X(n56812) );
  inv_x2_sg U54030 ( .A(\shifter_0/reg_w_10 [8]), .X(n56814) );
  inv_x2_sg U54031 ( .A(\shifter_0/reg_w_10 [13]), .X(n51370) );
  inv_x2_sg U54032 ( .A(\shifter_0/reg_w_11 [8]), .X(n51372) );
  inv_x2_sg U54033 ( .A(\shifter_0/reg_w_11 [13]), .X(n56820) );
  inv_x2_sg U54034 ( .A(\shifter_0/reg_w_14 [9]), .X(n51376) );
  inv_x2_sg U54035 ( .A(\shifter_0/reg_w_14 [12]), .X(n51378) );
  inv_x2_sg U54036 ( .A(\shifter_0/reg_i_0 [5]), .X(n51190) );
  inv_x2_sg U54037 ( .A(\shifter_0/reg_i_0 [14]), .X(n51192) );
  inv_x2_sg U54038 ( .A(\shifter_0/reg_i_0 [16]), .X(n55270) );
  inv_x2_sg U54039 ( .A(\shifter_0/reg_i_5 [7]), .X(n56824) );
  inv_x2_sg U54040 ( .A(\shifter_0/reg_i_5 [11]), .X(n56826) );
  inv_x2_sg U54041 ( .A(\shifter_0/reg_i_5 [14]), .X(n51386) );
  inv_x2_sg U54042 ( .A(\shifter_0/reg_i_12 [18]), .X(n56830) );
  inv_x2_sg U54043 ( .A(\shifter_0/reg_i_13 [18]), .X(n56832) );
  inv_x2_sg U54044 ( .A(\shifter_0/reg_i_14 [17]), .X(n51392) );
  inv_x2_sg U54045 ( .A(\shifter_0/reg_w_0 [5]), .X(n51194) );
  inv_x2_sg U54046 ( .A(\shifter_0/reg_w_0 [14]), .X(n51196) );
  inv_x2_sg U54047 ( .A(\shifter_0/reg_w_0 [16]), .X(n55282) );
  inv_x2_sg U54048 ( .A(\shifter_0/reg_w_5 [7]), .X(n56836) );
  inv_x2_sg U54049 ( .A(\shifter_0/reg_w_5 [11]), .X(n56838) );
  inv_x2_sg U54050 ( .A(\shifter_0/reg_w_5 [14]), .X(n51400) );
  inv_x2_sg U54051 ( .A(\shifter_0/reg_w_12 [17]), .X(n51402) );
  inv_x2_sg U54052 ( .A(\shifter_0/reg_w_13 [18]), .X(n56844) );
  inv_x2_sg U54053 ( .A(\shifter_0/reg_i_5 [19]), .X(n56846) );
  inv_x2_sg U54054 ( .A(\shifter_0/reg_w_5 [19]), .X(n56848) );
  inv_x2_sg U54055 ( .A(\shifter_0/reg_i_11 [18]), .X(n51410) );
  inv_x2_sg U54056 ( .A(\shifter_0/reg_i_10 [16]), .X(n51416) );
  inv_x2_sg U54057 ( .A(\shifter_0/reg_w_10 [16]), .X(n51420) );
  inv_x2_sg U54058 ( .A(\shifter_0/reg_w_14 [16]), .X(n51422) );
  inv_x2_sg U54059 ( .A(\shifter_0/reg_i_5 [16]), .X(n56864) );
  inv_x2_sg U54060 ( .A(\shifter_0/reg_w_5 [16]), .X(n56866) );
  inv_x2_sg U54061 ( .A(mask_input_ready), .X(n55070) );
  inv_x2_sg U54062 ( .A(\shifter_0/reg_i_2 [2]), .X(n55220) );
  inv_x2_sg U54063 ( .A(\shifter_0/reg_i_2 [9]), .X(n51156) );
  inv_x2_sg U54064 ( .A(\shifter_0/reg_i_2 [13]), .X(n51160) );
  inv_x2_sg U54065 ( .A(\shifter_0/reg_i_6 [14]), .X(n56874) );
  inv_x2_sg U54066 ( .A(\shifter_0/reg_w_2 [4]), .X(n51162) );
  inv_x2_sg U54067 ( .A(\shifter_0/reg_w_2 [13]), .X(n51170) );
  inv_x2_sg U54068 ( .A(\shifter_0/reg_w_6 [14]), .X(n56882) );
  inv_x2_sg U54069 ( .A(\shifter_0/reg_w_2 [9]), .X(n51166) );
  inv_x2_sg U54070 ( .A(\shifter_0/reg_i_2 [15]), .X(n51174) );
  inv_x2_sg U54071 ( .A(\shifter_0/reg_i_6 [4]), .X(n51440) );
  inv_x2_sg U54072 ( .A(\shifter_0/reg_i_6 [9]), .X(n51442) );
  inv_x2_sg U54073 ( .A(\shifter_0/reg_i_6 [13]), .X(n51444) );
  inv_x2_sg U54074 ( .A(\shifter_0/reg_w_2 [15]), .X(n51176) );
  inv_x2_sg U54075 ( .A(\shifter_0/reg_w_6 [4]), .X(n51446) );
  inv_x2_sg U54076 ( .A(\shifter_0/reg_w_6 [9]), .X(n51448) );
  inv_x2_sg U54077 ( .A(\shifter_0/reg_w_6 [13]), .X(n51450) );
  inv_x2_sg U54078 ( .A(\shifter_0/reg_i_3 [7]), .X(n56884) );
  inv_x2_sg U54079 ( .A(\shifter_0/reg_i_3 [11]), .X(n56886) );
  inv_x2_sg U54080 ( .A(\shifter_0/reg_i_3 [19]), .X(n56888) );
  inv_x2_sg U54081 ( .A(\shifter_0/reg_w_3 [7]), .X(n56890) );
  inv_x2_sg U54082 ( .A(\shifter_0/reg_w_3 [11]), .X(n56892) );
  inv_x2_sg U54083 ( .A(\shifter_0/reg_w_3 [19]), .X(n56894) );
  inv_x2_sg U54084 ( .A(\shifter_0/reg_i_3 [3]), .X(n51464) );
  inv_x2_sg U54085 ( .A(\shifter_0/reg_i_3 [8]), .X(n51466) );
  inv_x2_sg U54086 ( .A(\shifter_0/reg_i_3 [14]), .X(n51470) );
  inv_x2_sg U54087 ( .A(\shifter_0/reg_w_3 [12]), .X(n51478) );
  inv_x2_sg U54088 ( .A(\shifter_0/reg_w_3 [14]), .X(n51480) );
  inv_x2_sg U54089 ( .A(\shifter_0/reg_i_3 [18]), .X(n56912) );
  inv_x2_sg U54090 ( .A(\shifter_0/reg_w_3 [18]), .X(n56914) );
  inv_x2_sg U54091 ( .A(\shifter_0/pointer [1]), .X(n53716) );
  nor_x1_sg U54092 ( .A(n57308), .B(n26327), .X(n26325) );
  nor_x2_sg U54093 ( .A(n51067), .B(n57091), .X(n26327) );
  nor_x2_sg U54094 ( .A(n51509), .B(n57153), .X(n23076) );
  nor_x2_sg U54095 ( .A(n51497), .B(n57152), .X(n23054) );
  nor_x2_sg U54096 ( .A(n57031), .B(n22988), .X(n23032) );
  nor_x2_sg U54097 ( .A(n51515), .B(n57159), .X(n22849) );
  nor_x2_sg U54098 ( .A(n51491), .B(n57158), .X(n22827) );
  nor_x2_sg U54099 ( .A(n57015), .B(n22761), .X(n22805) );
  inv_x4_sg U54100 ( .A(n25780), .X(n67462) );
  inv_x4_sg U54101 ( .A(n25540), .X(n67470) );
  inv_x4_sg U54102 ( .A(n25328), .X(n67264) );
  inv_x4_sg U54103 ( .A(n25058), .X(n67273) );
  inv_x4_sg U54104 ( .A(n24908), .X(n67278) );
  nor_x4_sg U54105 ( .A(n35705), .B(n57779), .X(n35708) );
  nand_x2_sg U54106 ( .A(n58616), .B(n57100), .X(n57976) );
  inv_x4_sg U54107 ( .A(n58477), .X(n29332) );
  nand_x2_sg U54108 ( .A(n58479), .B(n57349), .X(n58477) );
  inv_x4_sg U54109 ( .A(n22590), .X(n67357) );
  inv_x4_sg U54110 ( .A(n22587), .X(n67360) );
  inv_x4_sg U54111 ( .A(n22584), .X(n67363) );
  inv_x4_sg U54112 ( .A(n22582), .X(n67365) );
  inv_x4_sg U54113 ( .A(n22580), .X(n67367) );
  inv_x4_sg U54114 ( .A(n22566), .X(n67142) );
  inv_x4_sg U54115 ( .A(n22564), .X(n67144) );
  inv_x4_sg U54116 ( .A(n22561), .X(n67147) );
  inv_x4_sg U54117 ( .A(n22558), .X(n67150) );
  inv_x4_sg U54118 ( .A(n22556), .X(n67152) );
  inv_x4_sg U54119 ( .A(n22554), .X(n67154) );
  inv_x4_sg U54120 ( .A(n22540), .X(n67338) );
  inv_x4_sg U54121 ( .A(n22517), .X(n67123) );
  inv_x4_sg U54122 ( .A(n22515), .X(n67125) );
  inv_x4_sg U54123 ( .A(n47759), .X(n67307) );
  inv_x2_sg U54124 ( .A(n47496), .X(n47497) );
  inv_x2_sg U54125 ( .A(n47498), .X(n47499) );
  inv_x2_sg U54126 ( .A(n47500), .X(n47501) );
  inv_x2_sg U54127 ( .A(n47502), .X(n47503) );
  inv_x4_sg U54128 ( .A(n47504), .X(n47505) );
  inv_x4_sg U54129 ( .A(n47506), .X(n47507) );
  inv_x4_sg U54130 ( .A(n47508), .X(n47509) );
  inv_x4_sg U54131 ( .A(n47510), .X(n47511) );
  inv_x4_sg U54132 ( .A(n47512), .X(n47513) );
  inv_x4_sg U54133 ( .A(n47514), .X(n47515) );
  inv_x4_sg U54134 ( .A(n47516), .X(n47517) );
  inv_x4_sg U54135 ( .A(n47518), .X(n47519) );
  nor_x8_sg U54136 ( .A(n57951), .B(n58613), .X(n31994) );
  nand_x8_sg U54137 ( .A(n57454), .B(n61910), .X(n58613) );
  inv_x4_sg U54138 ( .A(n47520), .X(n47521) );
  inv_x4_sg U54139 ( .A(n47522), .X(n47523) );
  inv_x4_sg U54140 ( .A(n47524), .X(n47525) );
  inv_x4_sg U54141 ( .A(n47526), .X(n47527) );
  inv_x4_sg U54142 ( .A(n47528), .X(n47529) );
  inv_x4_sg U54143 ( .A(n47530), .X(n47531) );
  inv_x4_sg U54144 ( .A(n47532), .X(n47533) );
  inv_x4_sg U54145 ( .A(n47534), .X(n47535) );
  inv_x4_sg U54146 ( .A(n47536), .X(n47537) );
  inv_x4_sg U54147 ( .A(n47538), .X(n47539) );
  inv_x4_sg U54148 ( .A(n47540), .X(n47541) );
  inv_x4_sg U54149 ( .A(n47542), .X(n47543) );
  inv_x4_sg U54150 ( .A(n47544), .X(n47545) );
  inv_x4_sg U54151 ( .A(n47546), .X(n47547) );
  inv_x4_sg U54152 ( .A(n47548), .X(n47549) );
  inv_x4_sg U54153 ( .A(n47550), .X(n47551) );
  inv_x4_sg U54154 ( .A(n47552), .X(n47553) );
  inv_x4_sg U54155 ( .A(n47554), .X(n47555) );
  inv_x4_sg U54156 ( .A(n47556), .X(n47557) );
  inv_x4_sg U54157 ( .A(n47558), .X(n47559) );
  inv_x4_sg U54158 ( .A(n47560), .X(n47561) );
  inv_x4_sg U54159 ( .A(n47562), .X(n47563) );
  inv_x4_sg U54160 ( .A(n47564), .X(n47565) );
  inv_x4_sg U54161 ( .A(n47566), .X(n47567) );
  inv_x4_sg U54162 ( .A(n47568), .X(n47569) );
  inv_x4_sg U54163 ( .A(n47570), .X(n47571) );
  inv_x8_sg U54164 ( .A(n57300), .X(n68572) );
  inv_x2_sg U54165 ( .A(n51543), .X(n58484) );
  inv_x2_sg U54166 ( .A(n51549), .X(n58535) );
  nor_x2_sg U54167 ( .A(n26080), .B(n68373), .X(n26079) );
  nor_x2_sg U54168 ( .A(n57069), .B(n26123), .X(n26078) );
  nand_x4_sg U54169 ( .A(n26077), .B(n67574), .X(n26060) );
  nand_x2_sg U54170 ( .A(n47485), .B(n57862), .X(n23047) );
  nand_x2_sg U54171 ( .A(n47489), .B(n57862), .X(n22952) );
  nand_x2_sg U54172 ( .A(n47487), .B(n57862), .X(n22842) );
  nand_x2_sg U54173 ( .A(n47483), .B(n57862), .X(n22820) );
  nand_x4_sg U54174 ( .A(n25844), .B(n25845), .X(n24126) );
  nand_x4_sg U54175 ( .A(n25604), .B(n25605), .X(n24086) );
  nand_x4_sg U54176 ( .A(n25484), .B(n25485), .X(n24066) );
  nand_x4_sg U54177 ( .A(n25122), .B(n25123), .X(n23996) );
  nand_x4_sg U54178 ( .A(n24882), .B(n24883), .X(n23956) );
  nor_x2_sg U54179 ( .A(n68574), .B(n23543), .X(n23541) );
  inv_x4_sg U54180 ( .A(n56993), .X(n68480) );
  nand_x2_sg U54181 ( .A(n68481), .B(n68482), .X(n32494) );
  inv_x4_sg U54182 ( .A(n57005), .X(n68481) );
  nand_x2_sg U54183 ( .A(n68485), .B(n68486), .X(n32506) );
  inv_x4_sg U54184 ( .A(n56973), .X(n68485) );
  nand_x2_sg U54185 ( .A(n68585), .B(n68586), .X(n32060) );
  inv_x4_sg U54186 ( .A(n56997), .X(n68585) );
  nand_x2_sg U54187 ( .A(n68483), .B(n68484), .X(n32500) );
  inv_x4_sg U54188 ( .A(n56999), .X(n68483) );
  nand_x2_sg U54189 ( .A(n68583), .B(n68584), .X(n32057) );
  inv_x4_sg U54190 ( .A(n57001), .X(n68583) );
  inv_x4_sg U54191 ( .A(n56981), .X(n68580) );
  nand_x2_sg U54192 ( .A(n68581), .B(n68582), .X(n32051) );
  inv_x4_sg U54193 ( .A(n57009), .X(n68581) );
  inv_x4_sg U54194 ( .A(n57047), .X(n58611) );
  inv_x4_sg U54195 ( .A(n57045), .X(n58650) );
  inv_x4_sg U54196 ( .A(state[1]), .X(n68271) );
  inv_x2_sg U54197 ( .A(\filter_0/reg_i_0 [0]), .X(n55316) );
  inv_x2_sg U54198 ( .A(\filter_0/reg_i_0 [1]), .X(n55318) );
  inv_x2_sg U54199 ( .A(\filter_0/reg_i_0 [2]), .X(n55320) );
  inv_x2_sg U54200 ( .A(\filter_0/reg_i_0 [3]), .X(n55322) );
  inv_x2_sg U54201 ( .A(\filter_0/reg_i_0 [4]), .X(n55324) );
  inv_x2_sg U54202 ( .A(\filter_0/reg_i_0 [5]), .X(n55326) );
  inv_x2_sg U54203 ( .A(\filter_0/reg_i_0 [6]), .X(n55328) );
  inv_x2_sg U54204 ( .A(\filter_0/reg_i_0 [7]), .X(n55330) );
  inv_x2_sg U54205 ( .A(\filter_0/reg_i_0 [8]), .X(n55332) );
  inv_x2_sg U54206 ( .A(\filter_0/reg_i_0 [9]), .X(n55334) );
  inv_x2_sg U54207 ( .A(\filter_0/reg_i_0 [10]), .X(n55336) );
  inv_x2_sg U54208 ( .A(\filter_0/reg_i_0 [11]), .X(n55338) );
  inv_x2_sg U54209 ( .A(\filter_0/reg_i_0 [12]), .X(n55340) );
  inv_x2_sg U54210 ( .A(\filter_0/reg_i_0 [13]), .X(n55342) );
  inv_x2_sg U54211 ( .A(\filter_0/reg_i_0 [14]), .X(n55344) );
  inv_x2_sg U54212 ( .A(\filter_0/reg_i_0 [15]), .X(n55346) );
  inv_x2_sg U54213 ( .A(\filter_0/reg_i_0 [16]), .X(n55348) );
  inv_x2_sg U54214 ( .A(\filter_0/reg_i_0 [17]), .X(n55350) );
  inv_x2_sg U54215 ( .A(\filter_0/reg_i_0 [18]), .X(n55352) );
  inv_x2_sg U54216 ( .A(\filter_0/reg_i_0 [19]), .X(n55354) );
  inv_x2_sg U54217 ( .A(\filter_0/reg_i_1 [0]), .X(n55356) );
  inv_x2_sg U54218 ( .A(\filter_0/reg_i_1 [1]), .X(n55358) );
  inv_x2_sg U54219 ( .A(\filter_0/reg_i_1 [2]), .X(n55360) );
  inv_x2_sg U54220 ( .A(\filter_0/reg_i_1 [3]), .X(n55362) );
  inv_x2_sg U54221 ( .A(\filter_0/reg_i_1 [4]), .X(n55364) );
  inv_x2_sg U54222 ( .A(\filter_0/reg_i_1 [5]), .X(n55366) );
  inv_x2_sg U54223 ( .A(\filter_0/reg_i_1 [6]), .X(n55368) );
  inv_x2_sg U54224 ( .A(\filter_0/reg_i_1 [7]), .X(n55370) );
  inv_x2_sg U54225 ( .A(\filter_0/reg_i_1 [8]), .X(n55372) );
  inv_x2_sg U54226 ( .A(\filter_0/reg_i_1 [9]), .X(n55374) );
  inv_x2_sg U54227 ( .A(\filter_0/reg_i_1 [10]), .X(n55376) );
  inv_x2_sg U54228 ( .A(\filter_0/reg_i_1 [11]), .X(n55378) );
  inv_x2_sg U54229 ( .A(\filter_0/reg_i_1 [12]), .X(n55380) );
  inv_x2_sg U54230 ( .A(\filter_0/reg_i_1 [13]), .X(n55382) );
  inv_x2_sg U54231 ( .A(\filter_0/reg_i_1 [14]), .X(n55384) );
  inv_x2_sg U54232 ( .A(\filter_0/reg_i_1 [15]), .X(n55386) );
  inv_x2_sg U54233 ( .A(\filter_0/reg_i_1 [16]), .X(n55388) );
  inv_x2_sg U54234 ( .A(\filter_0/reg_i_1 [17]), .X(n55390) );
  inv_x2_sg U54235 ( .A(\filter_0/reg_i_1 [18]), .X(n55392) );
  inv_x2_sg U54236 ( .A(\filter_0/reg_i_1 [19]), .X(n55394) );
  inv_x2_sg U54237 ( .A(\filter_0/reg_i_2 [0]), .X(n55396) );
  inv_x2_sg U54238 ( .A(\filter_0/reg_i_2 [1]), .X(n55398) );
  inv_x2_sg U54239 ( .A(\filter_0/reg_i_2 [2]), .X(n55400) );
  inv_x2_sg U54240 ( .A(\filter_0/reg_i_2 [3]), .X(n55402) );
  inv_x2_sg U54241 ( .A(\filter_0/reg_i_2 [4]), .X(n55404) );
  inv_x2_sg U54242 ( .A(\filter_0/reg_i_2 [5]), .X(n55406) );
  inv_x2_sg U54243 ( .A(\filter_0/reg_i_2 [6]), .X(n55408) );
  inv_x2_sg U54244 ( .A(\filter_0/reg_i_2 [7]), .X(n55410) );
  inv_x2_sg U54245 ( .A(\filter_0/reg_i_2 [8]), .X(n55412) );
  inv_x2_sg U54246 ( .A(\filter_0/reg_i_2 [9]), .X(n55414) );
  inv_x2_sg U54247 ( .A(\filter_0/reg_i_2 [10]), .X(n55416) );
  inv_x2_sg U54248 ( .A(\filter_0/reg_i_2 [11]), .X(n55418) );
  inv_x2_sg U54249 ( .A(\filter_0/reg_i_2 [12]), .X(n55420) );
  inv_x2_sg U54250 ( .A(\filter_0/reg_i_2 [13]), .X(n55422) );
  inv_x2_sg U54251 ( .A(\filter_0/reg_i_2 [14]), .X(n55424) );
  inv_x2_sg U54252 ( .A(\filter_0/reg_i_2 [15]), .X(n55426) );
  inv_x2_sg U54253 ( .A(\filter_0/reg_i_2 [16]), .X(n55428) );
  inv_x2_sg U54254 ( .A(\filter_0/reg_i_2 [17]), .X(n55430) );
  inv_x2_sg U54255 ( .A(\filter_0/reg_i_2 [18]), .X(n55432) );
  inv_x2_sg U54256 ( .A(\filter_0/reg_i_2 [19]), .X(n55434) );
  inv_x2_sg U54257 ( .A(\filter_0/reg_i_3 [0]), .X(n55436) );
  inv_x2_sg U54258 ( .A(\filter_0/reg_i_3 [1]), .X(n55438) );
  inv_x2_sg U54259 ( .A(\filter_0/reg_i_3 [2]), .X(n55440) );
  inv_x2_sg U54260 ( .A(\filter_0/reg_i_3 [3]), .X(n55442) );
  inv_x2_sg U54261 ( .A(\filter_0/reg_i_3 [4]), .X(n55444) );
  inv_x2_sg U54262 ( .A(\filter_0/reg_i_3 [5]), .X(n55446) );
  inv_x2_sg U54263 ( .A(\filter_0/reg_i_3 [6]), .X(n55448) );
  inv_x2_sg U54264 ( .A(\filter_0/reg_i_3 [7]), .X(n55450) );
  inv_x2_sg U54265 ( .A(\filter_0/reg_i_3 [8]), .X(n55452) );
  inv_x2_sg U54266 ( .A(\filter_0/reg_i_3 [9]), .X(n55454) );
  inv_x2_sg U54267 ( .A(\filter_0/reg_i_3 [10]), .X(n55456) );
  inv_x2_sg U54268 ( .A(\filter_0/reg_i_3 [11]), .X(n55458) );
  inv_x2_sg U54269 ( .A(\filter_0/reg_i_3 [12]), .X(n55460) );
  inv_x2_sg U54270 ( .A(\filter_0/reg_i_3 [13]), .X(n55462) );
  inv_x2_sg U54271 ( .A(\filter_0/reg_i_3 [14]), .X(n55464) );
  inv_x2_sg U54272 ( .A(\filter_0/reg_i_3 [15]), .X(n55466) );
  inv_x2_sg U54273 ( .A(\filter_0/reg_i_3 [16]), .X(n55468) );
  inv_x2_sg U54274 ( .A(\filter_0/reg_i_3 [17]), .X(n55470) );
  inv_x2_sg U54275 ( .A(\filter_0/reg_i_3 [18]), .X(n55472) );
  inv_x2_sg U54276 ( .A(\filter_0/reg_i_3 [19]), .X(n55474) );
  inv_x2_sg U54277 ( .A(\filter_0/reg_i_4 [0]), .X(n55476) );
  inv_x2_sg U54278 ( .A(\filter_0/reg_i_4 [1]), .X(n55478) );
  inv_x2_sg U54279 ( .A(\filter_0/reg_i_4 [2]), .X(n55480) );
  inv_x2_sg U54280 ( .A(\filter_0/reg_i_4 [3]), .X(n55482) );
  inv_x2_sg U54281 ( .A(\filter_0/reg_i_4 [4]), .X(n55484) );
  inv_x2_sg U54282 ( .A(\filter_0/reg_i_4 [5]), .X(n55486) );
  inv_x2_sg U54283 ( .A(\filter_0/reg_i_4 [6]), .X(n55488) );
  inv_x2_sg U54284 ( .A(\filter_0/reg_i_4 [7]), .X(n55490) );
  inv_x2_sg U54285 ( .A(\filter_0/reg_i_4 [8]), .X(n55492) );
  inv_x2_sg U54286 ( .A(\filter_0/reg_i_4 [9]), .X(n55494) );
  inv_x2_sg U54287 ( .A(\filter_0/reg_i_4 [10]), .X(n55496) );
  inv_x2_sg U54288 ( .A(\filter_0/reg_i_4 [11]), .X(n55498) );
  inv_x2_sg U54289 ( .A(\filter_0/reg_i_4 [12]), .X(n55500) );
  inv_x2_sg U54290 ( .A(\filter_0/reg_i_4 [13]), .X(n55502) );
  inv_x2_sg U54291 ( .A(\filter_0/reg_i_4 [14]), .X(n55504) );
  inv_x2_sg U54292 ( .A(\filter_0/reg_i_4 [15]), .X(n55506) );
  inv_x2_sg U54293 ( .A(\filter_0/reg_i_4 [16]), .X(n55508) );
  inv_x2_sg U54294 ( .A(\filter_0/reg_i_4 [17]), .X(n55510) );
  inv_x2_sg U54295 ( .A(\filter_0/reg_i_4 [18]), .X(n55512) );
  inv_x2_sg U54296 ( .A(\filter_0/reg_i_4 [19]), .X(n55514) );
  inv_x2_sg U54297 ( .A(\filter_0/reg_i_5 [0]), .X(n55516) );
  inv_x2_sg U54298 ( .A(\filter_0/reg_i_5 [1]), .X(n55518) );
  inv_x2_sg U54299 ( .A(\filter_0/reg_i_5 [2]), .X(n55520) );
  inv_x2_sg U54300 ( .A(\filter_0/reg_i_5 [3]), .X(n55522) );
  inv_x2_sg U54301 ( .A(\filter_0/reg_i_5 [4]), .X(n55524) );
  inv_x2_sg U54302 ( .A(\filter_0/reg_i_5 [5]), .X(n55526) );
  inv_x2_sg U54303 ( .A(\filter_0/reg_i_5 [6]), .X(n55528) );
  inv_x2_sg U54304 ( .A(\filter_0/reg_i_5 [7]), .X(n55530) );
  inv_x2_sg U54305 ( .A(\filter_0/reg_i_5 [8]), .X(n55532) );
  inv_x2_sg U54306 ( .A(\filter_0/reg_i_5 [9]), .X(n55534) );
  inv_x2_sg U54307 ( .A(\filter_0/reg_i_5 [10]), .X(n55536) );
  inv_x2_sg U54308 ( .A(\filter_0/reg_i_5 [11]), .X(n55538) );
  inv_x2_sg U54309 ( .A(\filter_0/reg_i_5 [12]), .X(n55540) );
  inv_x2_sg U54310 ( .A(\filter_0/reg_i_5 [13]), .X(n55542) );
  inv_x2_sg U54311 ( .A(\filter_0/reg_i_5 [14]), .X(n55544) );
  inv_x2_sg U54312 ( .A(\filter_0/reg_i_5 [15]), .X(n55546) );
  inv_x2_sg U54313 ( .A(\filter_0/reg_i_5 [16]), .X(n55548) );
  inv_x2_sg U54314 ( .A(\filter_0/reg_i_5 [17]), .X(n55550) );
  inv_x2_sg U54315 ( .A(\filter_0/reg_i_5 [18]), .X(n55552) );
  inv_x2_sg U54316 ( .A(\filter_0/reg_i_5 [19]), .X(n55554) );
  inv_x2_sg U54317 ( .A(\filter_0/reg_i_6 [0]), .X(n55556) );
  inv_x2_sg U54318 ( .A(\filter_0/reg_i_6 [1]), .X(n55558) );
  inv_x2_sg U54319 ( .A(\filter_0/reg_i_6 [2]), .X(n55560) );
  inv_x2_sg U54320 ( .A(\filter_0/reg_i_6 [3]), .X(n55562) );
  inv_x2_sg U54321 ( .A(\filter_0/reg_i_6 [4]), .X(n55564) );
  inv_x2_sg U54322 ( .A(\filter_0/reg_i_6 [5]), .X(n55566) );
  inv_x2_sg U54323 ( .A(\filter_0/reg_i_6 [6]), .X(n55568) );
  inv_x2_sg U54324 ( .A(\filter_0/reg_i_6 [7]), .X(n55570) );
  inv_x2_sg U54325 ( .A(\filter_0/reg_i_6 [8]), .X(n55572) );
  inv_x2_sg U54326 ( .A(\filter_0/reg_i_6 [9]), .X(n55574) );
  inv_x2_sg U54327 ( .A(\filter_0/reg_i_6 [10]), .X(n55576) );
  inv_x2_sg U54328 ( .A(\filter_0/reg_i_6 [11]), .X(n55578) );
  inv_x2_sg U54329 ( .A(\filter_0/reg_i_6 [12]), .X(n55580) );
  inv_x2_sg U54330 ( .A(\filter_0/reg_i_6 [13]), .X(n55582) );
  inv_x2_sg U54331 ( .A(\filter_0/reg_i_6 [14]), .X(n55584) );
  inv_x2_sg U54332 ( .A(\filter_0/reg_i_6 [15]), .X(n55586) );
  inv_x2_sg U54333 ( .A(\filter_0/reg_i_6 [16]), .X(n55588) );
  inv_x2_sg U54334 ( .A(\filter_0/reg_i_6 [17]), .X(n55590) );
  inv_x2_sg U54335 ( .A(\filter_0/reg_i_6 [18]), .X(n55592) );
  inv_x2_sg U54336 ( .A(\filter_0/reg_i_6 [19]), .X(n55594) );
  inv_x2_sg U54337 ( .A(\filter_0/reg_i_7 [0]), .X(n55596) );
  inv_x2_sg U54338 ( .A(\filter_0/reg_i_7 [1]), .X(n55598) );
  inv_x2_sg U54339 ( .A(\filter_0/reg_i_7 [2]), .X(n55600) );
  inv_x2_sg U54340 ( .A(\filter_0/reg_i_7 [3]), .X(n55602) );
  inv_x2_sg U54341 ( .A(\filter_0/reg_i_7 [4]), .X(n55604) );
  inv_x2_sg U54342 ( .A(\filter_0/reg_i_7 [5]), .X(n55606) );
  inv_x2_sg U54343 ( .A(\filter_0/reg_i_7 [6]), .X(n55608) );
  inv_x2_sg U54344 ( .A(\filter_0/reg_i_7 [7]), .X(n55610) );
  inv_x2_sg U54345 ( .A(\filter_0/reg_i_7 [8]), .X(n55612) );
  inv_x2_sg U54346 ( .A(\filter_0/reg_i_7 [9]), .X(n55614) );
  inv_x2_sg U54347 ( .A(\filter_0/reg_i_7 [10]), .X(n55616) );
  inv_x2_sg U54348 ( .A(\filter_0/reg_i_7 [11]), .X(n55618) );
  inv_x2_sg U54349 ( .A(\filter_0/reg_i_7 [12]), .X(n55620) );
  inv_x2_sg U54350 ( .A(\filter_0/reg_i_7 [13]), .X(n55622) );
  inv_x2_sg U54351 ( .A(\filter_0/reg_i_7 [14]), .X(n55624) );
  inv_x2_sg U54352 ( .A(\filter_0/reg_i_7 [15]), .X(n55626) );
  inv_x2_sg U54353 ( .A(\filter_0/reg_i_7 [16]), .X(n55628) );
  inv_x2_sg U54354 ( .A(\filter_0/reg_i_7 [17]), .X(n55630) );
  inv_x2_sg U54355 ( .A(\filter_0/reg_i_7 [18]), .X(n55632) );
  inv_x2_sg U54356 ( .A(\filter_0/reg_i_7 [19]), .X(n55634) );
  inv_x2_sg U54357 ( .A(\filter_0/reg_i_8 [0]), .X(n55636) );
  inv_x2_sg U54358 ( .A(\filter_0/reg_i_8 [1]), .X(n55638) );
  inv_x2_sg U54359 ( .A(\filter_0/reg_i_8 [2]), .X(n55640) );
  inv_x2_sg U54360 ( .A(\filter_0/reg_i_8 [3]), .X(n55642) );
  inv_x2_sg U54361 ( .A(\filter_0/reg_i_8 [4]), .X(n55644) );
  inv_x2_sg U54362 ( .A(\filter_0/reg_i_8 [5]), .X(n55646) );
  inv_x2_sg U54363 ( .A(\filter_0/reg_i_8 [6]), .X(n55648) );
  inv_x2_sg U54364 ( .A(\filter_0/reg_i_8 [7]), .X(n55650) );
  inv_x2_sg U54365 ( .A(\filter_0/reg_i_8 [8]), .X(n55652) );
  inv_x2_sg U54366 ( .A(\filter_0/reg_i_8 [9]), .X(n55654) );
  inv_x2_sg U54367 ( .A(\filter_0/reg_i_8 [10]), .X(n55656) );
  inv_x2_sg U54368 ( .A(\filter_0/reg_i_8 [11]), .X(n55658) );
  inv_x2_sg U54369 ( .A(\filter_0/reg_i_8 [12]), .X(n55660) );
  inv_x2_sg U54370 ( .A(\filter_0/reg_i_8 [13]), .X(n55662) );
  inv_x2_sg U54371 ( .A(\filter_0/reg_i_8 [14]), .X(n55664) );
  inv_x2_sg U54372 ( .A(\filter_0/reg_i_8 [15]), .X(n55666) );
  inv_x2_sg U54373 ( .A(\filter_0/reg_i_8 [16]), .X(n55668) );
  inv_x2_sg U54374 ( .A(\filter_0/reg_i_8 [17]), .X(n55670) );
  inv_x2_sg U54375 ( .A(\filter_0/reg_i_8 [18]), .X(n55672) );
  inv_x2_sg U54376 ( .A(\filter_0/reg_i_8 [19]), .X(n55674) );
  inv_x2_sg U54377 ( .A(\filter_0/reg_i_9 [0]), .X(n55676) );
  inv_x2_sg U54378 ( .A(\filter_0/reg_i_9 [1]), .X(n55678) );
  inv_x2_sg U54379 ( .A(\filter_0/reg_i_9 [2]), .X(n55680) );
  inv_x2_sg U54380 ( .A(\filter_0/reg_i_9 [3]), .X(n55682) );
  inv_x2_sg U54381 ( .A(\filter_0/reg_i_9 [4]), .X(n55684) );
  inv_x2_sg U54382 ( .A(\filter_0/reg_i_9 [5]), .X(n55686) );
  inv_x2_sg U54383 ( .A(\filter_0/reg_i_9 [6]), .X(n55688) );
  inv_x2_sg U54384 ( .A(\filter_0/reg_i_9 [7]), .X(n55690) );
  inv_x2_sg U54385 ( .A(\filter_0/reg_i_9 [8]), .X(n55692) );
  inv_x2_sg U54386 ( .A(\filter_0/reg_i_9 [9]), .X(n55694) );
  inv_x2_sg U54387 ( .A(\filter_0/reg_i_9 [10]), .X(n55696) );
  inv_x2_sg U54388 ( .A(\filter_0/reg_i_9 [11]), .X(n55698) );
  inv_x2_sg U54389 ( .A(\filter_0/reg_i_9 [12]), .X(n55700) );
  inv_x2_sg U54390 ( .A(\filter_0/reg_i_9 [13]), .X(n55702) );
  inv_x2_sg U54391 ( .A(\filter_0/reg_i_9 [14]), .X(n55704) );
  inv_x2_sg U54392 ( .A(\filter_0/reg_i_9 [15]), .X(n55706) );
  inv_x2_sg U54393 ( .A(\filter_0/reg_i_9 [16]), .X(n55708) );
  inv_x2_sg U54394 ( .A(\filter_0/reg_i_9 [17]), .X(n55710) );
  inv_x2_sg U54395 ( .A(\filter_0/reg_i_9 [18]), .X(n55712) );
  inv_x2_sg U54396 ( .A(\filter_0/reg_i_9 [19]), .X(n55714) );
  inv_x2_sg U54397 ( .A(\filter_0/reg_i_10 [0]), .X(n55716) );
  inv_x2_sg U54398 ( .A(\filter_0/reg_i_10 [1]), .X(n55718) );
  inv_x2_sg U54399 ( .A(\filter_0/reg_i_10 [2]), .X(n55720) );
  inv_x2_sg U54400 ( .A(\filter_0/reg_i_10 [3]), .X(n55722) );
  inv_x2_sg U54401 ( .A(\filter_0/reg_i_10 [4]), .X(n55724) );
  inv_x2_sg U54402 ( .A(\filter_0/reg_i_10 [5]), .X(n55726) );
  inv_x2_sg U54403 ( .A(\filter_0/reg_i_10 [6]), .X(n55728) );
  inv_x2_sg U54404 ( .A(\filter_0/reg_i_10 [7]), .X(n55730) );
  inv_x2_sg U54405 ( .A(\filter_0/reg_i_10 [8]), .X(n55732) );
  inv_x2_sg U54406 ( .A(\filter_0/reg_i_10 [9]), .X(n55734) );
  inv_x2_sg U54407 ( .A(\filter_0/reg_i_10 [10]), .X(n55736) );
  inv_x2_sg U54408 ( .A(\filter_0/reg_i_10 [11]), .X(n55738) );
  inv_x2_sg U54409 ( .A(\filter_0/reg_i_10 [12]), .X(n55740) );
  inv_x2_sg U54410 ( .A(\filter_0/reg_i_10 [13]), .X(n55742) );
  inv_x2_sg U54411 ( .A(\filter_0/reg_i_10 [14]), .X(n55744) );
  inv_x2_sg U54412 ( .A(\filter_0/reg_i_10 [15]), .X(n55746) );
  inv_x2_sg U54413 ( .A(\filter_0/reg_i_10 [16]), .X(n55748) );
  inv_x2_sg U54414 ( .A(\filter_0/reg_i_10 [17]), .X(n55750) );
  inv_x2_sg U54415 ( .A(\filter_0/reg_i_10 [18]), .X(n55752) );
  inv_x2_sg U54416 ( .A(\filter_0/reg_i_10 [19]), .X(n55754) );
  inv_x2_sg U54417 ( .A(\filter_0/reg_i_11 [0]), .X(n55756) );
  inv_x2_sg U54418 ( .A(\filter_0/reg_i_11 [1]), .X(n55758) );
  inv_x2_sg U54419 ( .A(\filter_0/reg_i_11 [2]), .X(n55760) );
  inv_x2_sg U54420 ( .A(\filter_0/reg_i_11 [3]), .X(n55762) );
  inv_x2_sg U54421 ( .A(\filter_0/reg_i_11 [4]), .X(n55764) );
  inv_x2_sg U54422 ( .A(\filter_0/reg_i_11 [5]), .X(n55766) );
  inv_x2_sg U54423 ( .A(\filter_0/reg_i_11 [6]), .X(n55768) );
  inv_x2_sg U54424 ( .A(\filter_0/reg_i_11 [7]), .X(n55770) );
  inv_x2_sg U54425 ( .A(\filter_0/reg_i_11 [8]), .X(n55772) );
  inv_x2_sg U54426 ( .A(\filter_0/reg_i_11 [9]), .X(n55774) );
  inv_x2_sg U54427 ( .A(\filter_0/reg_i_11 [10]), .X(n55776) );
  inv_x2_sg U54428 ( .A(\filter_0/reg_i_11 [11]), .X(n55778) );
  inv_x2_sg U54429 ( .A(\filter_0/reg_i_11 [12]), .X(n55780) );
  inv_x2_sg U54430 ( .A(\filter_0/reg_i_11 [14]), .X(n55784) );
  inv_x2_sg U54431 ( .A(\filter_0/reg_i_11 [15]), .X(n55786) );
  inv_x2_sg U54432 ( .A(\filter_0/reg_i_11 [16]), .X(n55788) );
  inv_x2_sg U54433 ( .A(\filter_0/reg_i_11 [17]), .X(n55790) );
  inv_x2_sg U54434 ( .A(\filter_0/reg_i_11 [18]), .X(n55792) );
  inv_x2_sg U54435 ( .A(\filter_0/reg_i_11 [19]), .X(n55794) );
  inv_x2_sg U54436 ( .A(\filter_0/reg_i_12 [0]), .X(n55796) );
  inv_x2_sg U54437 ( .A(\filter_0/reg_i_12 [1]), .X(n55798) );
  inv_x2_sg U54438 ( .A(\filter_0/reg_i_12 [2]), .X(n55800) );
  inv_x2_sg U54439 ( .A(\filter_0/reg_i_12 [3]), .X(n55802) );
  inv_x2_sg U54440 ( .A(\filter_0/reg_i_12 [4]), .X(n55804) );
  inv_x2_sg U54441 ( .A(\filter_0/reg_i_12 [5]), .X(n55806) );
  inv_x2_sg U54442 ( .A(\filter_0/reg_i_12 [6]), .X(n55808) );
  inv_x2_sg U54443 ( .A(\filter_0/reg_i_12 [7]), .X(n55810) );
  inv_x2_sg U54444 ( .A(\filter_0/reg_i_12 [8]), .X(n55812) );
  inv_x2_sg U54445 ( .A(\filter_0/reg_i_12 [9]), .X(n55814) );
  inv_x2_sg U54446 ( .A(\filter_0/reg_i_12 [10]), .X(n55816) );
  inv_x2_sg U54447 ( .A(\filter_0/reg_i_12 [11]), .X(n55818) );
  inv_x2_sg U54448 ( .A(\filter_0/reg_i_12 [12]), .X(n55820) );
  inv_x2_sg U54449 ( .A(\filter_0/reg_i_12 [13]), .X(n55822) );
  inv_x2_sg U54450 ( .A(\filter_0/reg_i_12 [14]), .X(n55824) );
  inv_x2_sg U54451 ( .A(\filter_0/reg_i_12 [15]), .X(n55826) );
  inv_x2_sg U54452 ( .A(\filter_0/reg_i_12 [16]), .X(n55828) );
  inv_x2_sg U54453 ( .A(\filter_0/reg_i_12 [17]), .X(n55830) );
  inv_x2_sg U54454 ( .A(\filter_0/reg_i_12 [18]), .X(n55832) );
  inv_x2_sg U54455 ( .A(\filter_0/reg_i_12 [19]), .X(n55834) );
  inv_x2_sg U54456 ( .A(\filter_0/reg_i_13 [0]), .X(n55836) );
  inv_x2_sg U54457 ( .A(\filter_0/reg_i_13 [1]), .X(n55838) );
  inv_x2_sg U54458 ( .A(\filter_0/reg_i_13 [2]), .X(n55840) );
  inv_x2_sg U54459 ( .A(\filter_0/reg_i_13 [3]), .X(n55842) );
  inv_x2_sg U54460 ( .A(\filter_0/reg_i_13 [4]), .X(n55844) );
  inv_x2_sg U54461 ( .A(\filter_0/reg_i_13 [5]), .X(n55846) );
  inv_x2_sg U54462 ( .A(\filter_0/reg_i_13 [6]), .X(n55848) );
  inv_x2_sg U54463 ( .A(\filter_0/reg_i_13 [7]), .X(n55850) );
  inv_x2_sg U54464 ( .A(\filter_0/reg_i_13 [8]), .X(n55852) );
  inv_x2_sg U54465 ( .A(\filter_0/reg_i_13 [9]), .X(n55854) );
  inv_x2_sg U54466 ( .A(\filter_0/reg_i_13 [10]), .X(n55856) );
  inv_x2_sg U54467 ( .A(\filter_0/reg_i_13 [11]), .X(n55858) );
  inv_x2_sg U54468 ( .A(\filter_0/reg_i_13 [12]), .X(n55860) );
  inv_x2_sg U54469 ( .A(\filter_0/reg_i_13 [13]), .X(n55862) );
  inv_x2_sg U54470 ( .A(\filter_0/reg_i_13 [14]), .X(n55864) );
  inv_x2_sg U54471 ( .A(\filter_0/reg_i_13 [15]), .X(n55866) );
  inv_x2_sg U54472 ( .A(\filter_0/reg_i_13 [16]), .X(n55868) );
  inv_x2_sg U54473 ( .A(\filter_0/reg_i_13 [17]), .X(n55870) );
  inv_x2_sg U54474 ( .A(\filter_0/reg_i_13 [18]), .X(n55872) );
  inv_x2_sg U54475 ( .A(\filter_0/reg_i_13 [19]), .X(n55874) );
  inv_x2_sg U54476 ( .A(\filter_0/reg_i_14 [0]), .X(n55876) );
  inv_x2_sg U54477 ( .A(\filter_0/reg_i_14 [1]), .X(n55878) );
  inv_x2_sg U54478 ( .A(\filter_0/reg_i_14 [2]), .X(n55880) );
  inv_x2_sg U54479 ( .A(\filter_0/reg_i_14 [3]), .X(n55882) );
  inv_x2_sg U54480 ( .A(\filter_0/reg_i_14 [4]), .X(n55884) );
  inv_x2_sg U54481 ( .A(\filter_0/reg_i_14 [5]), .X(n55886) );
  inv_x2_sg U54482 ( .A(\filter_0/reg_i_14 [6]), .X(n55888) );
  inv_x2_sg U54483 ( .A(\filter_0/reg_i_14 [7]), .X(n55890) );
  inv_x2_sg U54484 ( .A(\filter_0/reg_i_14 [8]), .X(n55892) );
  inv_x2_sg U54485 ( .A(\filter_0/reg_i_14 [9]), .X(n55894) );
  inv_x2_sg U54486 ( .A(\filter_0/reg_i_14 [10]), .X(n55896) );
  inv_x2_sg U54487 ( .A(\filter_0/reg_i_14 [11]), .X(n55898) );
  inv_x2_sg U54488 ( .A(\filter_0/reg_i_14 [12]), .X(n55900) );
  inv_x2_sg U54489 ( .A(\filter_0/reg_i_14 [13]), .X(n55902) );
  inv_x2_sg U54490 ( .A(\filter_0/reg_i_14 [14]), .X(n55904) );
  inv_x2_sg U54491 ( .A(\filter_0/reg_i_14 [15]), .X(n55906) );
  inv_x2_sg U54492 ( .A(\filter_0/reg_i_14 [16]), .X(n55908) );
  inv_x2_sg U54493 ( .A(\filter_0/reg_i_14 [17]), .X(n55910) );
  inv_x2_sg U54494 ( .A(\filter_0/reg_i_14 [18]), .X(n55912) );
  inv_x2_sg U54495 ( .A(\filter_0/reg_i_14 [19]), .X(n55914) );
  inv_x2_sg U54496 ( .A(\filter_0/reg_i_15 [0]), .X(n55916) );
  inv_x2_sg U54497 ( .A(\filter_0/reg_i_15 [1]), .X(n55918) );
  inv_x2_sg U54498 ( .A(\filter_0/reg_i_15 [2]), .X(n55920) );
  inv_x2_sg U54499 ( .A(\filter_0/reg_i_15 [3]), .X(n55922) );
  inv_x2_sg U54500 ( .A(\filter_0/reg_i_15 [4]), .X(n55924) );
  inv_x2_sg U54501 ( .A(\filter_0/reg_i_15 [5]), .X(n55926) );
  inv_x2_sg U54502 ( .A(\filter_0/reg_i_15 [6]), .X(n55928) );
  inv_x2_sg U54503 ( .A(\filter_0/reg_i_15 [7]), .X(n55930) );
  inv_x2_sg U54504 ( .A(\filter_0/reg_i_15 [8]), .X(n55932) );
  inv_x2_sg U54505 ( .A(\filter_0/reg_i_15 [9]), .X(n55934) );
  inv_x2_sg U54506 ( .A(\filter_0/reg_i_15 [10]), .X(n55936) );
  inv_x2_sg U54507 ( .A(\filter_0/reg_i_15 [11]), .X(n55938) );
  inv_x2_sg U54508 ( .A(\filter_0/reg_i_15 [12]), .X(n55940) );
  inv_x2_sg U54509 ( .A(\filter_0/reg_i_15 [13]), .X(n55942) );
  inv_x2_sg U54510 ( .A(\filter_0/reg_i_15 [14]), .X(n55944) );
  inv_x2_sg U54511 ( .A(\filter_0/reg_i_15 [15]), .X(n55946) );
  inv_x2_sg U54512 ( .A(\filter_0/reg_i_15 [16]), .X(n55948) );
  inv_x2_sg U54513 ( .A(\filter_0/reg_i_15 [17]), .X(n55950) );
  inv_x2_sg U54514 ( .A(\filter_0/reg_i_15 [18]), .X(n55952) );
  inv_x2_sg U54515 ( .A(\filter_0/reg_i_15 [19]), .X(n55954) );
  inv_x2_sg U54516 ( .A(\filter_0/reg_w_0 [0]), .X(n55956) );
  inv_x2_sg U54517 ( .A(\filter_0/reg_w_0 [1]), .X(n55958) );
  inv_x2_sg U54518 ( .A(\filter_0/reg_w_0 [2]), .X(n55960) );
  inv_x2_sg U54519 ( .A(\filter_0/reg_w_0 [3]), .X(n55962) );
  inv_x2_sg U54520 ( .A(\filter_0/reg_w_0 [4]), .X(n55964) );
  inv_x2_sg U54521 ( .A(\filter_0/reg_w_0 [5]), .X(n55966) );
  inv_x2_sg U54522 ( .A(\filter_0/reg_w_0 [6]), .X(n55968) );
  inv_x2_sg U54523 ( .A(\filter_0/reg_w_0 [7]), .X(n55970) );
  inv_x2_sg U54524 ( .A(\filter_0/reg_w_0 [8]), .X(n55972) );
  inv_x2_sg U54525 ( .A(\filter_0/reg_w_0 [9]), .X(n55974) );
  inv_x2_sg U54526 ( .A(\filter_0/reg_w_0 [10]), .X(n55976) );
  inv_x2_sg U54527 ( .A(\filter_0/reg_w_0 [11]), .X(n55978) );
  inv_x2_sg U54528 ( .A(\filter_0/reg_w_0 [12]), .X(n55980) );
  inv_x2_sg U54529 ( .A(\filter_0/reg_w_0 [13]), .X(n55982) );
  inv_x2_sg U54530 ( .A(\filter_0/reg_w_0 [14]), .X(n55984) );
  inv_x2_sg U54531 ( .A(\filter_0/reg_w_0 [15]), .X(n55986) );
  inv_x2_sg U54532 ( .A(\filter_0/reg_w_0 [16]), .X(n55988) );
  inv_x2_sg U54533 ( .A(\filter_0/reg_w_0 [17]), .X(n55990) );
  inv_x2_sg U54534 ( .A(\filter_0/reg_w_0 [18]), .X(n55992) );
  inv_x2_sg U54535 ( .A(\filter_0/reg_w_0 [19]), .X(n55994) );
  inv_x2_sg U54536 ( .A(\filter_0/reg_w_1 [0]), .X(n55996) );
  inv_x2_sg U54537 ( .A(\filter_0/reg_w_1 [1]), .X(n55998) );
  inv_x2_sg U54538 ( .A(\filter_0/reg_w_1 [2]), .X(n56000) );
  inv_x2_sg U54539 ( .A(\filter_0/reg_w_1 [3]), .X(n56002) );
  inv_x2_sg U54540 ( .A(\filter_0/reg_w_1 [4]), .X(n56004) );
  inv_x2_sg U54541 ( .A(\filter_0/reg_w_1 [5]), .X(n56006) );
  inv_x2_sg U54542 ( .A(\filter_0/reg_w_1 [6]), .X(n56008) );
  inv_x2_sg U54543 ( .A(\filter_0/reg_w_1 [7]), .X(n56010) );
  inv_x2_sg U54544 ( .A(\filter_0/reg_w_1 [8]), .X(n56012) );
  inv_x2_sg U54545 ( .A(\filter_0/reg_w_1 [9]), .X(n56014) );
  inv_x2_sg U54546 ( .A(\filter_0/reg_w_1 [10]), .X(n56016) );
  inv_x2_sg U54547 ( .A(\filter_0/reg_w_1 [11]), .X(n56018) );
  inv_x2_sg U54548 ( .A(\filter_0/reg_w_1 [12]), .X(n56020) );
  inv_x2_sg U54549 ( .A(\filter_0/reg_w_1 [13]), .X(n56022) );
  inv_x2_sg U54550 ( .A(\filter_0/reg_w_1 [14]), .X(n56024) );
  inv_x2_sg U54551 ( .A(\filter_0/reg_w_1 [15]), .X(n56026) );
  inv_x2_sg U54552 ( .A(\filter_0/reg_w_1 [16]), .X(n56028) );
  inv_x2_sg U54553 ( .A(\filter_0/reg_w_1 [17]), .X(n56030) );
  inv_x2_sg U54554 ( .A(\filter_0/reg_w_1 [18]), .X(n56032) );
  inv_x2_sg U54555 ( .A(\filter_0/reg_w_1 [19]), .X(n56034) );
  inv_x2_sg U54556 ( .A(\filter_0/reg_w_2 [0]), .X(n56036) );
  inv_x2_sg U54557 ( .A(\filter_0/reg_w_2 [1]), .X(n56038) );
  inv_x2_sg U54558 ( .A(\filter_0/reg_w_2 [2]), .X(n56040) );
  inv_x2_sg U54559 ( .A(\filter_0/reg_w_2 [3]), .X(n56042) );
  inv_x2_sg U54560 ( .A(\filter_0/reg_w_2 [4]), .X(n56044) );
  inv_x2_sg U54561 ( .A(\filter_0/reg_w_2 [5]), .X(n56046) );
  inv_x2_sg U54562 ( .A(\filter_0/reg_w_2 [6]), .X(n56048) );
  inv_x2_sg U54563 ( .A(\filter_0/reg_w_2 [7]), .X(n56050) );
  inv_x2_sg U54564 ( .A(\filter_0/reg_w_2 [8]), .X(n56052) );
  inv_x2_sg U54565 ( .A(\filter_0/reg_w_2 [9]), .X(n56054) );
  inv_x2_sg U54566 ( .A(\filter_0/reg_w_2 [10]), .X(n56056) );
  inv_x2_sg U54567 ( .A(\filter_0/reg_w_2 [11]), .X(n56058) );
  inv_x2_sg U54568 ( .A(\filter_0/reg_w_2 [12]), .X(n56060) );
  inv_x2_sg U54569 ( .A(\filter_0/reg_w_2 [13]), .X(n56062) );
  inv_x2_sg U54570 ( .A(\filter_0/reg_w_2 [14]), .X(n56064) );
  inv_x2_sg U54571 ( .A(\filter_0/reg_w_2 [15]), .X(n56066) );
  inv_x2_sg U54572 ( .A(\filter_0/reg_w_2 [16]), .X(n56068) );
  inv_x2_sg U54573 ( .A(\filter_0/reg_w_2 [17]), .X(n56070) );
  inv_x2_sg U54574 ( .A(\filter_0/reg_w_2 [18]), .X(n56072) );
  inv_x2_sg U54575 ( .A(\filter_0/reg_w_2 [19]), .X(n56074) );
  inv_x2_sg U54576 ( .A(\filter_0/reg_w_3 [0]), .X(n56076) );
  inv_x2_sg U54577 ( .A(\filter_0/reg_w_3 [1]), .X(n56078) );
  inv_x2_sg U54578 ( .A(\filter_0/reg_w_3 [2]), .X(n56080) );
  inv_x2_sg U54579 ( .A(\filter_0/reg_w_3 [3]), .X(n56082) );
  inv_x2_sg U54580 ( .A(\filter_0/reg_w_3 [4]), .X(n56084) );
  inv_x2_sg U54581 ( .A(\filter_0/reg_w_3 [5]), .X(n56086) );
  inv_x2_sg U54582 ( .A(\filter_0/reg_w_3 [6]), .X(n56088) );
  inv_x2_sg U54583 ( .A(\filter_0/reg_w_3 [7]), .X(n56090) );
  inv_x2_sg U54584 ( .A(\filter_0/reg_w_3 [8]), .X(n56092) );
  inv_x2_sg U54585 ( .A(\filter_0/reg_w_3 [9]), .X(n56094) );
  inv_x2_sg U54586 ( .A(\filter_0/reg_w_3 [10]), .X(n56096) );
  inv_x2_sg U54587 ( .A(\filter_0/reg_w_3 [11]), .X(n56098) );
  inv_x2_sg U54588 ( .A(\filter_0/reg_w_3 [12]), .X(n56100) );
  inv_x2_sg U54589 ( .A(\filter_0/reg_w_3 [13]), .X(n56102) );
  inv_x2_sg U54590 ( .A(\filter_0/reg_w_3 [14]), .X(n56104) );
  inv_x2_sg U54591 ( .A(\filter_0/reg_w_3 [15]), .X(n56106) );
  inv_x2_sg U54592 ( .A(\filter_0/reg_w_3 [16]), .X(n56108) );
  inv_x2_sg U54593 ( .A(\filter_0/reg_w_3 [17]), .X(n56110) );
  inv_x2_sg U54594 ( .A(\filter_0/reg_w_3 [18]), .X(n56112) );
  inv_x2_sg U54595 ( .A(\filter_0/reg_w_3 [19]), .X(n56114) );
  inv_x2_sg U54596 ( .A(\filter_0/reg_w_4 [0]), .X(n56116) );
  inv_x2_sg U54597 ( .A(\filter_0/reg_w_4 [1]), .X(n56118) );
  inv_x2_sg U54598 ( .A(\filter_0/reg_w_4 [2]), .X(n56120) );
  inv_x2_sg U54599 ( .A(\filter_0/reg_w_4 [3]), .X(n56122) );
  inv_x2_sg U54600 ( .A(\filter_0/reg_w_4 [4]), .X(n56124) );
  inv_x2_sg U54601 ( .A(\filter_0/reg_w_4 [5]), .X(n56126) );
  inv_x2_sg U54602 ( .A(\filter_0/reg_w_4 [6]), .X(n56128) );
  inv_x2_sg U54603 ( .A(\filter_0/reg_w_4 [7]), .X(n56130) );
  inv_x2_sg U54604 ( .A(\filter_0/reg_w_4 [8]), .X(n56132) );
  inv_x2_sg U54605 ( .A(\filter_0/reg_w_4 [9]), .X(n56134) );
  inv_x2_sg U54606 ( .A(\filter_0/reg_w_4 [10]), .X(n56136) );
  inv_x2_sg U54607 ( .A(\filter_0/reg_w_4 [11]), .X(n56138) );
  inv_x2_sg U54608 ( .A(\filter_0/reg_w_4 [12]), .X(n56140) );
  inv_x2_sg U54609 ( .A(\filter_0/reg_w_4 [13]), .X(n56142) );
  inv_x2_sg U54610 ( .A(\filter_0/reg_w_4 [14]), .X(n56144) );
  inv_x2_sg U54611 ( .A(\filter_0/reg_w_4 [15]), .X(n56146) );
  inv_x2_sg U54612 ( .A(\filter_0/reg_w_4 [16]), .X(n56148) );
  inv_x2_sg U54613 ( .A(\filter_0/reg_w_4 [17]), .X(n56150) );
  inv_x2_sg U54614 ( .A(\filter_0/reg_w_4 [18]), .X(n56152) );
  inv_x2_sg U54615 ( .A(\filter_0/reg_w_4 [19]), .X(n56154) );
  inv_x2_sg U54616 ( .A(\filter_0/reg_w_5 [0]), .X(n56156) );
  inv_x2_sg U54617 ( .A(\filter_0/reg_w_5 [1]), .X(n56158) );
  inv_x2_sg U54618 ( .A(\filter_0/reg_w_5 [2]), .X(n56160) );
  inv_x2_sg U54619 ( .A(\filter_0/reg_w_5 [3]), .X(n56162) );
  inv_x2_sg U54620 ( .A(\filter_0/reg_w_5 [4]), .X(n56164) );
  inv_x2_sg U54621 ( .A(\filter_0/reg_w_5 [5]), .X(n56166) );
  inv_x2_sg U54622 ( .A(\filter_0/reg_w_5 [6]), .X(n56168) );
  inv_x2_sg U54623 ( .A(\filter_0/reg_w_5 [7]), .X(n56170) );
  inv_x2_sg U54624 ( .A(\filter_0/reg_w_5 [8]), .X(n56172) );
  inv_x2_sg U54625 ( .A(\filter_0/reg_w_5 [9]), .X(n56174) );
  inv_x2_sg U54626 ( .A(\filter_0/reg_w_5 [10]), .X(n56176) );
  inv_x2_sg U54627 ( .A(\filter_0/reg_w_5 [11]), .X(n56178) );
  inv_x2_sg U54628 ( .A(\filter_0/reg_w_5 [12]), .X(n56180) );
  inv_x2_sg U54629 ( .A(\filter_0/reg_w_5 [13]), .X(n56182) );
  inv_x2_sg U54630 ( .A(\filter_0/reg_w_5 [14]), .X(n56184) );
  inv_x2_sg U54631 ( .A(\filter_0/reg_w_5 [15]), .X(n56186) );
  inv_x2_sg U54632 ( .A(\filter_0/reg_w_5 [16]), .X(n56188) );
  inv_x2_sg U54633 ( .A(\filter_0/reg_w_5 [17]), .X(n56190) );
  inv_x2_sg U54634 ( .A(\filter_0/reg_w_5 [18]), .X(n56192) );
  inv_x2_sg U54635 ( .A(\filter_0/reg_w_5 [19]), .X(n56194) );
  inv_x2_sg U54636 ( .A(\filter_0/reg_w_6 [0]), .X(n56196) );
  inv_x2_sg U54637 ( .A(\filter_0/reg_w_6 [1]), .X(n56198) );
  inv_x2_sg U54638 ( .A(\filter_0/reg_w_6 [2]), .X(n56200) );
  inv_x2_sg U54639 ( .A(\filter_0/reg_w_6 [3]), .X(n56202) );
  inv_x2_sg U54640 ( .A(\filter_0/reg_w_6 [4]), .X(n56204) );
  inv_x2_sg U54641 ( .A(\filter_0/reg_w_6 [5]), .X(n56206) );
  inv_x2_sg U54642 ( .A(\filter_0/reg_w_6 [6]), .X(n56208) );
  inv_x2_sg U54643 ( .A(\filter_0/reg_w_6 [7]), .X(n56210) );
  inv_x2_sg U54644 ( .A(\filter_0/reg_w_6 [8]), .X(n56212) );
  inv_x2_sg U54645 ( .A(\filter_0/reg_w_6 [9]), .X(n56214) );
  inv_x2_sg U54646 ( .A(\filter_0/reg_w_6 [10]), .X(n56216) );
  inv_x2_sg U54647 ( .A(\filter_0/reg_w_6 [11]), .X(n56218) );
  inv_x2_sg U54648 ( .A(\filter_0/reg_w_6 [12]), .X(n56220) );
  inv_x2_sg U54649 ( .A(\filter_0/reg_w_6 [13]), .X(n56222) );
  inv_x2_sg U54650 ( .A(\filter_0/reg_w_6 [14]), .X(n56224) );
  inv_x2_sg U54651 ( .A(\filter_0/reg_w_6 [15]), .X(n56226) );
  inv_x2_sg U54652 ( .A(\filter_0/reg_w_6 [16]), .X(n56228) );
  inv_x2_sg U54653 ( .A(\filter_0/reg_w_6 [17]), .X(n56230) );
  inv_x2_sg U54654 ( .A(\filter_0/reg_w_6 [18]), .X(n56232) );
  inv_x2_sg U54655 ( .A(\filter_0/reg_w_6 [19]), .X(n56234) );
  inv_x2_sg U54656 ( .A(\filter_0/reg_w_7 [0]), .X(n56236) );
  inv_x2_sg U54657 ( .A(\filter_0/reg_w_7 [1]), .X(n56238) );
  inv_x2_sg U54658 ( .A(\filter_0/reg_w_7 [2]), .X(n56240) );
  inv_x2_sg U54659 ( .A(\filter_0/reg_w_7 [3]), .X(n56242) );
  inv_x2_sg U54660 ( .A(\filter_0/reg_w_7 [4]), .X(n56244) );
  inv_x2_sg U54661 ( .A(\filter_0/reg_w_7 [5]), .X(n56246) );
  inv_x2_sg U54662 ( .A(\filter_0/reg_w_7 [6]), .X(n56248) );
  inv_x2_sg U54663 ( .A(\filter_0/reg_w_7 [7]), .X(n56250) );
  inv_x2_sg U54664 ( .A(\filter_0/reg_w_7 [8]), .X(n56252) );
  inv_x2_sg U54665 ( .A(\filter_0/reg_w_7 [9]), .X(n56254) );
  inv_x2_sg U54666 ( .A(\filter_0/reg_w_7 [10]), .X(n56256) );
  inv_x2_sg U54667 ( .A(\filter_0/reg_w_7 [11]), .X(n56258) );
  inv_x2_sg U54668 ( .A(\filter_0/reg_w_7 [12]), .X(n56260) );
  inv_x2_sg U54669 ( .A(\filter_0/reg_w_7 [13]), .X(n56262) );
  inv_x2_sg U54670 ( .A(\filter_0/reg_w_7 [14]), .X(n56264) );
  inv_x2_sg U54671 ( .A(\filter_0/reg_w_7 [15]), .X(n56266) );
  inv_x2_sg U54672 ( .A(\filter_0/reg_w_7 [16]), .X(n56268) );
  inv_x2_sg U54673 ( .A(\filter_0/reg_w_7 [17]), .X(n56270) );
  inv_x2_sg U54674 ( .A(\filter_0/reg_w_7 [18]), .X(n56272) );
  inv_x2_sg U54675 ( .A(\filter_0/reg_w_7 [19]), .X(n56274) );
  inv_x2_sg U54676 ( .A(\filter_0/reg_w_8 [0]), .X(n56276) );
  inv_x2_sg U54677 ( .A(\filter_0/reg_w_8 [1]), .X(n56278) );
  inv_x2_sg U54678 ( .A(\filter_0/reg_w_8 [2]), .X(n56280) );
  inv_x2_sg U54679 ( .A(\filter_0/reg_w_8 [3]), .X(n56282) );
  inv_x2_sg U54680 ( .A(\filter_0/reg_w_8 [4]), .X(n56284) );
  inv_x2_sg U54681 ( .A(\filter_0/reg_w_8 [5]), .X(n56286) );
  inv_x2_sg U54682 ( .A(\filter_0/reg_w_8 [6]), .X(n56288) );
  inv_x2_sg U54683 ( .A(\filter_0/reg_w_8 [7]), .X(n56290) );
  inv_x2_sg U54684 ( .A(\filter_0/reg_w_8 [8]), .X(n56292) );
  inv_x2_sg U54685 ( .A(\filter_0/reg_w_8 [9]), .X(n56294) );
  inv_x2_sg U54686 ( .A(\filter_0/reg_w_8 [10]), .X(n56296) );
  inv_x2_sg U54687 ( .A(\filter_0/reg_w_8 [11]), .X(n56298) );
  inv_x2_sg U54688 ( .A(\filter_0/reg_w_8 [12]), .X(n56300) );
  inv_x2_sg U54689 ( .A(\filter_0/reg_w_8 [13]), .X(n56302) );
  inv_x2_sg U54690 ( .A(\filter_0/reg_w_8 [14]), .X(n56304) );
  inv_x2_sg U54691 ( .A(\filter_0/reg_w_8 [15]), .X(n56306) );
  inv_x2_sg U54692 ( .A(\filter_0/reg_w_8 [16]), .X(n56308) );
  inv_x2_sg U54693 ( .A(\filter_0/reg_w_8 [17]), .X(n56310) );
  inv_x2_sg U54694 ( .A(\filter_0/reg_w_8 [18]), .X(n56312) );
  inv_x2_sg U54695 ( .A(\filter_0/reg_w_8 [19]), .X(n56314) );
  inv_x2_sg U54696 ( .A(\filter_0/reg_w_9 [0]), .X(n56316) );
  inv_x2_sg U54697 ( .A(\filter_0/reg_w_9 [1]), .X(n56318) );
  inv_x2_sg U54698 ( .A(\filter_0/reg_w_9 [2]), .X(n56320) );
  inv_x2_sg U54699 ( .A(\filter_0/reg_w_9 [3]), .X(n56322) );
  inv_x2_sg U54700 ( .A(\filter_0/reg_w_9 [4]), .X(n56324) );
  inv_x2_sg U54701 ( .A(\filter_0/reg_w_9 [5]), .X(n56326) );
  inv_x2_sg U54702 ( .A(\filter_0/reg_w_9 [6]), .X(n56328) );
  inv_x2_sg U54703 ( .A(\filter_0/reg_w_9 [7]), .X(n56330) );
  inv_x2_sg U54704 ( .A(\filter_0/reg_w_9 [8]), .X(n56332) );
  inv_x2_sg U54705 ( .A(\filter_0/reg_w_9 [9]), .X(n56334) );
  inv_x2_sg U54706 ( .A(\filter_0/reg_w_9 [10]), .X(n56336) );
  inv_x2_sg U54707 ( .A(\filter_0/reg_w_9 [11]), .X(n56338) );
  inv_x2_sg U54708 ( .A(\filter_0/reg_w_9 [12]), .X(n56340) );
  inv_x2_sg U54709 ( .A(\filter_0/reg_w_9 [13]), .X(n56342) );
  inv_x2_sg U54710 ( .A(\filter_0/reg_w_9 [14]), .X(n56344) );
  inv_x2_sg U54711 ( .A(\filter_0/reg_w_9 [15]), .X(n56346) );
  inv_x2_sg U54712 ( .A(\filter_0/reg_w_9 [16]), .X(n56348) );
  inv_x2_sg U54713 ( .A(\filter_0/reg_w_9 [17]), .X(n56350) );
  inv_x2_sg U54714 ( .A(\filter_0/reg_w_9 [18]), .X(n56352) );
  inv_x2_sg U54715 ( .A(\filter_0/reg_w_9 [19]), .X(n56354) );
  inv_x2_sg U54716 ( .A(\filter_0/reg_w_10 [0]), .X(n56356) );
  inv_x2_sg U54717 ( .A(\filter_0/reg_w_10 [1]), .X(n56358) );
  inv_x2_sg U54718 ( .A(\filter_0/reg_w_10 [2]), .X(n56360) );
  inv_x2_sg U54719 ( .A(\filter_0/reg_w_10 [3]), .X(n56362) );
  inv_x2_sg U54720 ( .A(\filter_0/reg_w_10 [4]), .X(n56364) );
  inv_x2_sg U54721 ( .A(\filter_0/reg_w_10 [5]), .X(n56366) );
  inv_x2_sg U54722 ( .A(\filter_0/reg_w_10 [6]), .X(n56368) );
  inv_x2_sg U54723 ( .A(\filter_0/reg_w_10 [7]), .X(n56370) );
  inv_x2_sg U54724 ( .A(\filter_0/reg_w_10 [8]), .X(n56372) );
  inv_x2_sg U54725 ( .A(\filter_0/reg_w_10 [9]), .X(n56374) );
  inv_x2_sg U54726 ( .A(\filter_0/reg_w_10 [10]), .X(n56376) );
  inv_x2_sg U54727 ( .A(\filter_0/reg_w_10 [11]), .X(n56378) );
  inv_x2_sg U54728 ( .A(\filter_0/reg_w_10 [12]), .X(n56380) );
  inv_x2_sg U54729 ( .A(\filter_0/reg_w_10 [13]), .X(n56382) );
  inv_x2_sg U54730 ( .A(\filter_0/reg_w_10 [14]), .X(n56384) );
  inv_x2_sg U54731 ( .A(\filter_0/reg_w_10 [15]), .X(n56386) );
  inv_x2_sg U54732 ( .A(\filter_0/reg_w_10 [16]), .X(n56388) );
  inv_x2_sg U54733 ( .A(\filter_0/reg_w_10 [17]), .X(n56390) );
  inv_x2_sg U54734 ( .A(\filter_0/reg_w_10 [18]), .X(n56392) );
  inv_x2_sg U54735 ( .A(\filter_0/reg_w_10 [19]), .X(n56394) );
  inv_x2_sg U54736 ( .A(\filter_0/reg_w_11 [0]), .X(n56396) );
  inv_x2_sg U54737 ( .A(\filter_0/reg_w_11 [1]), .X(n56398) );
  inv_x2_sg U54738 ( .A(\filter_0/reg_w_11 [2]), .X(n56400) );
  inv_x2_sg U54739 ( .A(\filter_0/reg_w_11 [3]), .X(n56402) );
  inv_x2_sg U54740 ( .A(\filter_0/reg_w_11 [4]), .X(n56404) );
  inv_x2_sg U54741 ( .A(\filter_0/reg_w_11 [5]), .X(n56406) );
  inv_x2_sg U54742 ( .A(\filter_0/reg_w_11 [6]), .X(n56408) );
  inv_x2_sg U54743 ( .A(\filter_0/reg_w_11 [7]), .X(n56410) );
  inv_x2_sg U54744 ( .A(\filter_0/reg_w_11 [8]), .X(n56412) );
  inv_x2_sg U54745 ( .A(\filter_0/reg_w_11 [9]), .X(n56414) );
  inv_x2_sg U54746 ( .A(\filter_0/reg_w_11 [10]), .X(n56416) );
  inv_x2_sg U54747 ( .A(\filter_0/reg_w_11 [11]), .X(n56418) );
  inv_x2_sg U54748 ( .A(\filter_0/reg_w_11 [12]), .X(n56420) );
  inv_x2_sg U54749 ( .A(\filter_0/reg_w_11 [13]), .X(n56422) );
  inv_x2_sg U54750 ( .A(\filter_0/reg_w_11 [14]), .X(n56424) );
  inv_x2_sg U54751 ( .A(\filter_0/reg_w_11 [15]), .X(n56426) );
  inv_x2_sg U54752 ( .A(\filter_0/reg_w_11 [16]), .X(n56428) );
  inv_x2_sg U54753 ( .A(\filter_0/reg_w_11 [17]), .X(n56430) );
  inv_x2_sg U54754 ( .A(\filter_0/reg_w_11 [18]), .X(n56432) );
  inv_x2_sg U54755 ( .A(\filter_0/reg_w_11 [19]), .X(n56434) );
  inv_x2_sg U54756 ( .A(\filter_0/reg_w_12 [0]), .X(n56436) );
  inv_x2_sg U54757 ( .A(\filter_0/reg_w_12 [1]), .X(n56438) );
  inv_x2_sg U54758 ( .A(\filter_0/reg_w_12 [2]), .X(n56440) );
  inv_x2_sg U54759 ( .A(\filter_0/reg_w_12 [3]), .X(n56442) );
  inv_x2_sg U54760 ( .A(\filter_0/reg_w_12 [4]), .X(n56444) );
  inv_x2_sg U54761 ( .A(\filter_0/reg_w_12 [5]), .X(n56446) );
  inv_x2_sg U54762 ( .A(\filter_0/reg_w_12 [6]), .X(n56448) );
  inv_x2_sg U54763 ( .A(\filter_0/reg_w_12 [7]), .X(n56450) );
  inv_x2_sg U54764 ( .A(\filter_0/reg_w_12 [8]), .X(n56452) );
  inv_x2_sg U54765 ( .A(\filter_0/reg_w_12 [9]), .X(n56454) );
  inv_x2_sg U54766 ( .A(\filter_0/reg_w_12 [10]), .X(n56456) );
  inv_x2_sg U54767 ( .A(\filter_0/reg_w_12 [11]), .X(n56458) );
  inv_x2_sg U54768 ( .A(\filter_0/reg_w_12 [12]), .X(n56460) );
  inv_x2_sg U54769 ( .A(\filter_0/reg_w_12 [13]), .X(n56462) );
  inv_x2_sg U54770 ( .A(\filter_0/reg_w_12 [14]), .X(n56464) );
  inv_x2_sg U54771 ( .A(\filter_0/reg_w_12 [15]), .X(n56466) );
  inv_x2_sg U54772 ( .A(\filter_0/reg_w_12 [16]), .X(n56468) );
  inv_x2_sg U54773 ( .A(\filter_0/reg_w_12 [17]), .X(n56470) );
  inv_x2_sg U54774 ( .A(\filter_0/reg_w_12 [18]), .X(n56472) );
  inv_x2_sg U54775 ( .A(\filter_0/reg_w_12 [19]), .X(n56474) );
  inv_x2_sg U54776 ( .A(\filter_0/reg_w_13 [0]), .X(n56476) );
  inv_x2_sg U54777 ( .A(\filter_0/reg_w_13 [1]), .X(n56478) );
  inv_x2_sg U54778 ( .A(\filter_0/reg_w_13 [2]), .X(n56480) );
  inv_x2_sg U54779 ( .A(\filter_0/reg_w_13 [3]), .X(n56482) );
  inv_x2_sg U54780 ( .A(\filter_0/reg_w_13 [4]), .X(n56484) );
  inv_x2_sg U54781 ( .A(\filter_0/reg_w_13 [5]), .X(n56486) );
  inv_x2_sg U54782 ( .A(\filter_0/reg_w_13 [6]), .X(n56488) );
  inv_x2_sg U54783 ( .A(\filter_0/reg_w_13 [7]), .X(n56490) );
  inv_x2_sg U54784 ( .A(\filter_0/reg_w_13 [8]), .X(n56492) );
  inv_x2_sg U54785 ( .A(\filter_0/reg_w_13 [9]), .X(n56494) );
  inv_x2_sg U54786 ( .A(\filter_0/reg_w_13 [10]), .X(n56496) );
  inv_x2_sg U54787 ( .A(\filter_0/reg_w_13 [11]), .X(n56498) );
  inv_x2_sg U54788 ( .A(\filter_0/reg_w_13 [12]), .X(n56500) );
  inv_x2_sg U54789 ( .A(\filter_0/reg_w_13 [13]), .X(n56502) );
  inv_x2_sg U54790 ( .A(\filter_0/reg_w_13 [14]), .X(n56504) );
  inv_x2_sg U54791 ( .A(\filter_0/reg_w_13 [15]), .X(n56506) );
  inv_x2_sg U54792 ( .A(\filter_0/reg_w_13 [16]), .X(n56508) );
  inv_x2_sg U54793 ( .A(\filter_0/reg_w_13 [17]), .X(n56510) );
  inv_x2_sg U54794 ( .A(\filter_0/reg_w_13 [18]), .X(n56512) );
  inv_x2_sg U54795 ( .A(\filter_0/reg_w_13 [19]), .X(n56514) );
  inv_x2_sg U54796 ( .A(\filter_0/reg_w_14 [0]), .X(n56516) );
  inv_x2_sg U54797 ( .A(\filter_0/reg_w_14 [1]), .X(n56518) );
  inv_x2_sg U54798 ( .A(\filter_0/reg_w_14 [2]), .X(n56520) );
  inv_x2_sg U54799 ( .A(\filter_0/reg_w_14 [3]), .X(n56522) );
  inv_x2_sg U54800 ( .A(\filter_0/reg_w_14 [4]), .X(n56524) );
  inv_x2_sg U54801 ( .A(\filter_0/reg_w_14 [5]), .X(n56526) );
  inv_x2_sg U54802 ( .A(\filter_0/reg_w_14 [6]), .X(n56528) );
  inv_x2_sg U54803 ( .A(\filter_0/reg_w_14 [7]), .X(n56530) );
  inv_x2_sg U54804 ( .A(\filter_0/reg_w_14 [8]), .X(n56532) );
  inv_x2_sg U54805 ( .A(\filter_0/reg_w_14 [9]), .X(n56534) );
  inv_x2_sg U54806 ( .A(\filter_0/reg_w_14 [10]), .X(n56536) );
  inv_x2_sg U54807 ( .A(\filter_0/reg_w_14 [11]), .X(n56538) );
  inv_x2_sg U54808 ( .A(\filter_0/reg_w_14 [12]), .X(n56540) );
  inv_x2_sg U54809 ( .A(\filter_0/reg_w_14 [13]), .X(n56542) );
  inv_x2_sg U54810 ( .A(\filter_0/reg_w_14 [14]), .X(n56544) );
  inv_x2_sg U54811 ( .A(\filter_0/reg_w_14 [15]), .X(n56546) );
  inv_x2_sg U54812 ( .A(\filter_0/reg_w_14 [16]), .X(n56548) );
  inv_x2_sg U54813 ( .A(\filter_0/reg_w_14 [17]), .X(n56550) );
  inv_x2_sg U54814 ( .A(\filter_0/reg_w_14 [18]), .X(n56552) );
  inv_x2_sg U54815 ( .A(\filter_0/reg_w_14 [19]), .X(n56554) );
  inv_x2_sg U54816 ( .A(\filter_0/reg_w_15 [0]), .X(n56556) );
  inv_x2_sg U54817 ( .A(\filter_0/reg_w_15 [1]), .X(n56558) );
  inv_x2_sg U54818 ( .A(\filter_0/reg_w_15 [2]), .X(n56560) );
  inv_x2_sg U54819 ( .A(\filter_0/reg_w_15 [3]), .X(n56562) );
  inv_x2_sg U54820 ( .A(\filter_0/reg_w_15 [4]), .X(n56564) );
  inv_x2_sg U54821 ( .A(\filter_0/reg_w_15 [5]), .X(n56566) );
  inv_x2_sg U54822 ( .A(\filter_0/reg_w_15 [6]), .X(n56568) );
  inv_x2_sg U54823 ( .A(\filter_0/reg_w_15 [7]), .X(n56570) );
  inv_x2_sg U54824 ( .A(\filter_0/reg_w_15 [8]), .X(n56572) );
  inv_x2_sg U54825 ( .A(\filter_0/reg_w_15 [9]), .X(n56574) );
  inv_x2_sg U54826 ( .A(\filter_0/reg_w_15 [10]), .X(n56576) );
  inv_x2_sg U54827 ( .A(\filter_0/reg_w_15 [11]), .X(n56578) );
  inv_x2_sg U54828 ( .A(\filter_0/reg_w_15 [12]), .X(n56580) );
  inv_x2_sg U54829 ( .A(\filter_0/reg_w_15 [13]), .X(n56582) );
  inv_x2_sg U54830 ( .A(\filter_0/reg_w_15 [14]), .X(n56584) );
  inv_x2_sg U54831 ( .A(\filter_0/reg_w_15 [15]), .X(n56586) );
  inv_x2_sg U54832 ( .A(\filter_0/reg_w_15 [16]), .X(n56588) );
  inv_x2_sg U54833 ( .A(\filter_0/reg_w_15 [17]), .X(n56590) );
  inv_x2_sg U54834 ( .A(\filter_0/reg_w_15 [18]), .X(n56592) );
  inv_x2_sg U54835 ( .A(\filter_0/reg_w_15 [19]), .X(n56594) );
  inv_x2_sg U54836 ( .A(\filter_0/reg_o_mask [0]), .X(n51066) );
  inv_x2_sg U54837 ( .A(\filter_0/reg_o_mask [1]), .X(n51068) );
  inv_x2_sg U54838 ( .A(\filter_0/reg_o_mask [18]), .X(n51058) );
  inv_x2_sg U54839 ( .A(\shifter_0/reg_w_9 [7]), .X(n51214) );
  inv_x2_sg U54840 ( .A(\shifter_0/reg_w_10 [7]), .X(n51216) );
  inv_x2_sg U54841 ( .A(\shifter_0/reg_i_4 [15]), .X(n55084) );
  inv_x2_sg U54842 ( .A(\shifter_0/reg_w_4 [15]), .X(n55086) );
  inv_x2_sg U54843 ( .A(\mask_0/reg_ii_mask [1]), .X(n55088) );
  inv_x2_sg U54844 ( .A(\mask_0/reg_ii_mask [2]), .X(n55090) );
  inv_x2_sg U54845 ( .A(\mask_0/reg_ii_mask [3]), .X(n55092) );
  inv_x2_sg U54846 ( .A(\mask_0/reg_ii_mask [6]), .X(n55094) );
  inv_x2_sg U54847 ( .A(\mask_0/reg_ii_mask [7]), .X(n55096) );
  inv_x2_sg U54848 ( .A(\mask_0/reg_ii_mask [8]), .X(n55098) );
  inv_x2_sg U54849 ( .A(\mask_0/reg_ii_mask [9]), .X(n55100) );
  inv_x2_sg U54850 ( .A(\mask_0/reg_ii_mask [10]), .X(n55102) );
  inv_x2_sg U54851 ( .A(\mask_0/reg_ii_mask [11]), .X(n55104) );
  inv_x2_sg U54852 ( .A(\mask_0/reg_ii_mask [12]), .X(n55106) );
  inv_x2_sg U54853 ( .A(\mask_0/reg_ii_mask [13]), .X(n55108) );
  inv_x2_sg U54854 ( .A(\mask_0/reg_ii_mask [14]), .X(n55110) );
  inv_x2_sg U54855 ( .A(\mask_0/reg_ii_mask [15]), .X(n55112) );
  inv_x2_sg U54856 ( .A(\mask_0/reg_ii_mask [16]), .X(n55114) );
  inv_x2_sg U54857 ( .A(\mask_0/reg_ii_mask [18]), .X(n55116) );
  inv_x2_sg U54858 ( .A(\mask_0/reg_ii_mask [19]), .X(n55118) );
  inv_x2_sg U54859 ( .A(\mask_0/reg_ii_mask [20]), .X(n55120) );
  inv_x2_sg U54860 ( .A(\mask_0/reg_ii_mask [21]), .X(n55122) );
  inv_x2_sg U54861 ( .A(\mask_0/reg_ii_mask [22]), .X(n55124) );
  inv_x2_sg U54862 ( .A(\mask_0/reg_ii_mask [23]), .X(n55126) );
  inv_x2_sg U54863 ( .A(\mask_0/reg_ii_mask [24]), .X(n55128) );
  inv_x2_sg U54864 ( .A(\mask_0/reg_ii_mask [25]), .X(n55130) );
  inv_x2_sg U54865 ( .A(\mask_0/reg_ii_mask [26]), .X(n55132) );
  inv_x2_sg U54866 ( .A(\mask_0/reg_ii_mask [27]), .X(n55134) );
  inv_x2_sg U54867 ( .A(\mask_0/reg_ww_mask [0]), .X(n55136) );
  inv_x2_sg U54868 ( .A(\mask_0/reg_ww_mask [4]), .X(n55138) );
  inv_x2_sg U54869 ( .A(\mask_0/reg_ww_mask [5]), .X(n55140) );
  inv_x2_sg U54870 ( .A(\mask_0/reg_ww_mask [17]), .X(n55142) );
  inv_x2_sg U54871 ( .A(\mask_0/reg_ww_mask [28]), .X(n55144) );
  inv_x2_sg U54872 ( .A(\mask_0/reg_ww_mask [29]), .X(n55146) );
  inv_x2_sg U54873 ( .A(\mask_0/reg_ww_mask [30]), .X(n55148) );
  inv_x2_sg U54874 ( .A(\mask_0/reg_ww_mask [31]), .X(n55150) );
  inv_x2_sg U54875 ( .A(\filter_0/reg_o_mask [2]), .X(n51060) );
  inv_x2_sg U54876 ( .A(\shifter_0/reg_i_0 [10]), .X(n55252) );
  inv_x2_sg U54877 ( .A(\shifter_0/reg_i_0 [19]), .X(n55254) );
  inv_x2_sg U54878 ( .A(\shifter_0/reg_w_0 [10]), .X(n55256) );
  inv_x2_sg U54879 ( .A(\shifter_0/reg_w_0 [19]), .X(n55258) );
  inv_x2_sg U54880 ( .A(\shifter_0/reg_i_4 [3]), .X(n54998) );
  inv_x2_sg U54881 ( .A(\shifter_0/reg_i_4 [4]), .X(n55000) );
  inv_x2_sg U54882 ( .A(\shifter_0/reg_i_4 [8]), .X(n55002) );
  inv_x2_sg U54883 ( .A(\shifter_0/reg_i_4 [9]), .X(n55004) );
  inv_x2_sg U54884 ( .A(\shifter_0/reg_i_4 [12]), .X(n55006) );
  inv_x2_sg U54885 ( .A(\shifter_0/reg_i_4 [13]), .X(n55008) );
  inv_x2_sg U54886 ( .A(\shifter_0/reg_w_4 [3]), .X(n55010) );
  inv_x2_sg U54887 ( .A(\shifter_0/reg_w_4 [4]), .X(n55012) );
  inv_x2_sg U54888 ( .A(\shifter_0/reg_w_4 [8]), .X(n55014) );
  inv_x2_sg U54889 ( .A(\shifter_0/reg_w_4 [9]), .X(n55016) );
  inv_x2_sg U54890 ( .A(\shifter_0/reg_w_4 [12]), .X(n55018) );
  inv_x2_sg U54891 ( .A(\shifter_0/reg_w_4 [13]), .X(n55020) );
  inv_x2_sg U54892 ( .A(\shifter_0/reg_i_14 [13]), .X(n56718) );
  inv_x2_sg U54893 ( .A(\shifter_0/reg_w_9 [4]), .X(n51258) );
  inv_x2_sg U54894 ( .A(\shifter_0/reg_w_14 [4]), .X(n56738) );
  inv_x2_sg U54895 ( .A(\shifter_0/reg_i_9 [7]), .X(n51278) );
  inv_x2_sg U54896 ( .A(\shifter_0/reg_i_9 [11]), .X(n51280) );
  inv_x2_sg U54897 ( .A(\shifter_0/reg_i_10 [7]), .X(n51284) );
  inv_x2_sg U54898 ( .A(\shifter_0/reg_i_10 [11]), .X(n51286) );
  inv_x2_sg U54899 ( .A(\shifter_0/reg_i_11 [14]), .X(n51296) );
  inv_x2_sg U54900 ( .A(\shifter_0/reg_w_9 [11]), .X(n51304) );
  inv_x2_sg U54901 ( .A(\shifter_0/reg_w_10 [11]), .X(n51308) );
  inv_x2_sg U54902 ( .A(\shifter_0/reg_w_11 [14]), .X(n51314) );
  inv_x2_sg U54903 ( .A(\shifter_0/reg_i_9 [19]), .X(n51320) );
  inv_x2_sg U54904 ( .A(\shifter_0/reg_w_9 [19]), .X(n51324) );
  inv_x2_sg U54905 ( .A(\shifter_0/reg_w_10 [19]), .X(n51326) );
  inv_x2_sg U54906 ( .A(\shifter_0/reg_i_0 [3]), .X(n55022) );
  inv_x2_sg U54907 ( .A(\shifter_0/reg_i_0 [4]), .X(n55024) );
  inv_x2_sg U54908 ( .A(\shifter_0/reg_i_0 [8]), .X(n55026) );
  inv_x2_sg U54909 ( .A(\shifter_0/reg_i_0 [9]), .X(n55028) );
  inv_x2_sg U54910 ( .A(\shifter_0/reg_i_0 [12]), .X(n55030) );
  inv_x2_sg U54911 ( .A(\shifter_0/reg_i_0 [13]), .X(n55032) );
  inv_x2_sg U54912 ( .A(\shifter_0/reg_i_0 [17]), .X(n55034) );
  inv_x2_sg U54913 ( .A(\shifter_0/reg_i_0 [18]), .X(n55036) );
  inv_x2_sg U54914 ( .A(\shifter_0/reg_i_4 [17]), .X(n55038) );
  inv_x2_sg U54915 ( .A(\shifter_0/reg_i_4 [18]), .X(n55040) );
  inv_x2_sg U54916 ( .A(\shifter_0/reg_w_0 [3]), .X(n55042) );
  inv_x2_sg U54917 ( .A(\shifter_0/reg_w_0 [4]), .X(n55044) );
  inv_x2_sg U54918 ( .A(\shifter_0/reg_w_0 [8]), .X(n55046) );
  inv_x2_sg U54919 ( .A(\shifter_0/reg_w_0 [9]), .X(n55048) );
  inv_x2_sg U54920 ( .A(\shifter_0/reg_w_0 [12]), .X(n55050) );
  inv_x2_sg U54921 ( .A(\shifter_0/reg_w_0 [13]), .X(n55052) );
  inv_x2_sg U54922 ( .A(\shifter_0/reg_w_0 [17]), .X(n55054) );
  inv_x2_sg U54923 ( .A(\shifter_0/reg_w_0 [18]), .X(n55056) );
  inv_x2_sg U54924 ( .A(\shifter_0/reg_w_4 [17]), .X(n55058) );
  inv_x2_sg U54925 ( .A(\shifter_0/reg_w_4 [18]), .X(n55060) );
  inv_x2_sg U54926 ( .A(\shifter_0/reg_i_5 [4]), .X(n56778) );
  inv_x2_sg U54927 ( .A(\shifter_0/reg_i_5 [9]), .X(n56780) );
  inv_x2_sg U54928 ( .A(\shifter_0/reg_i_5 [13]), .X(n56782) );
  inv_x2_sg U54929 ( .A(\shifter_0/reg_w_5 [4]), .X(n56784) );
  inv_x2_sg U54930 ( .A(\shifter_0/reg_w_5 [9]), .X(n56786) );
  inv_x2_sg U54931 ( .A(\shifter_0/reg_w_5 [13]), .X(n56788) );
  inv_x2_sg U54932 ( .A(\shifter_0/reg_i_9 [4]), .X(n51342) );
  inv_x2_sg U54933 ( .A(\shifter_0/reg_i_9 [9]), .X(n51344) );
  inv_x2_sg U54934 ( .A(\shifter_0/reg_i_9 [13]), .X(n51346) );
  inv_x2_sg U54935 ( .A(\shifter_0/reg_i_10 [9]), .X(n51350) );
  inv_x2_sg U54936 ( .A(\shifter_0/reg_i_14 [4]), .X(n56808) );
  inv_x2_sg U54937 ( .A(\shifter_0/reg_w_9 [9]), .X(n51364) );
  inv_x2_sg U54938 ( .A(\shifter_0/reg_w_9 [13]), .X(n51366) );
  inv_x2_sg U54939 ( .A(\shifter_0/reg_w_10 [9]), .X(n51368) );
  inv_x2_sg U54940 ( .A(\shifter_0/reg_w_14 [13]), .X(n56822) );
  inv_x2_sg U54941 ( .A(\shifter_0/reg_i_1 [3]), .X(n55284) );
  inv_x2_sg U54942 ( .A(\shifter_0/reg_i_1 [4]), .X(n55286) );
  inv_x2_sg U54943 ( .A(\shifter_0/reg_i_1 [8]), .X(n55288) );
  inv_x2_sg U54944 ( .A(\shifter_0/reg_i_1 [9]), .X(n55290) );
  inv_x2_sg U54945 ( .A(\shifter_0/reg_i_1 [12]), .X(n55292) );
  inv_x2_sg U54946 ( .A(\shifter_0/reg_i_1 [13]), .X(n55294) );
  inv_x2_sg U54947 ( .A(\shifter_0/reg_w_1 [3]), .X(n55296) );
  inv_x2_sg U54948 ( .A(\shifter_0/reg_w_1 [4]), .X(n55298) );
  inv_x2_sg U54949 ( .A(\shifter_0/reg_w_1 [8]), .X(n55300) );
  inv_x2_sg U54950 ( .A(\shifter_0/reg_w_1 [9]), .X(n55302) );
  inv_x2_sg U54951 ( .A(\shifter_0/reg_w_1 [12]), .X(n55304) );
  inv_x2_sg U54952 ( .A(\shifter_0/reg_w_1 [13]), .X(n55306) );
  inv_x2_sg U54953 ( .A(\shifter_0/reg_i_1 [17]), .X(n55308) );
  inv_x2_sg U54954 ( .A(\shifter_0/reg_i_1 [18]), .X(n55310) );
  inv_x2_sg U54955 ( .A(\shifter_0/reg_w_1 [17]), .X(n55312) );
  inv_x2_sg U54956 ( .A(\shifter_0/reg_w_1 [18]), .X(n55314) );
  inv_x2_sg U54957 ( .A(\shifter_0/reg_i_4 [16]), .X(n55152) );
  inv_x2_sg U54958 ( .A(\shifter_0/reg_w_4 [16]), .X(n55154) );
  inv_x2_sg U54959 ( .A(\shifter_0/reg_i_0 [2]), .X(n55260) );
  inv_x2_sg U54960 ( .A(\shifter_0/reg_i_0 [6]), .X(n55262) );
  inv_x2_sg U54961 ( .A(\shifter_0/reg_i_0 [7]), .X(n55264) );
  inv_x2_sg U54962 ( .A(\shifter_0/reg_i_0 [11]), .X(n55266) );
  inv_x2_sg U54963 ( .A(\shifter_0/reg_i_0 [15]), .X(n55268) );
  inv_x2_sg U54964 ( .A(\shifter_0/reg_i_5 [15]), .X(n56828) );
  inv_x2_sg U54965 ( .A(\shifter_0/reg_w_0 [2]), .X(n55272) );
  inv_x2_sg U54966 ( .A(\shifter_0/reg_w_0 [6]), .X(n55274) );
  inv_x2_sg U54967 ( .A(\shifter_0/reg_w_0 [7]), .X(n55276) );
  inv_x2_sg U54968 ( .A(\shifter_0/reg_w_0 [11]), .X(n55278) );
  inv_x2_sg U54969 ( .A(\shifter_0/reg_w_0 [15]), .X(n55280) );
  inv_x2_sg U54970 ( .A(\shifter_0/reg_w_5 [15]), .X(n56840) );
  inv_x2_sg U54971 ( .A(\mask_0/counter [1]), .X(n51198) );
  inv_x2_sg U54972 ( .A(\shifter_0/reg_i_9 [16]), .X(n51414) );
  inv_x2_sg U54973 ( .A(\shifter_0/reg_w_9 [16]), .X(n51418) );
  inv_x2_sg U54974 ( .A(\filter_0/reg_o_mask [3]), .X(n51062) );
  inv_x2_sg U54975 ( .A(\shifter_0/i_pointer [2]), .X(n51052) );
  inv_x2_sg U54976 ( .A(filter_input_ready), .X(n51064) );
  inv_x2_sg U54977 ( .A(\shifter_0/reg_i_2 [3]), .X(n55222) );
  inv_x2_sg U54978 ( .A(\shifter_0/reg_i_2 [7]), .X(n51154) );
  inv_x2_sg U54979 ( .A(\shifter_0/reg_i_2 [8]), .X(n55226) );
  inv_x2_sg U54980 ( .A(\shifter_0/reg_i_2 [11]), .X(n51158) );
  inv_x2_sg U54981 ( .A(\shifter_0/reg_i_2 [12]), .X(n55230) );
  inv_x2_sg U54982 ( .A(\shifter_0/reg_i_6 [7]), .X(n51424) );
  inv_x2_sg U54983 ( .A(\shifter_0/reg_i_6 [11]), .X(n51426) );
  inv_x2_sg U54984 ( .A(\shifter_0/reg_i_6 [15]), .X(n51428) );
  inv_x2_sg U54985 ( .A(\shifter_0/reg_i_6 [19]), .X(n51430) );
  inv_x2_sg U54986 ( .A(\shifter_0/reg_w_2 [7]), .X(n51164) );
  inv_x2_sg U54987 ( .A(\shifter_0/reg_w_2 [11]), .X(n51168) );
  inv_x2_sg U54988 ( .A(\shifter_0/reg_w_6 [7]), .X(n51432) );
  inv_x2_sg U54989 ( .A(\shifter_0/reg_w_6 [11]), .X(n51434) );
  inv_x2_sg U54990 ( .A(\shifter_0/reg_w_6 [15]), .X(n51436) );
  inv_x2_sg U54991 ( .A(\shifter_0/reg_w_6 [19]), .X(n51438) );
  inv_x2_sg U54992 ( .A(\shifter_0/reg_w_2 [3]), .X(n55234) );
  inv_x2_sg U54993 ( .A(\shifter_0/reg_w_2 [8]), .X(n55238) );
  inv_x2_sg U54994 ( .A(\shifter_0/reg_w_2 [12]), .X(n55242) );
  inv_x2_sg U54995 ( .A(\shifter_0/reg_w_2 [19]), .X(n51172) );
  inv_x2_sg U54996 ( .A(\shifter_0/reg_i_2 [14]), .X(n55244) );
  inv_x2_sg U54997 ( .A(\shifter_0/reg_w_2 [14]), .X(n55246) );
  inv_x2_sg U54998 ( .A(\shifter_0/reg_i_2 [18]), .X(n51178) );
  inv_x2_sg U54999 ( .A(\shifter_0/reg_i_3 [4]), .X(n56896) );
  inv_x2_sg U55000 ( .A(\shifter_0/reg_i_3 [9]), .X(n56898) );
  inv_x2_sg U55001 ( .A(\shifter_0/reg_i_3 [13]), .X(n56900) );
  inv_x2_sg U55002 ( .A(\shifter_0/reg_i_3 [15]), .X(n56902) );
  inv_x2_sg U55003 ( .A(\shifter_0/reg_w_2 [18]), .X(n51180) );
  inv_x2_sg U55004 ( .A(\shifter_0/reg_w_3 [4]), .X(n56904) );
  inv_x2_sg U55005 ( .A(\shifter_0/reg_w_3 [9]), .X(n56906) );
  inv_x2_sg U55006 ( .A(\shifter_0/reg_w_3 [13]), .X(n56908) );
  inv_x2_sg U55007 ( .A(\shifter_0/reg_w_3 [15]), .X(n56910) );
  inv_x2_sg U55008 ( .A(n55271), .X(n67488) );
  inv_x2_sg U55009 ( .A(n51193), .X(n67490) );
  inv_x2_sg U55010 ( .A(n51191), .X(n67495) );
  inv_x2_sg U55011 ( .A(n51185), .X(n67497) );
  inv_x2_sg U55012 ( .A(n51183), .X(n67498) );
  inv_x2_sg U55013 ( .A(n55283), .X(n67295) );
  inv_x2_sg U55014 ( .A(n51197), .X(n67297) );
  inv_x2_sg U55015 ( .A(n51195), .X(n67302) );
  inv_x2_sg U55016 ( .A(n51189), .X(n67304) );
  inv_x2_sg U55017 ( .A(n51187), .X(n67305) );
  nor_x2_sg U55018 ( .A(n51499), .B(n22988), .X(n23098) );
  nor_x2_sg U55019 ( .A(n51507), .B(n57152), .X(n23021) );
  nor_x2_sg U55020 ( .A(n51495), .B(n57153), .X(n23010) );
  nor_x2_sg U55021 ( .A(n51503), .B(n22761), .X(n22871) );
  nor_x2_sg U55022 ( .A(n51493), .B(n57158), .X(n22794) );
  nor_x2_sg U55023 ( .A(n51489), .B(n57159), .X(n22783) );
  nor_x4_sg U55024 ( .A(n57168), .B(n57170), .X(n32802) );
  nand_x4_sg U55025 ( .A(n33309), .B(n33094), .X(n34047) );
  nand_x4_sg U55026 ( .A(n33222), .B(n32965), .X(n34135) );
  nor_x4_sg U55027 ( .A(n57917), .B(n57925), .X(n58374) );
  nor_x4_sg U55028 ( .A(n57920), .B(n57922), .X(n58376) );
  inv_x4_sg U55029 ( .A(n58483), .X(n29333) );
  nand_x4_sg U55030 ( .A(n33396), .B(n33782), .X(n33781) );
  inv_x4_sg U55031 ( .A(n47572), .X(n47573) );
  nor_x4_sg U55032 ( .A(n57168), .B(n57557), .X(n34232) );
  inv_x4_sg U55033 ( .A(n22440), .X(n61900) );
  inv_x4_sg U55034 ( .A(n22592), .X(n67355) );
  inv_x4_sg U55035 ( .A(n22589), .X(n67358) );
  inv_x4_sg U55036 ( .A(n22586), .X(n67361) );
  inv_x4_sg U55037 ( .A(n22585), .X(n67362) );
  inv_x4_sg U55038 ( .A(n22583), .X(n67364) );
  inv_x4_sg U55039 ( .A(n22581), .X(n67366) );
  inv_x4_sg U55040 ( .A(n22579), .X(n67368) );
  inv_x4_sg U55041 ( .A(n22577), .X(n67370) );
  inv_x4_sg U55042 ( .A(n22576), .X(n67371) );
  inv_x4_sg U55043 ( .A(n22575), .X(n67372) );
  inv_x4_sg U55044 ( .A(n22563), .X(n67145) );
  inv_x4_sg U55045 ( .A(n22560), .X(n67148) );
  inv_x4_sg U55046 ( .A(n22559), .X(n67149) );
  inv_x4_sg U55047 ( .A(n22557), .X(n67151) );
  inv_x4_sg U55048 ( .A(n22555), .X(n67153) );
  inv_x4_sg U55049 ( .A(n22553), .X(n67155) );
  inv_x4_sg U55050 ( .A(n22551), .X(n67157) );
  inv_x4_sg U55051 ( .A(n22550), .X(n67158) );
  inv_x4_sg U55052 ( .A(n22549), .X(n67159) );
  inv_x4_sg U55053 ( .A(n22493), .X(n67315) );
  inv_x4_sg U55054 ( .A(n22542), .X(n67336) );
  inv_x4_sg U55055 ( .A(n22539), .X(n67339) );
  inv_x4_sg U55056 ( .A(n22535), .X(n67343) );
  inv_x4_sg U55057 ( .A(n22533), .X(n67345) );
  inv_x4_sg U55058 ( .A(n22531), .X(n67347) );
  inv_x4_sg U55059 ( .A(n22518), .X(n67122) );
  inv_x4_sg U55060 ( .A(n22514), .X(n67126) );
  inv_x4_sg U55061 ( .A(n22510), .X(n67130) );
  inv_x4_sg U55062 ( .A(n22508), .X(n67132) );
  inv_x4_sg U55063 ( .A(n22506), .X(n67134) );
  inv_x4_sg U55064 ( .A(n22491), .X(n67317) );
  inv_x4_sg U55065 ( .A(n22488), .X(n67320) );
  inv_x4_sg U55066 ( .A(n22487), .X(n67321) );
  inv_x4_sg U55067 ( .A(n22486), .X(n67322) );
  inv_x4_sg U55068 ( .A(n22484), .X(n67324) );
  inv_x4_sg U55069 ( .A(n22482), .X(n67326) );
  inv_x4_sg U55070 ( .A(n22480), .X(n67328) );
  inv_x4_sg U55071 ( .A(n22478), .X(n67330) );
  inv_x4_sg U55072 ( .A(n22477), .X(n67331) );
  inv_x4_sg U55073 ( .A(n22476), .X(n67332) );
  inv_x4_sg U55074 ( .A(n22465), .X(n67103) );
  inv_x4_sg U55075 ( .A(n22464), .X(n67104) );
  inv_x4_sg U55076 ( .A(n22461), .X(n67107) );
  inv_x4_sg U55077 ( .A(n22460), .X(n67108) );
  inv_x4_sg U55078 ( .A(n22459), .X(n67109) );
  inv_x4_sg U55079 ( .A(n22457), .X(n67111) );
  inv_x4_sg U55080 ( .A(n22455), .X(n67113) );
  inv_x4_sg U55081 ( .A(n22453), .X(n67115) );
  inv_x4_sg U55082 ( .A(n22451), .X(n67117) );
  inv_x4_sg U55083 ( .A(n22450), .X(n67118) );
  inv_x4_sg U55084 ( .A(n22449), .X(n67119) );
  inv_x4_sg U55085 ( .A(n22437), .X(n61897) );
  inv_x4_sg U55086 ( .A(n22433), .X(n61893) );
  inv_x4_sg U55087 ( .A(n22431), .X(n61891) );
  inv_x4_sg U55088 ( .A(n22429), .X(n61889) );
  inv_x4_sg U55089 ( .A(n22416), .X(n61881) );
  inv_x4_sg U55090 ( .A(n22412), .X(n61877) );
  inv_x4_sg U55091 ( .A(n22408), .X(n61873) );
  inv_x4_sg U55092 ( .A(n22406), .X(n61871) );
  inv_x4_sg U55093 ( .A(n22404), .X(n61869) );
  nor_x2_sg U55094 ( .A(n67097), .B(n68574), .X(n22417) );
  nor_x4_sg U55095 ( .A(n22746), .B(n57862), .X(n22974) );
  inv_x2_sg U55096 ( .A(n47574), .X(n47575) );
  inv_x2_sg U55097 ( .A(n47576), .X(n47577) );
  inv_x2_sg U55098 ( .A(n47578), .X(n47579) );
  inv_x2_sg U55099 ( .A(n47580), .X(n47581) );
  inv_x2_sg U55100 ( .A(n47582), .X(n47583) );
  inv_x2_sg U55101 ( .A(n47584), .X(n47585) );
  inv_x2_sg U55102 ( .A(n47586), .X(n47587) );
  inv_x2_sg U55103 ( .A(n47588), .X(n47589) );
  inv_x2_sg U55104 ( .A(n47590), .X(n47591) );
  inv_x2_sg U55105 ( .A(n47592), .X(n47593) );
  inv_x2_sg U55106 ( .A(n47594), .X(n47595) );
  inv_x2_sg U55107 ( .A(n47596), .X(n47597) );
  inv_x2_sg U55108 ( .A(n47598), .X(n47599) );
  inv_x4_sg U55109 ( .A(n22640), .X(n67379) );
  inv_x4_sg U55110 ( .A(n22639), .X(n67380) );
  inv_x4_sg U55111 ( .A(n22613), .X(n67166) );
  inv_x4_sg U55112 ( .A(n22612), .X(n67167) );
  nor_x4_sg U55113 ( .A(n67534), .B(n57091), .X(n26095) );
  inv_x4_sg U55114 ( .A(n23304), .X(n67099) );
  nor_x8_sg U55115 ( .A(n26303), .B(n26304), .X(n26122) );
  nand_x8_sg U55116 ( .A(n57308), .B(n57310), .X(n26304) );
  inv_x4_sg U55117 ( .A(n68268), .X(n61909) );
  nor_x4_sg U55118 ( .A(n31952), .B(n32063), .X(n31978) );
  nand_x8_sg U55119 ( .A(n32072), .B(n32073), .X(n31952) );
  nand_x4_sg U55120 ( .A(n32064), .B(n32065), .X(n32063) );
  inv_x4_sg U55121 ( .A(n47600), .X(n47601) );
  inv_x4_sg U55122 ( .A(n47602), .X(n47603) );
  inv_x4_sg U55123 ( .A(n47604), .X(n47605) );
  inv_x4_sg U55124 ( .A(n47606), .X(n47607) );
  inv_x4_sg U55125 ( .A(n47608), .X(n47609) );
  inv_x4_sg U55126 ( .A(n47610), .X(n47611) );
  inv_x4_sg U55127 ( .A(n47612), .X(n47613) );
  inv_x4_sg U55128 ( .A(n46893), .X(n47614) );
  inv_x8_sg U55129 ( .A(n47614), .X(n47615) );
  inv_x4_sg U55130 ( .A(n47615), .X(n61911) );
  inv_x4_sg U55131 ( .A(n47616), .X(n47617) );
  inv_x4_sg U55132 ( .A(n47618), .X(n47619) );
  inv_x4_sg U55133 ( .A(n47620), .X(n47621) );
  inv_x4_sg U55134 ( .A(n47622), .X(n47623) );
  inv_x4_sg U55135 ( .A(n47624), .X(n47625) );
  inv_x4_sg U55136 ( .A(n47626), .X(n47627) );
  inv_x4_sg U55137 ( .A(n47628), .X(n47629) );
  inv_x4_sg U55138 ( .A(n47630), .X(n47631) );
  inv_x4_sg U55139 ( .A(n47632), .X(n47633) );
  inv_x4_sg U55140 ( .A(n47634), .X(n47635) );
  inv_x4_sg U55141 ( .A(n47636), .X(n47637) );
  inv_x4_sg U55142 ( .A(n47638), .X(n47639) );
  inv_x4_sg U55143 ( .A(n47640), .X(n47641) );
  inv_x4_sg U55144 ( .A(n47642), .X(n47643) );
  inv_x4_sg U55145 ( .A(n47644), .X(n47645) );
  inv_x4_sg U55146 ( .A(n47646), .X(n47647) );
  inv_x4_sg U55147 ( .A(n47648), .X(n47649) );
  inv_x4_sg U55148 ( .A(n47650), .X(n47651) );
  inv_x4_sg U55149 ( .A(n47652), .X(n47653) );
  inv_x4_sg U55150 ( .A(n47654), .X(n47655) );
  inv_x4_sg U55151 ( .A(n47656), .X(n47657) );
  inv_x4_sg U55152 ( .A(n47658), .X(n47659) );
  inv_x4_sg U55153 ( .A(n47660), .X(n47661) );
  inv_x4_sg U55154 ( .A(n47662), .X(n47663) );
  inv_x4_sg U55155 ( .A(n47664), .X(n47665) );
  inv_x4_sg U55156 ( .A(n47666), .X(n47667) );
  inv_x4_sg U55157 ( .A(n47668), .X(n47669) );
  inv_x4_sg U55158 ( .A(n47670), .X(n47671) );
  inv_x4_sg U55159 ( .A(n47672), .X(n47673) );
  inv_x4_sg U55160 ( .A(n47674), .X(n47675) );
  inv_x4_sg U55161 ( .A(n47676), .X(n47677) );
  inv_x4_sg U55162 ( .A(n47678), .X(n47679) );
  inv_x4_sg U55163 ( .A(n47680), .X(n47681) );
  inv_x4_sg U55164 ( .A(n47682), .X(n47683) );
  inv_x4_sg U55165 ( .A(n47684), .X(n47685) );
  inv_x4_sg U55166 ( .A(n47686), .X(n47687) );
  inv_x4_sg U55167 ( .A(n47688), .X(n47689) );
  inv_x4_sg U55168 ( .A(n47690), .X(n47691) );
  inv_x4_sg U55169 ( .A(n47692), .X(n47693) );
  inv_x4_sg U55170 ( .A(n47694), .X(n47695) );
  inv_x4_sg U55171 ( .A(n47696), .X(n47697) );
  inv_x4_sg U55172 ( .A(n47698), .X(n47699) );
  inv_x4_sg U55173 ( .A(n47700), .X(n47701) );
  inv_x4_sg U55174 ( .A(n47702), .X(n47703) );
  inv_x4_sg U55175 ( .A(n47704), .X(n47705) );
  inv_x4_sg U55176 ( .A(n47706), .X(n47707) );
  inv_x4_sg U55177 ( .A(n47708), .X(n47709) );
  inv_x4_sg U55178 ( .A(n47710), .X(n47711) );
  inv_x4_sg U55179 ( .A(n47712), .X(n47713) );
  inv_x4_sg U55180 ( .A(n47714), .X(n47715) );
  inv_x4_sg U55181 ( .A(n47716), .X(n47717) );
  inv_x4_sg U55182 ( .A(n47718), .X(n47719) );
  inv_x4_sg U55183 ( .A(n47720), .X(n47721) );
  inv_x4_sg U55184 ( .A(n47722), .X(n47723) );
  inv_x4_sg U55185 ( .A(n47724), .X(n47725) );
  inv_x4_sg U55186 ( .A(n47726), .X(n47727) );
  inv_x4_sg U55187 ( .A(n47728), .X(n47729) );
  inv_x4_sg U55188 ( .A(n47730), .X(n47731) );
  inv_x4_sg U55189 ( .A(n47732), .X(n47733) );
  inv_x4_sg U55190 ( .A(n47734), .X(n47735) );
  inv_x4_sg U55191 ( .A(n47736), .X(n47737) );
  inv_x4_sg U55192 ( .A(n47738), .X(n47739) );
  inv_x4_sg U55193 ( .A(n47285), .X(n47740) );
  inv_x8_sg U55194 ( .A(n47740), .X(state[0]) );
  inv_x4_sg U55195 ( .A(n46977), .X(n47742) );
  inv_x8_sg U55196 ( .A(n47742), .X(n47743) );
  inv_x4_sg U55197 ( .A(n46975), .X(n47744) );
  inv_x8_sg U55198 ( .A(n47744), .X(n47745) );
  inv_x4_sg U55199 ( .A(n46967), .X(n47746) );
  inv_x8_sg U55200 ( .A(n47746), .X(n47747) );
  inv_x4_sg U55201 ( .A(n47121), .X(n47748) );
  inv_x8_sg U55202 ( .A(n47748), .X(n47749) );
  inv_x4_sg U55203 ( .A(n47119), .X(n47750) );
  inv_x8_sg U55204 ( .A(n47750), .X(n47751) );
  inv_x4_sg U55205 ( .A(n47111), .X(n47752) );
  inv_x8_sg U55206 ( .A(n47752), .X(n47753) );
  inv_x4_sg U55207 ( .A(n47093), .X(n47754) );
  inv_x8_sg U55208 ( .A(n47754), .X(n47755) );
  inv_x4_sg U55209 ( .A(n46949), .X(n47756) );
  inv_x8_sg U55210 ( .A(n47756), .X(n47757) );
  inv_x4_sg U55211 ( .A(n47045), .X(n47758) );
  inv_x8_sg U55212 ( .A(n47758), .X(n47759) );
  inv_x4_sg U55213 ( .A(n47161), .X(n47760) );
  inv_x8_sg U55214 ( .A(n47760), .X(n47761) );
  inv_x4_sg U55215 ( .A(n47159), .X(n47762) );
  inv_x8_sg U55216 ( .A(n47762), .X(n47763) );
  inv_x4_sg U55217 ( .A(n47151), .X(n47764) );
  inv_x8_sg U55218 ( .A(n47764), .X(n47765) );
  inv_x4_sg U55219 ( .A(n47017), .X(n47766) );
  inv_x8_sg U55220 ( .A(n47766), .X(n47767) );
  inv_x4_sg U55221 ( .A(n47015), .X(n47768) );
  inv_x8_sg U55222 ( .A(n47768), .X(n47769) );
  inv_x4_sg U55223 ( .A(n47007), .X(n47770) );
  inv_x8_sg U55224 ( .A(n47770), .X(n47771) );
  inv_x4_sg U55225 ( .A(n46931), .X(n47772) );
  inv_x8_sg U55226 ( .A(n47772), .X(n47773) );
  inv_x4_sg U55227 ( .A(n46937), .X(n47774) );
  inv_x8_sg U55228 ( .A(n47774), .X(n47775) );
  inv_x8_sg U55229 ( .A(n47775), .X(n68574) );
  inv_x2_sg U55230 ( .A(n57083), .X(n58496) );
  inv_x2_sg U55231 ( .A(n57077), .X(n58506) );
  inv_x2_sg U55232 ( .A(n57073), .X(n58527) );
  inv_x2_sg U55233 ( .A(n57087), .X(n58545) );
  inv_x2_sg U55234 ( .A(n57079), .X(n58555) );
  nand_x2_sg U55235 ( .A(n67096), .B(n57104), .X(n23807) );
  nand_x2_sg U55236 ( .A(n47493), .B(n57862), .X(n23135) );
  nand_x2_sg U55237 ( .A(n47495), .B(n57862), .X(n22908) );
  nand_x4_sg U55238 ( .A(n25574), .B(n25575), .X(n24081) );
  nand_x4_sg U55239 ( .A(n25152), .B(n25153), .X(n24001) );
  nand_x4_sg U55240 ( .A(n24972), .B(n24973), .X(n23971) );
  nand_x4_sg U55241 ( .A(n25995), .B(n25996), .X(n24151) );
  nand_x4_sg U55242 ( .A(n25393), .B(n25394), .X(n24041) );
  nand_x2_sg U55243 ( .A(n68373), .B(n26297), .X(n26261) );
  nand_x2_sg U55244 ( .A(n57069), .B(n26263), .X(n26262) );
  nor_x2_sg U55245 ( .A(n24829), .B(n68405), .X(n25940) );
  inv_x4_sg U55246 ( .A(n55035), .X(n68405) );
  nor_x2_sg U55247 ( .A(n68412), .B(n57102), .X(n25791) );
  inv_x4_sg U55248 ( .A(n55293), .X(n68412) );
  nor_x2_sg U55249 ( .A(n24829), .B(n68403), .X(n25790) );
  inv_x4_sg U55250 ( .A(n55031), .X(n68403) );
  nor_x2_sg U55251 ( .A(n68410), .B(n57102), .X(n25671) );
  inv_x4_sg U55252 ( .A(n55289), .X(n68410) );
  nor_x2_sg U55253 ( .A(n24829), .B(n68401), .X(n25670) );
  inv_x4_sg U55254 ( .A(n55027), .X(n68401) );
  nor_x2_sg U55255 ( .A(n68408), .B(n57102), .X(n25521) );
  inv_x4_sg U55256 ( .A(n55285), .X(n68408) );
  nor_x2_sg U55257 ( .A(n24829), .B(n68399), .X(n25520) );
  inv_x4_sg U55258 ( .A(n55023), .X(n68399) );
  nor_x2_sg U55259 ( .A(n24829), .B(n68494), .X(n25338) );
  inv_x4_sg U55260 ( .A(n55055), .X(n68494) );
  nor_x2_sg U55261 ( .A(n68501), .B(n57102), .X(n25189) );
  inv_x4_sg U55262 ( .A(n55305), .X(n68501) );
  nor_x2_sg U55263 ( .A(n24829), .B(n68492), .X(n25188) );
  inv_x4_sg U55264 ( .A(n55051), .X(n68492) );
  nor_x2_sg U55265 ( .A(n68499), .B(n57102), .X(n25069) );
  inv_x4_sg U55266 ( .A(n55301), .X(n68499) );
  nor_x2_sg U55267 ( .A(n24829), .B(n68490), .X(n25068) );
  inv_x4_sg U55268 ( .A(n55047), .X(n68490) );
  nor_x2_sg U55269 ( .A(n24829), .B(n68488), .X(n24918) );
  inv_x4_sg U55270 ( .A(n55043), .X(n68488) );
  nor_x2_sg U55271 ( .A(n68497), .B(n57102), .X(n24919) );
  inv_x4_sg U55272 ( .A(n55297), .X(n68497) );
  inv_x4_sg U55273 ( .A(n57007), .X(n68482) );
  inv_x4_sg U55274 ( .A(n56975), .X(n68486) );
  inv_x4_sg U55275 ( .A(n56995), .X(n68586) );
  nor_x2_sg U55276 ( .A(n68414), .B(n57102), .X(n25941) );
  inv_x4_sg U55277 ( .A(n55309), .X(n68414) );
  nor_x2_sg U55278 ( .A(n68503), .B(n57102), .X(n25339) );
  inv_x4_sg U55279 ( .A(n55313), .X(n68503) );
  inv_x4_sg U55280 ( .A(n56977), .X(n68484) );
  inv_x4_sg U55281 ( .A(n57003), .X(n68584) );
  inv_x4_sg U55282 ( .A(n57011), .X(n68582) );
  nor_x2_sg U55283 ( .A(n68433), .B(n58638), .X(n58142) );
  inv_x4_sg U55284 ( .A(n55041), .X(n68433) );
  nor_x2_sg U55285 ( .A(n68523), .B(n57104), .X(n58242) );
  inv_x4_sg U55286 ( .A(n55061), .X(n68523) );
  inv_x2_sg U55287 ( .A(\mask_0/reg_ii_mask [0]), .X(n55156) );
  inv_x2_sg U55288 ( .A(\mask_0/reg_ii_mask [4]), .X(n55158) );
  inv_x2_sg U55289 ( .A(\mask_0/reg_ii_mask [5]), .X(n55160) );
  inv_x2_sg U55290 ( .A(\mask_0/reg_ii_mask [17]), .X(n55162) );
  inv_x2_sg U55291 ( .A(\mask_0/reg_ii_mask [28]), .X(n55164) );
  inv_x2_sg U55292 ( .A(\mask_0/reg_ii_mask [29]), .X(n55166) );
  inv_x2_sg U55293 ( .A(\mask_0/reg_ii_mask [30]), .X(n55168) );
  inv_x2_sg U55294 ( .A(\mask_0/reg_ii_mask [31]), .X(n55170) );
  inv_x2_sg U55295 ( .A(\mask_0/reg_ww_mask [1]), .X(n55172) );
  inv_x2_sg U55296 ( .A(\mask_0/reg_ww_mask [2]), .X(n55174) );
  inv_x2_sg U55297 ( .A(\mask_0/reg_ww_mask [3]), .X(n55176) );
  inv_x2_sg U55298 ( .A(\mask_0/reg_ww_mask [6]), .X(n55178) );
  inv_x2_sg U55299 ( .A(\mask_0/reg_ww_mask [7]), .X(n55180) );
  inv_x2_sg U55300 ( .A(\mask_0/reg_ww_mask [8]), .X(n55182) );
  inv_x2_sg U55301 ( .A(\mask_0/reg_ww_mask [9]), .X(n55184) );
  inv_x2_sg U55302 ( .A(\mask_0/reg_ww_mask [10]), .X(n55186) );
  inv_x2_sg U55303 ( .A(\mask_0/reg_ww_mask [11]), .X(n55188) );
  inv_x2_sg U55304 ( .A(\mask_0/reg_ww_mask [12]), .X(n55190) );
  inv_x2_sg U55305 ( .A(\mask_0/reg_ww_mask [13]), .X(n55192) );
  inv_x2_sg U55306 ( .A(\mask_0/reg_ww_mask [14]), .X(n55194) );
  inv_x2_sg U55307 ( .A(\mask_0/reg_ww_mask [15]), .X(n55196) );
  inv_x2_sg U55308 ( .A(\mask_0/reg_ww_mask [16]), .X(n55198) );
  inv_x2_sg U55309 ( .A(\mask_0/reg_ww_mask [18]), .X(n55200) );
  inv_x2_sg U55310 ( .A(\mask_0/reg_ww_mask [19]), .X(n55202) );
  inv_x2_sg U55311 ( .A(\mask_0/reg_ww_mask [20]), .X(n55204) );
  inv_x2_sg U55312 ( .A(\mask_0/reg_ww_mask [21]), .X(n55206) );
  inv_x2_sg U55313 ( .A(\mask_0/reg_ww_mask [22]), .X(n55208) );
  inv_x2_sg U55314 ( .A(\mask_0/reg_ww_mask [23]), .X(n55210) );
  inv_x2_sg U55315 ( .A(\mask_0/reg_ww_mask [24]), .X(n55212) );
  inv_x2_sg U55316 ( .A(\mask_0/reg_ww_mask [25]), .X(n55214) );
  inv_x2_sg U55317 ( .A(\mask_0/reg_ww_mask [26]), .X(n55216) );
  inv_x2_sg U55318 ( .A(\mask_0/reg_ww_mask [27]), .X(n55218) );
  inv_x2_sg U55319 ( .A(\filter_0/reg_xor_i_mask [2]), .X(n55062) );
  inv_x2_sg U55320 ( .A(\filter_0/reg_xor_i_mask [18]), .X(n55064) );
  inv_x2_sg U55321 ( .A(\filter_0/reg_xor_w_mask [2]), .X(n55066) );
  inv_x2_sg U55322 ( .A(\filter_0/reg_xor_w_mask [18]), .X(n55068) );
  inv_x2_sg U55323 ( .A(n55255), .X(n67487) );
  inv_x2_sg U55324 ( .A(n55269), .X(n67489) );
  inv_x2_sg U55325 ( .A(n55267), .X(n67491) );
  inv_x2_sg U55326 ( .A(n55253), .X(n67492) );
  inv_x2_sg U55327 ( .A(n55265), .X(n67493) );
  inv_x2_sg U55328 ( .A(n55263), .X(n67494) );
  inv_x2_sg U55329 ( .A(n55261), .X(n67496) );
  inv_x2_sg U55330 ( .A(n55259), .X(n67294) );
  inv_x2_sg U55331 ( .A(n55281), .X(n67296) );
  inv_x2_sg U55332 ( .A(n55279), .X(n67298) );
  inv_x2_sg U55333 ( .A(n55257), .X(n67299) );
  inv_x2_sg U55334 ( .A(n55277), .X(n67300) );
  inv_x2_sg U55335 ( .A(n55275), .X(n67301) );
  inv_x2_sg U55336 ( .A(n55273), .X(n67303) );
  nor_x1_sg U55337 ( .A(n24485), .B(n46887), .X(n58131) );
  inv_x8_sg U55338 ( .A(n23308), .X(n67096) );
  inv_x4_sg U55339 ( .A(n25900), .X(n67458) );
  inv_x4_sg U55340 ( .A(n25298), .X(n67265) );
  inv_x4_sg U55341 ( .A(n24848), .X(n67280) );
  inv_x4_sg U55342 ( .A(n23412), .X(n67502) );
  nor_x4_sg U55343 ( .A(n57920), .B(n57951), .X(n58388) );
  nand_x2_sg U55344 ( .A(n58478), .B(n57100), .X(n58390) );
  nor_x4_sg U55345 ( .A(n68227), .B(n57527), .X(n38414) );
  inv_x4_sg U55346 ( .A(n22441), .X(n61901) );
  inv_x4_sg U55347 ( .A(n22588), .X(n67359) );
  inv_x4_sg U55348 ( .A(n22578), .X(n67369) );
  inv_x4_sg U55349 ( .A(n22574), .X(n67373) );
  inv_x4_sg U55350 ( .A(n22573), .X(n67374) );
  inv_x4_sg U55351 ( .A(n22562), .X(n67146) );
  inv_x4_sg U55352 ( .A(n22552), .X(n67156) );
  inv_x4_sg U55353 ( .A(n22547), .X(n67161) );
  inv_x4_sg U55354 ( .A(n22492), .X(n67316) );
  inv_x4_sg U55355 ( .A(n22543), .X(n67335) );
  inv_x4_sg U55356 ( .A(n22537), .X(n67341) );
  inv_x4_sg U55357 ( .A(n22528), .X(n67350) );
  inv_x4_sg U55358 ( .A(n22512), .X(n67128) );
  inv_x4_sg U55359 ( .A(n22503), .X(n67137) );
  inv_x4_sg U55360 ( .A(n22500), .X(n67140) );
  inv_x4_sg U55361 ( .A(n22490), .X(n67318) );
  inv_x4_sg U55362 ( .A(n22489), .X(n67319) );
  inv_x4_sg U55363 ( .A(n22485), .X(n67323) );
  inv_x4_sg U55364 ( .A(n22483), .X(n67325) );
  inv_x4_sg U55365 ( .A(n22481), .X(n67327) );
  inv_x4_sg U55366 ( .A(n22479), .X(n67329) );
  inv_x4_sg U55367 ( .A(n22475), .X(n67333) );
  inv_x4_sg U55368 ( .A(n22474), .X(n67334) );
  inv_x4_sg U55369 ( .A(n22466), .X(n67102) );
  inv_x4_sg U55370 ( .A(n22463), .X(n67105) );
  inv_x4_sg U55371 ( .A(n22462), .X(n67106) );
  inv_x4_sg U55372 ( .A(n22458), .X(n67110) );
  inv_x4_sg U55373 ( .A(n22456), .X(n67112) );
  inv_x4_sg U55374 ( .A(n22454), .X(n67114) );
  inv_x4_sg U55375 ( .A(n22452), .X(n67116) );
  inv_x4_sg U55376 ( .A(n22447), .X(n67121) );
  inv_x4_sg U55377 ( .A(n22435), .X(n61895) );
  inv_x4_sg U55378 ( .A(n22426), .X(n61886) );
  inv_x4_sg U55379 ( .A(n22415), .X(n61880) );
  inv_x4_sg U55380 ( .A(n22410), .X(n61875) );
  inv_x4_sg U55381 ( .A(n22401), .X(n61866) );
  inv_x4_sg U55382 ( .A(n22398), .X(n61863) );
  inv_x2_sg U55383 ( .A(n47776), .X(n47777) );
  inv_x2_sg U55384 ( .A(n47778), .X(n47779) );
  inv_x2_sg U55385 ( .A(n47780), .X(n47781) );
  inv_x2_sg U55386 ( .A(n47782), .X(n47783) );
  inv_x2_sg U55387 ( .A(n47784), .X(n47785) );
  inv_x2_sg U55388 ( .A(n47786), .X(n47787) );
  inv_x2_sg U55389 ( .A(n47788), .X(n47789) );
  inv_x2_sg U55390 ( .A(n47790), .X(n47791) );
  inv_x2_sg U55391 ( .A(n47792), .X(n47793) );
  inv_x2_sg U55392 ( .A(n47794), .X(n47795) );
  inv_x2_sg U55393 ( .A(n47796), .X(n47797) );
  inv_x2_sg U55394 ( .A(n47798), .X(n47799) );
  inv_x2_sg U55395 ( .A(n47800), .X(n47801) );
  inv_x2_sg U55396 ( .A(n47802), .X(n47803) );
  inv_x2_sg U55397 ( .A(n47804), .X(n47805) );
  inv_x2_sg U55398 ( .A(n47806), .X(n47807) );
  inv_x2_sg U55399 ( .A(n47808), .X(n47809) );
  inv_x2_sg U55400 ( .A(n47810), .X(n47811) );
  inv_x2_sg U55401 ( .A(n47812), .X(n47813) );
  inv_x2_sg U55402 ( .A(n47814), .X(n47815) );
  inv_x2_sg U55403 ( .A(n47816), .X(n47817) );
  inv_x2_sg U55404 ( .A(n47818), .X(n47819) );
  inv_x2_sg U55405 ( .A(n47820), .X(n47821) );
  inv_x2_sg U55406 ( .A(n47822), .X(n47823) );
  inv_x2_sg U55407 ( .A(n47824), .X(n47825) );
  inv_x2_sg U55408 ( .A(n47826), .X(n47827) );
  inv_x2_sg U55409 ( .A(n47828), .X(n47829) );
  inv_x2_sg U55410 ( .A(n47830), .X(n47831) );
  inv_x2_sg U55411 ( .A(n47832), .X(n47833) );
  inv_x2_sg U55412 ( .A(n47834), .X(n47835) );
  inv_x2_sg U55413 ( .A(n47836), .X(n47837) );
  inv_x2_sg U55414 ( .A(n47838), .X(n47839) );
  inv_x2_sg U55415 ( .A(n47840), .X(n47841) );
  inv_x2_sg U55416 ( .A(n47842), .X(n47843) );
  inv_x2_sg U55417 ( .A(n47844), .X(n47845) );
  inv_x2_sg U55418 ( .A(n47846), .X(n47847) );
  inv_x2_sg U55419 ( .A(n47848), .X(n47849) );
  inv_x2_sg U55420 ( .A(n47850), .X(n47851) );
  inv_x2_sg U55421 ( .A(n47852), .X(n47853) );
  inv_x2_sg U55422 ( .A(n47854), .X(n47855) );
  inv_x2_sg U55423 ( .A(n47856), .X(n47857) );
  inv_x2_sg U55424 ( .A(n47858), .X(n47859) );
  inv_x2_sg U55425 ( .A(n47860), .X(n47861) );
  inv_x2_sg U55426 ( .A(n47862), .X(n47863) );
  inv_x2_sg U55427 ( .A(n47864), .X(n47865) );
  inv_x2_sg U55428 ( .A(n47866), .X(n47867) );
  inv_x2_sg U55429 ( .A(n47868), .X(n47869) );
  inv_x2_sg U55430 ( .A(n47870), .X(n47871) );
  inv_x2_sg U55431 ( .A(n47872), .X(n47873) );
  inv_x2_sg U55432 ( .A(n47874), .X(n47875) );
  inv_x2_sg U55433 ( .A(n47876), .X(n47877) );
  inv_x2_sg U55434 ( .A(n47878), .X(n47879) );
  inv_x2_sg U55435 ( .A(n47880), .X(n47881) );
  inv_x2_sg U55436 ( .A(n47882), .X(n47883) );
  inv_x2_sg U55437 ( .A(n47884), .X(n47885) );
  inv_x2_sg U55438 ( .A(n47886), .X(n47887) );
  inv_x2_sg U55439 ( .A(n47888), .X(n47889) );
  inv_x2_sg U55440 ( .A(n47890), .X(n47891) );
  inv_x2_sg U55441 ( .A(n47892), .X(n47893) );
  inv_x2_sg U55442 ( .A(n47894), .X(n47895) );
  inv_x2_sg U55443 ( .A(n47896), .X(n47897) );
  inv_x2_sg U55444 ( .A(n47898), .X(n47899) );
  inv_x2_sg U55445 ( .A(n47900), .X(n47901) );
  inv_x2_sg U55446 ( .A(n47902), .X(n47903) );
  inv_x2_sg U55447 ( .A(n47904), .X(n47905) );
  inv_x2_sg U55448 ( .A(n47906), .X(n47907) );
  inv_x2_sg U55449 ( .A(n47908), .X(n47909) );
  inv_x2_sg U55450 ( .A(n47910), .X(n47911) );
  inv_x2_sg U55451 ( .A(n47912), .X(n47913) );
  inv_x2_sg U55452 ( .A(n47914), .X(n47915) );
  inv_x2_sg U55453 ( .A(n47916), .X(n47917) );
  inv_x2_sg U55454 ( .A(n47918), .X(n47919) );
  inv_x2_sg U55455 ( .A(n47920), .X(n47921) );
  inv_x2_sg U55456 ( .A(n47922), .X(n47923) );
  inv_x2_sg U55457 ( .A(n47924), .X(n47925) );
  inv_x2_sg U55458 ( .A(n47926), .X(n47927) );
  inv_x2_sg U55459 ( .A(n47928), .X(n47929) );
  inv_x2_sg U55460 ( .A(n47930), .X(n47931) );
  inv_x2_sg U55461 ( .A(n47932), .X(n47933) );
  inv_x2_sg U55462 ( .A(n47934), .X(n47935) );
  inv_x2_sg U55463 ( .A(n47936), .X(n47937) );
  inv_x2_sg U55464 ( .A(n47938), .X(n47939) );
  inv_x2_sg U55465 ( .A(n47940), .X(n47941) );
  inv_x2_sg U55466 ( .A(n47942), .X(n47943) );
  inv_x2_sg U55467 ( .A(n47944), .X(n47945) );
  inv_x2_sg U55468 ( .A(n47946), .X(n47947) );
  inv_x2_sg U55469 ( .A(n47948), .X(n47949) );
  inv_x2_sg U55470 ( .A(n47950), .X(n47951) );
  inv_x2_sg U55471 ( .A(n47952), .X(n47953) );
  inv_x2_sg U55472 ( .A(n47954), .X(n47955) );
  inv_x2_sg U55473 ( .A(n47956), .X(n47957) );
  inv_x2_sg U55474 ( .A(n47958), .X(n47959) );
  inv_x2_sg U55475 ( .A(n47960), .X(n47961) );
  inv_x2_sg U55476 ( .A(n47962), .X(n47963) );
  inv_x2_sg U55477 ( .A(n47964), .X(n47965) );
  inv_x2_sg U55478 ( .A(n47966), .X(n47967) );
  inv_x2_sg U55479 ( .A(n47968), .X(n47969) );
  inv_x2_sg U55480 ( .A(n47970), .X(n47971) );
  inv_x2_sg U55481 ( .A(n47972), .X(n47973) );
  inv_x2_sg U55482 ( .A(n47974), .X(n47975) );
  inv_x2_sg U55483 ( .A(n47976), .X(n47977) );
  inv_x2_sg U55484 ( .A(n47978), .X(n47979) );
  inv_x2_sg U55485 ( .A(n47980), .X(n47981) );
  inv_x2_sg U55486 ( .A(n47982), .X(n47983) );
  inv_x2_sg U55487 ( .A(n47984), .X(n47985) );
  inv_x2_sg U55488 ( .A(n47986), .X(n47987) );
  inv_x2_sg U55489 ( .A(n47988), .X(n47989) );
  inv_x2_sg U55490 ( .A(n47990), .X(n47991) );
  inv_x2_sg U55491 ( .A(n47992), .X(n47993) );
  inv_x2_sg U55492 ( .A(n47994), .X(n47995) );
  inv_x2_sg U55493 ( .A(n47996), .X(n47997) );
  inv_x2_sg U55494 ( .A(n47998), .X(n47999) );
  inv_x2_sg U55495 ( .A(n48000), .X(n48001) );
  inv_x2_sg U55496 ( .A(n48002), .X(n48003) );
  inv_x2_sg U55497 ( .A(n48004), .X(n48005) );
  inv_x2_sg U55498 ( .A(n48006), .X(n48007) );
  inv_x2_sg U55499 ( .A(n48008), .X(n48009) );
  inv_x2_sg U55500 ( .A(n48010), .X(n48011) );
  inv_x2_sg U55501 ( .A(n48012), .X(n48013) );
  inv_x2_sg U55502 ( .A(n48014), .X(n48015) );
  inv_x2_sg U55503 ( .A(n48016), .X(n48017) );
  inv_x2_sg U55504 ( .A(n48018), .X(n48019) );
  inv_x2_sg U55505 ( .A(n48020), .X(n48021) );
  inv_x2_sg U55506 ( .A(n48022), .X(n48023) );
  inv_x2_sg U55507 ( .A(n48024), .X(n48025) );
  inv_x2_sg U55508 ( .A(n48026), .X(n48027) );
  inv_x2_sg U55509 ( .A(n48028), .X(n48029) );
  inv_x2_sg U55510 ( .A(n48030), .X(n48031) );
  inv_x2_sg U55511 ( .A(n48032), .X(n48033) );
  inv_x2_sg U55512 ( .A(n48034), .X(n48035) );
  inv_x2_sg U55513 ( .A(n48036), .X(n48037) );
  inv_x2_sg U55514 ( .A(n48038), .X(n48039) );
  inv_x2_sg U55515 ( .A(n48040), .X(n48041) );
  inv_x2_sg U55516 ( .A(n48042), .X(n48043) );
  inv_x2_sg U55517 ( .A(n48044), .X(n48045) );
  inv_x2_sg U55518 ( .A(n48046), .X(n48047) );
  inv_x2_sg U55519 ( .A(n48048), .X(n48049) );
  inv_x2_sg U55520 ( .A(n48050), .X(n48051) );
  inv_x2_sg U55521 ( .A(n48052), .X(n48053) );
  inv_x2_sg U55522 ( .A(n48054), .X(n48055) );
  inv_x2_sg U55523 ( .A(n48056), .X(n48057) );
  inv_x2_sg U55524 ( .A(n48058), .X(n48059) );
  inv_x2_sg U55525 ( .A(n48060), .X(n48061) );
  inv_x2_sg U55526 ( .A(n48062), .X(n48063) );
  inv_x2_sg U55527 ( .A(n48064), .X(n48065) );
  inv_x2_sg U55528 ( .A(n48066), .X(n48067) );
  inv_x2_sg U55529 ( .A(n48068), .X(n48069) );
  inv_x2_sg U55530 ( .A(n48070), .X(n48071) );
  inv_x2_sg U55531 ( .A(n48072), .X(n48073) );
  inv_x2_sg U55532 ( .A(n48074), .X(n48075) );
  inv_x2_sg U55533 ( .A(n48076), .X(n48077) );
  inv_x2_sg U55534 ( .A(n48078), .X(n48079) );
  inv_x2_sg U55535 ( .A(n48080), .X(n48081) );
  inv_x2_sg U55536 ( .A(n48082), .X(n48083) );
  inv_x2_sg U55537 ( .A(n48084), .X(n48085) );
  inv_x2_sg U55538 ( .A(n48086), .X(n48087) );
  inv_x2_sg U55539 ( .A(n48088), .X(n48089) );
  inv_x2_sg U55540 ( .A(n48090), .X(n48091) );
  inv_x2_sg U55541 ( .A(n48092), .X(n48093) );
  inv_x2_sg U55542 ( .A(n48094), .X(n48095) );
  inv_x2_sg U55543 ( .A(n48096), .X(n48097) );
  inv_x2_sg U55544 ( .A(n48098), .X(n48099) );
  inv_x2_sg U55545 ( .A(n48100), .X(n48101) );
  inv_x2_sg U55546 ( .A(n48102), .X(n48103) );
  inv_x2_sg U55547 ( .A(n48104), .X(n48105) );
  inv_x2_sg U55548 ( .A(n48106), .X(n48107) );
  inv_x2_sg U55549 ( .A(n48108), .X(n48109) );
  inv_x2_sg U55550 ( .A(n48110), .X(n48111) );
  inv_x2_sg U55551 ( .A(n48112), .X(n48113) );
  inv_x2_sg U55552 ( .A(n48114), .X(n48115) );
  inv_x2_sg U55553 ( .A(n48116), .X(n48117) );
  inv_x2_sg U55554 ( .A(n48118), .X(n48119) );
  inv_x2_sg U55555 ( .A(n48120), .X(n48121) );
  inv_x2_sg U55556 ( .A(n48122), .X(n48123) );
  inv_x2_sg U55557 ( .A(n48124), .X(n48125) );
  inv_x2_sg U55558 ( .A(n48126), .X(n48127) );
  inv_x2_sg U55559 ( .A(n48128), .X(n48129) );
  inv_x2_sg U55560 ( .A(n48130), .X(n48131) );
  inv_x2_sg U55561 ( .A(n48132), .X(n48133) );
  inv_x2_sg U55562 ( .A(n48134), .X(n48135) );
  inv_x2_sg U55563 ( .A(n48136), .X(n48137) );
  inv_x2_sg U55564 ( .A(n48138), .X(n48139) );
  inv_x2_sg U55565 ( .A(n48140), .X(n48141) );
  inv_x2_sg U55566 ( .A(n48142), .X(n48143) );
  inv_x2_sg U55567 ( .A(n48144), .X(n48145) );
  inv_x2_sg U55568 ( .A(n48146), .X(n48147) );
  inv_x2_sg U55569 ( .A(n48148), .X(n48149) );
  inv_x2_sg U55570 ( .A(n48150), .X(n48151) );
  inv_x2_sg U55571 ( .A(n48152), .X(n48153) );
  inv_x2_sg U55572 ( .A(n48154), .X(n48155) );
  inv_x2_sg U55573 ( .A(n48156), .X(n48157) );
  inv_x2_sg U55574 ( .A(n48158), .X(n48159) );
  inv_x2_sg U55575 ( .A(n48160), .X(n48161) );
  inv_x2_sg U55576 ( .A(n48162), .X(n48163) );
  inv_x2_sg U55577 ( .A(n48164), .X(n48165) );
  inv_x2_sg U55578 ( .A(n48166), .X(n48167) );
  inv_x2_sg U55579 ( .A(n48168), .X(n48169) );
  inv_x2_sg U55580 ( .A(n48170), .X(n48171) );
  inv_x2_sg U55581 ( .A(n48172), .X(n48173) );
  inv_x2_sg U55582 ( .A(n48174), .X(n48175) );
  inv_x2_sg U55583 ( .A(n48176), .X(n48177) );
  inv_x2_sg U55584 ( .A(n48178), .X(n48179) );
  inv_x2_sg U55585 ( .A(n48180), .X(n48181) );
  inv_x2_sg U55586 ( .A(n48182), .X(n48183) );
  inv_x2_sg U55587 ( .A(n48184), .X(n48185) );
  inv_x2_sg U55588 ( .A(n48186), .X(n48187) );
  inv_x2_sg U55589 ( .A(n48188), .X(n48189) );
  inv_x2_sg U55590 ( .A(n48190), .X(n48191) );
  inv_x2_sg U55591 ( .A(n48192), .X(n48193) );
  inv_x2_sg U55592 ( .A(n48194), .X(n48195) );
  inv_x2_sg U55593 ( .A(n48196), .X(n48197) );
  inv_x2_sg U55594 ( .A(n48198), .X(n48199) );
  inv_x2_sg U55595 ( .A(n48200), .X(n48201) );
  inv_x2_sg U55596 ( .A(n48202), .X(n48203) );
  inv_x2_sg U55597 ( .A(n48204), .X(n48205) );
  inv_x2_sg U55598 ( .A(n48206), .X(n48207) );
  inv_x2_sg U55599 ( .A(n48208), .X(n48209) );
  inv_x2_sg U55600 ( .A(n48210), .X(n48211) );
  inv_x2_sg U55601 ( .A(n48212), .X(n48213) );
  inv_x2_sg U55602 ( .A(n48214), .X(n48215) );
  inv_x2_sg U55603 ( .A(n48216), .X(n48217) );
  inv_x2_sg U55604 ( .A(n48218), .X(n48219) );
  inv_x2_sg U55605 ( .A(n48220), .X(n48221) );
  inv_x2_sg U55606 ( .A(n48222), .X(n48223) );
  inv_x2_sg U55607 ( .A(n48224), .X(n48225) );
  inv_x2_sg U55608 ( .A(n48226), .X(n48227) );
  inv_x2_sg U55609 ( .A(n48228), .X(n48229) );
  inv_x2_sg U55610 ( .A(n48230), .X(n48231) );
  inv_x2_sg U55611 ( .A(n48232), .X(n48233) );
  inv_x2_sg U55612 ( .A(n48234), .X(n48235) );
  inv_x2_sg U55613 ( .A(n48236), .X(n48237) );
  inv_x2_sg U55614 ( .A(n48238), .X(n48239) );
  inv_x2_sg U55615 ( .A(n48240), .X(n48241) );
  inv_x2_sg U55616 ( .A(n48242), .X(n48243) );
  inv_x2_sg U55617 ( .A(n48244), .X(n48245) );
  inv_x2_sg U55618 ( .A(n48246), .X(n48247) );
  inv_x2_sg U55619 ( .A(n48248), .X(n48249) );
  inv_x2_sg U55620 ( .A(n48250), .X(n48251) );
  inv_x2_sg U55621 ( .A(n48252), .X(n48253) );
  inv_x2_sg U55622 ( .A(n48254), .X(n48255) );
  inv_x2_sg U55623 ( .A(n48256), .X(n48257) );
  inv_x2_sg U55624 ( .A(n48258), .X(n48259) );
  inv_x2_sg U55625 ( .A(n48260), .X(n48261) );
  inv_x2_sg U55626 ( .A(n48262), .X(n48263) );
  inv_x2_sg U55627 ( .A(n48264), .X(n48265) );
  inv_x2_sg U55628 ( .A(n48266), .X(n48267) );
  inv_x2_sg U55629 ( .A(n48268), .X(n48269) );
  inv_x2_sg U55630 ( .A(n48270), .X(n48271) );
  inv_x2_sg U55631 ( .A(n48272), .X(n48273) );
  inv_x2_sg U55632 ( .A(n48274), .X(n48275) );
  inv_x2_sg U55633 ( .A(n48276), .X(n48277) );
  inv_x2_sg U55634 ( .A(n48278), .X(n48279) );
  inv_x2_sg U55635 ( .A(n48280), .X(n48281) );
  inv_x2_sg U55636 ( .A(n48282), .X(n48283) );
  inv_x2_sg U55637 ( .A(n48284), .X(n48285) );
  inv_x2_sg U55638 ( .A(n48286), .X(n48287) );
  inv_x2_sg U55639 ( .A(n48288), .X(n48289) );
  inv_x2_sg U55640 ( .A(n48290), .X(n48291) );
  inv_x2_sg U55641 ( .A(n48292), .X(n48293) );
  inv_x2_sg U55642 ( .A(n48294), .X(n48295) );
  inv_x2_sg U55643 ( .A(n48296), .X(n48297) );
  inv_x2_sg U55644 ( .A(n48298), .X(n48299) );
  inv_x2_sg U55645 ( .A(n48300), .X(n48301) );
  inv_x2_sg U55646 ( .A(n48302), .X(n48303) );
  inv_x2_sg U55647 ( .A(n48304), .X(n48305) );
  inv_x2_sg U55648 ( .A(n48306), .X(n48307) );
  inv_x2_sg U55649 ( .A(n48308), .X(n48309) );
  inv_x2_sg U55650 ( .A(n48310), .X(n48311) );
  inv_x2_sg U55651 ( .A(n48312), .X(n48313) );
  inv_x2_sg U55652 ( .A(n48314), .X(n48315) );
  inv_x2_sg U55653 ( .A(n48316), .X(n48317) );
  inv_x2_sg U55654 ( .A(n48318), .X(n48319) );
  inv_x2_sg U55655 ( .A(n48320), .X(n48321) );
  inv_x2_sg U55656 ( .A(n48322), .X(n48323) );
  inv_x2_sg U55657 ( .A(n48324), .X(n48325) );
  inv_x2_sg U55658 ( .A(n48326), .X(n48327) );
  inv_x2_sg U55659 ( .A(n48328), .X(n48329) );
  inv_x2_sg U55660 ( .A(n48330), .X(n48331) );
  inv_x2_sg U55661 ( .A(n48332), .X(n48333) );
  inv_x2_sg U55662 ( .A(n48334), .X(n48335) );
  inv_x2_sg U55663 ( .A(n48336), .X(n48337) );
  inv_x2_sg U55664 ( .A(n48338), .X(n48339) );
  inv_x2_sg U55665 ( .A(n48340), .X(n48341) );
  inv_x2_sg U55666 ( .A(n48342), .X(n48343) );
  inv_x2_sg U55667 ( .A(n48344), .X(n48345) );
  inv_x2_sg U55668 ( .A(n48346), .X(n48347) );
  inv_x2_sg U55669 ( .A(n48348), .X(n48349) );
  inv_x2_sg U55670 ( .A(n48350), .X(n48351) );
  inv_x2_sg U55671 ( .A(n48352), .X(n48353) );
  inv_x2_sg U55672 ( .A(n48354), .X(n48355) );
  inv_x2_sg U55673 ( .A(n48356), .X(n48357) );
  inv_x2_sg U55674 ( .A(n48358), .X(n48359) );
  inv_x2_sg U55675 ( .A(n48360), .X(n48361) );
  inv_x2_sg U55676 ( .A(n48362), .X(n48363) );
  inv_x2_sg U55677 ( .A(n48364), .X(n48365) );
  inv_x2_sg U55678 ( .A(n48366), .X(n48367) );
  inv_x2_sg U55679 ( .A(n48368), .X(n48369) );
  inv_x2_sg U55680 ( .A(n48370), .X(n48371) );
  inv_x2_sg U55681 ( .A(n48372), .X(n48373) );
  inv_x2_sg U55682 ( .A(n48374), .X(n48375) );
  inv_x2_sg U55683 ( .A(n48376), .X(n48377) );
  inv_x2_sg U55684 ( .A(n48378), .X(n48379) );
  inv_x2_sg U55685 ( .A(n48380), .X(n48381) );
  inv_x2_sg U55686 ( .A(n48382), .X(n48383) );
  inv_x2_sg U55687 ( .A(n48384), .X(n48385) );
  inv_x2_sg U55688 ( .A(n48386), .X(n48387) );
  inv_x2_sg U55689 ( .A(n48388), .X(n48389) );
  inv_x2_sg U55690 ( .A(n48390), .X(n48391) );
  inv_x2_sg U55691 ( .A(n48392), .X(n48393) );
  inv_x2_sg U55692 ( .A(n48394), .X(n48395) );
  inv_x2_sg U55693 ( .A(n48396), .X(n48397) );
  inv_x2_sg U55694 ( .A(n48398), .X(n48399) );
  inv_x2_sg U55695 ( .A(n48400), .X(n48401) );
  inv_x2_sg U55696 ( .A(n48402), .X(n48403) );
  inv_x2_sg U55697 ( .A(n48404), .X(n48405) );
  inv_x2_sg U55698 ( .A(n48406), .X(n48407) );
  inv_x2_sg U55699 ( .A(n48408), .X(n48409) );
  inv_x2_sg U55700 ( .A(n48410), .X(n48411) );
  inv_x2_sg U55701 ( .A(n48412), .X(n48413) );
  inv_x2_sg U55702 ( .A(n48414), .X(n48415) );
  inv_x2_sg U55703 ( .A(n48416), .X(n48417) );
  inv_x2_sg U55704 ( .A(n48418), .X(n48419) );
  inv_x2_sg U55705 ( .A(n48420), .X(n48421) );
  inv_x2_sg U55706 ( .A(n48422), .X(n48423) );
  inv_x2_sg U55707 ( .A(n48424), .X(n48425) );
  inv_x2_sg U55708 ( .A(n48426), .X(n48427) );
  inv_x2_sg U55709 ( .A(n48428), .X(n48429) );
  inv_x2_sg U55710 ( .A(n48430), .X(n48431) );
  inv_x2_sg U55711 ( .A(n48432), .X(n48433) );
  inv_x2_sg U55712 ( .A(n48434), .X(n48435) );
  inv_x2_sg U55713 ( .A(n48436), .X(n48437) );
  inv_x2_sg U55714 ( .A(n48438), .X(n48439) );
  inv_x2_sg U55715 ( .A(n48440), .X(n48441) );
  inv_x2_sg U55716 ( .A(n48442), .X(n48443) );
  inv_x2_sg U55717 ( .A(n48444), .X(n48445) );
  inv_x2_sg U55718 ( .A(n48446), .X(n48447) );
  inv_x2_sg U55719 ( .A(n48448), .X(n48449) );
  inv_x2_sg U55720 ( .A(n48450), .X(n48451) );
  inv_x2_sg U55721 ( .A(n48452), .X(n48453) );
  inv_x2_sg U55722 ( .A(n48454), .X(n48455) );
  inv_x2_sg U55723 ( .A(n48456), .X(n48457) );
  inv_x2_sg U55724 ( .A(n48458), .X(n48459) );
  inv_x2_sg U55725 ( .A(n48460), .X(n48461) );
  inv_x2_sg U55726 ( .A(n48462), .X(n48463) );
  inv_x2_sg U55727 ( .A(n48464), .X(n48465) );
  inv_x2_sg U55728 ( .A(n48466), .X(n48467) );
  inv_x2_sg U55729 ( .A(n48468), .X(n48469) );
  inv_x2_sg U55730 ( .A(n48470), .X(n48471) );
  inv_x2_sg U55731 ( .A(n48472), .X(n48473) );
  inv_x2_sg U55732 ( .A(n48474), .X(n48475) );
  inv_x2_sg U55733 ( .A(n48476), .X(n48477) );
  inv_x2_sg U55734 ( .A(n48478), .X(n48479) );
  inv_x2_sg U55735 ( .A(n48480), .X(n48481) );
  inv_x2_sg U55736 ( .A(n48482), .X(n48483) );
  inv_x2_sg U55737 ( .A(n48484), .X(n48485) );
  inv_x2_sg U55738 ( .A(n48486), .X(n48487) );
  inv_x2_sg U55739 ( .A(n48488), .X(n48489) );
  inv_x2_sg U55740 ( .A(n48490), .X(n48491) );
  inv_x2_sg U55741 ( .A(n48492), .X(n48493) );
  inv_x2_sg U55742 ( .A(n48494), .X(n48495) );
  inv_x2_sg U55743 ( .A(n48496), .X(n48497) );
  inv_x2_sg U55744 ( .A(n48498), .X(n48499) );
  inv_x2_sg U55745 ( .A(n48500), .X(n48501) );
  inv_x2_sg U55746 ( .A(n48502), .X(n48503) );
  inv_x2_sg U55747 ( .A(n48504), .X(n48505) );
  inv_x2_sg U55748 ( .A(n48506), .X(n48507) );
  inv_x2_sg U55749 ( .A(n48508), .X(n48509) );
  inv_x2_sg U55750 ( .A(n48510), .X(n48511) );
  inv_x2_sg U55751 ( .A(n48512), .X(n48513) );
  inv_x2_sg U55752 ( .A(n48514), .X(n48515) );
  inv_x2_sg U55753 ( .A(n48516), .X(n48517) );
  inv_x2_sg U55754 ( .A(n48518), .X(n48519) );
  inv_x2_sg U55755 ( .A(n48520), .X(n48521) );
  inv_x2_sg U55756 ( .A(n48522), .X(n48523) );
  inv_x2_sg U55757 ( .A(n48524), .X(n48525) );
  inv_x2_sg U55758 ( .A(n48526), .X(n48527) );
  inv_x2_sg U55759 ( .A(n48528), .X(n48529) );
  inv_x2_sg U55760 ( .A(n48530), .X(n48531) );
  inv_x2_sg U55761 ( .A(n48532), .X(n48533) );
  inv_x2_sg U55762 ( .A(n48534), .X(n48535) );
  inv_x2_sg U55763 ( .A(n48536), .X(n48537) );
  inv_x2_sg U55764 ( .A(n48538), .X(n48539) );
  inv_x2_sg U55765 ( .A(n48540), .X(n48541) );
  inv_x2_sg U55766 ( .A(n48542), .X(n48543) );
  inv_x2_sg U55767 ( .A(n48544), .X(n48545) );
  inv_x2_sg U55768 ( .A(n48546), .X(n48547) );
  inv_x2_sg U55769 ( .A(n48548), .X(n48549) );
  inv_x2_sg U55770 ( .A(n48550), .X(n48551) );
  inv_x2_sg U55771 ( .A(n48552), .X(n48553) );
  inv_x2_sg U55772 ( .A(n48554), .X(n48555) );
  inv_x2_sg U55773 ( .A(n48556), .X(n48557) );
  inv_x2_sg U55774 ( .A(n48558), .X(n48559) );
  inv_x2_sg U55775 ( .A(n48560), .X(n48561) );
  inv_x2_sg U55776 ( .A(n48562), .X(n48563) );
  inv_x2_sg U55777 ( .A(n48564), .X(n48565) );
  inv_x2_sg U55778 ( .A(n48566), .X(n48567) );
  inv_x2_sg U55779 ( .A(n48568), .X(n48569) );
  inv_x2_sg U55780 ( .A(n48570), .X(n48571) );
  inv_x2_sg U55781 ( .A(n48572), .X(n48573) );
  inv_x2_sg U55782 ( .A(n48574), .X(n48575) );
  inv_x2_sg U55783 ( .A(n48576), .X(n48577) );
  inv_x2_sg U55784 ( .A(n48578), .X(n48579) );
  inv_x2_sg U55785 ( .A(n48580), .X(n48581) );
  inv_x2_sg U55786 ( .A(n48582), .X(n48583) );
  inv_x2_sg U55787 ( .A(n48584), .X(n48585) );
  inv_x2_sg U55788 ( .A(n48586), .X(n48587) );
  inv_x2_sg U55789 ( .A(n48588), .X(n48589) );
  inv_x2_sg U55790 ( .A(n48590), .X(n48591) );
  inv_x2_sg U55791 ( .A(n48592), .X(n48593) );
  inv_x2_sg U55792 ( .A(n48594), .X(n48595) );
  inv_x2_sg U55793 ( .A(n48596), .X(n48597) );
  inv_x2_sg U55794 ( .A(n48598), .X(n48599) );
  inv_x2_sg U55795 ( .A(n48600), .X(n48601) );
  inv_x2_sg U55796 ( .A(n48602), .X(n48603) );
  inv_x2_sg U55797 ( .A(n48604), .X(n48605) );
  inv_x2_sg U55798 ( .A(n48606), .X(n48607) );
  inv_x2_sg U55799 ( .A(n48608), .X(n48609) );
  inv_x2_sg U55800 ( .A(n48610), .X(n48611) );
  inv_x2_sg U55801 ( .A(n48612), .X(n48613) );
  inv_x2_sg U55802 ( .A(n48614), .X(n48615) );
  inv_x2_sg U55803 ( .A(n48616), .X(n48617) );
  inv_x2_sg U55804 ( .A(n48618), .X(n48619) );
  inv_x2_sg U55805 ( .A(n48620), .X(n48621) );
  inv_x2_sg U55806 ( .A(n48622), .X(n48623) );
  inv_x2_sg U55807 ( .A(n48624), .X(n48625) );
  inv_x2_sg U55808 ( .A(n48626), .X(n48627) );
  inv_x2_sg U55809 ( .A(n48628), .X(n48629) );
  inv_x2_sg U55810 ( .A(n48630), .X(n48631) );
  inv_x2_sg U55811 ( .A(n48632), .X(n48633) );
  inv_x2_sg U55812 ( .A(n48634), .X(n48635) );
  inv_x2_sg U55813 ( .A(n48636), .X(n48637) );
  inv_x2_sg U55814 ( .A(n48638), .X(n48639) );
  inv_x2_sg U55815 ( .A(n48640), .X(n48641) );
  inv_x2_sg U55816 ( .A(n48642), .X(n48643) );
  inv_x2_sg U55817 ( .A(n48644), .X(n48645) );
  inv_x2_sg U55818 ( .A(n48646), .X(n48647) );
  inv_x2_sg U55819 ( .A(n48648), .X(n48649) );
  inv_x2_sg U55820 ( .A(n48650), .X(n48651) );
  inv_x2_sg U55821 ( .A(n48652), .X(n48653) );
  inv_x2_sg U55822 ( .A(n48654), .X(n48655) );
  inv_x2_sg U55823 ( .A(n48656), .X(n48657) );
  inv_x2_sg U55824 ( .A(n48658), .X(n48659) );
  inv_x2_sg U55825 ( .A(n48660), .X(n48661) );
  inv_x2_sg U55826 ( .A(n48662), .X(n48663) );
  inv_x2_sg U55827 ( .A(n48664), .X(n48665) );
  inv_x2_sg U55828 ( .A(n48666), .X(n48667) );
  inv_x2_sg U55829 ( .A(n48668), .X(n48669) );
  inv_x2_sg U55830 ( .A(n48670), .X(n48671) );
  inv_x2_sg U55831 ( .A(n48672), .X(n48673) );
  inv_x2_sg U55832 ( .A(n48674), .X(n48675) );
  inv_x2_sg U55833 ( .A(n48676), .X(n48677) );
  inv_x2_sg U55834 ( .A(n48678), .X(n48679) );
  inv_x2_sg U55835 ( .A(n48680), .X(n48681) );
  inv_x2_sg U55836 ( .A(n48682), .X(n48683) );
  inv_x2_sg U55837 ( .A(n48684), .X(n48685) );
  inv_x2_sg U55838 ( .A(n48686), .X(n48687) );
  inv_x2_sg U55839 ( .A(n48688), .X(n48689) );
  inv_x2_sg U55840 ( .A(n48690), .X(n48691) );
  inv_x2_sg U55841 ( .A(n48692), .X(n48693) );
  inv_x2_sg U55842 ( .A(n48694), .X(n48695) );
  inv_x2_sg U55843 ( .A(n48696), .X(n48697) );
  inv_x2_sg U55844 ( .A(n48698), .X(n48699) );
  inv_x2_sg U55845 ( .A(n48700), .X(n48701) );
  inv_x2_sg U55846 ( .A(n48702), .X(n48703) );
  inv_x2_sg U55847 ( .A(n48704), .X(n48705) );
  inv_x2_sg U55848 ( .A(n48706), .X(n48707) );
  inv_x2_sg U55849 ( .A(n48708), .X(n48709) );
  inv_x2_sg U55850 ( .A(n48710), .X(n48711) );
  inv_x2_sg U55851 ( .A(n48712), .X(n48713) );
  inv_x2_sg U55852 ( .A(n48714), .X(n48715) );
  inv_x2_sg U55853 ( .A(n48716), .X(n48717) );
  inv_x2_sg U55854 ( .A(n48718), .X(n48719) );
  inv_x2_sg U55855 ( .A(n48720), .X(n48721) );
  inv_x2_sg U55856 ( .A(n48722), .X(n48723) );
  inv_x2_sg U55857 ( .A(n48724), .X(n48725) );
  inv_x2_sg U55858 ( .A(n48726), .X(n48727) );
  inv_x2_sg U55859 ( .A(n48728), .X(n48729) );
  inv_x2_sg U55860 ( .A(n48730), .X(n48731) );
  inv_x2_sg U55861 ( .A(n48732), .X(n48733) );
  inv_x2_sg U55862 ( .A(n48734), .X(n48735) );
  inv_x2_sg U55863 ( .A(n48736), .X(n48737) );
  inv_x2_sg U55864 ( .A(n48738), .X(n48739) );
  inv_x2_sg U55865 ( .A(n48740), .X(n48741) );
  inv_x2_sg U55866 ( .A(n48742), .X(n48743) );
  inv_x2_sg U55867 ( .A(n48744), .X(n48745) );
  inv_x2_sg U55868 ( .A(n48746), .X(n48747) );
  inv_x2_sg U55869 ( .A(n48748), .X(n48749) );
  inv_x2_sg U55870 ( .A(n48750), .X(n48751) );
  inv_x2_sg U55871 ( .A(n48752), .X(n48753) );
  inv_x2_sg U55872 ( .A(n48754), .X(n48755) );
  inv_x2_sg U55873 ( .A(n48756), .X(n48757) );
  inv_x2_sg U55874 ( .A(n48758), .X(n48759) );
  inv_x2_sg U55875 ( .A(n48760), .X(n48761) );
  inv_x2_sg U55876 ( .A(n48762), .X(n48763) );
  inv_x2_sg U55877 ( .A(n48764), .X(n48765) );
  inv_x2_sg U55878 ( .A(n48766), .X(n48767) );
  inv_x2_sg U55879 ( .A(n48768), .X(n48769) );
  inv_x2_sg U55880 ( .A(n48770), .X(n48771) );
  inv_x2_sg U55881 ( .A(n48772), .X(n48773) );
  inv_x2_sg U55882 ( .A(n48774), .X(n48775) );
  inv_x2_sg U55883 ( .A(n48776), .X(n48777) );
  inv_x2_sg U55884 ( .A(n48778), .X(n48779) );
  inv_x2_sg U55885 ( .A(n48780), .X(n48781) );
  inv_x2_sg U55886 ( .A(n48782), .X(n48783) );
  inv_x2_sg U55887 ( .A(n48784), .X(n48785) );
  inv_x2_sg U55888 ( .A(n48786), .X(n48787) );
  inv_x2_sg U55889 ( .A(n48788), .X(n48789) );
  inv_x2_sg U55890 ( .A(n48790), .X(n48791) );
  inv_x2_sg U55891 ( .A(n48792), .X(n48793) );
  inv_x2_sg U55892 ( .A(n48794), .X(n48795) );
  inv_x2_sg U55893 ( .A(n48796), .X(n48797) );
  inv_x2_sg U55894 ( .A(n48798), .X(n48799) );
  inv_x2_sg U55895 ( .A(n48800), .X(n48801) );
  inv_x2_sg U55896 ( .A(n48802), .X(n48803) );
  inv_x2_sg U55897 ( .A(n48804), .X(n48805) );
  inv_x2_sg U55898 ( .A(n48806), .X(n48807) );
  inv_x2_sg U55899 ( .A(n48808), .X(n48809) );
  inv_x2_sg U55900 ( .A(n48810), .X(n48811) );
  inv_x2_sg U55901 ( .A(n48812), .X(n48813) );
  inv_x2_sg U55902 ( .A(n48814), .X(n48815) );
  inv_x2_sg U55903 ( .A(n48816), .X(n48817) );
  inv_x2_sg U55904 ( .A(n48818), .X(n48819) );
  inv_x2_sg U55905 ( .A(n48820), .X(n48821) );
  inv_x2_sg U55906 ( .A(n48822), .X(n48823) );
  inv_x2_sg U55907 ( .A(n48824), .X(n48825) );
  inv_x2_sg U55908 ( .A(n48826), .X(n48827) );
  inv_x2_sg U55909 ( .A(n48828), .X(n48829) );
  inv_x2_sg U55910 ( .A(n48830), .X(n48831) );
  inv_x2_sg U55911 ( .A(n48832), .X(n48833) );
  inv_x2_sg U55912 ( .A(n48834), .X(n48835) );
  inv_x2_sg U55913 ( .A(n48836), .X(n48837) );
  inv_x2_sg U55914 ( .A(n48838), .X(n48839) );
  inv_x2_sg U55915 ( .A(n48840), .X(n48841) );
  inv_x2_sg U55916 ( .A(n48842), .X(n48843) );
  inv_x2_sg U55917 ( .A(n48844), .X(n48845) );
  inv_x2_sg U55918 ( .A(n48846), .X(n48847) );
  inv_x2_sg U55919 ( .A(n48848), .X(n48849) );
  inv_x2_sg U55920 ( .A(n48850), .X(n48851) );
  inv_x2_sg U55921 ( .A(n48852), .X(n48853) );
  inv_x2_sg U55922 ( .A(n48854), .X(n48855) );
  inv_x2_sg U55923 ( .A(n48856), .X(n48857) );
  inv_x2_sg U55924 ( .A(n48858), .X(n48859) );
  inv_x2_sg U55925 ( .A(n48860), .X(n48861) );
  inv_x2_sg U55926 ( .A(n48862), .X(n48863) );
  inv_x2_sg U55927 ( .A(n48864), .X(n48865) );
  inv_x2_sg U55928 ( .A(n48866), .X(n48867) );
  inv_x2_sg U55929 ( .A(n48868), .X(n48869) );
  inv_x2_sg U55930 ( .A(n48870), .X(n48871) );
  inv_x2_sg U55931 ( .A(n48872), .X(n48873) );
  inv_x2_sg U55932 ( .A(n48874), .X(n48875) );
  inv_x2_sg U55933 ( .A(n48876), .X(n48877) );
  inv_x2_sg U55934 ( .A(n48878), .X(n48879) );
  inv_x2_sg U55935 ( .A(n48880), .X(n48881) );
  inv_x2_sg U55936 ( .A(n48882), .X(n48883) );
  inv_x2_sg U55937 ( .A(n48884), .X(n48885) );
  inv_x2_sg U55938 ( .A(n48886), .X(n48887) );
  inv_x2_sg U55939 ( .A(n48888), .X(n48889) );
  inv_x2_sg U55940 ( .A(n48890), .X(n48891) );
  inv_x2_sg U55941 ( .A(n48892), .X(n48893) );
  inv_x2_sg U55942 ( .A(n48894), .X(n48895) );
  inv_x2_sg U55943 ( .A(n48896), .X(n48897) );
  inv_x2_sg U55944 ( .A(n48898), .X(n48899) );
  inv_x2_sg U55945 ( .A(n48900), .X(n48901) );
  inv_x2_sg U55946 ( .A(n48902), .X(n48903) );
  inv_x2_sg U55947 ( .A(n48904), .X(n48905) );
  inv_x2_sg U55948 ( .A(n48906), .X(n48907) );
  inv_x2_sg U55949 ( .A(n48908), .X(n48909) );
  inv_x2_sg U55950 ( .A(n48910), .X(n48911) );
  inv_x2_sg U55951 ( .A(n48912), .X(n48913) );
  inv_x2_sg U55952 ( .A(n48914), .X(n48915) );
  inv_x2_sg U55953 ( .A(n48916), .X(n48917) );
  inv_x2_sg U55954 ( .A(n48918), .X(n48919) );
  inv_x2_sg U55955 ( .A(n48920), .X(n48921) );
  inv_x2_sg U55956 ( .A(n48922), .X(n48923) );
  inv_x2_sg U55957 ( .A(n48924), .X(n48925) );
  inv_x2_sg U55958 ( .A(n48926), .X(n48927) );
  inv_x2_sg U55959 ( .A(n48928), .X(n48929) );
  inv_x2_sg U55960 ( .A(n48930), .X(n48931) );
  inv_x2_sg U55961 ( .A(n48932), .X(n48933) );
  inv_x2_sg U55962 ( .A(n48934), .X(n48935) );
  inv_x2_sg U55963 ( .A(n48936), .X(n48937) );
  inv_x2_sg U55964 ( .A(n48938), .X(n48939) );
  inv_x2_sg U55965 ( .A(n48940), .X(n48941) );
  inv_x2_sg U55966 ( .A(n48942), .X(n48943) );
  inv_x2_sg U55967 ( .A(n48944), .X(n48945) );
  inv_x2_sg U55968 ( .A(n48946), .X(n48947) );
  inv_x2_sg U55969 ( .A(n48948), .X(n48949) );
  inv_x2_sg U55970 ( .A(n48950), .X(n48951) );
  inv_x2_sg U55971 ( .A(n48952), .X(n48953) );
  inv_x2_sg U55972 ( .A(n48954), .X(n48955) );
  inv_x2_sg U55973 ( .A(n48956), .X(n48957) );
  inv_x2_sg U55974 ( .A(n48958), .X(n48959) );
  inv_x2_sg U55975 ( .A(n48960), .X(n48961) );
  inv_x2_sg U55976 ( .A(n48962), .X(n48963) );
  inv_x2_sg U55977 ( .A(n48964), .X(n48965) );
  inv_x2_sg U55978 ( .A(n48966), .X(n48967) );
  inv_x2_sg U55979 ( .A(n48968), .X(n48969) );
  inv_x2_sg U55980 ( .A(n48970), .X(n48971) );
  inv_x2_sg U55981 ( .A(n48972), .X(n48973) );
  inv_x2_sg U55982 ( .A(n48974), .X(n48975) );
  inv_x2_sg U55983 ( .A(n48976), .X(n48977) );
  inv_x2_sg U55984 ( .A(n48978), .X(n48979) );
  inv_x2_sg U55985 ( .A(n48980), .X(n48981) );
  inv_x2_sg U55986 ( .A(n48982), .X(n48983) );
  inv_x2_sg U55987 ( .A(n48984), .X(n48985) );
  inv_x2_sg U55988 ( .A(n48986), .X(n48987) );
  inv_x2_sg U55989 ( .A(n48988), .X(n48989) );
  inv_x2_sg U55990 ( .A(n48990), .X(n48991) );
  inv_x2_sg U55991 ( .A(n48992), .X(n48993) );
  inv_x2_sg U55992 ( .A(n48994), .X(n48995) );
  inv_x2_sg U55993 ( .A(n48996), .X(n48997) );
  inv_x2_sg U55994 ( .A(n48998), .X(n48999) );
  inv_x2_sg U55995 ( .A(n49000), .X(n49001) );
  inv_x2_sg U55996 ( .A(n49002), .X(n49003) );
  inv_x2_sg U55997 ( .A(n49004), .X(n49005) );
  inv_x2_sg U55998 ( .A(n49006), .X(n49007) );
  inv_x2_sg U55999 ( .A(n49008), .X(n49009) );
  inv_x2_sg U56000 ( .A(n49010), .X(n49011) );
  inv_x2_sg U56001 ( .A(n49012), .X(n49013) );
  inv_x2_sg U56002 ( .A(n49014), .X(n49015) );
  inv_x2_sg U56003 ( .A(n49016), .X(n49017) );
  inv_x2_sg U56004 ( .A(n49018), .X(n49019) );
  inv_x2_sg U56005 ( .A(n49020), .X(n49021) );
  inv_x2_sg U56006 ( .A(n49022), .X(n49023) );
  inv_x2_sg U56007 ( .A(n49024), .X(n49025) );
  inv_x2_sg U56008 ( .A(n49026), .X(n49027) );
  inv_x2_sg U56009 ( .A(n49028), .X(n49029) );
  inv_x2_sg U56010 ( .A(n49030), .X(n49031) );
  inv_x2_sg U56011 ( .A(n49032), .X(n49033) );
  inv_x2_sg U56012 ( .A(n49034), .X(n49035) );
  inv_x2_sg U56013 ( .A(n49036), .X(n49037) );
  inv_x2_sg U56014 ( .A(n49038), .X(n49039) );
  inv_x2_sg U56015 ( .A(n49040), .X(n49041) );
  inv_x2_sg U56016 ( .A(n49042), .X(n49043) );
  inv_x2_sg U56017 ( .A(n49044), .X(n49045) );
  inv_x2_sg U56018 ( .A(n49046), .X(n49047) );
  inv_x2_sg U56019 ( .A(n49048), .X(n49049) );
  inv_x2_sg U56020 ( .A(n49050), .X(n49051) );
  inv_x2_sg U56021 ( .A(n49052), .X(n49053) );
  inv_x2_sg U56022 ( .A(n49054), .X(n49055) );
  inv_x2_sg U56023 ( .A(n49056), .X(n49057) );
  inv_x2_sg U56024 ( .A(n49058), .X(n49059) );
  inv_x2_sg U56025 ( .A(n49060), .X(n49061) );
  inv_x2_sg U56026 ( .A(n49062), .X(n49063) );
  inv_x2_sg U56027 ( .A(n49064), .X(n49065) );
  inv_x2_sg U56028 ( .A(n49066), .X(n49067) );
  inv_x2_sg U56029 ( .A(n49068), .X(n49069) );
  inv_x2_sg U56030 ( .A(n49070), .X(n49071) );
  inv_x2_sg U56031 ( .A(n49072), .X(n49073) );
  inv_x2_sg U56032 ( .A(n49074), .X(n49075) );
  inv_x2_sg U56033 ( .A(n49076), .X(n49077) );
  inv_x2_sg U56034 ( .A(n49078), .X(n49079) );
  inv_x2_sg U56035 ( .A(n49080), .X(n49081) );
  inv_x2_sg U56036 ( .A(n49082), .X(n49083) );
  inv_x2_sg U56037 ( .A(n49084), .X(n49085) );
  inv_x2_sg U56038 ( .A(n49086), .X(n49087) );
  inv_x2_sg U56039 ( .A(n49088), .X(n49089) );
  inv_x2_sg U56040 ( .A(n49090), .X(n49091) );
  inv_x2_sg U56041 ( .A(n49092), .X(n49093) );
  inv_x2_sg U56042 ( .A(n49094), .X(n49095) );
  inv_x2_sg U56043 ( .A(n49096), .X(n49097) );
  inv_x2_sg U56044 ( .A(n49098), .X(n49099) );
  inv_x2_sg U56045 ( .A(n49100), .X(n49101) );
  inv_x2_sg U56046 ( .A(n49102), .X(n49103) );
  inv_x2_sg U56047 ( .A(n49104), .X(n49105) );
  inv_x2_sg U56048 ( .A(n49106), .X(n49107) );
  inv_x2_sg U56049 ( .A(n49108), .X(n49109) );
  inv_x2_sg U56050 ( .A(n49110), .X(n49111) );
  inv_x2_sg U56051 ( .A(n49112), .X(n49113) );
  inv_x2_sg U56052 ( .A(n49114), .X(n49115) );
  inv_x2_sg U56053 ( .A(n49116), .X(n49117) );
  inv_x2_sg U56054 ( .A(n49118), .X(n49119) );
  inv_x2_sg U56055 ( .A(n49120), .X(n49121) );
  inv_x2_sg U56056 ( .A(n49122), .X(n49123) );
  inv_x2_sg U56057 ( .A(n49124), .X(n49125) );
  inv_x2_sg U56058 ( .A(n49126), .X(n49127) );
  inv_x2_sg U56059 ( .A(n49128), .X(n49129) );
  inv_x2_sg U56060 ( .A(n49130), .X(n49131) );
  inv_x2_sg U56061 ( .A(n49132), .X(n49133) );
  inv_x2_sg U56062 ( .A(n49134), .X(n49135) );
  inv_x2_sg U56063 ( .A(n49136), .X(n49137) );
  inv_x2_sg U56064 ( .A(n49138), .X(n49139) );
  inv_x2_sg U56065 ( .A(n49140), .X(n49141) );
  inv_x2_sg U56066 ( .A(n49142), .X(n49143) );
  inv_x2_sg U56067 ( .A(n49144), .X(n49145) );
  inv_x2_sg U56068 ( .A(n49146), .X(n49147) );
  inv_x2_sg U56069 ( .A(n49148), .X(n49149) );
  inv_x2_sg U56070 ( .A(n49150), .X(n49151) );
  inv_x2_sg U56071 ( .A(n49152), .X(n49153) );
  inv_x2_sg U56072 ( .A(n49154), .X(n49155) );
  inv_x2_sg U56073 ( .A(n49156), .X(n49157) );
  inv_x2_sg U56074 ( .A(n49158), .X(n49159) );
  inv_x2_sg U56075 ( .A(n49160), .X(n49161) );
  inv_x2_sg U56076 ( .A(n49162), .X(n49163) );
  inv_x2_sg U56077 ( .A(n49164), .X(n49165) );
  inv_x2_sg U56078 ( .A(n49166), .X(n49167) );
  inv_x2_sg U56079 ( .A(n49168), .X(n49169) );
  inv_x2_sg U56080 ( .A(n49170), .X(n49171) );
  inv_x2_sg U56081 ( .A(n49172), .X(n49173) );
  inv_x2_sg U56082 ( .A(n49174), .X(n49175) );
  inv_x2_sg U56083 ( .A(n49176), .X(n49177) );
  inv_x2_sg U56084 ( .A(n49178), .X(n49179) );
  inv_x2_sg U56085 ( .A(n49180), .X(n49181) );
  inv_x2_sg U56086 ( .A(n49182), .X(n49183) );
  inv_x2_sg U56087 ( .A(n49184), .X(n49185) );
  inv_x2_sg U56088 ( .A(n49186), .X(n49187) );
  inv_x2_sg U56089 ( .A(n49188), .X(n49189) );
  inv_x2_sg U56090 ( .A(n49190), .X(n49191) );
  inv_x2_sg U56091 ( .A(n49192), .X(n49193) );
  inv_x2_sg U56092 ( .A(n49194), .X(n49195) );
  inv_x2_sg U56093 ( .A(n49196), .X(n49197) );
  inv_x2_sg U56094 ( .A(n49198), .X(n49199) );
  inv_x2_sg U56095 ( .A(n49200), .X(n49201) );
  inv_x2_sg U56096 ( .A(n49202), .X(n49203) );
  inv_x2_sg U56097 ( .A(n49204), .X(n49205) );
  inv_x2_sg U56098 ( .A(n49206), .X(n49207) );
  inv_x2_sg U56099 ( .A(n49208), .X(n49209) );
  inv_x2_sg U56100 ( .A(n49210), .X(n49211) );
  inv_x2_sg U56101 ( .A(n49212), .X(n49213) );
  inv_x2_sg U56102 ( .A(n49214), .X(n49215) );
  inv_x2_sg U56103 ( .A(n49216), .X(n49217) );
  inv_x2_sg U56104 ( .A(n49218), .X(n49219) );
  inv_x2_sg U56105 ( .A(n49220), .X(n49221) );
  inv_x2_sg U56106 ( .A(n49222), .X(n49223) );
  inv_x2_sg U56107 ( .A(n49224), .X(n49225) );
  inv_x2_sg U56108 ( .A(n49226), .X(n49227) );
  inv_x2_sg U56109 ( .A(n49228), .X(n49229) );
  inv_x2_sg U56110 ( .A(n49230), .X(n49231) );
  inv_x2_sg U56111 ( .A(n49232), .X(n49233) );
  inv_x2_sg U56112 ( .A(n49234), .X(n49235) );
  inv_x2_sg U56113 ( .A(n49236), .X(n49237) );
  inv_x2_sg U56114 ( .A(n49238), .X(n49239) );
  inv_x2_sg U56115 ( .A(n49240), .X(n49241) );
  inv_x2_sg U56116 ( .A(n49242), .X(n49243) );
  inv_x2_sg U56117 ( .A(n49244), .X(n49245) );
  inv_x2_sg U56118 ( .A(n49246), .X(n49247) );
  inv_x2_sg U56119 ( .A(n49248), .X(n49249) );
  inv_x2_sg U56120 ( .A(n49250), .X(n49251) );
  inv_x2_sg U56121 ( .A(n49252), .X(n49253) );
  inv_x2_sg U56122 ( .A(n49254), .X(n49255) );
  inv_x2_sg U56123 ( .A(n49256), .X(n49257) );
  inv_x2_sg U56124 ( .A(n49258), .X(n49259) );
  inv_x2_sg U56125 ( .A(n49260), .X(n49261) );
  inv_x2_sg U56126 ( .A(n49262), .X(n49263) );
  inv_x2_sg U56127 ( .A(n49264), .X(n49265) );
  inv_x2_sg U56128 ( .A(n49266), .X(n49267) );
  inv_x2_sg U56129 ( .A(n49268), .X(n49269) );
  inv_x2_sg U56130 ( .A(n49270), .X(n49271) );
  inv_x2_sg U56131 ( .A(n49272), .X(n49273) );
  inv_x2_sg U56132 ( .A(n49274), .X(n49275) );
  inv_x2_sg U56133 ( .A(n49276), .X(n49277) );
  inv_x2_sg U56134 ( .A(n49278), .X(n49279) );
  inv_x2_sg U56135 ( .A(n49280), .X(n49281) );
  inv_x2_sg U56136 ( .A(n49282), .X(n49283) );
  inv_x2_sg U56137 ( .A(n49284), .X(n49285) );
  inv_x2_sg U56138 ( .A(n49286), .X(n49287) );
  inv_x2_sg U56139 ( .A(n49288), .X(n49289) );
  inv_x2_sg U56140 ( .A(n49290), .X(n49291) );
  inv_x2_sg U56141 ( .A(n49292), .X(n49293) );
  inv_x2_sg U56142 ( .A(n49294), .X(n49295) );
  inv_x2_sg U56143 ( .A(n49296), .X(n49297) );
  inv_x2_sg U56144 ( .A(n49298), .X(n49299) );
  inv_x2_sg U56145 ( .A(n49300), .X(n49301) );
  inv_x2_sg U56146 ( .A(n49302), .X(n49303) );
  inv_x2_sg U56147 ( .A(n49304), .X(n49305) );
  inv_x2_sg U56148 ( .A(n49306), .X(n49307) );
  inv_x2_sg U56149 ( .A(n49308), .X(n49309) );
  inv_x2_sg U56150 ( .A(n49310), .X(n49311) );
  inv_x2_sg U56151 ( .A(n49312), .X(n49313) );
  inv_x2_sg U56152 ( .A(n49314), .X(n49315) );
  inv_x2_sg U56153 ( .A(n49316), .X(n49317) );
  inv_x2_sg U56154 ( .A(n49318), .X(n49319) );
  inv_x2_sg U56155 ( .A(n49320), .X(n49321) );
  inv_x2_sg U56156 ( .A(n49322), .X(n49323) );
  inv_x2_sg U56157 ( .A(n49324), .X(n49325) );
  inv_x2_sg U56158 ( .A(n49326), .X(n49327) );
  inv_x2_sg U56159 ( .A(n49328), .X(n49329) );
  inv_x2_sg U56160 ( .A(n49330), .X(n49331) );
  inv_x2_sg U56161 ( .A(n49332), .X(n49333) );
  inv_x2_sg U56162 ( .A(n49334), .X(n49335) );
  inv_x2_sg U56163 ( .A(n49336), .X(n49337) );
  inv_x2_sg U56164 ( .A(n49338), .X(n49339) );
  inv_x2_sg U56165 ( .A(n49340), .X(n49341) );
  inv_x2_sg U56166 ( .A(n49342), .X(n49343) );
  inv_x2_sg U56167 ( .A(n49344), .X(n49345) );
  inv_x2_sg U56168 ( .A(n49346), .X(n49347) );
  inv_x2_sg U56169 ( .A(n49348), .X(n49349) );
  inv_x2_sg U56170 ( .A(n49350), .X(n49351) );
  inv_x2_sg U56171 ( .A(n49352), .X(n49353) );
  inv_x2_sg U56172 ( .A(n49354), .X(n49355) );
  inv_x2_sg U56173 ( .A(n49356), .X(n49357) );
  inv_x2_sg U56174 ( .A(n49358), .X(n49359) );
  inv_x2_sg U56175 ( .A(n49360), .X(n49361) );
  inv_x2_sg U56176 ( .A(n49362), .X(n49363) );
  inv_x2_sg U56177 ( .A(n49364), .X(n49365) );
  inv_x2_sg U56178 ( .A(n49366), .X(n49367) );
  inv_x2_sg U56179 ( .A(n49368), .X(n49369) );
  inv_x2_sg U56180 ( .A(n49370), .X(n49371) );
  inv_x2_sg U56181 ( .A(n49372), .X(n49373) );
  inv_x2_sg U56182 ( .A(n49374), .X(n49375) );
  inv_x2_sg U56183 ( .A(n49376), .X(n49377) );
  inv_x2_sg U56184 ( .A(n49378), .X(n49379) );
  inv_x2_sg U56185 ( .A(n49380), .X(n49381) );
  inv_x2_sg U56186 ( .A(n49382), .X(n49383) );
  inv_x2_sg U56187 ( .A(n49384), .X(n49385) );
  inv_x2_sg U56188 ( .A(n49386), .X(n49387) );
  inv_x2_sg U56189 ( .A(n49388), .X(n49389) );
  inv_x2_sg U56190 ( .A(n49390), .X(n49391) );
  inv_x2_sg U56191 ( .A(n49392), .X(n49393) );
  inv_x2_sg U56192 ( .A(n49394), .X(n49395) );
  inv_x2_sg U56193 ( .A(n49396), .X(n49397) );
  inv_x2_sg U56194 ( .A(n49398), .X(n49399) );
  inv_x2_sg U56195 ( .A(n49400), .X(n49401) );
  inv_x2_sg U56196 ( .A(n49402), .X(n49403) );
  inv_x2_sg U56197 ( .A(n49404), .X(n49405) );
  inv_x2_sg U56198 ( .A(n49406), .X(n49407) );
  inv_x2_sg U56199 ( .A(n49408), .X(n49409) );
  inv_x2_sg U56200 ( .A(n49410), .X(n49411) );
  inv_x2_sg U56201 ( .A(n49412), .X(n49413) );
  inv_x2_sg U56202 ( .A(n49414), .X(n49415) );
  inv_x2_sg U56203 ( .A(n49416), .X(n49417) );
  inv_x2_sg U56204 ( .A(n49418), .X(n49419) );
  inv_x2_sg U56205 ( .A(n49420), .X(n49421) );
  inv_x2_sg U56206 ( .A(n49422), .X(n49423) );
  inv_x2_sg U56207 ( .A(n49424), .X(n49425) );
  inv_x2_sg U56208 ( .A(n49426), .X(n49427) );
  inv_x2_sg U56209 ( .A(n49428), .X(n49429) );
  inv_x2_sg U56210 ( .A(n49430), .X(n49431) );
  inv_x2_sg U56211 ( .A(n49432), .X(n49433) );
  inv_x2_sg U56212 ( .A(n49434), .X(n49435) );
  inv_x2_sg U56213 ( .A(n49436), .X(n49437) );
  inv_x2_sg U56214 ( .A(n49438), .X(n49439) );
  inv_x2_sg U56215 ( .A(n49440), .X(n49441) );
  inv_x2_sg U56216 ( .A(n49442), .X(n49443) );
  inv_x2_sg U56217 ( .A(n49444), .X(n49445) );
  inv_x2_sg U56218 ( .A(n49446), .X(n49447) );
  inv_x2_sg U56219 ( .A(n49448), .X(n49449) );
  inv_x2_sg U56220 ( .A(n49450), .X(n49451) );
  inv_x2_sg U56221 ( .A(n49452), .X(n49453) );
  inv_x2_sg U56222 ( .A(n49454), .X(n49455) );
  inv_x2_sg U56223 ( .A(n49456), .X(n49457) );
  inv_x2_sg U56224 ( .A(n49458), .X(n49459) );
  inv_x2_sg U56225 ( .A(n49460), .X(n49461) );
  inv_x2_sg U56226 ( .A(n49462), .X(n49463) );
  inv_x2_sg U56227 ( .A(n49464), .X(n49465) );
  inv_x2_sg U56228 ( .A(n49466), .X(n49467) );
  inv_x2_sg U56229 ( .A(n49468), .X(n49469) );
  inv_x2_sg U56230 ( .A(n49470), .X(n49471) );
  inv_x2_sg U56231 ( .A(n49472), .X(n49473) );
  inv_x2_sg U56232 ( .A(n49474), .X(n49475) );
  inv_x2_sg U56233 ( .A(n49476), .X(n49477) );
  inv_x2_sg U56234 ( .A(n49478), .X(n49479) );
  inv_x2_sg U56235 ( .A(n49480), .X(n49481) );
  inv_x2_sg U56236 ( .A(n49482), .X(n49483) );
  inv_x2_sg U56237 ( .A(n49484), .X(n49485) );
  inv_x2_sg U56238 ( .A(n49486), .X(n49487) );
  inv_x2_sg U56239 ( .A(n49488), .X(n49489) );
  inv_x2_sg U56240 ( .A(n49490), .X(n49491) );
  inv_x2_sg U56241 ( .A(n49492), .X(n49493) );
  inv_x2_sg U56242 ( .A(n49494), .X(n49495) );
  inv_x2_sg U56243 ( .A(n49496), .X(n49497) );
  inv_x2_sg U56244 ( .A(n49498), .X(n49499) );
  inv_x2_sg U56245 ( .A(n49500), .X(n49501) );
  inv_x2_sg U56246 ( .A(n49502), .X(n49503) );
  inv_x2_sg U56247 ( .A(n49504), .X(n49505) );
  inv_x2_sg U56248 ( .A(n49506), .X(n49507) );
  inv_x2_sg U56249 ( .A(n49508), .X(n49509) );
  inv_x2_sg U56250 ( .A(n49510), .X(n49511) );
  inv_x2_sg U56251 ( .A(n49512), .X(n49513) );
  inv_x2_sg U56252 ( .A(n49514), .X(n49515) );
  inv_x2_sg U56253 ( .A(n49516), .X(n49517) );
  inv_x2_sg U56254 ( .A(n49518), .X(n49519) );
  inv_x2_sg U56255 ( .A(n49520), .X(n49521) );
  inv_x2_sg U56256 ( .A(n49522), .X(n49523) );
  inv_x2_sg U56257 ( .A(n49524), .X(n49525) );
  inv_x2_sg U56258 ( .A(n49526), .X(n49527) );
  inv_x2_sg U56259 ( .A(n49528), .X(n49529) );
  inv_x2_sg U56260 ( .A(n49530), .X(n49531) );
  inv_x2_sg U56261 ( .A(n49532), .X(n49533) );
  inv_x2_sg U56262 ( .A(n49534), .X(n49535) );
  inv_x2_sg U56263 ( .A(n49536), .X(n49537) );
  inv_x2_sg U56264 ( .A(n49538), .X(n49539) );
  inv_x2_sg U56265 ( .A(n49540), .X(n49541) );
  inv_x2_sg U56266 ( .A(n49542), .X(n49543) );
  inv_x2_sg U56267 ( .A(n49544), .X(n49545) );
  inv_x2_sg U56268 ( .A(n49546), .X(n49547) );
  inv_x2_sg U56269 ( .A(n49548), .X(n49549) );
  inv_x2_sg U56270 ( .A(n49550), .X(n49551) );
  inv_x2_sg U56271 ( .A(n49552), .X(n49553) );
  inv_x2_sg U56272 ( .A(n49554), .X(n49555) );
  inv_x2_sg U56273 ( .A(n49556), .X(n49557) );
  inv_x2_sg U56274 ( .A(n49558), .X(n49559) );
  inv_x2_sg U56275 ( .A(n49560), .X(n49561) );
  inv_x2_sg U56276 ( .A(n49562), .X(n49563) );
  inv_x2_sg U56277 ( .A(n49564), .X(n49565) );
  inv_x2_sg U56278 ( .A(n49566), .X(n49567) );
  inv_x2_sg U56279 ( .A(n49568), .X(n49569) );
  inv_x2_sg U56280 ( .A(n49570), .X(n49571) );
  inv_x2_sg U56281 ( .A(n49572), .X(n49573) );
  inv_x2_sg U56282 ( .A(n49574), .X(n49575) );
  inv_x2_sg U56283 ( .A(n49576), .X(n49577) );
  inv_x2_sg U56284 ( .A(n49578), .X(n49579) );
  inv_x2_sg U56285 ( .A(n49580), .X(n49581) );
  inv_x2_sg U56286 ( .A(n49582), .X(n49583) );
  inv_x2_sg U56287 ( .A(n49584), .X(n49585) );
  inv_x2_sg U56288 ( .A(n49586), .X(n49587) );
  inv_x2_sg U56289 ( .A(n49588), .X(n49589) );
  inv_x2_sg U56290 ( .A(n49590), .X(n49591) );
  inv_x2_sg U56291 ( .A(n49592), .X(n49593) );
  inv_x2_sg U56292 ( .A(n49594), .X(n49595) );
  inv_x2_sg U56293 ( .A(n49596), .X(n49597) );
  inv_x2_sg U56294 ( .A(n49598), .X(n49599) );
  inv_x2_sg U56295 ( .A(n49600), .X(n49601) );
  inv_x2_sg U56296 ( .A(n49602), .X(n49603) );
  inv_x2_sg U56297 ( .A(n49604), .X(n49605) );
  inv_x2_sg U56298 ( .A(n49606), .X(n49607) );
  inv_x2_sg U56299 ( .A(n49608), .X(n49609) );
  inv_x2_sg U56300 ( .A(n49610), .X(n49611) );
  inv_x2_sg U56301 ( .A(n49612), .X(n49613) );
  inv_x2_sg U56302 ( .A(n49614), .X(n49615) );
  inv_x2_sg U56303 ( .A(n49616), .X(n49617) );
  inv_x2_sg U56304 ( .A(n49618), .X(n49619) );
  inv_x2_sg U56305 ( .A(n49620), .X(n49621) );
  inv_x2_sg U56306 ( .A(n49622), .X(n49623) );
  inv_x2_sg U56307 ( .A(n49624), .X(n49625) );
  inv_x2_sg U56308 ( .A(n49626), .X(n49627) );
  inv_x2_sg U56309 ( .A(n49628), .X(n49629) );
  inv_x2_sg U56310 ( .A(n49630), .X(n49631) );
  inv_x2_sg U56311 ( .A(n49632), .X(n49633) );
  inv_x2_sg U56312 ( .A(n49634), .X(n49635) );
  inv_x2_sg U56313 ( .A(n49636), .X(n49637) );
  inv_x2_sg U56314 ( .A(n49638), .X(n49639) );
  inv_x2_sg U56315 ( .A(n49640), .X(n49641) );
  inv_x2_sg U56316 ( .A(n49642), .X(n49643) );
  inv_x2_sg U56317 ( .A(n49644), .X(n49645) );
  inv_x2_sg U56318 ( .A(n49646), .X(n49647) );
  inv_x2_sg U56319 ( .A(n49648), .X(n49649) );
  inv_x2_sg U56320 ( .A(n49650), .X(n49651) );
  inv_x2_sg U56321 ( .A(n49652), .X(n49653) );
  inv_x2_sg U56322 ( .A(n49654), .X(n49655) );
  inv_x2_sg U56323 ( .A(n49656), .X(n49657) );
  inv_x2_sg U56324 ( .A(n49658), .X(n49659) );
  inv_x2_sg U56325 ( .A(n49660), .X(n49661) );
  inv_x2_sg U56326 ( .A(n49662), .X(n49663) );
  inv_x2_sg U56327 ( .A(n49664), .X(n49665) );
  inv_x2_sg U56328 ( .A(n49666), .X(n49667) );
  inv_x2_sg U56329 ( .A(n49668), .X(n49669) );
  inv_x2_sg U56330 ( .A(n49670), .X(n49671) );
  inv_x2_sg U56331 ( .A(n49672), .X(n49673) );
  inv_x2_sg U56332 ( .A(n49674), .X(n49675) );
  inv_x2_sg U56333 ( .A(n49676), .X(n49677) );
  inv_x2_sg U56334 ( .A(n49678), .X(n49679) );
  inv_x2_sg U56335 ( .A(n49680), .X(n49681) );
  inv_x2_sg U56336 ( .A(n49682), .X(n49683) );
  inv_x2_sg U56337 ( .A(n49684), .X(n49685) );
  inv_x2_sg U56338 ( .A(n49686), .X(n49687) );
  inv_x2_sg U56339 ( .A(n49688), .X(n49689) );
  inv_x2_sg U56340 ( .A(n49690), .X(n49691) );
  inv_x2_sg U56341 ( .A(n49692), .X(n49693) );
  inv_x2_sg U56342 ( .A(n49694), .X(n49695) );
  inv_x2_sg U56343 ( .A(n49696), .X(n49697) );
  inv_x2_sg U56344 ( .A(n49698), .X(n49699) );
  inv_x2_sg U56345 ( .A(n49700), .X(n49701) );
  inv_x2_sg U56346 ( .A(n49702), .X(n49703) );
  inv_x2_sg U56347 ( .A(n49704), .X(n49705) );
  inv_x2_sg U56348 ( .A(n49706), .X(n49707) );
  inv_x2_sg U56349 ( .A(n49708), .X(n49709) );
  inv_x2_sg U56350 ( .A(n49710), .X(n49711) );
  inv_x2_sg U56351 ( .A(n49712), .X(n49713) );
  inv_x2_sg U56352 ( .A(n49714), .X(n49715) );
  inv_x2_sg U56353 ( .A(n49716), .X(n49717) );
  inv_x2_sg U56354 ( .A(n49718), .X(n49719) );
  inv_x2_sg U56355 ( .A(n49720), .X(n49721) );
  inv_x2_sg U56356 ( .A(n49722), .X(n49723) );
  inv_x2_sg U56357 ( .A(n49724), .X(n49725) );
  inv_x2_sg U56358 ( .A(n49726), .X(n49727) );
  inv_x2_sg U56359 ( .A(n49728), .X(n49729) );
  inv_x2_sg U56360 ( .A(n49730), .X(n49731) );
  inv_x2_sg U56361 ( .A(n49732), .X(n49733) );
  inv_x2_sg U56362 ( .A(n49734), .X(n49735) );
  inv_x2_sg U56363 ( .A(n49736), .X(n49737) );
  inv_x2_sg U56364 ( .A(n49738), .X(n49739) );
  inv_x2_sg U56365 ( .A(n49740), .X(n49741) );
  inv_x2_sg U56366 ( .A(n49742), .X(n49743) );
  inv_x2_sg U56367 ( .A(n49744), .X(n49745) );
  inv_x2_sg U56368 ( .A(n49746), .X(n49747) );
  inv_x2_sg U56369 ( .A(n49748), .X(n49749) );
  inv_x2_sg U56370 ( .A(n49750), .X(n49751) );
  inv_x2_sg U56371 ( .A(n49752), .X(n49753) );
  inv_x2_sg U56372 ( .A(n49754), .X(n49755) );
  inv_x2_sg U56373 ( .A(n49756), .X(n49757) );
  inv_x2_sg U56374 ( .A(n49758), .X(n49759) );
  inv_x2_sg U56375 ( .A(n49760), .X(n49761) );
  inv_x2_sg U56376 ( .A(n49762), .X(n49763) );
  inv_x2_sg U56377 ( .A(n49764), .X(n49765) );
  inv_x2_sg U56378 ( .A(n49766), .X(n49767) );
  inv_x2_sg U56379 ( .A(n49768), .X(n49769) );
  inv_x2_sg U56380 ( .A(n49770), .X(n49771) );
  inv_x2_sg U56381 ( .A(n49772), .X(n49773) );
  inv_x2_sg U56382 ( .A(n49774), .X(n49775) );
  inv_x2_sg U56383 ( .A(n49776), .X(n49777) );
  inv_x2_sg U56384 ( .A(n49778), .X(n49779) );
  inv_x2_sg U56385 ( .A(n49780), .X(n49781) );
  inv_x2_sg U56386 ( .A(n49782), .X(n49783) );
  inv_x2_sg U56387 ( .A(n49784), .X(n49785) );
  inv_x2_sg U56388 ( .A(n49786), .X(n49787) );
  inv_x2_sg U56389 ( .A(n49788), .X(n49789) );
  inv_x2_sg U56390 ( .A(n49790), .X(n49791) );
  inv_x2_sg U56391 ( .A(n49792), .X(n49793) );
  inv_x2_sg U56392 ( .A(n49794), .X(n49795) );
  inv_x2_sg U56393 ( .A(n49796), .X(n49797) );
  inv_x2_sg U56394 ( .A(n49798), .X(n49799) );
  inv_x2_sg U56395 ( .A(n49800), .X(n49801) );
  inv_x2_sg U56396 ( .A(n49802), .X(n49803) );
  inv_x2_sg U56397 ( .A(n49804), .X(n49805) );
  inv_x2_sg U56398 ( .A(n49806), .X(n49807) );
  inv_x2_sg U56399 ( .A(n49808), .X(n49809) );
  inv_x2_sg U56400 ( .A(n49810), .X(n49811) );
  inv_x2_sg U56401 ( .A(n49812), .X(n49813) );
  inv_x2_sg U56402 ( .A(n49814), .X(n49815) );
  inv_x2_sg U56403 ( .A(n49816), .X(n49817) );
  inv_x2_sg U56404 ( .A(n49818), .X(n49819) );
  inv_x2_sg U56405 ( .A(n49820), .X(n49821) );
  inv_x2_sg U56406 ( .A(n49822), .X(n49823) );
  inv_x2_sg U56407 ( .A(n49824), .X(n49825) );
  inv_x2_sg U56408 ( .A(n49826), .X(n49827) );
  inv_x2_sg U56409 ( .A(n49828), .X(n49829) );
  inv_x2_sg U56410 ( .A(n49830), .X(n49831) );
  inv_x2_sg U56411 ( .A(n49832), .X(n49833) );
  inv_x2_sg U56412 ( .A(n49834), .X(n49835) );
  inv_x2_sg U56413 ( .A(n49836), .X(n49837) );
  inv_x2_sg U56414 ( .A(n49838), .X(n49839) );
  inv_x2_sg U56415 ( .A(n49840), .X(n49841) );
  inv_x2_sg U56416 ( .A(n49842), .X(n49843) );
  inv_x2_sg U56417 ( .A(n49844), .X(n49845) );
  inv_x2_sg U56418 ( .A(n49846), .X(n49847) );
  inv_x2_sg U56419 ( .A(n49848), .X(n49849) );
  inv_x2_sg U56420 ( .A(n49850), .X(n49851) );
  inv_x2_sg U56421 ( .A(n49852), .X(n49853) );
  inv_x2_sg U56422 ( .A(n49854), .X(n49855) );
  inv_x2_sg U56423 ( .A(n49856), .X(n49857) );
  inv_x2_sg U56424 ( .A(n49858), .X(n49859) );
  inv_x2_sg U56425 ( .A(n49860), .X(n49861) );
  inv_x2_sg U56426 ( .A(n49862), .X(n49863) );
  inv_x2_sg U56427 ( .A(n49864), .X(n49865) );
  inv_x2_sg U56428 ( .A(n49866), .X(n49867) );
  inv_x2_sg U56429 ( .A(n49868), .X(n49869) );
  inv_x2_sg U56430 ( .A(n49870), .X(n49871) );
  inv_x2_sg U56431 ( .A(n49872), .X(n49873) );
  inv_x2_sg U56432 ( .A(n49874), .X(n49875) );
  inv_x2_sg U56433 ( .A(n49876), .X(n49877) );
  inv_x2_sg U56434 ( .A(n49878), .X(n49879) );
  inv_x2_sg U56435 ( .A(n49880), .X(n49881) );
  inv_x2_sg U56436 ( .A(n49882), .X(n49883) );
  inv_x2_sg U56437 ( .A(n49884), .X(n49885) );
  inv_x2_sg U56438 ( .A(n49886), .X(n49887) );
  inv_x2_sg U56439 ( .A(n49888), .X(n49889) );
  inv_x2_sg U56440 ( .A(n49890), .X(n49891) );
  inv_x2_sg U56441 ( .A(n49892), .X(n49893) );
  inv_x2_sg U56442 ( .A(n49894), .X(n49895) );
  inv_x2_sg U56443 ( .A(n49896), .X(n49897) );
  inv_x2_sg U56444 ( .A(n49898), .X(n49899) );
  inv_x2_sg U56445 ( .A(n49900), .X(n49901) );
  inv_x2_sg U56446 ( .A(n49902), .X(n49903) );
  inv_x2_sg U56447 ( .A(n49904), .X(n49905) );
  inv_x2_sg U56448 ( .A(n49906), .X(n49907) );
  inv_x2_sg U56449 ( .A(n49908), .X(n49909) );
  inv_x2_sg U56450 ( .A(n49910), .X(n49911) );
  inv_x2_sg U56451 ( .A(n49912), .X(n49913) );
  inv_x2_sg U56452 ( .A(n49914), .X(n49915) );
  inv_x2_sg U56453 ( .A(n49916), .X(n49917) );
  inv_x2_sg U56454 ( .A(n49918), .X(n49919) );
  inv_x2_sg U56455 ( .A(n49920), .X(n49921) );
  inv_x2_sg U56456 ( .A(n49922), .X(n49923) );
  inv_x2_sg U56457 ( .A(n49924), .X(n49925) );
  inv_x2_sg U56458 ( .A(n49926), .X(n49927) );
  inv_x2_sg U56459 ( .A(n49928), .X(n49929) );
  inv_x2_sg U56460 ( .A(n49930), .X(n49931) );
  inv_x2_sg U56461 ( .A(n49932), .X(n49933) );
  inv_x2_sg U56462 ( .A(n49934), .X(n49935) );
  inv_x2_sg U56463 ( .A(n49936), .X(n49937) );
  inv_x2_sg U56464 ( .A(n49938), .X(n49939) );
  inv_x2_sg U56465 ( .A(n49940), .X(n49941) );
  inv_x2_sg U56466 ( .A(n49942), .X(n49943) );
  inv_x2_sg U56467 ( .A(n49944), .X(n49945) );
  inv_x2_sg U56468 ( .A(n49946), .X(n49947) );
  inv_x2_sg U56469 ( .A(n49948), .X(n49949) );
  inv_x2_sg U56470 ( .A(n49950), .X(n49951) );
  inv_x2_sg U56471 ( .A(n49952), .X(n49953) );
  inv_x2_sg U56472 ( .A(n49954), .X(n49955) );
  inv_x2_sg U56473 ( .A(n49956), .X(n49957) );
  inv_x2_sg U56474 ( .A(n49958), .X(n49959) );
  inv_x2_sg U56475 ( .A(n49960), .X(n49961) );
  inv_x2_sg U56476 ( .A(n49962), .X(n49963) );
  inv_x2_sg U56477 ( .A(n49964), .X(n49965) );
  inv_x2_sg U56478 ( .A(n49966), .X(n49967) );
  inv_x2_sg U56479 ( .A(n49968), .X(n49969) );
  inv_x2_sg U56480 ( .A(n49970), .X(n49971) );
  inv_x2_sg U56481 ( .A(n49972), .X(n49973) );
  inv_x2_sg U56482 ( .A(n49974), .X(n49975) );
  inv_x2_sg U56483 ( .A(n49976), .X(n49977) );
  inv_x2_sg U56484 ( .A(n49978), .X(n49979) );
  inv_x2_sg U56485 ( .A(n49980), .X(n49981) );
  inv_x2_sg U56486 ( .A(n49982), .X(n49983) );
  inv_x2_sg U56487 ( .A(n49984), .X(n49985) );
  inv_x2_sg U56488 ( .A(n49986), .X(n49987) );
  inv_x2_sg U56489 ( .A(n49988), .X(n49989) );
  inv_x2_sg U56490 ( .A(n49990), .X(n49991) );
  inv_x2_sg U56491 ( .A(n49992), .X(n49993) );
  inv_x2_sg U56492 ( .A(n49994), .X(n49995) );
  inv_x2_sg U56493 ( .A(n49996), .X(n49997) );
  inv_x2_sg U56494 ( .A(n49998), .X(n49999) );
  inv_x2_sg U56495 ( .A(n50000), .X(n50001) );
  inv_x2_sg U56496 ( .A(n50002), .X(n50003) );
  inv_x2_sg U56497 ( .A(n50004), .X(n50005) );
  inv_x2_sg U56498 ( .A(n50006), .X(n50007) );
  inv_x2_sg U56499 ( .A(n50008), .X(n50009) );
  inv_x2_sg U56500 ( .A(n50010), .X(n50011) );
  inv_x2_sg U56501 ( .A(n50012), .X(n50013) );
  inv_x2_sg U56502 ( .A(n50014), .X(n50015) );
  inv_x2_sg U56503 ( .A(n50016), .X(n50017) );
  inv_x2_sg U56504 ( .A(n50018), .X(n50019) );
  inv_x2_sg U56505 ( .A(n50020), .X(n50021) );
  inv_x2_sg U56506 ( .A(n50022), .X(n50023) );
  inv_x2_sg U56507 ( .A(n50024), .X(n50025) );
  inv_x2_sg U56508 ( .A(n50026), .X(n50027) );
  inv_x2_sg U56509 ( .A(n50028), .X(n50029) );
  inv_x2_sg U56510 ( .A(n50030), .X(n50031) );
  inv_x2_sg U56511 ( .A(n50032), .X(n50033) );
  inv_x2_sg U56512 ( .A(n50034), .X(n50035) );
  inv_x2_sg U56513 ( .A(n50036), .X(n50037) );
  inv_x2_sg U56514 ( .A(n50038), .X(n50039) );
  inv_x2_sg U56515 ( .A(n50040), .X(n50041) );
  inv_x2_sg U56516 ( .A(n50042), .X(n50043) );
  inv_x2_sg U56517 ( .A(n50044), .X(n50045) );
  inv_x2_sg U56518 ( .A(n50046), .X(n50047) );
  inv_x2_sg U56519 ( .A(n50048), .X(n50049) );
  inv_x2_sg U56520 ( .A(n50050), .X(n50051) );
  inv_x2_sg U56521 ( .A(n50052), .X(n50053) );
  inv_x2_sg U56522 ( .A(n50054), .X(n50055) );
  inv_x2_sg U56523 ( .A(n50056), .X(n50057) );
  inv_x2_sg U56524 ( .A(n50058), .X(n50059) );
  inv_x2_sg U56525 ( .A(n50060), .X(n50061) );
  inv_x2_sg U56526 ( .A(n50062), .X(n50063) );
  inv_x2_sg U56527 ( .A(n50064), .X(n50065) );
  inv_x2_sg U56528 ( .A(n50066), .X(n50067) );
  inv_x2_sg U56529 ( .A(n50068), .X(n50069) );
  inv_x2_sg U56530 ( .A(n50070), .X(n50071) );
  inv_x2_sg U56531 ( .A(n50072), .X(n50073) );
  inv_x2_sg U56532 ( .A(n50074), .X(n50075) );
  inv_x2_sg U56533 ( .A(n50076), .X(n50077) );
  inv_x2_sg U56534 ( .A(n50078), .X(n50079) );
  inv_x2_sg U56535 ( .A(n50080), .X(n50081) );
  inv_x2_sg U56536 ( .A(n50082), .X(n50083) );
  inv_x2_sg U56537 ( .A(n50084), .X(n50085) );
  inv_x2_sg U56538 ( .A(n50086), .X(n50087) );
  inv_x2_sg U56539 ( .A(n50088), .X(n50089) );
  inv_x2_sg U56540 ( .A(n50090), .X(n50091) );
  inv_x2_sg U56541 ( .A(n50092), .X(n50093) );
  inv_x2_sg U56542 ( .A(n50094), .X(n50095) );
  inv_x2_sg U56543 ( .A(n50096), .X(n50097) );
  inv_x2_sg U56544 ( .A(n50098), .X(n50099) );
  inv_x2_sg U56545 ( .A(n50100), .X(n50101) );
  inv_x2_sg U56546 ( .A(n50102), .X(n50103) );
  inv_x2_sg U56547 ( .A(n50104), .X(n50105) );
  inv_x2_sg U56548 ( .A(n50106), .X(n50107) );
  inv_x2_sg U56549 ( .A(n50108), .X(n50109) );
  inv_x2_sg U56550 ( .A(n50110), .X(n50111) );
  inv_x2_sg U56551 ( .A(n50112), .X(n50113) );
  inv_x2_sg U56552 ( .A(n50114), .X(n50115) );
  inv_x2_sg U56553 ( .A(n50116), .X(n50117) );
  inv_x2_sg U56554 ( .A(n50118), .X(n50119) );
  inv_x2_sg U56555 ( .A(n50120), .X(n50121) );
  inv_x2_sg U56556 ( .A(n50122), .X(n50123) );
  inv_x2_sg U56557 ( .A(n50124), .X(n50125) );
  inv_x2_sg U56558 ( .A(n50126), .X(n50127) );
  inv_x2_sg U56559 ( .A(n50128), .X(n50129) );
  inv_x2_sg U56560 ( .A(n50130), .X(n50131) );
  inv_x2_sg U56561 ( .A(n50132), .X(n50133) );
  inv_x2_sg U56562 ( .A(n50134), .X(n50135) );
  inv_x2_sg U56563 ( .A(n50136), .X(n50137) );
  inv_x2_sg U56564 ( .A(n50138), .X(n50139) );
  inv_x2_sg U56565 ( .A(n50140), .X(n50141) );
  inv_x2_sg U56566 ( .A(n50142), .X(n50143) );
  inv_x2_sg U56567 ( .A(n50144), .X(n50145) );
  inv_x2_sg U56568 ( .A(n50146), .X(n50147) );
  inv_x2_sg U56569 ( .A(n50148), .X(n50149) );
  inv_x2_sg U56570 ( .A(n50150), .X(n50151) );
  inv_x2_sg U56571 ( .A(n50152), .X(n50153) );
  inv_x2_sg U56572 ( .A(n50154), .X(n50155) );
  inv_x2_sg U56573 ( .A(n50156), .X(n50157) );
  inv_x2_sg U56574 ( .A(n50158), .X(n50159) );
  inv_x2_sg U56575 ( .A(n50160), .X(n50161) );
  inv_x2_sg U56576 ( .A(n50162), .X(n50163) );
  inv_x2_sg U56577 ( .A(n50164), .X(n50165) );
  inv_x2_sg U56578 ( .A(n50166), .X(n50167) );
  inv_x2_sg U56579 ( .A(n50168), .X(n50169) );
  inv_x2_sg U56580 ( .A(n50170), .X(n50171) );
  inv_x2_sg U56581 ( .A(n50172), .X(n50173) );
  inv_x2_sg U56582 ( .A(n50174), .X(n50175) );
  inv_x2_sg U56583 ( .A(n50176), .X(n50177) );
  inv_x2_sg U56584 ( .A(n50178), .X(n50179) );
  inv_x2_sg U56585 ( .A(n50180), .X(n50181) );
  inv_x2_sg U56586 ( .A(n50182), .X(n50183) );
  inv_x2_sg U56587 ( .A(n50184), .X(n50185) );
  inv_x2_sg U56588 ( .A(n50186), .X(n50187) );
  inv_x2_sg U56589 ( .A(n50188), .X(n50189) );
  inv_x2_sg U56590 ( .A(n50190), .X(n50191) );
  inv_x2_sg U56591 ( .A(n50192), .X(n50193) );
  inv_x2_sg U56592 ( .A(n50194), .X(n50195) );
  inv_x2_sg U56593 ( .A(n50196), .X(n50197) );
  inv_x2_sg U56594 ( .A(n50198), .X(n50199) );
  inv_x2_sg U56595 ( .A(n50200), .X(n50201) );
  inv_x2_sg U56596 ( .A(n50202), .X(n50203) );
  inv_x2_sg U56597 ( .A(n50204), .X(n50205) );
  inv_x2_sg U56598 ( .A(n50206), .X(n50207) );
  inv_x2_sg U56599 ( .A(n50208), .X(n50209) );
  inv_x2_sg U56600 ( .A(n50210), .X(n50211) );
  inv_x2_sg U56601 ( .A(n50212), .X(n50213) );
  inv_x2_sg U56602 ( .A(n50214), .X(n50215) );
  inv_x2_sg U56603 ( .A(n50216), .X(n50217) );
  inv_x2_sg U56604 ( .A(n50218), .X(n50219) );
  inv_x2_sg U56605 ( .A(n50220), .X(n50221) );
  inv_x2_sg U56606 ( .A(n50222), .X(n50223) );
  inv_x2_sg U56607 ( .A(n50224), .X(n50225) );
  inv_x2_sg U56608 ( .A(n50226), .X(n50227) );
  inv_x2_sg U56609 ( .A(n50228), .X(n50229) );
  inv_x2_sg U56610 ( .A(n50230), .X(n50231) );
  inv_x2_sg U56611 ( .A(n50232), .X(n50233) );
  inv_x2_sg U56612 ( .A(n50234), .X(n50235) );
  inv_x2_sg U56613 ( .A(n50236), .X(n50237) );
  inv_x2_sg U56614 ( .A(n50238), .X(n50239) );
  inv_x2_sg U56615 ( .A(n50240), .X(n50241) );
  inv_x2_sg U56616 ( .A(n50242), .X(n50243) );
  inv_x2_sg U56617 ( .A(n50244), .X(n50245) );
  inv_x2_sg U56618 ( .A(n50246), .X(n50247) );
  inv_x2_sg U56619 ( .A(n50248), .X(n50249) );
  inv_x2_sg U56620 ( .A(n50250), .X(n50251) );
  inv_x2_sg U56621 ( .A(n50252), .X(n50253) );
  inv_x2_sg U56622 ( .A(n50254), .X(n50255) );
  inv_x2_sg U56623 ( .A(n50256), .X(n50257) );
  inv_x2_sg U56624 ( .A(n50258), .X(n50259) );
  inv_x2_sg U56625 ( .A(n50260), .X(n50261) );
  inv_x2_sg U56626 ( .A(n50262), .X(n50263) );
  inv_x2_sg U56627 ( .A(n50264), .X(n50265) );
  inv_x2_sg U56628 ( .A(n50266), .X(n50267) );
  inv_x2_sg U56629 ( .A(n50268), .X(n50269) );
  inv_x2_sg U56630 ( .A(n50270), .X(n50271) );
  inv_x2_sg U56631 ( .A(n50272), .X(n50273) );
  inv_x2_sg U56632 ( .A(n50274), .X(n50275) );
  inv_x2_sg U56633 ( .A(n50276), .X(n50277) );
  inv_x2_sg U56634 ( .A(n50278), .X(n50279) );
  inv_x2_sg U56635 ( .A(n50280), .X(n50281) );
  inv_x2_sg U56636 ( .A(n50282), .X(n50283) );
  inv_x2_sg U56637 ( .A(n50284), .X(n50285) );
  inv_x2_sg U56638 ( .A(n50286), .X(n50287) );
  inv_x2_sg U56639 ( .A(n50288), .X(n50289) );
  inv_x2_sg U56640 ( .A(n50290), .X(n50291) );
  inv_x2_sg U56641 ( .A(n50292), .X(n50293) );
  inv_x2_sg U56642 ( .A(n50294), .X(n50295) );
  inv_x2_sg U56643 ( .A(n50296), .X(n50297) );
  inv_x2_sg U56644 ( .A(n50298), .X(n50299) );
  inv_x2_sg U56645 ( .A(n50300), .X(n50301) );
  inv_x2_sg U56646 ( .A(n50302), .X(n50303) );
  inv_x2_sg U56647 ( .A(n50304), .X(n50305) );
  inv_x2_sg U56648 ( .A(n50306), .X(n50307) );
  inv_x2_sg U56649 ( .A(n50308), .X(n50309) );
  inv_x2_sg U56650 ( .A(n50310), .X(n50311) );
  inv_x2_sg U56651 ( .A(n50312), .X(n50313) );
  inv_x2_sg U56652 ( .A(n50314), .X(n50315) );
  inv_x2_sg U56653 ( .A(n50316), .X(n50317) );
  inv_x2_sg U56654 ( .A(n50318), .X(n50319) );
  inv_x2_sg U56655 ( .A(n50320), .X(n50321) );
  inv_x2_sg U56656 ( .A(n50322), .X(n50323) );
  inv_x2_sg U56657 ( .A(n50324), .X(n50325) );
  inv_x2_sg U56658 ( .A(n50326), .X(n50327) );
  inv_x2_sg U56659 ( .A(n50328), .X(n50329) );
  inv_x2_sg U56660 ( .A(n50330), .X(n50331) );
  inv_x2_sg U56661 ( .A(n50332), .X(n50333) );
  inv_x2_sg U56662 ( .A(n50334), .X(n50335) );
  inv_x2_sg U56663 ( .A(n50336), .X(n50337) );
  inv_x2_sg U56664 ( .A(n50338), .X(n50339) );
  inv_x2_sg U56665 ( .A(n50340), .X(n50341) );
  inv_x2_sg U56666 ( .A(n50342), .X(n50343) );
  inv_x2_sg U56667 ( .A(n50344), .X(n50345) );
  inv_x2_sg U56668 ( .A(n50346), .X(n50347) );
  inv_x2_sg U56669 ( .A(n50348), .X(n50349) );
  inv_x2_sg U56670 ( .A(n50350), .X(n50351) );
  inv_x2_sg U56671 ( .A(n50352), .X(n50353) );
  inv_x2_sg U56672 ( .A(n50354), .X(n50355) );
  inv_x2_sg U56673 ( .A(n50356), .X(n50357) );
  inv_x2_sg U56674 ( .A(n50358), .X(n50359) );
  inv_x2_sg U56675 ( .A(n50360), .X(n50361) );
  inv_x2_sg U56676 ( .A(n50362), .X(n50363) );
  inv_x2_sg U56677 ( .A(n50364), .X(n50365) );
  inv_x2_sg U56678 ( .A(n50366), .X(n50367) );
  inv_x2_sg U56679 ( .A(n50368), .X(n50369) );
  inv_x2_sg U56680 ( .A(n50370), .X(n50371) );
  inv_x2_sg U56681 ( .A(n50372), .X(n50373) );
  inv_x2_sg U56682 ( .A(n50374), .X(n50375) );
  inv_x2_sg U56683 ( .A(n50376), .X(n50377) );
  inv_x2_sg U56684 ( .A(n50378), .X(n50379) );
  inv_x2_sg U56685 ( .A(n50380), .X(n50381) );
  inv_x2_sg U56686 ( .A(n50382), .X(n50383) );
  inv_x2_sg U56687 ( .A(n50384), .X(n50385) );
  inv_x2_sg U56688 ( .A(n50386), .X(n50387) );
  inv_x2_sg U56689 ( .A(n50388), .X(n50389) );
  inv_x2_sg U56690 ( .A(n50390), .X(n50391) );
  inv_x2_sg U56691 ( .A(n50392), .X(n50393) );
  inv_x2_sg U56692 ( .A(n50394), .X(n50395) );
  inv_x2_sg U56693 ( .A(n50396), .X(n50397) );
  inv_x2_sg U56694 ( .A(n50398), .X(n50399) );
  inv_x2_sg U56695 ( .A(n50400), .X(n50401) );
  inv_x2_sg U56696 ( .A(n50402), .X(n50403) );
  inv_x2_sg U56697 ( .A(n50404), .X(n50405) );
  inv_x2_sg U56698 ( .A(n50406), .X(n50407) );
  inv_x2_sg U56699 ( .A(n50408), .X(n50409) );
  inv_x2_sg U56700 ( .A(n50410), .X(n50411) );
  inv_x2_sg U56701 ( .A(n50412), .X(n50413) );
  inv_x2_sg U56702 ( .A(n50414), .X(n50415) );
  inv_x2_sg U56703 ( .A(n50416), .X(n50417) );
  inv_x2_sg U56704 ( .A(n50418), .X(n50419) );
  inv_x2_sg U56705 ( .A(n50420), .X(n50421) );
  inv_x2_sg U56706 ( .A(n50422), .X(n50423) );
  inv_x2_sg U56707 ( .A(n50424), .X(n50425) );
  inv_x2_sg U56708 ( .A(n50426), .X(n50427) );
  inv_x2_sg U56709 ( .A(n50428), .X(n50429) );
  inv_x2_sg U56710 ( .A(n50430), .X(n50431) );
  inv_x2_sg U56711 ( .A(n50432), .X(n50433) );
  inv_x2_sg U56712 ( .A(n50434), .X(n50435) );
  inv_x2_sg U56713 ( .A(n50436), .X(n50437) );
  inv_x2_sg U56714 ( .A(n50438), .X(n50439) );
  inv_x2_sg U56715 ( .A(n50440), .X(n50441) );
  inv_x2_sg U56716 ( .A(n50442), .X(n50443) );
  inv_x2_sg U56717 ( .A(n50444), .X(n50445) );
  inv_x2_sg U56718 ( .A(n50446), .X(n50447) );
  inv_x2_sg U56719 ( .A(n50448), .X(n50449) );
  inv_x2_sg U56720 ( .A(n50450), .X(n50451) );
  inv_x2_sg U56721 ( .A(n50452), .X(n50453) );
  inv_x2_sg U56722 ( .A(n50454), .X(n50455) );
  inv_x2_sg U56723 ( .A(n50456), .X(n50457) );
  inv_x2_sg U56724 ( .A(n50458), .X(n50459) );
  inv_x2_sg U56725 ( .A(n50460), .X(n50461) );
  inv_x2_sg U56726 ( .A(n50462), .X(n50463) );
  inv_x2_sg U56727 ( .A(n50464), .X(n50465) );
  inv_x2_sg U56728 ( .A(n50466), .X(n50467) );
  inv_x2_sg U56729 ( .A(n50468), .X(n50469) );
  inv_x2_sg U56730 ( .A(n50470), .X(n50471) );
  inv_x2_sg U56731 ( .A(n50472), .X(n50473) );
  inv_x2_sg U56732 ( .A(n50474), .X(n50475) );
  inv_x2_sg U56733 ( .A(n50476), .X(n50477) );
  inv_x2_sg U56734 ( .A(n50478), .X(n50479) );
  inv_x2_sg U56735 ( .A(n50480), .X(n50481) );
  inv_x2_sg U56736 ( .A(n50482), .X(n50483) );
  inv_x2_sg U56737 ( .A(n50484), .X(n50485) );
  inv_x2_sg U56738 ( .A(n50486), .X(n50487) );
  inv_x2_sg U56739 ( .A(n50488), .X(n50489) );
  inv_x2_sg U56740 ( .A(n50490), .X(n50491) );
  inv_x2_sg U56741 ( .A(n50492), .X(n50493) );
  inv_x2_sg U56742 ( .A(n50494), .X(n50495) );
  inv_x2_sg U56743 ( .A(n50496), .X(n50497) );
  inv_x2_sg U56744 ( .A(n50498), .X(n50499) );
  inv_x2_sg U56745 ( .A(n50500), .X(n50501) );
  inv_x2_sg U56746 ( .A(n50502), .X(n50503) );
  inv_x2_sg U56747 ( .A(n50504), .X(n50505) );
  inv_x2_sg U56748 ( .A(n50506), .X(n50507) );
  inv_x2_sg U56749 ( .A(n50508), .X(n50509) );
  inv_x2_sg U56750 ( .A(n50510), .X(n50511) );
  inv_x2_sg U56751 ( .A(n50512), .X(n50513) );
  inv_x2_sg U56752 ( .A(n50514), .X(n50515) );
  inv_x2_sg U56753 ( .A(n50516), .X(n50517) );
  inv_x2_sg U56754 ( .A(n50518), .X(n50519) );
  inv_x2_sg U56755 ( .A(n50520), .X(n50521) );
  inv_x2_sg U56756 ( .A(n50522), .X(n50523) );
  inv_x2_sg U56757 ( .A(n50524), .X(n50525) );
  inv_x2_sg U56758 ( .A(n50526), .X(n50527) );
  inv_x2_sg U56759 ( .A(n50528), .X(n50529) );
  inv_x2_sg U56760 ( .A(n50530), .X(n50531) );
  inv_x2_sg U56761 ( .A(n50532), .X(n50533) );
  inv_x2_sg U56762 ( .A(n50534), .X(n50535) );
  inv_x2_sg U56763 ( .A(n50536), .X(n50537) );
  inv_x2_sg U56764 ( .A(n50538), .X(n50539) );
  inv_x2_sg U56765 ( .A(n50540), .X(n50541) );
  inv_x2_sg U56766 ( .A(n50542), .X(n50543) );
  inv_x2_sg U56767 ( .A(n50544), .X(n50545) );
  inv_x2_sg U56768 ( .A(n50546), .X(n50547) );
  inv_x2_sg U56769 ( .A(n50548), .X(n50549) );
  inv_x2_sg U56770 ( .A(n50550), .X(n50551) );
  inv_x2_sg U56771 ( .A(n50552), .X(n50553) );
  inv_x2_sg U56772 ( .A(n50554), .X(n50555) );
  inv_x2_sg U56773 ( .A(n50556), .X(n50557) );
  inv_x2_sg U56774 ( .A(n50558), .X(n50559) );
  inv_x2_sg U56775 ( .A(n50560), .X(n50561) );
  inv_x2_sg U56776 ( .A(n50562), .X(n50563) );
  inv_x2_sg U56777 ( .A(n50564), .X(n50565) );
  inv_x2_sg U56778 ( .A(n50566), .X(n50567) );
  inv_x2_sg U56779 ( .A(n50568), .X(n50569) );
  inv_x2_sg U56780 ( .A(n50570), .X(n50571) );
  inv_x2_sg U56781 ( .A(n50572), .X(n50573) );
  inv_x2_sg U56782 ( .A(n50574), .X(n50575) );
  inv_x2_sg U56783 ( .A(n50576), .X(n50577) );
  inv_x2_sg U56784 ( .A(n50578), .X(n50579) );
  inv_x2_sg U56785 ( .A(n50580), .X(n50581) );
  inv_x2_sg U56786 ( .A(n50582), .X(n50583) );
  inv_x2_sg U56787 ( .A(n50584), .X(n50585) );
  inv_x2_sg U56788 ( .A(n50586), .X(n50587) );
  inv_x2_sg U56789 ( .A(n50588), .X(n50589) );
  inv_x2_sg U56790 ( .A(n50590), .X(n50591) );
  inv_x2_sg U56791 ( .A(n50592), .X(n50593) );
  inv_x2_sg U56792 ( .A(n50594), .X(n50595) );
  inv_x2_sg U56793 ( .A(n50596), .X(n50597) );
  inv_x2_sg U56794 ( .A(n50598), .X(n50599) );
  inv_x2_sg U56795 ( .A(n50600), .X(n50601) );
  inv_x2_sg U56796 ( .A(n50602), .X(n50603) );
  inv_x2_sg U56797 ( .A(n50604), .X(n50605) );
  inv_x2_sg U56798 ( .A(n50606), .X(n50607) );
  inv_x2_sg U56799 ( .A(n50608), .X(n50609) );
  inv_x2_sg U56800 ( .A(n50610), .X(n50611) );
  inv_x2_sg U56801 ( .A(n50612), .X(n50613) );
  inv_x2_sg U56802 ( .A(n50614), .X(n50615) );
  inv_x2_sg U56803 ( .A(n50616), .X(n50617) );
  inv_x2_sg U56804 ( .A(n50618), .X(n50619) );
  inv_x2_sg U56805 ( .A(n50620), .X(n50621) );
  inv_x2_sg U56806 ( .A(n50622), .X(n50623) );
  inv_x2_sg U56807 ( .A(n50624), .X(n50625) );
  inv_x2_sg U56808 ( .A(n50626), .X(n50627) );
  inv_x2_sg U56809 ( .A(n50628), .X(n50629) );
  inv_x2_sg U56810 ( .A(n50630), .X(n50631) );
  inv_x2_sg U56811 ( .A(n50632), .X(n50633) );
  inv_x2_sg U56812 ( .A(n50634), .X(n50635) );
  inv_x2_sg U56813 ( .A(n50636), .X(n50637) );
  inv_x2_sg U56814 ( .A(n50638), .X(n50639) );
  inv_x2_sg U56815 ( .A(n50640), .X(n50641) );
  inv_x2_sg U56816 ( .A(n50642), .X(n50643) );
  inv_x2_sg U56817 ( .A(n50644), .X(n50645) );
  inv_x2_sg U56818 ( .A(n50646), .X(n50647) );
  inv_x2_sg U56819 ( .A(n50648), .X(n50649) );
  inv_x2_sg U56820 ( .A(n50650), .X(n50651) );
  inv_x2_sg U56821 ( .A(n50652), .X(n50653) );
  inv_x2_sg U56822 ( .A(n50654), .X(n50655) );
  inv_x2_sg U56823 ( .A(n50656), .X(n50657) );
  inv_x2_sg U56824 ( .A(n50658), .X(n50659) );
  inv_x2_sg U56825 ( .A(n50660), .X(n50661) );
  inv_x2_sg U56826 ( .A(n50662), .X(n50663) );
  inv_x2_sg U56827 ( .A(n50664), .X(n50665) );
  inv_x2_sg U56828 ( .A(n50666), .X(n50667) );
  inv_x2_sg U56829 ( .A(n50668), .X(n50669) );
  inv_x2_sg U56830 ( .A(n50670), .X(n50671) );
  inv_x2_sg U56831 ( .A(n50672), .X(n50673) );
  inv_x2_sg U56832 ( .A(n50674), .X(n50675) );
  inv_x2_sg U56833 ( .A(n50676), .X(n50677) );
  inv_x2_sg U56834 ( .A(n50678), .X(n50679) );
  inv_x2_sg U56835 ( .A(n50680), .X(n50681) );
  inv_x2_sg U56836 ( .A(n50682), .X(n50683) );
  inv_x2_sg U56837 ( .A(n50684), .X(n50685) );
  inv_x2_sg U56838 ( .A(n50686), .X(n50687) );
  inv_x2_sg U56839 ( .A(n50688), .X(n50689) );
  inv_x2_sg U56840 ( .A(n50690), .X(n50691) );
  inv_x2_sg U56841 ( .A(n50692), .X(n50693) );
  inv_x2_sg U56842 ( .A(n50694), .X(n50695) );
  inv_x2_sg U56843 ( .A(n50696), .X(n50697) );
  inv_x2_sg U56844 ( .A(n50698), .X(n50699) );
  inv_x2_sg U56845 ( .A(n50700), .X(n50701) );
  inv_x2_sg U56846 ( .A(n50702), .X(n50703) );
  inv_x2_sg U56847 ( .A(n50704), .X(n50705) );
  inv_x2_sg U56848 ( .A(n50706), .X(n50707) );
  inv_x2_sg U56849 ( .A(n50708), .X(n50709) );
  inv_x2_sg U56850 ( .A(n50710), .X(n50711) );
  inv_x2_sg U56851 ( .A(n50712), .X(n50713) );
  inv_x2_sg U56852 ( .A(n50714), .X(n50715) );
  inv_x2_sg U56853 ( .A(n50716), .X(n50717) );
  inv_x2_sg U56854 ( .A(n50718), .X(n50719) );
  inv_x2_sg U56855 ( .A(n50720), .X(n50721) );
  inv_x2_sg U56856 ( .A(n50722), .X(n50723) );
  inv_x2_sg U56857 ( .A(n50724), .X(n50725) );
  inv_x2_sg U56858 ( .A(n50726), .X(n50727) );
  inv_x2_sg U56859 ( .A(n50728), .X(n50729) );
  inv_x2_sg U56860 ( .A(n50730), .X(n50731) );
  inv_x2_sg U56861 ( .A(n50732), .X(n50733) );
  inv_x2_sg U56862 ( .A(n50734), .X(n50735) );
  inv_x2_sg U56863 ( .A(n50736), .X(n50737) );
  inv_x2_sg U56864 ( .A(n50738), .X(n50739) );
  inv_x2_sg U56865 ( .A(n50740), .X(n50741) );
  inv_x2_sg U56866 ( .A(n50742), .X(n50743) );
  inv_x2_sg U56867 ( .A(n50744), .X(n50745) );
  inv_x2_sg U56868 ( .A(n50746), .X(n50747) );
  inv_x2_sg U56869 ( .A(n50748), .X(n50749) );
  inv_x2_sg U56870 ( .A(n50750), .X(n50751) );
  inv_x2_sg U56871 ( .A(n50752), .X(n50753) );
  inv_x2_sg U56872 ( .A(n50754), .X(n50755) );
  inv_x2_sg U56873 ( .A(n50756), .X(n50757) );
  inv_x2_sg U56874 ( .A(n50758), .X(n50759) );
  inv_x2_sg U56875 ( .A(n50760), .X(n50761) );
  inv_x2_sg U56876 ( .A(n50762), .X(n50763) );
  inv_x2_sg U56877 ( .A(n50764), .X(n50765) );
  inv_x2_sg U56878 ( .A(n50766), .X(n50767) );
  inv_x2_sg U56879 ( .A(n50768), .X(n50769) );
  inv_x2_sg U56880 ( .A(n50770), .X(n50771) );
  inv_x2_sg U56881 ( .A(n50772), .X(n50773) );
  inv_x2_sg U56882 ( .A(n50774), .X(n50775) );
  inv_x2_sg U56883 ( .A(n50776), .X(n50777) );
  inv_x2_sg U56884 ( .A(n50778), .X(n50779) );
  inv_x2_sg U56885 ( .A(n50780), .X(n50781) );
  inv_x2_sg U56886 ( .A(n50782), .X(n50783) );
  inv_x2_sg U56887 ( .A(n50784), .X(n50785) );
  inv_x2_sg U56888 ( .A(n50786), .X(n50787) );
  inv_x2_sg U56889 ( .A(n50788), .X(n50789) );
  inv_x2_sg U56890 ( .A(n50790), .X(n50791) );
  inv_x2_sg U56891 ( .A(n50792), .X(n50793) );
  inv_x2_sg U56892 ( .A(n50794), .X(n50795) );
  inv_x2_sg U56893 ( .A(n50796), .X(n50797) );
  inv_x2_sg U56894 ( .A(n50798), .X(n50799) );
  inv_x2_sg U56895 ( .A(n50800), .X(n50801) );
  inv_x2_sg U56896 ( .A(n50802), .X(n50803) );
  inv_x2_sg U56897 ( .A(n50804), .X(n50805) );
  inv_x2_sg U56898 ( .A(n50806), .X(n50807) );
  inv_x2_sg U56899 ( .A(n50808), .X(n50809) );
  inv_x2_sg U56900 ( .A(n50810), .X(n50811) );
  inv_x2_sg U56901 ( .A(n50812), .X(n50813) );
  inv_x2_sg U56902 ( .A(n50814), .X(n50815) );
  inv_x2_sg U56903 ( .A(n50816), .X(n50817) );
  inv_x2_sg U56904 ( .A(n50818), .X(n50819) );
  inv_x2_sg U56905 ( .A(n50820), .X(n50821) );
  inv_x2_sg U56906 ( .A(n50822), .X(n50823) );
  inv_x2_sg U56907 ( .A(n50824), .X(n50825) );
  inv_x2_sg U56908 ( .A(n50826), .X(n50827) );
  inv_x2_sg U56909 ( .A(n50828), .X(n50829) );
  inv_x2_sg U56910 ( .A(n50830), .X(n50831) );
  inv_x2_sg U56911 ( .A(n50832), .X(n50833) );
  inv_x2_sg U56912 ( .A(n50834), .X(n50835) );
  inv_x2_sg U56913 ( .A(n50836), .X(n50837) );
  inv_x2_sg U56914 ( .A(n50838), .X(n50839) );
  inv_x2_sg U56915 ( .A(n50840), .X(n50841) );
  inv_x2_sg U56916 ( .A(n50842), .X(n50843) );
  inv_x2_sg U56917 ( .A(n50844), .X(n50845) );
  inv_x2_sg U56918 ( .A(n50846), .X(n50847) );
  inv_x2_sg U56919 ( .A(n50848), .X(n50849) );
  inv_x2_sg U56920 ( .A(n50850), .X(n50851) );
  inv_x2_sg U56921 ( .A(n50852), .X(n50853) );
  inv_x2_sg U56922 ( .A(n50854), .X(n50855) );
  inv_x2_sg U56923 ( .A(n50856), .X(n50857) );
  inv_x2_sg U56924 ( .A(n50858), .X(n50859) );
  inv_x2_sg U56925 ( .A(n50860), .X(n50861) );
  inv_x2_sg U56926 ( .A(n50862), .X(n50863) );
  inv_x2_sg U56927 ( .A(n50864), .X(n50865) );
  inv_x2_sg U56928 ( .A(n50866), .X(n50867) );
  inv_x2_sg U56929 ( .A(n50868), .X(n50869) );
  inv_x2_sg U56930 ( .A(n50870), .X(n50871) );
  inv_x2_sg U56931 ( .A(n50872), .X(n50873) );
  inv_x2_sg U56932 ( .A(n50874), .X(n50875) );
  inv_x2_sg U56933 ( .A(n50876), .X(n50877) );
  inv_x2_sg U56934 ( .A(n50878), .X(n50879) );
  inv_x2_sg U56935 ( .A(n50880), .X(n50881) );
  inv_x2_sg U56936 ( .A(n50882), .X(n50883) );
  inv_x2_sg U56937 ( .A(n50884), .X(n50885) );
  inv_x2_sg U56938 ( .A(n50886), .X(n50887) );
  inv_x2_sg U56939 ( .A(n50888), .X(n50889) );
  inv_x2_sg U56940 ( .A(n50890), .X(n50891) );
  inv_x2_sg U56941 ( .A(n50892), .X(n50893) );
  inv_x2_sg U56942 ( .A(n50894), .X(n50895) );
  inv_x2_sg U56943 ( .A(n50896), .X(n50897) );
  inv_x2_sg U56944 ( .A(n50898), .X(n50899) );
  inv_x2_sg U56945 ( .A(n50900), .X(n50901) );
  inv_x2_sg U56946 ( .A(n50902), .X(n50903) );
  inv_x2_sg U56947 ( .A(n50904), .X(n50905) );
  inv_x2_sg U56948 ( .A(n50906), .X(n50907) );
  inv_x2_sg U56949 ( .A(n50908), .X(n50909) );
  inv_x2_sg U56950 ( .A(n50910), .X(n50911) );
  inv_x2_sg U56951 ( .A(n50912), .X(n50913) );
  inv_x2_sg U56952 ( .A(n50914), .X(n50915) );
  inv_x2_sg U56953 ( .A(n50916), .X(n50917) );
  inv_x2_sg U56954 ( .A(n50918), .X(n50919) );
  inv_x2_sg U56955 ( .A(n50920), .X(n50921) );
  inv_x2_sg U56956 ( .A(n50922), .X(n50923) );
  inv_x2_sg U56957 ( .A(n50924), .X(n50925) );
  inv_x2_sg U56958 ( .A(n50926), .X(n50927) );
  inv_x2_sg U56959 ( .A(n50928), .X(n50929) );
  inv_x2_sg U56960 ( .A(n50930), .X(n50931) );
  inv_x2_sg U56961 ( .A(n50932), .X(n50933) );
  inv_x2_sg U56962 ( .A(n50934), .X(n50935) );
  inv_x2_sg U56963 ( .A(n50936), .X(n50937) );
  inv_x2_sg U56964 ( .A(n50938), .X(n50939) );
  inv_x2_sg U56965 ( .A(n50940), .X(n50941) );
  inv_x2_sg U56966 ( .A(n50942), .X(n50943) );
  inv_x2_sg U56967 ( .A(n50944), .X(n50945) );
  inv_x2_sg U56968 ( .A(n50946), .X(n50947) );
  inv_x2_sg U56969 ( .A(n50948), .X(n50949) );
  inv_x2_sg U56970 ( .A(n50950), .X(n50951) );
  inv_x2_sg U56971 ( .A(n50952), .X(n50953) );
  inv_x2_sg U56972 ( .A(n50954), .X(n50955) );
  inv_x2_sg U56973 ( .A(n50956), .X(n50957) );
  inv_x2_sg U56974 ( .A(n50958), .X(n50959) );
  inv_x2_sg U56975 ( .A(n50960), .X(n50961) );
  inv_x2_sg U56976 ( .A(n50962), .X(n50963) );
  inv_x2_sg U56977 ( .A(n50964), .X(n50965) );
  inv_x2_sg U56978 ( .A(n50966), .X(n50967) );
  inv_x2_sg U56979 ( .A(n50968), .X(n50969) );
  inv_x2_sg U56980 ( .A(n50970), .X(n50971) );
  inv_x2_sg U56981 ( .A(n50972), .X(n50973) );
  inv_x2_sg U56982 ( .A(n50974), .X(n50975) );
  inv_x2_sg U56983 ( .A(n50976), .X(n50977) );
  inv_x2_sg U56984 ( .A(n50978), .X(n50979) );
  inv_x2_sg U56985 ( .A(n50980), .X(n50981) );
  inv_x2_sg U56986 ( .A(n50982), .X(n50983) );
  inv_x2_sg U56987 ( .A(n50984), .X(n50985) );
  inv_x2_sg U56988 ( .A(n50986), .X(n50987) );
  inv_x2_sg U56989 ( .A(n50988), .X(n50989) );
  inv_x2_sg U56990 ( .A(n50990), .X(n50991) );
  inv_x2_sg U56991 ( .A(n50992), .X(n50993) );
  inv_x2_sg U56992 ( .A(n50994), .X(n50995) );
  inv_x2_sg U56993 ( .A(n50996), .X(n50997) );
  inv_x2_sg U56994 ( .A(n50998), .X(n50999) );
  inv_x2_sg U56995 ( .A(n51000), .X(n51001) );
  inv_x2_sg U56996 ( .A(n51002), .X(n51003) );
  inv_x2_sg U56997 ( .A(n51004), .X(n51005) );
  inv_x2_sg U56998 ( .A(n51006), .X(n51007) );
  inv_x2_sg U56999 ( .A(n51008), .X(n51009) );
  inv_x2_sg U57000 ( .A(n51010), .X(n51011) );
  inv_x2_sg U57001 ( .A(n51012), .X(n51013) );
  inv_x2_sg U57002 ( .A(n51014), .X(n51015) );
  inv_x2_sg U57003 ( .A(n51016), .X(n51017) );
  inv_x2_sg U57004 ( .A(n51018), .X(n51019) );
  inv_x2_sg U57005 ( .A(n51020), .X(n51021) );
  inv_x2_sg U57006 ( .A(n51022), .X(n51023) );
  inv_x2_sg U57007 ( .A(n51024), .X(n51025) );
  inv_x2_sg U57008 ( .A(n51026), .X(n51027) );
  inv_x2_sg U57009 ( .A(n51028), .X(n51029) );
  inv_x2_sg U57010 ( .A(n51030), .X(n51031) );
  inv_x2_sg U57011 ( .A(n51032), .X(n51033) );
  inv_x2_sg U57012 ( .A(n51034), .X(n51035) );
  inv_x2_sg U57013 ( .A(n51036), .X(n51037) );
  inv_x2_sg U57014 ( .A(n51038), .X(n51039) );
  inv_x2_sg U57015 ( .A(n51040), .X(n51041) );
  inv_x2_sg U57016 ( .A(n51042), .X(n51043) );
  inv_x2_sg U57017 ( .A(n51044), .X(n51045) );
  inv_x2_sg U57018 ( .A(n51046), .X(n51047) );
  inv_x2_sg U57019 ( .A(n51048), .X(n51049) );
  inv_x2_sg U57020 ( .A(n51050), .X(n51051) );
  inv_x4_sg U57021 ( .A(n22643), .X(n67376) );
  inv_x4_sg U57022 ( .A(n22642), .X(n67377) );
  inv_x4_sg U57023 ( .A(n22637), .X(n67382) );
  inv_x4_sg U57024 ( .A(n22635), .X(n67384) );
  inv_x4_sg U57025 ( .A(n22633), .X(n67386) );
  inv_x4_sg U57026 ( .A(n22631), .X(n67388) );
  inv_x4_sg U57027 ( .A(n22628), .X(n67391) );
  inv_x4_sg U57028 ( .A(n22627), .X(n67392) );
  inv_x4_sg U57029 ( .A(n22616), .X(n67163) );
  inv_x4_sg U57030 ( .A(n22615), .X(n67164) );
  inv_x4_sg U57031 ( .A(n22610), .X(n67169) );
  inv_x4_sg U57032 ( .A(n22608), .X(n67171) );
  inv_x4_sg U57033 ( .A(n22606), .X(n67173) );
  inv_x4_sg U57034 ( .A(n22604), .X(n67175) );
  inv_x4_sg U57035 ( .A(n22601), .X(n67178) );
  inv_x4_sg U57036 ( .A(n22600), .X(n67179) );
  inv_x4_sg U57037 ( .A(n51052), .X(n51053) );
  nor_x4_sg U57038 ( .A(n67530), .B(n56935), .X(n26092) );
  inv_x4_sg U57039 ( .A(n51056), .X(n51057) );
  nand_x8_sg U57040 ( .A(n57862), .B(n22467), .X(n22693) );
  inv_x4_sg U57041 ( .A(n51058), .X(n51059) );
  inv_x4_sg U57042 ( .A(n51060), .X(n51061) );
  inv_x4_sg U57043 ( .A(n51062), .X(n51063) );
  inv_x4_sg U57044 ( .A(n51064), .X(n51065) );
  inv_x4_sg U57045 ( .A(n51066), .X(n51067) );
  inv_x4_sg U57046 ( .A(n51068), .X(n51069) );
  nor_x8_sg U57047 ( .A(n68386), .B(n57168), .X(n34220) );
  nor_x8_sg U57048 ( .A(n68380), .B(n57168), .X(n33912) );
  inv_x4_sg U57049 ( .A(n51070), .X(n51071) );
  inv_x4_sg U57050 ( .A(n51072), .X(n51073) );
  inv_x4_sg U57051 ( .A(n51074), .X(n51075) );
  inv_x4_sg U57052 ( .A(n51076), .X(n51077) );
  inv_x4_sg U57053 ( .A(n51078), .X(n51079) );
  inv_x4_sg U57054 ( .A(n51080), .X(n51081) );
  inv_x4_sg U57055 ( .A(n51082), .X(n51083) );
  inv_x4_sg U57056 ( .A(n51084), .X(n51085) );
  inv_x4_sg U57057 ( .A(n51086), .X(n51087) );
  inv_x4_sg U57058 ( .A(n51088), .X(n51089) );
  inv_x4_sg U57059 ( .A(n51090), .X(n51091) );
  inv_x4_sg U57060 ( .A(n51092), .X(n51093) );
  inv_x4_sg U57061 ( .A(n51094), .X(n51095) );
  inv_x4_sg U57062 ( .A(n51096), .X(n51097) );
  inv_x4_sg U57063 ( .A(n51098), .X(n51099) );
  inv_x4_sg U57064 ( .A(n51100), .X(n51101) );
  inv_x4_sg U57065 ( .A(n51102), .X(n51103) );
  inv_x4_sg U57066 ( .A(n51104), .X(n51105) );
  inv_x4_sg U57067 ( .A(n51106), .X(n51107) );
  inv_x4_sg U57068 ( .A(n51108), .X(n51109) );
  inv_x4_sg U57069 ( .A(n51110), .X(n51111) );
  inv_x4_sg U57070 ( .A(n51112), .X(n51113) );
  inv_x4_sg U57071 ( .A(n51114), .X(n51115) );
  inv_x4_sg U57072 ( .A(n51116), .X(n51117) );
  inv_x4_sg U57073 ( .A(n51118), .X(n51119) );
  inv_x4_sg U57074 ( .A(n51120), .X(n51121) );
  inv_x4_sg U57075 ( .A(n51122), .X(n51123) );
  inv_x4_sg U57076 ( .A(n51124), .X(n51125) );
  inv_x4_sg U57077 ( .A(n51126), .X(n51127) );
  inv_x4_sg U57078 ( .A(n51128), .X(n51129) );
  inv_x4_sg U57079 ( .A(n51130), .X(n51131) );
  inv_x4_sg U57080 ( .A(n51132), .X(n51133) );
  nand_x8_sg U57081 ( .A(n58482), .B(n68587), .X(n22522) );
  nor_x4_sg U57082 ( .A(n32429), .B(n32535), .X(n32378) );
  nand_x4_sg U57083 ( .A(n32536), .B(n32537), .X(n32535) );
  inv_x8_sg U57084 ( .A(reset), .X(n61908) );
  inv_x4_sg U57085 ( .A(n58617), .X(n58655) );
  nand_x2_sg U57086 ( .A(n57455), .B(n58616), .X(n58617) );
  inv_x4_sg U57087 ( .A(n51134), .X(n51135) );
  inv_x4_sg U57088 ( .A(n51136), .X(n51137) );
  inv_x4_sg U57089 ( .A(n51138), .X(n51139) );
  inv_x4_sg U57090 ( .A(n51140), .X(n51141) );
  inv_x4_sg U57091 ( .A(n51142), .X(n51143) );
  inv_x4_sg U57092 ( .A(n51144), .X(n51145) );
  inv_x4_sg U57093 ( .A(n51146), .X(n51147) );
  inv_x4_sg U57094 ( .A(n51148), .X(n51149) );
  inv_x4_sg U57095 ( .A(n51150), .X(n51151) );
  inv_x4_sg U57096 ( .A(n51152), .X(n51153) );
  inv_x4_sg U57097 ( .A(n51154), .X(n51155) );
  inv_x4_sg U57098 ( .A(n51156), .X(n51157) );
  inv_x4_sg U57099 ( .A(n51158), .X(n51159) );
  inv_x4_sg U57100 ( .A(n51160), .X(n51161) );
  inv_x4_sg U57101 ( .A(n51162), .X(n51163) );
  inv_x4_sg U57102 ( .A(n51164), .X(n51165) );
  inv_x4_sg U57103 ( .A(n51166), .X(n51167) );
  inv_x4_sg U57104 ( .A(n51168), .X(n51169) );
  inv_x4_sg U57105 ( .A(n51170), .X(n51171) );
  inv_x4_sg U57106 ( .A(n51172), .X(n51173) );
  inv_x4_sg U57107 ( .A(n51174), .X(n51175) );
  inv_x4_sg U57108 ( .A(n51176), .X(n51177) );
  inv_x4_sg U57109 ( .A(n51178), .X(n51179) );
  inv_x4_sg U57110 ( .A(n51180), .X(n51181) );
  inv_x4_sg U57111 ( .A(n51182), .X(n51183) );
  inv_x4_sg U57112 ( .A(n51184), .X(n51185) );
  inv_x4_sg U57113 ( .A(n51186), .X(n51187) );
  inv_x4_sg U57114 ( .A(n51188), .X(n51189) );
  inv_x4_sg U57115 ( .A(n51190), .X(n51191) );
  inv_x4_sg U57116 ( .A(n51192), .X(n51193) );
  inv_x4_sg U57117 ( .A(n51194), .X(n51195) );
  inv_x4_sg U57118 ( .A(n51196), .X(n51197) );
  inv_x4_sg U57119 ( .A(n51198), .X(n51199) );
  nor_x8_sg U57120 ( .A(n67535), .B(n26304), .X(n26121) );
  inv_x8_sg U57121 ( .A(n57111), .X(n67535) );
  inv_x8_sg U57122 ( .A(n26051), .X(n67532) );
  inv_x8_sg U57123 ( .A(n58476), .X(n58479) );
  nand_x4_sg U57124 ( .A(n58479), .B(n58616), .X(n58480) );
  inv_x4_sg U57125 ( .A(n51200), .X(n51201) );
  inv_x4_sg U57126 ( .A(n51202), .X(n51203) );
  inv_x4_sg U57127 ( .A(n51204), .X(n51205) );
  inv_x4_sg U57128 ( .A(n51206), .X(n51207) );
  inv_x4_sg U57129 ( .A(n51208), .X(n51209) );
  inv_x4_sg U57130 ( .A(n51210), .X(n51211) );
  inv_x4_sg U57131 ( .A(n51212), .X(n51213) );
  inv_x4_sg U57132 ( .A(n51214), .X(n51215) );
  inv_x4_sg U57133 ( .A(n51216), .X(n51217) );
  inv_x4_sg U57134 ( .A(n51218), .X(n51219) );
  inv_x4_sg U57135 ( .A(n51220), .X(n51221) );
  inv_x4_sg U57136 ( .A(n51222), .X(n51223) );
  inv_x4_sg U57137 ( .A(n51224), .X(n51225) );
  inv_x4_sg U57138 ( .A(n51226), .X(n51227) );
  inv_x4_sg U57139 ( .A(n51228), .X(n51229) );
  inv_x4_sg U57140 ( .A(n51230), .X(n51231) );
  inv_x4_sg U57141 ( .A(n51232), .X(n51233) );
  inv_x4_sg U57142 ( .A(n51234), .X(n51235) );
  inv_x4_sg U57143 ( .A(n51236), .X(n51237) );
  inv_x4_sg U57144 ( .A(n51238), .X(n51239) );
  inv_x4_sg U57145 ( .A(n51240), .X(n51241) );
  inv_x4_sg U57146 ( .A(n51242), .X(n51243) );
  inv_x4_sg U57147 ( .A(n51244), .X(n51245) );
  inv_x4_sg U57148 ( .A(n51246), .X(n51247) );
  inv_x4_sg U57149 ( .A(n51248), .X(n51249) );
  inv_x4_sg U57150 ( .A(n51250), .X(n51251) );
  inv_x4_sg U57151 ( .A(n51252), .X(n51253) );
  inv_x4_sg U57152 ( .A(n51254), .X(n51255) );
  inv_x4_sg U57153 ( .A(n51256), .X(n51257) );
  inv_x4_sg U57154 ( .A(n51258), .X(n51259) );
  inv_x4_sg U57155 ( .A(n51260), .X(n51261) );
  inv_x4_sg U57156 ( .A(n51262), .X(n51263) );
  inv_x4_sg U57157 ( .A(n51264), .X(n51265) );
  inv_x4_sg U57158 ( .A(n51266), .X(n51267) );
  inv_x4_sg U57159 ( .A(n51268), .X(n51269) );
  inv_x4_sg U57160 ( .A(n51270), .X(n51271) );
  inv_x4_sg U57161 ( .A(n51272), .X(n51273) );
  inv_x4_sg U57162 ( .A(n51274), .X(n51275) );
  inv_x4_sg U57163 ( .A(n51276), .X(n51277) );
  inv_x4_sg U57164 ( .A(n51278), .X(n51279) );
  inv_x4_sg U57165 ( .A(n51280), .X(n51281) );
  inv_x4_sg U57166 ( .A(n51282), .X(n51283) );
  inv_x4_sg U57167 ( .A(n51284), .X(n51285) );
  inv_x4_sg U57168 ( .A(n51286), .X(n51287) );
  inv_x4_sg U57169 ( .A(n51288), .X(n51289) );
  inv_x4_sg U57170 ( .A(n51290), .X(n51291) );
  inv_x4_sg U57171 ( .A(n51292), .X(n51293) );
  inv_x4_sg U57172 ( .A(n51294), .X(n51295) );
  inv_x4_sg U57173 ( .A(n51296), .X(n51297) );
  inv_x4_sg U57174 ( .A(n51298), .X(n51299) );
  inv_x4_sg U57175 ( .A(n51300), .X(n51301) );
  inv_x4_sg U57176 ( .A(n51302), .X(n51303) );
  inv_x4_sg U57177 ( .A(n51304), .X(n51305) );
  inv_x4_sg U57178 ( .A(n51306), .X(n51307) );
  inv_x4_sg U57179 ( .A(n51308), .X(n51309) );
  inv_x4_sg U57180 ( .A(n51310), .X(n51311) );
  inv_x4_sg U57181 ( .A(n51312), .X(n51313) );
  inv_x4_sg U57182 ( .A(n51314), .X(n51315) );
  inv_x4_sg U57183 ( .A(n51316), .X(n51317) );
  inv_x4_sg U57184 ( .A(n51318), .X(n51319) );
  inv_x4_sg U57185 ( .A(n51320), .X(n51321) );
  inv_x4_sg U57186 ( .A(n51322), .X(n51323) );
  inv_x4_sg U57187 ( .A(n51324), .X(n51325) );
  inv_x4_sg U57188 ( .A(n51326), .X(n51327) );
  inv_x4_sg U57189 ( .A(n51328), .X(n51329) );
  inv_x4_sg U57190 ( .A(n51330), .X(n51331) );
  inv_x4_sg U57191 ( .A(n51332), .X(n51333) );
  inv_x4_sg U57192 ( .A(n51334), .X(n51335) );
  inv_x4_sg U57193 ( .A(n51336), .X(n51337) );
  inv_x4_sg U57194 ( .A(n51338), .X(n51339) );
  inv_x4_sg U57195 ( .A(n51340), .X(n51341) );
  inv_x4_sg U57196 ( .A(n51342), .X(n51343) );
  inv_x4_sg U57197 ( .A(n51344), .X(n51345) );
  inv_x4_sg U57198 ( .A(n51346), .X(n51347) );
  inv_x4_sg U57199 ( .A(n51348), .X(n51349) );
  inv_x4_sg U57200 ( .A(n51350), .X(n51351) );
  inv_x4_sg U57201 ( .A(n51352), .X(n51353) );
  inv_x4_sg U57202 ( .A(n51354), .X(n51355) );
  inv_x4_sg U57203 ( .A(n51356), .X(n51357) );
  inv_x4_sg U57204 ( .A(n51358), .X(n51359) );
  inv_x4_sg U57205 ( .A(n51360), .X(n51361) );
  inv_x4_sg U57206 ( .A(n51362), .X(n51363) );
  inv_x4_sg U57207 ( .A(n51364), .X(n51365) );
  inv_x4_sg U57208 ( .A(n51366), .X(n51367) );
  inv_x4_sg U57209 ( .A(n51368), .X(n51369) );
  inv_x4_sg U57210 ( .A(n51370), .X(n51371) );
  inv_x4_sg U57211 ( .A(n51372), .X(n51373) );
  inv_x4_sg U57212 ( .A(n51374), .X(n51375) );
  inv_x4_sg U57213 ( .A(n51376), .X(n51377) );
  inv_x4_sg U57214 ( .A(n51378), .X(n51379) );
  inv_x4_sg U57215 ( .A(n51380), .X(n51381) );
  inv_x4_sg U57216 ( .A(n51382), .X(n51383) );
  inv_x4_sg U57217 ( .A(n51384), .X(n51385) );
  inv_x4_sg U57218 ( .A(n51386), .X(n51387) );
  inv_x4_sg U57219 ( .A(n51388), .X(n51389) );
  inv_x4_sg U57220 ( .A(n51390), .X(n51391) );
  inv_x4_sg U57221 ( .A(n51392), .X(n51393) );
  inv_x4_sg U57222 ( .A(n51394), .X(n51395) );
  inv_x4_sg U57223 ( .A(n51396), .X(n51397) );
  inv_x4_sg U57224 ( .A(n51398), .X(n51399) );
  inv_x4_sg U57225 ( .A(n51400), .X(n51401) );
  inv_x4_sg U57226 ( .A(n51402), .X(n51403) );
  inv_x4_sg U57227 ( .A(n51404), .X(n51405) );
  inv_x4_sg U57228 ( .A(n51406), .X(n51407) );
  inv_x4_sg U57229 ( .A(n51408), .X(n51409) );
  inv_x4_sg U57230 ( .A(n51410), .X(n51411) );
  inv_x4_sg U57231 ( .A(n51412), .X(n51413) );
  inv_x4_sg U57232 ( .A(n51414), .X(n51415) );
  inv_x4_sg U57233 ( .A(n51416), .X(n51417) );
  inv_x4_sg U57234 ( .A(n51418), .X(n51419) );
  inv_x4_sg U57235 ( .A(n51420), .X(n51421) );
  inv_x4_sg U57236 ( .A(n51422), .X(n51423) );
  inv_x4_sg U57237 ( .A(n51424), .X(n51425) );
  inv_x4_sg U57238 ( .A(n51426), .X(n51427) );
  inv_x4_sg U57239 ( .A(n51428), .X(n51429) );
  inv_x4_sg U57240 ( .A(n51430), .X(n51431) );
  inv_x4_sg U57241 ( .A(n51432), .X(n51433) );
  inv_x4_sg U57242 ( .A(n51434), .X(n51435) );
  inv_x4_sg U57243 ( .A(n51436), .X(n51437) );
  inv_x4_sg U57244 ( .A(n51438), .X(n51439) );
  inv_x4_sg U57245 ( .A(n51440), .X(n51441) );
  inv_x4_sg U57246 ( .A(n51442), .X(n51443) );
  inv_x4_sg U57247 ( .A(n51444), .X(n51445) );
  inv_x4_sg U57248 ( .A(n51446), .X(n51447) );
  inv_x4_sg U57249 ( .A(n51448), .X(n51449) );
  inv_x4_sg U57250 ( .A(n51450), .X(n51451) );
  inv_x4_sg U57251 ( .A(n51452), .X(n51453) );
  inv_x4_sg U57252 ( .A(n51454), .X(n51455) );
  inv_x4_sg U57253 ( .A(n51456), .X(n51457) );
  inv_x4_sg U57254 ( .A(n51458), .X(n51459) );
  inv_x4_sg U57255 ( .A(n51460), .X(n51461) );
  inv_x4_sg U57256 ( .A(n51462), .X(n51463) );
  inv_x4_sg U57257 ( .A(n51464), .X(n51465) );
  inv_x4_sg U57258 ( .A(n51466), .X(n51467) );
  inv_x4_sg U57259 ( .A(n51468), .X(n51469) );
  inv_x4_sg U57260 ( .A(n51470), .X(n51471) );
  inv_x4_sg U57261 ( .A(n51472), .X(n51473) );
  inv_x4_sg U57262 ( .A(n51474), .X(n51475) );
  inv_x4_sg U57263 ( .A(n51476), .X(n51477) );
  inv_x4_sg U57264 ( .A(n51478), .X(n51479) );
  inv_x4_sg U57265 ( .A(n51480), .X(n51481) );
  inv_x4_sg U57266 ( .A(n51482), .X(n51483) );
  inv_x4_sg U57267 ( .A(n51484), .X(n51485) );
  inv_x4_sg U57268 ( .A(n51486), .X(n51487) );
  inv_x4_sg U57269 ( .A(n46973), .X(n51488) );
  inv_x8_sg U57270 ( .A(n51488), .X(n51489) );
  inv_x4_sg U57271 ( .A(n46965), .X(n51490) );
  inv_x8_sg U57272 ( .A(n51490), .X(n51491) );
  inv_x4_sg U57273 ( .A(n46971), .X(n51492) );
  inv_x8_sg U57274 ( .A(n51492), .X(n51493) );
  inv_x4_sg U57275 ( .A(n47117), .X(n51494) );
  inv_x8_sg U57276 ( .A(n51494), .X(n51495) );
  inv_x4_sg U57277 ( .A(n47109), .X(n51496) );
  inv_x8_sg U57278 ( .A(n51496), .X(n51497) );
  inv_x4_sg U57279 ( .A(n47101), .X(n51498) );
  inv_x8_sg U57280 ( .A(n51498), .X(n51499) );
  inv_x4_sg U57281 ( .A(n47091), .X(n51500) );
  inv_x8_sg U57282 ( .A(n51500), .X(n51501) );
  inv_x4_sg U57283 ( .A(n46957), .X(n51502) );
  inv_x8_sg U57284 ( .A(n51502), .X(n51503) );
  inv_x4_sg U57285 ( .A(n46947), .X(n51504) );
  inv_x8_sg U57286 ( .A(n51504), .X(n51505) );
  inv_x4_sg U57287 ( .A(n47115), .X(n51506) );
  inv_x8_sg U57288 ( .A(n51506), .X(n51507) );
  inv_x4_sg U57289 ( .A(n47105), .X(n51508) );
  inv_x8_sg U57290 ( .A(n51508), .X(n51509) );
  inv_x4_sg U57291 ( .A(n47097), .X(n51510) );
  inv_x8_sg U57292 ( .A(n51510), .X(n51511) );
  inv_x4_sg U57293 ( .A(n47087), .X(n51512) );
  inv_x8_sg U57294 ( .A(n51512), .X(n51513) );
  inv_x4_sg U57295 ( .A(n46961), .X(n51514) );
  inv_x8_sg U57296 ( .A(n51514), .X(n51515) );
  inv_x4_sg U57297 ( .A(n46953), .X(n51516) );
  inv_x8_sg U57298 ( .A(n51516), .X(n51517) );
  inv_x4_sg U57299 ( .A(n46943), .X(n51518) );
  inv_x8_sg U57300 ( .A(n51518), .X(n51519) );
  inv_x4_sg U57301 ( .A(n47287), .X(n51520) );
  inv_x8_sg U57302 ( .A(n51520), .X(state[1]) );
  inv_x8_sg U57303 ( .A(n58612), .X(n61910) );
  inv_x4_sg U57304 ( .A(n47201), .X(n51522) );
  inv_x8_sg U57305 ( .A(n51522), .X(n51523) );
  inv_x8_sg U57306 ( .A(n51523), .X(n68380) );
  inv_x4_sg U57307 ( .A(n47193), .X(n51524) );
  inv_x8_sg U57308 ( .A(n51524), .X(n51525) );
  inv_x8_sg U57309 ( .A(n51525), .X(n68386) );
  inv_x4_sg U57310 ( .A(n47157), .X(n51526) );
  inv_x8_sg U57311 ( .A(n51526), .X(n51527) );
  inv_x4_sg U57312 ( .A(n47149), .X(n51528) );
  inv_x8_sg U57313 ( .A(n51528), .X(n51529) );
  inv_x4_sg U57314 ( .A(n47141), .X(n51530) );
  inv_x8_sg U57315 ( .A(n51530), .X(n51531) );
  inv_x4_sg U57316 ( .A(n47133), .X(n51532) );
  inv_x8_sg U57317 ( .A(n51532), .X(n51533) );
  inv_x4_sg U57318 ( .A(n47013), .X(n51534) );
  inv_x8_sg U57319 ( .A(n51534), .X(n51535) );
  inv_x4_sg U57320 ( .A(n47005), .X(n51536) );
  inv_x8_sg U57321 ( .A(n51536), .X(n51537) );
  inv_x4_sg U57322 ( .A(n46997), .X(n51538) );
  inv_x8_sg U57323 ( .A(n51538), .X(n51539) );
  inv_x4_sg U57324 ( .A(n46989), .X(n51540) );
  inv_x8_sg U57325 ( .A(n51540), .X(n51541) );
  inv_x4_sg U57326 ( .A(n47043), .X(n51542) );
  inv_x8_sg U57327 ( .A(n51542), .X(n51543) );
  inv_x4_sg U57328 ( .A(n46925), .X(n51544) );
  inv_x8_sg U57329 ( .A(n51544), .X(n51545) );
  inv_x4_sg U57330 ( .A(n47073), .X(n51546) );
  inv_x8_sg U57331 ( .A(n51546), .X(n51547) );
  inv_x4_sg U57332 ( .A(n46897), .X(n51548) );
  inv_x8_sg U57333 ( .A(n51548), .X(n51549) );
  inv_x4_sg U57334 ( .A(n47055), .X(n51550) );
  inv_x8_sg U57335 ( .A(n51550), .X(n51551) );
  inv_x4_sg U57336 ( .A(n46907), .X(n51552) );
  inv_x8_sg U57337 ( .A(n51552), .X(n51553) );
  inv_x8_sg U57338 ( .A(n33395), .X(n68231) );
  nand_x4_sg U57339 ( .A(n33396), .B(n33397), .X(n33395) );
  inv_x2_sg U57340 ( .A(n51554), .X(n51555) );
  inv_x8_sg U57341 ( .A(n38411), .X(n68227) );
  inv_x8_sg U57342 ( .A(state[0]), .X(n68272) );
  nor_x1_sg U57343 ( .A(n32417), .B(n32418), .X(n32392) );
  nor_x1_sg U57344 ( .A(n31949), .B(n31950), .X(n31924) );
  inv_x4_sg U57345 ( .A(n25570), .X(n67469) );
  inv_x4_sg U57346 ( .A(n25420), .X(n67474) );
  inv_x4_sg U57347 ( .A(n24816), .X(n67281) );
  nand_x4_sg U57348 ( .A(n68228), .B(n33094), .X(n34002) );
  inv_x8_sg U57349 ( .A(n34041), .X(n68228) );
  nand_x4_sg U57350 ( .A(n33955), .B(n33310), .X(n34180) );
  nor_x8_sg U57351 ( .A(n34087), .B(n34220), .X(n33955) );
  nand_x4_sg U57352 ( .A(n33265), .B(n32965), .X(n33872) );
  nor_x8_sg U57353 ( .A(n33911), .B(n33912), .X(n33265) );
  nand_x4_sg U57354 ( .A(n68229), .B(n33008), .X(n33742) );
  inv_x8_sg U57355 ( .A(n33781), .X(n68229) );
  inv_x4_sg U57356 ( .A(n24154), .X(n67501) );
  inv_x4_sg U57357 ( .A(n24044), .X(n67098) );
  nor_x4_sg U57358 ( .A(n57917), .B(n57949), .X(n58387) );
  inv_x4_sg U57359 ( .A(n58581), .X(n29329) );
  nand_x8_sg U57360 ( .A(n67530), .B(n67534), .X(n26303) );
  inv_x4_sg U57361 ( .A(n22591), .X(n67356) );
  inv_x4_sg U57362 ( .A(n22565), .X(n67143) );
  inv_x4_sg U57363 ( .A(n22541), .X(n67337) );
  inv_x4_sg U57364 ( .A(n22538), .X(n67340) );
  inv_x4_sg U57365 ( .A(n22536), .X(n67342) );
  inv_x4_sg U57366 ( .A(n22534), .X(n67344) );
  inv_x4_sg U57367 ( .A(n22532), .X(n67346) );
  inv_x4_sg U57368 ( .A(n22530), .X(n67348) );
  inv_x4_sg U57369 ( .A(n22529), .X(n67349) );
  inv_x4_sg U57370 ( .A(n22527), .X(n67351) );
  inv_x4_sg U57371 ( .A(n22526), .X(n67352) );
  inv_x4_sg U57372 ( .A(n22525), .X(n67353) );
  inv_x4_sg U57373 ( .A(n22524), .X(n67354) );
  inv_x4_sg U57374 ( .A(n22516), .X(n67124) );
  inv_x4_sg U57375 ( .A(n22513), .X(n67127) );
  inv_x4_sg U57376 ( .A(n22511), .X(n67129) );
  inv_x4_sg U57377 ( .A(n22509), .X(n67131) );
  inv_x4_sg U57378 ( .A(n22507), .X(n67133) );
  inv_x4_sg U57379 ( .A(n22505), .X(n67135) );
  inv_x4_sg U57380 ( .A(n22504), .X(n67136) );
  inv_x4_sg U57381 ( .A(n22502), .X(n67138) );
  inv_x4_sg U57382 ( .A(n22501), .X(n67139) );
  inv_x4_sg U57383 ( .A(n22499), .X(n67141) );
  inv_x4_sg U57384 ( .A(n22448), .X(n67120) );
  inv_x4_sg U57385 ( .A(n22439), .X(n61899) );
  inv_x4_sg U57386 ( .A(n22438), .X(n61898) );
  inv_x4_sg U57387 ( .A(n22436), .X(n61896) );
  inv_x4_sg U57388 ( .A(n22434), .X(n61894) );
  inv_x4_sg U57389 ( .A(n22432), .X(n61892) );
  inv_x4_sg U57390 ( .A(n22430), .X(n61890) );
  inv_x4_sg U57391 ( .A(n22428), .X(n61888) );
  inv_x4_sg U57392 ( .A(n22427), .X(n61887) );
  inv_x4_sg U57393 ( .A(n22425), .X(n61885) );
  inv_x4_sg U57394 ( .A(n22424), .X(n61884) );
  inv_x4_sg U57395 ( .A(n22423), .X(n61883) );
  inv_x4_sg U57396 ( .A(n22422), .X(n61882) );
  inv_x4_sg U57397 ( .A(n22414), .X(n61879) );
  inv_x4_sg U57398 ( .A(n22413), .X(n61878) );
  inv_x4_sg U57399 ( .A(n22411), .X(n61876) );
  inv_x4_sg U57400 ( .A(n22409), .X(n61874) );
  inv_x4_sg U57401 ( .A(n22407), .X(n61872) );
  inv_x4_sg U57402 ( .A(n22405), .X(n61870) );
  inv_x4_sg U57403 ( .A(n22403), .X(n61868) );
  inv_x4_sg U57404 ( .A(n22402), .X(n61867) );
  inv_x4_sg U57405 ( .A(n22400), .X(n61865) );
  inv_x4_sg U57406 ( .A(n22399), .X(n61864) );
  inv_x4_sg U57407 ( .A(n22397), .X(n61862) );
  inv_x2_sg U57408 ( .A(n51558), .X(input_taken) );
  inv_x2_sg U57409 ( .A(n51560), .X(n51561) );
  inv_x2_sg U57410 ( .A(n51562), .X(n51563) );
  inv_x2_sg U57411 ( .A(n51564), .X(n51565) );
  inv_x2_sg U57412 ( .A(n51566), .X(n51567) );
  inv_x2_sg U57413 ( .A(n51568), .X(n51569) );
  inv_x2_sg U57414 ( .A(n51570), .X(n51571) );
  inv_x2_sg U57415 ( .A(n51572), .X(n51573) );
  inv_x2_sg U57416 ( .A(n51574), .X(n51575) );
  inv_x2_sg U57417 ( .A(n51576), .X(n51577) );
  inv_x2_sg U57418 ( .A(n51578), .X(n51579) );
  inv_x2_sg U57419 ( .A(n51580), .X(n51581) );
  inv_x2_sg U57420 ( .A(n51582), .X(n51583) );
  inv_x2_sg U57421 ( .A(n51584), .X(n51585) );
  inv_x2_sg U57422 ( .A(n51586), .X(n51587) );
  inv_x2_sg U57423 ( .A(n51588), .X(n51589) );
  inv_x2_sg U57424 ( .A(n51590), .X(n51591) );
  inv_x2_sg U57425 ( .A(n51592), .X(n51593) );
  inv_x2_sg U57426 ( .A(n51594), .X(n51595) );
  inv_x2_sg U57427 ( .A(n51596), .X(n51597) );
  inv_x2_sg U57428 ( .A(n51598), .X(n51599) );
  inv_x2_sg U57429 ( .A(n51600), .X(n51601) );
  inv_x2_sg U57430 ( .A(n51602), .X(n51603) );
  inv_x2_sg U57431 ( .A(n51604), .X(n51605) );
  inv_x2_sg U57432 ( .A(n51606), .X(n51607) );
  inv_x2_sg U57433 ( .A(n51608), .X(n51609) );
  inv_x2_sg U57434 ( .A(n51610), .X(n51611) );
  inv_x2_sg U57435 ( .A(n51612), .X(n51613) );
  inv_x2_sg U57436 ( .A(n51614), .X(n51615) );
  inv_x2_sg U57437 ( .A(n51616), .X(n51617) );
  inv_x2_sg U57438 ( .A(n51618), .X(n51619) );
  inv_x2_sg U57439 ( .A(n51620), .X(n51621) );
  inv_x2_sg U57440 ( .A(n51622), .X(n51623) );
  inv_x2_sg U57441 ( .A(n51624), .X(n51625) );
  inv_x2_sg U57442 ( .A(n51626), .X(n51627) );
  inv_x2_sg U57443 ( .A(n51628), .X(n51629) );
  inv_x2_sg U57444 ( .A(n51630), .X(n51631) );
  inv_x2_sg U57445 ( .A(n51632), .X(n51633) );
  inv_x2_sg U57446 ( .A(n51634), .X(n51635) );
  inv_x2_sg U57447 ( .A(n51636), .X(n51637) );
  inv_x2_sg U57448 ( .A(n51638), .X(n51639) );
  inv_x2_sg U57449 ( .A(n51640), .X(n51641) );
  inv_x2_sg U57450 ( .A(n51642), .X(n51643) );
  inv_x2_sg U57451 ( .A(n51644), .X(n51645) );
  inv_x2_sg U57452 ( .A(n51646), .X(n51647) );
  inv_x2_sg U57453 ( .A(n51648), .X(n51649) );
  inv_x2_sg U57454 ( .A(n51650), .X(n51651) );
  inv_x2_sg U57455 ( .A(n51652), .X(n51653) );
  inv_x2_sg U57456 ( .A(n51654), .X(n51655) );
  inv_x2_sg U57457 ( .A(n51656), .X(n51657) );
  inv_x2_sg U57458 ( .A(n51658), .X(n51659) );
  inv_x2_sg U57459 ( .A(n51660), .X(n51661) );
  inv_x2_sg U57460 ( .A(n51662), .X(n51663) );
  inv_x2_sg U57461 ( .A(n51664), .X(n51665) );
  inv_x2_sg U57462 ( .A(n51666), .X(n51667) );
  inv_x2_sg U57463 ( .A(n51668), .X(n51669) );
  inv_x2_sg U57464 ( .A(n51670), .X(n51671) );
  inv_x2_sg U57465 ( .A(n51672), .X(n51673) );
  inv_x2_sg U57466 ( .A(n51674), .X(n51675) );
  inv_x2_sg U57467 ( .A(n51676), .X(n51677) );
  inv_x2_sg U57468 ( .A(n51678), .X(n51679) );
  inv_x2_sg U57469 ( .A(n51680), .X(n51681) );
  inv_x2_sg U57470 ( .A(n51682), .X(n51683) );
  inv_x2_sg U57471 ( .A(n51684), .X(n51685) );
  inv_x2_sg U57472 ( .A(n51686), .X(n51687) );
  inv_x2_sg U57473 ( .A(n51688), .X(n51689) );
  inv_x2_sg U57474 ( .A(n51690), .X(n51691) );
  inv_x2_sg U57475 ( .A(n51692), .X(n51693) );
  inv_x2_sg U57476 ( .A(n51694), .X(n51695) );
  inv_x2_sg U57477 ( .A(n51696), .X(n51697) );
  inv_x2_sg U57478 ( .A(n51698), .X(n51699) );
  inv_x2_sg U57479 ( .A(n51700), .X(n51701) );
  inv_x2_sg U57480 ( .A(n51702), .X(n51703) );
  inv_x2_sg U57481 ( .A(n51704), .X(n51705) );
  inv_x2_sg U57482 ( .A(n51706), .X(n51707) );
  inv_x2_sg U57483 ( .A(n51708), .X(n51709) );
  inv_x2_sg U57484 ( .A(n51710), .X(n51711) );
  inv_x2_sg U57485 ( .A(n51712), .X(n51713) );
  inv_x2_sg U57486 ( .A(n51714), .X(n51715) );
  inv_x2_sg U57487 ( .A(n51716), .X(n51717) );
  inv_x2_sg U57488 ( .A(n51718), .X(n51719) );
  inv_x2_sg U57489 ( .A(n51720), .X(n51721) );
  inv_x2_sg U57490 ( .A(n51722), .X(n51723) );
  inv_x2_sg U57491 ( .A(n51724), .X(n51725) );
  inv_x2_sg U57492 ( .A(n51726), .X(n51727) );
  inv_x2_sg U57493 ( .A(n51728), .X(n51729) );
  inv_x2_sg U57494 ( .A(n51730), .X(n51731) );
  inv_x2_sg U57495 ( .A(n51732), .X(n51733) );
  inv_x2_sg U57496 ( .A(n51734), .X(n51735) );
  inv_x2_sg U57497 ( .A(n51736), .X(n51737) );
  inv_x2_sg U57498 ( .A(n51738), .X(n51739) );
  inv_x2_sg U57499 ( .A(n51740), .X(n51741) );
  inv_x2_sg U57500 ( .A(n51742), .X(n51743) );
  inv_x2_sg U57501 ( .A(n51744), .X(n51745) );
  inv_x2_sg U57502 ( .A(n51746), .X(n51747) );
  inv_x2_sg U57503 ( .A(n51748), .X(n51749) );
  inv_x2_sg U57504 ( .A(n51750), .X(n51751) );
  inv_x2_sg U57505 ( .A(n51752), .X(n51753) );
  inv_x2_sg U57506 ( .A(n51754), .X(n51755) );
  inv_x2_sg U57507 ( .A(n51756), .X(n51757) );
  inv_x2_sg U57508 ( .A(n51758), .X(n51759) );
  inv_x2_sg U57509 ( .A(n51760), .X(n51761) );
  inv_x2_sg U57510 ( .A(n51762), .X(n51763) );
  inv_x2_sg U57511 ( .A(n51764), .X(n51765) );
  inv_x2_sg U57512 ( .A(n51766), .X(n51767) );
  inv_x2_sg U57513 ( .A(n51768), .X(n51769) );
  inv_x2_sg U57514 ( .A(n51770), .X(n51771) );
  inv_x2_sg U57515 ( .A(n51772), .X(n51773) );
  inv_x2_sg U57516 ( .A(n51774), .X(n51775) );
  inv_x2_sg U57517 ( .A(n51776), .X(n51777) );
  inv_x2_sg U57518 ( .A(n51778), .X(n51779) );
  inv_x2_sg U57519 ( .A(n51780), .X(n51781) );
  inv_x2_sg U57520 ( .A(n51782), .X(n51783) );
  inv_x2_sg U57521 ( .A(n51784), .X(n51785) );
  inv_x2_sg U57522 ( .A(n51786), .X(n51787) );
  inv_x2_sg U57523 ( .A(n51788), .X(n51789) );
  inv_x2_sg U57524 ( .A(n51790), .X(n51791) );
  inv_x2_sg U57525 ( .A(n51792), .X(n51793) );
  inv_x2_sg U57526 ( .A(n51794), .X(n51795) );
  inv_x2_sg U57527 ( .A(n51796), .X(n51797) );
  inv_x2_sg U57528 ( .A(n51798), .X(n51799) );
  inv_x2_sg U57529 ( .A(n51800), .X(n51801) );
  inv_x2_sg U57530 ( .A(n51802), .X(n51803) );
  inv_x2_sg U57531 ( .A(n51804), .X(n51805) );
  inv_x2_sg U57532 ( .A(n51806), .X(n51807) );
  inv_x2_sg U57533 ( .A(n51808), .X(n51809) );
  inv_x2_sg U57534 ( .A(n51810), .X(n51811) );
  inv_x2_sg U57535 ( .A(n51812), .X(n51813) );
  inv_x2_sg U57536 ( .A(n51814), .X(n51815) );
  inv_x2_sg U57537 ( .A(n51816), .X(n51817) );
  inv_x2_sg U57538 ( .A(n51818), .X(n51819) );
  inv_x2_sg U57539 ( .A(n51820), .X(n51821) );
  inv_x2_sg U57540 ( .A(n51822), .X(n51823) );
  inv_x2_sg U57541 ( .A(n51824), .X(n51825) );
  inv_x2_sg U57542 ( .A(n51826), .X(n51827) );
  inv_x2_sg U57543 ( .A(n51828), .X(n51829) );
  inv_x2_sg U57544 ( .A(n51830), .X(n51831) );
  inv_x2_sg U57545 ( .A(n51832), .X(n51833) );
  inv_x2_sg U57546 ( .A(n51834), .X(n51835) );
  inv_x2_sg U57547 ( .A(n51836), .X(n51837) );
  inv_x2_sg U57548 ( .A(n51838), .X(n51839) );
  inv_x2_sg U57549 ( .A(n51840), .X(n51841) );
  inv_x2_sg U57550 ( .A(n51842), .X(n51843) );
  inv_x2_sg U57551 ( .A(n51844), .X(n51845) );
  inv_x2_sg U57552 ( .A(n51846), .X(n51847) );
  inv_x2_sg U57553 ( .A(n51848), .X(n51849) );
  inv_x2_sg U57554 ( .A(n51850), .X(n51851) );
  inv_x2_sg U57555 ( .A(n51852), .X(n51853) );
  inv_x2_sg U57556 ( .A(n51854), .X(n51855) );
  inv_x2_sg U57557 ( .A(n51856), .X(n51857) );
  inv_x2_sg U57558 ( .A(n51858), .X(n51859) );
  inv_x2_sg U57559 ( .A(n51860), .X(n51861) );
  inv_x2_sg U57560 ( .A(n51862), .X(n51863) );
  inv_x2_sg U57561 ( .A(n51864), .X(n51865) );
  inv_x2_sg U57562 ( .A(n51866), .X(n51867) );
  inv_x2_sg U57563 ( .A(n51868), .X(n51869) );
  inv_x2_sg U57564 ( .A(n51870), .X(n51871) );
  inv_x2_sg U57565 ( .A(n51872), .X(n51873) );
  inv_x2_sg U57566 ( .A(n51874), .X(n51875) );
  inv_x2_sg U57567 ( .A(n51876), .X(n51877) );
  inv_x2_sg U57568 ( .A(n51878), .X(n51879) );
  inv_x2_sg U57569 ( .A(n51880), .X(n51881) );
  inv_x2_sg U57570 ( .A(n51882), .X(n51883) );
  inv_x2_sg U57571 ( .A(n51884), .X(n51885) );
  inv_x2_sg U57572 ( .A(n51886), .X(n51887) );
  inv_x2_sg U57573 ( .A(n51888), .X(n51889) );
  inv_x2_sg U57574 ( .A(n51890), .X(n51891) );
  inv_x2_sg U57575 ( .A(n51892), .X(n51893) );
  inv_x2_sg U57576 ( .A(n51894), .X(n51895) );
  inv_x2_sg U57577 ( .A(n51896), .X(n51897) );
  inv_x2_sg U57578 ( .A(n51898), .X(n51899) );
  inv_x2_sg U57579 ( .A(n51900), .X(n51901) );
  inv_x2_sg U57580 ( .A(n51902), .X(n51903) );
  inv_x2_sg U57581 ( .A(n51904), .X(n51905) );
  inv_x2_sg U57582 ( .A(n51906), .X(n51907) );
  inv_x2_sg U57583 ( .A(n51908), .X(n51909) );
  inv_x2_sg U57584 ( .A(n51910), .X(n51911) );
  inv_x2_sg U57585 ( .A(n51912), .X(n51913) );
  inv_x2_sg U57586 ( .A(n51914), .X(n51915) );
  inv_x2_sg U57587 ( .A(n51916), .X(n51917) );
  inv_x2_sg U57588 ( .A(n51918), .X(n51919) );
  inv_x2_sg U57589 ( .A(n51920), .X(n51921) );
  inv_x2_sg U57590 ( .A(n51922), .X(n51923) );
  inv_x2_sg U57591 ( .A(n51924), .X(n51925) );
  inv_x2_sg U57592 ( .A(n51926), .X(n51927) );
  inv_x2_sg U57593 ( .A(n51928), .X(n51929) );
  inv_x2_sg U57594 ( .A(n51930), .X(n51931) );
  inv_x2_sg U57595 ( .A(n51932), .X(n51933) );
  inv_x2_sg U57596 ( .A(n51934), .X(n51935) );
  inv_x2_sg U57597 ( .A(n51936), .X(n51937) );
  inv_x2_sg U57598 ( .A(n51938), .X(n51939) );
  inv_x2_sg U57599 ( .A(n51940), .X(n51941) );
  inv_x2_sg U57600 ( .A(n51942), .X(n51943) );
  inv_x2_sg U57601 ( .A(n51944), .X(n51945) );
  inv_x2_sg U57602 ( .A(n51946), .X(n51947) );
  inv_x2_sg U57603 ( .A(n51948), .X(n51949) );
  inv_x2_sg U57604 ( .A(n51950), .X(n51951) );
  inv_x2_sg U57605 ( .A(n51952), .X(n51953) );
  inv_x2_sg U57606 ( .A(n51954), .X(n51955) );
  inv_x2_sg U57607 ( .A(n51956), .X(n51957) );
  inv_x2_sg U57608 ( .A(n51958), .X(n51959) );
  inv_x2_sg U57609 ( .A(n51960), .X(n51961) );
  inv_x2_sg U57610 ( .A(n51962), .X(n51963) );
  inv_x2_sg U57611 ( .A(n51964), .X(n51965) );
  inv_x2_sg U57612 ( .A(n51966), .X(n51967) );
  inv_x2_sg U57613 ( .A(n51968), .X(n51969) );
  inv_x2_sg U57614 ( .A(n51970), .X(n51971) );
  inv_x2_sg U57615 ( .A(n51972), .X(n51973) );
  inv_x2_sg U57616 ( .A(n51974), .X(n51975) );
  inv_x2_sg U57617 ( .A(n51976), .X(n51977) );
  inv_x2_sg U57618 ( .A(n51978), .X(n51979) );
  inv_x2_sg U57619 ( .A(n51980), .X(n51981) );
  inv_x2_sg U57620 ( .A(n51982), .X(n51983) );
  inv_x2_sg U57621 ( .A(n51984), .X(n51985) );
  inv_x2_sg U57622 ( .A(n51986), .X(n51987) );
  inv_x2_sg U57623 ( .A(n51988), .X(n51989) );
  inv_x2_sg U57624 ( .A(n51990), .X(n51991) );
  inv_x2_sg U57625 ( .A(n51992), .X(n51993) );
  inv_x2_sg U57626 ( .A(n51994), .X(n51995) );
  inv_x2_sg U57627 ( .A(n51996), .X(n51997) );
  inv_x2_sg U57628 ( .A(n51998), .X(n51999) );
  inv_x2_sg U57629 ( .A(n52000), .X(n52001) );
  inv_x2_sg U57630 ( .A(n52002), .X(n52003) );
  inv_x2_sg U57631 ( .A(n52004), .X(n52005) );
  inv_x2_sg U57632 ( .A(n52006), .X(n52007) );
  inv_x2_sg U57633 ( .A(n52008), .X(n52009) );
  inv_x2_sg U57634 ( .A(n52010), .X(n52011) );
  inv_x2_sg U57635 ( .A(n52012), .X(n52013) );
  inv_x2_sg U57636 ( .A(n52014), .X(n52015) );
  inv_x2_sg U57637 ( .A(n52016), .X(n52017) );
  inv_x2_sg U57638 ( .A(n52018), .X(n52019) );
  inv_x2_sg U57639 ( .A(n52020), .X(n52021) );
  inv_x2_sg U57640 ( .A(n52022), .X(n52023) );
  inv_x2_sg U57641 ( .A(n52024), .X(n52025) );
  inv_x2_sg U57642 ( .A(n52026), .X(n52027) );
  inv_x2_sg U57643 ( .A(n52028), .X(n52029) );
  inv_x2_sg U57644 ( .A(n52030), .X(n52031) );
  inv_x2_sg U57645 ( .A(n52032), .X(n52033) );
  inv_x2_sg U57646 ( .A(n52034), .X(n52035) );
  inv_x2_sg U57647 ( .A(n52036), .X(n52037) );
  inv_x2_sg U57648 ( .A(n52038), .X(n52039) );
  inv_x2_sg U57649 ( .A(n52040), .X(n52041) );
  inv_x2_sg U57650 ( .A(n52042), .X(n52043) );
  inv_x2_sg U57651 ( .A(n52044), .X(n52045) );
  inv_x2_sg U57652 ( .A(n52046), .X(n52047) );
  inv_x2_sg U57653 ( .A(n52048), .X(n52049) );
  inv_x2_sg U57654 ( .A(n52050), .X(n52051) );
  inv_x2_sg U57655 ( .A(n52052), .X(n52053) );
  inv_x2_sg U57656 ( .A(n52054), .X(n52055) );
  inv_x2_sg U57657 ( .A(n52056), .X(n52057) );
  inv_x2_sg U57658 ( .A(n52058), .X(n52059) );
  inv_x2_sg U57659 ( .A(n52060), .X(n52061) );
  inv_x2_sg U57660 ( .A(n52062), .X(n52063) );
  inv_x2_sg U57661 ( .A(n52064), .X(n52065) );
  inv_x2_sg U57662 ( .A(n52066), .X(n52067) );
  inv_x2_sg U57663 ( .A(n52068), .X(n52069) );
  inv_x2_sg U57664 ( .A(n52070), .X(n52071) );
  inv_x2_sg U57665 ( .A(n52072), .X(n52073) );
  inv_x2_sg U57666 ( .A(n52074), .X(n52075) );
  inv_x2_sg U57667 ( .A(n52076), .X(n52077) );
  inv_x2_sg U57668 ( .A(n52078), .X(n52079) );
  inv_x2_sg U57669 ( .A(n52080), .X(n52081) );
  inv_x2_sg U57670 ( .A(n52082), .X(n52083) );
  inv_x2_sg U57671 ( .A(n52084), .X(n52085) );
  inv_x2_sg U57672 ( .A(n52086), .X(n52087) );
  inv_x2_sg U57673 ( .A(n52088), .X(n52089) );
  inv_x2_sg U57674 ( .A(n52090), .X(n52091) );
  inv_x2_sg U57675 ( .A(n52092), .X(n52093) );
  inv_x2_sg U57676 ( .A(n52094), .X(n52095) );
  inv_x2_sg U57677 ( .A(n52096), .X(n52097) );
  inv_x2_sg U57678 ( .A(n52098), .X(n52099) );
  inv_x2_sg U57679 ( .A(n52100), .X(n52101) );
  inv_x2_sg U57680 ( .A(n52102), .X(n52103) );
  inv_x2_sg U57681 ( .A(n52104), .X(n52105) );
  inv_x2_sg U57682 ( .A(n52106), .X(n52107) );
  inv_x2_sg U57683 ( .A(n52108), .X(n52109) );
  inv_x2_sg U57684 ( .A(n52110), .X(n52111) );
  inv_x2_sg U57685 ( .A(n52112), .X(n52113) );
  inv_x2_sg U57686 ( .A(n52114), .X(n52115) );
  inv_x2_sg U57687 ( .A(n52116), .X(n52117) );
  inv_x2_sg U57688 ( .A(n52118), .X(n52119) );
  inv_x2_sg U57689 ( .A(n52120), .X(n52121) );
  inv_x2_sg U57690 ( .A(n52122), .X(n52123) );
  inv_x2_sg U57691 ( .A(n52124), .X(n52125) );
  inv_x2_sg U57692 ( .A(n52126), .X(n52127) );
  inv_x2_sg U57693 ( .A(n52128), .X(n52129) );
  inv_x2_sg U57694 ( .A(n52130), .X(n52131) );
  inv_x2_sg U57695 ( .A(n52132), .X(n52133) );
  inv_x2_sg U57696 ( .A(n52134), .X(n52135) );
  inv_x2_sg U57697 ( .A(n52136), .X(n52137) );
  inv_x2_sg U57698 ( .A(n52138), .X(n52139) );
  inv_x2_sg U57699 ( .A(n52140), .X(n52141) );
  inv_x2_sg U57700 ( .A(n52142), .X(n52143) );
  inv_x2_sg U57701 ( .A(n52144), .X(n52145) );
  inv_x2_sg U57702 ( .A(n52146), .X(n52147) );
  inv_x2_sg U57703 ( .A(n52148), .X(n52149) );
  inv_x2_sg U57704 ( .A(n52150), .X(n52151) );
  inv_x2_sg U57705 ( .A(n52152), .X(n52153) );
  inv_x2_sg U57706 ( .A(n52154), .X(n52155) );
  inv_x2_sg U57707 ( .A(n52156), .X(n52157) );
  inv_x2_sg U57708 ( .A(n52158), .X(n52159) );
  inv_x2_sg U57709 ( .A(n52160), .X(n52161) );
  inv_x2_sg U57710 ( .A(n52162), .X(n52163) );
  inv_x2_sg U57711 ( .A(n52164), .X(n52165) );
  inv_x2_sg U57712 ( .A(n52166), .X(n52167) );
  inv_x2_sg U57713 ( .A(n52168), .X(n52169) );
  inv_x2_sg U57714 ( .A(n52170), .X(n52171) );
  inv_x2_sg U57715 ( .A(n52172), .X(n52173) );
  inv_x2_sg U57716 ( .A(n52174), .X(n52175) );
  inv_x2_sg U57717 ( .A(n52176), .X(n52177) );
  inv_x2_sg U57718 ( .A(n52178), .X(n52179) );
  inv_x2_sg U57719 ( .A(n52180), .X(n52181) );
  inv_x2_sg U57720 ( .A(n52182), .X(n52183) );
  inv_x2_sg U57721 ( .A(n52184), .X(n52185) );
  inv_x2_sg U57722 ( .A(n52186), .X(n52187) );
  inv_x2_sg U57723 ( .A(n52188), .X(n52189) );
  inv_x2_sg U57724 ( .A(n52190), .X(n52191) );
  inv_x2_sg U57725 ( .A(n52192), .X(n52193) );
  inv_x2_sg U57726 ( .A(n52194), .X(n52195) );
  inv_x2_sg U57727 ( .A(n52196), .X(n52197) );
  inv_x2_sg U57728 ( .A(n52198), .X(n52199) );
  inv_x2_sg U57729 ( .A(n52200), .X(n52201) );
  inv_x2_sg U57730 ( .A(n52202), .X(n52203) );
  inv_x2_sg U57731 ( .A(n52204), .X(n52205) );
  inv_x2_sg U57732 ( .A(n52206), .X(n52207) );
  inv_x2_sg U57733 ( .A(n52208), .X(n52209) );
  inv_x2_sg U57734 ( .A(n52210), .X(n52211) );
  inv_x2_sg U57735 ( .A(n52212), .X(n52213) );
  inv_x2_sg U57736 ( .A(n52214), .X(n52215) );
  inv_x2_sg U57737 ( .A(n52216), .X(n52217) );
  inv_x2_sg U57738 ( .A(n52218), .X(n52219) );
  inv_x2_sg U57739 ( .A(n52220), .X(n52221) );
  inv_x2_sg U57740 ( .A(n52222), .X(n52223) );
  inv_x2_sg U57741 ( .A(n52224), .X(n52225) );
  inv_x2_sg U57742 ( .A(n52226), .X(n52227) );
  inv_x2_sg U57743 ( .A(n52228), .X(n52229) );
  inv_x2_sg U57744 ( .A(n52230), .X(n52231) );
  inv_x2_sg U57745 ( .A(n52232), .X(n52233) );
  inv_x2_sg U57746 ( .A(n52234), .X(n52235) );
  inv_x2_sg U57747 ( .A(n52236), .X(n52237) );
  inv_x2_sg U57748 ( .A(n52238), .X(n52239) );
  inv_x2_sg U57749 ( .A(n52240), .X(n52241) );
  inv_x2_sg U57750 ( .A(n52242), .X(n52243) );
  inv_x2_sg U57751 ( .A(n52244), .X(n52245) );
  inv_x2_sg U57752 ( .A(n52246), .X(n52247) );
  inv_x2_sg U57753 ( .A(n52248), .X(n52249) );
  inv_x2_sg U57754 ( .A(n52250), .X(n52251) );
  inv_x2_sg U57755 ( .A(n52252), .X(n52253) );
  inv_x2_sg U57756 ( .A(n52254), .X(n52255) );
  inv_x2_sg U57757 ( .A(n52256), .X(n52257) );
  inv_x2_sg U57758 ( .A(n52258), .X(n52259) );
  inv_x2_sg U57759 ( .A(n52260), .X(n52261) );
  inv_x2_sg U57760 ( .A(n52262), .X(n52263) );
  inv_x2_sg U57761 ( .A(n52264), .X(n52265) );
  inv_x2_sg U57762 ( .A(n52266), .X(n52267) );
  inv_x2_sg U57763 ( .A(n52268), .X(n52269) );
  inv_x2_sg U57764 ( .A(n52270), .X(n52271) );
  inv_x2_sg U57765 ( .A(n52272), .X(n52273) );
  inv_x2_sg U57766 ( .A(n52274), .X(n52275) );
  inv_x2_sg U57767 ( .A(n52276), .X(n52277) );
  inv_x2_sg U57768 ( .A(n52278), .X(n52279) );
  inv_x2_sg U57769 ( .A(n52280), .X(n52281) );
  inv_x2_sg U57770 ( .A(n52282), .X(n52283) );
  inv_x2_sg U57771 ( .A(n52284), .X(n52285) );
  inv_x2_sg U57772 ( .A(n52286), .X(n52287) );
  inv_x2_sg U57773 ( .A(n52288), .X(n52289) );
  inv_x2_sg U57774 ( .A(n52290), .X(n52291) );
  inv_x2_sg U57775 ( .A(n52292), .X(n52293) );
  inv_x2_sg U57776 ( .A(n52294), .X(n52295) );
  inv_x2_sg U57777 ( .A(n52296), .X(n52297) );
  inv_x2_sg U57778 ( .A(n52298), .X(n52299) );
  inv_x2_sg U57779 ( .A(n52300), .X(n52301) );
  inv_x2_sg U57780 ( .A(n52302), .X(n52303) );
  inv_x2_sg U57781 ( .A(n52304), .X(n52305) );
  inv_x2_sg U57782 ( .A(n52306), .X(n52307) );
  inv_x2_sg U57783 ( .A(n52308), .X(n52309) );
  inv_x2_sg U57784 ( .A(n52310), .X(n52311) );
  inv_x2_sg U57785 ( .A(n52312), .X(n52313) );
  inv_x2_sg U57786 ( .A(n52314), .X(n52315) );
  inv_x2_sg U57787 ( .A(n52316), .X(n52317) );
  inv_x2_sg U57788 ( .A(n52318), .X(n52319) );
  inv_x2_sg U57789 ( .A(n52320), .X(n52321) );
  inv_x2_sg U57790 ( .A(n52322), .X(n52323) );
  inv_x2_sg U57791 ( .A(n52324), .X(n52325) );
  inv_x2_sg U57792 ( .A(n52326), .X(n52327) );
  inv_x2_sg U57793 ( .A(n52328), .X(n52329) );
  inv_x2_sg U57794 ( .A(n52330), .X(n52331) );
  inv_x2_sg U57795 ( .A(n52332), .X(n52333) );
  inv_x2_sg U57796 ( .A(n52334), .X(n52335) );
  inv_x2_sg U57797 ( .A(n52336), .X(n52337) );
  inv_x2_sg U57798 ( .A(n52338), .X(n52339) );
  inv_x2_sg U57799 ( .A(n52340), .X(n52341) );
  inv_x2_sg U57800 ( .A(n52342), .X(n52343) );
  inv_x2_sg U57801 ( .A(n52344), .X(n52345) );
  inv_x2_sg U57802 ( .A(n52346), .X(n52347) );
  inv_x2_sg U57803 ( .A(n52348), .X(n52349) );
  inv_x2_sg U57804 ( .A(n52350), .X(n52351) );
  inv_x2_sg U57805 ( .A(n52352), .X(n52353) );
  inv_x2_sg U57806 ( .A(n52354), .X(n52355) );
  inv_x2_sg U57807 ( .A(n52356), .X(n52357) );
  inv_x2_sg U57808 ( .A(n52358), .X(n52359) );
  inv_x2_sg U57809 ( .A(n52360), .X(n52361) );
  inv_x2_sg U57810 ( .A(n52362), .X(n52363) );
  inv_x2_sg U57811 ( .A(n52364), .X(n52365) );
  inv_x2_sg U57812 ( .A(n52366), .X(n52367) );
  inv_x2_sg U57813 ( .A(n52368), .X(n52369) );
  inv_x2_sg U57814 ( .A(n52370), .X(n52371) );
  inv_x2_sg U57815 ( .A(n52372), .X(n52373) );
  inv_x2_sg U57816 ( .A(n52374), .X(n52375) );
  inv_x2_sg U57817 ( .A(n52376), .X(n52377) );
  inv_x2_sg U57818 ( .A(n52378), .X(n52379) );
  inv_x2_sg U57819 ( .A(n52380), .X(n52381) );
  inv_x2_sg U57820 ( .A(n52382), .X(n52383) );
  inv_x2_sg U57821 ( .A(n52384), .X(n52385) );
  inv_x2_sg U57822 ( .A(n52386), .X(n52387) );
  inv_x2_sg U57823 ( .A(n52388), .X(n52389) );
  inv_x2_sg U57824 ( .A(n52390), .X(n52391) );
  inv_x2_sg U57825 ( .A(n52392), .X(n52393) );
  inv_x2_sg U57826 ( .A(n52394), .X(n52395) );
  inv_x2_sg U57827 ( .A(n52396), .X(n52397) );
  inv_x2_sg U57828 ( .A(n52398), .X(n52399) );
  inv_x2_sg U57829 ( .A(n52400), .X(n52401) );
  inv_x2_sg U57830 ( .A(n52402), .X(n52403) );
  inv_x2_sg U57831 ( .A(n52404), .X(n52405) );
  inv_x2_sg U57832 ( .A(n52406), .X(n52407) );
  inv_x2_sg U57833 ( .A(n52408), .X(n52409) );
  inv_x2_sg U57834 ( .A(n52410), .X(n52411) );
  inv_x2_sg U57835 ( .A(n52412), .X(n52413) );
  inv_x2_sg U57836 ( .A(n52414), .X(n52415) );
  inv_x2_sg U57837 ( .A(n52416), .X(n52417) );
  inv_x2_sg U57838 ( .A(n52418), .X(n52419) );
  inv_x2_sg U57839 ( .A(n52420), .X(n52421) );
  inv_x2_sg U57840 ( .A(n52422), .X(n52423) );
  inv_x2_sg U57841 ( .A(n52424), .X(n52425) );
  inv_x2_sg U57842 ( .A(n52426), .X(n52427) );
  inv_x2_sg U57843 ( .A(n52428), .X(n52429) );
  inv_x2_sg U57844 ( .A(n52430), .X(n52431) );
  inv_x2_sg U57845 ( .A(n52432), .X(n52433) );
  inv_x2_sg U57846 ( .A(n52434), .X(n52435) );
  inv_x2_sg U57847 ( .A(n52436), .X(n52437) );
  inv_x2_sg U57848 ( .A(n52438), .X(n52439) );
  inv_x2_sg U57849 ( .A(n52440), .X(n52441) );
  inv_x2_sg U57850 ( .A(n52442), .X(n52443) );
  inv_x2_sg U57851 ( .A(n52444), .X(n52445) );
  inv_x2_sg U57852 ( .A(n52446), .X(n52447) );
  inv_x2_sg U57853 ( .A(n52448), .X(n52449) );
  inv_x2_sg U57854 ( .A(n52450), .X(n52451) );
  inv_x2_sg U57855 ( .A(n52452), .X(n52453) );
  inv_x2_sg U57856 ( .A(n52454), .X(n52455) );
  inv_x2_sg U57857 ( .A(n52456), .X(n52457) );
  inv_x2_sg U57858 ( .A(n52458), .X(n52459) );
  inv_x2_sg U57859 ( .A(n52460), .X(n52461) );
  inv_x2_sg U57860 ( .A(n52462), .X(n52463) );
  inv_x2_sg U57861 ( .A(n52464), .X(n52465) );
  inv_x2_sg U57862 ( .A(n52466), .X(n52467) );
  inv_x2_sg U57863 ( .A(n52468), .X(n52469) );
  inv_x2_sg U57864 ( .A(n52470), .X(n52471) );
  inv_x2_sg U57865 ( .A(n52472), .X(n52473) );
  inv_x2_sg U57866 ( .A(n52474), .X(n52475) );
  inv_x2_sg U57867 ( .A(n52476), .X(n52477) );
  inv_x2_sg U57868 ( .A(n52478), .X(n52479) );
  inv_x2_sg U57869 ( .A(n52480), .X(n52481) );
  inv_x2_sg U57870 ( .A(n52482), .X(n52483) );
  inv_x2_sg U57871 ( .A(n52484), .X(n52485) );
  inv_x2_sg U57872 ( .A(n52486), .X(n52487) );
  inv_x2_sg U57873 ( .A(n52488), .X(n52489) );
  inv_x2_sg U57874 ( .A(n52490), .X(n52491) );
  inv_x2_sg U57875 ( .A(n52492), .X(n52493) );
  inv_x2_sg U57876 ( .A(n52494), .X(n52495) );
  inv_x2_sg U57877 ( .A(n52496), .X(n52497) );
  inv_x2_sg U57878 ( .A(n52498), .X(n52499) );
  inv_x2_sg U57879 ( .A(n52500), .X(n52501) );
  inv_x2_sg U57880 ( .A(n52502), .X(n52503) );
  inv_x2_sg U57881 ( .A(n52504), .X(n52505) );
  inv_x2_sg U57882 ( .A(n52506), .X(n52507) );
  inv_x2_sg U57883 ( .A(n52508), .X(n52509) );
  inv_x2_sg U57884 ( .A(n52510), .X(n52511) );
  inv_x2_sg U57885 ( .A(n52512), .X(n52513) );
  inv_x2_sg U57886 ( .A(n52514), .X(n52515) );
  inv_x2_sg U57887 ( .A(n52516), .X(n52517) );
  inv_x2_sg U57888 ( .A(n52518), .X(n52519) );
  inv_x2_sg U57889 ( .A(n52520), .X(n52521) );
  inv_x2_sg U57890 ( .A(n52522), .X(n52523) );
  inv_x2_sg U57891 ( .A(n52524), .X(n52525) );
  inv_x2_sg U57892 ( .A(n52526), .X(n52527) );
  inv_x2_sg U57893 ( .A(n52528), .X(n52529) );
  inv_x2_sg U57894 ( .A(n52530), .X(n52531) );
  inv_x2_sg U57895 ( .A(n52532), .X(n52533) );
  inv_x2_sg U57896 ( .A(n52534), .X(n52535) );
  inv_x2_sg U57897 ( .A(n52536), .X(n52537) );
  inv_x2_sg U57898 ( .A(n52538), .X(n52539) );
  inv_x2_sg U57899 ( .A(n52540), .X(n52541) );
  inv_x2_sg U57900 ( .A(n52542), .X(n52543) );
  inv_x2_sg U57901 ( .A(n52544), .X(n52545) );
  inv_x2_sg U57902 ( .A(n52546), .X(n52547) );
  inv_x2_sg U57903 ( .A(n52548), .X(n52549) );
  inv_x2_sg U57904 ( .A(n52550), .X(n52551) );
  inv_x2_sg U57905 ( .A(n52552), .X(n52553) );
  inv_x2_sg U57906 ( .A(n52554), .X(n52555) );
  inv_x2_sg U57907 ( .A(n52556), .X(n52557) );
  inv_x2_sg U57908 ( .A(n52558), .X(n52559) );
  inv_x2_sg U57909 ( .A(n52560), .X(n52561) );
  inv_x2_sg U57910 ( .A(n52562), .X(n52563) );
  inv_x2_sg U57911 ( .A(n52564), .X(n52565) );
  inv_x2_sg U57912 ( .A(n52566), .X(n52567) );
  inv_x2_sg U57913 ( .A(n52568), .X(n52569) );
  inv_x2_sg U57914 ( .A(n52570), .X(n52571) );
  inv_x2_sg U57915 ( .A(n52572), .X(n52573) );
  inv_x2_sg U57916 ( .A(n52574), .X(n52575) );
  inv_x2_sg U57917 ( .A(n52576), .X(n52577) );
  inv_x2_sg U57918 ( .A(n52578), .X(n52579) );
  inv_x2_sg U57919 ( .A(n52580), .X(n52581) );
  inv_x2_sg U57920 ( .A(n52582), .X(n52583) );
  inv_x2_sg U57921 ( .A(n52584), .X(n52585) );
  inv_x2_sg U57922 ( .A(n52586), .X(n52587) );
  inv_x2_sg U57923 ( .A(n52588), .X(n52589) );
  inv_x2_sg U57924 ( .A(n52590), .X(n52591) );
  inv_x2_sg U57925 ( .A(n52592), .X(n52593) );
  inv_x2_sg U57926 ( .A(n52594), .X(n52595) );
  inv_x2_sg U57927 ( .A(n52596), .X(n52597) );
  inv_x2_sg U57928 ( .A(n52598), .X(n52599) );
  inv_x2_sg U57929 ( .A(n52600), .X(n52601) );
  inv_x2_sg U57930 ( .A(n52602), .X(n52603) );
  inv_x2_sg U57931 ( .A(n52604), .X(n52605) );
  inv_x2_sg U57932 ( .A(n52606), .X(n52607) );
  inv_x2_sg U57933 ( .A(n52608), .X(n52609) );
  inv_x2_sg U57934 ( .A(n52610), .X(n52611) );
  inv_x2_sg U57935 ( .A(n52612), .X(n52613) );
  inv_x2_sg U57936 ( .A(n52614), .X(n52615) );
  inv_x2_sg U57937 ( .A(n52616), .X(n52617) );
  inv_x2_sg U57938 ( .A(n52618), .X(n52619) );
  inv_x2_sg U57939 ( .A(n52620), .X(n52621) );
  inv_x2_sg U57940 ( .A(n52622), .X(n52623) );
  inv_x2_sg U57941 ( .A(n52624), .X(n52625) );
  inv_x2_sg U57942 ( .A(n52626), .X(n52627) );
  inv_x2_sg U57943 ( .A(n52628), .X(n52629) );
  inv_x2_sg U57944 ( .A(n52630), .X(n52631) );
  inv_x2_sg U57945 ( .A(n52632), .X(n52633) );
  inv_x2_sg U57946 ( .A(n52634), .X(n52635) );
  inv_x2_sg U57947 ( .A(n52636), .X(n52637) );
  inv_x2_sg U57948 ( .A(n52638), .X(n52639) );
  inv_x2_sg U57949 ( .A(n52640), .X(n52641) );
  inv_x2_sg U57950 ( .A(n52642), .X(n52643) );
  inv_x2_sg U57951 ( .A(n52644), .X(n52645) );
  inv_x2_sg U57952 ( .A(n52646), .X(n52647) );
  inv_x2_sg U57953 ( .A(n52648), .X(n52649) );
  inv_x2_sg U57954 ( .A(n52650), .X(n52651) );
  inv_x2_sg U57955 ( .A(n52652), .X(n52653) );
  inv_x2_sg U57956 ( .A(n52654), .X(n52655) );
  inv_x2_sg U57957 ( .A(n52656), .X(n52657) );
  inv_x2_sg U57958 ( .A(n52658), .X(n52659) );
  inv_x2_sg U57959 ( .A(n52660), .X(n52661) );
  inv_x2_sg U57960 ( .A(n52662), .X(n52663) );
  inv_x2_sg U57961 ( .A(n52664), .X(n52665) );
  inv_x2_sg U57962 ( .A(n52666), .X(n52667) );
  inv_x2_sg U57963 ( .A(n52668), .X(n52669) );
  inv_x2_sg U57964 ( .A(n52670), .X(n52671) );
  inv_x2_sg U57965 ( .A(n52672), .X(n52673) );
  inv_x2_sg U57966 ( .A(n52674), .X(n52675) );
  inv_x2_sg U57967 ( .A(n52676), .X(n52677) );
  inv_x2_sg U57968 ( .A(n52678), .X(n52679) );
  inv_x2_sg U57969 ( .A(n52680), .X(n52681) );
  inv_x2_sg U57970 ( .A(n52682), .X(n52683) );
  inv_x2_sg U57971 ( .A(n52684), .X(n52685) );
  inv_x2_sg U57972 ( .A(n52686), .X(n52687) );
  inv_x2_sg U57973 ( .A(n52688), .X(n52689) );
  inv_x2_sg U57974 ( .A(n52690), .X(n52691) );
  inv_x2_sg U57975 ( .A(n52692), .X(n52693) );
  inv_x2_sg U57976 ( .A(n52694), .X(n52695) );
  inv_x2_sg U57977 ( .A(n52696), .X(n52697) );
  inv_x2_sg U57978 ( .A(n52698), .X(n52699) );
  inv_x2_sg U57979 ( .A(n52700), .X(n52701) );
  inv_x2_sg U57980 ( .A(n52702), .X(n52703) );
  inv_x2_sg U57981 ( .A(n52704), .X(n52705) );
  inv_x2_sg U57982 ( .A(n52706), .X(n52707) );
  inv_x2_sg U57983 ( .A(n52708), .X(n52709) );
  inv_x2_sg U57984 ( .A(n52710), .X(n52711) );
  inv_x2_sg U57985 ( .A(n52712), .X(n52713) );
  inv_x2_sg U57986 ( .A(n52714), .X(n52715) );
  inv_x2_sg U57987 ( .A(n52716), .X(n52717) );
  inv_x2_sg U57988 ( .A(n52718), .X(n52719) );
  inv_x2_sg U57989 ( .A(n52720), .X(n52721) );
  inv_x2_sg U57990 ( .A(n52722), .X(n52723) );
  inv_x2_sg U57991 ( .A(n52724), .X(n52725) );
  inv_x2_sg U57992 ( .A(n52726), .X(n52727) );
  inv_x2_sg U57993 ( .A(n52728), .X(n52729) );
  inv_x2_sg U57994 ( .A(n52730), .X(n52731) );
  inv_x2_sg U57995 ( .A(n52732), .X(n52733) );
  inv_x2_sg U57996 ( .A(n52734), .X(n52735) );
  inv_x2_sg U57997 ( .A(n52736), .X(n52737) );
  inv_x2_sg U57998 ( .A(n52738), .X(n52739) );
  inv_x2_sg U57999 ( .A(n52740), .X(n52741) );
  inv_x2_sg U58000 ( .A(n52742), .X(n52743) );
  inv_x2_sg U58001 ( .A(n52744), .X(n52745) );
  inv_x2_sg U58002 ( .A(n52746), .X(n52747) );
  inv_x2_sg U58003 ( .A(n52748), .X(n52749) );
  inv_x2_sg U58004 ( .A(n52750), .X(n52751) );
  inv_x2_sg U58005 ( .A(n52752), .X(n52753) );
  inv_x2_sg U58006 ( .A(n52754), .X(n52755) );
  inv_x2_sg U58007 ( .A(n52756), .X(n52757) );
  inv_x2_sg U58008 ( .A(n52758), .X(n52759) );
  inv_x2_sg U58009 ( .A(n52760), .X(n52761) );
  inv_x2_sg U58010 ( .A(n52762), .X(n52763) );
  inv_x2_sg U58011 ( .A(n52764), .X(n52765) );
  inv_x2_sg U58012 ( .A(n52766), .X(n52767) );
  inv_x2_sg U58013 ( .A(n52768), .X(n52769) );
  inv_x2_sg U58014 ( .A(n52770), .X(n52771) );
  inv_x2_sg U58015 ( .A(n52772), .X(n52773) );
  inv_x2_sg U58016 ( .A(n52774), .X(n52775) );
  inv_x2_sg U58017 ( .A(n52776), .X(n52777) );
  inv_x2_sg U58018 ( .A(n52778), .X(n52779) );
  inv_x2_sg U58019 ( .A(n52780), .X(n52781) );
  inv_x2_sg U58020 ( .A(n52782), .X(n52783) );
  inv_x2_sg U58021 ( .A(n52784), .X(n52785) );
  inv_x2_sg U58022 ( .A(n52786), .X(n52787) );
  inv_x2_sg U58023 ( .A(n52788), .X(n52789) );
  inv_x2_sg U58024 ( .A(n52790), .X(n52791) );
  inv_x2_sg U58025 ( .A(n52792), .X(n52793) );
  inv_x2_sg U58026 ( .A(n52794), .X(n52795) );
  inv_x2_sg U58027 ( .A(n52796), .X(n52797) );
  inv_x2_sg U58028 ( .A(n52798), .X(n52799) );
  inv_x2_sg U58029 ( .A(n52800), .X(n52801) );
  inv_x2_sg U58030 ( .A(n52802), .X(n52803) );
  inv_x2_sg U58031 ( .A(n52804), .X(n52805) );
  inv_x2_sg U58032 ( .A(n52806), .X(n52807) );
  inv_x2_sg U58033 ( .A(n52808), .X(n52809) );
  inv_x2_sg U58034 ( .A(n52810), .X(n52811) );
  inv_x2_sg U58035 ( .A(n52812), .X(n52813) );
  inv_x2_sg U58036 ( .A(n52814), .X(n52815) );
  inv_x2_sg U58037 ( .A(n52816), .X(n52817) );
  inv_x2_sg U58038 ( .A(n52818), .X(n52819) );
  inv_x2_sg U58039 ( .A(n52820), .X(n52821) );
  inv_x2_sg U58040 ( .A(n52822), .X(n52823) );
  inv_x2_sg U58041 ( .A(n52824), .X(n52825) );
  inv_x2_sg U58042 ( .A(n52826), .X(n52827) );
  inv_x2_sg U58043 ( .A(n52828), .X(n52829) );
  inv_x2_sg U58044 ( .A(n52830), .X(n52831) );
  inv_x2_sg U58045 ( .A(n52832), .X(n52833) );
  inv_x2_sg U58046 ( .A(n52834), .X(n52835) );
  inv_x2_sg U58047 ( .A(n52836), .X(n52837) );
  inv_x2_sg U58048 ( .A(n52838), .X(n52839) );
  inv_x2_sg U58049 ( .A(n52840), .X(n52841) );
  inv_x2_sg U58050 ( .A(n52842), .X(n52843) );
  inv_x2_sg U58051 ( .A(n52844), .X(n52845) );
  inv_x2_sg U58052 ( .A(n52846), .X(n52847) );
  inv_x2_sg U58053 ( .A(n52848), .X(n52849) );
  inv_x2_sg U58054 ( .A(n52850), .X(n52851) );
  inv_x2_sg U58055 ( .A(n52852), .X(n52853) );
  inv_x2_sg U58056 ( .A(n52854), .X(n52855) );
  inv_x2_sg U58057 ( .A(n52856), .X(n52857) );
  inv_x2_sg U58058 ( .A(n52858), .X(n52859) );
  inv_x2_sg U58059 ( .A(n52860), .X(n52861) );
  inv_x2_sg U58060 ( .A(n52862), .X(n52863) );
  inv_x2_sg U58061 ( .A(n52864), .X(n52865) );
  inv_x2_sg U58062 ( .A(n52866), .X(n52867) );
  inv_x2_sg U58063 ( .A(n52868), .X(n52869) );
  inv_x2_sg U58064 ( .A(n52870), .X(n52871) );
  inv_x2_sg U58065 ( .A(n52872), .X(n52873) );
  inv_x2_sg U58066 ( .A(n52874), .X(n52875) );
  inv_x2_sg U58067 ( .A(n52876), .X(n52877) );
  inv_x2_sg U58068 ( .A(n52878), .X(n52879) );
  inv_x2_sg U58069 ( .A(n52880), .X(n52881) );
  inv_x2_sg U58070 ( .A(n52882), .X(n52883) );
  inv_x2_sg U58071 ( .A(n52884), .X(n52885) );
  inv_x2_sg U58072 ( .A(n52886), .X(n52887) );
  inv_x2_sg U58073 ( .A(n52888), .X(n52889) );
  inv_x2_sg U58074 ( .A(n52890), .X(n52891) );
  inv_x2_sg U58075 ( .A(n52892), .X(n52893) );
  inv_x2_sg U58076 ( .A(n52894), .X(n52895) );
  inv_x2_sg U58077 ( .A(n52896), .X(n52897) );
  inv_x2_sg U58078 ( .A(n52898), .X(n52899) );
  inv_x2_sg U58079 ( .A(n52900), .X(n52901) );
  inv_x2_sg U58080 ( .A(n52902), .X(n52903) );
  inv_x2_sg U58081 ( .A(n52904), .X(n52905) );
  inv_x2_sg U58082 ( .A(n52906), .X(n52907) );
  inv_x2_sg U58083 ( .A(n52908), .X(n52909) );
  inv_x2_sg U58084 ( .A(n52910), .X(n52911) );
  inv_x2_sg U58085 ( .A(n52912), .X(n52913) );
  inv_x2_sg U58086 ( .A(n52914), .X(n52915) );
  inv_x2_sg U58087 ( .A(n52916), .X(n52917) );
  inv_x2_sg U58088 ( .A(n52918), .X(n52919) );
  inv_x2_sg U58089 ( .A(n52920), .X(n52921) );
  inv_x2_sg U58090 ( .A(n52922), .X(n52923) );
  inv_x2_sg U58091 ( .A(n52924), .X(n52925) );
  inv_x2_sg U58092 ( .A(n52926), .X(n52927) );
  inv_x2_sg U58093 ( .A(n52928), .X(n52929) );
  inv_x2_sg U58094 ( .A(n52930), .X(n52931) );
  inv_x2_sg U58095 ( .A(n52932), .X(n52933) );
  inv_x2_sg U58096 ( .A(n52934), .X(n52935) );
  inv_x2_sg U58097 ( .A(n52936), .X(n52937) );
  inv_x2_sg U58098 ( .A(n52938), .X(n52939) );
  inv_x2_sg U58099 ( .A(n52940), .X(n52941) );
  inv_x2_sg U58100 ( .A(n52942), .X(n52943) );
  inv_x2_sg U58101 ( .A(n52944), .X(n52945) );
  inv_x2_sg U58102 ( .A(n52946), .X(n52947) );
  inv_x2_sg U58103 ( .A(n52948), .X(n52949) );
  inv_x2_sg U58104 ( .A(n52950), .X(n52951) );
  inv_x2_sg U58105 ( .A(n52952), .X(n52953) );
  inv_x2_sg U58106 ( .A(n52954), .X(n52955) );
  inv_x2_sg U58107 ( .A(n52956), .X(n52957) );
  inv_x2_sg U58108 ( .A(n52958), .X(n52959) );
  inv_x2_sg U58109 ( .A(n52960), .X(n52961) );
  inv_x2_sg U58110 ( .A(n52962), .X(n52963) );
  inv_x2_sg U58111 ( .A(n52964), .X(n52965) );
  inv_x2_sg U58112 ( .A(n52966), .X(n52967) );
  inv_x2_sg U58113 ( .A(n52968), .X(n52969) );
  inv_x2_sg U58114 ( .A(n52970), .X(n52971) );
  inv_x2_sg U58115 ( .A(n52972), .X(n52973) );
  inv_x2_sg U58116 ( .A(n52974), .X(n52975) );
  inv_x2_sg U58117 ( .A(n52976), .X(n52977) );
  inv_x2_sg U58118 ( .A(n52978), .X(n52979) );
  inv_x2_sg U58119 ( .A(n52980), .X(n52981) );
  inv_x2_sg U58120 ( .A(n52982), .X(n52983) );
  inv_x2_sg U58121 ( .A(n52984), .X(n52985) );
  inv_x2_sg U58122 ( .A(n52986), .X(n52987) );
  inv_x2_sg U58123 ( .A(n52988), .X(n52989) );
  inv_x2_sg U58124 ( .A(n52990), .X(n52991) );
  inv_x2_sg U58125 ( .A(n52992), .X(n52993) );
  inv_x2_sg U58126 ( .A(n52994), .X(n52995) );
  inv_x2_sg U58127 ( .A(n52996), .X(n52997) );
  inv_x2_sg U58128 ( .A(n52998), .X(n52999) );
  inv_x2_sg U58129 ( .A(n53000), .X(n53001) );
  inv_x2_sg U58130 ( .A(n53002), .X(n53003) );
  inv_x2_sg U58131 ( .A(n53004), .X(n53005) );
  inv_x2_sg U58132 ( .A(n53006), .X(n53007) );
  inv_x2_sg U58133 ( .A(n53008), .X(n53009) );
  inv_x2_sg U58134 ( .A(n53010), .X(n53011) );
  inv_x2_sg U58135 ( .A(n53012), .X(n53013) );
  inv_x2_sg U58136 ( .A(n53014), .X(n53015) );
  inv_x2_sg U58137 ( .A(n53016), .X(n53017) );
  inv_x2_sg U58138 ( .A(n53018), .X(n53019) );
  inv_x2_sg U58139 ( .A(n53020), .X(n53021) );
  inv_x2_sg U58140 ( .A(n53022), .X(n53023) );
  inv_x2_sg U58141 ( .A(n53024), .X(n53025) );
  inv_x2_sg U58142 ( .A(n53026), .X(n53027) );
  inv_x2_sg U58143 ( .A(n53028), .X(n53029) );
  inv_x2_sg U58144 ( .A(n53030), .X(n53031) );
  inv_x2_sg U58145 ( .A(n53032), .X(n53033) );
  inv_x2_sg U58146 ( .A(n53034), .X(n53035) );
  inv_x2_sg U58147 ( .A(n53036), .X(n53037) );
  inv_x2_sg U58148 ( .A(n53038), .X(n53039) );
  inv_x2_sg U58149 ( .A(n53040), .X(n53041) );
  inv_x2_sg U58150 ( .A(n53042), .X(n53043) );
  inv_x2_sg U58151 ( .A(n53044), .X(n53045) );
  inv_x2_sg U58152 ( .A(n53046), .X(n53047) );
  inv_x2_sg U58153 ( .A(n53048), .X(n53049) );
  inv_x2_sg U58154 ( .A(n53050), .X(n53051) );
  inv_x2_sg U58155 ( .A(n53052), .X(n53053) );
  inv_x2_sg U58156 ( .A(n53054), .X(n53055) );
  inv_x2_sg U58157 ( .A(n53056), .X(n53057) );
  inv_x2_sg U58158 ( .A(n53058), .X(n53059) );
  inv_x2_sg U58159 ( .A(n53060), .X(n53061) );
  inv_x2_sg U58160 ( .A(n53062), .X(n53063) );
  inv_x2_sg U58161 ( .A(n53064), .X(n53065) );
  inv_x2_sg U58162 ( .A(n53066), .X(n53067) );
  inv_x2_sg U58163 ( .A(n53068), .X(n53069) );
  inv_x2_sg U58164 ( .A(n53070), .X(n53071) );
  inv_x2_sg U58165 ( .A(n53072), .X(n53073) );
  inv_x2_sg U58166 ( .A(n53074), .X(n53075) );
  inv_x2_sg U58167 ( .A(n53076), .X(n53077) );
  inv_x2_sg U58168 ( .A(n53078), .X(n53079) );
  inv_x2_sg U58169 ( .A(n53080), .X(n53081) );
  inv_x2_sg U58170 ( .A(n53082), .X(n53083) );
  inv_x2_sg U58171 ( .A(n53084), .X(n53085) );
  inv_x2_sg U58172 ( .A(n53086), .X(n53087) );
  inv_x2_sg U58173 ( .A(n53088), .X(n53089) );
  inv_x2_sg U58174 ( .A(n53090), .X(n53091) );
  inv_x2_sg U58175 ( .A(n53092), .X(n53093) );
  inv_x2_sg U58176 ( .A(n53094), .X(n53095) );
  inv_x2_sg U58177 ( .A(n53096), .X(n53097) );
  inv_x2_sg U58178 ( .A(n53098), .X(n53099) );
  inv_x2_sg U58179 ( .A(n53100), .X(n53101) );
  inv_x2_sg U58180 ( .A(n53102), .X(n53103) );
  inv_x2_sg U58181 ( .A(n53104), .X(n53105) );
  inv_x2_sg U58182 ( .A(n53106), .X(n53107) );
  inv_x2_sg U58183 ( .A(n53108), .X(n53109) );
  inv_x2_sg U58184 ( .A(n53110), .X(n53111) );
  inv_x2_sg U58185 ( .A(n53112), .X(n53113) );
  inv_x2_sg U58186 ( .A(n53114), .X(n53115) );
  inv_x2_sg U58187 ( .A(n53116), .X(n53117) );
  inv_x2_sg U58188 ( .A(n53118), .X(n53119) );
  inv_x2_sg U58189 ( .A(n53120), .X(n53121) );
  inv_x2_sg U58190 ( .A(n53122), .X(n53123) );
  inv_x2_sg U58191 ( .A(n53124), .X(n53125) );
  inv_x2_sg U58192 ( .A(n53126), .X(n53127) );
  inv_x2_sg U58193 ( .A(n53128), .X(n53129) );
  inv_x2_sg U58194 ( .A(n53130), .X(n53131) );
  inv_x2_sg U58195 ( .A(n53132), .X(n53133) );
  inv_x2_sg U58196 ( .A(n53134), .X(n53135) );
  inv_x2_sg U58197 ( .A(n53136), .X(n53137) );
  inv_x2_sg U58198 ( .A(n53138), .X(n53139) );
  inv_x2_sg U58199 ( .A(n53140), .X(n53141) );
  inv_x2_sg U58200 ( .A(n53142), .X(n53143) );
  inv_x2_sg U58201 ( .A(n53144), .X(n53145) );
  inv_x2_sg U58202 ( .A(n53146), .X(n53147) );
  inv_x2_sg U58203 ( .A(n53148), .X(n53149) );
  inv_x2_sg U58204 ( .A(n53150), .X(n53151) );
  inv_x2_sg U58205 ( .A(n53152), .X(n53153) );
  inv_x2_sg U58206 ( .A(n53154), .X(n53155) );
  inv_x2_sg U58207 ( .A(n53156), .X(n53157) );
  inv_x2_sg U58208 ( .A(n53158), .X(n53159) );
  inv_x2_sg U58209 ( .A(n53160), .X(n53161) );
  inv_x2_sg U58210 ( .A(n53162), .X(n53163) );
  inv_x2_sg U58211 ( .A(n53164), .X(n53165) );
  inv_x2_sg U58212 ( .A(n53166), .X(n53167) );
  inv_x2_sg U58213 ( .A(n53168), .X(n53169) );
  inv_x2_sg U58214 ( .A(n53170), .X(n53171) );
  inv_x2_sg U58215 ( .A(n53172), .X(n53173) );
  inv_x2_sg U58216 ( .A(n53174), .X(n53175) );
  inv_x2_sg U58217 ( .A(n53176), .X(n53177) );
  inv_x2_sg U58218 ( .A(n53178), .X(n53179) );
  inv_x2_sg U58219 ( .A(n53180), .X(n53181) );
  inv_x2_sg U58220 ( .A(n53182), .X(n53183) );
  inv_x2_sg U58221 ( .A(n53184), .X(n53185) );
  inv_x2_sg U58222 ( .A(n53186), .X(n53187) );
  inv_x2_sg U58223 ( .A(n53188), .X(n53189) );
  inv_x2_sg U58224 ( .A(n53190), .X(n53191) );
  inv_x2_sg U58225 ( .A(n53192), .X(n53193) );
  inv_x2_sg U58226 ( .A(n53194), .X(n53195) );
  inv_x2_sg U58227 ( .A(n53196), .X(n53197) );
  inv_x2_sg U58228 ( .A(n53198), .X(n53199) );
  inv_x2_sg U58229 ( .A(n53200), .X(n53201) );
  inv_x2_sg U58230 ( .A(n53202), .X(n53203) );
  inv_x2_sg U58231 ( .A(n53204), .X(n53205) );
  inv_x2_sg U58232 ( .A(n53206), .X(n53207) );
  inv_x2_sg U58233 ( .A(n53208), .X(n53209) );
  inv_x2_sg U58234 ( .A(n53210), .X(n53211) );
  inv_x2_sg U58235 ( .A(n53212), .X(n53213) );
  inv_x2_sg U58236 ( .A(n53214), .X(n53215) );
  inv_x2_sg U58237 ( .A(n53216), .X(n53217) );
  inv_x2_sg U58238 ( .A(n53218), .X(n53219) );
  inv_x2_sg U58239 ( .A(n53220), .X(n53221) );
  inv_x2_sg U58240 ( .A(n53222), .X(n53223) );
  inv_x2_sg U58241 ( .A(n53224), .X(n53225) );
  inv_x2_sg U58242 ( .A(n53226), .X(n53227) );
  inv_x2_sg U58243 ( .A(n53228), .X(n53229) );
  inv_x2_sg U58244 ( .A(n53230), .X(n53231) );
  inv_x2_sg U58245 ( .A(n53232), .X(n53233) );
  inv_x2_sg U58246 ( .A(n53234), .X(n53235) );
  inv_x2_sg U58247 ( .A(n53236), .X(n53237) );
  inv_x2_sg U58248 ( .A(n53238), .X(n53239) );
  inv_x2_sg U58249 ( .A(n53240), .X(n53241) );
  inv_x2_sg U58250 ( .A(n53242), .X(n53243) );
  inv_x2_sg U58251 ( .A(n53244), .X(n53245) );
  inv_x2_sg U58252 ( .A(n53246), .X(n53247) );
  inv_x2_sg U58253 ( .A(n53248), .X(n53249) );
  inv_x2_sg U58254 ( .A(n53250), .X(n53251) );
  inv_x2_sg U58255 ( .A(n53252), .X(n53253) );
  inv_x2_sg U58256 ( .A(n53254), .X(n53255) );
  inv_x2_sg U58257 ( .A(n53256), .X(n53257) );
  inv_x2_sg U58258 ( .A(n53258), .X(n53259) );
  inv_x2_sg U58259 ( .A(n53260), .X(n53261) );
  inv_x2_sg U58260 ( .A(n53262), .X(n53263) );
  inv_x2_sg U58261 ( .A(n53264), .X(n53265) );
  inv_x2_sg U58262 ( .A(n53266), .X(n53267) );
  inv_x2_sg U58263 ( .A(n53268), .X(n53269) );
  inv_x2_sg U58264 ( .A(n53270), .X(n53271) );
  inv_x2_sg U58265 ( .A(n53272), .X(n53273) );
  inv_x2_sg U58266 ( .A(n53274), .X(n53275) );
  inv_x2_sg U58267 ( .A(n53276), .X(n53277) );
  inv_x2_sg U58268 ( .A(n53278), .X(n53279) );
  inv_x2_sg U58269 ( .A(n53280), .X(n53281) );
  inv_x2_sg U58270 ( .A(n53282), .X(n53283) );
  inv_x2_sg U58271 ( .A(n53284), .X(n53285) );
  inv_x2_sg U58272 ( .A(n53286), .X(n53287) );
  inv_x2_sg U58273 ( .A(n53288), .X(n53289) );
  inv_x2_sg U58274 ( .A(n53290), .X(n53291) );
  inv_x2_sg U58275 ( .A(n53292), .X(n53293) );
  inv_x2_sg U58276 ( .A(n53294), .X(n53295) );
  inv_x2_sg U58277 ( .A(n53296), .X(n53297) );
  inv_x2_sg U58278 ( .A(n53298), .X(n53299) );
  inv_x2_sg U58279 ( .A(n53300), .X(n53301) );
  inv_x2_sg U58280 ( .A(n53302), .X(n53303) );
  inv_x2_sg U58281 ( .A(n53304), .X(n53305) );
  inv_x2_sg U58282 ( .A(n53306), .X(n53307) );
  inv_x2_sg U58283 ( .A(n53308), .X(n53309) );
  inv_x2_sg U58284 ( .A(n53310), .X(n53311) );
  inv_x2_sg U58285 ( .A(n53312), .X(n53313) );
  inv_x2_sg U58286 ( .A(n53314), .X(n53315) );
  inv_x2_sg U58287 ( .A(n53316), .X(n53317) );
  inv_x2_sg U58288 ( .A(n53318), .X(n53319) );
  inv_x2_sg U58289 ( .A(n53320), .X(n53321) );
  inv_x2_sg U58290 ( .A(n53322), .X(n53323) );
  inv_x2_sg U58291 ( .A(n53324), .X(n53325) );
  inv_x2_sg U58292 ( .A(n53326), .X(n53327) );
  inv_x2_sg U58293 ( .A(n53328), .X(n53329) );
  inv_x2_sg U58294 ( .A(n53330), .X(n53331) );
  inv_x2_sg U58295 ( .A(n53332), .X(n53333) );
  inv_x2_sg U58296 ( .A(n53334), .X(n53335) );
  inv_x2_sg U58297 ( .A(n53336), .X(n53337) );
  inv_x2_sg U58298 ( .A(n53338), .X(n53339) );
  inv_x2_sg U58299 ( .A(n53340), .X(n53341) );
  inv_x2_sg U58300 ( .A(n53342), .X(n53343) );
  inv_x2_sg U58301 ( .A(n53344), .X(n53345) );
  inv_x2_sg U58302 ( .A(n53346), .X(n53347) );
  inv_x2_sg U58303 ( .A(n53348), .X(n53349) );
  inv_x2_sg U58304 ( .A(n53350), .X(n53351) );
  inv_x2_sg U58305 ( .A(n53352), .X(n53353) );
  inv_x2_sg U58306 ( .A(n53354), .X(n53355) );
  inv_x2_sg U58307 ( .A(n53356), .X(n53357) );
  inv_x2_sg U58308 ( .A(n53358), .X(n53359) );
  inv_x2_sg U58309 ( .A(n53360), .X(n53361) );
  inv_x2_sg U58310 ( .A(n53362), .X(n53363) );
  inv_x2_sg U58311 ( .A(n53364), .X(n53365) );
  inv_x2_sg U58312 ( .A(n53366), .X(n53367) );
  inv_x2_sg U58313 ( .A(n53368), .X(n53369) );
  inv_x2_sg U58314 ( .A(n53370), .X(n53371) );
  inv_x2_sg U58315 ( .A(n53372), .X(n53373) );
  inv_x2_sg U58316 ( .A(n53374), .X(n53375) );
  inv_x2_sg U58317 ( .A(n53376), .X(n53377) );
  inv_x2_sg U58318 ( .A(n53378), .X(n53379) );
  inv_x2_sg U58319 ( .A(n53380), .X(n53381) );
  inv_x2_sg U58320 ( .A(n53382), .X(n53383) );
  inv_x2_sg U58321 ( .A(n53384), .X(n53385) );
  inv_x2_sg U58322 ( .A(n53386), .X(n53387) );
  inv_x2_sg U58323 ( .A(n53388), .X(n53389) );
  inv_x2_sg U58324 ( .A(n53390), .X(n53391) );
  inv_x2_sg U58325 ( .A(n53392), .X(n53393) );
  inv_x2_sg U58326 ( .A(n53394), .X(n53395) );
  inv_x2_sg U58327 ( .A(n53396), .X(n53397) );
  inv_x2_sg U58328 ( .A(n53398), .X(n53399) );
  inv_x2_sg U58329 ( .A(n53400), .X(n53401) );
  inv_x2_sg U58330 ( .A(n53402), .X(n53403) );
  inv_x2_sg U58331 ( .A(n53404), .X(n53405) );
  inv_x2_sg U58332 ( .A(n53406), .X(n53407) );
  inv_x2_sg U58333 ( .A(n53408), .X(n53409) );
  inv_x2_sg U58334 ( .A(n53410), .X(n53411) );
  inv_x2_sg U58335 ( .A(n53412), .X(n53413) );
  inv_x2_sg U58336 ( .A(n53414), .X(n53415) );
  inv_x2_sg U58337 ( .A(n53416), .X(n53417) );
  inv_x2_sg U58338 ( .A(n53418), .X(n53419) );
  inv_x2_sg U58339 ( .A(n53420), .X(n53421) );
  inv_x2_sg U58340 ( .A(n53422), .X(n53423) );
  inv_x2_sg U58341 ( .A(n53424), .X(n53425) );
  inv_x2_sg U58342 ( .A(n53426), .X(n53427) );
  inv_x2_sg U58343 ( .A(n53428), .X(n53429) );
  inv_x2_sg U58344 ( .A(n53430), .X(n53431) );
  inv_x2_sg U58345 ( .A(n53432), .X(n53433) );
  inv_x2_sg U58346 ( .A(n53434), .X(n53435) );
  inv_x2_sg U58347 ( .A(n53436), .X(n53437) );
  inv_x2_sg U58348 ( .A(n53438), .X(n53439) );
  inv_x2_sg U58349 ( .A(n53440), .X(n53441) );
  inv_x2_sg U58350 ( .A(n53442), .X(n53443) );
  inv_x2_sg U58351 ( .A(n53444), .X(n53445) );
  inv_x2_sg U58352 ( .A(n53446), .X(n53447) );
  inv_x2_sg U58353 ( .A(n53448), .X(n53449) );
  inv_x2_sg U58354 ( .A(n53450), .X(n53451) );
  inv_x2_sg U58355 ( .A(n53452), .X(n53453) );
  inv_x2_sg U58356 ( .A(n53454), .X(n53455) );
  inv_x2_sg U58357 ( .A(n53456), .X(n53457) );
  inv_x2_sg U58358 ( .A(n53458), .X(n53459) );
  inv_x2_sg U58359 ( .A(n53460), .X(n53461) );
  inv_x2_sg U58360 ( .A(n53462), .X(n53463) );
  inv_x2_sg U58361 ( .A(n53464), .X(n53465) );
  inv_x2_sg U58362 ( .A(n53466), .X(n53467) );
  inv_x2_sg U58363 ( .A(n53468), .X(n53469) );
  inv_x2_sg U58364 ( .A(n53470), .X(n53471) );
  inv_x2_sg U58365 ( .A(n53472), .X(n53473) );
  inv_x2_sg U58366 ( .A(n53474), .X(n53475) );
  inv_x2_sg U58367 ( .A(n53476), .X(n53477) );
  inv_x2_sg U58368 ( .A(n53478), .X(n53479) );
  inv_x2_sg U58369 ( .A(n53480), .X(n53481) );
  inv_x2_sg U58370 ( .A(n53482), .X(n53483) );
  inv_x2_sg U58371 ( .A(n53484), .X(n53485) );
  inv_x2_sg U58372 ( .A(n53486), .X(n53487) );
  inv_x2_sg U58373 ( .A(n53488), .X(n53489) );
  inv_x2_sg U58374 ( .A(n53490), .X(n53491) );
  inv_x2_sg U58375 ( .A(n53492), .X(n53493) );
  inv_x2_sg U58376 ( .A(n53494), .X(n53495) );
  inv_x2_sg U58377 ( .A(n53496), .X(n53497) );
  inv_x2_sg U58378 ( .A(n53498), .X(n53499) );
  inv_x2_sg U58379 ( .A(n53500), .X(n53501) );
  inv_x2_sg U58380 ( .A(n53502), .X(n53503) );
  inv_x2_sg U58381 ( .A(n53504), .X(n53505) );
  inv_x2_sg U58382 ( .A(n53506), .X(n53507) );
  inv_x2_sg U58383 ( .A(n53508), .X(n53509) );
  inv_x2_sg U58384 ( .A(n53510), .X(n53511) );
  inv_x2_sg U58385 ( .A(n53512), .X(n53513) );
  inv_x2_sg U58386 ( .A(n53514), .X(n53515) );
  inv_x2_sg U58387 ( .A(n53516), .X(n53517) );
  inv_x2_sg U58388 ( .A(n53518), .X(n53519) );
  inv_x2_sg U58389 ( .A(n53520), .X(n53521) );
  inv_x2_sg U58390 ( .A(n53522), .X(n53523) );
  inv_x2_sg U58391 ( .A(n53524), .X(n53525) );
  inv_x2_sg U58392 ( .A(n53526), .X(n53527) );
  inv_x2_sg U58393 ( .A(n53528), .X(n53529) );
  inv_x2_sg U58394 ( .A(n53530), .X(n53531) );
  inv_x2_sg U58395 ( .A(n53532), .X(n53533) );
  inv_x2_sg U58396 ( .A(n53534), .X(n53535) );
  inv_x2_sg U58397 ( .A(n53536), .X(n53537) );
  inv_x2_sg U58398 ( .A(n53538), .X(n53539) );
  inv_x2_sg U58399 ( .A(n53540), .X(n53541) );
  inv_x2_sg U58400 ( .A(n53542), .X(n53543) );
  inv_x2_sg U58401 ( .A(n53544), .X(n53545) );
  inv_x2_sg U58402 ( .A(n53546), .X(n53547) );
  inv_x2_sg U58403 ( .A(n53548), .X(n53549) );
  inv_x2_sg U58404 ( .A(n53550), .X(n53551) );
  inv_x2_sg U58405 ( .A(n53552), .X(n53553) );
  inv_x2_sg U58406 ( .A(n53554), .X(n53555) );
  inv_x2_sg U58407 ( .A(n53556), .X(n53557) );
  inv_x2_sg U58408 ( .A(n53558), .X(n53559) );
  inv_x2_sg U58409 ( .A(n53560), .X(n53561) );
  inv_x2_sg U58410 ( .A(n53562), .X(n53563) );
  inv_x2_sg U58411 ( .A(n53564), .X(n53565) );
  inv_x2_sg U58412 ( .A(n53566), .X(n53567) );
  inv_x2_sg U58413 ( .A(n53568), .X(n53569) );
  inv_x2_sg U58414 ( .A(n53570), .X(n53571) );
  inv_x2_sg U58415 ( .A(n53572), .X(n53573) );
  inv_x2_sg U58416 ( .A(n53574), .X(n53575) );
  inv_x2_sg U58417 ( .A(n53576), .X(n53577) );
  inv_x2_sg U58418 ( .A(n53578), .X(n53579) );
  inv_x2_sg U58419 ( .A(n53580), .X(n53581) );
  inv_x2_sg U58420 ( .A(n53582), .X(n53583) );
  inv_x2_sg U58421 ( .A(n53584), .X(n53585) );
  inv_x2_sg U58422 ( .A(n53586), .X(n53587) );
  inv_x2_sg U58423 ( .A(n53588), .X(n53589) );
  inv_x2_sg U58424 ( .A(n53590), .X(n53591) );
  inv_x2_sg U58425 ( .A(n53592), .X(n53593) );
  inv_x2_sg U58426 ( .A(n53594), .X(n53595) );
  inv_x2_sg U58427 ( .A(n53596), .X(n53597) );
  inv_x2_sg U58428 ( .A(n53598), .X(n53599) );
  inv_x2_sg U58429 ( .A(n53600), .X(n53601) );
  inv_x2_sg U58430 ( .A(n53602), .X(n53603) );
  inv_x2_sg U58431 ( .A(n53604), .X(n53605) );
  inv_x2_sg U58432 ( .A(n53606), .X(n53607) );
  inv_x2_sg U58433 ( .A(n53608), .X(n53609) );
  inv_x2_sg U58434 ( .A(n53610), .X(n53611) );
  inv_x2_sg U58435 ( .A(n53612), .X(n53613) );
  inv_x2_sg U58436 ( .A(n53614), .X(n53615) );
  inv_x2_sg U58437 ( .A(n53616), .X(n53617) );
  inv_x2_sg U58438 ( .A(n53618), .X(n53619) );
  inv_x2_sg U58439 ( .A(n53620), .X(n53621) );
  inv_x2_sg U58440 ( .A(n53622), .X(n53623) );
  inv_x2_sg U58441 ( .A(n53624), .X(n53625) );
  inv_x2_sg U58442 ( .A(n53626), .X(n53627) );
  inv_x2_sg U58443 ( .A(n53628), .X(n53629) );
  inv_x2_sg U58444 ( .A(n53630), .X(n53631) );
  inv_x2_sg U58445 ( .A(n53632), .X(n53633) );
  inv_x2_sg U58446 ( .A(n53634), .X(n53635) );
  inv_x2_sg U58447 ( .A(n53636), .X(n53637) );
  inv_x2_sg U58448 ( .A(n53638), .X(n53639) );
  inv_x2_sg U58449 ( .A(n53640), .X(n53641) );
  inv_x2_sg U58450 ( .A(n53642), .X(n53643) );
  inv_x2_sg U58451 ( .A(n53644), .X(n53645) );
  inv_x2_sg U58452 ( .A(n53646), .X(n53647) );
  inv_x4_sg U58453 ( .A(n22644), .X(n67375) );
  inv_x4_sg U58454 ( .A(n22641), .X(n67378) );
  inv_x4_sg U58455 ( .A(n22638), .X(n67381) );
  inv_x4_sg U58456 ( .A(n22636), .X(n67383) );
  inv_x4_sg U58457 ( .A(n22634), .X(n67385) );
  inv_x4_sg U58458 ( .A(n22632), .X(n67387) );
  inv_x4_sg U58459 ( .A(n22630), .X(n67389) );
  inv_x4_sg U58460 ( .A(n22629), .X(n67390) );
  inv_x4_sg U58461 ( .A(n22626), .X(n67393) );
  inv_x4_sg U58462 ( .A(n22625), .X(n67394) );
  inv_x4_sg U58463 ( .A(n22617), .X(n67162) );
  inv_x4_sg U58464 ( .A(n22614), .X(n67165) );
  inv_x4_sg U58465 ( .A(n22611), .X(n67168) );
  inv_x4_sg U58466 ( .A(n22609), .X(n67170) );
  inv_x4_sg U58467 ( .A(n22607), .X(n67172) );
  inv_x4_sg U58468 ( .A(n22605), .X(n67174) );
  inv_x4_sg U58469 ( .A(n22603), .X(n67176) );
  inv_x4_sg U58470 ( .A(n22602), .X(n67177) );
  inv_x4_sg U58471 ( .A(n22599), .X(n67180) );
  inv_x4_sg U58472 ( .A(n22598), .X(n67181) );
  inv_x2_sg U58473 ( .A(n53648), .X(n53649) );
  inv_x2_sg U58474 ( .A(n53650), .X(n53651) );
  inv_x2_sg U58475 ( .A(n53652), .X(n53653) );
  inv_x2_sg U58476 ( .A(n53654), .X(n53655) );
  inv_x2_sg U58477 ( .A(n53656), .X(n53657) );
  inv_x2_sg U58478 ( .A(n53658), .X(n53659) );
  inv_x2_sg U58479 ( .A(n53660), .X(n53661) );
  inv_x2_sg U58480 ( .A(n53662), .X(n53663) );
  inv_x2_sg U58481 ( .A(n53664), .X(n53665) );
  inv_x2_sg U58482 ( .A(n53666), .X(n53667) );
  inv_x2_sg U58483 ( .A(n53668), .X(n53669) );
  inv_x2_sg U58484 ( .A(n53670), .X(n53671) );
  inv_x2_sg U58485 ( .A(n53672), .X(n53673) );
  inv_x2_sg U58486 ( .A(n53674), .X(n53675) );
  inv_x2_sg U58487 ( .A(n53676), .X(n53677) );
  inv_x2_sg U58488 ( .A(n53678), .X(n53679) );
  inv_x2_sg U58489 ( .A(n53680), .X(n53681) );
  inv_x2_sg U58490 ( .A(n53682), .X(n53683) );
  inv_x2_sg U58491 ( .A(n53684), .X(n53685) );
  inv_x2_sg U58492 ( .A(n53686), .X(n53687) );
  inv_x2_sg U58493 ( .A(n53688), .X(n53689) );
  inv_x2_sg U58494 ( .A(n53690), .X(n53691) );
  inv_x2_sg U58495 ( .A(n53692), .X(n53693) );
  inv_x2_sg U58496 ( .A(n53694), .X(n53695) );
  inv_x2_sg U58497 ( .A(n53696), .X(n53697) );
  inv_x2_sg U58498 ( .A(n53698), .X(n53699) );
  inv_x2_sg U58499 ( .A(n53700), .X(n53701) );
  inv_x2_sg U58500 ( .A(n53702), .X(n53703) );
  inv_x2_sg U58501 ( .A(n53704), .X(n53705) );
  inv_x2_sg U58502 ( .A(n53706), .X(n53707) );
  inv_x2_sg U58503 ( .A(n53708), .X(n53709) );
  inv_x2_sg U58504 ( .A(n53710), .X(n53711) );
  inv_x4_sg U58505 ( .A(n53714), .X(n53715) );
  nor_x4_sg U58506 ( .A(n67530), .B(n67534), .X(n26091) );
  inv_x4_sg U58507 ( .A(n53716), .X(n53717) );
  nand_x8_sg U58508 ( .A(n24261), .B(n23308), .X(n24260) );
  nor_x2_sg U58509 ( .A(n57918), .B(n68571), .X(n24261) );
  inv_x8_sg U58510 ( .A(n29336), .X(n68571) );
  inv_x2_sg U58511 ( .A(n53718), .X(ow_14[0]) );
  inv_x2_sg U58512 ( .A(n53720), .X(ow_14[1]) );
  inv_x2_sg U58513 ( .A(n53722), .X(ow_14[2]) );
  inv_x2_sg U58514 ( .A(n53724), .X(ow_14[3]) );
  inv_x2_sg U58515 ( .A(n53726), .X(ow_14[4]) );
  inv_x2_sg U58516 ( .A(n53728), .X(ow_14[5]) );
  inv_x2_sg U58517 ( .A(n53730), .X(ow_14[6]) );
  inv_x2_sg U58518 ( .A(n53732), .X(ow_14[7]) );
  inv_x2_sg U58519 ( .A(n53734), .X(ow_14[8]) );
  inv_x2_sg U58520 ( .A(n53736), .X(ow_14[9]) );
  inv_x2_sg U58521 ( .A(n53738), .X(ow_14[10]) );
  inv_x2_sg U58522 ( .A(n53740), .X(ow_14[11]) );
  inv_x2_sg U58523 ( .A(n53742), .X(ow_14[12]) );
  inv_x2_sg U58524 ( .A(n53744), .X(ow_14[13]) );
  inv_x2_sg U58525 ( .A(n53746), .X(ow_14[14]) );
  inv_x2_sg U58526 ( .A(n53748), .X(ow_14[15]) );
  inv_x2_sg U58527 ( .A(n53750), .X(ow_14[16]) );
  inv_x2_sg U58528 ( .A(n53752), .X(ow_14[17]) );
  inv_x2_sg U58529 ( .A(n53754), .X(ow_14[18]) );
  inv_x2_sg U58530 ( .A(n53756), .X(ow_14[19]) );
  inv_x2_sg U58531 ( .A(n53758), .X(ow_13[0]) );
  inv_x2_sg U58532 ( .A(n53760), .X(ow_13[1]) );
  inv_x2_sg U58533 ( .A(n53762), .X(ow_13[2]) );
  inv_x2_sg U58534 ( .A(n53764), .X(ow_13[3]) );
  inv_x2_sg U58535 ( .A(n53766), .X(ow_13[4]) );
  inv_x2_sg U58536 ( .A(n53768), .X(ow_13[5]) );
  inv_x2_sg U58537 ( .A(n53770), .X(ow_13[6]) );
  inv_x2_sg U58538 ( .A(n53772), .X(ow_13[7]) );
  inv_x2_sg U58539 ( .A(n53774), .X(ow_13[8]) );
  inv_x2_sg U58540 ( .A(n53776), .X(ow_13[9]) );
  inv_x2_sg U58541 ( .A(n53778), .X(ow_13[10]) );
  inv_x2_sg U58542 ( .A(n53780), .X(ow_13[11]) );
  inv_x2_sg U58543 ( .A(n53782), .X(ow_13[12]) );
  inv_x2_sg U58544 ( .A(n53784), .X(ow_13[13]) );
  inv_x2_sg U58545 ( .A(n53786), .X(ow_13[14]) );
  inv_x2_sg U58546 ( .A(n53788), .X(ow_13[15]) );
  inv_x2_sg U58547 ( .A(n53790), .X(ow_13[16]) );
  inv_x2_sg U58548 ( .A(n53792), .X(ow_13[17]) );
  inv_x2_sg U58549 ( .A(n53794), .X(ow_13[18]) );
  inv_x2_sg U58550 ( .A(n53796), .X(ow_13[19]) );
  inv_x2_sg U58551 ( .A(n53798), .X(ow_12[0]) );
  inv_x2_sg U58552 ( .A(n53800), .X(ow_12[1]) );
  inv_x2_sg U58553 ( .A(n53802), .X(ow_12[2]) );
  inv_x2_sg U58554 ( .A(n53804), .X(ow_12[3]) );
  inv_x2_sg U58555 ( .A(n53806), .X(ow_12[4]) );
  inv_x2_sg U58556 ( .A(n53808), .X(ow_12[5]) );
  inv_x2_sg U58557 ( .A(n53810), .X(ow_12[6]) );
  inv_x2_sg U58558 ( .A(n53812), .X(ow_12[7]) );
  inv_x2_sg U58559 ( .A(n53814), .X(ow_12[8]) );
  inv_x2_sg U58560 ( .A(n53816), .X(ow_12[9]) );
  inv_x2_sg U58561 ( .A(n53818), .X(ow_12[10]) );
  inv_x2_sg U58562 ( .A(n53820), .X(ow_12[11]) );
  inv_x2_sg U58563 ( .A(n53822), .X(ow_12[12]) );
  inv_x2_sg U58564 ( .A(n53824), .X(ow_12[13]) );
  inv_x2_sg U58565 ( .A(n53826), .X(ow_12[14]) );
  inv_x2_sg U58566 ( .A(n53828), .X(ow_12[15]) );
  inv_x2_sg U58567 ( .A(n53830), .X(ow_12[16]) );
  inv_x2_sg U58568 ( .A(n53832), .X(ow_12[17]) );
  inv_x2_sg U58569 ( .A(n53834), .X(ow_12[18]) );
  inv_x2_sg U58570 ( .A(n53836), .X(ow_12[19]) );
  inv_x2_sg U58571 ( .A(n53838), .X(ow_11[0]) );
  inv_x2_sg U58572 ( .A(n53840), .X(ow_11[1]) );
  inv_x2_sg U58573 ( .A(n53842), .X(ow_11[2]) );
  inv_x2_sg U58574 ( .A(n53844), .X(ow_11[3]) );
  inv_x2_sg U58575 ( .A(n53846), .X(ow_11[4]) );
  inv_x2_sg U58576 ( .A(n53848), .X(ow_11[5]) );
  inv_x2_sg U58577 ( .A(n53850), .X(ow_11[6]) );
  inv_x2_sg U58578 ( .A(n53852), .X(ow_11[7]) );
  inv_x2_sg U58579 ( .A(n53854), .X(ow_11[8]) );
  inv_x2_sg U58580 ( .A(n53856), .X(ow_11[9]) );
  inv_x2_sg U58581 ( .A(n53858), .X(ow_11[10]) );
  inv_x2_sg U58582 ( .A(n53860), .X(ow_11[11]) );
  inv_x2_sg U58583 ( .A(n53862), .X(ow_11[12]) );
  inv_x2_sg U58584 ( .A(n53864), .X(ow_11[13]) );
  inv_x2_sg U58585 ( .A(n53866), .X(ow_11[14]) );
  inv_x2_sg U58586 ( .A(n53868), .X(ow_11[15]) );
  inv_x2_sg U58587 ( .A(n53870), .X(ow_11[16]) );
  inv_x2_sg U58588 ( .A(n53872), .X(ow_11[17]) );
  inv_x2_sg U58589 ( .A(n53874), .X(ow_11[18]) );
  inv_x2_sg U58590 ( .A(n53876), .X(ow_11[19]) );
  inv_x2_sg U58591 ( .A(n53878), .X(ow_10[0]) );
  inv_x2_sg U58592 ( .A(n53880), .X(ow_10[1]) );
  inv_x2_sg U58593 ( .A(n53882), .X(ow_10[2]) );
  inv_x2_sg U58594 ( .A(n53884), .X(ow_10[3]) );
  inv_x2_sg U58595 ( .A(n53886), .X(ow_10[4]) );
  inv_x2_sg U58596 ( .A(n53888), .X(ow_10[5]) );
  inv_x2_sg U58597 ( .A(n53890), .X(ow_10[6]) );
  inv_x2_sg U58598 ( .A(n53892), .X(ow_10[7]) );
  inv_x2_sg U58599 ( .A(n53894), .X(ow_10[8]) );
  inv_x2_sg U58600 ( .A(n53896), .X(ow_10[9]) );
  inv_x2_sg U58601 ( .A(n53898), .X(ow_10[10]) );
  inv_x2_sg U58602 ( .A(n53900), .X(ow_10[11]) );
  inv_x2_sg U58603 ( .A(n53902), .X(ow_10[12]) );
  inv_x2_sg U58604 ( .A(n53904), .X(ow_10[13]) );
  inv_x2_sg U58605 ( .A(n53906), .X(ow_10[14]) );
  inv_x2_sg U58606 ( .A(n53908), .X(ow_10[15]) );
  inv_x2_sg U58607 ( .A(n53910), .X(ow_10[16]) );
  inv_x2_sg U58608 ( .A(n53912), .X(ow_10[17]) );
  inv_x2_sg U58609 ( .A(n53914), .X(ow_10[18]) );
  inv_x2_sg U58610 ( .A(n53916), .X(ow_10[19]) );
  inv_x2_sg U58611 ( .A(n53918), .X(ow_9[0]) );
  inv_x2_sg U58612 ( .A(n53920), .X(ow_9[1]) );
  inv_x2_sg U58613 ( .A(n53922), .X(ow_9[2]) );
  inv_x2_sg U58614 ( .A(n53924), .X(ow_9[3]) );
  inv_x2_sg U58615 ( .A(n53926), .X(ow_9[4]) );
  inv_x2_sg U58616 ( .A(n53928), .X(ow_9[5]) );
  inv_x2_sg U58617 ( .A(n53930), .X(ow_9[6]) );
  inv_x2_sg U58618 ( .A(n53932), .X(ow_9[7]) );
  inv_x2_sg U58619 ( .A(n53934), .X(ow_9[8]) );
  inv_x2_sg U58620 ( .A(n53936), .X(ow_9[9]) );
  inv_x2_sg U58621 ( .A(n53938), .X(ow_9[10]) );
  inv_x2_sg U58622 ( .A(n53940), .X(ow_9[11]) );
  inv_x2_sg U58623 ( .A(n53942), .X(ow_9[12]) );
  inv_x2_sg U58624 ( .A(n53944), .X(ow_9[13]) );
  inv_x2_sg U58625 ( .A(n53946), .X(ow_9[14]) );
  inv_x2_sg U58626 ( .A(n53948), .X(ow_9[15]) );
  inv_x2_sg U58627 ( .A(n53950), .X(ow_9[16]) );
  inv_x2_sg U58628 ( .A(n53952), .X(ow_9[17]) );
  inv_x2_sg U58629 ( .A(n53954), .X(ow_9[18]) );
  inv_x2_sg U58630 ( .A(n53956), .X(ow_9[19]) );
  inv_x2_sg U58631 ( .A(n53958), .X(ow_8[0]) );
  inv_x2_sg U58632 ( .A(n53960), .X(ow_8[1]) );
  inv_x2_sg U58633 ( .A(n53962), .X(ow_8[2]) );
  inv_x2_sg U58634 ( .A(n53964), .X(ow_8[3]) );
  inv_x2_sg U58635 ( .A(n53966), .X(ow_8[4]) );
  inv_x2_sg U58636 ( .A(n53968), .X(ow_8[5]) );
  inv_x2_sg U58637 ( .A(n53970), .X(ow_8[6]) );
  inv_x2_sg U58638 ( .A(n53972), .X(ow_8[7]) );
  inv_x2_sg U58639 ( .A(n53974), .X(ow_8[8]) );
  inv_x2_sg U58640 ( .A(n53976), .X(ow_8[9]) );
  inv_x2_sg U58641 ( .A(n53978), .X(ow_8[10]) );
  inv_x2_sg U58642 ( .A(n53980), .X(ow_8[11]) );
  inv_x2_sg U58643 ( .A(n53982), .X(ow_8[12]) );
  inv_x2_sg U58644 ( .A(n53984), .X(ow_8[13]) );
  inv_x2_sg U58645 ( .A(n53986), .X(ow_8[14]) );
  inv_x2_sg U58646 ( .A(n53988), .X(ow_8[15]) );
  inv_x2_sg U58647 ( .A(n53990), .X(ow_8[16]) );
  inv_x2_sg U58648 ( .A(n53992), .X(ow_8[17]) );
  inv_x2_sg U58649 ( .A(n53994), .X(ow_8[18]) );
  inv_x2_sg U58650 ( .A(n53996), .X(ow_8[19]) );
  inv_x2_sg U58651 ( .A(n53998), .X(ow_7[0]) );
  inv_x2_sg U58652 ( .A(n54000), .X(ow_7[1]) );
  inv_x2_sg U58653 ( .A(n54002), .X(ow_7[2]) );
  inv_x2_sg U58654 ( .A(n54004), .X(ow_7[3]) );
  inv_x2_sg U58655 ( .A(n54006), .X(ow_7[4]) );
  inv_x2_sg U58656 ( .A(n54008), .X(ow_7[5]) );
  inv_x2_sg U58657 ( .A(n54010), .X(ow_7[6]) );
  inv_x2_sg U58658 ( .A(n54012), .X(ow_7[7]) );
  inv_x2_sg U58659 ( .A(n54014), .X(ow_7[8]) );
  inv_x2_sg U58660 ( .A(n54016), .X(ow_7[9]) );
  inv_x2_sg U58661 ( .A(n54018), .X(ow_7[10]) );
  inv_x2_sg U58662 ( .A(n54020), .X(ow_7[11]) );
  inv_x2_sg U58663 ( .A(n54022), .X(ow_7[12]) );
  inv_x2_sg U58664 ( .A(n54024), .X(ow_7[13]) );
  inv_x2_sg U58665 ( .A(n54026), .X(ow_7[14]) );
  inv_x2_sg U58666 ( .A(n54028), .X(ow_7[15]) );
  inv_x2_sg U58667 ( .A(n54030), .X(ow_7[16]) );
  inv_x2_sg U58668 ( .A(n54032), .X(ow_7[17]) );
  inv_x2_sg U58669 ( .A(n54034), .X(ow_7[18]) );
  inv_x2_sg U58670 ( .A(n54036), .X(ow_7[19]) );
  inv_x2_sg U58671 ( .A(n54038), .X(ow_6[0]) );
  inv_x2_sg U58672 ( .A(n54040), .X(ow_6[1]) );
  inv_x2_sg U58673 ( .A(n54042), .X(ow_6[2]) );
  inv_x2_sg U58674 ( .A(n54044), .X(ow_6[3]) );
  inv_x2_sg U58675 ( .A(n54046), .X(ow_6[4]) );
  inv_x2_sg U58676 ( .A(n54048), .X(ow_6[5]) );
  inv_x2_sg U58677 ( .A(n54050), .X(ow_6[6]) );
  inv_x2_sg U58678 ( .A(n54052), .X(ow_6[7]) );
  inv_x2_sg U58679 ( .A(n54054), .X(ow_6[8]) );
  inv_x2_sg U58680 ( .A(n54056), .X(ow_6[9]) );
  inv_x2_sg U58681 ( .A(n54058), .X(ow_6[10]) );
  inv_x2_sg U58682 ( .A(n54060), .X(ow_6[11]) );
  inv_x2_sg U58683 ( .A(n54062), .X(ow_6[12]) );
  inv_x2_sg U58684 ( .A(n54064), .X(ow_6[13]) );
  inv_x2_sg U58685 ( .A(n54066), .X(ow_6[14]) );
  inv_x2_sg U58686 ( .A(n54068), .X(ow_6[15]) );
  inv_x2_sg U58687 ( .A(n54070), .X(ow_6[16]) );
  inv_x2_sg U58688 ( .A(n54072), .X(ow_6[17]) );
  inv_x2_sg U58689 ( .A(n54074), .X(ow_6[18]) );
  inv_x2_sg U58690 ( .A(n54076), .X(ow_6[19]) );
  inv_x2_sg U58691 ( .A(n54078), .X(ow_5[0]) );
  inv_x2_sg U58692 ( .A(n54080), .X(ow_5[1]) );
  inv_x2_sg U58693 ( .A(n54082), .X(ow_5[2]) );
  inv_x2_sg U58694 ( .A(n54084), .X(ow_5[3]) );
  inv_x2_sg U58695 ( .A(n54086), .X(ow_5[4]) );
  inv_x2_sg U58696 ( .A(n54088), .X(ow_5[5]) );
  inv_x2_sg U58697 ( .A(n54090), .X(ow_5[6]) );
  inv_x2_sg U58698 ( .A(n54092), .X(ow_5[7]) );
  inv_x2_sg U58699 ( .A(n54094), .X(ow_5[8]) );
  inv_x2_sg U58700 ( .A(n54096), .X(ow_5[9]) );
  inv_x2_sg U58701 ( .A(n54098), .X(ow_5[10]) );
  inv_x2_sg U58702 ( .A(n54100), .X(ow_5[11]) );
  inv_x2_sg U58703 ( .A(n54102), .X(ow_5[12]) );
  inv_x2_sg U58704 ( .A(n54104), .X(ow_5[13]) );
  inv_x2_sg U58705 ( .A(n54106), .X(ow_5[14]) );
  inv_x2_sg U58706 ( .A(n54108), .X(ow_5[15]) );
  inv_x2_sg U58707 ( .A(n54110), .X(ow_5[16]) );
  inv_x2_sg U58708 ( .A(n54112), .X(ow_5[17]) );
  inv_x2_sg U58709 ( .A(n54114), .X(ow_5[18]) );
  inv_x2_sg U58710 ( .A(n54116), .X(ow_5[19]) );
  inv_x2_sg U58711 ( .A(n54118), .X(ow_4[0]) );
  inv_x2_sg U58712 ( .A(n54120), .X(ow_4[1]) );
  inv_x2_sg U58713 ( .A(n54122), .X(ow_4[2]) );
  inv_x2_sg U58714 ( .A(n54124), .X(ow_4[3]) );
  inv_x2_sg U58715 ( .A(n54126), .X(ow_4[4]) );
  inv_x2_sg U58716 ( .A(n54128), .X(ow_4[5]) );
  inv_x2_sg U58717 ( .A(n54130), .X(ow_4[6]) );
  inv_x2_sg U58718 ( .A(n54132), .X(ow_4[7]) );
  inv_x2_sg U58719 ( .A(n54134), .X(ow_4[8]) );
  inv_x2_sg U58720 ( .A(n54136), .X(ow_4[9]) );
  inv_x2_sg U58721 ( .A(n54138), .X(ow_4[10]) );
  inv_x2_sg U58722 ( .A(n54140), .X(ow_4[11]) );
  inv_x2_sg U58723 ( .A(n54142), .X(ow_4[12]) );
  inv_x2_sg U58724 ( .A(n54144), .X(ow_4[13]) );
  inv_x2_sg U58725 ( .A(n54146), .X(ow_4[14]) );
  inv_x2_sg U58726 ( .A(n54148), .X(ow_4[15]) );
  inv_x2_sg U58727 ( .A(n54150), .X(ow_4[16]) );
  inv_x2_sg U58728 ( .A(n54152), .X(ow_4[17]) );
  inv_x2_sg U58729 ( .A(n54154), .X(ow_4[18]) );
  inv_x2_sg U58730 ( .A(n54156), .X(ow_4[19]) );
  inv_x2_sg U58731 ( .A(n54158), .X(ow_3[0]) );
  inv_x2_sg U58732 ( .A(n54160), .X(ow_3[1]) );
  inv_x2_sg U58733 ( .A(n54162), .X(ow_3[2]) );
  inv_x2_sg U58734 ( .A(n54164), .X(ow_3[3]) );
  inv_x2_sg U58735 ( .A(n54166), .X(ow_3[4]) );
  inv_x2_sg U58736 ( .A(n54168), .X(ow_3[5]) );
  inv_x2_sg U58737 ( .A(n54170), .X(ow_3[6]) );
  inv_x2_sg U58738 ( .A(n54172), .X(ow_3[7]) );
  inv_x2_sg U58739 ( .A(n54174), .X(ow_3[8]) );
  inv_x2_sg U58740 ( .A(n54176), .X(ow_3[9]) );
  inv_x2_sg U58741 ( .A(n54178), .X(ow_3[10]) );
  inv_x2_sg U58742 ( .A(n54180), .X(ow_3[11]) );
  inv_x2_sg U58743 ( .A(n54182), .X(ow_3[12]) );
  inv_x2_sg U58744 ( .A(n54184), .X(ow_3[13]) );
  inv_x2_sg U58745 ( .A(n54186), .X(ow_3[14]) );
  inv_x2_sg U58746 ( .A(n54188), .X(ow_3[15]) );
  inv_x2_sg U58747 ( .A(n54190), .X(ow_3[16]) );
  inv_x2_sg U58748 ( .A(n54192), .X(ow_3[17]) );
  inv_x2_sg U58749 ( .A(n54194), .X(ow_3[18]) );
  inv_x2_sg U58750 ( .A(n54196), .X(ow_3[19]) );
  inv_x2_sg U58751 ( .A(n54198), .X(ow_2[0]) );
  inv_x2_sg U58752 ( .A(n54200), .X(ow_2[1]) );
  inv_x2_sg U58753 ( .A(n54202), .X(ow_2[2]) );
  inv_x2_sg U58754 ( .A(n54204), .X(ow_2[3]) );
  inv_x2_sg U58755 ( .A(n54206), .X(ow_2[4]) );
  inv_x2_sg U58756 ( .A(n54208), .X(ow_2[5]) );
  inv_x2_sg U58757 ( .A(n54210), .X(ow_2[6]) );
  inv_x2_sg U58758 ( .A(n54212), .X(ow_2[7]) );
  inv_x2_sg U58759 ( .A(n54214), .X(ow_2[8]) );
  inv_x2_sg U58760 ( .A(n54216), .X(ow_2[9]) );
  inv_x2_sg U58761 ( .A(n54218), .X(ow_2[10]) );
  inv_x2_sg U58762 ( .A(n54220), .X(ow_2[11]) );
  inv_x2_sg U58763 ( .A(n54222), .X(ow_2[12]) );
  inv_x2_sg U58764 ( .A(n54224), .X(ow_2[13]) );
  inv_x2_sg U58765 ( .A(n54226), .X(ow_2[14]) );
  inv_x2_sg U58766 ( .A(n54228), .X(ow_2[15]) );
  inv_x2_sg U58767 ( .A(n54230), .X(ow_2[16]) );
  inv_x2_sg U58768 ( .A(n54232), .X(ow_2[17]) );
  inv_x2_sg U58769 ( .A(n54234), .X(ow_2[18]) );
  inv_x2_sg U58770 ( .A(n54236), .X(ow_2[19]) );
  inv_x2_sg U58771 ( .A(n54238), .X(ow_1[0]) );
  inv_x2_sg U58772 ( .A(n54240), .X(ow_1[1]) );
  inv_x2_sg U58773 ( .A(n54242), .X(ow_1[2]) );
  inv_x2_sg U58774 ( .A(n54244), .X(ow_1[3]) );
  inv_x2_sg U58775 ( .A(n54246), .X(ow_1[4]) );
  inv_x2_sg U58776 ( .A(n54248), .X(ow_1[5]) );
  inv_x2_sg U58777 ( .A(n54250), .X(ow_1[6]) );
  inv_x2_sg U58778 ( .A(n54252), .X(ow_1[7]) );
  inv_x2_sg U58779 ( .A(n54254), .X(ow_1[8]) );
  inv_x2_sg U58780 ( .A(n54256), .X(ow_1[9]) );
  inv_x2_sg U58781 ( .A(n54258), .X(ow_1[10]) );
  inv_x2_sg U58782 ( .A(n54260), .X(ow_1[11]) );
  inv_x2_sg U58783 ( .A(n54262), .X(ow_1[12]) );
  inv_x2_sg U58784 ( .A(n54264), .X(ow_1[13]) );
  inv_x2_sg U58785 ( .A(n54266), .X(ow_1[14]) );
  inv_x2_sg U58786 ( .A(n54268), .X(ow_1[15]) );
  inv_x2_sg U58787 ( .A(n54270), .X(ow_1[16]) );
  inv_x2_sg U58788 ( .A(n54272), .X(ow_1[17]) );
  inv_x2_sg U58789 ( .A(n54274), .X(ow_1[18]) );
  inv_x2_sg U58790 ( .A(n54276), .X(ow_1[19]) );
  inv_x2_sg U58791 ( .A(n54278), .X(ow_0[0]) );
  inv_x2_sg U58792 ( .A(n54280), .X(ow_0[1]) );
  inv_x2_sg U58793 ( .A(n54282), .X(ow_0[2]) );
  inv_x2_sg U58794 ( .A(n54284), .X(ow_0[3]) );
  inv_x2_sg U58795 ( .A(n54286), .X(ow_0[4]) );
  inv_x2_sg U58796 ( .A(n54288), .X(ow_0[5]) );
  inv_x2_sg U58797 ( .A(n54290), .X(ow_0[6]) );
  inv_x2_sg U58798 ( .A(n54292), .X(ow_0[7]) );
  inv_x2_sg U58799 ( .A(n54294), .X(ow_0[8]) );
  inv_x2_sg U58800 ( .A(n54296), .X(ow_0[9]) );
  inv_x2_sg U58801 ( .A(n54298), .X(ow_0[10]) );
  inv_x2_sg U58802 ( .A(n54300), .X(ow_0[11]) );
  inv_x2_sg U58803 ( .A(n54302), .X(ow_0[12]) );
  inv_x2_sg U58804 ( .A(n54304), .X(ow_0[13]) );
  inv_x2_sg U58805 ( .A(n54306), .X(ow_0[14]) );
  inv_x2_sg U58806 ( .A(n54308), .X(ow_0[15]) );
  inv_x2_sg U58807 ( .A(n54310), .X(ow_0[16]) );
  inv_x2_sg U58808 ( .A(n54312), .X(ow_0[17]) );
  inv_x2_sg U58809 ( .A(n54314), .X(ow_0[18]) );
  inv_x2_sg U58810 ( .A(n54316), .X(ow_0[19]) );
  inv_x2_sg U58811 ( .A(n54318), .X(oi_15[0]) );
  inv_x2_sg U58812 ( .A(n54320), .X(oi_15[1]) );
  inv_x2_sg U58813 ( .A(n54322), .X(oi_15[2]) );
  inv_x2_sg U58814 ( .A(n54324), .X(oi_15[3]) );
  inv_x2_sg U58815 ( .A(n54326), .X(oi_15[4]) );
  inv_x2_sg U58816 ( .A(n54328), .X(oi_15[5]) );
  inv_x2_sg U58817 ( .A(n54330), .X(oi_15[6]) );
  inv_x2_sg U58818 ( .A(n54332), .X(oi_15[7]) );
  inv_x2_sg U58819 ( .A(n54334), .X(oi_15[8]) );
  inv_x2_sg U58820 ( .A(n54336), .X(oi_15[9]) );
  inv_x2_sg U58821 ( .A(n54338), .X(oi_15[10]) );
  inv_x2_sg U58822 ( .A(n54340), .X(oi_15[11]) );
  inv_x2_sg U58823 ( .A(n54342), .X(oi_15[12]) );
  inv_x2_sg U58824 ( .A(n54344), .X(oi_15[13]) );
  inv_x2_sg U58825 ( .A(n54346), .X(oi_15[14]) );
  inv_x2_sg U58826 ( .A(n54348), .X(oi_15[15]) );
  inv_x2_sg U58827 ( .A(n54350), .X(oi_15[16]) );
  inv_x2_sg U58828 ( .A(n54352), .X(oi_15[17]) );
  inv_x2_sg U58829 ( .A(n54354), .X(oi_15[18]) );
  inv_x2_sg U58830 ( .A(n54356), .X(oi_15[19]) );
  inv_x2_sg U58831 ( .A(n54358), .X(oi_14[0]) );
  inv_x2_sg U58832 ( .A(n54360), .X(oi_14[1]) );
  inv_x2_sg U58833 ( .A(n54362), .X(oi_14[2]) );
  inv_x2_sg U58834 ( .A(n54364), .X(oi_14[3]) );
  inv_x2_sg U58835 ( .A(n54366), .X(oi_14[4]) );
  inv_x2_sg U58836 ( .A(n54368), .X(oi_14[5]) );
  inv_x2_sg U58837 ( .A(n54370), .X(oi_14[6]) );
  inv_x2_sg U58838 ( .A(n54372), .X(oi_14[7]) );
  inv_x2_sg U58839 ( .A(n54374), .X(oi_14[8]) );
  inv_x2_sg U58840 ( .A(n54376), .X(oi_14[9]) );
  inv_x2_sg U58841 ( .A(n54378), .X(oi_14[10]) );
  inv_x2_sg U58842 ( .A(n54380), .X(oi_14[11]) );
  inv_x2_sg U58843 ( .A(n54382), .X(oi_14[12]) );
  inv_x2_sg U58844 ( .A(n54384), .X(oi_14[13]) );
  inv_x2_sg U58845 ( .A(n54386), .X(oi_14[14]) );
  inv_x2_sg U58846 ( .A(n54388), .X(oi_14[15]) );
  inv_x2_sg U58847 ( .A(n54390), .X(oi_14[16]) );
  inv_x2_sg U58848 ( .A(n54392), .X(oi_14[17]) );
  inv_x2_sg U58849 ( .A(n54394), .X(oi_14[18]) );
  inv_x2_sg U58850 ( .A(n54396), .X(oi_14[19]) );
  inv_x2_sg U58851 ( .A(n54398), .X(oi_13[0]) );
  inv_x2_sg U58852 ( .A(n54400), .X(oi_13[1]) );
  inv_x2_sg U58853 ( .A(n54402), .X(oi_13[2]) );
  inv_x2_sg U58854 ( .A(n54404), .X(oi_13[3]) );
  inv_x2_sg U58855 ( .A(n54406), .X(oi_13[4]) );
  inv_x2_sg U58856 ( .A(n54408), .X(oi_13[5]) );
  inv_x2_sg U58857 ( .A(n54410), .X(oi_13[6]) );
  inv_x2_sg U58858 ( .A(n54412), .X(oi_13[7]) );
  inv_x2_sg U58859 ( .A(n54414), .X(oi_13[8]) );
  inv_x2_sg U58860 ( .A(n54416), .X(oi_13[9]) );
  inv_x2_sg U58861 ( .A(n54418), .X(oi_13[10]) );
  inv_x2_sg U58862 ( .A(n54420), .X(oi_13[11]) );
  inv_x2_sg U58863 ( .A(n54422), .X(oi_13[12]) );
  inv_x2_sg U58864 ( .A(n54424), .X(oi_13[13]) );
  inv_x2_sg U58865 ( .A(n54426), .X(oi_13[14]) );
  inv_x2_sg U58866 ( .A(n54428), .X(oi_13[15]) );
  inv_x2_sg U58867 ( .A(n54430), .X(oi_13[16]) );
  inv_x2_sg U58868 ( .A(n54432), .X(oi_13[17]) );
  inv_x2_sg U58869 ( .A(n54434), .X(oi_13[18]) );
  inv_x2_sg U58870 ( .A(n54436), .X(oi_13[19]) );
  inv_x2_sg U58871 ( .A(n54438), .X(oi_12[0]) );
  inv_x2_sg U58872 ( .A(n54440), .X(oi_12[1]) );
  inv_x2_sg U58873 ( .A(n54442), .X(oi_12[2]) );
  inv_x2_sg U58874 ( .A(n54444), .X(oi_12[3]) );
  inv_x2_sg U58875 ( .A(n54446), .X(oi_12[4]) );
  inv_x2_sg U58876 ( .A(n54448), .X(oi_12[5]) );
  inv_x2_sg U58877 ( .A(n54450), .X(oi_12[6]) );
  inv_x2_sg U58878 ( .A(n54452), .X(oi_12[7]) );
  inv_x2_sg U58879 ( .A(n54454), .X(oi_12[8]) );
  inv_x2_sg U58880 ( .A(n54456), .X(oi_12[9]) );
  inv_x2_sg U58881 ( .A(n54458), .X(oi_12[10]) );
  inv_x2_sg U58882 ( .A(n54460), .X(oi_12[11]) );
  inv_x2_sg U58883 ( .A(n54462), .X(oi_12[12]) );
  inv_x2_sg U58884 ( .A(n54464), .X(oi_12[13]) );
  inv_x2_sg U58885 ( .A(n54466), .X(oi_12[14]) );
  inv_x2_sg U58886 ( .A(n54468), .X(oi_12[15]) );
  inv_x2_sg U58887 ( .A(n54470), .X(oi_12[16]) );
  inv_x2_sg U58888 ( .A(n54472), .X(oi_12[17]) );
  inv_x2_sg U58889 ( .A(n54474), .X(oi_12[18]) );
  inv_x2_sg U58890 ( .A(n54476), .X(oi_12[19]) );
  inv_x2_sg U58891 ( .A(n54478), .X(oi_11[0]) );
  inv_x2_sg U58892 ( .A(n54480), .X(oi_11[1]) );
  inv_x2_sg U58893 ( .A(n54482), .X(oi_11[2]) );
  inv_x2_sg U58894 ( .A(n54484), .X(oi_11[3]) );
  inv_x2_sg U58895 ( .A(n54486), .X(oi_11[4]) );
  inv_x2_sg U58896 ( .A(n54488), .X(oi_11[5]) );
  inv_x2_sg U58897 ( .A(n54490), .X(oi_11[6]) );
  inv_x2_sg U58898 ( .A(n54492), .X(oi_11[7]) );
  inv_x2_sg U58899 ( .A(n54494), .X(oi_11[8]) );
  inv_x2_sg U58900 ( .A(n54496), .X(oi_11[9]) );
  inv_x2_sg U58901 ( .A(n54498), .X(oi_11[10]) );
  inv_x2_sg U58902 ( .A(n54500), .X(oi_11[11]) );
  inv_x2_sg U58903 ( .A(n54502), .X(oi_11[12]) );
  inv_x2_sg U58904 ( .A(n54504), .X(oi_11[13]) );
  inv_x2_sg U58905 ( .A(n54506), .X(oi_11[14]) );
  inv_x2_sg U58906 ( .A(n54508), .X(oi_11[15]) );
  inv_x2_sg U58907 ( .A(n54510), .X(oi_11[16]) );
  inv_x2_sg U58908 ( .A(n54512), .X(oi_11[17]) );
  inv_x2_sg U58909 ( .A(n54514), .X(oi_11[18]) );
  inv_x2_sg U58910 ( .A(n54516), .X(oi_11[19]) );
  inv_x2_sg U58911 ( .A(n54518), .X(oi_10[0]) );
  inv_x2_sg U58912 ( .A(n54520), .X(oi_10[1]) );
  inv_x2_sg U58913 ( .A(n54522), .X(oi_10[2]) );
  inv_x2_sg U58914 ( .A(n54524), .X(oi_10[3]) );
  inv_x2_sg U58915 ( .A(n54526), .X(oi_10[4]) );
  inv_x2_sg U58916 ( .A(n54528), .X(oi_10[5]) );
  inv_x2_sg U58917 ( .A(n54530), .X(oi_10[6]) );
  inv_x2_sg U58918 ( .A(n54532), .X(oi_10[7]) );
  inv_x2_sg U58919 ( .A(n54534), .X(oi_10[8]) );
  inv_x2_sg U58920 ( .A(n54536), .X(oi_10[9]) );
  inv_x2_sg U58921 ( .A(n54538), .X(oi_10[10]) );
  inv_x2_sg U58922 ( .A(n54540), .X(oi_10[11]) );
  inv_x2_sg U58923 ( .A(n54542), .X(oi_10[12]) );
  inv_x2_sg U58924 ( .A(n54544), .X(oi_10[13]) );
  inv_x2_sg U58925 ( .A(n54546), .X(oi_10[14]) );
  inv_x2_sg U58926 ( .A(n54548), .X(oi_10[15]) );
  inv_x2_sg U58927 ( .A(n54550), .X(oi_10[16]) );
  inv_x2_sg U58928 ( .A(n54552), .X(oi_10[17]) );
  inv_x2_sg U58929 ( .A(n54554), .X(oi_10[18]) );
  inv_x2_sg U58930 ( .A(n54556), .X(oi_10[19]) );
  inv_x2_sg U58931 ( .A(n54558), .X(oi_9[0]) );
  inv_x2_sg U58932 ( .A(n54560), .X(oi_9[1]) );
  inv_x2_sg U58933 ( .A(n54562), .X(oi_9[2]) );
  inv_x2_sg U58934 ( .A(n54564), .X(oi_9[3]) );
  inv_x2_sg U58935 ( .A(n54566), .X(oi_9[4]) );
  inv_x2_sg U58936 ( .A(n54568), .X(oi_9[5]) );
  inv_x2_sg U58937 ( .A(n54570), .X(oi_9[6]) );
  inv_x2_sg U58938 ( .A(n54572), .X(oi_9[7]) );
  inv_x2_sg U58939 ( .A(n54574), .X(oi_9[8]) );
  inv_x2_sg U58940 ( .A(n54576), .X(oi_9[9]) );
  inv_x2_sg U58941 ( .A(n54578), .X(oi_9[10]) );
  inv_x2_sg U58942 ( .A(n54580), .X(oi_9[11]) );
  inv_x2_sg U58943 ( .A(n54582), .X(oi_9[12]) );
  inv_x2_sg U58944 ( .A(n54584), .X(oi_9[13]) );
  inv_x2_sg U58945 ( .A(n54586), .X(oi_9[14]) );
  inv_x2_sg U58946 ( .A(n54588), .X(oi_9[15]) );
  inv_x2_sg U58947 ( .A(n54590), .X(oi_9[16]) );
  inv_x2_sg U58948 ( .A(n54592), .X(oi_9[17]) );
  inv_x2_sg U58949 ( .A(n54594), .X(oi_9[18]) );
  inv_x2_sg U58950 ( .A(n54596), .X(oi_9[19]) );
  inv_x2_sg U58951 ( .A(n54598), .X(oi_8[0]) );
  inv_x2_sg U58952 ( .A(n54600), .X(oi_8[1]) );
  inv_x2_sg U58953 ( .A(n54602), .X(oi_8[2]) );
  inv_x2_sg U58954 ( .A(n54604), .X(oi_8[3]) );
  inv_x2_sg U58955 ( .A(n54606), .X(oi_8[4]) );
  inv_x2_sg U58956 ( .A(n54608), .X(oi_8[5]) );
  inv_x2_sg U58957 ( .A(n54610), .X(oi_8[6]) );
  inv_x2_sg U58958 ( .A(n54612), .X(oi_8[7]) );
  inv_x2_sg U58959 ( .A(n54614), .X(oi_8[8]) );
  inv_x2_sg U58960 ( .A(n54616), .X(oi_8[9]) );
  inv_x2_sg U58961 ( .A(n54618), .X(oi_8[10]) );
  inv_x2_sg U58962 ( .A(n54620), .X(oi_8[11]) );
  inv_x2_sg U58963 ( .A(n54622), .X(oi_8[12]) );
  inv_x2_sg U58964 ( .A(n54624), .X(oi_8[13]) );
  inv_x2_sg U58965 ( .A(n54626), .X(oi_8[14]) );
  inv_x2_sg U58966 ( .A(n54628), .X(oi_8[15]) );
  inv_x2_sg U58967 ( .A(n54630), .X(oi_8[16]) );
  inv_x2_sg U58968 ( .A(n54632), .X(oi_8[17]) );
  inv_x2_sg U58969 ( .A(n54634), .X(oi_8[18]) );
  inv_x2_sg U58970 ( .A(n54636), .X(oi_8[19]) );
  inv_x2_sg U58971 ( .A(n54638), .X(oi_7[0]) );
  inv_x2_sg U58972 ( .A(n54640), .X(oi_7[1]) );
  inv_x2_sg U58973 ( .A(n54642), .X(oi_7[2]) );
  inv_x2_sg U58974 ( .A(n54644), .X(oi_7[3]) );
  inv_x2_sg U58975 ( .A(n54646), .X(oi_7[4]) );
  inv_x2_sg U58976 ( .A(n54648), .X(oi_7[5]) );
  inv_x2_sg U58977 ( .A(n54650), .X(oi_7[6]) );
  inv_x2_sg U58978 ( .A(n54652), .X(oi_7[7]) );
  inv_x2_sg U58979 ( .A(n54654), .X(oi_7[8]) );
  inv_x2_sg U58980 ( .A(n54656), .X(oi_7[9]) );
  inv_x2_sg U58981 ( .A(n54658), .X(oi_7[10]) );
  inv_x2_sg U58982 ( .A(n54660), .X(oi_7[11]) );
  inv_x2_sg U58983 ( .A(n54662), .X(oi_7[12]) );
  inv_x2_sg U58984 ( .A(n54664), .X(oi_7[13]) );
  inv_x2_sg U58985 ( .A(n54666), .X(oi_7[14]) );
  inv_x2_sg U58986 ( .A(n54668), .X(oi_7[15]) );
  inv_x2_sg U58987 ( .A(n54670), .X(oi_7[16]) );
  inv_x2_sg U58988 ( .A(n54672), .X(oi_7[17]) );
  inv_x2_sg U58989 ( .A(n54674), .X(oi_7[18]) );
  inv_x2_sg U58990 ( .A(n54676), .X(oi_7[19]) );
  inv_x2_sg U58991 ( .A(n54678), .X(oi_6[0]) );
  inv_x2_sg U58992 ( .A(n54680), .X(oi_6[1]) );
  inv_x2_sg U58993 ( .A(n54682), .X(oi_6[2]) );
  inv_x2_sg U58994 ( .A(n54684), .X(oi_6[3]) );
  inv_x2_sg U58995 ( .A(n54686), .X(oi_6[4]) );
  inv_x2_sg U58996 ( .A(n54688), .X(oi_6[5]) );
  inv_x2_sg U58997 ( .A(n54690), .X(oi_6[6]) );
  inv_x2_sg U58998 ( .A(n54692), .X(oi_6[7]) );
  inv_x2_sg U58999 ( .A(n54694), .X(oi_6[8]) );
  inv_x2_sg U59000 ( .A(n54696), .X(oi_6[9]) );
  inv_x2_sg U59001 ( .A(n54698), .X(oi_6[10]) );
  inv_x2_sg U59002 ( .A(n54700), .X(oi_6[11]) );
  inv_x2_sg U59003 ( .A(n54702), .X(oi_6[12]) );
  inv_x2_sg U59004 ( .A(n54704), .X(oi_6[13]) );
  inv_x2_sg U59005 ( .A(n54706), .X(oi_6[14]) );
  inv_x2_sg U59006 ( .A(n54708), .X(oi_6[15]) );
  inv_x2_sg U59007 ( .A(n54710), .X(oi_6[16]) );
  inv_x2_sg U59008 ( .A(n54712), .X(oi_6[17]) );
  inv_x2_sg U59009 ( .A(n54714), .X(oi_6[18]) );
  inv_x2_sg U59010 ( .A(n54716), .X(oi_6[19]) );
  inv_x2_sg U59011 ( .A(n54718), .X(oi_5[0]) );
  inv_x2_sg U59012 ( .A(n54720), .X(oi_5[1]) );
  inv_x2_sg U59013 ( .A(n54722), .X(oi_5[2]) );
  inv_x2_sg U59014 ( .A(n54724), .X(oi_5[3]) );
  inv_x2_sg U59015 ( .A(n54726), .X(oi_5[4]) );
  inv_x2_sg U59016 ( .A(n54728), .X(oi_5[5]) );
  inv_x2_sg U59017 ( .A(n54730), .X(oi_5[6]) );
  inv_x2_sg U59018 ( .A(n54732), .X(oi_5[7]) );
  inv_x2_sg U59019 ( .A(n54734), .X(oi_5[8]) );
  inv_x2_sg U59020 ( .A(n54736), .X(oi_5[9]) );
  inv_x2_sg U59021 ( .A(n54738), .X(oi_5[10]) );
  inv_x2_sg U59022 ( .A(n54740), .X(oi_5[11]) );
  inv_x2_sg U59023 ( .A(n54742), .X(oi_5[12]) );
  inv_x2_sg U59024 ( .A(n54744), .X(oi_5[13]) );
  inv_x2_sg U59025 ( .A(n54746), .X(oi_5[14]) );
  inv_x2_sg U59026 ( .A(n54748), .X(oi_5[15]) );
  inv_x2_sg U59027 ( .A(n54750), .X(oi_5[16]) );
  inv_x2_sg U59028 ( .A(n54752), .X(oi_5[17]) );
  inv_x2_sg U59029 ( .A(n54754), .X(oi_5[18]) );
  inv_x2_sg U59030 ( .A(n54756), .X(oi_5[19]) );
  inv_x2_sg U59031 ( .A(n54758), .X(oi_4[0]) );
  inv_x2_sg U59032 ( .A(n54760), .X(oi_4[1]) );
  inv_x2_sg U59033 ( .A(n54762), .X(oi_4[2]) );
  inv_x2_sg U59034 ( .A(n54764), .X(oi_4[3]) );
  inv_x2_sg U59035 ( .A(n54766), .X(oi_4[4]) );
  inv_x2_sg U59036 ( .A(n54768), .X(oi_4[5]) );
  inv_x2_sg U59037 ( .A(n54770), .X(oi_4[6]) );
  inv_x2_sg U59038 ( .A(n54772), .X(oi_4[7]) );
  inv_x2_sg U59039 ( .A(n54774), .X(oi_4[8]) );
  inv_x2_sg U59040 ( .A(n54776), .X(oi_4[9]) );
  inv_x2_sg U59041 ( .A(n54778), .X(oi_4[10]) );
  inv_x2_sg U59042 ( .A(n54780), .X(oi_4[11]) );
  inv_x2_sg U59043 ( .A(n54782), .X(oi_4[12]) );
  inv_x2_sg U59044 ( .A(n54784), .X(oi_4[13]) );
  inv_x2_sg U59045 ( .A(n54786), .X(oi_4[14]) );
  inv_x2_sg U59046 ( .A(n54788), .X(oi_4[15]) );
  inv_x2_sg U59047 ( .A(n54790), .X(oi_4[16]) );
  inv_x2_sg U59048 ( .A(n54792), .X(oi_4[17]) );
  inv_x2_sg U59049 ( .A(n54794), .X(oi_4[18]) );
  inv_x2_sg U59050 ( .A(n54796), .X(oi_4[19]) );
  inv_x2_sg U59051 ( .A(n54798), .X(oi_3[0]) );
  inv_x2_sg U59052 ( .A(n54800), .X(oi_3[1]) );
  inv_x2_sg U59053 ( .A(n54802), .X(oi_3[2]) );
  inv_x2_sg U59054 ( .A(n54804), .X(oi_3[3]) );
  inv_x2_sg U59055 ( .A(n54806), .X(oi_3[4]) );
  inv_x2_sg U59056 ( .A(n54808), .X(oi_3[5]) );
  inv_x2_sg U59057 ( .A(n54810), .X(oi_3[6]) );
  inv_x2_sg U59058 ( .A(n54812), .X(oi_3[7]) );
  inv_x2_sg U59059 ( .A(n54814), .X(oi_3[8]) );
  inv_x2_sg U59060 ( .A(n54816), .X(oi_3[9]) );
  inv_x2_sg U59061 ( .A(n54818), .X(oi_3[10]) );
  inv_x2_sg U59062 ( .A(n54820), .X(oi_3[11]) );
  inv_x2_sg U59063 ( .A(n54822), .X(oi_3[12]) );
  inv_x2_sg U59064 ( .A(n54824), .X(oi_3[13]) );
  inv_x2_sg U59065 ( .A(n54826), .X(oi_3[14]) );
  inv_x2_sg U59066 ( .A(n54828), .X(oi_3[15]) );
  inv_x2_sg U59067 ( .A(n54830), .X(oi_3[16]) );
  inv_x2_sg U59068 ( .A(n54832), .X(oi_3[17]) );
  inv_x2_sg U59069 ( .A(n54834), .X(oi_3[18]) );
  inv_x2_sg U59070 ( .A(n54836), .X(oi_3[19]) );
  inv_x2_sg U59071 ( .A(n54838), .X(oi_2[0]) );
  inv_x2_sg U59072 ( .A(n54840), .X(oi_2[1]) );
  inv_x2_sg U59073 ( .A(n54842), .X(oi_2[2]) );
  inv_x2_sg U59074 ( .A(n54844), .X(oi_2[3]) );
  inv_x2_sg U59075 ( .A(n54846), .X(oi_2[4]) );
  inv_x2_sg U59076 ( .A(n54848), .X(oi_2[5]) );
  inv_x2_sg U59077 ( .A(n54850), .X(oi_2[6]) );
  inv_x2_sg U59078 ( .A(n54852), .X(oi_2[7]) );
  inv_x2_sg U59079 ( .A(n54854), .X(oi_2[8]) );
  inv_x2_sg U59080 ( .A(n54856), .X(oi_2[9]) );
  inv_x2_sg U59081 ( .A(n54858), .X(oi_2[10]) );
  inv_x2_sg U59082 ( .A(n54860), .X(oi_2[11]) );
  inv_x2_sg U59083 ( .A(n54862), .X(oi_2[12]) );
  inv_x2_sg U59084 ( .A(n54864), .X(oi_2[13]) );
  inv_x2_sg U59085 ( .A(n54866), .X(oi_2[14]) );
  inv_x2_sg U59086 ( .A(n54868), .X(oi_2[15]) );
  inv_x2_sg U59087 ( .A(n54870), .X(oi_2[16]) );
  inv_x2_sg U59088 ( .A(n54872), .X(oi_2[17]) );
  inv_x2_sg U59089 ( .A(n54874), .X(oi_2[18]) );
  inv_x2_sg U59090 ( .A(n54876), .X(oi_2[19]) );
  inv_x2_sg U59091 ( .A(n54878), .X(oi_1[0]) );
  inv_x2_sg U59092 ( .A(n54880), .X(oi_1[1]) );
  inv_x2_sg U59093 ( .A(n54882), .X(oi_1[2]) );
  inv_x2_sg U59094 ( .A(n54884), .X(oi_1[3]) );
  inv_x2_sg U59095 ( .A(n54886), .X(oi_1[4]) );
  inv_x2_sg U59096 ( .A(n54888), .X(oi_1[5]) );
  inv_x2_sg U59097 ( .A(n54890), .X(oi_1[6]) );
  inv_x2_sg U59098 ( .A(n54892), .X(oi_1[7]) );
  inv_x2_sg U59099 ( .A(n54894), .X(oi_1[8]) );
  inv_x2_sg U59100 ( .A(n54896), .X(oi_1[9]) );
  inv_x2_sg U59101 ( .A(n54898), .X(oi_1[10]) );
  inv_x2_sg U59102 ( .A(n54900), .X(oi_1[11]) );
  inv_x2_sg U59103 ( .A(n54902), .X(oi_1[12]) );
  inv_x2_sg U59104 ( .A(n54904), .X(oi_1[13]) );
  inv_x2_sg U59105 ( .A(n54906), .X(oi_1[14]) );
  inv_x2_sg U59106 ( .A(n54908), .X(oi_1[15]) );
  inv_x2_sg U59107 ( .A(n54910), .X(oi_1[16]) );
  inv_x2_sg U59108 ( .A(n54912), .X(oi_1[17]) );
  inv_x2_sg U59109 ( .A(n54914), .X(oi_1[18]) );
  inv_x2_sg U59110 ( .A(n54916), .X(oi_1[19]) );
  inv_x2_sg U59111 ( .A(n54918), .X(oi_0[0]) );
  inv_x2_sg U59112 ( .A(n54920), .X(oi_0[1]) );
  inv_x2_sg U59113 ( .A(n54922), .X(oi_0[2]) );
  inv_x2_sg U59114 ( .A(n54924), .X(oi_0[3]) );
  inv_x2_sg U59115 ( .A(n54926), .X(oi_0[4]) );
  inv_x2_sg U59116 ( .A(n54928), .X(oi_0[5]) );
  inv_x2_sg U59117 ( .A(n54930), .X(oi_0[6]) );
  inv_x2_sg U59118 ( .A(n54932), .X(oi_0[7]) );
  inv_x2_sg U59119 ( .A(n54934), .X(oi_0[8]) );
  inv_x2_sg U59120 ( .A(n54936), .X(oi_0[9]) );
  inv_x2_sg U59121 ( .A(n54938), .X(oi_0[10]) );
  inv_x2_sg U59122 ( .A(n54940), .X(oi_0[11]) );
  inv_x2_sg U59123 ( .A(n54942), .X(oi_0[12]) );
  inv_x2_sg U59124 ( .A(n54944), .X(oi_0[13]) );
  inv_x2_sg U59125 ( .A(n54946), .X(oi_0[14]) );
  inv_x2_sg U59126 ( .A(n54948), .X(oi_0[15]) );
  inv_x2_sg U59127 ( .A(n54950), .X(oi_0[16]) );
  inv_x2_sg U59128 ( .A(n54952), .X(oi_0[17]) );
  inv_x2_sg U59129 ( .A(n54954), .X(oi_0[18]) );
  inv_x2_sg U59130 ( .A(n54956), .X(oi_0[19]) );
  inv_x2_sg U59131 ( .A(n54958), .X(ow_15[1]) );
  inv_x2_sg U59132 ( .A(n54960), .X(ow_15[2]) );
  inv_x2_sg U59133 ( .A(n54962), .X(ow_15[3]) );
  inv_x2_sg U59134 ( .A(n54964), .X(ow_15[4]) );
  inv_x2_sg U59135 ( .A(n54966), .X(ow_15[5]) );
  inv_x2_sg U59136 ( .A(n54968), .X(ow_15[6]) );
  inv_x2_sg U59137 ( .A(n54970), .X(ow_15[7]) );
  inv_x2_sg U59138 ( .A(n54972), .X(ow_15[8]) );
  inv_x2_sg U59139 ( .A(n54974), .X(ow_15[9]) );
  inv_x2_sg U59140 ( .A(n54976), .X(ow_15[10]) );
  inv_x2_sg U59141 ( .A(n54978), .X(ow_15[11]) );
  inv_x2_sg U59142 ( .A(n54980), .X(ow_15[12]) );
  inv_x2_sg U59143 ( .A(n54982), .X(ow_15[13]) );
  inv_x2_sg U59144 ( .A(n54984), .X(ow_15[14]) );
  inv_x2_sg U59145 ( .A(n54986), .X(ow_15[15]) );
  inv_x2_sg U59146 ( .A(n54988), .X(ow_15[16]) );
  inv_x2_sg U59147 ( .A(n54990), .X(ow_15[17]) );
  inv_x2_sg U59148 ( .A(n54992), .X(ow_15[18]) );
  inv_x2_sg U59149 ( .A(n54994), .X(ow_15[19]) );
  inv_x2_sg U59150 ( .A(n54996), .X(ow_15[0]) );
  inv_x4_sg U59151 ( .A(n54998), .X(n54999) );
  inv_x4_sg U59152 ( .A(n55000), .X(n55001) );
  inv_x4_sg U59153 ( .A(n55002), .X(n55003) );
  inv_x4_sg U59154 ( .A(n55004), .X(n55005) );
  inv_x4_sg U59155 ( .A(n55006), .X(n55007) );
  inv_x4_sg U59156 ( .A(n55008), .X(n55009) );
  inv_x4_sg U59157 ( .A(n55010), .X(n55011) );
  inv_x4_sg U59158 ( .A(n55012), .X(n55013) );
  inv_x4_sg U59159 ( .A(n55014), .X(n55015) );
  inv_x4_sg U59160 ( .A(n55016), .X(n55017) );
  inv_x4_sg U59161 ( .A(n55018), .X(n55019) );
  inv_x4_sg U59162 ( .A(n55020), .X(n55021) );
  inv_x4_sg U59163 ( .A(n55022), .X(n55023) );
  inv_x4_sg U59164 ( .A(n55024), .X(n55025) );
  inv_x4_sg U59165 ( .A(n55026), .X(n55027) );
  inv_x4_sg U59166 ( .A(n55028), .X(n55029) );
  inv_x4_sg U59167 ( .A(n55030), .X(n55031) );
  inv_x4_sg U59168 ( .A(n55032), .X(n55033) );
  inv_x4_sg U59169 ( .A(n55034), .X(n55035) );
  inv_x4_sg U59170 ( .A(n55036), .X(n55037) );
  inv_x4_sg U59171 ( .A(n55038), .X(n55039) );
  inv_x4_sg U59172 ( .A(n55040), .X(n55041) );
  inv_x4_sg U59173 ( .A(n55042), .X(n55043) );
  inv_x4_sg U59174 ( .A(n55044), .X(n55045) );
  inv_x4_sg U59175 ( .A(n55046), .X(n55047) );
  inv_x4_sg U59176 ( .A(n55048), .X(n55049) );
  inv_x4_sg U59177 ( .A(n55050), .X(n55051) );
  inv_x4_sg U59178 ( .A(n55052), .X(n55053) );
  inv_x4_sg U59179 ( .A(n55054), .X(n55055) );
  inv_x4_sg U59180 ( .A(n55056), .X(n55057) );
  inv_x4_sg U59181 ( .A(n55058), .X(n55059) );
  inv_x4_sg U59182 ( .A(n55060), .X(n55061) );
  inv_x4_sg U59183 ( .A(n55062), .X(n55063) );
  inv_x4_sg U59184 ( .A(n55064), .X(n55065) );
  inv_x4_sg U59185 ( .A(n55066), .X(n55067) );
  inv_x4_sg U59186 ( .A(n55068), .X(n55069) );
  inv_x4_sg U59187 ( .A(n55070), .X(n55071) );
  nand_x4_sg U59188 ( .A(n39705), .B(n55071), .X(n35839) );
  nor_x2_sg U59189 ( .A(n68389), .B(n57303), .X(n32799) );
  nor_x8_sg U59190 ( .A(n67535), .B(n57307), .X(n26113) );
  nor_x4_sg U59191 ( .A(n31962), .B(n32090), .X(n31979) );
  nand_x4_sg U59192 ( .A(n32091), .B(n32092), .X(n32090) );
  inv_x4_sg U59193 ( .A(n55072), .X(n55073) );
  inv_x4_sg U59194 ( .A(n55074), .X(n55075) );
  inv_x4_sg U59195 ( .A(n55076), .X(n55077) );
  inv_x4_sg U59196 ( .A(n55078), .X(n55079) );
  inv_x4_sg U59197 ( .A(n55080), .X(n55081) );
  inv_x4_sg U59198 ( .A(n55082), .X(n55083) );
  inv_x4_sg U59199 ( .A(n55084), .X(n55085) );
  inv_x4_sg U59200 ( .A(n55086), .X(n55087) );
  inv_x4_sg U59201 ( .A(n55088), .X(n55089) );
  inv_x4_sg U59202 ( .A(n55090), .X(n55091) );
  inv_x4_sg U59203 ( .A(n55092), .X(n55093) );
  inv_x4_sg U59204 ( .A(n55094), .X(n55095) );
  inv_x4_sg U59205 ( .A(n55096), .X(n55097) );
  inv_x4_sg U59206 ( .A(n55098), .X(n55099) );
  inv_x4_sg U59207 ( .A(n55100), .X(n55101) );
  inv_x4_sg U59208 ( .A(n55102), .X(n55103) );
  inv_x4_sg U59209 ( .A(n55104), .X(n55105) );
  inv_x4_sg U59210 ( .A(n55106), .X(n55107) );
  inv_x4_sg U59211 ( .A(n55108), .X(n55109) );
  inv_x4_sg U59212 ( .A(n55110), .X(n55111) );
  inv_x4_sg U59213 ( .A(n55112), .X(n55113) );
  inv_x4_sg U59214 ( .A(n55114), .X(n55115) );
  inv_x4_sg U59215 ( .A(n55116), .X(n55117) );
  inv_x4_sg U59216 ( .A(n55118), .X(n55119) );
  inv_x4_sg U59217 ( .A(n55120), .X(n55121) );
  inv_x4_sg U59218 ( .A(n55122), .X(n55123) );
  inv_x4_sg U59219 ( .A(n55124), .X(n55125) );
  inv_x4_sg U59220 ( .A(n55126), .X(n55127) );
  inv_x4_sg U59221 ( .A(n55128), .X(n55129) );
  inv_x4_sg U59222 ( .A(n55130), .X(n55131) );
  inv_x4_sg U59223 ( .A(n55132), .X(n55133) );
  inv_x4_sg U59224 ( .A(n55134), .X(n55135) );
  inv_x4_sg U59225 ( .A(n55136), .X(n55137) );
  inv_x4_sg U59226 ( .A(n55138), .X(n55139) );
  inv_x4_sg U59227 ( .A(n55140), .X(n55141) );
  inv_x4_sg U59228 ( .A(n55142), .X(n55143) );
  inv_x4_sg U59229 ( .A(n55144), .X(n55145) );
  inv_x4_sg U59230 ( .A(n55146), .X(n55147) );
  inv_x4_sg U59231 ( .A(n55148), .X(n55149) );
  inv_x4_sg U59232 ( .A(n55150), .X(n55151) );
  inv_x4_sg U59233 ( .A(n55152), .X(n55153) );
  inv_x4_sg U59234 ( .A(n55154), .X(n55155) );
  inv_x4_sg U59235 ( .A(n55156), .X(n55157) );
  inv_x4_sg U59236 ( .A(n55158), .X(n55159) );
  inv_x4_sg U59237 ( .A(n55160), .X(n55161) );
  inv_x4_sg U59238 ( .A(n55162), .X(n55163) );
  inv_x4_sg U59239 ( .A(n55164), .X(n55165) );
  inv_x4_sg U59240 ( .A(n55166), .X(n55167) );
  inv_x4_sg U59241 ( .A(n55168), .X(n55169) );
  inv_x4_sg U59242 ( .A(n55170), .X(n55171) );
  inv_x4_sg U59243 ( .A(n55172), .X(n55173) );
  inv_x4_sg U59244 ( .A(n55174), .X(n55175) );
  inv_x4_sg U59245 ( .A(n55176), .X(n55177) );
  inv_x4_sg U59246 ( .A(n55178), .X(n55179) );
  inv_x4_sg U59247 ( .A(n55180), .X(n55181) );
  inv_x4_sg U59248 ( .A(n55182), .X(n55183) );
  inv_x4_sg U59249 ( .A(n55184), .X(n55185) );
  inv_x4_sg U59250 ( .A(n55186), .X(n55187) );
  inv_x4_sg U59251 ( .A(n55188), .X(n55189) );
  inv_x4_sg U59252 ( .A(n55190), .X(n55191) );
  inv_x4_sg U59253 ( .A(n55192), .X(n55193) );
  inv_x4_sg U59254 ( .A(n55194), .X(n55195) );
  inv_x4_sg U59255 ( .A(n55196), .X(n55197) );
  inv_x4_sg U59256 ( .A(n55198), .X(n55199) );
  inv_x4_sg U59257 ( .A(n55200), .X(n55201) );
  inv_x4_sg U59258 ( .A(n55202), .X(n55203) );
  inv_x4_sg U59259 ( .A(n55204), .X(n55205) );
  inv_x4_sg U59260 ( .A(n55206), .X(n55207) );
  inv_x4_sg U59261 ( .A(n55208), .X(n55209) );
  inv_x4_sg U59262 ( .A(n55210), .X(n55211) );
  inv_x4_sg U59263 ( .A(n55212), .X(n55213) );
  inv_x4_sg U59264 ( .A(n55214), .X(n55215) );
  inv_x4_sg U59265 ( .A(n55216), .X(n55217) );
  inv_x4_sg U59266 ( .A(n55218), .X(n55219) );
  inv_x4_sg U59267 ( .A(n55220), .X(n55221) );
  inv_x4_sg U59268 ( .A(n55222), .X(n55223) );
  inv_x4_sg U59269 ( .A(n55224), .X(n55225) );
  inv_x4_sg U59270 ( .A(n55226), .X(n55227) );
  inv_x4_sg U59271 ( .A(n55228), .X(n55229) );
  inv_x4_sg U59272 ( .A(n55230), .X(n55231) );
  inv_x4_sg U59273 ( .A(n55232), .X(n55233) );
  inv_x4_sg U59274 ( .A(n55234), .X(n55235) );
  inv_x4_sg U59275 ( .A(n55236), .X(n55237) );
  inv_x4_sg U59276 ( .A(n55238), .X(n55239) );
  inv_x4_sg U59277 ( .A(n55240), .X(n55241) );
  inv_x4_sg U59278 ( .A(n55242), .X(n55243) );
  inv_x4_sg U59279 ( .A(n55244), .X(n55245) );
  inv_x4_sg U59280 ( .A(n55246), .X(n55247) );
  inv_x4_sg U59281 ( .A(n55248), .X(n55249) );
  inv_x4_sg U59282 ( .A(n55250), .X(n55251) );
  inv_x4_sg U59283 ( .A(n55252), .X(n55253) );
  inv_x4_sg U59284 ( .A(n55254), .X(n55255) );
  inv_x4_sg U59285 ( .A(n55256), .X(n55257) );
  inv_x4_sg U59286 ( .A(n55258), .X(n55259) );
  inv_x4_sg U59287 ( .A(n55260), .X(n55261) );
  inv_x4_sg U59288 ( .A(n55262), .X(n55263) );
  inv_x4_sg U59289 ( .A(n55264), .X(n55265) );
  inv_x4_sg U59290 ( .A(n55266), .X(n55267) );
  inv_x4_sg U59291 ( .A(n55268), .X(n55269) );
  inv_x4_sg U59292 ( .A(n55270), .X(n55271) );
  inv_x4_sg U59293 ( .A(n55272), .X(n55273) );
  inv_x4_sg U59294 ( .A(n55274), .X(n55275) );
  inv_x4_sg U59295 ( .A(n55276), .X(n55277) );
  inv_x4_sg U59296 ( .A(n55278), .X(n55279) );
  inv_x4_sg U59297 ( .A(n55280), .X(n55281) );
  inv_x4_sg U59298 ( .A(n55282), .X(n55283) );
  inv_x4_sg U59299 ( .A(n55284), .X(n55285) );
  inv_x4_sg U59300 ( .A(n55286), .X(n55287) );
  inv_x4_sg U59301 ( .A(n55288), .X(n55289) );
  inv_x4_sg U59302 ( .A(n55290), .X(n55291) );
  inv_x4_sg U59303 ( .A(n55292), .X(n55293) );
  inv_x4_sg U59304 ( .A(n55294), .X(n55295) );
  inv_x4_sg U59305 ( .A(n55296), .X(n55297) );
  inv_x4_sg U59306 ( .A(n55298), .X(n55299) );
  inv_x4_sg U59307 ( .A(n55300), .X(n55301) );
  inv_x4_sg U59308 ( .A(n55302), .X(n55303) );
  inv_x4_sg U59309 ( .A(n55304), .X(n55305) );
  inv_x4_sg U59310 ( .A(n55306), .X(n55307) );
  inv_x4_sg U59311 ( .A(n55308), .X(n55309) );
  inv_x4_sg U59312 ( .A(n55310), .X(n55311) );
  inv_x4_sg U59313 ( .A(n55312), .X(n55313) );
  inv_x4_sg U59314 ( .A(n55314), .X(n55315) );
  inv_x4_sg U59315 ( .A(n55316), .X(n55317) );
  inv_x4_sg U59316 ( .A(n55318), .X(n55319) );
  inv_x4_sg U59317 ( .A(n55320), .X(n55321) );
  inv_x4_sg U59318 ( .A(n55322), .X(n55323) );
  inv_x4_sg U59319 ( .A(n55324), .X(n55325) );
  inv_x4_sg U59320 ( .A(n55326), .X(n55327) );
  inv_x4_sg U59321 ( .A(n55328), .X(n55329) );
  inv_x4_sg U59322 ( .A(n55330), .X(n55331) );
  inv_x4_sg U59323 ( .A(n55332), .X(n55333) );
  inv_x4_sg U59324 ( .A(n55334), .X(n55335) );
  inv_x4_sg U59325 ( .A(n55336), .X(n55337) );
  inv_x4_sg U59326 ( .A(n55338), .X(n55339) );
  inv_x4_sg U59327 ( .A(n55340), .X(n55341) );
  inv_x4_sg U59328 ( .A(n55342), .X(n55343) );
  inv_x4_sg U59329 ( .A(n55344), .X(n55345) );
  inv_x4_sg U59330 ( .A(n55346), .X(n55347) );
  inv_x4_sg U59331 ( .A(n55348), .X(n55349) );
  inv_x4_sg U59332 ( .A(n55350), .X(n55351) );
  inv_x4_sg U59333 ( .A(n55352), .X(n55353) );
  inv_x4_sg U59334 ( .A(n55354), .X(n55355) );
  inv_x4_sg U59335 ( .A(n55356), .X(n55357) );
  inv_x4_sg U59336 ( .A(n55358), .X(n55359) );
  inv_x4_sg U59337 ( .A(n55360), .X(n55361) );
  inv_x4_sg U59338 ( .A(n55362), .X(n55363) );
  inv_x4_sg U59339 ( .A(n55364), .X(n55365) );
  inv_x4_sg U59340 ( .A(n55366), .X(n55367) );
  inv_x4_sg U59341 ( .A(n55368), .X(n55369) );
  inv_x4_sg U59342 ( .A(n55370), .X(n55371) );
  inv_x4_sg U59343 ( .A(n55372), .X(n55373) );
  inv_x4_sg U59344 ( .A(n55374), .X(n55375) );
  inv_x4_sg U59345 ( .A(n55376), .X(n55377) );
  inv_x4_sg U59346 ( .A(n55378), .X(n55379) );
  inv_x4_sg U59347 ( .A(n55380), .X(n55381) );
  inv_x4_sg U59348 ( .A(n55382), .X(n55383) );
  inv_x4_sg U59349 ( .A(n55384), .X(n55385) );
  inv_x4_sg U59350 ( .A(n55386), .X(n55387) );
  inv_x4_sg U59351 ( .A(n55388), .X(n55389) );
  inv_x4_sg U59352 ( .A(n55390), .X(n55391) );
  inv_x4_sg U59353 ( .A(n55392), .X(n55393) );
  inv_x4_sg U59354 ( .A(n55394), .X(n55395) );
  inv_x4_sg U59355 ( .A(n55396), .X(n55397) );
  inv_x4_sg U59356 ( .A(n55398), .X(n55399) );
  inv_x4_sg U59357 ( .A(n55400), .X(n55401) );
  inv_x4_sg U59358 ( .A(n55402), .X(n55403) );
  inv_x4_sg U59359 ( .A(n55404), .X(n55405) );
  inv_x4_sg U59360 ( .A(n55406), .X(n55407) );
  inv_x4_sg U59361 ( .A(n55408), .X(n55409) );
  inv_x4_sg U59362 ( .A(n55410), .X(n55411) );
  inv_x4_sg U59363 ( .A(n55412), .X(n55413) );
  inv_x4_sg U59364 ( .A(n55414), .X(n55415) );
  inv_x4_sg U59365 ( .A(n55416), .X(n55417) );
  inv_x4_sg U59366 ( .A(n55418), .X(n55419) );
  inv_x4_sg U59367 ( .A(n55420), .X(n55421) );
  inv_x4_sg U59368 ( .A(n55422), .X(n55423) );
  inv_x4_sg U59369 ( .A(n55424), .X(n55425) );
  inv_x4_sg U59370 ( .A(n55426), .X(n55427) );
  inv_x4_sg U59371 ( .A(n55428), .X(n55429) );
  inv_x4_sg U59372 ( .A(n55430), .X(n55431) );
  inv_x4_sg U59373 ( .A(n55432), .X(n55433) );
  inv_x4_sg U59374 ( .A(n55434), .X(n55435) );
  inv_x4_sg U59375 ( .A(n55436), .X(n55437) );
  inv_x4_sg U59376 ( .A(n55438), .X(n55439) );
  inv_x4_sg U59377 ( .A(n55440), .X(n55441) );
  inv_x4_sg U59378 ( .A(n55442), .X(n55443) );
  inv_x4_sg U59379 ( .A(n55444), .X(n55445) );
  inv_x4_sg U59380 ( .A(n55446), .X(n55447) );
  inv_x4_sg U59381 ( .A(n55448), .X(n55449) );
  inv_x4_sg U59382 ( .A(n55450), .X(n55451) );
  inv_x4_sg U59383 ( .A(n55452), .X(n55453) );
  inv_x4_sg U59384 ( .A(n55454), .X(n55455) );
  inv_x4_sg U59385 ( .A(n55456), .X(n55457) );
  inv_x4_sg U59386 ( .A(n55458), .X(n55459) );
  inv_x4_sg U59387 ( .A(n55460), .X(n55461) );
  inv_x4_sg U59388 ( .A(n55462), .X(n55463) );
  inv_x4_sg U59389 ( .A(n55464), .X(n55465) );
  inv_x4_sg U59390 ( .A(n55466), .X(n55467) );
  inv_x4_sg U59391 ( .A(n55468), .X(n55469) );
  inv_x4_sg U59392 ( .A(n55470), .X(n55471) );
  inv_x4_sg U59393 ( .A(n55472), .X(n55473) );
  inv_x4_sg U59394 ( .A(n55474), .X(n55475) );
  inv_x4_sg U59395 ( .A(n55476), .X(n55477) );
  inv_x4_sg U59396 ( .A(n55478), .X(n55479) );
  inv_x4_sg U59397 ( .A(n55480), .X(n55481) );
  inv_x4_sg U59398 ( .A(n55482), .X(n55483) );
  inv_x4_sg U59399 ( .A(n55484), .X(n55485) );
  inv_x4_sg U59400 ( .A(n55486), .X(n55487) );
  inv_x4_sg U59401 ( .A(n55488), .X(n55489) );
  inv_x4_sg U59402 ( .A(n55490), .X(n55491) );
  inv_x4_sg U59403 ( .A(n55492), .X(n55493) );
  inv_x4_sg U59404 ( .A(n55494), .X(n55495) );
  inv_x4_sg U59405 ( .A(n55496), .X(n55497) );
  inv_x4_sg U59406 ( .A(n55498), .X(n55499) );
  inv_x4_sg U59407 ( .A(n55500), .X(n55501) );
  inv_x4_sg U59408 ( .A(n55502), .X(n55503) );
  inv_x4_sg U59409 ( .A(n55504), .X(n55505) );
  inv_x4_sg U59410 ( .A(n55506), .X(n55507) );
  inv_x4_sg U59411 ( .A(n55508), .X(n55509) );
  inv_x4_sg U59412 ( .A(n55510), .X(n55511) );
  inv_x4_sg U59413 ( .A(n55512), .X(n55513) );
  inv_x4_sg U59414 ( .A(n55514), .X(n55515) );
  inv_x4_sg U59415 ( .A(n55516), .X(n55517) );
  inv_x4_sg U59416 ( .A(n55518), .X(n55519) );
  inv_x4_sg U59417 ( .A(n55520), .X(n55521) );
  inv_x4_sg U59418 ( .A(n55522), .X(n55523) );
  inv_x4_sg U59419 ( .A(n55524), .X(n55525) );
  inv_x4_sg U59420 ( .A(n55526), .X(n55527) );
  inv_x4_sg U59421 ( .A(n55528), .X(n55529) );
  inv_x4_sg U59422 ( .A(n55530), .X(n55531) );
  inv_x4_sg U59423 ( .A(n55532), .X(n55533) );
  inv_x4_sg U59424 ( .A(n55534), .X(n55535) );
  inv_x4_sg U59425 ( .A(n55536), .X(n55537) );
  inv_x4_sg U59426 ( .A(n55538), .X(n55539) );
  inv_x4_sg U59427 ( .A(n55540), .X(n55541) );
  inv_x4_sg U59428 ( .A(n55542), .X(n55543) );
  inv_x4_sg U59429 ( .A(n55544), .X(n55545) );
  inv_x4_sg U59430 ( .A(n55546), .X(n55547) );
  inv_x4_sg U59431 ( .A(n55548), .X(n55549) );
  inv_x4_sg U59432 ( .A(n55550), .X(n55551) );
  inv_x4_sg U59433 ( .A(n55552), .X(n55553) );
  inv_x4_sg U59434 ( .A(n55554), .X(n55555) );
  inv_x4_sg U59435 ( .A(n55556), .X(n55557) );
  inv_x4_sg U59436 ( .A(n55558), .X(n55559) );
  inv_x4_sg U59437 ( .A(n55560), .X(n55561) );
  inv_x4_sg U59438 ( .A(n55562), .X(n55563) );
  inv_x4_sg U59439 ( .A(n55564), .X(n55565) );
  inv_x4_sg U59440 ( .A(n55566), .X(n55567) );
  inv_x4_sg U59441 ( .A(n55568), .X(n55569) );
  inv_x4_sg U59442 ( .A(n55570), .X(n55571) );
  inv_x4_sg U59443 ( .A(n55572), .X(n55573) );
  inv_x4_sg U59444 ( .A(n55574), .X(n55575) );
  inv_x4_sg U59445 ( .A(n55576), .X(n55577) );
  inv_x4_sg U59446 ( .A(n55578), .X(n55579) );
  inv_x4_sg U59447 ( .A(n55580), .X(n55581) );
  inv_x4_sg U59448 ( .A(n55582), .X(n55583) );
  inv_x4_sg U59449 ( .A(n55584), .X(n55585) );
  inv_x4_sg U59450 ( .A(n55586), .X(n55587) );
  inv_x4_sg U59451 ( .A(n55588), .X(n55589) );
  inv_x4_sg U59452 ( .A(n55590), .X(n55591) );
  inv_x4_sg U59453 ( .A(n55592), .X(n55593) );
  inv_x4_sg U59454 ( .A(n55594), .X(n55595) );
  inv_x4_sg U59455 ( .A(n55596), .X(n55597) );
  inv_x4_sg U59456 ( .A(n55598), .X(n55599) );
  inv_x4_sg U59457 ( .A(n55600), .X(n55601) );
  inv_x4_sg U59458 ( .A(n55602), .X(n55603) );
  inv_x4_sg U59459 ( .A(n55604), .X(n55605) );
  inv_x4_sg U59460 ( .A(n55606), .X(n55607) );
  inv_x4_sg U59461 ( .A(n55608), .X(n55609) );
  inv_x4_sg U59462 ( .A(n55610), .X(n55611) );
  inv_x4_sg U59463 ( .A(n55612), .X(n55613) );
  inv_x4_sg U59464 ( .A(n55614), .X(n55615) );
  inv_x4_sg U59465 ( .A(n55616), .X(n55617) );
  inv_x4_sg U59466 ( .A(n55618), .X(n55619) );
  inv_x4_sg U59467 ( .A(n55620), .X(n55621) );
  inv_x4_sg U59468 ( .A(n55622), .X(n55623) );
  inv_x4_sg U59469 ( .A(n55624), .X(n55625) );
  inv_x4_sg U59470 ( .A(n55626), .X(n55627) );
  inv_x4_sg U59471 ( .A(n55628), .X(n55629) );
  inv_x4_sg U59472 ( .A(n55630), .X(n55631) );
  inv_x4_sg U59473 ( .A(n55632), .X(n55633) );
  inv_x4_sg U59474 ( .A(n55634), .X(n55635) );
  inv_x4_sg U59475 ( .A(n55636), .X(n55637) );
  inv_x4_sg U59476 ( .A(n55638), .X(n55639) );
  inv_x4_sg U59477 ( .A(n55640), .X(n55641) );
  inv_x4_sg U59478 ( .A(n55642), .X(n55643) );
  inv_x4_sg U59479 ( .A(n55644), .X(n55645) );
  inv_x4_sg U59480 ( .A(n55646), .X(n55647) );
  inv_x4_sg U59481 ( .A(n55648), .X(n55649) );
  inv_x4_sg U59482 ( .A(n55650), .X(n55651) );
  inv_x4_sg U59483 ( .A(n55652), .X(n55653) );
  inv_x4_sg U59484 ( .A(n55654), .X(n55655) );
  inv_x4_sg U59485 ( .A(n55656), .X(n55657) );
  inv_x4_sg U59486 ( .A(n55658), .X(n55659) );
  inv_x4_sg U59487 ( .A(n55660), .X(n55661) );
  inv_x4_sg U59488 ( .A(n55662), .X(n55663) );
  inv_x4_sg U59489 ( .A(n55664), .X(n55665) );
  inv_x4_sg U59490 ( .A(n55666), .X(n55667) );
  inv_x4_sg U59491 ( .A(n55668), .X(n55669) );
  inv_x4_sg U59492 ( .A(n55670), .X(n55671) );
  inv_x4_sg U59493 ( .A(n55672), .X(n55673) );
  inv_x4_sg U59494 ( .A(n55674), .X(n55675) );
  inv_x4_sg U59495 ( .A(n55676), .X(n55677) );
  inv_x4_sg U59496 ( .A(n55678), .X(n55679) );
  inv_x4_sg U59497 ( .A(n55680), .X(n55681) );
  inv_x4_sg U59498 ( .A(n55682), .X(n55683) );
  inv_x4_sg U59499 ( .A(n55684), .X(n55685) );
  inv_x4_sg U59500 ( .A(n55686), .X(n55687) );
  inv_x4_sg U59501 ( .A(n55688), .X(n55689) );
  inv_x4_sg U59502 ( .A(n55690), .X(n55691) );
  inv_x4_sg U59503 ( .A(n55692), .X(n55693) );
  inv_x4_sg U59504 ( .A(n55694), .X(n55695) );
  inv_x4_sg U59505 ( .A(n55696), .X(n55697) );
  inv_x4_sg U59506 ( .A(n55698), .X(n55699) );
  inv_x4_sg U59507 ( .A(n55700), .X(n55701) );
  inv_x4_sg U59508 ( .A(n55702), .X(n55703) );
  inv_x4_sg U59509 ( .A(n55704), .X(n55705) );
  inv_x4_sg U59510 ( .A(n55706), .X(n55707) );
  inv_x4_sg U59511 ( .A(n55708), .X(n55709) );
  inv_x4_sg U59512 ( .A(n55710), .X(n55711) );
  inv_x4_sg U59513 ( .A(n55712), .X(n55713) );
  inv_x4_sg U59514 ( .A(n55714), .X(n55715) );
  inv_x4_sg U59515 ( .A(n55716), .X(n55717) );
  inv_x4_sg U59516 ( .A(n55718), .X(n55719) );
  inv_x4_sg U59517 ( .A(n55720), .X(n55721) );
  inv_x4_sg U59518 ( .A(n55722), .X(n55723) );
  inv_x4_sg U59519 ( .A(n55724), .X(n55725) );
  inv_x4_sg U59520 ( .A(n55726), .X(n55727) );
  inv_x4_sg U59521 ( .A(n55728), .X(n55729) );
  inv_x4_sg U59522 ( .A(n55730), .X(n55731) );
  inv_x4_sg U59523 ( .A(n55732), .X(n55733) );
  inv_x4_sg U59524 ( .A(n55734), .X(n55735) );
  inv_x4_sg U59525 ( .A(n55736), .X(n55737) );
  inv_x4_sg U59526 ( .A(n55738), .X(n55739) );
  inv_x4_sg U59527 ( .A(n55740), .X(n55741) );
  inv_x4_sg U59528 ( .A(n55742), .X(n55743) );
  inv_x4_sg U59529 ( .A(n55744), .X(n55745) );
  inv_x4_sg U59530 ( .A(n55746), .X(n55747) );
  inv_x4_sg U59531 ( .A(n55748), .X(n55749) );
  inv_x4_sg U59532 ( .A(n55750), .X(n55751) );
  inv_x4_sg U59533 ( .A(n55752), .X(n55753) );
  inv_x4_sg U59534 ( .A(n55754), .X(n55755) );
  inv_x4_sg U59535 ( .A(n55756), .X(n55757) );
  inv_x4_sg U59536 ( .A(n55758), .X(n55759) );
  inv_x4_sg U59537 ( .A(n55760), .X(n55761) );
  inv_x4_sg U59538 ( .A(n55762), .X(n55763) );
  inv_x4_sg U59539 ( .A(n55764), .X(n55765) );
  inv_x4_sg U59540 ( .A(n55766), .X(n55767) );
  inv_x4_sg U59541 ( .A(n55768), .X(n55769) );
  inv_x4_sg U59542 ( .A(n55770), .X(n55771) );
  inv_x4_sg U59543 ( .A(n55772), .X(n55773) );
  inv_x4_sg U59544 ( .A(n55774), .X(n55775) );
  inv_x4_sg U59545 ( .A(n55776), .X(n55777) );
  inv_x4_sg U59546 ( .A(n55778), .X(n55779) );
  inv_x4_sg U59547 ( .A(n55780), .X(n55781) );
  inv_x4_sg U59548 ( .A(n55782), .X(n55783) );
  inv_x4_sg U59549 ( .A(n55784), .X(n55785) );
  inv_x4_sg U59550 ( .A(n55786), .X(n55787) );
  inv_x4_sg U59551 ( .A(n55788), .X(n55789) );
  inv_x4_sg U59552 ( .A(n55790), .X(n55791) );
  inv_x4_sg U59553 ( .A(n55792), .X(n55793) );
  inv_x4_sg U59554 ( .A(n55794), .X(n55795) );
  inv_x4_sg U59555 ( .A(n55796), .X(n55797) );
  inv_x4_sg U59556 ( .A(n55798), .X(n55799) );
  inv_x4_sg U59557 ( .A(n55800), .X(n55801) );
  inv_x4_sg U59558 ( .A(n55802), .X(n55803) );
  inv_x4_sg U59559 ( .A(n55804), .X(n55805) );
  inv_x4_sg U59560 ( .A(n55806), .X(n55807) );
  inv_x4_sg U59561 ( .A(n55808), .X(n55809) );
  inv_x4_sg U59562 ( .A(n55810), .X(n55811) );
  inv_x4_sg U59563 ( .A(n55812), .X(n55813) );
  inv_x4_sg U59564 ( .A(n55814), .X(n55815) );
  inv_x4_sg U59565 ( .A(n55816), .X(n55817) );
  inv_x4_sg U59566 ( .A(n55818), .X(n55819) );
  inv_x4_sg U59567 ( .A(n55820), .X(n55821) );
  inv_x4_sg U59568 ( .A(n55822), .X(n55823) );
  inv_x4_sg U59569 ( .A(n55824), .X(n55825) );
  inv_x4_sg U59570 ( .A(n55826), .X(n55827) );
  inv_x4_sg U59571 ( .A(n55828), .X(n55829) );
  inv_x4_sg U59572 ( .A(n55830), .X(n55831) );
  inv_x4_sg U59573 ( .A(n55832), .X(n55833) );
  inv_x4_sg U59574 ( .A(n55834), .X(n55835) );
  inv_x4_sg U59575 ( .A(n55836), .X(n55837) );
  inv_x4_sg U59576 ( .A(n55838), .X(n55839) );
  inv_x4_sg U59577 ( .A(n55840), .X(n55841) );
  inv_x4_sg U59578 ( .A(n55842), .X(n55843) );
  inv_x4_sg U59579 ( .A(n55844), .X(n55845) );
  inv_x4_sg U59580 ( .A(n55846), .X(n55847) );
  inv_x4_sg U59581 ( .A(n55848), .X(n55849) );
  inv_x4_sg U59582 ( .A(n55850), .X(n55851) );
  inv_x4_sg U59583 ( .A(n55852), .X(n55853) );
  inv_x4_sg U59584 ( .A(n55854), .X(n55855) );
  inv_x4_sg U59585 ( .A(n55856), .X(n55857) );
  inv_x4_sg U59586 ( .A(n55858), .X(n55859) );
  inv_x4_sg U59587 ( .A(n55860), .X(n55861) );
  inv_x4_sg U59588 ( .A(n55862), .X(n55863) );
  inv_x4_sg U59589 ( .A(n55864), .X(n55865) );
  inv_x4_sg U59590 ( .A(n55866), .X(n55867) );
  inv_x4_sg U59591 ( .A(n55868), .X(n55869) );
  inv_x4_sg U59592 ( .A(n55870), .X(n55871) );
  inv_x4_sg U59593 ( .A(n55872), .X(n55873) );
  inv_x4_sg U59594 ( .A(n55874), .X(n55875) );
  inv_x4_sg U59595 ( .A(n55876), .X(n55877) );
  inv_x4_sg U59596 ( .A(n55878), .X(n55879) );
  inv_x4_sg U59597 ( .A(n55880), .X(n55881) );
  inv_x4_sg U59598 ( .A(n55882), .X(n55883) );
  inv_x4_sg U59599 ( .A(n55884), .X(n55885) );
  inv_x4_sg U59600 ( .A(n55886), .X(n55887) );
  inv_x4_sg U59601 ( .A(n55888), .X(n55889) );
  inv_x4_sg U59602 ( .A(n55890), .X(n55891) );
  inv_x4_sg U59603 ( .A(n55892), .X(n55893) );
  inv_x4_sg U59604 ( .A(n55894), .X(n55895) );
  inv_x4_sg U59605 ( .A(n55896), .X(n55897) );
  inv_x4_sg U59606 ( .A(n55898), .X(n55899) );
  inv_x4_sg U59607 ( .A(n55900), .X(n55901) );
  inv_x4_sg U59608 ( .A(n55902), .X(n55903) );
  inv_x4_sg U59609 ( .A(n55904), .X(n55905) );
  inv_x4_sg U59610 ( .A(n55906), .X(n55907) );
  inv_x4_sg U59611 ( .A(n55908), .X(n55909) );
  inv_x4_sg U59612 ( .A(n55910), .X(n55911) );
  inv_x4_sg U59613 ( .A(n55912), .X(n55913) );
  inv_x4_sg U59614 ( .A(n55914), .X(n55915) );
  inv_x4_sg U59615 ( .A(n55916), .X(n55917) );
  inv_x4_sg U59616 ( .A(n55918), .X(n55919) );
  inv_x4_sg U59617 ( .A(n55920), .X(n55921) );
  inv_x4_sg U59618 ( .A(n55922), .X(n55923) );
  inv_x4_sg U59619 ( .A(n55924), .X(n55925) );
  inv_x4_sg U59620 ( .A(n55926), .X(n55927) );
  inv_x4_sg U59621 ( .A(n55928), .X(n55929) );
  inv_x4_sg U59622 ( .A(n55930), .X(n55931) );
  inv_x4_sg U59623 ( .A(n55932), .X(n55933) );
  inv_x4_sg U59624 ( .A(n55934), .X(n55935) );
  inv_x4_sg U59625 ( .A(n55936), .X(n55937) );
  inv_x4_sg U59626 ( .A(n55938), .X(n55939) );
  inv_x4_sg U59627 ( .A(n55940), .X(n55941) );
  inv_x4_sg U59628 ( .A(n55942), .X(n55943) );
  inv_x4_sg U59629 ( .A(n55944), .X(n55945) );
  inv_x4_sg U59630 ( .A(n55946), .X(n55947) );
  inv_x4_sg U59631 ( .A(n55948), .X(n55949) );
  inv_x4_sg U59632 ( .A(n55950), .X(n55951) );
  inv_x4_sg U59633 ( .A(n55952), .X(n55953) );
  inv_x4_sg U59634 ( .A(n55954), .X(n55955) );
  inv_x4_sg U59635 ( .A(n55956), .X(n55957) );
  inv_x4_sg U59636 ( .A(n55958), .X(n55959) );
  inv_x4_sg U59637 ( .A(n55960), .X(n55961) );
  inv_x4_sg U59638 ( .A(n55962), .X(n55963) );
  inv_x4_sg U59639 ( .A(n55964), .X(n55965) );
  inv_x4_sg U59640 ( .A(n55966), .X(n55967) );
  inv_x4_sg U59641 ( .A(n55968), .X(n55969) );
  inv_x4_sg U59642 ( .A(n55970), .X(n55971) );
  inv_x4_sg U59643 ( .A(n55972), .X(n55973) );
  inv_x4_sg U59644 ( .A(n55974), .X(n55975) );
  inv_x4_sg U59645 ( .A(n55976), .X(n55977) );
  inv_x4_sg U59646 ( .A(n55978), .X(n55979) );
  inv_x4_sg U59647 ( .A(n55980), .X(n55981) );
  inv_x4_sg U59648 ( .A(n55982), .X(n55983) );
  inv_x4_sg U59649 ( .A(n55984), .X(n55985) );
  inv_x4_sg U59650 ( .A(n55986), .X(n55987) );
  inv_x4_sg U59651 ( .A(n55988), .X(n55989) );
  inv_x4_sg U59652 ( .A(n55990), .X(n55991) );
  inv_x4_sg U59653 ( .A(n55992), .X(n55993) );
  inv_x4_sg U59654 ( .A(n55994), .X(n55995) );
  inv_x4_sg U59655 ( .A(n55996), .X(n55997) );
  inv_x4_sg U59656 ( .A(n55998), .X(n55999) );
  inv_x4_sg U59657 ( .A(n56000), .X(n56001) );
  inv_x4_sg U59658 ( .A(n56002), .X(n56003) );
  inv_x4_sg U59659 ( .A(n56004), .X(n56005) );
  inv_x4_sg U59660 ( .A(n56006), .X(n56007) );
  inv_x4_sg U59661 ( .A(n56008), .X(n56009) );
  inv_x4_sg U59662 ( .A(n56010), .X(n56011) );
  inv_x4_sg U59663 ( .A(n56012), .X(n56013) );
  inv_x4_sg U59664 ( .A(n56014), .X(n56015) );
  inv_x4_sg U59665 ( .A(n56016), .X(n56017) );
  inv_x4_sg U59666 ( .A(n56018), .X(n56019) );
  inv_x4_sg U59667 ( .A(n56020), .X(n56021) );
  inv_x4_sg U59668 ( .A(n56022), .X(n56023) );
  inv_x4_sg U59669 ( .A(n56024), .X(n56025) );
  inv_x4_sg U59670 ( .A(n56026), .X(n56027) );
  inv_x4_sg U59671 ( .A(n56028), .X(n56029) );
  inv_x4_sg U59672 ( .A(n56030), .X(n56031) );
  inv_x4_sg U59673 ( .A(n56032), .X(n56033) );
  inv_x4_sg U59674 ( .A(n56034), .X(n56035) );
  inv_x4_sg U59675 ( .A(n56036), .X(n56037) );
  inv_x4_sg U59676 ( .A(n56038), .X(n56039) );
  inv_x4_sg U59677 ( .A(n56040), .X(n56041) );
  inv_x4_sg U59678 ( .A(n56042), .X(n56043) );
  inv_x4_sg U59679 ( .A(n56044), .X(n56045) );
  inv_x4_sg U59680 ( .A(n56046), .X(n56047) );
  inv_x4_sg U59681 ( .A(n56048), .X(n56049) );
  inv_x4_sg U59682 ( .A(n56050), .X(n56051) );
  inv_x4_sg U59683 ( .A(n56052), .X(n56053) );
  inv_x4_sg U59684 ( .A(n56054), .X(n56055) );
  inv_x4_sg U59685 ( .A(n56056), .X(n56057) );
  inv_x4_sg U59686 ( .A(n56058), .X(n56059) );
  inv_x4_sg U59687 ( .A(n56060), .X(n56061) );
  inv_x4_sg U59688 ( .A(n56062), .X(n56063) );
  inv_x4_sg U59689 ( .A(n56064), .X(n56065) );
  inv_x4_sg U59690 ( .A(n56066), .X(n56067) );
  inv_x4_sg U59691 ( .A(n56068), .X(n56069) );
  inv_x4_sg U59692 ( .A(n56070), .X(n56071) );
  inv_x4_sg U59693 ( .A(n56072), .X(n56073) );
  inv_x4_sg U59694 ( .A(n56074), .X(n56075) );
  inv_x4_sg U59695 ( .A(n56076), .X(n56077) );
  inv_x4_sg U59696 ( .A(n56078), .X(n56079) );
  inv_x4_sg U59697 ( .A(n56080), .X(n56081) );
  inv_x4_sg U59698 ( .A(n56082), .X(n56083) );
  inv_x4_sg U59699 ( .A(n56084), .X(n56085) );
  inv_x4_sg U59700 ( .A(n56086), .X(n56087) );
  inv_x4_sg U59701 ( .A(n56088), .X(n56089) );
  inv_x4_sg U59702 ( .A(n56090), .X(n56091) );
  inv_x4_sg U59703 ( .A(n56092), .X(n56093) );
  inv_x4_sg U59704 ( .A(n56094), .X(n56095) );
  inv_x4_sg U59705 ( .A(n56096), .X(n56097) );
  inv_x4_sg U59706 ( .A(n56098), .X(n56099) );
  inv_x4_sg U59707 ( .A(n56100), .X(n56101) );
  inv_x4_sg U59708 ( .A(n56102), .X(n56103) );
  inv_x4_sg U59709 ( .A(n56104), .X(n56105) );
  inv_x4_sg U59710 ( .A(n56106), .X(n56107) );
  inv_x4_sg U59711 ( .A(n56108), .X(n56109) );
  inv_x4_sg U59712 ( .A(n56110), .X(n56111) );
  inv_x4_sg U59713 ( .A(n56112), .X(n56113) );
  inv_x4_sg U59714 ( .A(n56114), .X(n56115) );
  inv_x4_sg U59715 ( .A(n56116), .X(n56117) );
  inv_x4_sg U59716 ( .A(n56118), .X(n56119) );
  inv_x4_sg U59717 ( .A(n56120), .X(n56121) );
  inv_x4_sg U59718 ( .A(n56122), .X(n56123) );
  inv_x4_sg U59719 ( .A(n56124), .X(n56125) );
  inv_x4_sg U59720 ( .A(n56126), .X(n56127) );
  inv_x4_sg U59721 ( .A(n56128), .X(n56129) );
  inv_x4_sg U59722 ( .A(n56130), .X(n56131) );
  inv_x4_sg U59723 ( .A(n56132), .X(n56133) );
  inv_x4_sg U59724 ( .A(n56134), .X(n56135) );
  inv_x4_sg U59725 ( .A(n56136), .X(n56137) );
  inv_x4_sg U59726 ( .A(n56138), .X(n56139) );
  inv_x4_sg U59727 ( .A(n56140), .X(n56141) );
  inv_x4_sg U59728 ( .A(n56142), .X(n56143) );
  inv_x4_sg U59729 ( .A(n56144), .X(n56145) );
  inv_x4_sg U59730 ( .A(n56146), .X(n56147) );
  inv_x4_sg U59731 ( .A(n56148), .X(n56149) );
  inv_x4_sg U59732 ( .A(n56150), .X(n56151) );
  inv_x4_sg U59733 ( .A(n56152), .X(n56153) );
  inv_x4_sg U59734 ( .A(n56154), .X(n56155) );
  inv_x4_sg U59735 ( .A(n56156), .X(n56157) );
  inv_x4_sg U59736 ( .A(n56158), .X(n56159) );
  inv_x4_sg U59737 ( .A(n56160), .X(n56161) );
  inv_x4_sg U59738 ( .A(n56162), .X(n56163) );
  inv_x4_sg U59739 ( .A(n56164), .X(n56165) );
  inv_x4_sg U59740 ( .A(n56166), .X(n56167) );
  inv_x4_sg U59741 ( .A(n56168), .X(n56169) );
  inv_x4_sg U59742 ( .A(n56170), .X(n56171) );
  inv_x4_sg U59743 ( .A(n56172), .X(n56173) );
  inv_x4_sg U59744 ( .A(n56174), .X(n56175) );
  inv_x4_sg U59745 ( .A(n56176), .X(n56177) );
  inv_x4_sg U59746 ( .A(n56178), .X(n56179) );
  inv_x4_sg U59747 ( .A(n56180), .X(n56181) );
  inv_x4_sg U59748 ( .A(n56182), .X(n56183) );
  inv_x4_sg U59749 ( .A(n56184), .X(n56185) );
  inv_x4_sg U59750 ( .A(n56186), .X(n56187) );
  inv_x4_sg U59751 ( .A(n56188), .X(n56189) );
  inv_x4_sg U59752 ( .A(n56190), .X(n56191) );
  inv_x4_sg U59753 ( .A(n56192), .X(n56193) );
  inv_x4_sg U59754 ( .A(n56194), .X(n56195) );
  inv_x4_sg U59755 ( .A(n56196), .X(n56197) );
  inv_x4_sg U59756 ( .A(n56198), .X(n56199) );
  inv_x4_sg U59757 ( .A(n56200), .X(n56201) );
  inv_x4_sg U59758 ( .A(n56202), .X(n56203) );
  inv_x4_sg U59759 ( .A(n56204), .X(n56205) );
  inv_x4_sg U59760 ( .A(n56206), .X(n56207) );
  inv_x4_sg U59761 ( .A(n56208), .X(n56209) );
  inv_x4_sg U59762 ( .A(n56210), .X(n56211) );
  inv_x4_sg U59763 ( .A(n56212), .X(n56213) );
  inv_x4_sg U59764 ( .A(n56214), .X(n56215) );
  inv_x4_sg U59765 ( .A(n56216), .X(n56217) );
  inv_x4_sg U59766 ( .A(n56218), .X(n56219) );
  inv_x4_sg U59767 ( .A(n56220), .X(n56221) );
  inv_x4_sg U59768 ( .A(n56222), .X(n56223) );
  inv_x4_sg U59769 ( .A(n56224), .X(n56225) );
  inv_x4_sg U59770 ( .A(n56226), .X(n56227) );
  inv_x4_sg U59771 ( .A(n56228), .X(n56229) );
  inv_x4_sg U59772 ( .A(n56230), .X(n56231) );
  inv_x4_sg U59773 ( .A(n56232), .X(n56233) );
  inv_x4_sg U59774 ( .A(n56234), .X(n56235) );
  inv_x4_sg U59775 ( .A(n56236), .X(n56237) );
  inv_x4_sg U59776 ( .A(n56238), .X(n56239) );
  inv_x4_sg U59777 ( .A(n56240), .X(n56241) );
  inv_x4_sg U59778 ( .A(n56242), .X(n56243) );
  inv_x4_sg U59779 ( .A(n56244), .X(n56245) );
  inv_x4_sg U59780 ( .A(n56246), .X(n56247) );
  inv_x4_sg U59781 ( .A(n56248), .X(n56249) );
  inv_x4_sg U59782 ( .A(n56250), .X(n56251) );
  inv_x4_sg U59783 ( .A(n56252), .X(n56253) );
  inv_x4_sg U59784 ( .A(n56254), .X(n56255) );
  inv_x4_sg U59785 ( .A(n56256), .X(n56257) );
  inv_x4_sg U59786 ( .A(n56258), .X(n56259) );
  inv_x4_sg U59787 ( .A(n56260), .X(n56261) );
  inv_x4_sg U59788 ( .A(n56262), .X(n56263) );
  inv_x4_sg U59789 ( .A(n56264), .X(n56265) );
  inv_x4_sg U59790 ( .A(n56266), .X(n56267) );
  inv_x4_sg U59791 ( .A(n56268), .X(n56269) );
  inv_x4_sg U59792 ( .A(n56270), .X(n56271) );
  inv_x4_sg U59793 ( .A(n56272), .X(n56273) );
  inv_x4_sg U59794 ( .A(n56274), .X(n56275) );
  inv_x4_sg U59795 ( .A(n56276), .X(n56277) );
  inv_x4_sg U59796 ( .A(n56278), .X(n56279) );
  inv_x4_sg U59797 ( .A(n56280), .X(n56281) );
  inv_x4_sg U59798 ( .A(n56282), .X(n56283) );
  inv_x4_sg U59799 ( .A(n56284), .X(n56285) );
  inv_x4_sg U59800 ( .A(n56286), .X(n56287) );
  inv_x4_sg U59801 ( .A(n56288), .X(n56289) );
  inv_x4_sg U59802 ( .A(n56290), .X(n56291) );
  inv_x4_sg U59803 ( .A(n56292), .X(n56293) );
  inv_x4_sg U59804 ( .A(n56294), .X(n56295) );
  inv_x4_sg U59805 ( .A(n56296), .X(n56297) );
  inv_x4_sg U59806 ( .A(n56298), .X(n56299) );
  inv_x4_sg U59807 ( .A(n56300), .X(n56301) );
  inv_x4_sg U59808 ( .A(n56302), .X(n56303) );
  inv_x4_sg U59809 ( .A(n56304), .X(n56305) );
  inv_x4_sg U59810 ( .A(n56306), .X(n56307) );
  inv_x4_sg U59811 ( .A(n56308), .X(n56309) );
  inv_x4_sg U59812 ( .A(n56310), .X(n56311) );
  inv_x4_sg U59813 ( .A(n56312), .X(n56313) );
  inv_x4_sg U59814 ( .A(n56314), .X(n56315) );
  inv_x4_sg U59815 ( .A(n56316), .X(n56317) );
  inv_x4_sg U59816 ( .A(n56318), .X(n56319) );
  inv_x4_sg U59817 ( .A(n56320), .X(n56321) );
  inv_x4_sg U59818 ( .A(n56322), .X(n56323) );
  inv_x4_sg U59819 ( .A(n56324), .X(n56325) );
  inv_x4_sg U59820 ( .A(n56326), .X(n56327) );
  inv_x4_sg U59821 ( .A(n56328), .X(n56329) );
  inv_x4_sg U59822 ( .A(n56330), .X(n56331) );
  inv_x4_sg U59823 ( .A(n56332), .X(n56333) );
  inv_x4_sg U59824 ( .A(n56334), .X(n56335) );
  inv_x4_sg U59825 ( .A(n56336), .X(n56337) );
  inv_x4_sg U59826 ( .A(n56338), .X(n56339) );
  inv_x4_sg U59827 ( .A(n56340), .X(n56341) );
  inv_x4_sg U59828 ( .A(n56342), .X(n56343) );
  inv_x4_sg U59829 ( .A(n56344), .X(n56345) );
  inv_x4_sg U59830 ( .A(n56346), .X(n56347) );
  inv_x4_sg U59831 ( .A(n56348), .X(n56349) );
  inv_x4_sg U59832 ( .A(n56350), .X(n56351) );
  inv_x4_sg U59833 ( .A(n56352), .X(n56353) );
  inv_x4_sg U59834 ( .A(n56354), .X(n56355) );
  inv_x4_sg U59835 ( .A(n56356), .X(n56357) );
  inv_x4_sg U59836 ( .A(n56358), .X(n56359) );
  inv_x4_sg U59837 ( .A(n56360), .X(n56361) );
  inv_x4_sg U59838 ( .A(n56362), .X(n56363) );
  inv_x4_sg U59839 ( .A(n56364), .X(n56365) );
  inv_x4_sg U59840 ( .A(n56366), .X(n56367) );
  inv_x4_sg U59841 ( .A(n56368), .X(n56369) );
  inv_x4_sg U59842 ( .A(n56370), .X(n56371) );
  inv_x4_sg U59843 ( .A(n56372), .X(n56373) );
  inv_x4_sg U59844 ( .A(n56374), .X(n56375) );
  inv_x4_sg U59845 ( .A(n56376), .X(n56377) );
  inv_x4_sg U59846 ( .A(n56378), .X(n56379) );
  inv_x4_sg U59847 ( .A(n56380), .X(n56381) );
  inv_x4_sg U59848 ( .A(n56382), .X(n56383) );
  inv_x4_sg U59849 ( .A(n56384), .X(n56385) );
  inv_x4_sg U59850 ( .A(n56386), .X(n56387) );
  inv_x4_sg U59851 ( .A(n56388), .X(n56389) );
  inv_x4_sg U59852 ( .A(n56390), .X(n56391) );
  inv_x4_sg U59853 ( .A(n56392), .X(n56393) );
  inv_x4_sg U59854 ( .A(n56394), .X(n56395) );
  inv_x4_sg U59855 ( .A(n56396), .X(n56397) );
  inv_x4_sg U59856 ( .A(n56398), .X(n56399) );
  inv_x4_sg U59857 ( .A(n56400), .X(n56401) );
  inv_x4_sg U59858 ( .A(n56402), .X(n56403) );
  inv_x4_sg U59859 ( .A(n56404), .X(n56405) );
  inv_x4_sg U59860 ( .A(n56406), .X(n56407) );
  inv_x4_sg U59861 ( .A(n56408), .X(n56409) );
  inv_x4_sg U59862 ( .A(n56410), .X(n56411) );
  inv_x4_sg U59863 ( .A(n56412), .X(n56413) );
  inv_x4_sg U59864 ( .A(n56414), .X(n56415) );
  inv_x4_sg U59865 ( .A(n56416), .X(n56417) );
  inv_x4_sg U59866 ( .A(n56418), .X(n56419) );
  inv_x4_sg U59867 ( .A(n56420), .X(n56421) );
  inv_x4_sg U59868 ( .A(n56422), .X(n56423) );
  inv_x4_sg U59869 ( .A(n56424), .X(n56425) );
  inv_x4_sg U59870 ( .A(n56426), .X(n56427) );
  inv_x4_sg U59871 ( .A(n56428), .X(n56429) );
  inv_x4_sg U59872 ( .A(n56430), .X(n56431) );
  inv_x4_sg U59873 ( .A(n56432), .X(n56433) );
  inv_x4_sg U59874 ( .A(n56434), .X(n56435) );
  inv_x4_sg U59875 ( .A(n56436), .X(n56437) );
  inv_x4_sg U59876 ( .A(n56438), .X(n56439) );
  inv_x4_sg U59877 ( .A(n56440), .X(n56441) );
  inv_x4_sg U59878 ( .A(n56442), .X(n56443) );
  inv_x4_sg U59879 ( .A(n56444), .X(n56445) );
  inv_x4_sg U59880 ( .A(n56446), .X(n56447) );
  inv_x4_sg U59881 ( .A(n56448), .X(n56449) );
  inv_x4_sg U59882 ( .A(n56450), .X(n56451) );
  inv_x4_sg U59883 ( .A(n56452), .X(n56453) );
  inv_x4_sg U59884 ( .A(n56454), .X(n56455) );
  inv_x4_sg U59885 ( .A(n56456), .X(n56457) );
  inv_x4_sg U59886 ( .A(n56458), .X(n56459) );
  inv_x4_sg U59887 ( .A(n56460), .X(n56461) );
  inv_x4_sg U59888 ( .A(n56462), .X(n56463) );
  inv_x4_sg U59889 ( .A(n56464), .X(n56465) );
  inv_x4_sg U59890 ( .A(n56466), .X(n56467) );
  inv_x4_sg U59891 ( .A(n56468), .X(n56469) );
  inv_x4_sg U59892 ( .A(n56470), .X(n56471) );
  inv_x4_sg U59893 ( .A(n56472), .X(n56473) );
  inv_x4_sg U59894 ( .A(n56474), .X(n56475) );
  inv_x4_sg U59895 ( .A(n56476), .X(n56477) );
  inv_x4_sg U59896 ( .A(n56478), .X(n56479) );
  inv_x4_sg U59897 ( .A(n56480), .X(n56481) );
  inv_x4_sg U59898 ( .A(n56482), .X(n56483) );
  inv_x4_sg U59899 ( .A(n56484), .X(n56485) );
  inv_x4_sg U59900 ( .A(n56486), .X(n56487) );
  inv_x4_sg U59901 ( .A(n56488), .X(n56489) );
  inv_x4_sg U59902 ( .A(n56490), .X(n56491) );
  inv_x4_sg U59903 ( .A(n56492), .X(n56493) );
  inv_x4_sg U59904 ( .A(n56494), .X(n56495) );
  inv_x4_sg U59905 ( .A(n56496), .X(n56497) );
  inv_x4_sg U59906 ( .A(n56498), .X(n56499) );
  inv_x4_sg U59907 ( .A(n56500), .X(n56501) );
  inv_x4_sg U59908 ( .A(n56502), .X(n56503) );
  inv_x4_sg U59909 ( .A(n56504), .X(n56505) );
  inv_x4_sg U59910 ( .A(n56506), .X(n56507) );
  inv_x4_sg U59911 ( .A(n56508), .X(n56509) );
  inv_x4_sg U59912 ( .A(n56510), .X(n56511) );
  inv_x4_sg U59913 ( .A(n56512), .X(n56513) );
  inv_x4_sg U59914 ( .A(n56514), .X(n56515) );
  inv_x4_sg U59915 ( .A(n56516), .X(n56517) );
  inv_x4_sg U59916 ( .A(n56518), .X(n56519) );
  inv_x4_sg U59917 ( .A(n56520), .X(n56521) );
  inv_x4_sg U59918 ( .A(n56522), .X(n56523) );
  inv_x4_sg U59919 ( .A(n56524), .X(n56525) );
  inv_x4_sg U59920 ( .A(n56526), .X(n56527) );
  inv_x4_sg U59921 ( .A(n56528), .X(n56529) );
  inv_x4_sg U59922 ( .A(n56530), .X(n56531) );
  inv_x4_sg U59923 ( .A(n56532), .X(n56533) );
  inv_x4_sg U59924 ( .A(n56534), .X(n56535) );
  inv_x4_sg U59925 ( .A(n56536), .X(n56537) );
  inv_x4_sg U59926 ( .A(n56538), .X(n56539) );
  inv_x4_sg U59927 ( .A(n56540), .X(n56541) );
  inv_x4_sg U59928 ( .A(n56542), .X(n56543) );
  inv_x4_sg U59929 ( .A(n56544), .X(n56545) );
  inv_x4_sg U59930 ( .A(n56546), .X(n56547) );
  inv_x4_sg U59931 ( .A(n56548), .X(n56549) );
  inv_x4_sg U59932 ( .A(n56550), .X(n56551) );
  inv_x4_sg U59933 ( .A(n56552), .X(n56553) );
  inv_x4_sg U59934 ( .A(n56554), .X(n56555) );
  inv_x4_sg U59935 ( .A(n56556), .X(n56557) );
  inv_x4_sg U59936 ( .A(n56558), .X(n56559) );
  inv_x4_sg U59937 ( .A(n56560), .X(n56561) );
  inv_x4_sg U59938 ( .A(n56562), .X(n56563) );
  inv_x4_sg U59939 ( .A(n56564), .X(n56565) );
  inv_x4_sg U59940 ( .A(n56566), .X(n56567) );
  inv_x4_sg U59941 ( .A(n56568), .X(n56569) );
  inv_x4_sg U59942 ( .A(n56570), .X(n56571) );
  inv_x4_sg U59943 ( .A(n56572), .X(n56573) );
  inv_x4_sg U59944 ( .A(n56574), .X(n56575) );
  inv_x4_sg U59945 ( .A(n56576), .X(n56577) );
  inv_x4_sg U59946 ( .A(n56578), .X(n56579) );
  inv_x4_sg U59947 ( .A(n56580), .X(n56581) );
  inv_x4_sg U59948 ( .A(n56582), .X(n56583) );
  inv_x4_sg U59949 ( .A(n56584), .X(n56585) );
  inv_x4_sg U59950 ( .A(n56586), .X(n56587) );
  inv_x4_sg U59951 ( .A(n56588), .X(n56589) );
  inv_x4_sg U59952 ( .A(n56590), .X(n56591) );
  inv_x4_sg U59953 ( .A(n56592), .X(n56593) );
  inv_x4_sg U59954 ( .A(n56594), .X(n56595) );
  inv_x4_sg U59955 ( .A(n47283), .X(n56596) );
  inv_x8_sg U59956 ( .A(n56596), .X(o_mask[0]) );
  inv_x8_sg U59957 ( .A(o_mask[0]), .X(n68337) );
  inv_x4_sg U59958 ( .A(n47281), .X(n56598) );
  inv_x8_sg U59959 ( .A(n56598), .X(o_mask[1]) );
  inv_x8_sg U59960 ( .A(o_mask[1]), .X(n68338) );
  inv_x4_sg U59961 ( .A(n47279), .X(n56600) );
  inv_x8_sg U59962 ( .A(n56600), .X(o_mask[2]) );
  inv_x8_sg U59963 ( .A(o_mask[2]), .X(n68339) );
  inv_x4_sg U59964 ( .A(n47277), .X(n56602) );
  inv_x8_sg U59965 ( .A(n56602), .X(o_mask[3]) );
  inv_x8_sg U59966 ( .A(o_mask[3]), .X(n68340) );
  inv_x4_sg U59967 ( .A(n47275), .X(n56604) );
  inv_x8_sg U59968 ( .A(n56604), .X(o_mask[4]) );
  inv_x8_sg U59969 ( .A(o_mask[4]), .X(n68341) );
  inv_x4_sg U59970 ( .A(n47273), .X(n56606) );
  inv_x8_sg U59971 ( .A(n56606), .X(o_mask[5]) );
  inv_x8_sg U59972 ( .A(o_mask[5]), .X(n68342) );
  inv_x4_sg U59973 ( .A(n47271), .X(n56608) );
  inv_x8_sg U59974 ( .A(n56608), .X(o_mask[6]) );
  inv_x8_sg U59975 ( .A(o_mask[6]), .X(n68343) );
  inv_x4_sg U59976 ( .A(n47269), .X(n56610) );
  inv_x8_sg U59977 ( .A(n56610), .X(o_mask[7]) );
  inv_x8_sg U59978 ( .A(o_mask[7]), .X(n68344) );
  inv_x4_sg U59979 ( .A(n47267), .X(n56612) );
  inv_x8_sg U59980 ( .A(n56612), .X(o_mask[8]) );
  inv_x8_sg U59981 ( .A(o_mask[8]), .X(n68345) );
  inv_x4_sg U59982 ( .A(n47265), .X(n56614) );
  inv_x8_sg U59983 ( .A(n56614), .X(o_mask[9]) );
  inv_x8_sg U59984 ( .A(o_mask[9]), .X(n68346) );
  inv_x4_sg U59985 ( .A(n47263), .X(n56616) );
  inv_x8_sg U59986 ( .A(n56616), .X(o_mask[10]) );
  inv_x8_sg U59987 ( .A(o_mask[10]), .X(n68347) );
  inv_x4_sg U59988 ( .A(n47261), .X(n56618) );
  inv_x8_sg U59989 ( .A(n56618), .X(o_mask[11]) );
  inv_x8_sg U59990 ( .A(o_mask[11]), .X(n68348) );
  inv_x4_sg U59991 ( .A(n47259), .X(n56620) );
  inv_x8_sg U59992 ( .A(n56620), .X(o_mask[12]) );
  inv_x8_sg U59993 ( .A(o_mask[12]), .X(n68349) );
  inv_x4_sg U59994 ( .A(n47257), .X(n56622) );
  inv_x8_sg U59995 ( .A(n56622), .X(o_mask[13]) );
  inv_x8_sg U59996 ( .A(o_mask[13]), .X(n68350) );
  inv_x4_sg U59997 ( .A(n47255), .X(n56624) );
  inv_x8_sg U59998 ( .A(n56624), .X(o_mask[14]) );
  inv_x8_sg U59999 ( .A(o_mask[14]), .X(n68351) );
  inv_x4_sg U60000 ( .A(n47253), .X(n56626) );
  inv_x8_sg U60001 ( .A(n56626), .X(o_mask[15]) );
  inv_x8_sg U60002 ( .A(o_mask[15]), .X(n68352) );
  inv_x4_sg U60003 ( .A(n47251), .X(n56628) );
  inv_x8_sg U60004 ( .A(n56628), .X(o_mask[16]) );
  inv_x8_sg U60005 ( .A(o_mask[16]), .X(n68353) );
  inv_x4_sg U60006 ( .A(n47249), .X(n56630) );
  inv_x8_sg U60007 ( .A(n56630), .X(o_mask[17]) );
  inv_x8_sg U60008 ( .A(o_mask[17]), .X(n68354) );
  inv_x4_sg U60009 ( .A(n47247), .X(n56632) );
  inv_x8_sg U60010 ( .A(n56632), .X(o_mask[18]) );
  inv_x8_sg U60011 ( .A(o_mask[18]), .X(n68355) );
  inv_x4_sg U60012 ( .A(n47245), .X(n56634) );
  inv_x8_sg U60013 ( .A(n56634), .X(o_mask[19]) );
  inv_x8_sg U60014 ( .A(o_mask[19]), .X(n68356) );
  inv_x4_sg U60015 ( .A(n47243), .X(n56636) );
  inv_x8_sg U60016 ( .A(n56636), .X(o_mask[20]) );
  inv_x8_sg U60017 ( .A(o_mask[20]), .X(n68357) );
  inv_x4_sg U60018 ( .A(n47241), .X(n56638) );
  inv_x8_sg U60019 ( .A(n56638), .X(o_mask[21]) );
  inv_x8_sg U60020 ( .A(o_mask[21]), .X(n68358) );
  inv_x4_sg U60021 ( .A(n47239), .X(n56640) );
  inv_x8_sg U60022 ( .A(n56640), .X(o_mask[22]) );
  inv_x8_sg U60023 ( .A(o_mask[22]), .X(n68359) );
  inv_x4_sg U60024 ( .A(n47237), .X(n56642) );
  inv_x8_sg U60025 ( .A(n56642), .X(o_mask[23]) );
  inv_x8_sg U60026 ( .A(o_mask[23]), .X(n68360) );
  inv_x4_sg U60027 ( .A(n47235), .X(n56644) );
  inv_x8_sg U60028 ( .A(n56644), .X(o_mask[24]) );
  inv_x8_sg U60029 ( .A(o_mask[24]), .X(n68361) );
  inv_x4_sg U60030 ( .A(n47233), .X(n56646) );
  inv_x8_sg U60031 ( .A(n56646), .X(o_mask[25]) );
  inv_x8_sg U60032 ( .A(o_mask[25]), .X(n68362) );
  inv_x4_sg U60033 ( .A(n47231), .X(n56648) );
  inv_x8_sg U60034 ( .A(n56648), .X(o_mask[26]) );
  inv_x8_sg U60035 ( .A(o_mask[26]), .X(n68363) );
  inv_x4_sg U60036 ( .A(n47229), .X(n56650) );
  inv_x8_sg U60037 ( .A(n56650), .X(o_mask[27]) );
  inv_x8_sg U60038 ( .A(o_mask[27]), .X(n68364) );
  inv_x4_sg U60039 ( .A(n47227), .X(n56652) );
  inv_x8_sg U60040 ( .A(n56652), .X(o_mask[28]) );
  inv_x8_sg U60041 ( .A(o_mask[28]), .X(n68365) );
  inv_x4_sg U60042 ( .A(n47225), .X(n56654) );
  inv_x8_sg U60043 ( .A(n56654), .X(o_mask[29]) );
  inv_x8_sg U60044 ( .A(o_mask[29]), .X(n68366) );
  inv_x4_sg U60045 ( .A(n47223), .X(n56656) );
  inv_x8_sg U60046 ( .A(n56656), .X(o_mask[30]) );
  inv_x8_sg U60047 ( .A(o_mask[30]), .X(n68367) );
  inv_x4_sg U60048 ( .A(n47221), .X(n56658) );
  inv_x8_sg U60049 ( .A(n56658), .X(o_mask[31]) );
  inv_x8_sg U60050 ( .A(o_mask[31]), .X(n68368) );
  inv_x4_sg U60051 ( .A(n56660), .X(n56661) );
  inv_x4_sg U60052 ( .A(n56662), .X(n56663) );
  inv_x4_sg U60053 ( .A(n56664), .X(n56665) );
  inv_x4_sg U60054 ( .A(n56666), .X(n56667) );
  inv_x4_sg U60055 ( .A(n56668), .X(n56669) );
  inv_x4_sg U60056 ( .A(n56670), .X(n56671) );
  inv_x4_sg U60057 ( .A(n56672), .X(n56673) );
  inv_x4_sg U60058 ( .A(n56674), .X(n56675) );
  inv_x4_sg U60059 ( .A(n56676), .X(n56677) );
  inv_x4_sg U60060 ( .A(n56678), .X(n56679) );
  inv_x4_sg U60061 ( .A(n56680), .X(n56681) );
  inv_x4_sg U60062 ( .A(n56682), .X(n56683) );
  inv_x4_sg U60063 ( .A(n56684), .X(n56685) );
  inv_x4_sg U60064 ( .A(n56686), .X(n56687) );
  inv_x4_sg U60065 ( .A(n56688), .X(n56689) );
  inv_x4_sg U60066 ( .A(n56690), .X(n56691) );
  inv_x4_sg U60067 ( .A(n56692), .X(n56693) );
  inv_x4_sg U60068 ( .A(n56694), .X(n56695) );
  inv_x4_sg U60069 ( .A(n56696), .X(n56697) );
  inv_x4_sg U60070 ( .A(n56698), .X(n56699) );
  inv_x4_sg U60071 ( .A(n56700), .X(n56701) );
  inv_x4_sg U60072 ( .A(n56702), .X(n56703) );
  inv_x4_sg U60073 ( .A(n56704), .X(n56705) );
  inv_x4_sg U60074 ( .A(n56706), .X(n56707) );
  inv_x4_sg U60075 ( .A(n56708), .X(n56709) );
  inv_x4_sg U60076 ( .A(n56710), .X(n56711) );
  inv_x4_sg U60077 ( .A(n56712), .X(n56713) );
  inv_x4_sg U60078 ( .A(n56714), .X(n56715) );
  inv_x4_sg U60079 ( .A(n56716), .X(n56717) );
  inv_x4_sg U60080 ( .A(n56718), .X(n56719) );
  inv_x4_sg U60081 ( .A(n56720), .X(n56721) );
  inv_x4_sg U60082 ( .A(n56722), .X(n56723) );
  inv_x4_sg U60083 ( .A(n56724), .X(n56725) );
  inv_x4_sg U60084 ( .A(n56726), .X(n56727) );
  inv_x4_sg U60085 ( .A(n56728), .X(n56729) );
  inv_x4_sg U60086 ( .A(n56730), .X(n56731) );
  inv_x4_sg U60087 ( .A(n56732), .X(n56733) );
  inv_x4_sg U60088 ( .A(n56734), .X(n56735) );
  inv_x4_sg U60089 ( .A(n56736), .X(n56737) );
  inv_x4_sg U60090 ( .A(n56738), .X(n56739) );
  inv_x4_sg U60091 ( .A(n56740), .X(n56741) );
  inv_x4_sg U60092 ( .A(n56742), .X(n56743) );
  inv_x4_sg U60093 ( .A(n56744), .X(n56745) );
  inv_x4_sg U60094 ( .A(n56746), .X(n56747) );
  inv_x4_sg U60095 ( .A(n56748), .X(n56749) );
  inv_x4_sg U60096 ( .A(n56750), .X(n56751) );
  inv_x4_sg U60097 ( .A(n56752), .X(n56753) );
  inv_x4_sg U60098 ( .A(n56754), .X(n56755) );
  inv_x4_sg U60099 ( .A(n56756), .X(n56757) );
  inv_x4_sg U60100 ( .A(n56758), .X(n56759) );
  inv_x4_sg U60101 ( .A(n56760), .X(n56761) );
  inv_x4_sg U60102 ( .A(n56762), .X(n56763) );
  inv_x4_sg U60103 ( .A(n56764), .X(n56765) );
  inv_x4_sg U60104 ( .A(n56766), .X(n56767) );
  inv_x4_sg U60105 ( .A(n56768), .X(n56769) );
  inv_x4_sg U60106 ( .A(n56770), .X(n56771) );
  inv_x4_sg U60107 ( .A(n56772), .X(n56773) );
  inv_x4_sg U60108 ( .A(n56774), .X(n56775) );
  inv_x4_sg U60109 ( .A(n56776), .X(n56777) );
  inv_x4_sg U60110 ( .A(n56778), .X(n56779) );
  inv_x4_sg U60111 ( .A(n56780), .X(n56781) );
  inv_x4_sg U60112 ( .A(n56782), .X(n56783) );
  inv_x4_sg U60113 ( .A(n56784), .X(n56785) );
  inv_x4_sg U60114 ( .A(n56786), .X(n56787) );
  inv_x4_sg U60115 ( .A(n56788), .X(n56789) );
  inv_x4_sg U60116 ( .A(n56790), .X(n56791) );
  inv_x4_sg U60117 ( .A(n56792), .X(n56793) );
  inv_x4_sg U60118 ( .A(n56794), .X(n56795) );
  inv_x4_sg U60119 ( .A(n56796), .X(n56797) );
  inv_x4_sg U60120 ( .A(n56798), .X(n56799) );
  inv_x4_sg U60121 ( .A(n56800), .X(n56801) );
  inv_x4_sg U60122 ( .A(n56802), .X(n56803) );
  inv_x4_sg U60123 ( .A(n56804), .X(n56805) );
  inv_x4_sg U60124 ( .A(n56806), .X(n56807) );
  inv_x4_sg U60125 ( .A(n56808), .X(n56809) );
  inv_x4_sg U60126 ( .A(n56810), .X(n56811) );
  inv_x4_sg U60127 ( .A(n56812), .X(n56813) );
  inv_x4_sg U60128 ( .A(n56814), .X(n56815) );
  inv_x4_sg U60129 ( .A(n56816), .X(n56817) );
  inv_x4_sg U60130 ( .A(n56818), .X(n56819) );
  inv_x4_sg U60131 ( .A(n56820), .X(n56821) );
  inv_x4_sg U60132 ( .A(n56822), .X(n56823) );
  inv_x4_sg U60133 ( .A(n56824), .X(n56825) );
  inv_x4_sg U60134 ( .A(n56826), .X(n56827) );
  inv_x4_sg U60135 ( .A(n56828), .X(n56829) );
  inv_x4_sg U60136 ( .A(n56830), .X(n56831) );
  inv_x4_sg U60137 ( .A(n56832), .X(n56833) );
  inv_x4_sg U60138 ( .A(n56834), .X(n56835) );
  inv_x4_sg U60139 ( .A(n56836), .X(n56837) );
  inv_x4_sg U60140 ( .A(n56838), .X(n56839) );
  inv_x4_sg U60141 ( .A(n56840), .X(n56841) );
  inv_x4_sg U60142 ( .A(n56842), .X(n56843) );
  inv_x4_sg U60143 ( .A(n56844), .X(n56845) );
  inv_x4_sg U60144 ( .A(n56846), .X(n56847) );
  inv_x4_sg U60145 ( .A(n56848), .X(n56849) );
  inv_x4_sg U60146 ( .A(n56850), .X(n56851) );
  inv_x4_sg U60147 ( .A(n56852), .X(n56853) );
  inv_x4_sg U60148 ( .A(n56854), .X(n56855) );
  inv_x4_sg U60149 ( .A(n56856), .X(n56857) );
  inv_x4_sg U60150 ( .A(n56858), .X(n56859) );
  inv_x4_sg U60151 ( .A(n56860), .X(n56861) );
  inv_x4_sg U60152 ( .A(n56862), .X(n56863) );
  inv_x4_sg U60153 ( .A(n56864), .X(n56865) );
  inv_x4_sg U60154 ( .A(n56866), .X(n56867) );
  inv_x4_sg U60155 ( .A(n56868), .X(n56869) );
  inv_x4_sg U60156 ( .A(n56870), .X(n56871) );
  inv_x4_sg U60157 ( .A(n56872), .X(n56873) );
  inv_x4_sg U60158 ( .A(n56874), .X(n56875) );
  inv_x4_sg U60159 ( .A(n56876), .X(n56877) );
  inv_x4_sg U60160 ( .A(n56878), .X(n56879) );
  inv_x4_sg U60161 ( .A(n56880), .X(n56881) );
  inv_x4_sg U60162 ( .A(n56882), .X(n56883) );
  inv_x4_sg U60163 ( .A(n56884), .X(n56885) );
  inv_x4_sg U60164 ( .A(n56886), .X(n56887) );
  inv_x4_sg U60165 ( .A(n56888), .X(n56889) );
  inv_x4_sg U60166 ( .A(n56890), .X(n56891) );
  inv_x4_sg U60167 ( .A(n56892), .X(n56893) );
  inv_x4_sg U60168 ( .A(n56894), .X(n56895) );
  inv_x4_sg U60169 ( .A(n56896), .X(n56897) );
  inv_x4_sg U60170 ( .A(n56898), .X(n56899) );
  inv_x4_sg U60171 ( .A(n56900), .X(n56901) );
  inv_x4_sg U60172 ( .A(n56902), .X(n56903) );
  inv_x4_sg U60173 ( .A(n56904), .X(n56905) );
  inv_x4_sg U60174 ( .A(n56906), .X(n56907) );
  inv_x4_sg U60175 ( .A(n56908), .X(n56909) );
  inv_x4_sg U60176 ( .A(n56910), .X(n56911) );
  inv_x4_sg U60177 ( .A(n56912), .X(n56913) );
  inv_x4_sg U60178 ( .A(n56914), .X(n56915) );
  inv_x4_sg U60179 ( .A(n47181), .X(n56916) );
  inv_x4_sg U60180 ( .A(n47175), .X(n56918) );
  inv_x4_sg U60181 ( .A(n47171), .X(n56920) );
  inv_x4_sg U60182 ( .A(n47037), .X(n56922) );
  inv_x4_sg U60183 ( .A(n47031), .X(n56924) );
  inv_x4_sg U60184 ( .A(n47027), .X(n56926) );
  inv_x4_sg U60185 ( .A(n47215), .X(n56928) );
  inv_x4_sg U60186 ( .A(n47165), .X(n56930) );
  inv_x4_sg U60187 ( .A(n47021), .X(n56932) );
  inv_x4_sg U60188 ( .A(n47211), .X(n56934) );
  inv_x8_sg U60189 ( .A(n56934), .X(n56935) );
  inv_x8_sg U60190 ( .A(n56935), .X(n67534) );
  inv_x8_sg U60191 ( .A(n58640), .X(n58478) );
  inv_x4_sg U60192 ( .A(n47155), .X(n56936) );
  inv_x4_sg U60193 ( .A(n47153), .X(n56938) );
  inv_x4_sg U60194 ( .A(n47145), .X(n56940) );
  inv_x4_sg U60195 ( .A(n47143), .X(n56942) );
  inv_x4_sg U60196 ( .A(n47137), .X(n56944) );
  inv_x4_sg U60197 ( .A(n47135), .X(n56946) );
  inv_x4_sg U60198 ( .A(n47127), .X(n56948) );
  inv_x4_sg U60199 ( .A(n47125), .X(n56950) );
  inv_x4_sg U60200 ( .A(n47011), .X(n56952) );
  inv_x4_sg U60201 ( .A(n47009), .X(n56954) );
  inv_x4_sg U60202 ( .A(n47001), .X(n56956) );
  inv_x4_sg U60203 ( .A(n46999), .X(n56958) );
  inv_x4_sg U60204 ( .A(n46993), .X(n56960) );
  inv_x4_sg U60205 ( .A(n46991), .X(n56962) );
  inv_x4_sg U60206 ( .A(n46983), .X(n56964) );
  inv_x4_sg U60207 ( .A(n46981), .X(n56966) );
  inv_x4_sg U60208 ( .A(n47203), .X(n56968) );
  inv_x8_sg U60209 ( .A(n56968), .X(n56969) );
  inv_x4_sg U60210 ( .A(n47195), .X(n56970) );
  inv_x8_sg U60211 ( .A(n56970), .X(n56971) );
  inv_x8_sg U60212 ( .A(n26047), .X(n67536) );
  inv_x4_sg U60213 ( .A(n47049), .X(n56972) );
  inv_x8_sg U60214 ( .A(n56972), .X(n56973) );
  inv_x4_sg U60215 ( .A(n47047), .X(n56974) );
  inv_x8_sg U60216 ( .A(n56974), .X(n56975) );
  inv_x4_sg U60217 ( .A(n47057), .X(n56976) );
  inv_x8_sg U60218 ( .A(n56976), .X(n56977) );
  inv_x4_sg U60219 ( .A(n46923), .X(n56978) );
  inv_x8_sg U60220 ( .A(n56978), .X(n56979) );
  inv_x4_sg U60221 ( .A(n46921), .X(n56980) );
  inv_x8_sg U60222 ( .A(n56980), .X(n56981) );
  inv_x4_sg U60223 ( .A(n46929), .X(n56982) );
  inv_x8_sg U60224 ( .A(n56982), .X(n56983) );
  inv_x4_sg U60225 ( .A(n46927), .X(n56984) );
  inv_x8_sg U60226 ( .A(n56984), .X(n56985) );
  inv_x4_sg U60227 ( .A(n47077), .X(n56986) );
  inv_x8_sg U60228 ( .A(n56986), .X(n56987) );
  inv_x4_sg U60229 ( .A(n47075), .X(n56988) );
  inv_x8_sg U60230 ( .A(n56988), .X(n56989) );
  inv_x4_sg U60231 ( .A(n47071), .X(n56990) );
  inv_x8_sg U60232 ( .A(n56990), .X(n56991) );
  inv_x4_sg U60233 ( .A(n47069), .X(n56992) );
  inv_x8_sg U60234 ( .A(n56992), .X(n56993) );
  inv_x4_sg U60235 ( .A(n46899), .X(n56994) );
  inv_x8_sg U60236 ( .A(n56994), .X(n56995) );
  inv_x4_sg U60237 ( .A(n46901), .X(n56996) );
  inv_x8_sg U60238 ( .A(n56996), .X(n56997) );
  inv_x4_sg U60239 ( .A(n47059), .X(n56998) );
  inv_x8_sg U60240 ( .A(n56998), .X(n56999) );
  inv_x4_sg U60241 ( .A(n46911), .X(n57000) );
  inv_x8_sg U60242 ( .A(n57000), .X(n57001) );
  inv_x4_sg U60243 ( .A(n46909), .X(n57002) );
  inv_x8_sg U60244 ( .A(n57002), .X(n57003) );
  inv_x4_sg U60245 ( .A(n47065), .X(n57004) );
  inv_x8_sg U60246 ( .A(n57004), .X(n57005) );
  inv_x4_sg U60247 ( .A(n47063), .X(n57006) );
  inv_x8_sg U60248 ( .A(n57006), .X(n57007) );
  inv_x4_sg U60249 ( .A(n46917), .X(n57008) );
  inv_x8_sg U60250 ( .A(n57008), .X(n57009) );
  inv_x4_sg U60251 ( .A(n46915), .X(n57010) );
  inv_x8_sg U60252 ( .A(n57010), .X(n57011) );
  inv_x4_sg U60253 ( .A(n46963), .X(n57012) );
  inv_x8_sg U60254 ( .A(n57012), .X(n57013) );
  inv_x4_sg U60255 ( .A(n46969), .X(n57014) );
  inv_x8_sg U60256 ( .A(n57014), .X(n57015) );
  inv_x4_sg U60257 ( .A(n47107), .X(n57016) );
  inv_x8_sg U60258 ( .A(n57016), .X(n57017) );
  inv_x4_sg U60259 ( .A(n47099), .X(n57018) );
  inv_x8_sg U60260 ( .A(n57018), .X(n57019) );
  inv_x4_sg U60261 ( .A(n46955), .X(n57020) );
  inv_x8_sg U60262 ( .A(n57020), .X(n57021) );
  inv_x4_sg U60263 ( .A(n47089), .X(n57022) );
  inv_x8_sg U60264 ( .A(n57022), .X(n57023) );
  inv_x4_sg U60265 ( .A(n47083), .X(n57024) );
  inv_x8_sg U60266 ( .A(n57024), .X(n57025) );
  inv_x4_sg U60267 ( .A(n46945), .X(n57026) );
  inv_x8_sg U60268 ( .A(n57026), .X(n57027) );
  inv_x4_sg U60269 ( .A(n46939), .X(n57028) );
  inv_x8_sg U60270 ( .A(n57028), .X(n57029) );
  inv_x4_sg U60271 ( .A(n47113), .X(n57030) );
  inv_x8_sg U60272 ( .A(n57030), .X(n57031) );
  inv_x4_sg U60273 ( .A(n47103), .X(n57032) );
  inv_x8_sg U60274 ( .A(n57032), .X(n57033) );
  inv_x4_sg U60275 ( .A(n47095), .X(n57034) );
  inv_x8_sg U60276 ( .A(n57034), .X(n57035) );
  inv_x4_sg U60277 ( .A(n47085), .X(n57036) );
  inv_x8_sg U60278 ( .A(n57036), .X(n57037) );
  inv_x4_sg U60279 ( .A(n46959), .X(n57038) );
  inv_x8_sg U60280 ( .A(n57038), .X(n57039) );
  inv_x4_sg U60281 ( .A(n46951), .X(n57040) );
  inv_x8_sg U60282 ( .A(n57040), .X(n57041) );
  inv_x4_sg U60283 ( .A(n46941), .X(n57042) );
  inv_x8_sg U60284 ( .A(n57042), .X(n57043) );
  inv_x4_sg U60285 ( .A(n46933), .X(n57044) );
  inv_x8_sg U60286 ( .A(n57044), .X(n57045) );
  inv_x4_sg U60287 ( .A(n47081), .X(n57046) );
  inv_x8_sg U60288 ( .A(n57046), .X(n57047) );
  inv_x8_sg U60289 ( .A(n30624), .X(n61905) );
  nand_x2_sg U60290 ( .A(n57962), .B(n61905), .X(n57963) );
  inv_x4_sg U60291 ( .A(n47147), .X(n57048) );
  inv_x8_sg U60292 ( .A(n57048), .X(n57049) );
  inv_x4_sg U60293 ( .A(n47139), .X(n57050) );
  inv_x8_sg U60294 ( .A(n57050), .X(n57051) );
  inv_x4_sg U60295 ( .A(n47131), .X(n57052) );
  inv_x8_sg U60296 ( .A(n57052), .X(n57053) );
  inv_x4_sg U60297 ( .A(n47123), .X(n57054) );
  inv_x8_sg U60298 ( .A(n57054), .X(n57055) );
  inv_x4_sg U60299 ( .A(n47003), .X(n57056) );
  inv_x8_sg U60300 ( .A(n57056), .X(n57057) );
  inv_x4_sg U60301 ( .A(n46995), .X(n57058) );
  inv_x8_sg U60302 ( .A(n57058), .X(n57059) );
  inv_x4_sg U60303 ( .A(n46987), .X(n57060) );
  inv_x8_sg U60304 ( .A(n57060), .X(n57061) );
  inv_x4_sg U60305 ( .A(n46979), .X(n57062) );
  inv_x8_sg U60306 ( .A(n57062), .X(n57063) );
  inv_x4_sg U60307 ( .A(n47129), .X(n57064) );
  inv_x8_sg U60308 ( .A(n57064), .X(n57065) );
  inv_x4_sg U60309 ( .A(n46985), .X(n57066) );
  inv_x8_sg U60310 ( .A(n57066), .X(n57067) );
  inv_x8_sg U60311 ( .A(n22445), .X(n67499) );
  nand_x8_sg U60312 ( .A(n57862), .B(n67499), .X(n22740) );
  nor_x8_sg U60313 ( .A(n68576), .B(n68575), .X(n22467) );
  inv_x8_sg U60314 ( .A(n57298), .X(n68575) );
  inv_x4_sg U60315 ( .A(n47213), .X(n57068) );
  inv_x8_sg U60316 ( .A(n57068), .X(n57069) );
  inv_x8_sg U60317 ( .A(n57069), .X(n68373) );
  inv_x4_sg U60318 ( .A(n46919), .X(n57070) );
  inv_x8_sg U60319 ( .A(n57070), .X(n57071) );
  inv_x4_sg U60320 ( .A(n47079), .X(n57072) );
  inv_x8_sg U60321 ( .A(n57072), .X(n57073) );
  inv_x4_sg U60322 ( .A(n47067), .X(n57074) );
  inv_x8_sg U60323 ( .A(n57074), .X(n57075) );
  inv_x4_sg U60324 ( .A(n47061), .X(n57076) );
  inv_x8_sg U60325 ( .A(n57076), .X(n57077) );
  inv_x4_sg U60326 ( .A(n46913), .X(n57078) );
  inv_x8_sg U60327 ( .A(n57078), .X(n57079) );
  inv_x4_sg U60328 ( .A(n46895), .X(n57080) );
  inv_x8_sg U60329 ( .A(n57080), .X(n57081) );
  inv_x4_sg U60330 ( .A(n47053), .X(n57082) );
  inv_x8_sg U60331 ( .A(n57082), .X(n57083) );
  inv_x4_sg U60332 ( .A(n47051), .X(n57084) );
  inv_x8_sg U60333 ( .A(n57084), .X(n57085) );
  inv_x4_sg U60334 ( .A(n46905), .X(n57086) );
  inv_x8_sg U60335 ( .A(n57086), .X(n57087) );
  inv_x4_sg U60336 ( .A(n46903), .X(n57088) );
  inv_x8_sg U60337 ( .A(n57088), .X(n57089) );
  inv_x8_sg U60338 ( .A(n57099), .X(n58616) );
  inv_x8_sg U60339 ( .A(n57302), .X(n68397) );
  inv_x4_sg U60340 ( .A(n47209), .X(n57090) );
  inv_x8_sg U60341 ( .A(n57090), .X(n57091) );
  inv_x8_sg U60342 ( .A(n57091), .X(n67530) );
  inv_x4_sg U60343 ( .A(n34088), .X(n57092) );
  inv_x8_sg U60344 ( .A(n57092), .X(n57093) );
  nor_x8_sg U60345 ( .A(n34087), .B(n57093), .X(n33309) );
  nand_x8_sg U60346 ( .A(n33396), .B(n34221), .X(n34087) );
  inv_x4_sg U60347 ( .A(n34175), .X(n57094) );
  inv_x8_sg U60348 ( .A(n57094), .X(n57095) );
  nor_x8_sg U60349 ( .A(n33911), .B(n57095), .X(n33222) );
  nand_x8_sg U60350 ( .A(n33396), .B(n34176), .X(n33911) );
  inv_x8_sg U60351 ( .A(n33652), .X(n68230) );
  nand_x4_sg U60352 ( .A(n33396), .B(n33653), .X(n33652) );
  inv_x4_sg U60353 ( .A(n46935), .X(n57096) );
  inv_x8_sg U60354 ( .A(n57096), .X(n57097) );
  inv_x8_sg U60355 ( .A(n57097), .X(n68576) );
  nor_x8_sg U60356 ( .A(n57298), .B(n57097), .X(n23308) );
  nand_x1_sg U60357 ( .A(n26044), .B(n57114), .X(n26045) );
  inv_x1_sg U60358 ( .A(n68509), .X(n58643) );
  inv_x1_sg U60359 ( .A(n68420), .X(n58605) );
  nand_x1_sg U60360 ( .A(n57107), .B(n51015), .X(n26293) );
  nand_x1_sg U60361 ( .A(n57107), .B(n51021), .X(n26279) );
  nand_x1_sg U60362 ( .A(n57107), .B(n51005), .X(n26315) );
  nand_x1_sg U60363 ( .A(n57109), .B(n51011), .X(n26314) );
  nand_x1_sg U60364 ( .A(n26092), .B(n51023), .X(n26277) );
  nand_x1_sg U60365 ( .A(n57106), .B(n51007), .X(n26313) );
  nand_x1_sg U60366 ( .A(n57111), .B(n51017), .X(n26294) );
  inv_x1_sg U60367 ( .A(n47355), .X(n57955) );
  nand_x1_sg U60368 ( .A(n57111), .B(n51009), .X(n26316) );
  nand_x2_sg U60369 ( .A(n56964), .B(n56966), .X(n32115) );
  nand_x2_sg U60370 ( .A(n56948), .B(n56950), .X(n32560) );
  nand_x2_sg U60371 ( .A(n56952), .B(n56954), .X(n32104) );
  nand_x2_sg U60372 ( .A(n56956), .B(n56958), .X(n32107) );
  nand_x2_sg U60373 ( .A(n56960), .B(n56962), .X(n32112) );
  nand_x2_sg U60374 ( .A(n56936), .B(n56938), .X(n32549) );
  nand_x2_sg U60375 ( .A(n56940), .B(n56942), .X(n32552) );
  nand_x2_sg U60376 ( .A(n56944), .B(n56946), .X(n32557) );
  nand_x1_sg U60377 ( .A(n35572), .B(n35573), .X(n44136) );
  nand_x1_sg U60378 ( .A(n35570), .B(n35571), .X(n44135) );
  nand_x1_sg U60379 ( .A(n35578), .B(n35579), .X(n44139) );
  nand_x1_sg U60380 ( .A(n35576), .B(n35577), .X(n44138) );
  nand_x1_sg U60381 ( .A(n35609), .B(n35610), .X(n44154) );
  nand_x1_sg U60382 ( .A(n35607), .B(n35608), .X(n44153) );
  nand_x1_sg U60383 ( .A(n35615), .B(n35616), .X(n44157) );
  nand_x1_sg U60384 ( .A(n35613), .B(n35614), .X(n44156) );
  nand_x1_sg U60385 ( .A(n35597), .B(n35598), .X(n44148) );
  nand_x1_sg U60386 ( .A(n35595), .B(n35596), .X(n44147) );
  nand_x1_sg U60387 ( .A(n35601), .B(n35602), .X(n44150) );
  nand_x1_sg U60388 ( .A(n35531), .B(n35532), .X(n44118) );
  nand_x1_sg U60389 ( .A(n35529), .B(n35530), .X(n44117) );
  nand_x1_sg U60390 ( .A(n35538), .B(n35539), .X(n44121) );
  nand_x1_sg U60391 ( .A(n35536), .B(n35537), .X(n44120) );
  nand_x1_sg U60392 ( .A(n35517), .B(n35518), .X(n44112) );
  nand_x1_sg U60393 ( .A(n35515), .B(n35516), .X(n44111) );
  nand_x1_sg U60394 ( .A(n35524), .B(n35525), .X(n44115) );
  nand_x1_sg U60395 ( .A(n35522), .B(n35523), .X(n44114) );
  nand_x1_sg U60396 ( .A(n35560), .B(n35561), .X(n44130) );
  nand_x1_sg U60397 ( .A(n35558), .B(n35559), .X(n44129) );
  nand_x1_sg U60398 ( .A(n35545), .B(n35546), .X(n44124) );
  nand_x1_sg U60399 ( .A(n35543), .B(n35544), .X(n44123) );
  nand_x1_sg U60400 ( .A(n35553), .B(n35554), .X(n44127) );
  nand_x1_sg U60401 ( .A(n35535), .B(n35677), .X(n44190) );
  nand_x1_sg U60402 ( .A(n35528), .B(n35676), .X(n44189) );
  nand_x1_sg U60403 ( .A(n35521), .B(n35681), .X(n44193) );
  nand_x1_sg U60404 ( .A(n35513), .B(n35680), .X(n44192) );
  nand_x1_sg U60405 ( .A(n35588), .B(n35692), .X(n44199) );
  nand_x1_sg U60406 ( .A(n35557), .B(n35661), .X(n44181) );
  nand_x1_sg U60407 ( .A(n35549), .B(n35660), .X(n44180) );
  nand_x1_sg U60408 ( .A(n35542), .B(n35649), .X(n44174) );
  nand_x1_sg U60409 ( .A(n26095), .B(n53595), .X(n26134) );
  nand_x1_sg U60410 ( .A(n57107), .B(n53593), .X(n26133) );
  nand_x1_sg U60411 ( .A(n57111), .B(n53609), .X(n26094) );
  nand_x1_sg U60412 ( .A(n57107), .B(n53607), .X(n26093) );
  nand_x1_sg U60413 ( .A(n57111), .B(n53623), .X(n26226) );
  nand_x1_sg U60414 ( .A(n57107), .B(n53621), .X(n26225) );
  nand_x1_sg U60415 ( .A(n57111), .B(n53637), .X(n26192) );
  nand_x1_sg U60416 ( .A(n57107), .B(n53635), .X(n26191) );
  nand_x2_sg U60417 ( .A(n57975), .B(n68268), .X(n57981) );
  nand_x2_sg U60418 ( .A(n53663), .B(n57786), .X(n35535) );
  nand_x2_sg U60419 ( .A(n53661), .B(n57786), .X(n35528) );
  nand_x2_sg U60420 ( .A(n53659), .B(n57786), .X(n35521) );
  nand_x2_sg U60421 ( .A(n53657), .B(n57786), .X(n35513) );
  nand_x2_sg U60422 ( .A(n57786), .B(n53703), .X(n35609) );
  nand_x2_sg U60423 ( .A(n57786), .B(n53701), .X(n35607) );
  nand_x2_sg U60424 ( .A(n57786), .B(n53693), .X(n35595) );
  nand_x2_sg U60425 ( .A(n57786), .B(n53673), .X(n35560) );
  nand_x2_sg U60426 ( .A(n57786), .B(n53671), .X(n35558) );
  nand_x2_sg U60427 ( .A(n57786), .B(n53669), .X(n35545) );
  nand_x2_sg U60428 ( .A(n57786), .B(n53667), .X(n35543) );
  nand_x2_sg U60429 ( .A(n57786), .B(n53699), .X(n35615) );
  nand_x2_sg U60430 ( .A(n57786), .B(n53697), .X(n35613) );
  nand_x2_sg U60431 ( .A(n57786), .B(n53695), .X(n35597) );
  nand_x2_sg U60432 ( .A(n57786), .B(n53685), .X(n35538) );
  nand_x2_sg U60433 ( .A(n57786), .B(n53683), .X(n35536) );
  nand_x2_sg U60434 ( .A(n57786), .B(n53681), .X(n35517) );
  nand_x2_sg U60435 ( .A(n57786), .B(n53679), .X(n35515) );
  nand_x2_sg U60436 ( .A(n57786), .B(n53675), .X(n35522) );
  nand_x2_sg U60437 ( .A(n53653), .B(n57786), .X(n35557) );
  nand_x2_sg U60438 ( .A(n53651), .B(n57786), .X(n35549) );
  nand_x2_sg U60439 ( .A(n57786), .B(n53707), .X(n35578) );
  nand_x2_sg U60440 ( .A(n57786), .B(n53705), .X(n35576) );
  nand_x2_sg U60441 ( .A(n57786), .B(n53689), .X(n35531) );
  nand_x2_sg U60442 ( .A(n47297), .B(n53687), .X(n35529) );
  nand_x2_sg U60443 ( .A(n47297), .B(n53677), .X(n35524) );
  nand_x2_sg U60444 ( .A(n53649), .B(n57786), .X(n35542) );
  nand_x2_sg U60445 ( .A(n57786), .B(n53709), .X(n35570) );
  nand_x2_sg U60446 ( .A(n53655), .B(n57786), .X(n35588) );
  nand_x2_sg U60447 ( .A(n57786), .B(n53691), .X(n35601) );
  nand_x2_sg U60448 ( .A(n57786), .B(n53665), .X(n35553) );
  nand_x2_sg U60449 ( .A(n57786), .B(n53711), .X(n35572) );
  nand_x2_sg U60450 ( .A(n58329), .B(n58328), .X(n58375) );
  nand_x2_sg U60451 ( .A(n58324), .B(n58323), .X(n58372) );
  nand_x2_sg U60452 ( .A(n58319), .B(n58318), .X(n58371) );
  nand_x2_sg U60453 ( .A(n58304), .B(n58303), .X(n58368) );
  nand_x2_sg U60454 ( .A(n58299), .B(n58298), .X(n58367) );
  nand_x2_sg U60455 ( .A(n58294), .B(n58293), .X(n58366) );
  nand_x2_sg U60456 ( .A(n58279), .B(n58278), .X(n58363) );
  nand_x2_sg U60457 ( .A(n58274), .B(n58273), .X(n58362) );
  nand_x2_sg U60458 ( .A(n58259), .B(n58258), .X(n58359) );
  nand_x2_sg U60459 ( .A(n58254), .B(n58253), .X(n58358) );
  nand_x2_sg U60460 ( .A(n58249), .B(n58248), .X(n58357) );
  nand_x2_sg U60461 ( .A(n58234), .B(n58233), .X(n58354) );
  nand_x2_sg U60462 ( .A(n58229), .B(n58228), .X(n58353) );
  nand_x2_sg U60463 ( .A(n58224), .B(n58223), .X(n58351) );
  nand_x2_sg U60464 ( .A(n58219), .B(n58218), .X(n58350) );
  nand_x2_sg U60465 ( .A(n58204), .B(n58203), .X(n58347) );
  nand_x2_sg U60466 ( .A(n58199), .B(n58198), .X(n58346) );
  nand_x2_sg U60467 ( .A(n58194), .B(n58193), .X(n58345) );
  nand_x2_sg U60468 ( .A(n58179), .B(n58178), .X(n58342) );
  nand_x2_sg U60469 ( .A(n58174), .B(n58173), .X(n58341) );
  nand_x2_sg U60470 ( .A(n58159), .B(n58158), .X(n58338) );
  nand_x2_sg U60471 ( .A(n58154), .B(n58153), .X(n58337) );
  nand_x2_sg U60472 ( .A(n58149), .B(n58148), .X(n58336) );
  nand_x2_sg U60473 ( .A(n58134), .B(n58133), .X(n58333) );
  nand_x2_sg U60474 ( .A(n58314), .B(n58313), .X(n58370) );
  nand_x2_sg U60475 ( .A(n58309), .B(n58308), .X(n58369) );
  nand_x2_sg U60476 ( .A(n58289), .B(n58288), .X(n58365) );
  nand_x2_sg U60477 ( .A(n58284), .B(n58283), .X(n58364) );
  nand_x2_sg U60478 ( .A(n58269), .B(n58268), .X(n58361) );
  nand_x2_sg U60479 ( .A(n58264), .B(n58263), .X(n58360) );
  nand_x2_sg U60480 ( .A(n58244), .B(n58243), .X(n58356) );
  nand_x2_sg U60481 ( .A(n58239), .B(n58238), .X(n58355) );
  nand_x2_sg U60482 ( .A(n58214), .B(n58213), .X(n58349) );
  nand_x2_sg U60483 ( .A(n58209), .B(n58208), .X(n58348) );
  nand_x2_sg U60484 ( .A(n58189), .B(n58188), .X(n58344) );
  nand_x2_sg U60485 ( .A(n58184), .B(n58183), .X(n58343) );
  nand_x2_sg U60486 ( .A(n58169), .B(n58168), .X(n58340) );
  nand_x2_sg U60487 ( .A(n58164), .B(n58163), .X(n58339) );
  nand_x2_sg U60488 ( .A(n58144), .B(n58143), .X(n58335) );
  nand_x2_sg U60489 ( .A(n58139), .B(n58138), .X(n58334) );
  nand_x2_sg U60490 ( .A(n58124), .B(n58123), .X(n24383) );
  nand_x2_sg U60491 ( .A(n58119), .B(n58118), .X(n24388) );
  nand_x2_sg U60492 ( .A(n58116), .B(n58115), .X(n24393) );
  nand_x2_sg U60493 ( .A(n58112), .B(n58111), .X(n24398) );
  nand_x2_sg U60494 ( .A(n58108), .B(n58107), .X(n24403) );
  nand_x2_sg U60495 ( .A(n58105), .B(n58104), .X(n24408) );
  nand_x2_sg U60496 ( .A(n58102), .B(n58101), .X(n24413) );
  nand_x2_sg U60497 ( .A(n58099), .B(n58098), .X(n24418) );
  nand_x2_sg U60498 ( .A(n58095), .B(n58094), .X(n24423) );
  nand_x2_sg U60499 ( .A(n58091), .B(n58090), .X(n24428) );
  nand_x2_sg U60500 ( .A(n58088), .B(n58087), .X(n24433) );
  nand_x2_sg U60501 ( .A(n58085), .B(n58084), .X(n24438) );
  nand_x2_sg U60502 ( .A(n58081), .B(n58080), .X(n24443) );
  nand_x2_sg U60503 ( .A(n58077), .B(n58076), .X(n24448) );
  nand_x2_sg U60504 ( .A(n58074), .B(n58073), .X(n24453) );
  nand_x2_sg U60505 ( .A(n58071), .B(n58070), .X(n24458) );
  nand_x2_sg U60506 ( .A(n58068), .B(n58067), .X(n24463) );
  nand_x2_sg U60507 ( .A(n58064), .B(n58063), .X(n24468) );
  nand_x2_sg U60508 ( .A(n58060), .B(n58059), .X(n24473) );
  nand_x2_sg U60509 ( .A(n58057), .B(n58056), .X(n24489) );
  nand_x2_sg U60510 ( .A(n58054), .B(n58053), .X(n24495) );
  nand_x2_sg U60511 ( .A(n58049), .B(n58048), .X(n24500) );
  nand_x2_sg U60512 ( .A(n58046), .B(n58045), .X(n24505) );
  nand_x2_sg U60513 ( .A(n58042), .B(n58041), .X(n24510) );
  nand_x2_sg U60514 ( .A(n58038), .B(n58037), .X(n24515) );
  nand_x2_sg U60515 ( .A(n58035), .B(n58034), .X(n24520) );
  nand_x2_sg U60516 ( .A(n58032), .B(n58031), .X(n24525) );
  nand_x2_sg U60517 ( .A(n58029), .B(n58028), .X(n24530) );
  nand_x2_sg U60518 ( .A(n58025), .B(n58024), .X(n24535) );
  nand_x2_sg U60519 ( .A(n58021), .B(n58020), .X(n24540) );
  nand_x2_sg U60520 ( .A(n58018), .B(n58017), .X(n24545) );
  nand_x2_sg U60521 ( .A(n58015), .B(n58014), .X(n24550) );
  nand_x2_sg U60522 ( .A(n58011), .B(n58010), .X(n24555) );
  nand_x2_sg U60523 ( .A(n58007), .B(n58006), .X(n24560) );
  nand_x2_sg U60524 ( .A(n58004), .B(n58003), .X(n24565) );
  nand_x2_sg U60525 ( .A(n58001), .B(n58000), .X(n24570) );
  nand_x2_sg U60526 ( .A(n57998), .B(n57997), .X(n24575) );
  nand_x2_sg U60527 ( .A(n57994), .B(n57993), .X(n24580) );
  nand_x2_sg U60528 ( .A(n57990), .B(n57989), .X(n24585) );
  nand_x2_sg U60529 ( .A(n57986), .B(n57985), .X(n24601) );
  inv_x4_sg U60530 ( .A(n58480), .X(n57347) );
  nand_x1_sg U60531 ( .A(n57461), .B(n58616), .X(n57979) );
  inv_x2_sg U60532 ( .A(n68591), .X(n57451) );
  inv_x2_sg U60533 ( .A(n68591), .X(n57452) );
  inv_x4_sg U60534 ( .A(n57868), .X(n57867) );
  inv_x4_sg U60535 ( .A(n57976), .X(n57324) );
  inv_x4_sg U60536 ( .A(n57495), .X(n57494) );
  inv_x4_sg U60537 ( .A(n57479), .X(n57478) );
  inv_x4_sg U60538 ( .A(n57475), .X(n57474) );
  inv_x4_sg U60539 ( .A(n57491), .X(n57490) );
  inv_x4_sg U60540 ( .A(n58390), .X(n57501) );
  inv_x4_sg U60541 ( .A(n57987), .X(n57313) );
  inv_x4_sg U60542 ( .A(n58389), .X(n57498) );
  inv_x4_sg U60543 ( .A(n58391), .X(n57504) );
  nand_x4_sg U60544 ( .A(n57922), .B(n57926), .X(n58644) );
  nand_x4_sg U60545 ( .A(n57453), .B(n57917), .X(n58483) );
  nand_x4_sg U60546 ( .A(n58481), .B(n57917), .X(n58581) );
  nand_x4_sg U60547 ( .A(n57920), .B(n57100), .X(n58476) );
  nand_x1_sg U60548 ( .A(n67499), .B(n57345), .X(n22594) );
  nand_x1_sg U60549 ( .A(n57864), .B(n67499), .X(n22646) );
  nand_x2_sg U60550 ( .A(n57455), .B(n57923), .X(n57987) );
  nand_x2_sg U60551 ( .A(n57349), .B(n57100), .X(n58389) );
  nand_x2_sg U60552 ( .A(n57327), .B(n57100), .X(n58391) );
  inv_x4_sg U60553 ( .A(n57487), .X(n57486) );
  inv_x4_sg U60554 ( .A(n57483), .X(n57482) );
  nand_x1_sg U60555 ( .A(n57166), .B(n68379), .X(n33653) );
  nand_x1_sg U60556 ( .A(n57166), .B(n68385), .X(n33397) );
  nor_x1_sg U60557 ( .A(n31978), .B(n68575), .X(n31986) );
  nor_x1_sg U60558 ( .A(n31979), .B(n68570), .X(n31985) );
  nor_x1_sg U60559 ( .A(n32377), .B(n68397), .X(n32508) );
  nor_x1_sg U60560 ( .A(n32440), .B(n32378), .X(n32507) );
  nor_x1_sg U60561 ( .A(n32377), .B(n57303), .X(n32385) );
  nor_x1_sg U60562 ( .A(n32378), .B(n68388), .X(n32384) );
  nand_x4_sg U60563 ( .A(n32211), .B(n32212), .X(n31962) );
  nor_x1_sg U60564 ( .A(n68546), .B(n32295), .X(n32211) );
  nor_x1_sg U60565 ( .A(n58633), .B(n58632), .X(n32212) );
  nand_x4_sg U60566 ( .A(n32656), .B(n32657), .X(n32429) );
  nor_x1_sg U60567 ( .A(n68453), .B(n32740), .X(n32656) );
  nor_x1_sg U60568 ( .A(n58598), .B(n58597), .X(n32657) );
  nand_x2_sg U60569 ( .A(n31963), .B(n31964), .X(n31958) );
  nand_x2_sg U60570 ( .A(n68535), .B(n31960), .X(n31959) );
  nand_x2_sg U60571 ( .A(n32430), .B(n32431), .X(n32425) );
  nand_x2_sg U60572 ( .A(n68442), .B(n32427), .X(n32426) );
  nand_x2_sg U60573 ( .A(n31954), .B(n31955), .X(n31953) );
  nand_x1_sg U60574 ( .A(n68509), .B(n58655), .X(n31955) );
  nand_x2_sg U60575 ( .A(n32422), .B(n32423), .X(n32421) );
  nand_x1_sg U60576 ( .A(n68420), .B(n58655), .X(n32423) );
  nand_x1_sg U60577 ( .A(n68407), .B(n57349), .X(n58608) );
  nor_x1_sg U60578 ( .A(n57099), .B(n32433), .X(n58606) );
  nand_x1_sg U60579 ( .A(n68496), .B(n57349), .X(n58647) );
  nor_x1_sg U60580 ( .A(n57099), .B(n31966), .X(n58645) );
  inv_x4_sg U60581 ( .A(n57560), .X(n57559) );
  nor_x1_sg U60582 ( .A(n32407), .B(n32408), .X(n32395) );
  nor_x1_sg U60583 ( .A(n58621), .B(n58620), .X(n32396) );
  nor_x1_sg U60584 ( .A(n31939), .B(n31940), .X(n31927) );
  nor_x1_sg U60585 ( .A(n58659), .B(n58658), .X(n31928) );
  nor_x1_sg U60586 ( .A(n57100), .B(n68571), .X(n24265) );
  nand_x4_sg U60587 ( .A(n24370), .B(n23416), .X(n24369) );
  nor_x1_sg U60588 ( .A(n57918), .B(n68389), .X(n24370) );
  nor_x1_sg U60589 ( .A(n23416), .B(n24158), .X(n24157) );
  nand_x1_sg U60590 ( .A(n23416), .B(n68389), .X(n24375) );
  nor_x1_sg U60591 ( .A(n68397), .B(n68389), .X(n22596) );
  nand_x2_sg U60592 ( .A(n23413), .B(n23414), .X(n23412) );
  nand_x1_sg U60593 ( .A(n29339), .B(n57917), .X(n23413) );
  nand_x1_sg U60594 ( .A(n58616), .B(n58431), .X(n23414) );
  nand_x2_sg U60595 ( .A(n24155), .B(n24156), .X(n24154) );
  nand_x1_sg U60596 ( .A(n24159), .B(n57920), .X(n24155) );
  nand_x1_sg U60597 ( .A(n26047), .B(n67537), .X(n26046) );
  nor_x1_sg U60598 ( .A(n57100), .B(n68389), .X(n24374) );
  nand_x1_sg U60599 ( .A(n24374), .B(n23416), .X(n24373) );
  nor_x1_sg U60600 ( .A(n57865), .B(n68572), .X(n22420) );
  nor_x1_sg U60601 ( .A(n57865), .B(n68390), .X(n22444) );
  nand_x1_sg U60602 ( .A(n68397), .B(n68390), .X(n23680) );
  inv_x4_sg U60603 ( .A(n57471), .X(n57470) );
  inv_x4_sg U60604 ( .A(n57467), .X(n57466) );
  nor_x1_sg U60605 ( .A(n31982), .B(n46871), .X(n31980) );
  nor_x1_sg U60606 ( .A(n68570), .B(n31974), .X(n31983) );
  nor_x1_sg U60607 ( .A(n32381), .B(n32382), .X(n32379) );
  nor_x1_sg U60608 ( .A(n32438), .B(n32439), .X(n32434) );
  nand_x1_sg U60609 ( .A(n31994), .B(n68487), .X(n31993) );
  nand_x1_sg U60610 ( .A(n68398), .B(n31994), .X(n32436) );
  nand_x2_sg U60611 ( .A(n57856), .B(n32922), .X(n32921) );
  nand_x2_sg U60612 ( .A(n57856), .B(n32877), .X(n32876) );
  nand_x2_sg U60613 ( .A(n58631), .B(n58630), .X(n58632) );
  nand_x2_sg U60614 ( .A(n58596), .B(n58630), .X(n58597) );
  nand_x2_sg U60615 ( .A(n32296), .B(n32297), .X(n32295) );
  nand_x2_sg U60616 ( .A(n32741), .B(n32742), .X(n32740) );
  nor_x1_sg U60617 ( .A(n32521), .B(n32522), .X(n32520) );
  nor_x1_sg U60618 ( .A(n32076), .B(n32077), .X(n32075) );
  nand_x2_sg U60619 ( .A(n32085), .B(n32086), .X(n32084) );
  nand_x2_sg U60620 ( .A(n32530), .B(n32531), .X(n32529) );
  nand_x2_sg U60621 ( .A(n32080), .B(n32081), .X(n32074) );
  nand_x1_sg U60622 ( .A(n47319), .B(n61902), .X(n32081) );
  nand_x2_sg U60623 ( .A(n32525), .B(n32526), .X(n32519) );
  nand_x1_sg U60624 ( .A(n47300), .B(n61902), .X(n32526) );
  nand_x1_sg U60625 ( .A(n29336), .B(n68575), .X(n31988) );
  nand_x1_sg U60626 ( .A(n57298), .B(n68571), .X(n31989) );
  nand_x2_sg U60627 ( .A(n32387), .B(n32388), .X(n32386) );
  nand_x1_sg U60628 ( .A(n29338), .B(n57303), .X(n32387) );
  nand_x1_sg U60629 ( .A(n58643), .B(n58655), .X(n31963) );
  nand_x1_sg U60630 ( .A(n58605), .B(n58655), .X(n32430) );
  inv_x4_sg U60631 ( .A(n57885), .X(n57884) );
  nor_x1_sg U60632 ( .A(n57099), .B(n58634), .X(n58635) );
  nor_x1_sg U60633 ( .A(n57099), .B(n58599), .X(n58600) );
  inv_x4_sg U60634 ( .A(n39839), .X(n57561) );
  nand_x1_sg U60635 ( .A(n57324), .B(n61910), .X(n57977) );
  nand_x4_sg U60636 ( .A(n32539), .B(n32540), .X(n32513) );
  nor_x1_sg U60637 ( .A(n32579), .B(n32580), .X(n32539) );
  nor_x1_sg U60638 ( .A(n58604), .B(n58603), .X(n32540) );
  nand_x4_sg U60639 ( .A(n32094), .B(n32095), .X(n32067) );
  nor_x1_sg U60640 ( .A(n32134), .B(n32135), .X(n32094) );
  nor_x1_sg U60641 ( .A(n58642), .B(n58641), .X(n32095) );
  nor_x1_sg U60642 ( .A(n57099), .B(n58622), .X(n58623) );
  nor_x1_sg U60643 ( .A(n57099), .B(n58588), .X(n58589) );
  nand_x1_sg U60644 ( .A(n61910), .B(n58644), .X(n57975) );
  nand_x1_sg U60645 ( .A(n61910), .B(n57980), .X(n57983) );
  nand_x2_sg U60646 ( .A(n68534), .B(n31932), .X(n31931) );
  nand_x2_sg U60647 ( .A(n68395), .B(n32400), .X(n32399) );
  nand_x1_sg U60648 ( .A(n57924), .B(n61909), .X(n57973) );
  nand_x1_sg U60649 ( .A(n61910), .B(n57972), .X(n57974) );
  inv_x4_sg U60650 ( .A(n38415), .X(n57529) );
  nand_x2_sg U60651 ( .A(n68393), .B(n32410), .X(n32409) );
  nand_x2_sg U60652 ( .A(n68524), .B(n31942), .X(n31941) );
  nand_x2_sg U60653 ( .A(n68515), .B(n31946), .X(n31945) );
  nand_x2_sg U60654 ( .A(n68392), .B(n32414), .X(n32413) );
  nor_x1_sg U60655 ( .A(n58618), .B(n57928), .X(n58619) );
  nand_x2_sg U60656 ( .A(n57454), .B(n32437), .X(n58618) );
  nor_x1_sg U60657 ( .A(n58653), .B(n57926), .X(n58654) );
  nand_x2_sg U60658 ( .A(n57455), .B(n31995), .X(n58653) );
  nand_x2_sg U60659 ( .A(n68394), .B(n32404), .X(n32403) );
  nand_x2_sg U60660 ( .A(n68529), .B(n31936), .X(n31935) );
  nor_x1_sg U60661 ( .A(n32401), .B(n57306), .X(n32402) );
  nor_x1_sg U60662 ( .A(n31933), .B(n57300), .X(n31934) );
  nor_x1_sg U60663 ( .A(n32411), .B(n57306), .X(n32412) );
  nor_x1_sg U60664 ( .A(n31943), .B(n57300), .X(n31944) );
  nor_x1_sg U60665 ( .A(n32405), .B(n57306), .X(n32406) );
  nor_x1_sg U60666 ( .A(n31937), .B(n57300), .X(n31938) );
  nor_x1_sg U60667 ( .A(n31947), .B(n57300), .X(n31948) );
  nor_x1_sg U60668 ( .A(n32415), .B(n57306), .X(n32416) );
  nand_x1_sg U60669 ( .A(n22467), .B(n57345), .X(n22568) );
  nand_x1_sg U60670 ( .A(n57864), .B(n22467), .X(n22619) );
  nand_x2_sg U60671 ( .A(n24045), .B(n24046), .X(n24044) );
  nand_x1_sg U60672 ( .A(n24050), .B(n57920), .X(n24045) );
  nor_x1_sg U60673 ( .A(n67086), .B(n22623), .X(n22622) );
  nor_x1_sg U60674 ( .A(n67086), .B(n22650), .X(n22649) );
  nor_x1_sg U60675 ( .A(n57298), .B(n67086), .X(n22698) );
  nor_x1_sg U60676 ( .A(n57304), .B(n67086), .X(n22745) );
  nor_x1_sg U60677 ( .A(n57298), .B(n22572), .X(n22571) );
  nor_x1_sg U60678 ( .A(n57304), .B(n22572), .X(n22597) );
  nand_x2_sg U60679 ( .A(n24780), .B(n24781), .X(n24779) );
  nand_x1_sg U60680 ( .A(n67523), .B(n57296), .X(n24781) );
  nand_x2_sg U60681 ( .A(n24686), .B(n24687), .X(n24685) );
  nand_x1_sg U60682 ( .A(n67101), .B(n57296), .X(n24687) );
  nor_x1_sg U60683 ( .A(n23416), .B(n23417), .X(n23415) );
  nor_x1_sg U60684 ( .A(n67116), .B(n22446), .X(\shifter_0/n12505 ) );
  nor_x1_sg U60685 ( .A(n67115), .B(n22446), .X(\shifter_0/n12501 ) );
  nor_x1_sg U60686 ( .A(n67114), .B(n22446), .X(\shifter_0/n12497 ) );
  nor_x1_sg U60687 ( .A(n67113), .B(n22446), .X(\shifter_0/n12493 ) );
  nor_x1_sg U60688 ( .A(n67112), .B(n22446), .X(\shifter_0/n12489 ) );
  nor_x1_sg U60689 ( .A(n67111), .B(n22446), .X(\shifter_0/n12485 ) );
  nor_x1_sg U60690 ( .A(n67110), .B(n22446), .X(\shifter_0/n12481 ) );
  nor_x1_sg U60691 ( .A(n67109), .B(n22446), .X(\shifter_0/n12477 ) );
  nor_x1_sg U60692 ( .A(n67108), .B(n22446), .X(\shifter_0/n12473 ) );
  nor_x1_sg U60693 ( .A(n67107), .B(n22446), .X(\shifter_0/n12469 ) );
  nor_x1_sg U60694 ( .A(n67106), .B(n22446), .X(\shifter_0/n12465 ) );
  nor_x1_sg U60695 ( .A(n67105), .B(n22446), .X(\shifter_0/n12461 ) );
  nor_x1_sg U60696 ( .A(n67104), .B(n22446), .X(\shifter_0/n12457 ) );
  nor_x1_sg U60697 ( .A(n67136), .B(n22498), .X(\shifter_0/n12345 ) );
  nor_x1_sg U60698 ( .A(n67135), .B(n22498), .X(\shifter_0/n12341 ) );
  nor_x1_sg U60699 ( .A(n67134), .B(n22498), .X(\shifter_0/n12337 ) );
  nor_x1_sg U60700 ( .A(n67133), .B(n22498), .X(\shifter_0/n12333 ) );
  nor_x1_sg U60701 ( .A(n67132), .B(n22498), .X(\shifter_0/n12329 ) );
  nor_x1_sg U60702 ( .A(n67131), .B(n22498), .X(\shifter_0/n12325 ) );
  nor_x1_sg U60703 ( .A(n67130), .B(n22498), .X(\shifter_0/n12321 ) );
  nor_x1_sg U60704 ( .A(n67129), .B(n22498), .X(\shifter_0/n12317 ) );
  nor_x1_sg U60705 ( .A(n67128), .B(n22498), .X(\shifter_0/n12313 ) );
  nor_x1_sg U60706 ( .A(n67127), .B(n22498), .X(\shifter_0/n12309 ) );
  nor_x1_sg U60707 ( .A(n67126), .B(n22498), .X(\shifter_0/n12305 ) );
  nor_x1_sg U60708 ( .A(n67125), .B(n22498), .X(\shifter_0/n12301 ) );
  nor_x1_sg U60709 ( .A(n67124), .B(n22498), .X(\shifter_0/n12297 ) );
  nor_x1_sg U60710 ( .A(n67329), .B(n22473), .X(\shifter_0/n12425 ) );
  nor_x1_sg U60711 ( .A(n67328), .B(n22473), .X(\shifter_0/n12421 ) );
  nor_x1_sg U60712 ( .A(n67327), .B(n22473), .X(\shifter_0/n12417 ) );
  nor_x1_sg U60713 ( .A(n67326), .B(n22473), .X(\shifter_0/n12413 ) );
  nor_x1_sg U60714 ( .A(n67325), .B(n22473), .X(\shifter_0/n12409 ) );
  nor_x1_sg U60715 ( .A(n67324), .B(n22473), .X(\shifter_0/n12405 ) );
  nor_x1_sg U60716 ( .A(n67323), .B(n22473), .X(\shifter_0/n12401 ) );
  nor_x1_sg U60717 ( .A(n67322), .B(n22473), .X(\shifter_0/n12397 ) );
  nor_x1_sg U60718 ( .A(n67321), .B(n22473), .X(\shifter_0/n12393 ) );
  nor_x1_sg U60719 ( .A(n67320), .B(n22473), .X(\shifter_0/n12389 ) );
  nor_x1_sg U60720 ( .A(n67319), .B(n22473), .X(\shifter_0/n12385 ) );
  nor_x1_sg U60721 ( .A(n67318), .B(n22473), .X(\shifter_0/n12381 ) );
  nor_x1_sg U60722 ( .A(n67317), .B(n22473), .X(\shifter_0/n12377 ) );
  nor_x1_sg U60723 ( .A(n67349), .B(n22523), .X(\shifter_0/n12265 ) );
  nor_x1_sg U60724 ( .A(n67348), .B(n22523), .X(\shifter_0/n12261 ) );
  nor_x1_sg U60725 ( .A(n67347), .B(n22523), .X(\shifter_0/n12257 ) );
  nor_x1_sg U60726 ( .A(n67346), .B(n22523), .X(\shifter_0/n12253 ) );
  nor_x1_sg U60727 ( .A(n67345), .B(n22523), .X(\shifter_0/n12249 ) );
  nor_x1_sg U60728 ( .A(n67344), .B(n22523), .X(\shifter_0/n12245 ) );
  nor_x1_sg U60729 ( .A(n67343), .B(n22523), .X(\shifter_0/n12241 ) );
  nor_x1_sg U60730 ( .A(n67342), .B(n22523), .X(\shifter_0/n12237 ) );
  nor_x1_sg U60731 ( .A(n67341), .B(n22523), .X(\shifter_0/n12233 ) );
  nor_x1_sg U60732 ( .A(n67340), .B(n22523), .X(\shifter_0/n12229 ) );
  nor_x1_sg U60733 ( .A(n67339), .B(n22523), .X(\shifter_0/n12225 ) );
  nor_x1_sg U60734 ( .A(n67338), .B(n22523), .X(\shifter_0/n12221 ) );
  nor_x1_sg U60735 ( .A(n67337), .B(n22523), .X(\shifter_0/n12217 ) );
  nor_x1_sg U60736 ( .A(n61867), .B(n22396), .X(\shifter_0/n12665 ) );
  nor_x1_sg U60737 ( .A(n61868), .B(n22396), .X(\shifter_0/n12661 ) );
  nor_x1_sg U60738 ( .A(n61869), .B(n22396), .X(\shifter_0/n12657 ) );
  nor_x1_sg U60739 ( .A(n61870), .B(n22396), .X(\shifter_0/n12653 ) );
  nor_x1_sg U60740 ( .A(n61871), .B(n22396), .X(\shifter_0/n12649 ) );
  nor_x1_sg U60741 ( .A(n61872), .B(n22396), .X(\shifter_0/n12645 ) );
  nor_x1_sg U60742 ( .A(n61873), .B(n22396), .X(\shifter_0/n12641 ) );
  nor_x1_sg U60743 ( .A(n61874), .B(n22396), .X(\shifter_0/n12637 ) );
  nor_x1_sg U60744 ( .A(n61875), .B(n22396), .X(\shifter_0/n12633 ) );
  nor_x1_sg U60745 ( .A(n61876), .B(n22396), .X(\shifter_0/n12629 ) );
  nor_x1_sg U60746 ( .A(n61877), .B(n22396), .X(\shifter_0/n12625 ) );
  nor_x1_sg U60747 ( .A(n61878), .B(n22396), .X(\shifter_0/n12621 ) );
  nor_x1_sg U60748 ( .A(n61879), .B(n22396), .X(\shifter_0/n12617 ) );
  nor_x1_sg U60749 ( .A(n61887), .B(n22421), .X(\shifter_0/n12585 ) );
  nor_x1_sg U60750 ( .A(n61888), .B(n22421), .X(\shifter_0/n12581 ) );
  nor_x1_sg U60751 ( .A(n61889), .B(n22421), .X(\shifter_0/n12577 ) );
  nor_x1_sg U60752 ( .A(n61890), .B(n22421), .X(\shifter_0/n12573 ) );
  nor_x1_sg U60753 ( .A(n61891), .B(n22421), .X(\shifter_0/n12569 ) );
  nor_x1_sg U60754 ( .A(n61892), .B(n22421), .X(\shifter_0/n12565 ) );
  nor_x1_sg U60755 ( .A(n61893), .B(n22421), .X(\shifter_0/n12561 ) );
  nor_x1_sg U60756 ( .A(n61894), .B(n22421), .X(\shifter_0/n12557 ) );
  nor_x1_sg U60757 ( .A(n61895), .B(n22421), .X(\shifter_0/n12553 ) );
  nor_x1_sg U60758 ( .A(n61896), .B(n22421), .X(\shifter_0/n12549 ) );
  nor_x1_sg U60759 ( .A(n61897), .B(n22421), .X(\shifter_0/n12545 ) );
  nor_x1_sg U60760 ( .A(n61898), .B(n22421), .X(\shifter_0/n12541 ) );
  nor_x1_sg U60761 ( .A(n61899), .B(n22421), .X(\shifter_0/n12537 ) );
  nor_x1_sg U60762 ( .A(n67121), .B(n22446), .X(\shifter_0/n12525 ) );
  nor_x1_sg U60763 ( .A(n67120), .B(n22446), .X(\shifter_0/n12521 ) );
  nor_x1_sg U60764 ( .A(n67119), .B(n22446), .X(\shifter_0/n12517 ) );
  nor_x1_sg U60765 ( .A(n67118), .B(n22446), .X(\shifter_0/n12513 ) );
  nor_x1_sg U60766 ( .A(n67117), .B(n22446), .X(\shifter_0/n12509 ) );
  nor_x1_sg U60767 ( .A(n67141), .B(n22498), .X(\shifter_0/n12365 ) );
  nor_x1_sg U60768 ( .A(n67140), .B(n22498), .X(\shifter_0/n12361 ) );
  nor_x1_sg U60769 ( .A(n67139), .B(n22498), .X(\shifter_0/n12357 ) );
  nor_x1_sg U60770 ( .A(n67138), .B(n22498), .X(\shifter_0/n12353 ) );
  nor_x1_sg U60771 ( .A(n67137), .B(n22498), .X(\shifter_0/n12349 ) );
  nor_x1_sg U60772 ( .A(n57510), .B(n67156), .X(\shifter_0/n12185 ) );
  nor_x1_sg U60773 ( .A(n57510), .B(n67155), .X(\shifter_0/n12181 ) );
  nor_x1_sg U60774 ( .A(n57510), .B(n67154), .X(\shifter_0/n12177 ) );
  nor_x1_sg U60775 ( .A(n57510), .B(n67153), .X(\shifter_0/n12173 ) );
  nor_x1_sg U60776 ( .A(n57510), .B(n67152), .X(\shifter_0/n12169 ) );
  nor_x1_sg U60777 ( .A(n57510), .B(n67151), .X(\shifter_0/n12165 ) );
  nor_x1_sg U60778 ( .A(n57510), .B(n67150), .X(\shifter_0/n12161 ) );
  nor_x1_sg U60779 ( .A(n57510), .B(n67149), .X(\shifter_0/n12157 ) );
  nor_x1_sg U60780 ( .A(n57510), .B(n67148), .X(\shifter_0/n12153 ) );
  nor_x1_sg U60781 ( .A(n57507), .B(n67176), .X(\shifter_0/n12025 ) );
  nor_x1_sg U60782 ( .A(n57507), .B(n67175), .X(\shifter_0/n12021 ) );
  nor_x1_sg U60783 ( .A(n57507), .B(n67174), .X(\shifter_0/n12017 ) );
  nor_x1_sg U60784 ( .A(n57507), .B(n67173), .X(\shifter_0/n12013 ) );
  nor_x1_sg U60785 ( .A(n57507), .B(n67172), .X(\shifter_0/n12009 ) );
  nor_x1_sg U60786 ( .A(n57507), .B(n67171), .X(\shifter_0/n12005 ) );
  nor_x1_sg U60787 ( .A(n57507), .B(n67170), .X(\shifter_0/n12001 ) );
  nor_x1_sg U60788 ( .A(n57507), .B(n67169), .X(\shifter_0/n11997 ) );
  nor_x1_sg U60789 ( .A(n57507), .B(n67168), .X(\shifter_0/n11993 ) );
  nor_x1_sg U60790 ( .A(n57516), .B(n67369), .X(\shifter_0/n12105 ) );
  nor_x1_sg U60791 ( .A(n57516), .B(n67368), .X(\shifter_0/n12101 ) );
  nor_x1_sg U60792 ( .A(n57516), .B(n67367), .X(\shifter_0/n12097 ) );
  nor_x1_sg U60793 ( .A(n57516), .B(n67366), .X(\shifter_0/n12093 ) );
  nor_x1_sg U60794 ( .A(n57516), .B(n67365), .X(\shifter_0/n12089 ) );
  nor_x1_sg U60795 ( .A(n57516), .B(n67364), .X(\shifter_0/n12085 ) );
  nor_x1_sg U60796 ( .A(n57516), .B(n67363), .X(\shifter_0/n12081 ) );
  nor_x1_sg U60797 ( .A(n57516), .B(n67362), .X(\shifter_0/n12077 ) );
  nor_x1_sg U60798 ( .A(n57516), .B(n67361), .X(\shifter_0/n12073 ) );
  nor_x1_sg U60799 ( .A(n57513), .B(n67389), .X(\shifter_0/n11945 ) );
  nor_x1_sg U60800 ( .A(n57513), .B(n67388), .X(\shifter_0/n11941 ) );
  nor_x1_sg U60801 ( .A(n57513), .B(n67387), .X(\shifter_0/n11937 ) );
  nor_x1_sg U60802 ( .A(n57513), .B(n67386), .X(\shifter_0/n11933 ) );
  nor_x1_sg U60803 ( .A(n57513), .B(n67385), .X(\shifter_0/n11929 ) );
  nor_x1_sg U60804 ( .A(n57513), .B(n67384), .X(\shifter_0/n11925 ) );
  nor_x1_sg U60805 ( .A(n57513), .B(n67383), .X(\shifter_0/n11921 ) );
  nor_x1_sg U60806 ( .A(n57513), .B(n67382), .X(\shifter_0/n11917 ) );
  nor_x1_sg U60807 ( .A(n57513), .B(n67381), .X(\shifter_0/n11913 ) );
  nor_x1_sg U60808 ( .A(n57510), .B(n67147), .X(\shifter_0/n12149 ) );
  nor_x1_sg U60809 ( .A(n57510), .B(n67146), .X(\shifter_0/n12145 ) );
  nor_x1_sg U60810 ( .A(n57510), .B(n67145), .X(\shifter_0/n12141 ) );
  nor_x1_sg U60811 ( .A(n57510), .B(n67144), .X(\shifter_0/n12137 ) );
  nor_x1_sg U60812 ( .A(n57507), .B(n67167), .X(\shifter_0/n11989 ) );
  nor_x1_sg U60813 ( .A(n57507), .B(n67166), .X(\shifter_0/n11985 ) );
  nor_x1_sg U60814 ( .A(n57507), .B(n67165), .X(\shifter_0/n11981 ) );
  nor_x1_sg U60815 ( .A(n57507), .B(n67164), .X(\shifter_0/n11977 ) );
  nor_x1_sg U60816 ( .A(n57516), .B(n67360), .X(\shifter_0/n12069 ) );
  nor_x1_sg U60817 ( .A(n57516), .B(n67359), .X(\shifter_0/n12065 ) );
  nor_x1_sg U60818 ( .A(n57516), .B(n67358), .X(\shifter_0/n12061 ) );
  nor_x1_sg U60819 ( .A(n57516), .B(n67357), .X(\shifter_0/n12057 ) );
  nor_x1_sg U60820 ( .A(n57513), .B(n67380), .X(\shifter_0/n11909 ) );
  nor_x1_sg U60821 ( .A(n57513), .B(n67379), .X(\shifter_0/n11905 ) );
  nor_x1_sg U60822 ( .A(n57513), .B(n67378), .X(\shifter_0/n11901 ) );
  nor_x1_sg U60823 ( .A(n57513), .B(n67377), .X(\shifter_0/n11897 ) );
  nor_x1_sg U60824 ( .A(n67334), .B(n22473), .X(\shifter_0/n12445 ) );
  nor_x1_sg U60825 ( .A(n67333), .B(n22473), .X(\shifter_0/n12441 ) );
  nor_x1_sg U60826 ( .A(n67332), .B(n22473), .X(\shifter_0/n12437 ) );
  nor_x1_sg U60827 ( .A(n67331), .B(n22473), .X(\shifter_0/n12433 ) );
  nor_x1_sg U60828 ( .A(n67330), .B(n22473), .X(\shifter_0/n12429 ) );
  nor_x1_sg U60829 ( .A(n67354), .B(n22523), .X(\shifter_0/n12285 ) );
  nor_x1_sg U60830 ( .A(n67353), .B(n22523), .X(\shifter_0/n12281 ) );
  nor_x1_sg U60831 ( .A(n67352), .B(n22523), .X(\shifter_0/n12277 ) );
  nor_x1_sg U60832 ( .A(n67351), .B(n22523), .X(\shifter_0/n12273 ) );
  nor_x1_sg U60833 ( .A(n67350), .B(n22523), .X(\shifter_0/n12269 ) );
  nor_x1_sg U60834 ( .A(n61862), .B(n22396), .X(\shifter_0/n12685 ) );
  nor_x1_sg U60835 ( .A(n61863), .B(n22396), .X(\shifter_0/n12681 ) );
  nor_x1_sg U60836 ( .A(n61864), .B(n22396), .X(\shifter_0/n12677 ) );
  nor_x1_sg U60837 ( .A(n61865), .B(n22396), .X(\shifter_0/n12673 ) );
  nor_x1_sg U60838 ( .A(n61866), .B(n22396), .X(\shifter_0/n12669 ) );
  nor_x1_sg U60839 ( .A(n61882), .B(n22421), .X(\shifter_0/n12605 ) );
  nor_x1_sg U60840 ( .A(n61883), .B(n22421), .X(\shifter_0/n12601 ) );
  nor_x1_sg U60841 ( .A(n61884), .B(n22421), .X(\shifter_0/n12597 ) );
  nor_x1_sg U60842 ( .A(n61885), .B(n22421), .X(\shifter_0/n12593 ) );
  nor_x1_sg U60843 ( .A(n61886), .B(n22421), .X(\shifter_0/n12589 ) );
  nor_x1_sg U60844 ( .A(n57128), .B(n24378), .X(\shifter_0/n10765 ) );
  nor_x1_sg U60845 ( .A(n57128), .B(n24384), .X(\shifter_0/n10761 ) );
  nor_x1_sg U60846 ( .A(n57128), .B(n24389), .X(\shifter_0/n10757 ) );
  nor_x1_sg U60847 ( .A(n57128), .B(n24394), .X(\shifter_0/n10753 ) );
  nor_x1_sg U60848 ( .A(n57128), .B(n24399), .X(\shifter_0/n10749 ) );
  nor_x1_sg U60849 ( .A(n57128), .B(n24404), .X(\shifter_0/n10745 ) );
  nor_x1_sg U60850 ( .A(n57128), .B(n24409), .X(\shifter_0/n10741 ) );
  nor_x1_sg U60851 ( .A(n57128), .B(n24414), .X(\shifter_0/n10737 ) );
  nor_x1_sg U60852 ( .A(n57128), .B(n24419), .X(\shifter_0/n10733 ) );
  nor_x1_sg U60853 ( .A(n57128), .B(n24424), .X(\shifter_0/n10729 ) );
  nor_x1_sg U60854 ( .A(n57128), .B(n24429), .X(\shifter_0/n10725 ) );
  nor_x1_sg U60855 ( .A(n57128), .B(n24434), .X(\shifter_0/n10721 ) );
  nor_x1_sg U60856 ( .A(n57128), .B(n24439), .X(\shifter_0/n10717 ) );
  nor_x1_sg U60857 ( .A(n57128), .B(n24444), .X(\shifter_0/n10713 ) );
  nor_x1_sg U60858 ( .A(n57128), .B(n24449), .X(\shifter_0/n10709 ) );
  nor_x1_sg U60859 ( .A(n57128), .B(n24454), .X(\shifter_0/n10705 ) );
  nor_x1_sg U60860 ( .A(n57128), .B(n24459), .X(\shifter_0/n10701 ) );
  nor_x1_sg U60861 ( .A(n57128), .B(n24464), .X(\shifter_0/n10697 ) );
  nor_x1_sg U60862 ( .A(n57128), .B(n24469), .X(\shifter_0/n10693 ) );
  nor_x1_sg U60863 ( .A(n57128), .B(n24474), .X(\shifter_0/n10689 ) );
  nor_x1_sg U60864 ( .A(n57125), .B(n24490), .X(\shifter_0/n10685 ) );
  nor_x1_sg U60865 ( .A(n57125), .B(n24496), .X(\shifter_0/n10681 ) );
  nor_x1_sg U60866 ( .A(n57125), .B(n24501), .X(\shifter_0/n10677 ) );
  nor_x1_sg U60867 ( .A(n57125), .B(n24506), .X(\shifter_0/n10673 ) );
  nor_x1_sg U60868 ( .A(n57125), .B(n24511), .X(\shifter_0/n10669 ) );
  nor_x1_sg U60869 ( .A(n57125), .B(n24516), .X(\shifter_0/n10665 ) );
  nor_x1_sg U60870 ( .A(n57125), .B(n24521), .X(\shifter_0/n10661 ) );
  nor_x1_sg U60871 ( .A(n57125), .B(n24526), .X(\shifter_0/n10657 ) );
  nor_x1_sg U60872 ( .A(n57125), .B(n24531), .X(\shifter_0/n10653 ) );
  nor_x1_sg U60873 ( .A(n57125), .B(n24536), .X(\shifter_0/n10649 ) );
  nor_x1_sg U60874 ( .A(n57125), .B(n24541), .X(\shifter_0/n10645 ) );
  nor_x1_sg U60875 ( .A(n57125), .B(n24546), .X(\shifter_0/n10641 ) );
  nor_x1_sg U60876 ( .A(n57125), .B(n24551), .X(\shifter_0/n10637 ) );
  nor_x1_sg U60877 ( .A(n57125), .B(n24556), .X(\shifter_0/n10633 ) );
  nor_x1_sg U60878 ( .A(n57125), .B(n24561), .X(\shifter_0/n10629 ) );
  nor_x1_sg U60879 ( .A(n57125), .B(n24566), .X(\shifter_0/n10625 ) );
  nor_x1_sg U60880 ( .A(n57125), .B(n24571), .X(\shifter_0/n10621 ) );
  nor_x1_sg U60881 ( .A(n57125), .B(n24576), .X(\shifter_0/n10617 ) );
  nor_x1_sg U60882 ( .A(n57125), .B(n24581), .X(\shifter_0/n10613 ) );
  nor_x1_sg U60883 ( .A(n57125), .B(n24586), .X(\shifter_0/n10609 ) );
  nor_x1_sg U60884 ( .A(n57118), .B(n24791), .X(\shifter_0/n10445 ) );
  nor_x1_sg U60885 ( .A(n57118), .B(n24830), .X(\shifter_0/n10441 ) );
  nor_x1_sg U60886 ( .A(n57118), .B(n24860), .X(\shifter_0/n10437 ) );
  nor_x1_sg U60887 ( .A(n57118), .B(n24890), .X(\shifter_0/n10433 ) );
  nor_x1_sg U60888 ( .A(n57118), .B(n24920), .X(\shifter_0/n10429 ) );
  nor_x1_sg U60889 ( .A(n57118), .B(n24950), .X(\shifter_0/n10425 ) );
  nor_x1_sg U60890 ( .A(n57118), .B(n24980), .X(\shifter_0/n10421 ) );
  nor_x1_sg U60891 ( .A(n57118), .B(n25010), .X(\shifter_0/n10417 ) );
  nor_x1_sg U60892 ( .A(n57118), .B(n25040), .X(\shifter_0/n10413 ) );
  nor_x1_sg U60893 ( .A(n57118), .B(n25070), .X(\shifter_0/n10409 ) );
  nor_x1_sg U60894 ( .A(n57118), .B(n25100), .X(\shifter_0/n10405 ) );
  nor_x1_sg U60895 ( .A(n57118), .B(n25130), .X(\shifter_0/n10401 ) );
  nor_x1_sg U60896 ( .A(n57118), .B(n25160), .X(\shifter_0/n10397 ) );
  nor_x1_sg U60897 ( .A(n57118), .B(n25190), .X(\shifter_0/n10393 ) );
  nor_x1_sg U60898 ( .A(n57118), .B(n25220), .X(\shifter_0/n10389 ) );
  nor_x1_sg U60899 ( .A(n57118), .B(n25250), .X(\shifter_0/n10385 ) );
  nor_x1_sg U60900 ( .A(n57118), .B(n25280), .X(\shifter_0/n10381 ) );
  nor_x1_sg U60901 ( .A(n57118), .B(n25310), .X(\shifter_0/n10377 ) );
  nor_x1_sg U60902 ( .A(n57118), .B(n25340), .X(\shifter_0/n10373 ) );
  nor_x1_sg U60903 ( .A(n57118), .B(n25370), .X(\shifter_0/n10369 ) );
  nor_x1_sg U60904 ( .A(n57116), .B(n25402), .X(\shifter_0/n10365 ) );
  nor_x1_sg U60905 ( .A(n57116), .B(n25432), .X(\shifter_0/n10361 ) );
  nor_x1_sg U60906 ( .A(n57116), .B(n25462), .X(\shifter_0/n10357 ) );
  nor_x1_sg U60907 ( .A(n57116), .B(n25492), .X(\shifter_0/n10353 ) );
  nor_x1_sg U60908 ( .A(n57116), .B(n25522), .X(\shifter_0/n10349 ) );
  nor_x1_sg U60909 ( .A(n57116), .B(n25552), .X(\shifter_0/n10345 ) );
  nor_x1_sg U60910 ( .A(n57116), .B(n25582), .X(\shifter_0/n10341 ) );
  nor_x1_sg U60911 ( .A(n57116), .B(n25612), .X(\shifter_0/n10337 ) );
  nor_x1_sg U60912 ( .A(n57116), .B(n25642), .X(\shifter_0/n10333 ) );
  nor_x1_sg U60913 ( .A(n57116), .B(n25672), .X(\shifter_0/n10329 ) );
  nor_x1_sg U60914 ( .A(n57116), .B(n25702), .X(\shifter_0/n10325 ) );
  nor_x1_sg U60915 ( .A(n57116), .B(n25732), .X(\shifter_0/n10321 ) );
  nor_x1_sg U60916 ( .A(n57116), .B(n25762), .X(\shifter_0/n10317 ) );
  nor_x1_sg U60917 ( .A(n57116), .B(n25792), .X(\shifter_0/n10313 ) );
  nor_x1_sg U60918 ( .A(n57116), .B(n25822), .X(\shifter_0/n10309 ) );
  nor_x1_sg U60919 ( .A(n57116), .B(n25852), .X(\shifter_0/n10305 ) );
  nor_x1_sg U60920 ( .A(n57116), .B(n25882), .X(\shifter_0/n10301 ) );
  nor_x1_sg U60921 ( .A(n57116), .B(n25912), .X(\shifter_0/n10297 ) );
  nor_x1_sg U60922 ( .A(n57116), .B(n25942), .X(\shifter_0/n10293 ) );
  nor_x1_sg U60923 ( .A(n57116), .B(n25972), .X(\shifter_0/n10289 ) );
  nor_x1_sg U60924 ( .A(n57510), .B(n67161), .X(\shifter_0/n12205 ) );
  nor_x1_sg U60925 ( .A(n57510), .B(n67160), .X(\shifter_0/n12201 ) );
  nor_x1_sg U60926 ( .A(n57510), .B(n67159), .X(\shifter_0/n12197 ) );
  nor_x1_sg U60927 ( .A(n57510), .B(n67158), .X(\shifter_0/n12193 ) );
  nor_x1_sg U60928 ( .A(n57510), .B(n67157), .X(\shifter_0/n12189 ) );
  nor_x1_sg U60929 ( .A(n67181), .B(n57507), .X(\shifter_0/n12045 ) );
  nor_x1_sg U60930 ( .A(n57507), .B(n67180), .X(\shifter_0/n12041 ) );
  nor_x1_sg U60931 ( .A(n57507), .B(n67179), .X(\shifter_0/n12037 ) );
  nor_x1_sg U60932 ( .A(n57507), .B(n67178), .X(\shifter_0/n12033 ) );
  nor_x1_sg U60933 ( .A(n57507), .B(n67177), .X(\shifter_0/n12029 ) );
  nor_x1_sg U60934 ( .A(n57516), .B(n67374), .X(\shifter_0/n12125 ) );
  nor_x1_sg U60935 ( .A(n57516), .B(n67373), .X(\shifter_0/n12121 ) );
  nor_x1_sg U60936 ( .A(n57516), .B(n67372), .X(\shifter_0/n12117 ) );
  nor_x1_sg U60937 ( .A(n57516), .B(n67371), .X(\shifter_0/n12113 ) );
  nor_x1_sg U60938 ( .A(n57516), .B(n67370), .X(\shifter_0/n12109 ) );
  nor_x1_sg U60939 ( .A(n67394), .B(n57513), .X(\shifter_0/n11965 ) );
  nor_x1_sg U60940 ( .A(n57513), .B(n67393), .X(\shifter_0/n11961 ) );
  nor_x1_sg U60941 ( .A(n57513), .B(n67392), .X(\shifter_0/n11957 ) );
  nor_x1_sg U60942 ( .A(n57513), .B(n67391), .X(\shifter_0/n11953 ) );
  nor_x1_sg U60943 ( .A(n57513), .B(n67390), .X(\shifter_0/n11949 ) );
  nor_x1_sg U60944 ( .A(n57113), .B(n26044), .X(\filter_0/n8284 ) );
  nor_x1_sg U60945 ( .A(n57113), .B(n26053), .X(\filter_0/n8276 ) );
  nor_x1_sg U60946 ( .A(n57113), .B(n26061), .X(\filter_0/n8264 ) );
  nor_x1_sg U60947 ( .A(n57113), .B(n26157), .X(\filter_0/n8252 ) );
  nor_x1_sg U60948 ( .A(n24567), .B(n24568), .X(\shifter_0/n10624 ) );
  nor_x1_sg U60949 ( .A(n24572), .B(n24573), .X(\shifter_0/n10620 ) );
  nor_x1_sg U60950 ( .A(n24577), .B(n24578), .X(\shifter_0/n10616 ) );
  nor_x1_sg U60951 ( .A(n24582), .B(n24583), .X(\shifter_0/n10612 ) );
  nor_x1_sg U60952 ( .A(n24587), .B(n24588), .X(\shifter_0/n10608 ) );
  nor_x1_sg U60953 ( .A(n25853), .B(n25854), .X(\shifter_0/n10304 ) );
  nor_x1_sg U60954 ( .A(n25883), .B(n25884), .X(\shifter_0/n10300 ) );
  nor_x1_sg U60955 ( .A(n25913), .B(n25914), .X(\shifter_0/n10296 ) );
  nor_x1_sg U60956 ( .A(n25943), .B(n25944), .X(\shifter_0/n10292 ) );
  nor_x1_sg U60957 ( .A(n25973), .B(n25974), .X(\shifter_0/n10288 ) );
  nor_x1_sg U60958 ( .A(n24385), .B(n24386), .X(\shifter_0/n10760 ) );
  nor_x1_sg U60959 ( .A(n24390), .B(n24391), .X(\shifter_0/n10756 ) );
  nor_x1_sg U60960 ( .A(n24395), .B(n24396), .X(\shifter_0/n10752 ) );
  nor_x1_sg U60961 ( .A(n24400), .B(n24401), .X(\shifter_0/n10748 ) );
  nor_x1_sg U60962 ( .A(n24405), .B(n24406), .X(\shifter_0/n10744 ) );
  nor_x1_sg U60963 ( .A(n24410), .B(n24411), .X(\shifter_0/n10740 ) );
  nor_x1_sg U60964 ( .A(n24415), .B(n24416), .X(\shifter_0/n10736 ) );
  nor_x1_sg U60965 ( .A(n24420), .B(n24421), .X(\shifter_0/n10732 ) );
  nor_x1_sg U60966 ( .A(n24425), .B(n24426), .X(\shifter_0/n10728 ) );
  nor_x1_sg U60967 ( .A(n24430), .B(n24431), .X(\shifter_0/n10724 ) );
  nor_x1_sg U60968 ( .A(n24435), .B(n24436), .X(\shifter_0/n10720 ) );
  nor_x1_sg U60969 ( .A(n24440), .B(n24441), .X(\shifter_0/n10716 ) );
  nor_x1_sg U60970 ( .A(n24445), .B(n24446), .X(\shifter_0/n10712 ) );
  nor_x1_sg U60971 ( .A(n24450), .B(n24451), .X(\shifter_0/n10708 ) );
  nor_x1_sg U60972 ( .A(n24455), .B(n24456), .X(\shifter_0/n10704 ) );
  nor_x1_sg U60973 ( .A(n24460), .B(n24461), .X(\shifter_0/n10700 ) );
  nor_x1_sg U60974 ( .A(n24465), .B(n24466), .X(\shifter_0/n10696 ) );
  nor_x1_sg U60975 ( .A(n24470), .B(n24471), .X(\shifter_0/n10692 ) );
  nor_x1_sg U60976 ( .A(n24475), .B(n24476), .X(\shifter_0/n10688 ) );
  nor_x1_sg U60977 ( .A(n24491), .B(n24492), .X(\shifter_0/n10684 ) );
  nor_x1_sg U60978 ( .A(n24497), .B(n24498), .X(\shifter_0/n10680 ) );
  nor_x1_sg U60979 ( .A(n24502), .B(n24503), .X(\shifter_0/n10676 ) );
  nor_x1_sg U60980 ( .A(n24507), .B(n24508), .X(\shifter_0/n10672 ) );
  nor_x1_sg U60981 ( .A(n24512), .B(n24513), .X(\shifter_0/n10668 ) );
  nor_x1_sg U60982 ( .A(n24517), .B(n24518), .X(\shifter_0/n10664 ) );
  nor_x1_sg U60983 ( .A(n24522), .B(n24523), .X(\shifter_0/n10660 ) );
  nor_x1_sg U60984 ( .A(n24527), .B(n24528), .X(\shifter_0/n10656 ) );
  nor_x1_sg U60985 ( .A(n24532), .B(n24533), .X(\shifter_0/n10652 ) );
  nor_x1_sg U60986 ( .A(n24537), .B(n24538), .X(\shifter_0/n10648 ) );
  nor_x1_sg U60987 ( .A(n24542), .B(n24543), .X(\shifter_0/n10644 ) );
  nor_x1_sg U60988 ( .A(n24547), .B(n24548), .X(\shifter_0/n10640 ) );
  nor_x1_sg U60989 ( .A(n24552), .B(n24553), .X(\shifter_0/n10636 ) );
  nor_x1_sg U60990 ( .A(n24557), .B(n24558), .X(\shifter_0/n10632 ) );
  nor_x1_sg U60991 ( .A(n24562), .B(n24563), .X(\shifter_0/n10628 ) );
  nor_x1_sg U60992 ( .A(n24831), .B(n24832), .X(\shifter_0/n10440 ) );
  nor_x1_sg U60993 ( .A(n24861), .B(n24862), .X(\shifter_0/n10436 ) );
  nor_x1_sg U60994 ( .A(n24891), .B(n24892), .X(\shifter_0/n10432 ) );
  nor_x1_sg U60995 ( .A(n24921), .B(n24922), .X(\shifter_0/n10428 ) );
  nor_x1_sg U60996 ( .A(n24951), .B(n24952), .X(\shifter_0/n10424 ) );
  nor_x1_sg U60997 ( .A(n24981), .B(n24982), .X(\shifter_0/n10420 ) );
  nor_x1_sg U60998 ( .A(n25011), .B(n25012), .X(\shifter_0/n10416 ) );
  nor_x1_sg U60999 ( .A(n25041), .B(n25042), .X(\shifter_0/n10412 ) );
  nor_x1_sg U61000 ( .A(n25071), .B(n25072), .X(\shifter_0/n10408 ) );
  nor_x1_sg U61001 ( .A(n25101), .B(n25102), .X(\shifter_0/n10404 ) );
  nor_x1_sg U61002 ( .A(n25131), .B(n25132), .X(\shifter_0/n10400 ) );
  nor_x1_sg U61003 ( .A(n25161), .B(n25162), .X(\shifter_0/n10396 ) );
  nor_x1_sg U61004 ( .A(n25191), .B(n25192), .X(\shifter_0/n10392 ) );
  nor_x1_sg U61005 ( .A(n25221), .B(n25222), .X(\shifter_0/n10388 ) );
  nor_x1_sg U61006 ( .A(n25251), .B(n25252), .X(\shifter_0/n10384 ) );
  nor_x1_sg U61007 ( .A(n25281), .B(n25282), .X(\shifter_0/n10380 ) );
  nor_x1_sg U61008 ( .A(n25311), .B(n25312), .X(\shifter_0/n10376 ) );
  nor_x1_sg U61009 ( .A(n25341), .B(n25342), .X(\shifter_0/n10372 ) );
  nor_x1_sg U61010 ( .A(n25371), .B(n25372), .X(\shifter_0/n10368 ) );
  nor_x1_sg U61011 ( .A(n25403), .B(n25404), .X(\shifter_0/n10364 ) );
  nor_x1_sg U61012 ( .A(n25433), .B(n25434), .X(\shifter_0/n10360 ) );
  nor_x1_sg U61013 ( .A(n25463), .B(n25464), .X(\shifter_0/n10356 ) );
  nor_x1_sg U61014 ( .A(n25493), .B(n25494), .X(\shifter_0/n10352 ) );
  nor_x1_sg U61015 ( .A(n25523), .B(n25524), .X(\shifter_0/n10348 ) );
  nor_x1_sg U61016 ( .A(n25553), .B(n25554), .X(\shifter_0/n10344 ) );
  nor_x1_sg U61017 ( .A(n25583), .B(n25584), .X(\shifter_0/n10340 ) );
  nor_x1_sg U61018 ( .A(n25613), .B(n25614), .X(\shifter_0/n10336 ) );
  nor_x1_sg U61019 ( .A(n25643), .B(n25644), .X(\shifter_0/n10332 ) );
  nor_x1_sg U61020 ( .A(n25673), .B(n25674), .X(\shifter_0/n10328 ) );
  nor_x1_sg U61021 ( .A(n25703), .B(n25704), .X(\shifter_0/n10324 ) );
  nor_x1_sg U61022 ( .A(n25733), .B(n25734), .X(\shifter_0/n10320 ) );
  nor_x1_sg U61023 ( .A(n25763), .B(n25764), .X(\shifter_0/n10316 ) );
  nor_x1_sg U61024 ( .A(n25793), .B(n25794), .X(\shifter_0/n10312 ) );
  nor_x1_sg U61025 ( .A(n25823), .B(n25824), .X(\shifter_0/n10308 ) );
  nor_x1_sg U61026 ( .A(n24379), .B(n24380), .X(\shifter_0/n10764 ) );
  nor_x1_sg U61027 ( .A(n24792), .B(n24793), .X(\shifter_0/n10444 ) );
  nor_x1_sg U61028 ( .A(n57510), .B(n67143), .X(\shifter_0/n12133 ) );
  nor_x1_sg U61029 ( .A(n57510), .B(n67142), .X(\shifter_0/n12129 ) );
  nor_x1_sg U61030 ( .A(n57516), .B(n67356), .X(\shifter_0/n12053 ) );
  nor_x1_sg U61031 ( .A(n57516), .B(n67355), .X(\shifter_0/n12049 ) );
  nor_x1_sg U61032 ( .A(n57507), .B(n67163), .X(\shifter_0/n11973 ) );
  nor_x1_sg U61033 ( .A(n57507), .B(n67162), .X(\shifter_0/n11969 ) );
  nor_x1_sg U61034 ( .A(n57513), .B(n67376), .X(\shifter_0/n11893 ) );
  nor_x1_sg U61035 ( .A(n57513), .B(n67375), .X(\shifter_0/n11889 ) );
  nor_x1_sg U61036 ( .A(n67123), .B(n22498), .X(\shifter_0/n12293 ) );
  nor_x1_sg U61037 ( .A(n67122), .B(n22498), .X(\shifter_0/n12289 ) );
  nor_x1_sg U61038 ( .A(n67336), .B(n22523), .X(\shifter_0/n12213 ) );
  nor_x1_sg U61039 ( .A(n67335), .B(n22523), .X(\shifter_0/n12209 ) );
  nor_x1_sg U61040 ( .A(n67103), .B(n22446), .X(\shifter_0/n12453 ) );
  nor_x1_sg U61041 ( .A(n67102), .B(n22446), .X(\shifter_0/n12449 ) );
  nor_x1_sg U61042 ( .A(n67316), .B(n22473), .X(\shifter_0/n12373 ) );
  nor_x1_sg U61043 ( .A(n67315), .B(n22473), .X(\shifter_0/n12369 ) );
  nor_x1_sg U61044 ( .A(n61880), .B(n22396), .X(\shifter_0/n12613 ) );
  nor_x1_sg U61045 ( .A(n61881), .B(n22396), .X(\shifter_0/n12609 ) );
  nor_x1_sg U61046 ( .A(n61900), .B(n22421), .X(\shifter_0/n12533 ) );
  nor_x1_sg U61047 ( .A(n61901), .B(n22421), .X(\shifter_0/n12529 ) );
  nor_x1_sg U61048 ( .A(n58122), .B(n58121), .X(n24689) );
  nand_x1_sg U61049 ( .A(n67101), .B(n58478), .X(n24690) );
  nor_x1_sg U61050 ( .A(n58052), .B(n58051), .X(n24783) );
  nand_x1_sg U61051 ( .A(n67523), .B(n58478), .X(n24784) );
  nand_x2_sg U61052 ( .A(n26286), .B(n67568), .X(n26282) );
  nand_x2_sg U61053 ( .A(n26284), .B(n26285), .X(n26283) );
  nor_x1_sg U61054 ( .A(n67564), .B(n26266), .X(n26265) );
  nor_x1_sg U61055 ( .A(n26270), .B(n26271), .X(n26264) );
  nand_x2_sg U61056 ( .A(n26267), .B(n26268), .X(n26266) );
  nor_x1_sg U61057 ( .A(n26306), .B(n26307), .X(n26298) );
  nand_x2_sg U61058 ( .A(n26308), .B(n26309), .X(n26307) );
  nand_x1_sg U61059 ( .A(n26085), .B(n67570), .X(n26308) );
  nand_x2_sg U61060 ( .A(n26331), .B(n26332), .X(n26318) );
  nand_x2_sg U61061 ( .A(n26320), .B(n26321), .X(n26319) );
  nand_x1_sg U61062 ( .A(n26333), .B(n57307), .X(n26332) );
  nand_x1_sg U61063 ( .A(n57166), .B(n33783), .X(n33782) );
  nand_x1_sg U61064 ( .A(n57166), .B(n34043), .X(n34042) );
  nor_x1_sg U61065 ( .A(n57394), .B(n46214), .X(n58757) );
  nor_x1_sg U61066 ( .A(n57394), .B(n46215), .X(n58752) );
  nor_x1_sg U61067 ( .A(n57444), .B(n46216), .X(n58747) );
  nor_x1_sg U61068 ( .A(n57439), .B(n46217), .X(n58742) );
  nor_x1_sg U61069 ( .A(n57445), .B(n46218), .X(n58737) );
  nor_x1_sg U61070 ( .A(n57443), .B(n46219), .X(n58732) );
  nor_x1_sg U61071 ( .A(n57439), .B(n46220), .X(n58727) );
  nor_x1_sg U61072 ( .A(n57441), .B(n46221), .X(n58722) );
  nor_x1_sg U61073 ( .A(n57445), .B(n46222), .X(n58717) );
  nor_x1_sg U61074 ( .A(n57439), .B(n46223), .X(n58712) );
  nor_x1_sg U61075 ( .A(n57394), .B(n46224), .X(n58707) );
  nor_x1_sg U61076 ( .A(n57440), .B(n46225), .X(n58702) );
  nor_x1_sg U61077 ( .A(n57397), .B(n46226), .X(n58697) );
  nor_x1_sg U61078 ( .A(n57439), .B(n46227), .X(n58692) );
  nor_x1_sg U61079 ( .A(n57441), .B(n46228), .X(n58687) );
  nor_x1_sg U61080 ( .A(n57441), .B(n46229), .X(n58682) );
  nor_x1_sg U61081 ( .A(n57440), .B(n46230), .X(n58677) );
  nor_x1_sg U61082 ( .A(n57442), .B(n46231), .X(n58672) );
  nor_x1_sg U61083 ( .A(n57396), .B(n46232), .X(n58667) );
  nor_x1_sg U61084 ( .A(n57443), .B(n46233), .X(n61859) );
  nor_x1_sg U61085 ( .A(n57415), .B(n46234), .X(n61852) );
  nor_x1_sg U61086 ( .A(n57415), .B(n46235), .X(n61847) );
  nor_x1_sg U61087 ( .A(n57415), .B(n46236), .X(n61842) );
  nor_x1_sg U61088 ( .A(n57415), .B(n46237), .X(n61837) );
  nor_x1_sg U61089 ( .A(n57415), .B(n46238), .X(n61832) );
  nor_x1_sg U61090 ( .A(n57414), .B(n46239), .X(n61827) );
  nor_x1_sg U61091 ( .A(n57414), .B(n46240), .X(n61822) );
  nor_x1_sg U61092 ( .A(n57414), .B(n46241), .X(n61817) );
  nor_x1_sg U61093 ( .A(n57414), .B(n46242), .X(n61812) );
  nor_x1_sg U61094 ( .A(n57414), .B(n46243), .X(n61807) );
  nor_x1_sg U61095 ( .A(n57414), .B(n46244), .X(n61802) );
  nor_x1_sg U61096 ( .A(n57414), .B(n46245), .X(n61797) );
  nor_x1_sg U61097 ( .A(n57414), .B(n46246), .X(n61792) );
  nor_x1_sg U61098 ( .A(n57414), .B(n46247), .X(n61787) );
  nor_x1_sg U61099 ( .A(n57413), .B(n46248), .X(n61782) );
  nor_x1_sg U61100 ( .A(n57413), .B(n46249), .X(n61777) );
  nor_x1_sg U61101 ( .A(n57413), .B(n46250), .X(n61772) );
  nor_x1_sg U61102 ( .A(n57413), .B(n46251), .X(n61767) );
  nor_x1_sg U61103 ( .A(n57413), .B(n46252), .X(n61762) );
  nor_x1_sg U61104 ( .A(n57413), .B(n46253), .X(n61757) );
  nor_x1_sg U61105 ( .A(n57413), .B(n46254), .X(n61752) );
  nor_x1_sg U61106 ( .A(n57413), .B(n46255), .X(n61747) );
  nor_x1_sg U61107 ( .A(n57413), .B(n46256), .X(n61742) );
  nor_x1_sg U61108 ( .A(n57412), .B(n46257), .X(n61737) );
  nor_x1_sg U61109 ( .A(n57412), .B(n46258), .X(n61732) );
  nor_x1_sg U61110 ( .A(n57412), .B(n46259), .X(n61727) );
  nor_x1_sg U61111 ( .A(n57412), .B(n46260), .X(n61722) );
  nor_x1_sg U61112 ( .A(n57412), .B(n46261), .X(n61717) );
  nor_x1_sg U61113 ( .A(n57412), .B(n46262), .X(n61712) );
  nor_x1_sg U61114 ( .A(n57412), .B(n46263), .X(n61707) );
  nor_x1_sg U61115 ( .A(n57412), .B(n46264), .X(n61702) );
  nor_x1_sg U61116 ( .A(n57412), .B(n46265), .X(n61697) );
  nor_x1_sg U61117 ( .A(n57411), .B(n46266), .X(n61692) );
  nor_x1_sg U61118 ( .A(n57411), .B(n46267), .X(n61687) );
  nor_x1_sg U61119 ( .A(n57411), .B(n46268), .X(n61682) );
  nor_x1_sg U61120 ( .A(n57411), .B(n46269), .X(n61677) );
  nor_x1_sg U61121 ( .A(n57411), .B(n46270), .X(n61672) );
  nor_x1_sg U61122 ( .A(n57411), .B(n46271), .X(n61667) );
  nor_x1_sg U61123 ( .A(n57411), .B(n46272), .X(n61662) );
  nor_x1_sg U61124 ( .A(n57411), .B(n46273), .X(n61657) );
  nor_x1_sg U61125 ( .A(n57411), .B(n46274), .X(n61652) );
  nor_x1_sg U61126 ( .A(n57410), .B(n46275), .X(n61647) );
  nor_x1_sg U61127 ( .A(n57410), .B(n46276), .X(n61642) );
  nor_x1_sg U61128 ( .A(n57410), .B(n46277), .X(n61637) );
  nor_x1_sg U61129 ( .A(n57410), .B(n46278), .X(n61632) );
  nor_x1_sg U61130 ( .A(n57410), .B(n46279), .X(n61627) );
  nor_x1_sg U61131 ( .A(n57410), .B(n46280), .X(n61622) );
  nor_x1_sg U61132 ( .A(n57410), .B(n46281), .X(n61617) );
  nor_x1_sg U61133 ( .A(n57410), .B(n46282), .X(n61612) );
  nor_x1_sg U61134 ( .A(n57410), .B(n46283), .X(n61607) );
  nor_x1_sg U61135 ( .A(n57409), .B(n46284), .X(n61602) );
  nor_x1_sg U61136 ( .A(n57409), .B(n46285), .X(n61597) );
  nor_x1_sg U61137 ( .A(n57409), .B(n46286), .X(n61592) );
  nor_x1_sg U61138 ( .A(n57409), .B(n46287), .X(n61587) );
  nor_x1_sg U61139 ( .A(n57409), .B(n46288), .X(n61582) );
  nor_x1_sg U61140 ( .A(n57409), .B(n46289), .X(n61577) );
  nor_x1_sg U61141 ( .A(n57409), .B(n46290), .X(n61572) );
  nor_x1_sg U61142 ( .A(n57409), .B(n46291), .X(n61567) );
  nor_x1_sg U61143 ( .A(n57409), .B(n46292), .X(n61562) );
  nor_x1_sg U61144 ( .A(n57408), .B(n46293), .X(n61557) );
  nor_x1_sg U61145 ( .A(n57408), .B(n46294), .X(n61552) );
  nor_x1_sg U61146 ( .A(n57408), .B(n46295), .X(n61547) );
  nor_x1_sg U61147 ( .A(n57408), .B(n46296), .X(n61542) );
  nor_x1_sg U61148 ( .A(n57408), .B(n46297), .X(n61537) );
  nor_x1_sg U61149 ( .A(n57408), .B(n46298), .X(n61532) );
  nor_x1_sg U61150 ( .A(n57408), .B(n46299), .X(n61527) );
  nor_x1_sg U61151 ( .A(n57408), .B(n46300), .X(n61522) );
  nor_x1_sg U61152 ( .A(n57408), .B(n46301), .X(n61517) );
  nor_x1_sg U61153 ( .A(n57407), .B(n46302), .X(n61512) );
  nor_x1_sg U61154 ( .A(n57407), .B(n46303), .X(n61507) );
  nor_x1_sg U61155 ( .A(n57407), .B(n46304), .X(n61502) );
  nor_x1_sg U61156 ( .A(n57407), .B(n46305), .X(n61497) );
  nor_x1_sg U61157 ( .A(n57407), .B(n46306), .X(n61492) );
  nor_x1_sg U61158 ( .A(n57407), .B(n46307), .X(n61487) );
  nor_x1_sg U61159 ( .A(n57407), .B(n46308), .X(n61482) );
  nor_x1_sg U61160 ( .A(n57407), .B(n46309), .X(n61477) );
  nor_x1_sg U61161 ( .A(n57407), .B(n46310), .X(n61472) );
  nor_x1_sg U61162 ( .A(n57406), .B(n46311), .X(n61467) );
  nor_x1_sg U61163 ( .A(n57406), .B(n46312), .X(n61462) );
  nor_x1_sg U61164 ( .A(n57406), .B(n46313), .X(n61457) );
  nor_x1_sg U61165 ( .A(n57406), .B(n46314), .X(n61452) );
  nor_x1_sg U61166 ( .A(n57406), .B(n46315), .X(n61447) );
  nor_x1_sg U61167 ( .A(n57406), .B(n46316), .X(n61442) );
  nor_x1_sg U61168 ( .A(n57406), .B(n46317), .X(n61437) );
  nor_x1_sg U61169 ( .A(n57406), .B(n46318), .X(n61432) );
  nor_x1_sg U61170 ( .A(n57405), .B(n46319), .X(n61427) );
  nor_x1_sg U61171 ( .A(n57405), .B(n46320), .X(n61422) );
  nor_x1_sg U61172 ( .A(n57405), .B(n46321), .X(n61417) );
  nor_x1_sg U61173 ( .A(n57405), .B(n46322), .X(n61412) );
  nor_x1_sg U61174 ( .A(n57405), .B(n46323), .X(n61407) );
  nor_x1_sg U61175 ( .A(n57405), .B(n46324), .X(n61402) );
  nor_x1_sg U61176 ( .A(n57405), .B(n46325), .X(n61397) );
  nor_x1_sg U61177 ( .A(n57405), .B(n46326), .X(n61392) );
  nor_x1_sg U61178 ( .A(n57405), .B(n46327), .X(n61387) );
  nor_x1_sg U61179 ( .A(n57404), .B(n46328), .X(n61382) );
  nor_x1_sg U61180 ( .A(n57404), .B(n46329), .X(n61377) );
  nor_x1_sg U61181 ( .A(n57404), .B(n46330), .X(n61372) );
  nor_x1_sg U61182 ( .A(n57404), .B(n46331), .X(n61367) );
  nor_x1_sg U61183 ( .A(n57404), .B(n46332), .X(n61362) );
  nor_x1_sg U61184 ( .A(n57404), .B(n46333), .X(n61357) );
  nor_x1_sg U61185 ( .A(n57404), .B(n46334), .X(n61352) );
  nor_x1_sg U61186 ( .A(n57404), .B(n46335), .X(n61347) );
  nor_x1_sg U61187 ( .A(n57404), .B(n46336), .X(n61342) );
  nor_x1_sg U61188 ( .A(n57403), .B(n46337), .X(n61337) );
  nor_x1_sg U61189 ( .A(n57403), .B(n46338), .X(n61332) );
  nor_x1_sg U61190 ( .A(n57403), .B(n46339), .X(n61327) );
  nor_x1_sg U61191 ( .A(n57403), .B(n46340), .X(n61322) );
  nor_x1_sg U61192 ( .A(n57403), .B(n46341), .X(n61317) );
  nor_x1_sg U61193 ( .A(n57403), .B(n46342), .X(n61312) );
  nor_x1_sg U61194 ( .A(n57403), .B(n46343), .X(n61307) );
  nor_x1_sg U61195 ( .A(n57403), .B(n46344), .X(n61302) );
  nor_x1_sg U61196 ( .A(n57403), .B(n46345), .X(n61297) );
  nor_x1_sg U61197 ( .A(n57402), .B(n46346), .X(n61292) );
  nor_x1_sg U61198 ( .A(n57402), .B(n46347), .X(n61287) );
  nor_x1_sg U61199 ( .A(n57402), .B(n46348), .X(n61282) );
  nor_x1_sg U61200 ( .A(n57402), .B(n46349), .X(n61277) );
  nor_x1_sg U61201 ( .A(n57402), .B(n46350), .X(n61272) );
  nor_x1_sg U61202 ( .A(n57402), .B(n46351), .X(n61267) );
  nor_x1_sg U61203 ( .A(n57402), .B(n46352), .X(n61262) );
  nor_x1_sg U61204 ( .A(n57402), .B(n46353), .X(n61257) );
  nor_x1_sg U61205 ( .A(n57402), .B(n46354), .X(n61252) );
  nor_x1_sg U61206 ( .A(n57401), .B(n46355), .X(n61247) );
  nor_x1_sg U61207 ( .A(n57401), .B(n46356), .X(n61242) );
  nor_x1_sg U61208 ( .A(n57401), .B(n46357), .X(n61237) );
  nor_x1_sg U61209 ( .A(n57401), .B(n46358), .X(n61232) );
  nor_x1_sg U61210 ( .A(n57401), .B(n46359), .X(n61227) );
  nor_x1_sg U61211 ( .A(n57401), .B(n46360), .X(n61222) );
  nor_x1_sg U61212 ( .A(n57401), .B(n46361), .X(n61217) );
  nor_x1_sg U61213 ( .A(n57401), .B(n46362), .X(n61212) );
  nor_x1_sg U61214 ( .A(n57401), .B(n46363), .X(n61207) );
  nor_x1_sg U61215 ( .A(n57400), .B(n46364), .X(n61202) );
  nor_x1_sg U61216 ( .A(n57400), .B(n46365), .X(n61197) );
  nor_x1_sg U61217 ( .A(n57400), .B(n46366), .X(n61192) );
  nor_x1_sg U61218 ( .A(n57400), .B(n46367), .X(n61187) );
  nor_x1_sg U61219 ( .A(n57400), .B(n46368), .X(n61182) );
  nor_x1_sg U61220 ( .A(n57400), .B(n46369), .X(n61177) );
  nor_x1_sg U61221 ( .A(n57400), .B(n46370), .X(n61172) );
  nor_x1_sg U61222 ( .A(n57400), .B(n46371), .X(n61167) );
  nor_x1_sg U61223 ( .A(n57400), .B(n46372), .X(n61162) );
  nor_x1_sg U61224 ( .A(n57399), .B(n46373), .X(n61157) );
  nor_x1_sg U61225 ( .A(n57399), .B(n46374), .X(n61152) );
  nor_x1_sg U61226 ( .A(n57399), .B(n46375), .X(n61147) );
  nor_x1_sg U61227 ( .A(n57399), .B(n46376), .X(n61142) );
  nor_x1_sg U61228 ( .A(n57399), .B(n46377), .X(n61137) );
  nor_x1_sg U61229 ( .A(n57399), .B(n46378), .X(n61132) );
  nor_x1_sg U61230 ( .A(n57399), .B(n46379), .X(n61127) );
  nor_x1_sg U61231 ( .A(n57399), .B(n46380), .X(n61122) );
  nor_x1_sg U61232 ( .A(n57399), .B(n46381), .X(n61117) );
  nor_x1_sg U61233 ( .A(n57398), .B(n46382), .X(n61112) );
  nor_x1_sg U61234 ( .A(n57398), .B(n46383), .X(n61107) );
  nor_x1_sg U61235 ( .A(n57398), .B(n46384), .X(n61102) );
  nor_x1_sg U61236 ( .A(n57398), .B(n46385), .X(n61097) );
  nor_x1_sg U61237 ( .A(n57398), .B(n46386), .X(n61092) );
  nor_x1_sg U61238 ( .A(n57398), .B(n46387), .X(n61087) );
  nor_x1_sg U61239 ( .A(n57398), .B(n46388), .X(n61082) );
  nor_x1_sg U61240 ( .A(n57398), .B(n46389), .X(n61077) );
  nor_x1_sg U61241 ( .A(n57398), .B(n46390), .X(n61072) );
  nor_x1_sg U61242 ( .A(n57413), .B(n46391), .X(n61067) );
  nor_x1_sg U61243 ( .A(n57410), .B(n46392), .X(n61062) );
  nor_x1_sg U61244 ( .A(n57406), .B(n46393), .X(n61057) );
  nor_x1_sg U61245 ( .A(n57430), .B(n46394), .X(n61052) );
  nor_x1_sg U61246 ( .A(n57430), .B(n46395), .X(n61047) );
  nor_x1_sg U61247 ( .A(n57430), .B(n46396), .X(n61042) );
  nor_x1_sg U61248 ( .A(n57446), .B(n46397), .X(n61037) );
  nor_x1_sg U61249 ( .A(n57446), .B(n46398), .X(n61032) );
  nor_x1_sg U61250 ( .A(n57440), .B(n46399), .X(n61027) );
  nor_x1_sg U61251 ( .A(n57439), .B(n46400), .X(n61022) );
  nor_x1_sg U61252 ( .A(n57439), .B(n46401), .X(n61017) );
  nor_x1_sg U61253 ( .A(n57439), .B(n46402), .X(n61012) );
  nor_x1_sg U61254 ( .A(n57396), .B(n46403), .X(n61007) );
  nor_x1_sg U61255 ( .A(n57440), .B(n46404), .X(n61002) );
  nor_x1_sg U61256 ( .A(n57444), .B(n46405), .X(n60997) );
  nor_x1_sg U61257 ( .A(n57394), .B(n46406), .X(n60992) );
  nor_x1_sg U61258 ( .A(n57394), .B(n46407), .X(n60987) );
  nor_x1_sg U61259 ( .A(n57444), .B(n46408), .X(n60982) );
  nor_x1_sg U61260 ( .A(n57439), .B(n46409), .X(n60977) );
  nor_x1_sg U61261 ( .A(n57440), .B(n46410), .X(n60972) );
  nor_x1_sg U61262 ( .A(n57441), .B(n46411), .X(n60967) );
  nor_x1_sg U61263 ( .A(n57441), .B(n46412), .X(n60962) );
  nor_x1_sg U61264 ( .A(n57394), .B(n46413), .X(n60957) );
  nor_x1_sg U61265 ( .A(n57396), .B(n46414), .X(n60952) );
  nor_x1_sg U61266 ( .A(n57444), .B(n46415), .X(n60947) );
  nor_x1_sg U61267 ( .A(n57445), .B(n46416), .X(n60942) );
  nor_x1_sg U61268 ( .A(n57440), .B(n46417), .X(n60937) );
  nor_x1_sg U61269 ( .A(n57439), .B(n46418), .X(n60932) );
  nor_x1_sg U61270 ( .A(n57397), .B(n46419), .X(n60927) );
  nor_x1_sg U61271 ( .A(n57443), .B(n46420), .X(n60922) );
  nor_x1_sg U61272 ( .A(n57446), .B(n46421), .X(n60917) );
  nor_x1_sg U61273 ( .A(n57396), .B(n46422), .X(n60912) );
  nor_x1_sg U61274 ( .A(n57442), .B(n46423), .X(n60907) );
  nor_x1_sg U61275 ( .A(n57429), .B(n46424), .X(n60902) );
  nor_x1_sg U61276 ( .A(n57429), .B(n46425), .X(n60897) );
  nor_x1_sg U61277 ( .A(n57429), .B(n46426), .X(n60892) );
  nor_x1_sg U61278 ( .A(n57429), .B(n46427), .X(n60887) );
  nor_x1_sg U61279 ( .A(n57429), .B(n46428), .X(n60882) );
  nor_x1_sg U61280 ( .A(n57429), .B(n46429), .X(n60877) );
  nor_x1_sg U61281 ( .A(n57429), .B(n46430), .X(n60872) );
  nor_x1_sg U61282 ( .A(n57429), .B(n46431), .X(n60867) );
  nor_x1_sg U61283 ( .A(n57429), .B(n46432), .X(n60862) );
  nor_x1_sg U61284 ( .A(n57428), .B(n46433), .X(n60857) );
  nor_x1_sg U61285 ( .A(n57428), .B(n46434), .X(n60852) );
  nor_x1_sg U61286 ( .A(n57428), .B(n46435), .X(n60847) );
  nor_x1_sg U61287 ( .A(n57428), .B(n46436), .X(n60842) );
  nor_x1_sg U61288 ( .A(n57428), .B(n46437), .X(n60837) );
  nor_x1_sg U61289 ( .A(n57428), .B(n46438), .X(n60832) );
  nor_x1_sg U61290 ( .A(n57428), .B(n46439), .X(n60827) );
  nor_x1_sg U61291 ( .A(n57428), .B(n46440), .X(n60822) );
  nor_x1_sg U61292 ( .A(n57428), .B(n46441), .X(n60817) );
  nor_x1_sg U61293 ( .A(n57427), .B(n46442), .X(n60812) );
  nor_x1_sg U61294 ( .A(n57427), .B(n46443), .X(n60807) );
  nor_x1_sg U61295 ( .A(n57427), .B(n46444), .X(n60802) );
  nor_x1_sg U61296 ( .A(n57427), .B(n46445), .X(n60797) );
  nor_x1_sg U61297 ( .A(n57427), .B(n46446), .X(n60792) );
  nor_x1_sg U61298 ( .A(n57427), .B(n46447), .X(n60787) );
  nor_x1_sg U61299 ( .A(n57427), .B(n46448), .X(n60782) );
  nor_x1_sg U61300 ( .A(n57427), .B(n46449), .X(n60777) );
  nor_x1_sg U61301 ( .A(n57427), .B(n46450), .X(n60772) );
  nor_x1_sg U61302 ( .A(n57426), .B(n46451), .X(n60767) );
  nor_x1_sg U61303 ( .A(n57426), .B(n46452), .X(n60762) );
  nor_x1_sg U61304 ( .A(n57426), .B(n46453), .X(n60757) );
  nor_x1_sg U61305 ( .A(n57426), .B(n46454), .X(n60752) );
  nor_x1_sg U61306 ( .A(n57426), .B(n46455), .X(n60747) );
  nor_x1_sg U61307 ( .A(n57426), .B(n46456), .X(n60742) );
  nor_x1_sg U61308 ( .A(n57426), .B(n46457), .X(n60737) );
  nor_x1_sg U61309 ( .A(n57426), .B(n46458), .X(n60732) );
  nor_x1_sg U61310 ( .A(n57426), .B(n46459), .X(n60727) );
  nor_x1_sg U61311 ( .A(n57425), .B(n46460), .X(n60722) );
  nor_x1_sg U61312 ( .A(n57425), .B(n46461), .X(n60717) );
  nor_x1_sg U61313 ( .A(n57425), .B(n46462), .X(n60712) );
  nor_x1_sg U61314 ( .A(n57425), .B(n46463), .X(n60707) );
  nor_x1_sg U61315 ( .A(n57425), .B(n46464), .X(n60702) );
  nor_x1_sg U61316 ( .A(n57425), .B(n46465), .X(n60697) );
  nor_x1_sg U61317 ( .A(n57425), .B(n46466), .X(n60692) );
  nor_x1_sg U61318 ( .A(n57425), .B(n46467), .X(n60687) );
  nor_x1_sg U61319 ( .A(n57425), .B(n46468), .X(n60682) );
  nor_x1_sg U61320 ( .A(n57424), .B(n46469), .X(n60677) );
  nor_x1_sg U61321 ( .A(n57424), .B(n46470), .X(n60672) );
  nor_x1_sg U61322 ( .A(n57424), .B(n46471), .X(n60667) );
  nor_x1_sg U61323 ( .A(n57424), .B(n46472), .X(n60662) );
  nor_x1_sg U61324 ( .A(n57424), .B(n46473), .X(n60657) );
  nor_x1_sg U61325 ( .A(n57424), .B(n46474), .X(n60652) );
  nor_x1_sg U61326 ( .A(n57424), .B(n46475), .X(n60647) );
  nor_x1_sg U61327 ( .A(n57424), .B(n46476), .X(n60642) );
  nor_x1_sg U61328 ( .A(n57423), .B(n46477), .X(n60637) );
  nor_x1_sg U61329 ( .A(n57423), .B(n46478), .X(n60632) );
  nor_x1_sg U61330 ( .A(n57423), .B(n46479), .X(n60627) );
  nor_x1_sg U61331 ( .A(n57423), .B(n46480), .X(n60622) );
  nor_x1_sg U61332 ( .A(n57423), .B(n46481), .X(n60617) );
  nor_x1_sg U61333 ( .A(n57423), .B(n46482), .X(n60612) );
  nor_x1_sg U61334 ( .A(n57423), .B(n46483), .X(n60607) );
  nor_x1_sg U61335 ( .A(n57423), .B(n46484), .X(n60602) );
  nor_x1_sg U61336 ( .A(n57423), .B(n46485), .X(n60597) );
  nor_x1_sg U61337 ( .A(n57422), .B(n46486), .X(n60592) );
  nor_x1_sg U61338 ( .A(n57422), .B(n46487), .X(n60587) );
  nor_x1_sg U61339 ( .A(n57422), .B(n46488), .X(n60582) );
  nor_x1_sg U61340 ( .A(n57422), .B(n46489), .X(n60577) );
  nor_x1_sg U61341 ( .A(n57422), .B(n46490), .X(n60572) );
  nor_x1_sg U61342 ( .A(n57422), .B(n46491), .X(n60567) );
  nor_x1_sg U61343 ( .A(n57422), .B(n46492), .X(n60562) );
  nor_x1_sg U61344 ( .A(n57422), .B(n46493), .X(n60557) );
  nor_x1_sg U61345 ( .A(n57422), .B(n46494), .X(n60552) );
  nor_x1_sg U61346 ( .A(n57421), .B(n46495), .X(n60547) );
  nor_x1_sg U61347 ( .A(n57421), .B(n46496), .X(n60542) );
  nor_x1_sg U61348 ( .A(n57421), .B(n46497), .X(n60537) );
  nor_x1_sg U61349 ( .A(n57421), .B(n46498), .X(n60532) );
  nor_x1_sg U61350 ( .A(n57421), .B(n46499), .X(n60527) );
  nor_x1_sg U61351 ( .A(n57421), .B(n46500), .X(n60522) );
  nor_x1_sg U61352 ( .A(n57421), .B(n46501), .X(n60517) );
  nor_x1_sg U61353 ( .A(n57421), .B(n46502), .X(n60512) );
  nor_x1_sg U61354 ( .A(n57421), .B(n46503), .X(n60507) );
  nor_x1_sg U61355 ( .A(n57420), .B(n46504), .X(n60502) );
  nor_x1_sg U61356 ( .A(n57420), .B(n46505), .X(n60497) );
  nor_x1_sg U61357 ( .A(n57420), .B(n46506), .X(n60492) );
  nor_x1_sg U61358 ( .A(n57420), .B(n46507), .X(n60487) );
  nor_x1_sg U61359 ( .A(n57420), .B(n46508), .X(n60482) );
  nor_x1_sg U61360 ( .A(n57420), .B(n46509), .X(n60477) );
  nor_x1_sg U61361 ( .A(n57420), .B(n46510), .X(n60472) );
  nor_x1_sg U61362 ( .A(n57420), .B(n46511), .X(n60467) );
  nor_x1_sg U61363 ( .A(n57420), .B(n46512), .X(n60462) );
  nor_x1_sg U61364 ( .A(n57419), .B(n46513), .X(n60457) );
  nor_x1_sg U61365 ( .A(n57419), .B(n46514), .X(n60452) );
  nor_x1_sg U61366 ( .A(n57419), .B(n46515), .X(n60447) );
  nor_x1_sg U61367 ( .A(n57419), .B(n46516), .X(n60442) );
  nor_x1_sg U61368 ( .A(n57419), .B(n46517), .X(n60437) );
  nor_x1_sg U61369 ( .A(n57419), .B(n46518), .X(n60432) );
  nor_x1_sg U61370 ( .A(n57419), .B(n46519), .X(n60427) );
  nor_x1_sg U61371 ( .A(n57419), .B(n46520), .X(n60422) );
  nor_x1_sg U61372 ( .A(n57419), .B(n46521), .X(n60417) );
  nor_x1_sg U61373 ( .A(n57418), .B(n46522), .X(n60412) );
  nor_x1_sg U61374 ( .A(n57418), .B(n46523), .X(n60407) );
  nor_x1_sg U61375 ( .A(n57418), .B(n46524), .X(n60402) );
  nor_x1_sg U61376 ( .A(n57418), .B(n46525), .X(n60397) );
  nor_x1_sg U61377 ( .A(n57418), .B(n46526), .X(n60392) );
  nor_x1_sg U61378 ( .A(n57418), .B(n46527), .X(n60387) );
  nor_x1_sg U61379 ( .A(n57418), .B(n46528), .X(n60382) );
  nor_x1_sg U61380 ( .A(n57418), .B(n46529), .X(n60377) );
  nor_x1_sg U61381 ( .A(n57418), .B(n46530), .X(n60372) );
  nor_x1_sg U61382 ( .A(n57417), .B(n46531), .X(n60367) );
  nor_x1_sg U61383 ( .A(n57417), .B(n46532), .X(n60362) );
  nor_x1_sg U61384 ( .A(n57417), .B(n46533), .X(n60357) );
  nor_x1_sg U61385 ( .A(n57417), .B(n46534), .X(n60352) );
  nor_x1_sg U61386 ( .A(n57417), .B(n46535), .X(n60347) );
  nor_x1_sg U61387 ( .A(n57417), .B(n46536), .X(n60342) );
  nor_x1_sg U61388 ( .A(n57417), .B(n46537), .X(n60337) );
  nor_x1_sg U61389 ( .A(n57417), .B(n46538), .X(n60332) );
  nor_x1_sg U61390 ( .A(n57417), .B(n46539), .X(n60327) );
  nor_x1_sg U61391 ( .A(n57416), .B(n46540), .X(n60322) );
  nor_x1_sg U61392 ( .A(n57416), .B(n46541), .X(n60317) );
  nor_x1_sg U61393 ( .A(n57416), .B(n46542), .X(n60312) );
  nor_x1_sg U61394 ( .A(n57416), .B(n46543), .X(n60307) );
  nor_x1_sg U61395 ( .A(n57416), .B(n46544), .X(n60302) );
  nor_x1_sg U61396 ( .A(n57416), .B(n46545), .X(n60297) );
  nor_x1_sg U61397 ( .A(n57416), .B(n46546), .X(n60292) );
  nor_x1_sg U61398 ( .A(n57416), .B(n46547), .X(n60287) );
  nor_x1_sg U61399 ( .A(n57416), .B(n46548), .X(n60282) );
  nor_x1_sg U61400 ( .A(n57415), .B(n46549), .X(n60277) );
  nor_x1_sg U61401 ( .A(n57415), .B(n46550), .X(n60272) );
  nor_x1_sg U61402 ( .A(n57415), .B(n46551), .X(n60267) );
  nor_x1_sg U61403 ( .A(n57415), .B(n46552), .X(n60262) );
  nor_x1_sg U61404 ( .A(n57424), .B(n46553), .X(n60257) );
  nor_x1_sg U61405 ( .A(n57394), .B(n46554), .X(n60252) );
  nor_x1_sg U61406 ( .A(n57396), .B(n46555), .X(n60247) );
  nor_x1_sg U61407 ( .A(n57396), .B(n46556), .X(n60242) );
  nor_x1_sg U61408 ( .A(n57394), .B(n46557), .X(n60237) );
  nor_x1_sg U61409 ( .A(n57440), .B(n46558), .X(n60232) );
  nor_x1_sg U61410 ( .A(n57446), .B(n46559), .X(n60227) );
  nor_x1_sg U61411 ( .A(n57394), .B(n46560), .X(n60222) );
  nor_x1_sg U61412 ( .A(n57396), .B(n46561), .X(n60217) );
  nor_x1_sg U61413 ( .A(n57396), .B(n46562), .X(n60212) );
  nor_x1_sg U61414 ( .A(n57394), .B(n46563), .X(n60207) );
  nor_x1_sg U61415 ( .A(n57443), .B(n46564), .X(n60202) );
  nor_x1_sg U61416 ( .A(n57394), .B(n46565), .X(n60197) );
  nor_x1_sg U61417 ( .A(n57440), .B(n46566), .X(n60192) );
  nor_x1_sg U61418 ( .A(n57442), .B(n46567), .X(n60187) );
  nor_x1_sg U61419 ( .A(n57439), .B(n46568), .X(n60182) );
  nor_x1_sg U61420 ( .A(n57439), .B(n46569), .X(n60177) );
  nor_x1_sg U61421 ( .A(n57440), .B(n46570), .X(n60172) );
  nor_x1_sg U61422 ( .A(n57411), .B(n46571), .X(n60167) );
  nor_x1_sg U61423 ( .A(n57396), .B(n46572), .X(n60162) );
  nor_x1_sg U61424 ( .A(n57439), .B(n46573), .X(n60157) );
  nor_x1_sg U61425 ( .A(n57442), .B(n46574), .X(n60152) );
  nor_x1_sg U61426 ( .A(n57446), .B(n46575), .X(n60147) );
  nor_x1_sg U61427 ( .A(n57441), .B(n46576), .X(n60142) );
  nor_x1_sg U61428 ( .A(n57444), .B(n46577), .X(n60137) );
  nor_x1_sg U61429 ( .A(n57444), .B(n46578), .X(n60132) );
  nor_x1_sg U61430 ( .A(n57445), .B(n46579), .X(n60127) );
  nor_x1_sg U61431 ( .A(n57442), .B(n46580), .X(n60122) );
  nor_x1_sg U61432 ( .A(n57440), .B(n46581), .X(n60117) );
  nor_x1_sg U61433 ( .A(n57394), .B(n46582), .X(n60112) );
  nor_x1_sg U61434 ( .A(n57439), .B(n46583), .X(n60107) );
  nor_x1_sg U61435 ( .A(n57443), .B(n46584), .X(n60102) );
  nor_x1_sg U61436 ( .A(n57439), .B(n46585), .X(n60097) );
  nor_x1_sg U61437 ( .A(n57446), .B(n46586), .X(n60092) );
  nor_x1_sg U61438 ( .A(n57441), .B(n46587), .X(n60087) );
  nor_x1_sg U61439 ( .A(n57396), .B(n46588), .X(n60082) );
  nor_x1_sg U61440 ( .A(n57442), .B(n46589), .X(n60077) );
  nor_x1_sg U61441 ( .A(n57444), .B(n46590), .X(n60072) );
  nor_x1_sg U61442 ( .A(n57445), .B(n46591), .X(n60067) );
  nor_x1_sg U61443 ( .A(n57440), .B(n46592), .X(n60062) );
  nor_x1_sg U61444 ( .A(n57445), .B(n46593), .X(n60057) );
  nor_x1_sg U61445 ( .A(n57397), .B(n46594), .X(n60052) );
  nor_x1_sg U61446 ( .A(n57443), .B(n46595), .X(n60047) );
  nor_x1_sg U61447 ( .A(n57439), .B(n46596), .X(n60042) );
  nor_x1_sg U61448 ( .A(n57410), .B(n46597), .X(n60037) );
  nor_x1_sg U61449 ( .A(n57413), .B(n46598), .X(n60032) );
  nor_x1_sg U61450 ( .A(n57446), .B(n46599), .X(n60027) );
  nor_x1_sg U61451 ( .A(n57441), .B(n46600), .X(n60022) );
  nor_x1_sg U61452 ( .A(n57394), .B(n46601), .X(n60017) );
  nor_x1_sg U61453 ( .A(n57444), .B(n46602), .X(n60012) );
  nor_x1_sg U61454 ( .A(n57445), .B(n46603), .X(n60007) );
  nor_x1_sg U61455 ( .A(n57439), .B(n46604), .X(n60002) );
  nor_x1_sg U61456 ( .A(n57443), .B(n46605), .X(n59997) );
  nor_x1_sg U61457 ( .A(n57440), .B(n46606), .X(n59992) );
  nor_x1_sg U61458 ( .A(n57446), .B(n46607), .X(n59987) );
  nor_x1_sg U61459 ( .A(n57443), .B(n46608), .X(n59982) );
  nor_x1_sg U61460 ( .A(n57441), .B(n46609), .X(n59977) );
  nor_x1_sg U61461 ( .A(n57445), .B(n46610), .X(n59972) );
  nor_x1_sg U61462 ( .A(n57442), .B(n46611), .X(n59967) );
  nor_x1_sg U61463 ( .A(n57439), .B(n46612), .X(n59962) );
  nor_x1_sg U61464 ( .A(n57444), .B(n46613), .X(n59957) );
  nor_x1_sg U61465 ( .A(n57443), .B(n46614), .X(n59952) );
  nor_x1_sg U61466 ( .A(n57412), .B(n46615), .X(n59947) );
  nor_x1_sg U61467 ( .A(n57439), .B(n46616), .X(n59942) );
  nor_x1_sg U61468 ( .A(n57394), .B(n46617), .X(n59937) );
  nor_x1_sg U61469 ( .A(n57439), .B(n46618), .X(n59932) );
  nor_x1_sg U61470 ( .A(n57440), .B(n46619), .X(n59927) );
  nor_x1_sg U61471 ( .A(n57442), .B(n46620), .X(n59922) );
  nor_x1_sg U61472 ( .A(n57446), .B(n46621), .X(n59917) );
  nor_x1_sg U61473 ( .A(n57439), .B(n46622), .X(n59912) );
  nor_x1_sg U61474 ( .A(n57443), .B(n46623), .X(n59907) );
  nor_x1_sg U61475 ( .A(n57439), .B(n46624), .X(n59902) );
  nor_x1_sg U61476 ( .A(n57446), .B(n46625), .X(n59897) );
  nor_x1_sg U61477 ( .A(n57440), .B(n46626), .X(n59892) );
  nor_x1_sg U61478 ( .A(n57443), .B(n46627), .X(n59887) );
  nor_x1_sg U61479 ( .A(n57412), .B(n46628), .X(n59882) );
  nor_x1_sg U61480 ( .A(n57413), .B(n46629), .X(n59877) );
  nor_x1_sg U61481 ( .A(n57410), .B(n46630), .X(n59872) );
  nor_x1_sg U61482 ( .A(n57411), .B(n46631), .X(n59867) );
  nor_x1_sg U61483 ( .A(n57442), .B(n46632), .X(n59862) );
  nor_x1_sg U61484 ( .A(n57446), .B(n46633), .X(n59857) );
  nor_x1_sg U61485 ( .A(n57439), .B(n46634), .X(n59852) );
  nor_x1_sg U61486 ( .A(n57441), .B(n46635), .X(n59847) );
  nor_x1_sg U61487 ( .A(n57439), .B(n46636), .X(n59842) );
  nor_x1_sg U61488 ( .A(n57440), .B(n46637), .X(n59837) );
  nor_x1_sg U61489 ( .A(n57445), .B(n46638), .X(n59832) );
  nor_x1_sg U61490 ( .A(n57412), .B(n46639), .X(n59827) );
  nor_x1_sg U61491 ( .A(n57413), .B(n46640), .X(n59822) );
  nor_x1_sg U61492 ( .A(n57394), .B(n46641), .X(n59817) );
  nor_x1_sg U61493 ( .A(n57444), .B(n46642), .X(n59812) );
  nor_x1_sg U61494 ( .A(n57445), .B(n46643), .X(n59807) );
  nor_x1_sg U61495 ( .A(n57443), .B(n46644), .X(n59802) );
  nor_x1_sg U61496 ( .A(n57444), .B(n46645), .X(n59797) );
  nor_x1_sg U61497 ( .A(n57445), .B(n46646), .X(n59792) );
  nor_x1_sg U61498 ( .A(n57446), .B(n46647), .X(n59787) );
  nor_x1_sg U61499 ( .A(n57443), .B(n46648), .X(n59782) );
  nor_x1_sg U61500 ( .A(n57444), .B(n46649), .X(n59777) );
  nor_x1_sg U61501 ( .A(n57445), .B(n46650), .X(n59772) );
  nor_x1_sg U61502 ( .A(n57443), .B(n46651), .X(n59767) );
  nor_x1_sg U61503 ( .A(n57446), .B(n46652), .X(n59762) );
  nor_x1_sg U61504 ( .A(n57446), .B(n46653), .X(n59757) );
  nor_x1_sg U61505 ( .A(n57443), .B(n46654), .X(n59752) );
  nor_x1_sg U61506 ( .A(n57444), .B(n46655), .X(n59747) );
  nor_x1_sg U61507 ( .A(n57445), .B(n46656), .X(n59742) );
  nor_x1_sg U61508 ( .A(n57446), .B(n46657), .X(n59737) );
  nor_x1_sg U61509 ( .A(n57441), .B(n46658), .X(n59732) );
  nor_x1_sg U61510 ( .A(n57410), .B(n46659), .X(n59727) );
  nor_x1_sg U61511 ( .A(n57396), .B(n46660), .X(n59722) );
  nor_x1_sg U61512 ( .A(n57411), .B(n46661), .X(n59717) );
  nor_x1_sg U61513 ( .A(n57443), .B(n46662), .X(n59712) );
  nor_x1_sg U61514 ( .A(n57443), .B(n46663), .X(n59707) );
  nor_x1_sg U61515 ( .A(n57443), .B(n46664), .X(n59702) );
  nor_x1_sg U61516 ( .A(n57443), .B(n46665), .X(n59697) );
  nor_x1_sg U61517 ( .A(n57394), .B(n46666), .X(n59692) );
  nor_x1_sg U61518 ( .A(n57396), .B(n46667), .X(n59687) );
  nor_x1_sg U61519 ( .A(n57394), .B(n46668), .X(n59682) );
  nor_x1_sg U61520 ( .A(n57444), .B(n46669), .X(n59677) );
  nor_x1_sg U61521 ( .A(n57445), .B(n46670), .X(n59672) );
  nor_x1_sg U61522 ( .A(n57441), .B(n46671), .X(n59667) );
  nor_x1_sg U61523 ( .A(n57445), .B(n46672), .X(n59662) );
  nor_x1_sg U61524 ( .A(n57394), .B(n46673), .X(n59657) );
  nor_x1_sg U61525 ( .A(n57396), .B(n46674), .X(n59652) );
  nor_x1_sg U61526 ( .A(n57441), .B(n46675), .X(n59647) );
  nor_x1_sg U61527 ( .A(n57446), .B(n46676), .X(n59642) );
  nor_x1_sg U61528 ( .A(n57412), .B(n46677), .X(n59637) );
  nor_x1_sg U61529 ( .A(n57445), .B(n46678), .X(n59632) );
  nor_x1_sg U61530 ( .A(n57442), .B(n46679), .X(n59627) );
  nor_x1_sg U61531 ( .A(n57444), .B(n46680), .X(n59622) );
  nor_x1_sg U61532 ( .A(n57444), .B(n46681), .X(n59617) );
  nor_x1_sg U61533 ( .A(n57440), .B(n46682), .X(n59612) );
  nor_x1_sg U61534 ( .A(n57442), .B(n46683), .X(n59607) );
  nor_x1_sg U61535 ( .A(n57441), .B(n46684), .X(n59602) );
  nor_x1_sg U61536 ( .A(n57446), .B(n46685), .X(n59597) );
  nor_x1_sg U61537 ( .A(n57441), .B(n46686), .X(n59592) );
  nor_x1_sg U61538 ( .A(n57445), .B(n46687), .X(n59587) );
  nor_x1_sg U61539 ( .A(n57442), .B(n46688), .X(n59582) );
  nor_x1_sg U61540 ( .A(n57439), .B(n46689), .X(n59577) );
  nor_x1_sg U61541 ( .A(n57397), .B(n46690), .X(n59572) );
  nor_x1_sg U61542 ( .A(n57439), .B(n46691), .X(n59567) );
  nor_x1_sg U61543 ( .A(n57444), .B(n46692), .X(n59562) );
  nor_x1_sg U61544 ( .A(n57443), .B(n46693), .X(n59557) );
  nor_x1_sg U61545 ( .A(n57444), .B(n46694), .X(n59552) );
  nor_x1_sg U61546 ( .A(n57441), .B(n46695), .X(n59547) );
  nor_x1_sg U61547 ( .A(n57440), .B(n46696), .X(n59542) );
  nor_x1_sg U61548 ( .A(n57442), .B(n46697), .X(n59537) );
  nor_x1_sg U61549 ( .A(n57441), .B(n46698), .X(n59532) );
  nor_x1_sg U61550 ( .A(n57444), .B(n46699), .X(n59527) );
  nor_x1_sg U61551 ( .A(n57440), .B(n46700), .X(n59522) );
  nor_x1_sg U61552 ( .A(n57442), .B(n46701), .X(n59517) );
  nor_x1_sg U61553 ( .A(n57446), .B(n46702), .X(n59512) );
  nor_x1_sg U61554 ( .A(n57441), .B(n46703), .X(n59507) );
  nor_x1_sg U61555 ( .A(n57440), .B(n46704), .X(n59502) );
  nor_x1_sg U61556 ( .A(n57445), .B(n46705), .X(n59497) );
  nor_x1_sg U61557 ( .A(n57445), .B(n46706), .X(n59492) );
  nor_x1_sg U61558 ( .A(n57440), .B(n46707), .X(n59487) );
  nor_x1_sg U61559 ( .A(n57442), .B(n46708), .X(n59482) );
  nor_x1_sg U61560 ( .A(n57440), .B(n46709), .X(n59477) );
  nor_x1_sg U61561 ( .A(n57446), .B(n46710), .X(n59472) );
  nor_x1_sg U61562 ( .A(n57441), .B(n46711), .X(n59467) );
  nor_x1_sg U61563 ( .A(n57445), .B(n46712), .X(n59462) );
  nor_x1_sg U61564 ( .A(n57439), .B(n46713), .X(n59457) );
  nor_x1_sg U61565 ( .A(n57411), .B(n46714), .X(n59452) );
  nor_x1_sg U61566 ( .A(n57430), .B(n46715), .X(n59447) );
  nor_x1_sg U61567 ( .A(n57440), .B(n46716), .X(n59442) );
  nor_x1_sg U61568 ( .A(n57397), .B(n46717), .X(n59437) );
  nor_x1_sg U61569 ( .A(n57413), .B(n46718), .X(n59432) );
  nor_x1_sg U61570 ( .A(n57410), .B(n46719), .X(n59427) );
  nor_x1_sg U61571 ( .A(n57411), .B(n46720), .X(n59422) );
  nor_x1_sg U61572 ( .A(n57397), .B(n46721), .X(n59417) );
  nor_x1_sg U61573 ( .A(n57397), .B(n46722), .X(n59412) );
  nor_x1_sg U61574 ( .A(n57397), .B(n46723), .X(n59407) );
  nor_x1_sg U61575 ( .A(n57397), .B(n46724), .X(n59402) );
  nor_x1_sg U61576 ( .A(n57397), .B(n46725), .X(n59397) );
  nor_x1_sg U61577 ( .A(n57397), .B(n46726), .X(n59392) );
  nor_x1_sg U61578 ( .A(n57397), .B(n46727), .X(n59387) );
  nor_x1_sg U61579 ( .A(n57397), .B(n46728), .X(n59382) );
  nor_x1_sg U61580 ( .A(n57397), .B(n46729), .X(n59377) );
  nor_x1_sg U61581 ( .A(n57406), .B(n46730), .X(n59372) );
  nor_x1_sg U61582 ( .A(n57406), .B(n46731), .X(n59367) );
  nor_x1_sg U61583 ( .A(n57407), .B(n46732), .X(n59362) );
  nor_x1_sg U61584 ( .A(n57430), .B(n46733), .X(n59357) );
  nor_x1_sg U61585 ( .A(n57430), .B(n46734), .X(n59352) );
  nor_x1_sg U61586 ( .A(n57410), .B(n46735), .X(n59347) );
  nor_x1_sg U61587 ( .A(n57395), .B(n46736), .X(n59342) );
  nor_x1_sg U61588 ( .A(n57408), .B(n46737), .X(n59337) );
  nor_x1_sg U61589 ( .A(n57409), .B(n46738), .X(n59332) );
  nor_x1_sg U61590 ( .A(n57446), .B(n46739), .X(n59327) );
  nor_x1_sg U61591 ( .A(n57394), .B(n46740), .X(n59322) );
  nor_x1_sg U61592 ( .A(n57444), .B(n46741), .X(n59317) );
  nor_x1_sg U61593 ( .A(n57445), .B(n46742), .X(n59312) );
  nor_x1_sg U61594 ( .A(n57443), .B(n46743), .X(n59307) );
  nor_x1_sg U61595 ( .A(n57441), .B(n46744), .X(n59302) );
  nor_x1_sg U61596 ( .A(n57396), .B(n46745), .X(n59297) );
  nor_x1_sg U61597 ( .A(n57412), .B(n46746), .X(n59292) );
  nor_x1_sg U61598 ( .A(n57413), .B(n46747), .X(n59287) );
  nor_x1_sg U61599 ( .A(n57397), .B(n46748), .X(n59282) );
  nor_x1_sg U61600 ( .A(n57397), .B(n46749), .X(n59277) );
  nor_x1_sg U61601 ( .A(n57397), .B(n46750), .X(n59272) );
  nor_x1_sg U61602 ( .A(n57397), .B(n46751), .X(n59267) );
  nor_x1_sg U61603 ( .A(n57397), .B(n46752), .X(n59262) );
  nor_x1_sg U61604 ( .A(n57397), .B(n46753), .X(n59257) );
  nor_x1_sg U61605 ( .A(n57397), .B(n46754), .X(n59252) );
  nor_x1_sg U61606 ( .A(n57397), .B(n46755), .X(n59247) );
  nor_x1_sg U61607 ( .A(n57397), .B(n46756), .X(n59242) );
  nor_x1_sg U61608 ( .A(n57396), .B(n46757), .X(n59237) );
  nor_x1_sg U61609 ( .A(n57396), .B(n46758), .X(n59232) );
  nor_x1_sg U61610 ( .A(n57396), .B(n46759), .X(n59227) );
  nor_x1_sg U61611 ( .A(n57396), .B(n46760), .X(n59222) );
  nor_x1_sg U61612 ( .A(n57396), .B(n46761), .X(n59217) );
  nor_x1_sg U61613 ( .A(n57396), .B(n46762), .X(n59212) );
  nor_x1_sg U61614 ( .A(n57396), .B(n46763), .X(n59207) );
  nor_x1_sg U61615 ( .A(n57396), .B(n46764), .X(n59202) );
  nor_x1_sg U61616 ( .A(n57396), .B(n46765), .X(n59197) );
  nor_x1_sg U61617 ( .A(n57444), .B(n46766), .X(n59192) );
  nor_x1_sg U61618 ( .A(n57396), .B(n46767), .X(n59187) );
  nor_x1_sg U61619 ( .A(n57440), .B(n46768), .X(n59182) );
  nor_x1_sg U61620 ( .A(n57444), .B(n46769), .X(n59177) );
  nor_x1_sg U61621 ( .A(n57445), .B(n46770), .X(n59172) );
  nor_x1_sg U61622 ( .A(n57439), .B(n46771), .X(n59167) );
  nor_x1_sg U61623 ( .A(n57439), .B(n46772), .X(n59162) );
  nor_x1_sg U61624 ( .A(n57441), .B(n46773), .X(n59157) );
  nor_x1_sg U61625 ( .A(n57444), .B(n46774), .X(n59152) );
  nor_x1_sg U61626 ( .A(n57446), .B(n46775), .X(n59147) );
  nor_x1_sg U61627 ( .A(n57412), .B(n46776), .X(n59142) );
  nor_x1_sg U61628 ( .A(n57413), .B(n46777), .X(n59137) );
  nor_x1_sg U61629 ( .A(n57410), .B(n46778), .X(n59132) );
  nor_x1_sg U61630 ( .A(n57411), .B(n46779), .X(n59127) );
  nor_x1_sg U61631 ( .A(n57442), .B(n46780), .X(n59122) );
  nor_x1_sg U61632 ( .A(n57443), .B(n46781), .X(n59117) );
  nor_x1_sg U61633 ( .A(n57394), .B(n46782), .X(n59112) );
  nor_x1_sg U61634 ( .A(n57446), .B(n46783), .X(n59107) );
  nor_x1_sg U61635 ( .A(n57443), .B(n46784), .X(n59102) );
  nor_x1_sg U61636 ( .A(n57442), .B(n46785), .X(n59097) );
  nor_x1_sg U61637 ( .A(n57443), .B(n46786), .X(n59092) );
  nor_x1_sg U61638 ( .A(n57444), .B(n46787), .X(n59087) );
  nor_x1_sg U61639 ( .A(n57445), .B(n46788), .X(n59082) );
  nor_x1_sg U61640 ( .A(n57446), .B(n46789), .X(n59077) );
  nor_x1_sg U61641 ( .A(n57394), .B(n46790), .X(n59072) );
  nor_x1_sg U61642 ( .A(n57442), .B(n46791), .X(n59067) );
  nor_x1_sg U61643 ( .A(n57443), .B(n46792), .X(n59062) );
  nor_x1_sg U61644 ( .A(n57394), .B(n46793), .X(n59057) );
  nor_x1_sg U61645 ( .A(n57439), .B(n46794), .X(n59052) );
  nor_x1_sg U61646 ( .A(n57439), .B(n46795), .X(n59047) );
  nor_x1_sg U61647 ( .A(n57441), .B(n46796), .X(n59042) );
  nor_x1_sg U61648 ( .A(n57440), .B(n46797), .X(n59037) );
  nor_x1_sg U61649 ( .A(n57445), .B(n46798), .X(n59032) );
  nor_x1_sg U61650 ( .A(n57443), .B(n46799), .X(n59027) );
  nor_x1_sg U61651 ( .A(n57446), .B(n46800), .X(n59022) );
  nor_x1_sg U61652 ( .A(n57407), .B(n46801), .X(n59017) );
  nor_x1_sg U61653 ( .A(n57440), .B(n46802), .X(n59012) );
  nor_x1_sg U61654 ( .A(n57397), .B(n46803), .X(n59007) );
  nor_x1_sg U61655 ( .A(n57430), .B(n46804), .X(n59002) );
  nor_x1_sg U61656 ( .A(n57412), .B(n46805), .X(n58997) );
  nor_x1_sg U61657 ( .A(n57411), .B(n46806), .X(n58992) );
  nor_x1_sg U61658 ( .A(n57446), .B(n46807), .X(n58987) );
  nor_x1_sg U61659 ( .A(n61858), .B(n46808), .X(n58982) );
  nor_x1_sg U61660 ( .A(n61858), .B(n46809), .X(n58977) );
  nor_x1_sg U61661 ( .A(n57395), .B(n46810), .X(n58972) );
  nor_x1_sg U61662 ( .A(n57395), .B(n46811), .X(n58967) );
  nor_x1_sg U61663 ( .A(n57395), .B(n46812), .X(n58962) );
  nor_x1_sg U61664 ( .A(n57395), .B(n46813), .X(n58957) );
  nor_x1_sg U61665 ( .A(n57395), .B(n46814), .X(n58952) );
  nor_x1_sg U61666 ( .A(n57395), .B(n46815), .X(n58947) );
  nor_x1_sg U61667 ( .A(n57395), .B(n46816), .X(n58942) );
  nor_x1_sg U61668 ( .A(n57395), .B(n46817), .X(n58937) );
  nor_x1_sg U61669 ( .A(n57395), .B(n46818), .X(n58932) );
  nor_x1_sg U61670 ( .A(n57394), .B(n46819), .X(n58927) );
  nor_x1_sg U61671 ( .A(n57396), .B(n46820), .X(n58922) );
  nor_x1_sg U61672 ( .A(n57439), .B(n46821), .X(n58917) );
  nor_x1_sg U61673 ( .A(n57440), .B(n46822), .X(n58912) );
  nor_x1_sg U61674 ( .A(n57394), .B(n46823), .X(n58907) );
  nor_x1_sg U61675 ( .A(n57397), .B(n46824), .X(n58902) );
  nor_x1_sg U61676 ( .A(n57396), .B(n46825), .X(n58897) );
  nor_x1_sg U61677 ( .A(n57444), .B(n46826), .X(n58892) );
  nor_x1_sg U61678 ( .A(n57442), .B(n46827), .X(n58887) );
  nor_x1_sg U61679 ( .A(n57394), .B(n46828), .X(n58882) );
  nor_x1_sg U61680 ( .A(n57444), .B(n46829), .X(n58877) );
  nor_x1_sg U61681 ( .A(n57396), .B(n46830), .X(n58872) );
  nor_x1_sg U61682 ( .A(n57396), .B(n46831), .X(n58867) );
  nor_x1_sg U61683 ( .A(n57445), .B(n46832), .X(n58862) );
  nor_x1_sg U61684 ( .A(n57394), .B(n46833), .X(n58857) );
  nor_x1_sg U61685 ( .A(n57446), .B(n46834), .X(n58852) );
  nor_x1_sg U61686 ( .A(n57396), .B(n46835), .X(n58847) );
  nor_x1_sg U61687 ( .A(n57441), .B(n46836), .X(n58842) );
  nor_x1_sg U61688 ( .A(n57396), .B(n46837), .X(n58837) );
  nor_x1_sg U61689 ( .A(n57445), .B(n46838), .X(n58832) );
  nor_x1_sg U61690 ( .A(n57396), .B(n46839), .X(n58827) );
  nor_x1_sg U61691 ( .A(n57441), .B(n46840), .X(n58822) );
  nor_x1_sg U61692 ( .A(n57396), .B(n46841), .X(n58817) );
  nor_x1_sg U61693 ( .A(n57397), .B(n46842), .X(n58812) );
  nor_x1_sg U61694 ( .A(n57439), .B(n46843), .X(n58807) );
  nor_x1_sg U61695 ( .A(n57439), .B(n46844), .X(n58802) );
  nor_x1_sg U61696 ( .A(n57396), .B(n46845), .X(n58797) );
  nor_x1_sg U61697 ( .A(n57394), .B(n46846), .X(n58792) );
  nor_x1_sg U61698 ( .A(n57394), .B(n46847), .X(n58787) );
  nor_x1_sg U61699 ( .A(n57394), .B(n46848), .X(n58782) );
  nor_x1_sg U61700 ( .A(n57394), .B(n46849), .X(n58777) );
  nor_x1_sg U61701 ( .A(n57394), .B(n46850), .X(n58772) );
  nor_x1_sg U61702 ( .A(n57394), .B(n46851), .X(n58767) );
  nor_x1_sg U61703 ( .A(n57394), .B(n46852), .X(n58762) );
  nor_x1_sg U61704 ( .A(n32044), .B(n32045), .X(n32043) );
  nor_x1_sg U61705 ( .A(n31978), .B(n68574), .X(n31977) );
  nor_x1_sg U61706 ( .A(n31979), .B(n31973), .X(n31976) );
  nor_x1_sg U61707 ( .A(n31978), .B(n68576), .X(n32062) );
  nor_x1_sg U61708 ( .A(n31998), .B(n31979), .X(n32061) );
  nor_x1_sg U61709 ( .A(n26288), .B(n57308), .X(n26287) );
  nand_x2_sg U61710 ( .A(n26293), .B(n26294), .X(n26289) );
  nand_x2_sg U61711 ( .A(n32483), .B(n68268), .X(n32482) );
  nor_x1_sg U61712 ( .A(n32487), .B(n32488), .X(n32486) );
  nor_x1_sg U61713 ( .A(n32377), .B(n68396), .X(n32376) );
  nor_x1_sg U61714 ( .A(n32378), .B(n32371), .X(n32375) );
  nor_x1_sg U61715 ( .A(n57446), .B(n46853), .X(n58662) );
  nor_x1_sg U61716 ( .A(n26311), .B(n26312), .X(n26310) );
  nand_x2_sg U61717 ( .A(n26315), .B(n26316), .X(n26311) );
  nand_x2_sg U61718 ( .A(n26313), .B(n26314), .X(n26312) );
  nand_x1_sg U61719 ( .A(n67534), .B(n26322), .X(n26320) );
  nor_x1_sg U61720 ( .A(n26328), .B(n26329), .X(n26323) );
  nor_x1_sg U61721 ( .A(n61907), .B(n57962), .X(n57959) );
  nor_x1_sg U61722 ( .A(n47317), .B(n57963), .X(n57965) );
  nand_x1_sg U61723 ( .A(n30627), .B(n61907), .X(n57957) );
  nor_x1_sg U61724 ( .A(n30624), .B(n47317), .X(n57958) );
  nor_x1_sg U61725 ( .A(n61911), .B(n57962), .X(n57961) );
  nor_x1_sg U61726 ( .A(n47299), .B(n38412), .X(n45553) );
  nor_x1_sg U61727 ( .A(n68373), .B(n68374), .X(\filter_0/N1845 ) );
  nand_x4_sg U61728 ( .A(n58612), .B(n61905), .X(n68268) );
  nand_x2_sg U61729 ( .A(n32558), .B(n32559), .X(n32553) );
  nand_x2_sg U61730 ( .A(n32113), .B(n32114), .X(n32108) );
  nor_x1_sg U61731 ( .A(n32287), .B(n32288), .X(n32277) );
  nor_x1_sg U61732 ( .A(n32279), .B(n32280), .X(n32278) );
  nor_x1_sg U61733 ( .A(n32732), .B(n32733), .X(n32722) );
  nor_x1_sg U61734 ( .A(n32724), .B(n32725), .X(n32723) );
  nand_x2_sg U61735 ( .A(n32596), .B(n32597), .X(n32591) );
  nand_x2_sg U61736 ( .A(n32151), .B(n32152), .X(n32146) );
  nand_x2_sg U61737 ( .A(n32131), .B(n32132), .X(n32126) );
  nand_x2_sg U61738 ( .A(n32576), .B(n32577), .X(n32571) );
  nand_x4_sg U61739 ( .A(n32175), .B(n32176), .X(n31966) );
  nor_x1_sg U61740 ( .A(n32185), .B(n32186), .X(n32175) );
  nor_x1_sg U61741 ( .A(n32177), .B(n32178), .X(n32176) );
  nand_x2_sg U61742 ( .A(n32190), .B(n32191), .X(n32185) );
  nand_x4_sg U61743 ( .A(n32620), .B(n32621), .X(n32433) );
  nor_x1_sg U61744 ( .A(n32630), .B(n32631), .X(n32620) );
  nor_x1_sg U61745 ( .A(n32622), .B(n32623), .X(n32621) );
  nand_x2_sg U61746 ( .A(n32635), .B(n32636), .X(n32630) );
  nand_x4_sg U61747 ( .A(n32703), .B(n32704), .X(n32533) );
  nor_x1_sg U61748 ( .A(n32713), .B(n32714), .X(n32703) );
  nor_x1_sg U61749 ( .A(n32705), .B(n32706), .X(n32704) );
  nand_x2_sg U61750 ( .A(n32718), .B(n32719), .X(n32713) );
  nand_x4_sg U61751 ( .A(n32258), .B(n32259), .X(n32088) );
  nor_x1_sg U61752 ( .A(n32268), .B(n32269), .X(n32258) );
  nor_x1_sg U61753 ( .A(n32260), .B(n32261), .X(n32259) );
  nand_x2_sg U61754 ( .A(n32273), .B(n32274), .X(n32268) );
  nand_x1_sg U61755 ( .A(n57929), .B(n61909), .X(n57970) );
  nor_x1_sg U61756 ( .A(n57927), .B(n58612), .X(n57969) );
  nand_x4_sg U61757 ( .A(n32667), .B(n32668), .X(n32524) );
  nor_x1_sg U61758 ( .A(n32677), .B(n32678), .X(n32667) );
  nor_x1_sg U61759 ( .A(n32669), .B(n32670), .X(n32668) );
  nand_x2_sg U61760 ( .A(n32682), .B(n32683), .X(n32677) );
  nand_x4_sg U61761 ( .A(n32222), .B(n32223), .X(n32079) );
  nor_x1_sg U61762 ( .A(n32232), .B(n32233), .X(n32222) );
  nor_x1_sg U61763 ( .A(n32224), .B(n32225), .X(n32223) );
  nand_x2_sg U61764 ( .A(n32237), .B(n32238), .X(n32232) );
  nor_x1_sg U61765 ( .A(n32695), .B(n32696), .X(n32685) );
  nor_x1_sg U61766 ( .A(n32687), .B(n32688), .X(n32686) );
  nand_x2_sg U61767 ( .A(n32700), .B(n32701), .X(n32695) );
  nor_x1_sg U61768 ( .A(n32250), .B(n32251), .X(n32240) );
  nor_x1_sg U61769 ( .A(n32242), .B(n32243), .X(n32241) );
  nand_x2_sg U61770 ( .A(n32255), .B(n32256), .X(n32250) );
  nand_x4_sg U61771 ( .A(n32316), .B(n32317), .X(n32078) );
  nor_x1_sg U61772 ( .A(n32326), .B(n32327), .X(n32316) );
  nor_x1_sg U61773 ( .A(n32318), .B(n32319), .X(n32317) );
  nand_x2_sg U61774 ( .A(n32331), .B(n32332), .X(n32326) );
  nand_x4_sg U61775 ( .A(n32761), .B(n32762), .X(n32523) );
  nor_x1_sg U61776 ( .A(n32771), .B(n32772), .X(n32761) );
  nor_x1_sg U61777 ( .A(n32763), .B(n32764), .X(n32762) );
  nand_x2_sg U61778 ( .A(n32776), .B(n32777), .X(n32771) );
  nor_x1_sg U61779 ( .A(n32308), .B(n32309), .X(n32298) );
  nor_x1_sg U61780 ( .A(n32300), .B(n32301), .X(n32299) );
  nand_x2_sg U61781 ( .A(n32313), .B(n32314), .X(n32308) );
  nor_x1_sg U61782 ( .A(n32753), .B(n32754), .X(n32743) );
  nor_x1_sg U61783 ( .A(n32745), .B(n32746), .X(n32744) );
  nand_x2_sg U61784 ( .A(n32758), .B(n32759), .X(n32753) );
  nand_x2_sg U61785 ( .A(n32169), .B(n32170), .X(n32164) );
  nand_x2_sg U61786 ( .A(n32614), .B(n32615), .X(n32609) );
  nand_x4_sg U61787 ( .A(n32335), .B(n32336), .X(n32089) );
  nor_x1_sg U61788 ( .A(n32345), .B(n32346), .X(n32335) );
  nor_x1_sg U61789 ( .A(n32337), .B(n32338), .X(n32336) );
  nand_x2_sg U61790 ( .A(n32350), .B(n32351), .X(n32345) );
  nand_x4_sg U61791 ( .A(n32780), .B(n32781), .X(n32534) );
  nor_x1_sg U61792 ( .A(n32790), .B(n32791), .X(n32780) );
  nor_x1_sg U61793 ( .A(n32782), .B(n32783), .X(n32781) );
  nand_x2_sg U61794 ( .A(n32795), .B(n32796), .X(n32790) );
  nand_x4_sg U61795 ( .A(n32193), .B(n32194), .X(n31961) );
  nor_x1_sg U61796 ( .A(n32203), .B(n32204), .X(n32193) );
  nor_x1_sg U61797 ( .A(n32195), .B(n32196), .X(n32194) );
  nand_x2_sg U61798 ( .A(n32208), .B(n32209), .X(n32203) );
  nand_x4_sg U61799 ( .A(n32638), .B(n32639), .X(n32428) );
  nor_x1_sg U61800 ( .A(n32648), .B(n32649), .X(n32638) );
  nor_x1_sg U61801 ( .A(n32640), .B(n32641), .X(n32639) );
  nand_x2_sg U61802 ( .A(n32653), .B(n32654), .X(n32648) );
  nor_x1_sg U61803 ( .A(n68369), .B(n35837), .X(n44271) );
  nor_x1_sg U61804 ( .A(n32012), .B(n32013), .X(n32002) );
  nor_x1_sg U61805 ( .A(n32004), .B(n32005), .X(n32003) );
  nand_x2_sg U61806 ( .A(n32017), .B(n32018), .X(n32012) );
  nor_x1_sg U61807 ( .A(n32454), .B(n32455), .X(n32444) );
  nor_x1_sg U61808 ( .A(n32446), .B(n32447), .X(n32445) );
  nand_x2_sg U61809 ( .A(n32459), .B(n32460), .X(n32454) );
  nand_x1_sg U61810 ( .A(n35839), .B(n68370), .X(n39702) );
  nand_x2_sg U61811 ( .A(n68271), .B(n61906), .X(n38416) );
  nand_x2_sg U61812 ( .A(n22469), .B(n22470), .X(n22468) );
  nand_x1_sg U61813 ( .A(n22471), .B(n58585), .X(n22470) );
  nand_x1_sg U61814 ( .A(n57463), .B(n68573), .X(n22469) );
  nand_x2_sg U61815 ( .A(n57859), .B(n22520), .X(n22519) );
  nand_x1_sg U61816 ( .A(n22521), .B(n22522), .X(n22520) );
  nand_x1_sg U61817 ( .A(n23308), .B(n68571), .X(n24266) );
  nor_x1_sg U61818 ( .A(n68576), .B(n68571), .X(n22570) );
  nor_x1_sg U61819 ( .A(n68576), .B(n68574), .X(n22621) );
  nor_x1_sg U61820 ( .A(n23308), .B(n24049), .X(n24047) );
  nand_x2_sg U61821 ( .A(n22495), .B(n22496), .X(n22494) );
  nand_x1_sg U61822 ( .A(n22497), .B(n58585), .X(n22496) );
  nand_x1_sg U61823 ( .A(n57463), .B(n68391), .X(n22495) );
  nand_x2_sg U61824 ( .A(n57861), .B(n22545), .X(n22544) );
  nand_x1_sg U61825 ( .A(n22546), .B(n22522), .X(n22545) );
  nor_x1_sg U61826 ( .A(n68397), .B(n68396), .X(n22648) );
  nor_x1_sg U61827 ( .A(n33738), .B(n67528), .X(n26065) );
  nor_x1_sg U61828 ( .A(n34219), .B(n67525), .X(n26161) );
  nor_x1_sg U61829 ( .A(n57113), .B(n67530), .X(\filter_0/n8271 ) );
  nand_x1_sg U61830 ( .A(n26085), .B(n67560), .X(n26127) );
  nor_x1_sg U61831 ( .A(n26129), .B(n26130), .X(n26128) );
  nand_x2_sg U61832 ( .A(n26133), .B(n26134), .X(n26129) );
  nand_x1_sg U61833 ( .A(n26085), .B(n67554), .X(n26084) );
  nor_x1_sg U61834 ( .A(n26087), .B(n26088), .X(n26086) );
  nand_x2_sg U61835 ( .A(n26093), .B(n26094), .X(n26087) );
  nand_x1_sg U61836 ( .A(n26085), .B(n67548), .X(n26219) );
  nor_x1_sg U61837 ( .A(n26221), .B(n26222), .X(n26220) );
  nand_x2_sg U61838 ( .A(n26225), .B(n26226), .X(n26221) );
  nand_x1_sg U61839 ( .A(n26085), .B(n67542), .X(n26185) );
  nor_x1_sg U61840 ( .A(n26187), .B(n26188), .X(n26186) );
  nand_x2_sg U61841 ( .A(n26191), .B(n26192), .X(n26187) );
  nand_x2_sg U61842 ( .A(n23305), .B(n23306), .X(n23304) );
  nand_x1_sg U61843 ( .A(n29337), .B(n57917), .X(n23305) );
  nand_x1_sg U61844 ( .A(n58616), .B(n58473), .X(n23306) );
  nand_x2_sg U61845 ( .A(n22973), .B(n22521), .X(n22972) );
  nor_x1_sg U61846 ( .A(n57298), .B(n22974), .X(n22973) );
  nand_x2_sg U61847 ( .A(n23200), .B(n22546), .X(n23199) );
  nor_x1_sg U61848 ( .A(n57304), .B(n22974), .X(n23200) );
  nand_x2_sg U61849 ( .A(n24164), .B(n24817), .X(n24816) );
  nand_x2_sg U61850 ( .A(n24169), .B(n24849), .X(n24848) );
  nand_x2_sg U61851 ( .A(n24174), .B(n24879), .X(n24878) );
  nand_x2_sg U61852 ( .A(n24179), .B(n24909), .X(n24908) );
  nand_x2_sg U61853 ( .A(n24184), .B(n24939), .X(n24938) );
  nand_x2_sg U61854 ( .A(n24189), .B(n24969), .X(n24968) );
  nand_x2_sg U61855 ( .A(n24194), .B(n24999), .X(n24998) );
  nand_x2_sg U61856 ( .A(n24199), .B(n25029), .X(n25028) );
  nand_x2_sg U61857 ( .A(n24204), .B(n25059), .X(n25058) );
  nand_x2_sg U61858 ( .A(n24209), .B(n25089), .X(n25088) );
  nand_x2_sg U61859 ( .A(n24214), .B(n25119), .X(n25118) );
  nand_x2_sg U61860 ( .A(n24219), .B(n25149), .X(n25148) );
  nand_x2_sg U61861 ( .A(n24224), .B(n25179), .X(n25178) );
  nand_x2_sg U61862 ( .A(n24229), .B(n25209), .X(n25208) );
  nand_x2_sg U61863 ( .A(n24244), .B(n25299), .X(n25298) );
  nand_x2_sg U61864 ( .A(n24249), .B(n25329), .X(n25328) );
  nand_x2_sg U61865 ( .A(n24254), .B(n25359), .X(n25358) );
  nand_x2_sg U61866 ( .A(n24267), .B(n25390), .X(n25389) );
  nand_x2_sg U61867 ( .A(n24273), .B(n25421), .X(n25420) );
  nand_x2_sg U61868 ( .A(n24278), .B(n25451), .X(n25450) );
  nand_x2_sg U61869 ( .A(n24283), .B(n25481), .X(n25480) );
  nand_x2_sg U61870 ( .A(n24288), .B(n25511), .X(n25510) );
  nand_x2_sg U61871 ( .A(n24293), .B(n25541), .X(n25540) );
  nand_x2_sg U61872 ( .A(n24298), .B(n25571), .X(n25570) );
  nand_x2_sg U61873 ( .A(n24303), .B(n25601), .X(n25600) );
  nand_x2_sg U61874 ( .A(n24308), .B(n25631), .X(n25630) );
  nand_x2_sg U61875 ( .A(n24313), .B(n25661), .X(n25660) );
  nand_x2_sg U61876 ( .A(n24318), .B(n25691), .X(n25690) );
  nand_x2_sg U61877 ( .A(n24323), .B(n25721), .X(n25720) );
  nand_x2_sg U61878 ( .A(n24333), .B(n25781), .X(n25780) );
  nand_x2_sg U61879 ( .A(n24338), .B(n25811), .X(n25810) );
  nand_x2_sg U61880 ( .A(n24343), .B(n25841), .X(n25840) );
  nand_x2_sg U61881 ( .A(n24348), .B(n25871), .X(n25870) );
  nand_x2_sg U61882 ( .A(n24353), .B(n25901), .X(n25900) );
  nand_x2_sg U61883 ( .A(n24358), .B(n25931), .X(n25930) );
  nand_x2_sg U61884 ( .A(n24363), .B(n25961), .X(n25960) );
  nand_x4_sg U61885 ( .A(n26052), .B(n26055), .X(n26053) );
  nand_x1_sg U61886 ( .A(n67530), .B(n57307), .X(n26055) );
  nand_x2_sg U61887 ( .A(n24263), .B(n24264), .X(n24262) );
  nand_x1_sg U61888 ( .A(n24265), .B(n23308), .X(n24264) );
  nand_x4_sg U61889 ( .A(n57459), .B(n23945), .X(n24164) );
  nand_x4_sg U61890 ( .A(n57459), .B(n23951), .X(n24169) );
  nand_x4_sg U61891 ( .A(n57459), .B(n23956), .X(n24174) );
  nand_x4_sg U61892 ( .A(n57459), .B(n23961), .X(n24179) );
  nand_x4_sg U61893 ( .A(n57459), .B(n23966), .X(n24184) );
  nand_x4_sg U61894 ( .A(n57459), .B(n23971), .X(n24189) );
  nand_x4_sg U61895 ( .A(n57459), .B(n23976), .X(n24194) );
  nand_x4_sg U61896 ( .A(n57459), .B(n23981), .X(n24199) );
  nand_x4_sg U61897 ( .A(n57459), .B(n23986), .X(n24204) );
  nand_x4_sg U61898 ( .A(n57459), .B(n23991), .X(n24209) );
  nand_x4_sg U61899 ( .A(n57459), .B(n23996), .X(n24214) );
  nand_x4_sg U61900 ( .A(n57459), .B(n24001), .X(n24219) );
  nand_x4_sg U61901 ( .A(n57459), .B(n24006), .X(n24224) );
  nand_x4_sg U61902 ( .A(n57459), .B(n24011), .X(n24229) );
  nand_x4_sg U61903 ( .A(n57459), .B(n24016), .X(n24234) );
  nand_x4_sg U61904 ( .A(n57459), .B(n24021), .X(n24239) );
  nand_x4_sg U61905 ( .A(n57459), .B(n24026), .X(n24244) );
  nand_x4_sg U61906 ( .A(n57459), .B(n24031), .X(n24249) );
  nand_x4_sg U61907 ( .A(n57459), .B(n24036), .X(n24254) );
  nand_x4_sg U61908 ( .A(n57459), .B(n24041), .X(n24267) );
  nand_x4_sg U61909 ( .A(n57459), .B(n24055), .X(n24273) );
  nand_x4_sg U61910 ( .A(n57459), .B(n24061), .X(n24278) );
  nand_x4_sg U61911 ( .A(n57459), .B(n24066), .X(n24283) );
  nand_x4_sg U61912 ( .A(n57459), .B(n24071), .X(n24288) );
  nand_x4_sg U61913 ( .A(n57459), .B(n24076), .X(n24293) );
  nand_x4_sg U61914 ( .A(n57459), .B(n24081), .X(n24298) );
  nand_x4_sg U61915 ( .A(n57459), .B(n24086), .X(n24303) );
  nand_x4_sg U61916 ( .A(n57459), .B(n24091), .X(n24308) );
  nand_x4_sg U61917 ( .A(n57459), .B(n24096), .X(n24313) );
  nand_x4_sg U61918 ( .A(n57459), .B(n24101), .X(n24318) );
  nand_x4_sg U61919 ( .A(n57459), .B(n24106), .X(n24323) );
  nand_x4_sg U61920 ( .A(n57459), .B(n24111), .X(n24328) );
  nand_x4_sg U61921 ( .A(n57459), .B(n24116), .X(n24333) );
  nand_x4_sg U61922 ( .A(n57459), .B(n24121), .X(n24338) );
  nand_x4_sg U61923 ( .A(n57459), .B(n24126), .X(n24343) );
  nand_x4_sg U61924 ( .A(n57459), .B(n24131), .X(n24348) );
  nand_x4_sg U61925 ( .A(n57459), .B(n24136), .X(n24353) );
  nand_x4_sg U61926 ( .A(n57459), .B(n24141), .X(n24358) );
  nand_x4_sg U61927 ( .A(n57459), .B(n24146), .X(n24363) );
  nand_x4_sg U61928 ( .A(n57459), .B(n24151), .X(n24376) );
  nand_x2_sg U61929 ( .A(n22743), .B(n22744), .X(n22742) );
  nand_x1_sg U61930 ( .A(n22745), .B(n22497), .X(n22744) );
  nand_x1_sg U61931 ( .A(n57862), .B(n68391), .X(n22743) );
  nand_x2_sg U61932 ( .A(n67096), .B(n57924), .X(n58382) );
  nand_x2_sg U61933 ( .A(n24481), .B(n24482), .X(n24480) );
  nand_x1_sg U61934 ( .A(n24479), .B(n57296), .X(n24482) );
  nand_x2_sg U61935 ( .A(n24593), .B(n24594), .X(n24592) );
  nand_x1_sg U61936 ( .A(n58132), .B(n58129), .X(n24593) );
  nand_x1_sg U61937 ( .A(n24591), .B(n57296), .X(n24594) );
  nand_x2_sg U61938 ( .A(n67500), .B(n57924), .X(n58377) );
  nand_x4_sg U61939 ( .A(n24815), .B(n67281), .X(n24792) );
  nor_x1_sg U61940 ( .A(n24827), .B(n67293), .X(n24815) );
  nand_x4_sg U61941 ( .A(n24847), .B(n67280), .X(n24831) );
  nor_x1_sg U61942 ( .A(n24858), .B(n67292), .X(n24847) );
  nand_x4_sg U61943 ( .A(n24877), .B(n67279), .X(n24861) );
  nor_x1_sg U61944 ( .A(n24888), .B(n67291), .X(n24877) );
  nand_x4_sg U61945 ( .A(n24907), .B(n67278), .X(n24891) );
  nor_x1_sg U61946 ( .A(n24918), .B(n24919), .X(n24907) );
  nand_x4_sg U61947 ( .A(n24937), .B(n67277), .X(n24921) );
  nor_x1_sg U61948 ( .A(n24948), .B(n24949), .X(n24937) );
  nand_x4_sg U61949 ( .A(n24967), .B(n67276), .X(n24951) );
  nor_x1_sg U61950 ( .A(n24978), .B(n67290), .X(n24967) );
  nand_x4_sg U61951 ( .A(n24997), .B(n67275), .X(n24981) );
  nor_x1_sg U61952 ( .A(n25008), .B(n67289), .X(n24997) );
  nand_x4_sg U61953 ( .A(n25027), .B(n67274), .X(n25011) );
  nor_x1_sg U61954 ( .A(n25038), .B(n67288), .X(n25027) );
  nand_x4_sg U61955 ( .A(n25057), .B(n67273), .X(n25041) );
  nor_x1_sg U61956 ( .A(n25068), .B(n25069), .X(n25057) );
  nand_x4_sg U61957 ( .A(n25087), .B(n67272), .X(n25071) );
  nor_x1_sg U61958 ( .A(n25098), .B(n25099), .X(n25087) );
  nand_x4_sg U61959 ( .A(n25117), .B(n67271), .X(n25101) );
  nor_x1_sg U61960 ( .A(n25128), .B(n67287), .X(n25117) );
  nand_x4_sg U61961 ( .A(n25147), .B(n67270), .X(n25131) );
  nor_x1_sg U61962 ( .A(n25158), .B(n67286), .X(n25147) );
  nand_x4_sg U61963 ( .A(n25177), .B(n67269), .X(n25161) );
  nor_x1_sg U61964 ( .A(n25188), .B(n25189), .X(n25177) );
  nand_x4_sg U61965 ( .A(n25207), .B(n67268), .X(n25191) );
  nor_x1_sg U61966 ( .A(n25218), .B(n25219), .X(n25207) );
  nand_x4_sg U61967 ( .A(n25237), .B(n47395), .X(n25221) );
  nor_x1_sg U61968 ( .A(n25248), .B(n67285), .X(n25237) );
  nand_x4_sg U61969 ( .A(n25267), .B(n47333), .X(n25251) );
  nor_x1_sg U61970 ( .A(n25278), .B(n67284), .X(n25267) );
  nand_x4_sg U61971 ( .A(n25297), .B(n67265), .X(n25281) );
  nor_x1_sg U61972 ( .A(n25308), .B(n67283), .X(n25297) );
  nand_x4_sg U61973 ( .A(n25327), .B(n67264), .X(n25311) );
  nor_x1_sg U61974 ( .A(n25338), .B(n25339), .X(n25327) );
  nand_x4_sg U61975 ( .A(n25357), .B(n67263), .X(n25341) );
  nor_x1_sg U61976 ( .A(n25368), .B(n25369), .X(n25357) );
  nand_x4_sg U61977 ( .A(n25388), .B(n67262), .X(n25371) );
  nor_x1_sg U61978 ( .A(n25399), .B(n67282), .X(n25388) );
  nand_x4_sg U61979 ( .A(n25419), .B(n67474), .X(n25403) );
  nor_x1_sg U61980 ( .A(n25430), .B(n67486), .X(n25419) );
  nand_x4_sg U61981 ( .A(n25449), .B(n67473), .X(n25433) );
  nor_x1_sg U61982 ( .A(n25460), .B(n67485), .X(n25449) );
  nand_x4_sg U61983 ( .A(n25479), .B(n67472), .X(n25463) );
  nor_x1_sg U61984 ( .A(n25490), .B(n67484), .X(n25479) );
  nand_x4_sg U61985 ( .A(n25509), .B(n67471), .X(n25493) );
  nor_x1_sg U61986 ( .A(n25520), .B(n25521), .X(n25509) );
  nand_x4_sg U61987 ( .A(n25539), .B(n67470), .X(n25523) );
  nor_x1_sg U61988 ( .A(n25550), .B(n25551), .X(n25539) );
  nand_x4_sg U61989 ( .A(n25569), .B(n67469), .X(n25553) );
  nor_x1_sg U61990 ( .A(n25580), .B(n67483), .X(n25569) );
  nand_x4_sg U61991 ( .A(n25599), .B(n67468), .X(n25583) );
  nor_x1_sg U61992 ( .A(n25610), .B(n67482), .X(n25599) );
  nand_x4_sg U61993 ( .A(n25629), .B(n67467), .X(n25613) );
  nor_x1_sg U61994 ( .A(n25640), .B(n67481), .X(n25629) );
  nand_x4_sg U61995 ( .A(n25659), .B(n67466), .X(n25643) );
  nor_x1_sg U61996 ( .A(n25670), .B(n25671), .X(n25659) );
  nand_x4_sg U61997 ( .A(n25689), .B(n67465), .X(n25673) );
  nor_x1_sg U61998 ( .A(n25700), .B(n25701), .X(n25689) );
  nand_x4_sg U61999 ( .A(n25719), .B(n67464), .X(n25703) );
  nor_x1_sg U62000 ( .A(n25730), .B(n67480), .X(n25719) );
  nand_x4_sg U62001 ( .A(n25749), .B(n47394), .X(n25733) );
  nor_x1_sg U62002 ( .A(n25760), .B(n67479), .X(n25749) );
  nand_x4_sg U62003 ( .A(n25779), .B(n67462), .X(n25763) );
  nor_x1_sg U62004 ( .A(n25790), .B(n25791), .X(n25779) );
  nand_x4_sg U62005 ( .A(n25809), .B(n67461), .X(n25793) );
  nor_x1_sg U62006 ( .A(n25820), .B(n25821), .X(n25809) );
  nand_x4_sg U62007 ( .A(n25839), .B(n67460), .X(n25823) );
  nor_x1_sg U62008 ( .A(n25850), .B(n67478), .X(n25839) );
  nand_x4_sg U62009 ( .A(n25869), .B(n67459), .X(n25853) );
  nor_x1_sg U62010 ( .A(n25880), .B(n67477), .X(n25869) );
  nand_x4_sg U62011 ( .A(n25899), .B(n67458), .X(n25883) );
  nor_x1_sg U62012 ( .A(n25910), .B(n67476), .X(n25899) );
  nand_x4_sg U62013 ( .A(n25929), .B(n67457), .X(n25913) );
  nor_x1_sg U62014 ( .A(n25940), .B(n25941), .X(n25929) );
  nand_x4_sg U62015 ( .A(n25959), .B(n67456), .X(n25943) );
  nor_x1_sg U62016 ( .A(n25970), .B(n25971), .X(n25959) );
  nand_x4_sg U62017 ( .A(n25990), .B(n47332), .X(n25973) );
  nor_x1_sg U62018 ( .A(n26001), .B(n67475), .X(n25990) );
  nor_x1_sg U62019 ( .A(n22395), .B(n68477), .X(\shifter_0/n12757 ) );
  nor_x1_sg U62020 ( .A(n22395), .B(n68478), .X(\shifter_0/n12753 ) );
  nor_x1_sg U62021 ( .A(n22395), .B(n68479), .X(\shifter_0/n12745 ) );
  nor_x1_sg U62022 ( .A(n22395), .B(n68480), .X(\shifter_0/n12741 ) );
  nor_x1_sg U62023 ( .A(n22395), .B(n68481), .X(\shifter_0/n12733 ) );
  nor_x1_sg U62024 ( .A(n22395), .B(n68482), .X(\shifter_0/n12729 ) );
  nor_x1_sg U62025 ( .A(n22395), .B(n68483), .X(\shifter_0/n12721 ) );
  nor_x1_sg U62026 ( .A(n22395), .B(n68484), .X(\shifter_0/n12717 ) );
  nor_x1_sg U62027 ( .A(n22395), .B(n68485), .X(\shifter_0/n12701 ) );
  nor_x1_sg U62028 ( .A(n22395), .B(n68486), .X(\shifter_0/n12697 ) );
  nor_x1_sg U62029 ( .A(n68577), .B(n26003), .X(\shifter_0/n10277 ) );
  nor_x1_sg U62030 ( .A(n68578), .B(n26003), .X(\shifter_0/n10273 ) );
  nor_x1_sg U62031 ( .A(n68579), .B(n26003), .X(\shifter_0/n10265 ) );
  nor_x1_sg U62032 ( .A(n68580), .B(n26003), .X(\shifter_0/n10261 ) );
  nor_x1_sg U62033 ( .A(n68581), .B(n26003), .X(\shifter_0/n10253 ) );
  nor_x1_sg U62034 ( .A(n68582), .B(n26003), .X(\shifter_0/n10249 ) );
  nor_x1_sg U62035 ( .A(n68583), .B(n26003), .X(\shifter_0/n10241 ) );
  nor_x1_sg U62036 ( .A(n68584), .B(n26003), .X(\shifter_0/n10237 ) );
  nor_x1_sg U62037 ( .A(n68585), .B(n26003), .X(\shifter_0/n10221 ) );
  nor_x1_sg U62038 ( .A(n68586), .B(n26003), .X(\shifter_0/n10217 ) );
  nand_x1_sg U62039 ( .A(n68576), .B(n68572), .X(n23549) );
  nor_x1_sg U62040 ( .A(n67558), .B(n26135), .X(n26126) );
  nor_x1_sg U62041 ( .A(n67552), .B(n26096), .X(n26083) );
  nor_x1_sg U62042 ( .A(n67546), .B(n26227), .X(n26218) );
  nor_x1_sg U62043 ( .A(n67540), .B(n26193), .X(n26184) );
  nand_x2_sg U62044 ( .A(n67559), .B(n26153), .X(n26124) );
  nand_x2_sg U62045 ( .A(n26126), .B(n26127), .X(n26125) );
  nand_x2_sg U62046 ( .A(n67553), .B(n26116), .X(n26081) );
  nand_x2_sg U62047 ( .A(n26083), .B(n26084), .X(n26082) );
  nand_x2_sg U62048 ( .A(n67547), .B(n26245), .X(n26216) );
  nand_x2_sg U62049 ( .A(n26218), .B(n26219), .X(n26217) );
  nand_x2_sg U62050 ( .A(n67541), .B(n26211), .X(n26182) );
  nand_x2_sg U62051 ( .A(n26184), .B(n26185), .X(n26183) );
  nor_x1_sg U62052 ( .A(n22446), .B(n22451), .X(\shifter_0/n12508 ) );
  nor_x1_sg U62053 ( .A(n22446), .B(n22452), .X(\shifter_0/n12504 ) );
  nor_x1_sg U62054 ( .A(n22446), .B(n22453), .X(\shifter_0/n12500 ) );
  nor_x1_sg U62055 ( .A(n22446), .B(n22454), .X(\shifter_0/n12496 ) );
  nor_x1_sg U62056 ( .A(n22446), .B(n22455), .X(\shifter_0/n12492 ) );
  nor_x1_sg U62057 ( .A(n22446), .B(n22456), .X(\shifter_0/n12488 ) );
  nor_x1_sg U62058 ( .A(n22446), .B(n22457), .X(\shifter_0/n12484 ) );
  nor_x1_sg U62059 ( .A(n22446), .B(n22458), .X(\shifter_0/n12480 ) );
  nor_x1_sg U62060 ( .A(n22446), .B(n22459), .X(\shifter_0/n12476 ) );
  nor_x1_sg U62061 ( .A(n22446), .B(n22460), .X(\shifter_0/n12472 ) );
  nor_x1_sg U62062 ( .A(n22446), .B(n22461), .X(\shifter_0/n12468 ) );
  nor_x1_sg U62063 ( .A(n22446), .B(n22462), .X(\shifter_0/n12464 ) );
  nor_x1_sg U62064 ( .A(n22446), .B(n22463), .X(\shifter_0/n12460 ) );
  nor_x1_sg U62065 ( .A(n22446), .B(n22464), .X(\shifter_0/n12456 ) );
  nor_x1_sg U62066 ( .A(n22498), .B(n22503), .X(\shifter_0/n12348 ) );
  nor_x1_sg U62067 ( .A(n22498), .B(n22504), .X(\shifter_0/n12344 ) );
  nor_x1_sg U62068 ( .A(n22498), .B(n22505), .X(\shifter_0/n12340 ) );
  nor_x1_sg U62069 ( .A(n22498), .B(n22506), .X(\shifter_0/n12336 ) );
  nor_x1_sg U62070 ( .A(n22498), .B(n22507), .X(\shifter_0/n12332 ) );
  nor_x1_sg U62071 ( .A(n22498), .B(n22508), .X(\shifter_0/n12328 ) );
  nor_x1_sg U62072 ( .A(n22498), .B(n22509), .X(\shifter_0/n12324 ) );
  nor_x1_sg U62073 ( .A(n22498), .B(n22510), .X(\shifter_0/n12320 ) );
  nor_x1_sg U62074 ( .A(n22498), .B(n22511), .X(\shifter_0/n12316 ) );
  nor_x1_sg U62075 ( .A(n22498), .B(n22512), .X(\shifter_0/n12312 ) );
  nor_x1_sg U62076 ( .A(n22498), .B(n22513), .X(\shifter_0/n12308 ) );
  nor_x1_sg U62077 ( .A(n22498), .B(n22514), .X(\shifter_0/n12304 ) );
  nor_x1_sg U62078 ( .A(n22498), .B(n22515), .X(\shifter_0/n12300 ) );
  nor_x1_sg U62079 ( .A(n22498), .B(n22516), .X(\shifter_0/n12296 ) );
  nand_x4_sg U62080 ( .A(n26063), .B(n26064), .X(n26061) );
  nand_x1_sg U62081 ( .A(n67529), .B(n26067), .X(n26063) );
  nand_x1_sg U62082 ( .A(n26065), .B(n26066), .X(n26064) );
  nand_x1_sg U62083 ( .A(n33738), .B(n26066), .X(n26067) );
  nand_x4_sg U62084 ( .A(n26159), .B(n26160), .X(n26157) );
  nand_x1_sg U62085 ( .A(n67526), .B(n26163), .X(n26159) );
  nand_x1_sg U62086 ( .A(n26161), .B(n26162), .X(n26160) );
  nand_x1_sg U62087 ( .A(n26162), .B(n34219), .X(n26163) );
  nor_x1_sg U62088 ( .A(n22473), .B(n22478), .X(\shifter_0/n12428 ) );
  nor_x1_sg U62089 ( .A(n22473), .B(n22479), .X(\shifter_0/n12424 ) );
  nor_x1_sg U62090 ( .A(n22473), .B(n22480), .X(\shifter_0/n12420 ) );
  nor_x1_sg U62091 ( .A(n22473), .B(n22481), .X(\shifter_0/n12416 ) );
  nor_x1_sg U62092 ( .A(n22473), .B(n22482), .X(\shifter_0/n12412 ) );
  nor_x1_sg U62093 ( .A(n22473), .B(n22483), .X(\shifter_0/n12408 ) );
  nor_x1_sg U62094 ( .A(n22473), .B(n22484), .X(\shifter_0/n12404 ) );
  nor_x1_sg U62095 ( .A(n22473), .B(n22485), .X(\shifter_0/n12400 ) );
  nor_x1_sg U62096 ( .A(n22473), .B(n22486), .X(\shifter_0/n12396 ) );
  nor_x1_sg U62097 ( .A(n22473), .B(n22487), .X(\shifter_0/n12392 ) );
  nor_x1_sg U62098 ( .A(n22473), .B(n22488), .X(\shifter_0/n12388 ) );
  nor_x1_sg U62099 ( .A(n22473), .B(n22489), .X(\shifter_0/n12384 ) );
  nor_x1_sg U62100 ( .A(n22473), .B(n22490), .X(\shifter_0/n12380 ) );
  nor_x1_sg U62101 ( .A(n22473), .B(n22491), .X(\shifter_0/n12376 ) );
  nor_x1_sg U62102 ( .A(n22523), .B(n22528), .X(\shifter_0/n12268 ) );
  nor_x1_sg U62103 ( .A(n22523), .B(n22529), .X(\shifter_0/n12264 ) );
  nor_x1_sg U62104 ( .A(n22523), .B(n22530), .X(\shifter_0/n12260 ) );
  nor_x1_sg U62105 ( .A(n22523), .B(n22531), .X(\shifter_0/n12256 ) );
  nor_x1_sg U62106 ( .A(n22523), .B(n22532), .X(\shifter_0/n12252 ) );
  nor_x1_sg U62107 ( .A(n22523), .B(n22533), .X(\shifter_0/n12248 ) );
  nor_x1_sg U62108 ( .A(n22523), .B(n22534), .X(\shifter_0/n12244 ) );
  nor_x1_sg U62109 ( .A(n22523), .B(n22535), .X(\shifter_0/n12240 ) );
  nor_x1_sg U62110 ( .A(n22523), .B(n22536), .X(\shifter_0/n12236 ) );
  nor_x1_sg U62111 ( .A(n22523), .B(n22537), .X(\shifter_0/n12232 ) );
  nor_x1_sg U62112 ( .A(n22523), .B(n22538), .X(\shifter_0/n12228 ) );
  nor_x1_sg U62113 ( .A(n22523), .B(n22539), .X(\shifter_0/n12224 ) );
  nor_x1_sg U62114 ( .A(n22523), .B(n22540), .X(\shifter_0/n12220 ) );
  nor_x1_sg U62115 ( .A(n22523), .B(n22541), .X(\shifter_0/n12216 ) );
  nor_x1_sg U62116 ( .A(n22396), .B(n22401), .X(\shifter_0/n12668 ) );
  nor_x1_sg U62117 ( .A(n22396), .B(n22402), .X(\shifter_0/n12664 ) );
  nor_x1_sg U62118 ( .A(n22396), .B(n22403), .X(\shifter_0/n12660 ) );
  nor_x1_sg U62119 ( .A(n22396), .B(n22404), .X(\shifter_0/n12656 ) );
  nor_x1_sg U62120 ( .A(n22396), .B(n22405), .X(\shifter_0/n12652 ) );
  nor_x1_sg U62121 ( .A(n22396), .B(n22406), .X(\shifter_0/n12648 ) );
  nor_x1_sg U62122 ( .A(n22396), .B(n22407), .X(\shifter_0/n12644 ) );
  nor_x1_sg U62123 ( .A(n22396), .B(n22408), .X(\shifter_0/n12640 ) );
  nor_x1_sg U62124 ( .A(n22396), .B(n22409), .X(\shifter_0/n12636 ) );
  nor_x1_sg U62125 ( .A(n22396), .B(n22410), .X(\shifter_0/n12632 ) );
  nor_x1_sg U62126 ( .A(n22396), .B(n22411), .X(\shifter_0/n12628 ) );
  nor_x1_sg U62127 ( .A(n22396), .B(n22412), .X(\shifter_0/n12624 ) );
  nor_x1_sg U62128 ( .A(n22396), .B(n22413), .X(\shifter_0/n12620 ) );
  nor_x1_sg U62129 ( .A(n22396), .B(n22414), .X(\shifter_0/n12616 ) );
  nor_x1_sg U62130 ( .A(n22421), .B(n22426), .X(\shifter_0/n12588 ) );
  nor_x1_sg U62131 ( .A(n22421), .B(n22427), .X(\shifter_0/n12584 ) );
  nor_x1_sg U62132 ( .A(n22421), .B(n22428), .X(\shifter_0/n12580 ) );
  nor_x1_sg U62133 ( .A(n22421), .B(n22429), .X(\shifter_0/n12576 ) );
  nor_x1_sg U62134 ( .A(n22421), .B(n22430), .X(\shifter_0/n12572 ) );
  nor_x1_sg U62135 ( .A(n22421), .B(n22431), .X(\shifter_0/n12568 ) );
  nor_x1_sg U62136 ( .A(n22421), .B(n22432), .X(\shifter_0/n12564 ) );
  nor_x1_sg U62137 ( .A(n22421), .B(n22433), .X(\shifter_0/n12560 ) );
  nor_x1_sg U62138 ( .A(n22421), .B(n22434), .X(\shifter_0/n12556 ) );
  nor_x1_sg U62139 ( .A(n22421), .B(n22435), .X(\shifter_0/n12552 ) );
  nor_x1_sg U62140 ( .A(n22421), .B(n22436), .X(\shifter_0/n12548 ) );
  nor_x1_sg U62141 ( .A(n22421), .B(n22437), .X(\shifter_0/n12544 ) );
  nor_x1_sg U62142 ( .A(n22421), .B(n22438), .X(\shifter_0/n12540 ) );
  nor_x1_sg U62143 ( .A(n22421), .B(n22439), .X(\shifter_0/n12536 ) );
  nor_x1_sg U62144 ( .A(n22446), .B(n22447), .X(\shifter_0/n12524 ) );
  nor_x1_sg U62145 ( .A(n22446), .B(n22448), .X(\shifter_0/n12520 ) );
  nor_x1_sg U62146 ( .A(n22446), .B(n22449), .X(\shifter_0/n12516 ) );
  nor_x1_sg U62147 ( .A(n22446), .B(n22450), .X(\shifter_0/n12512 ) );
  nor_x1_sg U62148 ( .A(n22498), .B(n22499), .X(\shifter_0/n12364 ) );
  nor_x1_sg U62149 ( .A(n22498), .B(n22500), .X(\shifter_0/n12360 ) );
  nor_x1_sg U62150 ( .A(n22498), .B(n22501), .X(\shifter_0/n12356 ) );
  nor_x1_sg U62151 ( .A(n22498), .B(n22502), .X(\shifter_0/n12352 ) );
  nor_x1_sg U62152 ( .A(n57510), .B(n22551), .X(\shifter_0/n12188 ) );
  nor_x1_sg U62153 ( .A(n57510), .B(n22552), .X(\shifter_0/n12184 ) );
  nor_x1_sg U62154 ( .A(n57510), .B(n22553), .X(\shifter_0/n12180 ) );
  nor_x1_sg U62155 ( .A(n57510), .B(n22554), .X(\shifter_0/n12176 ) );
  nor_x1_sg U62156 ( .A(n57510), .B(n22555), .X(\shifter_0/n12172 ) );
  nor_x1_sg U62157 ( .A(n57510), .B(n22556), .X(\shifter_0/n12168 ) );
  nor_x1_sg U62158 ( .A(n57510), .B(n22557), .X(\shifter_0/n12164 ) );
  nor_x1_sg U62159 ( .A(n57510), .B(n22558), .X(\shifter_0/n12160 ) );
  nor_x1_sg U62160 ( .A(n57510), .B(n22559), .X(\shifter_0/n12156 ) );
  nor_x1_sg U62161 ( .A(n57507), .B(n22602), .X(\shifter_0/n12028 ) );
  nor_x1_sg U62162 ( .A(n57507), .B(n22603), .X(\shifter_0/n12024 ) );
  nor_x1_sg U62163 ( .A(n57507), .B(n22604), .X(\shifter_0/n12020 ) );
  nor_x1_sg U62164 ( .A(n57507), .B(n22605), .X(\shifter_0/n12016 ) );
  nor_x1_sg U62165 ( .A(n57507), .B(n22606), .X(\shifter_0/n12012 ) );
  nor_x1_sg U62166 ( .A(n57507), .B(n22607), .X(\shifter_0/n12008 ) );
  nor_x1_sg U62167 ( .A(n57507), .B(n22608), .X(\shifter_0/n12004 ) );
  nor_x1_sg U62168 ( .A(n57507), .B(n22609), .X(\shifter_0/n12000 ) );
  nor_x1_sg U62169 ( .A(n57507), .B(n22610), .X(\shifter_0/n11996 ) );
  nor_x1_sg U62170 ( .A(n57516), .B(n22577), .X(\shifter_0/n12108 ) );
  nor_x1_sg U62171 ( .A(n57516), .B(n22578), .X(\shifter_0/n12104 ) );
  nor_x1_sg U62172 ( .A(n57516), .B(n22579), .X(\shifter_0/n12100 ) );
  nor_x1_sg U62173 ( .A(n57516), .B(n22580), .X(\shifter_0/n12096 ) );
  nor_x1_sg U62174 ( .A(n57516), .B(n22581), .X(\shifter_0/n12092 ) );
  nor_x1_sg U62175 ( .A(n57516), .B(n22582), .X(\shifter_0/n12088 ) );
  nor_x1_sg U62176 ( .A(n57516), .B(n22583), .X(\shifter_0/n12084 ) );
  nor_x1_sg U62177 ( .A(n57516), .B(n22584), .X(\shifter_0/n12080 ) );
  nor_x1_sg U62178 ( .A(n57516), .B(n22585), .X(\shifter_0/n12076 ) );
  nor_x1_sg U62179 ( .A(n57513), .B(n22629), .X(\shifter_0/n11948 ) );
  nor_x1_sg U62180 ( .A(n57513), .B(n22630), .X(\shifter_0/n11944 ) );
  nor_x1_sg U62181 ( .A(n57513), .B(n22631), .X(\shifter_0/n11940 ) );
  nor_x1_sg U62182 ( .A(n57513), .B(n22632), .X(\shifter_0/n11936 ) );
  nor_x1_sg U62183 ( .A(n57513), .B(n22633), .X(\shifter_0/n11932 ) );
  nor_x1_sg U62184 ( .A(n57513), .B(n22634), .X(\shifter_0/n11928 ) );
  nor_x1_sg U62185 ( .A(n57513), .B(n22635), .X(\shifter_0/n11924 ) );
  nor_x1_sg U62186 ( .A(n57513), .B(n22636), .X(\shifter_0/n11920 ) );
  nor_x1_sg U62187 ( .A(n57513), .B(n22637), .X(\shifter_0/n11916 ) );
  nor_x1_sg U62188 ( .A(n57510), .B(n22560), .X(\shifter_0/n12152 ) );
  nor_x1_sg U62189 ( .A(n57510), .B(n22561), .X(\shifter_0/n12148 ) );
  nor_x1_sg U62190 ( .A(n57510), .B(n22562), .X(\shifter_0/n12144 ) );
  nor_x1_sg U62191 ( .A(n57510), .B(n22563), .X(\shifter_0/n12140 ) );
  nor_x1_sg U62192 ( .A(n57510), .B(n22564), .X(\shifter_0/n12136 ) );
  nor_x1_sg U62193 ( .A(n57507), .B(n22611), .X(\shifter_0/n11992 ) );
  nor_x1_sg U62194 ( .A(n57507), .B(n22612), .X(\shifter_0/n11988 ) );
  nor_x1_sg U62195 ( .A(n57507), .B(n22613), .X(\shifter_0/n11984 ) );
  nor_x1_sg U62196 ( .A(n57507), .B(n22614), .X(\shifter_0/n11980 ) );
  nor_x1_sg U62197 ( .A(n57507), .B(n22615), .X(\shifter_0/n11976 ) );
  nor_x1_sg U62198 ( .A(n57516), .B(n22586), .X(\shifter_0/n12072 ) );
  nor_x1_sg U62199 ( .A(n57516), .B(n22587), .X(\shifter_0/n12068 ) );
  nor_x1_sg U62200 ( .A(n57516), .B(n22588), .X(\shifter_0/n12064 ) );
  nor_x1_sg U62201 ( .A(n57516), .B(n22589), .X(\shifter_0/n12060 ) );
  nor_x1_sg U62202 ( .A(n57516), .B(n22590), .X(\shifter_0/n12056 ) );
  nor_x1_sg U62203 ( .A(n57513), .B(n22638), .X(\shifter_0/n11912 ) );
  nor_x1_sg U62204 ( .A(n57513), .B(n22639), .X(\shifter_0/n11908 ) );
  nor_x1_sg U62205 ( .A(n57513), .B(n22640), .X(\shifter_0/n11904 ) );
  nor_x1_sg U62206 ( .A(n57513), .B(n22641), .X(\shifter_0/n11900 ) );
  nor_x1_sg U62207 ( .A(n57513), .B(n22642), .X(\shifter_0/n11896 ) );
  nor_x1_sg U62208 ( .A(n22473), .B(n22474), .X(\shifter_0/n12444 ) );
  nor_x1_sg U62209 ( .A(n22473), .B(n22475), .X(\shifter_0/n12440 ) );
  nor_x1_sg U62210 ( .A(n22473), .B(n22476), .X(\shifter_0/n12436 ) );
  nor_x1_sg U62211 ( .A(n22473), .B(n22477), .X(\shifter_0/n12432 ) );
  nor_x1_sg U62212 ( .A(n22523), .B(n22524), .X(\shifter_0/n12284 ) );
  nor_x1_sg U62213 ( .A(n22523), .B(n22525), .X(\shifter_0/n12280 ) );
  nor_x1_sg U62214 ( .A(n22523), .B(n22526), .X(\shifter_0/n12276 ) );
  nor_x1_sg U62215 ( .A(n22523), .B(n22527), .X(\shifter_0/n12272 ) );
  nor_x1_sg U62216 ( .A(n22396), .B(n22397), .X(\shifter_0/n12684 ) );
  nor_x1_sg U62217 ( .A(n22396), .B(n22398), .X(\shifter_0/n12680 ) );
  nor_x1_sg U62218 ( .A(n22396), .B(n22399), .X(\shifter_0/n12676 ) );
  nor_x1_sg U62219 ( .A(n22396), .B(n22400), .X(\shifter_0/n12672 ) );
  nor_x1_sg U62220 ( .A(n22421), .B(n22422), .X(\shifter_0/n12604 ) );
  nor_x1_sg U62221 ( .A(n22421), .B(n22423), .X(\shifter_0/n12600 ) );
  nor_x1_sg U62222 ( .A(n22421), .B(n22424), .X(\shifter_0/n12596 ) );
  nor_x1_sg U62223 ( .A(n22421), .B(n22425), .X(\shifter_0/n12592 ) );
  nor_x1_sg U62224 ( .A(n57145), .B(n23418), .X(\shifter_0/n11405 ) );
  nor_x1_sg U62225 ( .A(n57145), .B(n23427), .X(\shifter_0/n11401 ) );
  nor_x1_sg U62226 ( .A(n57145), .B(n23433), .X(\shifter_0/n11397 ) );
  nor_x1_sg U62227 ( .A(n57145), .B(n23439), .X(\shifter_0/n11393 ) );
  nor_x1_sg U62228 ( .A(n57145), .B(n23445), .X(\shifter_0/n11389 ) );
  nor_x1_sg U62229 ( .A(n57145), .B(n23451), .X(\shifter_0/n11385 ) );
  nor_x1_sg U62230 ( .A(n57145), .B(n23457), .X(\shifter_0/n11381 ) );
  nor_x1_sg U62231 ( .A(n57145), .B(n23463), .X(\shifter_0/n11377 ) );
  nor_x1_sg U62232 ( .A(n57145), .B(n23469), .X(\shifter_0/n11373 ) );
  nor_x1_sg U62233 ( .A(n57145), .B(n23475), .X(\shifter_0/n11369 ) );
  nor_x1_sg U62234 ( .A(n57145), .B(n23481), .X(\shifter_0/n11365 ) );
  nor_x1_sg U62235 ( .A(n57145), .B(n23487), .X(\shifter_0/n11361 ) );
  nor_x1_sg U62236 ( .A(n57145), .B(n23493), .X(\shifter_0/n11357 ) );
  nor_x1_sg U62237 ( .A(n57145), .B(n23499), .X(\shifter_0/n11353 ) );
  nor_x1_sg U62238 ( .A(n57145), .B(n23505), .X(\shifter_0/n11349 ) );
  nor_x1_sg U62239 ( .A(n57145), .B(n23511), .X(\shifter_0/n11345 ) );
  nor_x1_sg U62240 ( .A(n57145), .B(n23517), .X(\shifter_0/n11341 ) );
  nor_x1_sg U62241 ( .A(n57145), .B(n23523), .X(\shifter_0/n11337 ) );
  nor_x1_sg U62242 ( .A(n57145), .B(n23529), .X(\shifter_0/n11333 ) );
  nor_x1_sg U62243 ( .A(n57145), .B(n23535), .X(\shifter_0/n11329 ) );
  nor_x1_sg U62244 ( .A(n57142), .B(n23552), .X(\shifter_0/n11325 ) );
  nor_x1_sg U62245 ( .A(n57142), .B(n23559), .X(\shifter_0/n11321 ) );
  nor_x1_sg U62246 ( .A(n57142), .B(n23565), .X(\shifter_0/n11317 ) );
  nor_x1_sg U62247 ( .A(n57142), .B(n23571), .X(\shifter_0/n11313 ) );
  nor_x1_sg U62248 ( .A(n57142), .B(n23577), .X(\shifter_0/n11309 ) );
  nor_x1_sg U62249 ( .A(n57142), .B(n23583), .X(\shifter_0/n11305 ) );
  nor_x1_sg U62250 ( .A(n57142), .B(n23589), .X(\shifter_0/n11301 ) );
  nor_x1_sg U62251 ( .A(n57142), .B(n23595), .X(\shifter_0/n11297 ) );
  nor_x1_sg U62252 ( .A(n57142), .B(n23601), .X(\shifter_0/n11293 ) );
  nor_x1_sg U62253 ( .A(n57142), .B(n23607), .X(\shifter_0/n11289 ) );
  nor_x1_sg U62254 ( .A(n57142), .B(n23613), .X(\shifter_0/n11285 ) );
  nor_x1_sg U62255 ( .A(n57142), .B(n23619), .X(\shifter_0/n11281 ) );
  nor_x1_sg U62256 ( .A(n57142), .B(n23625), .X(\shifter_0/n11277 ) );
  nor_x1_sg U62257 ( .A(n57142), .B(n23631), .X(\shifter_0/n11273 ) );
  nor_x1_sg U62258 ( .A(n57142), .B(n23637), .X(\shifter_0/n11269 ) );
  nor_x1_sg U62259 ( .A(n57142), .B(n23643), .X(\shifter_0/n11265 ) );
  nor_x1_sg U62260 ( .A(n57142), .B(n23649), .X(\shifter_0/n11261 ) );
  nor_x1_sg U62261 ( .A(n57142), .B(n23655), .X(\shifter_0/n11257 ) );
  nor_x1_sg U62262 ( .A(n57142), .B(n23661), .X(\shifter_0/n11253 ) );
  nor_x1_sg U62263 ( .A(n57142), .B(n23667), .X(\shifter_0/n11249 ) );
  nor_x1_sg U62264 ( .A(n57139), .B(n23683), .X(\shifter_0/n11245 ) );
  nor_x1_sg U62265 ( .A(n57139), .B(n23691), .X(\shifter_0/n11241 ) );
  nor_x1_sg U62266 ( .A(n57139), .B(n23697), .X(\shifter_0/n11237 ) );
  nor_x1_sg U62267 ( .A(n57139), .B(n23703), .X(\shifter_0/n11233 ) );
  nor_x1_sg U62268 ( .A(n57139), .B(n23709), .X(\shifter_0/n11229 ) );
  nor_x1_sg U62269 ( .A(n57139), .B(n23715), .X(\shifter_0/n11225 ) );
  nor_x1_sg U62270 ( .A(n57139), .B(n23721), .X(\shifter_0/n11221 ) );
  nor_x1_sg U62271 ( .A(n57139), .B(n23727), .X(\shifter_0/n11217 ) );
  nor_x1_sg U62272 ( .A(n57139), .B(n23733), .X(\shifter_0/n11213 ) );
  nor_x1_sg U62273 ( .A(n57139), .B(n23739), .X(\shifter_0/n11209 ) );
  nor_x1_sg U62274 ( .A(n57139), .B(n23745), .X(\shifter_0/n11205 ) );
  nor_x1_sg U62275 ( .A(n57139), .B(n23751), .X(\shifter_0/n11201 ) );
  nor_x1_sg U62276 ( .A(n57139), .B(n23757), .X(\shifter_0/n11197 ) );
  nor_x1_sg U62277 ( .A(n57139), .B(n23763), .X(\shifter_0/n11193 ) );
  nor_x1_sg U62278 ( .A(n57139), .B(n23769), .X(\shifter_0/n11189 ) );
  nor_x1_sg U62279 ( .A(n57139), .B(n23775), .X(\shifter_0/n11185 ) );
  nor_x1_sg U62280 ( .A(n57139), .B(n23781), .X(\shifter_0/n11181 ) );
  nor_x1_sg U62281 ( .A(n57139), .B(n23787), .X(\shifter_0/n11177 ) );
  nor_x1_sg U62282 ( .A(n57139), .B(n23793), .X(\shifter_0/n11173 ) );
  nor_x1_sg U62283 ( .A(n57139), .B(n23799), .X(\shifter_0/n11169 ) );
  nor_x1_sg U62284 ( .A(n57136), .B(n23813), .X(\shifter_0/n11165 ) );
  nor_x1_sg U62285 ( .A(n57136), .B(n23820), .X(\shifter_0/n11161 ) );
  nor_x1_sg U62286 ( .A(n57136), .B(n23826), .X(\shifter_0/n11157 ) );
  nor_x1_sg U62287 ( .A(n57136), .B(n23832), .X(\shifter_0/n11153 ) );
  nor_x1_sg U62288 ( .A(n57136), .B(n23838), .X(\shifter_0/n11149 ) );
  nor_x1_sg U62289 ( .A(n57136), .B(n23844), .X(\shifter_0/n11145 ) );
  nor_x1_sg U62290 ( .A(n57136), .B(n23850), .X(\shifter_0/n11141 ) );
  nor_x1_sg U62291 ( .A(n57136), .B(n23856), .X(\shifter_0/n11137 ) );
  nor_x1_sg U62292 ( .A(n57136), .B(n23862), .X(\shifter_0/n11133 ) );
  nor_x1_sg U62293 ( .A(n57136), .B(n23868), .X(\shifter_0/n11129 ) );
  nor_x1_sg U62294 ( .A(n57136), .B(n23874), .X(\shifter_0/n11125 ) );
  nor_x1_sg U62295 ( .A(n57136), .B(n23880), .X(\shifter_0/n11121 ) );
  nor_x1_sg U62296 ( .A(n57136), .B(n23886), .X(\shifter_0/n11117 ) );
  nor_x1_sg U62297 ( .A(n57136), .B(n23892), .X(\shifter_0/n11113 ) );
  nor_x1_sg U62298 ( .A(n57136), .B(n23898), .X(\shifter_0/n11109 ) );
  nor_x1_sg U62299 ( .A(n57136), .B(n23904), .X(\shifter_0/n11105 ) );
  nor_x1_sg U62300 ( .A(n57136), .B(n23910), .X(\shifter_0/n11101 ) );
  nor_x1_sg U62301 ( .A(n57136), .B(n23916), .X(\shifter_0/n11097 ) );
  nor_x1_sg U62302 ( .A(n57136), .B(n23922), .X(\shifter_0/n11093 ) );
  nor_x1_sg U62303 ( .A(n57136), .B(n23928), .X(\shifter_0/n11089 ) );
  nor_x1_sg U62304 ( .A(n57133), .B(n24160), .X(\shifter_0/n10925 ) );
  nor_x1_sg U62305 ( .A(n57133), .B(n24166), .X(\shifter_0/n10921 ) );
  nor_x1_sg U62306 ( .A(n57133), .B(n24171), .X(\shifter_0/n10917 ) );
  nor_x1_sg U62307 ( .A(n57133), .B(n24176), .X(\shifter_0/n10913 ) );
  nor_x1_sg U62308 ( .A(n57133), .B(n24181), .X(\shifter_0/n10909 ) );
  nor_x1_sg U62309 ( .A(n57133), .B(n24186), .X(\shifter_0/n10905 ) );
  nor_x1_sg U62310 ( .A(n57133), .B(n24191), .X(\shifter_0/n10901 ) );
  nor_x1_sg U62311 ( .A(n57133), .B(n24196), .X(\shifter_0/n10897 ) );
  nor_x1_sg U62312 ( .A(n57133), .B(n24201), .X(\shifter_0/n10893 ) );
  nor_x1_sg U62313 ( .A(n57133), .B(n24206), .X(\shifter_0/n10889 ) );
  nor_x1_sg U62314 ( .A(n57133), .B(n24211), .X(\shifter_0/n10885 ) );
  nor_x1_sg U62315 ( .A(n57133), .B(n24216), .X(\shifter_0/n10881 ) );
  nor_x1_sg U62316 ( .A(n57133), .B(n24221), .X(\shifter_0/n10877 ) );
  nor_x1_sg U62317 ( .A(n57133), .B(n24226), .X(\shifter_0/n10873 ) );
  nor_x1_sg U62318 ( .A(n57133), .B(n24231), .X(\shifter_0/n10869 ) );
  nor_x1_sg U62319 ( .A(n57133), .B(n24236), .X(\shifter_0/n10865 ) );
  nor_x1_sg U62320 ( .A(n57133), .B(n24241), .X(\shifter_0/n10861 ) );
  nor_x1_sg U62321 ( .A(n57133), .B(n24246), .X(\shifter_0/n10857 ) );
  nor_x1_sg U62322 ( .A(n57133), .B(n24251), .X(\shifter_0/n10853 ) );
  nor_x1_sg U62323 ( .A(n57133), .B(n24256), .X(\shifter_0/n10849 ) );
  nor_x1_sg U62324 ( .A(n57131), .B(n24269), .X(\shifter_0/n10845 ) );
  nor_x1_sg U62325 ( .A(n57131), .B(n24275), .X(\shifter_0/n10841 ) );
  nor_x1_sg U62326 ( .A(n57131), .B(n24280), .X(\shifter_0/n10837 ) );
  nor_x1_sg U62327 ( .A(n57131), .B(n24285), .X(\shifter_0/n10833 ) );
  nor_x1_sg U62328 ( .A(n57131), .B(n24290), .X(\shifter_0/n10829 ) );
  nor_x1_sg U62329 ( .A(n57131), .B(n24295), .X(\shifter_0/n10825 ) );
  nor_x1_sg U62330 ( .A(n57131), .B(n24300), .X(\shifter_0/n10821 ) );
  nor_x1_sg U62331 ( .A(n57131), .B(n24305), .X(\shifter_0/n10817 ) );
  nor_x1_sg U62332 ( .A(n57131), .B(n24310), .X(\shifter_0/n10813 ) );
  nor_x1_sg U62333 ( .A(n57131), .B(n24315), .X(\shifter_0/n10809 ) );
  nor_x1_sg U62334 ( .A(n57131), .B(n24320), .X(\shifter_0/n10805 ) );
  nor_x1_sg U62335 ( .A(n57131), .B(n24325), .X(\shifter_0/n10801 ) );
  nor_x1_sg U62336 ( .A(n57131), .B(n24330), .X(\shifter_0/n10797 ) );
  nor_x1_sg U62337 ( .A(n57131), .B(n24335), .X(\shifter_0/n10793 ) );
  nor_x1_sg U62338 ( .A(n57131), .B(n24340), .X(\shifter_0/n10789 ) );
  nor_x1_sg U62339 ( .A(n57131), .B(n24345), .X(\shifter_0/n10785 ) );
  nor_x1_sg U62340 ( .A(n57131), .B(n24350), .X(\shifter_0/n10781 ) );
  nor_x1_sg U62341 ( .A(n57131), .B(n24355), .X(\shifter_0/n10777 ) );
  nor_x1_sg U62342 ( .A(n57131), .B(n24360), .X(\shifter_0/n10773 ) );
  nor_x1_sg U62343 ( .A(n57131), .B(n24365), .X(\shifter_0/n10769 ) );
  nor_x1_sg U62344 ( .A(n57122), .B(n24602), .X(\shifter_0/n10605 ) );
  nor_x1_sg U62345 ( .A(n57122), .B(n24608), .X(\shifter_0/n10601 ) );
  nor_x1_sg U62346 ( .A(n57122), .B(n24612), .X(\shifter_0/n10597 ) );
  nor_x1_sg U62347 ( .A(n57122), .B(n24616), .X(\shifter_0/n10593 ) );
  nor_x1_sg U62348 ( .A(n57122), .B(n24620), .X(\shifter_0/n10589 ) );
  nor_x1_sg U62349 ( .A(n57122), .B(n24624), .X(\shifter_0/n10585 ) );
  nor_x1_sg U62350 ( .A(n57122), .B(n24628), .X(\shifter_0/n10581 ) );
  nor_x1_sg U62351 ( .A(n57122), .B(n24632), .X(\shifter_0/n10577 ) );
  nor_x1_sg U62352 ( .A(n57122), .B(n24636), .X(\shifter_0/n10573 ) );
  nor_x1_sg U62353 ( .A(n57122), .B(n24640), .X(\shifter_0/n10569 ) );
  nor_x1_sg U62354 ( .A(n57122), .B(n24644), .X(\shifter_0/n10565 ) );
  nor_x1_sg U62355 ( .A(n57122), .B(n24648), .X(\shifter_0/n10561 ) );
  nor_x1_sg U62356 ( .A(n57122), .B(n24652), .X(\shifter_0/n10557 ) );
  nor_x1_sg U62357 ( .A(n57122), .B(n24656), .X(\shifter_0/n10553 ) );
  nor_x1_sg U62358 ( .A(n57122), .B(n24660), .X(\shifter_0/n10549 ) );
  nor_x1_sg U62359 ( .A(n57122), .B(n24664), .X(\shifter_0/n10545 ) );
  nor_x1_sg U62360 ( .A(n57122), .B(n24668), .X(\shifter_0/n10541 ) );
  nor_x1_sg U62361 ( .A(n57122), .B(n24672), .X(\shifter_0/n10537 ) );
  nor_x1_sg U62362 ( .A(n57122), .B(n24676), .X(\shifter_0/n10533 ) );
  nor_x1_sg U62363 ( .A(n57122), .B(n24680), .X(\shifter_0/n10529 ) );
  nor_x1_sg U62364 ( .A(n57119), .B(n24697), .X(\shifter_0/n10525 ) );
  nor_x1_sg U62365 ( .A(n57119), .B(n24702), .X(\shifter_0/n10521 ) );
  nor_x1_sg U62366 ( .A(n57119), .B(n24706), .X(\shifter_0/n10517 ) );
  nor_x1_sg U62367 ( .A(n57119), .B(n24710), .X(\shifter_0/n10513 ) );
  nor_x1_sg U62368 ( .A(n57119), .B(n24714), .X(\shifter_0/n10509 ) );
  nor_x1_sg U62369 ( .A(n57119), .B(n24718), .X(\shifter_0/n10505 ) );
  nor_x1_sg U62370 ( .A(n57119), .B(n24722), .X(\shifter_0/n10501 ) );
  nor_x1_sg U62371 ( .A(n57119), .B(n24726), .X(\shifter_0/n10497 ) );
  nor_x1_sg U62372 ( .A(n57119), .B(n24730), .X(\shifter_0/n10493 ) );
  nor_x1_sg U62373 ( .A(n57119), .B(n24734), .X(\shifter_0/n10489 ) );
  nor_x1_sg U62374 ( .A(n57119), .B(n24738), .X(\shifter_0/n10485 ) );
  nor_x1_sg U62375 ( .A(n57119), .B(n24742), .X(\shifter_0/n10481 ) );
  nor_x1_sg U62376 ( .A(n57119), .B(n24746), .X(\shifter_0/n10477 ) );
  nor_x1_sg U62377 ( .A(n57119), .B(n24750), .X(\shifter_0/n10473 ) );
  nor_x1_sg U62378 ( .A(n57119), .B(n24754), .X(\shifter_0/n10469 ) );
  nor_x1_sg U62379 ( .A(n57119), .B(n24758), .X(\shifter_0/n10465 ) );
  nor_x1_sg U62380 ( .A(n57119), .B(n24762), .X(\shifter_0/n10461 ) );
  nor_x1_sg U62381 ( .A(n57119), .B(n24766), .X(\shifter_0/n10457 ) );
  nor_x1_sg U62382 ( .A(n57119), .B(n24770), .X(\shifter_0/n10453 ) );
  nor_x1_sg U62383 ( .A(n57119), .B(n24774), .X(\shifter_0/n10449 ) );
  nor_x1_sg U62384 ( .A(n57510), .B(n22547), .X(\shifter_0/n12204 ) );
  nor_x1_sg U62385 ( .A(n57510), .B(n22548), .X(\shifter_0/n12200 ) );
  nor_x1_sg U62386 ( .A(n57510), .B(n22549), .X(\shifter_0/n12196 ) );
  nor_x1_sg U62387 ( .A(n57510), .B(n22550), .X(\shifter_0/n12192 ) );
  nor_x1_sg U62388 ( .A(n57507), .B(n22598), .X(\shifter_0/n12044 ) );
  nor_x1_sg U62389 ( .A(n57507), .B(n22599), .X(\shifter_0/n12040 ) );
  nor_x1_sg U62390 ( .A(n57507), .B(n22600), .X(\shifter_0/n12036 ) );
  nor_x1_sg U62391 ( .A(n57507), .B(n22601), .X(\shifter_0/n12032 ) );
  nor_x1_sg U62392 ( .A(n57516), .B(n22573), .X(\shifter_0/n12124 ) );
  nor_x1_sg U62393 ( .A(n57516), .B(n22574), .X(\shifter_0/n12120 ) );
  nor_x1_sg U62394 ( .A(n57516), .B(n22575), .X(\shifter_0/n12116 ) );
  nor_x1_sg U62395 ( .A(n57516), .B(n22576), .X(\shifter_0/n12112 ) );
  nor_x1_sg U62396 ( .A(n57513), .B(n22625), .X(\shifter_0/n11964 ) );
  nor_x1_sg U62397 ( .A(n57513), .B(n22626), .X(\shifter_0/n11960 ) );
  nor_x1_sg U62398 ( .A(n57513), .B(n22627), .X(\shifter_0/n11956 ) );
  nor_x1_sg U62399 ( .A(n57513), .B(n22628), .X(\shifter_0/n11952 ) );
  nor_x1_sg U62400 ( .A(n57113), .B(n26073), .X(\filter_0/n8255 ) );
  nor_x1_sg U62401 ( .A(n57113), .B(n26165), .X(\filter_0/n8247 ) );
  nor_x1_sg U62402 ( .A(n57113), .B(n26173), .X(\filter_0/n8240 ) );
  nand_x2_sg U62403 ( .A(n24843), .B(n24844), .X(n24842) );
  nand_x2_sg U62404 ( .A(n24933), .B(n24934), .X(n24932) );
  nand_x2_sg U62405 ( .A(n25023), .B(n25024), .X(n25022) );
  nand_x2_sg U62406 ( .A(n25113), .B(n25114), .X(n25112) );
  nand_x2_sg U62407 ( .A(n25203), .B(n25204), .X(n25202) );
  nand_x2_sg U62408 ( .A(n25233), .B(n25234), .X(n25232) );
  nand_x2_sg U62409 ( .A(n25263), .B(n25264), .X(n25262) );
  nand_x2_sg U62410 ( .A(n25353), .B(n25354), .X(n25352) );
  nand_x2_sg U62411 ( .A(n25384), .B(n25385), .X(n25383) );
  nand_x2_sg U62412 ( .A(n25445), .B(n25446), .X(n25444) );
  nand_x2_sg U62413 ( .A(n25535), .B(n25536), .X(n25534) );
  nand_x2_sg U62414 ( .A(n25625), .B(n25626), .X(n25624) );
  nand_x2_sg U62415 ( .A(n25715), .B(n25716), .X(n25714) );
  nand_x2_sg U62416 ( .A(n25805), .B(n25806), .X(n25804) );
  nand_x2_sg U62417 ( .A(n25835), .B(n25836), .X(n25834) );
  nand_x2_sg U62418 ( .A(n25865), .B(n25866), .X(n25864) );
  nand_x2_sg U62419 ( .A(n25955), .B(n25956), .X(n25954) );
  nand_x2_sg U62420 ( .A(n25986), .B(n25987), .X(n25985) );
  nand_x2_sg U62421 ( .A(n24807), .B(n24808), .X(n24806) );
  nand_x2_sg U62422 ( .A(n24873), .B(n24874), .X(n24872) );
  nand_x2_sg U62423 ( .A(n24903), .B(n24904), .X(n24902) );
  nand_x2_sg U62424 ( .A(n24963), .B(n24964), .X(n24962) );
  nand_x2_sg U62425 ( .A(n24993), .B(n24994), .X(n24992) );
  nand_x2_sg U62426 ( .A(n25053), .B(n25054), .X(n25052) );
  nand_x2_sg U62427 ( .A(n25083), .B(n25084), .X(n25082) );
  nand_x2_sg U62428 ( .A(n25143), .B(n25144), .X(n25142) );
  nand_x2_sg U62429 ( .A(n25173), .B(n25174), .X(n25172) );
  nand_x2_sg U62430 ( .A(n25293), .B(n25294), .X(n25292) );
  nand_x2_sg U62431 ( .A(n25323), .B(n25324), .X(n25322) );
  nand_x2_sg U62432 ( .A(n25415), .B(n25416), .X(n25414) );
  nand_x2_sg U62433 ( .A(n25475), .B(n25476), .X(n25474) );
  nand_x2_sg U62434 ( .A(n25505), .B(n25506), .X(n25504) );
  nand_x2_sg U62435 ( .A(n25565), .B(n25566), .X(n25564) );
  nand_x2_sg U62436 ( .A(n25595), .B(n25596), .X(n25594) );
  nand_x2_sg U62437 ( .A(n25655), .B(n25656), .X(n25654) );
  nand_x2_sg U62438 ( .A(n25685), .B(n25686), .X(n25684) );
  nand_x2_sg U62439 ( .A(n25745), .B(n25746), .X(n25744) );
  nand_x2_sg U62440 ( .A(n25775), .B(n25776), .X(n25774) );
  nand_x2_sg U62441 ( .A(n25895), .B(n25896), .X(n25894) );
  nand_x2_sg U62442 ( .A(n25925), .B(n25926), .X(n25924) );
  nand_x4_sg U62443 ( .A(n24164), .B(n24382), .X(n24379) );
  nand_x4_sg U62444 ( .A(n24169), .B(n24387), .X(n24385) );
  nand_x4_sg U62445 ( .A(n24174), .B(n24392), .X(n24390) );
  nand_x4_sg U62446 ( .A(n24179), .B(n24397), .X(n24395) );
  nand_x4_sg U62447 ( .A(n24184), .B(n24402), .X(n24400) );
  nand_x4_sg U62448 ( .A(n24189), .B(n24407), .X(n24405) );
  nand_x4_sg U62449 ( .A(n24194), .B(n24412), .X(n24410) );
  nand_x4_sg U62450 ( .A(n24199), .B(n24417), .X(n24415) );
  nand_x4_sg U62451 ( .A(n24204), .B(n24422), .X(n24420) );
  nand_x4_sg U62452 ( .A(n24209), .B(n24427), .X(n24425) );
  nand_x4_sg U62453 ( .A(n24214), .B(n24432), .X(n24430) );
  nand_x4_sg U62454 ( .A(n24219), .B(n24437), .X(n24435) );
  nand_x4_sg U62455 ( .A(n24224), .B(n24442), .X(n24440) );
  nand_x4_sg U62456 ( .A(n24229), .B(n24447), .X(n24445) );
  nand_x4_sg U62457 ( .A(n24234), .B(n24452), .X(n24450) );
  nand_x4_sg U62458 ( .A(n24239), .B(n24457), .X(n24455) );
  nand_x4_sg U62459 ( .A(n24244), .B(n24462), .X(n24460) );
  nand_x4_sg U62460 ( .A(n24249), .B(n24467), .X(n24465) );
  nand_x4_sg U62461 ( .A(n24254), .B(n24472), .X(n24470) );
  nand_x4_sg U62462 ( .A(n24267), .B(n24488), .X(n24475) );
  nand_x4_sg U62463 ( .A(n24273), .B(n24494), .X(n24491) );
  nand_x4_sg U62464 ( .A(n24278), .B(n24499), .X(n24497) );
  nand_x4_sg U62465 ( .A(n24283), .B(n24504), .X(n24502) );
  nand_x4_sg U62466 ( .A(n24288), .B(n24509), .X(n24507) );
  nand_x4_sg U62467 ( .A(n24293), .B(n24514), .X(n24512) );
  nand_x4_sg U62468 ( .A(n24298), .B(n24519), .X(n24517) );
  nand_x4_sg U62469 ( .A(n24303), .B(n24524), .X(n24522) );
  nand_x4_sg U62470 ( .A(n24308), .B(n24529), .X(n24527) );
  nand_x4_sg U62471 ( .A(n24313), .B(n24534), .X(n24532) );
  nand_x4_sg U62472 ( .A(n24318), .B(n24539), .X(n24537) );
  nand_x4_sg U62473 ( .A(n24323), .B(n24544), .X(n24542) );
  nand_x4_sg U62474 ( .A(n24328), .B(n24549), .X(n24547) );
  nand_x4_sg U62475 ( .A(n24333), .B(n24554), .X(n24552) );
  nand_x4_sg U62476 ( .A(n24338), .B(n24559), .X(n24557) );
  nand_x4_sg U62477 ( .A(n24343), .B(n24564), .X(n24562) );
  nand_x4_sg U62478 ( .A(n24348), .B(n24569), .X(n24567) );
  nand_x4_sg U62479 ( .A(n24353), .B(n24574), .X(n24572) );
  nand_x4_sg U62480 ( .A(n24358), .B(n24579), .X(n24577) );
  nand_x4_sg U62481 ( .A(n24363), .B(n24584), .X(n24582) );
  nand_x4_sg U62482 ( .A(n24376), .B(n24600), .X(n24587) );
  nor_x1_sg U62483 ( .A(n57113), .B(n26040), .X(\filter_0/n8287 ) );
  nor_x1_sg U62484 ( .A(n57113), .B(n26049), .X(\filter_0/n8279 ) );
  nor_x1_sg U62485 ( .A(n57113), .B(n26056), .X(\filter_0/n8268 ) );
  nor_x1_sg U62486 ( .A(n57113), .B(n26069), .X(\filter_0/n8259 ) );
  nor_x1_sg U62487 ( .A(n57113), .B(n26169), .X(\filter_0/n8243 ) );
  nor_x1_sg U62488 ( .A(n23645), .B(n23646), .X(\shifter_0/n11264 ) );
  nor_x1_sg U62489 ( .A(n23651), .B(n23652), .X(\shifter_0/n11260 ) );
  nor_x1_sg U62490 ( .A(n23657), .B(n23658), .X(\shifter_0/n11256 ) );
  nor_x1_sg U62491 ( .A(n23663), .B(n23664), .X(\shifter_0/n11252 ) );
  nor_x1_sg U62492 ( .A(n23669), .B(n23670), .X(\shifter_0/n11248 ) );
  nor_x1_sg U62493 ( .A(n23905), .B(n23906), .X(\shifter_0/n11104 ) );
  nor_x1_sg U62494 ( .A(n23911), .B(n23912), .X(\shifter_0/n11100 ) );
  nor_x1_sg U62495 ( .A(n23917), .B(n23918), .X(\shifter_0/n11096 ) );
  nor_x1_sg U62496 ( .A(n23923), .B(n23924), .X(\shifter_0/n11092 ) );
  nor_x1_sg U62497 ( .A(n23929), .B(n23930), .X(\shifter_0/n11088 ) );
  nor_x1_sg U62498 ( .A(n24346), .B(n24347), .X(\shifter_0/n10784 ) );
  nor_x1_sg U62499 ( .A(n24351), .B(n24352), .X(\shifter_0/n10780 ) );
  nor_x1_sg U62500 ( .A(n24356), .B(n24357), .X(\shifter_0/n10776 ) );
  nor_x1_sg U62501 ( .A(n24361), .B(n24362), .X(\shifter_0/n10772 ) );
  nor_x1_sg U62502 ( .A(n24366), .B(n24367), .X(\shifter_0/n10768 ) );
  nor_x1_sg U62503 ( .A(n24759), .B(n24760), .X(\shifter_0/n10464 ) );
  nor_x1_sg U62504 ( .A(n24763), .B(n24764), .X(\shifter_0/n10460 ) );
  nor_x1_sg U62505 ( .A(n24767), .B(n24768), .X(\shifter_0/n10456 ) );
  nor_x1_sg U62506 ( .A(n24771), .B(n24772), .X(\shifter_0/n10452 ) );
  nor_x1_sg U62507 ( .A(n24775), .B(n24776), .X(\shifter_0/n10448 ) );
  nor_x1_sg U62508 ( .A(n23429), .B(n23430), .X(\shifter_0/n11400 ) );
  nor_x1_sg U62509 ( .A(n23435), .B(n23436), .X(\shifter_0/n11396 ) );
  nor_x1_sg U62510 ( .A(n23441), .B(n23442), .X(\shifter_0/n11392 ) );
  nor_x1_sg U62511 ( .A(n23447), .B(n23448), .X(\shifter_0/n11388 ) );
  nor_x1_sg U62512 ( .A(n23453), .B(n23454), .X(\shifter_0/n11384 ) );
  nor_x1_sg U62513 ( .A(n23459), .B(n23460), .X(\shifter_0/n11380 ) );
  nor_x1_sg U62514 ( .A(n23465), .B(n23466), .X(\shifter_0/n11376 ) );
  nor_x1_sg U62515 ( .A(n23471), .B(n23472), .X(\shifter_0/n11372 ) );
  nor_x1_sg U62516 ( .A(n23477), .B(n23478), .X(\shifter_0/n11368 ) );
  nor_x1_sg U62517 ( .A(n23483), .B(n23484), .X(\shifter_0/n11364 ) );
  nor_x1_sg U62518 ( .A(n23489), .B(n23490), .X(\shifter_0/n11360 ) );
  nor_x1_sg U62519 ( .A(n23495), .B(n23496), .X(\shifter_0/n11356 ) );
  nor_x1_sg U62520 ( .A(n23501), .B(n23502), .X(\shifter_0/n11352 ) );
  nor_x1_sg U62521 ( .A(n23507), .B(n23508), .X(\shifter_0/n11348 ) );
  nor_x1_sg U62522 ( .A(n23513), .B(n23514), .X(\shifter_0/n11344 ) );
  nor_x1_sg U62523 ( .A(n23519), .B(n23520), .X(\shifter_0/n11340 ) );
  nor_x1_sg U62524 ( .A(n23525), .B(n23526), .X(\shifter_0/n11336 ) );
  nor_x1_sg U62525 ( .A(n23531), .B(n23532), .X(\shifter_0/n11332 ) );
  nor_x1_sg U62526 ( .A(n23537), .B(n23538), .X(\shifter_0/n11328 ) );
  nor_x1_sg U62527 ( .A(n23554), .B(n23555), .X(\shifter_0/n11324 ) );
  nor_x1_sg U62528 ( .A(n23561), .B(n23562), .X(\shifter_0/n11320 ) );
  nor_x1_sg U62529 ( .A(n23567), .B(n23568), .X(\shifter_0/n11316 ) );
  nor_x1_sg U62530 ( .A(n23573), .B(n23574), .X(\shifter_0/n11312 ) );
  nor_x1_sg U62531 ( .A(n23579), .B(n23580), .X(\shifter_0/n11308 ) );
  nor_x1_sg U62532 ( .A(n23585), .B(n23586), .X(\shifter_0/n11304 ) );
  nor_x1_sg U62533 ( .A(n23591), .B(n23592), .X(\shifter_0/n11300 ) );
  nor_x1_sg U62534 ( .A(n23597), .B(n23598), .X(\shifter_0/n11296 ) );
  nor_x1_sg U62535 ( .A(n23603), .B(n23604), .X(\shifter_0/n11292 ) );
  nor_x1_sg U62536 ( .A(n23609), .B(n23610), .X(\shifter_0/n11288 ) );
  nor_x1_sg U62537 ( .A(n23615), .B(n23616), .X(\shifter_0/n11284 ) );
  nor_x1_sg U62538 ( .A(n23621), .B(n23622), .X(\shifter_0/n11280 ) );
  nor_x1_sg U62539 ( .A(n23627), .B(n23628), .X(\shifter_0/n11276 ) );
  nor_x1_sg U62540 ( .A(n23633), .B(n23634), .X(\shifter_0/n11272 ) );
  nor_x1_sg U62541 ( .A(n23639), .B(n23640), .X(\shifter_0/n11268 ) );
  nor_x1_sg U62542 ( .A(n23692), .B(n23693), .X(\shifter_0/n11240 ) );
  nor_x1_sg U62543 ( .A(n23698), .B(n23699), .X(\shifter_0/n11236 ) );
  nor_x1_sg U62544 ( .A(n23704), .B(n23705), .X(\shifter_0/n11232 ) );
  nor_x1_sg U62545 ( .A(n23710), .B(n23711), .X(\shifter_0/n11228 ) );
  nor_x1_sg U62546 ( .A(n23716), .B(n23717), .X(\shifter_0/n11224 ) );
  nor_x1_sg U62547 ( .A(n23722), .B(n23723), .X(\shifter_0/n11220 ) );
  nor_x1_sg U62548 ( .A(n23728), .B(n23729), .X(\shifter_0/n11216 ) );
  nor_x1_sg U62549 ( .A(n23734), .B(n23735), .X(\shifter_0/n11212 ) );
  nor_x1_sg U62550 ( .A(n23740), .B(n23741), .X(\shifter_0/n11208 ) );
  nor_x1_sg U62551 ( .A(n23746), .B(n23747), .X(\shifter_0/n11204 ) );
  nor_x1_sg U62552 ( .A(n23752), .B(n23753), .X(\shifter_0/n11200 ) );
  nor_x1_sg U62553 ( .A(n23758), .B(n23759), .X(\shifter_0/n11196 ) );
  nor_x1_sg U62554 ( .A(n23764), .B(n23765), .X(\shifter_0/n11192 ) );
  nor_x1_sg U62555 ( .A(n23770), .B(n23771), .X(\shifter_0/n11188 ) );
  nor_x1_sg U62556 ( .A(n23776), .B(n23777), .X(\shifter_0/n11184 ) );
  nor_x1_sg U62557 ( .A(n23782), .B(n23783), .X(\shifter_0/n11180 ) );
  nor_x1_sg U62558 ( .A(n23788), .B(n23789), .X(\shifter_0/n11176 ) );
  nor_x1_sg U62559 ( .A(n23794), .B(n23795), .X(\shifter_0/n11172 ) );
  nor_x1_sg U62560 ( .A(n23800), .B(n23801), .X(\shifter_0/n11168 ) );
  nor_x1_sg U62561 ( .A(n23814), .B(n23815), .X(\shifter_0/n11164 ) );
  nor_x1_sg U62562 ( .A(n23821), .B(n23822), .X(\shifter_0/n11160 ) );
  nor_x1_sg U62563 ( .A(n23827), .B(n23828), .X(\shifter_0/n11156 ) );
  nor_x1_sg U62564 ( .A(n23833), .B(n23834), .X(\shifter_0/n11152 ) );
  nor_x1_sg U62565 ( .A(n23839), .B(n23840), .X(\shifter_0/n11148 ) );
  nor_x1_sg U62566 ( .A(n23845), .B(n23846), .X(\shifter_0/n11144 ) );
  nor_x1_sg U62567 ( .A(n23851), .B(n23852), .X(\shifter_0/n11140 ) );
  nor_x1_sg U62568 ( .A(n23857), .B(n23858), .X(\shifter_0/n11136 ) );
  nor_x1_sg U62569 ( .A(n23863), .B(n23864), .X(\shifter_0/n11132 ) );
  nor_x1_sg U62570 ( .A(n23869), .B(n23870), .X(\shifter_0/n11128 ) );
  nor_x1_sg U62571 ( .A(n23875), .B(n23876), .X(\shifter_0/n11124 ) );
  nor_x1_sg U62572 ( .A(n23881), .B(n23882), .X(\shifter_0/n11120 ) );
  nor_x1_sg U62573 ( .A(n23887), .B(n23888), .X(\shifter_0/n11116 ) );
  nor_x1_sg U62574 ( .A(n23893), .B(n23894), .X(\shifter_0/n11112 ) );
  nor_x1_sg U62575 ( .A(n23899), .B(n23900), .X(\shifter_0/n11108 ) );
  nor_x1_sg U62576 ( .A(n24167), .B(n24168), .X(\shifter_0/n10920 ) );
  nor_x1_sg U62577 ( .A(n24172), .B(n24173), .X(\shifter_0/n10916 ) );
  nor_x1_sg U62578 ( .A(n24177), .B(n24178), .X(\shifter_0/n10912 ) );
  nor_x1_sg U62579 ( .A(n24182), .B(n24183), .X(\shifter_0/n10908 ) );
  nor_x1_sg U62580 ( .A(n24187), .B(n24188), .X(\shifter_0/n10904 ) );
  nor_x1_sg U62581 ( .A(n24192), .B(n24193), .X(\shifter_0/n10900 ) );
  nor_x1_sg U62582 ( .A(n24197), .B(n24198), .X(\shifter_0/n10896 ) );
  nor_x1_sg U62583 ( .A(n24202), .B(n24203), .X(\shifter_0/n10892 ) );
  nor_x1_sg U62584 ( .A(n24207), .B(n24208), .X(\shifter_0/n10888 ) );
  nor_x1_sg U62585 ( .A(n24212), .B(n24213), .X(\shifter_0/n10884 ) );
  nor_x1_sg U62586 ( .A(n24217), .B(n24218), .X(\shifter_0/n10880 ) );
  nor_x1_sg U62587 ( .A(n24222), .B(n24223), .X(\shifter_0/n10876 ) );
  nor_x1_sg U62588 ( .A(n24227), .B(n24228), .X(\shifter_0/n10872 ) );
  nor_x1_sg U62589 ( .A(n24232), .B(n24233), .X(\shifter_0/n10868 ) );
  nor_x1_sg U62590 ( .A(n24237), .B(n24238), .X(\shifter_0/n10864 ) );
  nor_x1_sg U62591 ( .A(n24242), .B(n24243), .X(\shifter_0/n10860 ) );
  nor_x1_sg U62592 ( .A(n24247), .B(n24248), .X(\shifter_0/n10856 ) );
  nor_x1_sg U62593 ( .A(n24252), .B(n24253), .X(\shifter_0/n10852 ) );
  nor_x1_sg U62594 ( .A(n24257), .B(n24258), .X(\shifter_0/n10848 ) );
  nor_x1_sg U62595 ( .A(n24270), .B(n24271), .X(\shifter_0/n10844 ) );
  nor_x1_sg U62596 ( .A(n24276), .B(n24277), .X(\shifter_0/n10840 ) );
  nor_x1_sg U62597 ( .A(n24281), .B(n24282), .X(\shifter_0/n10836 ) );
  nor_x1_sg U62598 ( .A(n24286), .B(n24287), .X(\shifter_0/n10832 ) );
  nor_x1_sg U62599 ( .A(n24291), .B(n24292), .X(\shifter_0/n10828 ) );
  nor_x1_sg U62600 ( .A(n24296), .B(n24297), .X(\shifter_0/n10824 ) );
  nor_x1_sg U62601 ( .A(n24301), .B(n24302), .X(\shifter_0/n10820 ) );
  nor_x1_sg U62602 ( .A(n24306), .B(n24307), .X(\shifter_0/n10816 ) );
  nor_x1_sg U62603 ( .A(n24311), .B(n24312), .X(\shifter_0/n10812 ) );
  nor_x1_sg U62604 ( .A(n24316), .B(n24317), .X(\shifter_0/n10808 ) );
  nor_x1_sg U62605 ( .A(n24321), .B(n24322), .X(\shifter_0/n10804 ) );
  nor_x1_sg U62606 ( .A(n24326), .B(n24327), .X(\shifter_0/n10800 ) );
  nor_x1_sg U62607 ( .A(n24331), .B(n24332), .X(\shifter_0/n10796 ) );
  nor_x1_sg U62608 ( .A(n24336), .B(n24337), .X(\shifter_0/n10792 ) );
  nor_x1_sg U62609 ( .A(n24341), .B(n24342), .X(\shifter_0/n10788 ) );
  nor_x1_sg U62610 ( .A(n24609), .B(n24610), .X(\shifter_0/n10600 ) );
  nor_x1_sg U62611 ( .A(n24613), .B(n24614), .X(\shifter_0/n10596 ) );
  nor_x1_sg U62612 ( .A(n24617), .B(n24618), .X(\shifter_0/n10592 ) );
  nor_x1_sg U62613 ( .A(n24621), .B(n24622), .X(\shifter_0/n10588 ) );
  nor_x1_sg U62614 ( .A(n24625), .B(n24626), .X(\shifter_0/n10584 ) );
  nor_x1_sg U62615 ( .A(n24629), .B(n24630), .X(\shifter_0/n10580 ) );
  nor_x1_sg U62616 ( .A(n24633), .B(n24634), .X(\shifter_0/n10576 ) );
  nor_x1_sg U62617 ( .A(n24637), .B(n24638), .X(\shifter_0/n10572 ) );
  nor_x1_sg U62618 ( .A(n24641), .B(n24642), .X(\shifter_0/n10568 ) );
  nor_x1_sg U62619 ( .A(n24645), .B(n24646), .X(\shifter_0/n10564 ) );
  nor_x1_sg U62620 ( .A(n24649), .B(n24650), .X(\shifter_0/n10560 ) );
  nor_x1_sg U62621 ( .A(n24653), .B(n24654), .X(\shifter_0/n10556 ) );
  nor_x1_sg U62622 ( .A(n24657), .B(n24658), .X(\shifter_0/n10552 ) );
  nor_x1_sg U62623 ( .A(n24661), .B(n24662), .X(\shifter_0/n10548 ) );
  nor_x1_sg U62624 ( .A(n24665), .B(n24666), .X(\shifter_0/n10544 ) );
  nor_x1_sg U62625 ( .A(n24669), .B(n24670), .X(\shifter_0/n10540 ) );
  nor_x1_sg U62626 ( .A(n24673), .B(n24674), .X(\shifter_0/n10536 ) );
  nor_x1_sg U62627 ( .A(n24677), .B(n24678), .X(\shifter_0/n10532 ) );
  nor_x1_sg U62628 ( .A(n24681), .B(n24682), .X(\shifter_0/n10528 ) );
  nor_x1_sg U62629 ( .A(n24698), .B(n24699), .X(\shifter_0/n10524 ) );
  nor_x1_sg U62630 ( .A(n24703), .B(n24704), .X(\shifter_0/n10520 ) );
  nor_x1_sg U62631 ( .A(n24707), .B(n24708), .X(\shifter_0/n10516 ) );
  nor_x1_sg U62632 ( .A(n24711), .B(n24712), .X(\shifter_0/n10512 ) );
  nor_x1_sg U62633 ( .A(n24715), .B(n24716), .X(\shifter_0/n10508 ) );
  nor_x1_sg U62634 ( .A(n24719), .B(n24720), .X(\shifter_0/n10504 ) );
  nor_x1_sg U62635 ( .A(n24723), .B(n24724), .X(\shifter_0/n10500 ) );
  nor_x1_sg U62636 ( .A(n24727), .B(n24728), .X(\shifter_0/n10496 ) );
  nor_x1_sg U62637 ( .A(n24731), .B(n24732), .X(\shifter_0/n10492 ) );
  nor_x1_sg U62638 ( .A(n24735), .B(n24736), .X(\shifter_0/n10488 ) );
  nor_x1_sg U62639 ( .A(n24739), .B(n24740), .X(\shifter_0/n10484 ) );
  nor_x1_sg U62640 ( .A(n24743), .B(n24744), .X(\shifter_0/n10480 ) );
  nor_x1_sg U62641 ( .A(n24747), .B(n24748), .X(\shifter_0/n10476 ) );
  nor_x1_sg U62642 ( .A(n24751), .B(n24752), .X(\shifter_0/n10472 ) );
  nor_x1_sg U62643 ( .A(n24755), .B(n24756), .X(\shifter_0/n10468 ) );
  nor_x1_sg U62644 ( .A(n23420), .B(n23421), .X(\shifter_0/n11404 ) );
  nor_x1_sg U62645 ( .A(n23684), .B(n23685), .X(\shifter_0/n11244 ) );
  nor_x1_sg U62646 ( .A(n24161), .B(n24162), .X(\shifter_0/n10924 ) );
  nor_x1_sg U62647 ( .A(n24603), .B(n24604), .X(\shifter_0/n10604 ) );
  nor_x1_sg U62648 ( .A(n57165), .B(n22654), .X(\shifter_0/n11884 ) );
  nor_x1_sg U62649 ( .A(n57165), .B(n22656), .X(\shifter_0/n11880 ) );
  nor_x1_sg U62650 ( .A(n57165), .B(n22660), .X(\shifter_0/n11872 ) );
  nor_x1_sg U62651 ( .A(n57165), .B(n22662), .X(\shifter_0/n11868 ) );
  nor_x1_sg U62652 ( .A(n57165), .B(n22666), .X(\shifter_0/n11860 ) );
  nor_x1_sg U62653 ( .A(n57165), .B(n22668), .X(\shifter_0/n11856 ) );
  nor_x1_sg U62654 ( .A(n57165), .B(n22672), .X(\shifter_0/n11848 ) );
  nor_x1_sg U62655 ( .A(n57165), .B(n22674), .X(\shifter_0/n11844 ) );
  nor_x1_sg U62656 ( .A(n57165), .B(n22678), .X(\shifter_0/n11836 ) );
  nor_x1_sg U62657 ( .A(n57165), .B(n22680), .X(\shifter_0/n11832 ) );
  nor_x1_sg U62658 ( .A(n57165), .B(n22684), .X(\shifter_0/n11824 ) );
  nor_x1_sg U62659 ( .A(n57165), .B(n22686), .X(\shifter_0/n11820 ) );
  nor_x1_sg U62660 ( .A(n57165), .B(n22690), .X(\shifter_0/n11812 ) );
  nor_x1_sg U62661 ( .A(n57165), .B(n22692), .X(\shifter_0/n11808 ) );
  nor_x1_sg U62662 ( .A(n57162), .B(n22701), .X(\shifter_0/n11804 ) );
  nor_x1_sg U62663 ( .A(n57162), .B(n22703), .X(\shifter_0/n11800 ) );
  nor_x1_sg U62664 ( .A(n57162), .B(n22707), .X(\shifter_0/n11792 ) );
  nor_x1_sg U62665 ( .A(n57162), .B(n22709), .X(\shifter_0/n11788 ) );
  nor_x1_sg U62666 ( .A(n57162), .B(n22713), .X(\shifter_0/n11780 ) );
  nor_x1_sg U62667 ( .A(n57162), .B(n22715), .X(\shifter_0/n11776 ) );
  nor_x1_sg U62668 ( .A(n57162), .B(n22719), .X(\shifter_0/n11768 ) );
  nor_x1_sg U62669 ( .A(n57162), .B(n22721), .X(\shifter_0/n11764 ) );
  nor_x1_sg U62670 ( .A(n57162), .B(n22725), .X(\shifter_0/n11756 ) );
  nor_x1_sg U62671 ( .A(n57162), .B(n22727), .X(\shifter_0/n11752 ) );
  nor_x1_sg U62672 ( .A(n57162), .B(n22731), .X(\shifter_0/n11744 ) );
  nor_x1_sg U62673 ( .A(n57162), .B(n22733), .X(\shifter_0/n11740 ) );
  nor_x1_sg U62674 ( .A(n57162), .B(n22737), .X(\shifter_0/n11732 ) );
  nor_x1_sg U62675 ( .A(n57162), .B(n22739), .X(\shifter_0/n11728 ) );
  nor_x1_sg U62676 ( .A(n57165), .B(n22658), .X(\shifter_0/n11876 ) );
  nor_x1_sg U62677 ( .A(n57165), .B(n22664), .X(\shifter_0/n11864 ) );
  nor_x1_sg U62678 ( .A(n57165), .B(n22670), .X(\shifter_0/n11852 ) );
  nor_x1_sg U62679 ( .A(n57165), .B(n22676), .X(\shifter_0/n11840 ) );
  nor_x1_sg U62680 ( .A(n57165), .B(n22682), .X(\shifter_0/n11828 ) );
  nor_x1_sg U62681 ( .A(n57165), .B(n22688), .X(\shifter_0/n11816 ) );
  nor_x1_sg U62682 ( .A(n57162), .B(n22705), .X(\shifter_0/n11796 ) );
  nor_x1_sg U62683 ( .A(n57162), .B(n22711), .X(\shifter_0/n11784 ) );
  nor_x1_sg U62684 ( .A(n57162), .B(n22717), .X(\shifter_0/n11772 ) );
  nor_x1_sg U62685 ( .A(n57162), .B(n22723), .X(\shifter_0/n11760 ) );
  nor_x1_sg U62686 ( .A(n57162), .B(n22729), .X(\shifter_0/n11748 ) );
  nor_x1_sg U62687 ( .A(n57162), .B(n22735), .X(\shifter_0/n11736 ) );
  nor_x1_sg U62688 ( .A(n22446), .B(n22465), .X(\shifter_0/n12452 ) );
  nor_x1_sg U62689 ( .A(n22446), .B(n22466), .X(\shifter_0/n12448 ) );
  nor_x1_sg U62690 ( .A(n22498), .B(n22517), .X(\shifter_0/n12292 ) );
  nor_x1_sg U62691 ( .A(n22498), .B(n22518), .X(\shifter_0/n12288 ) );
  nor_x1_sg U62692 ( .A(n22473), .B(n22492), .X(\shifter_0/n12372 ) );
  nor_x1_sg U62693 ( .A(n22473), .B(n22493), .X(\shifter_0/n12368 ) );
  nor_x1_sg U62694 ( .A(n22523), .B(n22542), .X(\shifter_0/n12212 ) );
  nor_x1_sg U62695 ( .A(n22523), .B(n22543), .X(\shifter_0/n12208 ) );
  nor_x1_sg U62696 ( .A(n22396), .B(n22415), .X(\shifter_0/n12612 ) );
  nor_x1_sg U62697 ( .A(n22396), .B(n22416), .X(\shifter_0/n12608 ) );
  nor_x1_sg U62698 ( .A(n22421), .B(n22440), .X(\shifter_0/n12532 ) );
  nor_x1_sg U62699 ( .A(n22421), .B(n22441), .X(\shifter_0/n12528 ) );
  nor_x1_sg U62700 ( .A(n57510), .B(n22565), .X(\shifter_0/n12132 ) );
  nor_x1_sg U62701 ( .A(n57510), .B(n22566), .X(\shifter_0/n12128 ) );
  nor_x1_sg U62702 ( .A(n57507), .B(n22616), .X(\shifter_0/n11972 ) );
  nor_x1_sg U62703 ( .A(n57507), .B(n22617), .X(\shifter_0/n11968 ) );
  nor_x1_sg U62704 ( .A(n57516), .B(n22591), .X(\shifter_0/n12052 ) );
  nor_x1_sg U62705 ( .A(n57516), .B(n22592), .X(\shifter_0/n12048 ) );
  nor_x1_sg U62706 ( .A(n57513), .B(n22643), .X(\shifter_0/n11892 ) );
  nor_x1_sg U62707 ( .A(n57513), .B(n22644), .X(\shifter_0/n11888 ) );
  nand_x2_sg U62708 ( .A(n26141), .B(n67563), .X(n26137) );
  nor_x1_sg U62709 ( .A(n26150), .B(n67561), .X(n26141) );
  nor_x1_sg U62710 ( .A(n26143), .B(n57308), .X(n26142) );
  nand_x2_sg U62711 ( .A(n26102), .B(n67557), .X(n26098) );
  nor_x1_sg U62712 ( .A(n26111), .B(n67555), .X(n26102) );
  nor_x1_sg U62713 ( .A(n26104), .B(n57308), .X(n26103) );
  nand_x2_sg U62714 ( .A(n26233), .B(n67551), .X(n26229) );
  nor_x1_sg U62715 ( .A(n26242), .B(n67549), .X(n26233) );
  nor_x1_sg U62716 ( .A(n26235), .B(n57308), .X(n26234) );
  nand_x2_sg U62717 ( .A(n26199), .B(n67545), .X(n26195) );
  nor_x1_sg U62718 ( .A(n26208), .B(n67543), .X(n26199) );
  nor_x1_sg U62719 ( .A(n26201), .B(n57308), .X(n26200) );
  nand_x1_sg U62720 ( .A(n67234), .B(n57468), .X(n23222) );
  nand_x1_sg U62721 ( .A(n67232), .B(n57468), .X(n23227) );
  nand_x1_sg U62722 ( .A(n67224), .B(n57468), .X(n23247) );
  nand_x1_sg U62723 ( .A(n67222), .B(n57468), .X(n23252) );
  nand_x1_sg U62724 ( .A(n67216), .B(n57468), .X(n23267) );
  nand_x1_sg U62725 ( .A(n67214), .B(n57468), .X(n23272) );
  nand_x1_sg U62726 ( .A(n67206), .B(n57468), .X(n23292) );
  nand_x1_sg U62727 ( .A(n67204), .B(n57468), .X(n23297) );
  nand_x1_sg U62728 ( .A(n67427), .B(n57476), .X(n23330) );
  nand_x1_sg U62729 ( .A(n67425), .B(n57476), .X(n23335) );
  nand_x1_sg U62730 ( .A(n67417), .B(n57476), .X(n23355) );
  nand_x1_sg U62731 ( .A(n67415), .B(n57476), .X(n23360) );
  nand_x1_sg U62732 ( .A(n67409), .B(n57476), .X(n23375) );
  nand_x1_sg U62733 ( .A(n67407), .B(n57476), .X(n23380) );
  nand_x1_sg U62734 ( .A(n67399), .B(n57476), .X(n23400) );
  nand_x1_sg U62735 ( .A(n67397), .B(n57476), .X(n23405) );
  nand_x1_sg U62736 ( .A(n57484), .B(n67240), .X(n23947) );
  nand_x1_sg U62737 ( .A(n57484), .B(n67238), .X(n23952) );
  nand_x1_sg U62738 ( .A(n57484), .B(n67236), .X(n23957) );
  nand_x1_sg U62739 ( .A(n57484), .B(n67234), .X(n23962) );
  nand_x1_sg U62740 ( .A(n57484), .B(n67232), .X(n23967) );
  nand_x1_sg U62741 ( .A(n57484), .B(n67230), .X(n23972) );
  nand_x1_sg U62742 ( .A(n57484), .B(n67228), .X(n23977) );
  nand_x1_sg U62743 ( .A(n57484), .B(n67226), .X(n23982) );
  nand_x1_sg U62744 ( .A(n57484), .B(n67224), .X(n23987) );
  nand_x1_sg U62745 ( .A(n57484), .B(n67222), .X(n23992) );
  nand_x1_sg U62746 ( .A(n57484), .B(n67220), .X(n23997) );
  nand_x1_sg U62747 ( .A(n57484), .B(n67218), .X(n24002) );
  nand_x1_sg U62748 ( .A(n57484), .B(n67216), .X(n24007) );
  nand_x1_sg U62749 ( .A(n57484), .B(n67214), .X(n24012) );
  nand_x1_sg U62750 ( .A(n57484), .B(n67212), .X(n24017) );
  nand_x1_sg U62751 ( .A(n57484), .B(n67210), .X(n24022) );
  nand_x1_sg U62752 ( .A(n57484), .B(n67208), .X(n24027) );
  nand_x1_sg U62753 ( .A(n57484), .B(n67206), .X(n24032) );
  nand_x1_sg U62754 ( .A(n57484), .B(n67204), .X(n24037) );
  nand_x1_sg U62755 ( .A(n57484), .B(n67202), .X(n24042) );
  nand_x1_sg U62756 ( .A(n57492), .B(n67433), .X(n24057) );
  nand_x1_sg U62757 ( .A(n57492), .B(n67431), .X(n24062) );
  nand_x1_sg U62758 ( .A(n57492), .B(n67429), .X(n24067) );
  nand_x1_sg U62759 ( .A(n57492), .B(n67427), .X(n24072) );
  nand_x1_sg U62760 ( .A(n57492), .B(n67425), .X(n24077) );
  nand_x1_sg U62761 ( .A(n57492), .B(n67423), .X(n24082) );
  nand_x1_sg U62762 ( .A(n57492), .B(n67421), .X(n24087) );
  nand_x1_sg U62763 ( .A(n57492), .B(n67419), .X(n24092) );
  nand_x1_sg U62764 ( .A(n57492), .B(n67417), .X(n24097) );
  nand_x1_sg U62765 ( .A(n57492), .B(n67415), .X(n24102) );
  nand_x1_sg U62766 ( .A(n57492), .B(n67413), .X(n24107) );
  nand_x1_sg U62767 ( .A(n57492), .B(n67411), .X(n24112) );
  nand_x1_sg U62768 ( .A(n57492), .B(n67409), .X(n24117) );
  nand_x1_sg U62769 ( .A(n57492), .B(n67407), .X(n24122) );
  nand_x1_sg U62770 ( .A(n57492), .B(n67405), .X(n24127) );
  nand_x1_sg U62771 ( .A(n57492), .B(n67403), .X(n24132) );
  nand_x1_sg U62772 ( .A(n57492), .B(n67401), .X(n24137) );
  nand_x1_sg U62773 ( .A(n57492), .B(n67399), .X(n24142) );
  nand_x1_sg U62774 ( .A(n57492), .B(n67397), .X(n24147) );
  nand_x1_sg U62775 ( .A(n57492), .B(n67395), .X(n24152) );
  nand_x1_sg U62776 ( .A(n51051), .B(n67536), .X(n26285) );
  nand_x1_sg U62777 ( .A(n50727), .B(n57199), .X(n33879) );
  nand_x1_sg U62778 ( .A(n50725), .B(n57199), .X(n33889) );
  nand_x1_sg U62779 ( .A(n50723), .B(n57199), .X(n33891) );
  nand_x1_sg U62780 ( .A(n53251), .B(n57199), .X(n33883) );
  nand_x1_sg U62781 ( .A(n50721), .B(n57199), .X(n33869) );
  nand_x1_sg U62782 ( .A(n50719), .B(n33872), .X(n33873) );
  nand_x1_sg U62783 ( .A(n50717), .B(n57199), .X(n33893) );
  nand_x1_sg U62784 ( .A(n50713), .B(n57199), .X(n33897) );
  nand_x1_sg U62785 ( .A(n50711), .B(n57199), .X(n33875) );
  nand_x1_sg U62786 ( .A(n50709), .B(n57199), .X(n33899) );
  nand_x1_sg U62787 ( .A(n50707), .B(n57199), .X(n33881) );
  nand_x1_sg U62788 ( .A(n53249), .B(n57199), .X(n33901) );
  nand_x1_sg U62789 ( .A(n53247), .B(n57199), .X(n33907) );
  nand_x1_sg U62790 ( .A(n53245), .B(n57199), .X(n33909) );
  nand_x1_sg U62791 ( .A(n50999), .B(n57176), .X(n34156) );
  nand_x1_sg U62792 ( .A(n50997), .B(n57176), .X(n34136) );
  nand_x1_sg U62793 ( .A(n50995), .B(n57176), .X(n34146) );
  nand_x1_sg U62794 ( .A(n53581), .B(n57176), .X(n34160) );
  nand_x1_sg U62795 ( .A(n53579), .B(n57176), .X(n34144) );
  nand_x1_sg U62796 ( .A(n50991), .B(n34135), .X(n34154) );
  nand_x1_sg U62797 ( .A(n50989), .B(n57176), .X(n34162) );
  nand_x1_sg U62798 ( .A(n53577), .B(n57176), .X(n34164) );
  nand_x1_sg U62799 ( .A(n50983), .B(n57176), .X(n34132) );
  nand_x1_sg U62800 ( .A(n53575), .B(n57176), .X(n34152) );
  nand_x1_sg U62801 ( .A(n53573), .B(n57176), .X(n34170) );
  nand_x1_sg U62802 ( .A(n50981), .B(n57176), .X(n34142) );
  nand_x1_sg U62803 ( .A(n50977), .B(n57176), .X(n34138) );
  nand_x1_sg U62804 ( .A(n53571), .B(n57176), .X(n34172) );
  nand_x1_sg U62805 ( .A(n52957), .B(n57183), .X(n34044) );
  nand_x1_sg U62806 ( .A(n52955), .B(n57183), .X(n34064) );
  nand_x1_sg U62807 ( .A(n52953), .B(n57183), .X(n34066) );
  nand_x1_sg U62808 ( .A(n50461), .B(n57183), .X(n34058) );
  nand_x1_sg U62809 ( .A(n52951), .B(n57183), .X(n34056) );
  nand_x1_sg U62810 ( .A(n50459), .B(n57183), .X(n34050) );
  nand_x1_sg U62811 ( .A(n52949), .B(n57183), .X(n34068) );
  nand_x1_sg U62812 ( .A(n52947), .B(n57183), .X(n34072) );
  nand_x1_sg U62813 ( .A(n50455), .B(n57183), .X(n34074) );
  nand_x1_sg U62814 ( .A(n52945), .B(n57183), .X(n34076) );
  nand_x1_sg U62815 ( .A(n50453), .B(n34047), .X(n34048) );
  nand_x1_sg U62816 ( .A(n50449), .B(n57183), .X(n34054) );
  nand_x1_sg U62817 ( .A(n52939), .B(n57183), .X(n34082) );
  nand_x1_sg U62818 ( .A(n52937), .B(n57183), .X(n34084) );
  nand_x1_sg U62819 ( .A(n51003), .B(n67536), .X(n26321) );
  nand_x1_sg U62820 ( .A(n50641), .B(n57172), .X(n34201) );
  nand_x1_sg U62821 ( .A(n50639), .B(n57172), .X(n34181) );
  nand_x1_sg U62822 ( .A(n50637), .B(n57172), .X(n34205) );
  nand_x1_sg U62823 ( .A(n50635), .B(n57172), .X(n34207) );
  nand_x1_sg U62824 ( .A(n53179), .B(n57172), .X(n34189) );
  nand_x1_sg U62825 ( .A(n50633), .B(n57172), .X(n34199) );
  nand_x1_sg U62826 ( .A(n50631), .B(n57172), .X(n34191) );
  nand_x1_sg U62827 ( .A(n50629), .B(n57172), .X(n34209) );
  nand_x1_sg U62828 ( .A(n50623), .B(n34180), .X(n34177) );
  nand_x1_sg U62829 ( .A(n53175), .B(n57172), .X(n34197) );
  nand_x1_sg U62830 ( .A(n50621), .B(n57172), .X(n34187) );
  nand_x1_sg U62831 ( .A(n53171), .B(n57172), .X(n34183) );
  nand_x1_sg U62832 ( .A(n53169), .B(n57172), .X(n34215) );
  nand_x1_sg U62833 ( .A(n53167), .B(n57172), .X(n34217) );
  nand_x2_sg U62834 ( .A(n26272), .B(n26273), .X(n26271) );
  nand_x1_sg U62835 ( .A(n26085), .B(n67565), .X(n26272) );
  nand_x1_sg U62836 ( .A(n47341), .B(n26043), .X(n26273) );
  nand_x1_sg U62837 ( .A(n50731), .B(n57199), .X(n33877) );
  nand_x1_sg U62838 ( .A(n50729), .B(n57199), .X(n33885) );
  nand_x1_sg U62839 ( .A(n50715), .B(n57199), .X(n33895) );
  nand_x1_sg U62840 ( .A(n50705), .B(n57199), .X(n33903) );
  nand_x1_sg U62841 ( .A(n50703), .B(n57199), .X(n33887) );
  nand_x1_sg U62842 ( .A(n50701), .B(n57199), .X(n33905) );
  nand_x1_sg U62843 ( .A(n53583), .B(n57176), .X(n34140) );
  nand_x1_sg U62844 ( .A(n50993), .B(n57176), .X(n34150) );
  nand_x1_sg U62845 ( .A(n50987), .B(n57176), .X(n34166) );
  nand_x1_sg U62846 ( .A(n50985), .B(n57176), .X(n34168) );
  nand_x1_sg U62847 ( .A(n50979), .B(n57176), .X(n34158) );
  nand_x1_sg U62848 ( .A(n53569), .B(n57176), .X(n34148) );
  nand_x1_sg U62849 ( .A(n50643), .B(n57172), .X(n34185) );
  nand_x1_sg U62850 ( .A(n53177), .B(n57172), .X(n34195) );
  nand_x1_sg U62851 ( .A(n50627), .B(n57172), .X(n34211) );
  nand_x1_sg U62852 ( .A(n50625), .B(n57172), .X(n34193) );
  nand_x1_sg U62853 ( .A(n53173), .B(n57172), .X(n34213) );
  nand_x1_sg U62854 ( .A(n50619), .B(n57172), .X(n34203) );
  nand_x1_sg U62855 ( .A(n52959), .B(n57183), .X(n34052) );
  nand_x1_sg U62856 ( .A(n50463), .B(n57183), .X(n34060) );
  nand_x1_sg U62857 ( .A(n50457), .B(n57183), .X(n34070) );
  nand_x1_sg U62858 ( .A(n52943), .B(n57183), .X(n34078) );
  nand_x1_sg U62859 ( .A(n52941), .B(n57183), .X(n34080) );
  nand_x1_sg U62860 ( .A(n50451), .B(n57183), .X(n34062) );
  nand_x1_sg U62861 ( .A(n47339), .B(n26043), .X(n26309) );
  nand_x1_sg U62862 ( .A(n53297), .B(n33787), .X(n33784) );
  nand_x1_sg U62863 ( .A(n53293), .B(n33787), .X(n33806) );
  nand_x1_sg U62864 ( .A(n50761), .B(n33787), .X(n33798) );
  nand_x1_sg U62865 ( .A(n50759), .B(n33787), .X(n33790) );
  nand_x1_sg U62866 ( .A(n50755), .B(n33787), .X(n33814) );
  nand_x1_sg U62867 ( .A(n50749), .B(n33787), .X(n33794) );
  nand_x1_sg U62868 ( .A(n53279), .B(n33787), .X(n33822) );
  nand_x1_sg U62869 ( .A(n53055), .B(n33528), .X(n33535) );
  nand_x1_sg U62870 ( .A(n50523), .B(n33528), .X(n33547) );
  nand_x1_sg U62871 ( .A(n53051), .B(n33528), .X(n33539) );
  nand_x1_sg U62872 ( .A(n50521), .B(n33528), .X(n33525) );
  nand_x1_sg U62873 ( .A(n53045), .B(n33528), .X(n33531) );
  nand_x1_sg U62874 ( .A(n50515), .B(n33528), .X(n33555) );
  nand_x1_sg U62875 ( .A(n53035), .B(n33528), .X(n33563) );
  nand_x1_sg U62876 ( .A(n53295), .B(n57205), .X(n33804) );
  nand_x1_sg U62877 ( .A(n53291), .B(n57205), .X(n33796) );
  nand_x1_sg U62878 ( .A(n53289), .B(n57205), .X(n33808) );
  nand_x1_sg U62879 ( .A(n53287), .B(n57205), .X(n33812) );
  nand_x1_sg U62880 ( .A(n53285), .B(n57205), .X(n33816) );
  nand_x1_sg U62881 ( .A(n50753), .B(n57205), .X(n33788) );
  nand_x1_sg U62882 ( .A(n53277), .B(n57205), .X(n33824) );
  nand_x1_sg U62883 ( .A(n53053), .B(n57227), .X(n33545) );
  nand_x1_sg U62884 ( .A(n53049), .B(n57227), .X(n33529) );
  nand_x1_sg U62885 ( .A(n50519), .B(n57227), .X(n33549) );
  nand_x1_sg U62886 ( .A(n50517), .B(n57227), .X(n33553) );
  nand_x1_sg U62887 ( .A(n53043), .B(n57227), .X(n33537) );
  nand_x1_sg U62888 ( .A(n53041), .B(n57227), .X(n33557) );
  nand_x1_sg U62889 ( .A(n53033), .B(n57227), .X(n33565) );
  nand_x1_sg U62890 ( .A(n50743), .B(n57202), .X(n33846) );
  nand_x1_sg U62891 ( .A(n53269), .B(n57202), .X(n33830) );
  nand_x1_sg U62892 ( .A(n50739), .B(n57202), .X(n33850) );
  nand_x1_sg U62893 ( .A(n50737), .B(n57202), .X(n33854) );
  nand_x1_sg U62894 ( .A(n53263), .B(n57202), .X(n33838) );
  nand_x1_sg U62895 ( .A(n53261), .B(n57202), .X(n33858) );
  nand_x1_sg U62896 ( .A(n53253), .B(n57202), .X(n33866) );
  nand_x1_sg U62897 ( .A(n53029), .B(n57179), .X(n34109) );
  nand_x1_sg U62898 ( .A(n50505), .B(n57179), .X(n34101) );
  nand_x1_sg U62899 ( .A(n50503), .B(n57179), .X(n34113) );
  nand_x1_sg U62900 ( .A(n50501), .B(n57179), .X(n34117) );
  nand_x1_sg U62901 ( .A(n50499), .B(n57179), .X(n34121) );
  nand_x1_sg U62902 ( .A(n53019), .B(n57179), .X(n34093) );
  nand_x1_sg U62903 ( .A(n53009), .B(n57179), .X(n34129) );
  nand_x1_sg U62904 ( .A(n53275), .B(n33829), .X(n33836) );
  nand_x1_sg U62905 ( .A(n53273), .B(n33829), .X(n33848) );
  nand_x1_sg U62906 ( .A(n53271), .B(n33829), .X(n33840) );
  nand_x1_sg U62907 ( .A(n50741), .B(n33829), .X(n33826) );
  nand_x1_sg U62908 ( .A(n53265), .B(n33829), .X(n33832) );
  nand_x1_sg U62909 ( .A(n50735), .B(n33829), .X(n33856) );
  nand_x1_sg U62910 ( .A(n53255), .B(n33829), .X(n33864) );
  nand_x1_sg U62911 ( .A(n53031), .B(n34092), .X(n34089) );
  nand_x1_sg U62912 ( .A(n50507), .B(n34092), .X(n34111) );
  nand_x1_sg U62913 ( .A(n53027), .B(n34092), .X(n34103) );
  nand_x1_sg U62914 ( .A(n53025), .B(n34092), .X(n34095) );
  nand_x1_sg U62915 ( .A(n53021), .B(n34092), .X(n34119) );
  nand_x1_sg U62916 ( .A(n53013), .B(n34092), .X(n34099) );
  nand_x1_sg U62917 ( .A(n53011), .B(n34092), .X(n34127) );
  nand_x1_sg U62918 ( .A(n50779), .B(n57209), .X(n33739) );
  nand_x1_sg U62919 ( .A(n53319), .B(n57209), .X(n33759) );
  nand_x1_sg U62920 ( .A(n50777), .B(n57209), .X(n33761) );
  nand_x1_sg U62921 ( .A(n53317), .B(n57209), .X(n33753) );
  nand_x1_sg U62922 ( .A(n53315), .B(n57209), .X(n33751) );
  nand_x1_sg U62923 ( .A(n50775), .B(n57209), .X(n33745) );
  nand_x1_sg U62924 ( .A(n53313), .B(n57209), .X(n33763) );
  nand_x1_sg U62925 ( .A(n53311), .B(n57209), .X(n33767) );
  nand_x1_sg U62926 ( .A(n50771), .B(n57209), .X(n33769) );
  nand_x1_sg U62927 ( .A(n53309), .B(n57209), .X(n33771) );
  nand_x1_sg U62928 ( .A(n50769), .B(n33742), .X(n33743) );
  nand_x1_sg U62929 ( .A(n50765), .B(n57209), .X(n33749) );
  nand_x1_sg U62930 ( .A(n53303), .B(n57209), .X(n33777) );
  nand_x1_sg U62931 ( .A(n53301), .B(n57209), .X(n33779) );
  nand_x1_sg U62932 ( .A(n50479), .B(n57187), .X(n33999) );
  nand_x1_sg U62933 ( .A(n52979), .B(n57187), .X(n34019) );
  nand_x1_sg U62934 ( .A(n50477), .B(n57187), .X(n34021) );
  nand_x1_sg U62935 ( .A(n52977), .B(n57187), .X(n34013) );
  nand_x1_sg U62936 ( .A(n52975), .B(n57187), .X(n34011) );
  nand_x1_sg U62937 ( .A(n50475), .B(n57187), .X(n34005) );
  nand_x1_sg U62938 ( .A(n52973), .B(n57187), .X(n34023) );
  nand_x1_sg U62939 ( .A(n52971), .B(n57187), .X(n34027) );
  nand_x1_sg U62940 ( .A(n50471), .B(n57187), .X(n34029) );
  nand_x1_sg U62941 ( .A(n52969), .B(n57187), .X(n34031) );
  nand_x1_sg U62942 ( .A(n50469), .B(n34002), .X(n34003) );
  nand_x1_sg U62943 ( .A(n50465), .B(n57187), .X(n34009) );
  nand_x1_sg U62944 ( .A(n52963), .B(n57187), .X(n34037) );
  nand_x1_sg U62945 ( .A(n52961), .B(n57187), .X(n34039) );
  nand_x1_sg U62946 ( .A(n53299), .B(n57205), .X(n33792) );
  nand_x1_sg U62947 ( .A(n50763), .B(n57205), .X(n33800) );
  nand_x1_sg U62948 ( .A(n53281), .B(n57205), .X(n33820) );
  nand_x1_sg U62949 ( .A(n50527), .B(n57227), .X(n33533) );
  nand_x1_sg U62950 ( .A(n50525), .B(n57227), .X(n33541) );
  nand_x1_sg U62951 ( .A(n53037), .B(n57227), .X(n33561) );
  nand_x1_sg U62952 ( .A(n50757), .B(n33787), .X(n33810) );
  nand_x1_sg U62953 ( .A(n53283), .B(n33787), .X(n33818) );
  nand_x1_sg U62954 ( .A(n50751), .B(n33787), .X(n33802) );
  nand_x1_sg U62955 ( .A(n53047), .B(n33528), .X(n33551) );
  nand_x1_sg U62956 ( .A(n50513), .B(n33528), .X(n33559) );
  nand_x1_sg U62957 ( .A(n53039), .B(n33528), .X(n33543) );
  nand_x1_sg U62958 ( .A(n53267), .B(n33829), .X(n33852) );
  nand_x1_sg U62959 ( .A(n50733), .B(n33829), .X(n33860) );
  nand_x1_sg U62960 ( .A(n53259), .B(n33829), .X(n33844) );
  nand_x1_sg U62961 ( .A(n53023), .B(n34092), .X(n34115) );
  nand_x1_sg U62962 ( .A(n53017), .B(n34092), .X(n34123) );
  nand_x1_sg U62963 ( .A(n53015), .B(n34092), .X(n34107) );
  nand_x1_sg U62964 ( .A(n53323), .B(n57209), .X(n33747) );
  nand_x1_sg U62965 ( .A(n53321), .B(n57209), .X(n33755) );
  nand_x1_sg U62966 ( .A(n50773), .B(n57209), .X(n33765) );
  nand_x1_sg U62967 ( .A(n53307), .B(n57209), .X(n33773) );
  nand_x1_sg U62968 ( .A(n53305), .B(n57209), .X(n33775) );
  nand_x1_sg U62969 ( .A(n50767), .B(n57209), .X(n33757) );
  nand_x1_sg U62970 ( .A(n50747), .B(n57202), .X(n33834) );
  nand_x1_sg U62971 ( .A(n50745), .B(n57202), .X(n33842) );
  nand_x1_sg U62972 ( .A(n53257), .B(n57202), .X(n33862) );
  nand_x1_sg U62973 ( .A(n50511), .B(n57179), .X(n34097) );
  nand_x1_sg U62974 ( .A(n50509), .B(n57179), .X(n34105) );
  nand_x1_sg U62975 ( .A(n50497), .B(n57179), .X(n34125) );
  nand_x1_sg U62976 ( .A(n52983), .B(n57187), .X(n34007) );
  nand_x1_sg U62977 ( .A(n52981), .B(n57187), .X(n34015) );
  nand_x1_sg U62978 ( .A(n50473), .B(n57187), .X(n34025) );
  nand_x1_sg U62979 ( .A(n52967), .B(n57187), .X(n34033) );
  nand_x1_sg U62980 ( .A(n52965), .B(n57187), .X(n34035) );
  nand_x1_sg U62981 ( .A(n50467), .B(n57187), .X(n34017) );
  nand_x1_sg U62982 ( .A(n53475), .B(n57224), .X(n33587) );
  nand_x1_sg U62983 ( .A(n53469), .B(n57224), .X(n33571) );
  nand_x1_sg U62984 ( .A(n53467), .B(n57224), .X(n33591) );
  nand_x1_sg U62985 ( .A(n53465), .B(n57224), .X(n33595) );
  nand_x1_sg U62986 ( .A(n50897), .B(n57224), .X(n33579) );
  nand_x1_sg U62987 ( .A(n53459), .B(n57224), .X(n33599) );
  nand_x1_sg U62988 ( .A(n53451), .B(n57224), .X(n33607) );
  nand_x1_sg U62989 ( .A(n53083), .B(n57230), .X(n33502) );
  nand_x1_sg U62990 ( .A(n50533), .B(n57230), .X(n33494) );
  nand_x1_sg U62991 ( .A(n53075), .B(n57230), .X(n33506) );
  nand_x1_sg U62992 ( .A(n53071), .B(n57230), .X(n33510) );
  nand_x1_sg U62993 ( .A(n53067), .B(n57230), .X(n33514) );
  nand_x1_sg U62994 ( .A(n53065), .B(n57230), .X(n33486) );
  nand_x1_sg U62995 ( .A(n53057), .B(n57230), .X(n33522) );
  nand_x1_sg U62996 ( .A(n53477), .B(n33570), .X(n33577) );
  nand_x1_sg U62997 ( .A(n53473), .B(n33570), .X(n33589) );
  nand_x1_sg U62998 ( .A(n50901), .B(n33570), .X(n33581) );
  nand_x1_sg U62999 ( .A(n53471), .B(n33570), .X(n33567) );
  nand_x1_sg U63000 ( .A(n53463), .B(n33570), .X(n33573) );
  nand_x1_sg U63001 ( .A(n53461), .B(n33570), .X(n33597) );
  nand_x1_sg U63002 ( .A(n53453), .B(n33570), .X(n33605) );
  nand_x1_sg U63003 ( .A(n53085), .B(n33485), .X(n33482) );
  nand_x1_sg U63004 ( .A(n53081), .B(n33485), .X(n33504) );
  nand_x1_sg U63005 ( .A(n53079), .B(n33485), .X(n33496) );
  nand_x1_sg U63006 ( .A(n53077), .B(n33485), .X(n33488) );
  nand_x1_sg U63007 ( .A(n53069), .B(n33485), .X(n33512) );
  nand_x1_sg U63008 ( .A(n53059), .B(n33485), .X(n33492) );
  nand_x1_sg U63009 ( .A(n50529), .B(n33485), .X(n33520) );
  nand_x1_sg U63010 ( .A(n53481), .B(n57224), .X(n33575) );
  nand_x1_sg U63011 ( .A(n53479), .B(n57224), .X(n33583) );
  nand_x1_sg U63012 ( .A(n50895), .B(n57224), .X(n33603) );
  nand_x1_sg U63013 ( .A(n53087), .B(n57230), .X(n33490) );
  nand_x1_sg U63014 ( .A(n50535), .B(n57230), .X(n33498) );
  nand_x1_sg U63015 ( .A(n50531), .B(n57230), .X(n33518) );
  nand_x1_sg U63016 ( .A(n50899), .B(n33570), .X(n33593) );
  nand_x1_sg U63017 ( .A(n53457), .B(n33570), .X(n33601) );
  nand_x1_sg U63018 ( .A(n53455), .B(n33570), .X(n33585) );
  nand_x1_sg U63019 ( .A(n53073), .B(n33485), .X(n33508) );
  nand_x1_sg U63020 ( .A(n53063), .B(n33485), .X(n33516) );
  nand_x1_sg U63021 ( .A(n53061), .B(n33485), .X(n33500) );
  nand_x1_sg U63022 ( .A(n47599), .B(n67532), .X(n26284) );
  nand_x1_sg U63023 ( .A(n26117), .B(n47399), .X(n26269) );
  nand_x1_sg U63024 ( .A(n26117), .B(n47397), .X(n26305) );
  nand_x2_sg U63025 ( .A(n26301), .B(n26302), .X(n26300) );
  nand_x1_sg U63026 ( .A(n47575), .B(n26122), .X(n26302) );
  nand_x1_sg U63027 ( .A(n53503), .B(n57213), .X(n33696) );
  nand_x1_sg U63028 ( .A(n50915), .B(n57213), .X(n33716) );
  nand_x1_sg U63029 ( .A(n50913), .B(n57212), .X(n33718) );
  nand_x1_sg U63030 ( .A(n53501), .B(n57213), .X(n33710) );
  nand_x1_sg U63031 ( .A(n50911), .B(n33699), .X(n33708) );
  nand_x1_sg U63032 ( .A(n53499), .B(n33699), .X(n33702) );
  nand_x1_sg U63033 ( .A(n50909), .B(n33699), .X(n33720) );
  nand_x1_sg U63034 ( .A(n50907), .B(n57212), .X(n33724) );
  nand_x1_sg U63035 ( .A(n53495), .B(n33699), .X(n33726) );
  nand_x1_sg U63036 ( .A(n50905), .B(n57213), .X(n33728) );
  nand_x1_sg U63037 ( .A(n53493), .B(n57212), .X(n33700) );
  nand_x1_sg U63038 ( .A(n53487), .B(n57212), .X(n33706) );
  nand_x1_sg U63039 ( .A(n53485), .B(n57213), .X(n33734) );
  nand_x1_sg U63040 ( .A(n53483), .B(n57212), .X(n33736) );
  nand_x1_sg U63041 ( .A(n53395), .B(n57257), .X(n33190) );
  nand_x1_sg U63042 ( .A(n53393), .B(n57258), .X(n33200) );
  nand_x1_sg U63043 ( .A(n50823), .B(n57257), .X(n33202) );
  nand_x1_sg U63044 ( .A(n53391), .B(n57258), .X(n33194) );
  nand_x1_sg U63045 ( .A(n50821), .B(n57258), .X(n33180) );
  nand_x1_sg U63046 ( .A(n53389), .B(n57257), .X(n33184) );
  nand_x1_sg U63047 ( .A(n50819), .B(n33183), .X(n33204) );
  nand_x1_sg U63048 ( .A(n50817), .B(n57257), .X(n33208) );
  nand_x1_sg U63049 ( .A(n53385), .B(n33183), .X(n33186) );
  nand_x1_sg U63050 ( .A(n50815), .B(n33183), .X(n33210) );
  nand_x1_sg U63051 ( .A(n53383), .B(n33183), .X(n33192) );
  nand_x1_sg U63052 ( .A(n53381), .B(n57258), .X(n33212) );
  nand_x1_sg U63053 ( .A(n53375), .B(n57258), .X(n33218) );
  nand_x1_sg U63054 ( .A(n53373), .B(n57257), .X(n33220) );
  nand_x1_sg U63055 ( .A(n50697), .B(n57238), .X(n33398) );
  nand_x1_sg U63056 ( .A(n50695), .B(n57238), .X(n33418) );
  nand_x1_sg U63057 ( .A(n53241), .B(n57237), .X(n33420) );
  nand_x1_sg U63058 ( .A(n53239), .B(n57238), .X(n33412) );
  nand_x1_sg U63059 ( .A(n50693), .B(n33401), .X(n33410) );
  nand_x1_sg U63060 ( .A(n50691), .B(n33401), .X(n33404) );
  nand_x1_sg U63061 ( .A(n50689), .B(n33401), .X(n33422) );
  nand_x1_sg U63062 ( .A(n50687), .B(n57237), .X(n33426) );
  nand_x1_sg U63063 ( .A(n50685), .B(n33401), .X(n33428) );
  nand_x1_sg U63064 ( .A(n50683), .B(n57238), .X(n33430) );
  nand_x1_sg U63065 ( .A(n53235), .B(n57237), .X(n33402) );
  nand_x1_sg U63066 ( .A(n50677), .B(n57237), .X(n33408) );
  nand_x1_sg U63067 ( .A(n53231), .B(n57238), .X(n33436) );
  nand_x1_sg U63068 ( .A(n53229), .B(n57237), .X(n33438) );
  nand_x1_sg U63069 ( .A(n53163), .B(n57250), .X(n33267) );
  nand_x1_sg U63070 ( .A(n50615), .B(n57250), .X(n33287) );
  nand_x1_sg U63071 ( .A(n50613), .B(n57249), .X(n33289) );
  nand_x1_sg U63072 ( .A(n53161), .B(n57250), .X(n33281) );
  nand_x1_sg U63073 ( .A(n50611), .B(n33270), .X(n33279) );
  nand_x1_sg U63074 ( .A(n53159), .B(n33270), .X(n33273) );
  nand_x1_sg U63075 ( .A(n50609), .B(n33270), .X(n33291) );
  nand_x1_sg U63076 ( .A(n50607), .B(n57249), .X(n33295) );
  nand_x1_sg U63077 ( .A(n53155), .B(n33270), .X(n33297) );
  nand_x1_sg U63078 ( .A(n50605), .B(n57250), .X(n33299) );
  nand_x1_sg U63079 ( .A(n53153), .B(n57249), .X(n33271) );
  nand_x1_sg U63080 ( .A(n53147), .B(n57249), .X(n33277) );
  nand_x1_sg U63081 ( .A(n53145), .B(n57250), .X(n33305) );
  nand_x1_sg U63082 ( .A(n53143), .B(n57249), .X(n33307) );
  nand_x1_sg U63083 ( .A(n50939), .B(n57217), .X(n33654) );
  nand_x1_sg U63084 ( .A(n50937), .B(n57217), .X(n33674) );
  nand_x1_sg U63085 ( .A(n50935), .B(n57216), .X(n33676) );
  nand_x1_sg U63086 ( .A(n53519), .B(n57217), .X(n33668) );
  nand_x1_sg U63087 ( .A(n50933), .B(n33657), .X(n33666) );
  nand_x1_sg U63088 ( .A(n50931), .B(n33657), .X(n33660) );
  nand_x1_sg U63089 ( .A(n50929), .B(n33657), .X(n33678) );
  nand_x1_sg U63090 ( .A(n50927), .B(n57216), .X(n33682) );
  nand_x1_sg U63091 ( .A(n50925), .B(n33657), .X(n33684) );
  nand_x1_sg U63092 ( .A(n50923), .B(n57217), .X(n33686) );
  nand_x1_sg U63093 ( .A(n53515), .B(n57216), .X(n33658) );
  nand_x1_sg U63094 ( .A(n53511), .B(n57216), .X(n33664) );
  nand_x1_sg U63095 ( .A(n53509), .B(n57217), .X(n33692) );
  nand_x1_sg U63096 ( .A(n53507), .B(n57216), .X(n33694) );
  nand_x1_sg U63097 ( .A(n53371), .B(n57254), .X(n33223) );
  nand_x1_sg U63098 ( .A(n53369), .B(n57254), .X(n33243) );
  nand_x1_sg U63099 ( .A(n50807), .B(n57253), .X(n33245) );
  nand_x1_sg U63100 ( .A(n53367), .B(n57254), .X(n33237) );
  nand_x1_sg U63101 ( .A(n50805), .B(n33226), .X(n33235) );
  nand_x1_sg U63102 ( .A(n53365), .B(n33226), .X(n33229) );
  nand_x1_sg U63103 ( .A(n50803), .B(n33226), .X(n33247) );
  nand_x1_sg U63104 ( .A(n50801), .B(n57253), .X(n33251) );
  nand_x1_sg U63105 ( .A(n53361), .B(n33226), .X(n33253) );
  nand_x1_sg U63106 ( .A(n50799), .B(n57254), .X(n33255) );
  nand_x1_sg U63107 ( .A(n53359), .B(n57253), .X(n33227) );
  nand_x1_sg U63108 ( .A(n53353), .B(n57253), .X(n33233) );
  nand_x1_sg U63109 ( .A(n53351), .B(n57254), .X(n33261) );
  nand_x1_sg U63110 ( .A(n53349), .B(n57253), .X(n33263) );
  nand_x1_sg U63111 ( .A(n52935), .B(n57194), .X(n33923) );
  nand_x1_sg U63112 ( .A(n50443), .B(n57195), .X(n33933) );
  nand_x1_sg U63113 ( .A(n52933), .B(n57194), .X(n33935) );
  nand_x1_sg U63114 ( .A(n52931), .B(n57195), .X(n33927) );
  nand_x1_sg U63115 ( .A(n50441), .B(n57195), .X(n33913) );
  nand_x1_sg U63116 ( .A(n52929), .B(n57194), .X(n33917) );
  nand_x1_sg U63117 ( .A(n50439), .B(n33916), .X(n33937) );
  nand_x1_sg U63118 ( .A(n50437), .B(n57194), .X(n33941) );
  nand_x1_sg U63119 ( .A(n52925), .B(n33916), .X(n33919) );
  nand_x1_sg U63120 ( .A(n50435), .B(n33916), .X(n33943) );
  nand_x1_sg U63121 ( .A(n52923), .B(n33916), .X(n33925) );
  nand_x1_sg U63122 ( .A(n52921), .B(n57195), .X(n33945) );
  nand_x1_sg U63123 ( .A(n52915), .B(n57195), .X(n33951) );
  nand_x1_sg U63124 ( .A(n52913), .B(n57194), .X(n33953) );
  nand_x1_sg U63125 ( .A(n50427), .B(n57190), .X(n33966) );
  nand_x1_sg U63126 ( .A(n50425), .B(n57191), .X(n33976) );
  nand_x1_sg U63127 ( .A(n50423), .B(n57190), .X(n33978) );
  nand_x1_sg U63128 ( .A(n52911), .B(n57191), .X(n33970) );
  nand_x1_sg U63129 ( .A(n50421), .B(n57191), .X(n33956) );
  nand_x1_sg U63130 ( .A(n50419), .B(n57190), .X(n33960) );
  nand_x1_sg U63131 ( .A(n50417), .B(n33959), .X(n33980) );
  nand_x1_sg U63132 ( .A(n50413), .B(n57190), .X(n33984) );
  nand_x1_sg U63133 ( .A(n50411), .B(n33959), .X(n33962) );
  nand_x1_sg U63134 ( .A(n50409), .B(n33959), .X(n33986) );
  nand_x1_sg U63135 ( .A(n50407), .B(n33959), .X(n33968) );
  nand_x1_sg U63136 ( .A(n52909), .B(n57191), .X(n33988) );
  nand_x1_sg U63137 ( .A(n52907), .B(n57191), .X(n33994) );
  nand_x1_sg U63138 ( .A(n52905), .B(n57190), .X(n33996) );
  nand_x1_sg U63139 ( .A(n50903), .B(n33699), .X(n33732) );
  nand_x1_sg U63140 ( .A(n53489), .B(n33699), .X(n33714) );
  nand_x1_sg U63141 ( .A(n53379), .B(n33183), .X(n33198) );
  nand_x1_sg U63142 ( .A(n53377), .B(n33183), .X(n33216) );
  nand_x1_sg U63143 ( .A(n50681), .B(n33401), .X(n33434) );
  nand_x1_sg U63144 ( .A(n50679), .B(n33401), .X(n33416) );
  nand_x1_sg U63145 ( .A(n50603), .B(n33270), .X(n33303) );
  nand_x1_sg U63146 ( .A(n53149), .B(n33270), .X(n33285) );
  nand_x1_sg U63147 ( .A(n50917), .B(n57213), .X(n33704) );
  nand_x1_sg U63148 ( .A(n53505), .B(n57212), .X(n33712) );
  nand_x1_sg U63149 ( .A(n53497), .B(n57213), .X(n33722) );
  nand_x1_sg U63150 ( .A(n53491), .B(n57212), .X(n33730) );
  nand_x1_sg U63151 ( .A(n50827), .B(n57258), .X(n33188) );
  nand_x1_sg U63152 ( .A(n50825), .B(n57257), .X(n33196) );
  nand_x1_sg U63153 ( .A(n53387), .B(n57258), .X(n33206) );
  nand_x1_sg U63154 ( .A(n50813), .B(n57257), .X(n33214) );
  nand_x1_sg U63155 ( .A(n53243), .B(n57238), .X(n33406) );
  nand_x1_sg U63156 ( .A(n50699), .B(n57237), .X(n33414) );
  nand_x1_sg U63157 ( .A(n53237), .B(n57238), .X(n33424) );
  nand_x1_sg U63158 ( .A(n53233), .B(n57237), .X(n33432) );
  nand_x1_sg U63159 ( .A(n50617), .B(n57250), .X(n33275) );
  nand_x1_sg U63160 ( .A(n53165), .B(n57249), .X(n33283) );
  nand_x1_sg U63161 ( .A(n53157), .B(n57250), .X(n33293) );
  nand_x1_sg U63162 ( .A(n53151), .B(n57249), .X(n33301) );
  nand_x1_sg U63163 ( .A(n50943), .B(n57217), .X(n33662) );
  nand_x1_sg U63164 ( .A(n50941), .B(n57216), .X(n33670) );
  nand_x1_sg U63165 ( .A(n53517), .B(n57217), .X(n33680) );
  nand_x1_sg U63166 ( .A(n53513), .B(n57216), .X(n33688) );
  nand_x1_sg U63167 ( .A(n50921), .B(n33657), .X(n33690) );
  nand_x1_sg U63168 ( .A(n50919), .B(n33657), .X(n33672) );
  nand_x1_sg U63169 ( .A(n50811), .B(n57254), .X(n33231) );
  nand_x1_sg U63170 ( .A(n50809), .B(n57253), .X(n33239) );
  nand_x1_sg U63171 ( .A(n53363), .B(n57254), .X(n33249) );
  nand_x1_sg U63172 ( .A(n53357), .B(n57253), .X(n33257) );
  nand_x1_sg U63173 ( .A(n50797), .B(n33226), .X(n33259) );
  nand_x1_sg U63174 ( .A(n53355), .B(n33226), .X(n33241) );
  nand_x1_sg U63175 ( .A(n50447), .B(n57195), .X(n33921) );
  nand_x1_sg U63176 ( .A(n50445), .B(n57194), .X(n33929) );
  nand_x1_sg U63177 ( .A(n52927), .B(n57195), .X(n33939) );
  nand_x1_sg U63178 ( .A(n50433), .B(n57194), .X(n33947) );
  nand_x1_sg U63179 ( .A(n52919), .B(n33916), .X(n33931) );
  nand_x1_sg U63180 ( .A(n52917), .B(n33916), .X(n33949) );
  nand_x1_sg U63181 ( .A(n50431), .B(n57191), .X(n33964) );
  nand_x1_sg U63182 ( .A(n50429), .B(n57190), .X(n33972) );
  nand_x1_sg U63183 ( .A(n50415), .B(n57191), .X(n33982) );
  nand_x1_sg U63184 ( .A(n50405), .B(n57190), .X(n33990) );
  nand_x1_sg U63185 ( .A(n50403), .B(n33959), .X(n33974) );
  nand_x1_sg U63186 ( .A(n50401), .B(n33959), .X(n33992) );
  nand_x2_sg U63187 ( .A(n47615), .B(n57955), .X(n57956) );
  nor_x1_sg U63188 ( .A(n57380), .B(n58755), .X(n58756) );
  nor_x1_sg U63189 ( .A(n57372), .B(n58750), .X(n58751) );
  nor_x1_sg U63190 ( .A(n57381), .B(n58745), .X(n58746) );
  nor_x1_sg U63191 ( .A(n57371), .B(n58740), .X(n58741) );
  nor_x1_sg U63192 ( .A(n57378), .B(n58735), .X(n58736) );
  nor_x1_sg U63193 ( .A(n57379), .B(n58730), .X(n58731) );
  nor_x1_sg U63194 ( .A(n57377), .B(n58725), .X(n58726) );
  nor_x1_sg U63195 ( .A(n57367), .B(n58720), .X(n58721) );
  nor_x1_sg U63196 ( .A(n57368), .B(n58715), .X(n58716) );
  nor_x1_sg U63197 ( .A(n57365), .B(n58710), .X(n58711) );
  nor_x1_sg U63198 ( .A(n57381), .B(n58705), .X(n58706) );
  nor_x1_sg U63199 ( .A(n57381), .B(n58700), .X(n58701) );
  nor_x1_sg U63200 ( .A(n57381), .B(n58695), .X(n58696) );
  nor_x1_sg U63201 ( .A(n57381), .B(n58690), .X(n58691) );
  nor_x1_sg U63202 ( .A(n57381), .B(n58685), .X(n58686) );
  nor_x1_sg U63203 ( .A(n57381), .B(n58680), .X(n58681) );
  nor_x1_sg U63204 ( .A(n57381), .B(n58675), .X(n58676) );
  nor_x1_sg U63205 ( .A(n57381), .B(n58670), .X(n58671) );
  nor_x1_sg U63206 ( .A(n57381), .B(n58665), .X(n58666) );
  nor_x1_sg U63207 ( .A(n57372), .B(n61855), .X(n61857) );
  nor_x1_sg U63208 ( .A(n57381), .B(n61850), .X(n61851) );
  nor_x1_sg U63209 ( .A(n57372), .B(n61845), .X(n61846) );
  nor_x1_sg U63210 ( .A(n57371), .B(n61840), .X(n61841) );
  nor_x1_sg U63211 ( .A(n57381), .B(n61835), .X(n61836) );
  nor_x1_sg U63212 ( .A(n57371), .B(n61830), .X(n61831) );
  nor_x1_sg U63213 ( .A(n57372), .B(n61825), .X(n61826) );
  nor_x1_sg U63214 ( .A(n57381), .B(n61820), .X(n61821) );
  nor_x1_sg U63215 ( .A(n57381), .B(n61815), .X(n61816) );
  nor_x1_sg U63216 ( .A(n57372), .B(n61810), .X(n61811) );
  nor_x1_sg U63217 ( .A(n57381), .B(n61805), .X(n61806) );
  nor_x1_sg U63218 ( .A(n57371), .B(n61800), .X(n61801) );
  nor_x1_sg U63219 ( .A(n57372), .B(n61795), .X(n61796) );
  nor_x1_sg U63220 ( .A(n57381), .B(n61790), .X(n61791) );
  nor_x1_sg U63221 ( .A(n57358), .B(n61785), .X(n61786) );
  nor_x1_sg U63222 ( .A(n57371), .B(n61780), .X(n61781) );
  nor_x1_sg U63223 ( .A(n57371), .B(n61775), .X(n61776) );
  nor_x1_sg U63224 ( .A(n57372), .B(n61770), .X(n61771) );
  nor_x1_sg U63225 ( .A(n57371), .B(n61765), .X(n61766) );
  nor_x1_sg U63226 ( .A(n57372), .B(n61760), .X(n61761) );
  nor_x1_sg U63227 ( .A(n57381), .B(n61755), .X(n61756) );
  nor_x1_sg U63228 ( .A(n57371), .B(n61750), .X(n61751) );
  nor_x1_sg U63229 ( .A(n57372), .B(n61745), .X(n61746) );
  nor_x1_sg U63230 ( .A(n57381), .B(n61740), .X(n61741) );
  nor_x1_sg U63231 ( .A(n57387), .B(n61735), .X(n61736) );
  nor_x1_sg U63232 ( .A(n57372), .B(n61730), .X(n61731) );
  nor_x1_sg U63233 ( .A(n57381), .B(n61725), .X(n61726) );
  nor_x1_sg U63234 ( .A(n57372), .B(n61720), .X(n61721) );
  nor_x1_sg U63235 ( .A(n57371), .B(n61715), .X(n61716) );
  nor_x1_sg U63236 ( .A(n57372), .B(n61710), .X(n61711) );
  nor_x1_sg U63237 ( .A(n57381), .B(n61705), .X(n61706) );
  nor_x1_sg U63238 ( .A(n57371), .B(n61700), .X(n61701) );
  nor_x1_sg U63239 ( .A(n57371), .B(n61695), .X(n61696) );
  nor_x1_sg U63240 ( .A(n57372), .B(n61690), .X(n61691) );
  nor_x1_sg U63241 ( .A(n57381), .B(n61685), .X(n61686) );
  nor_x1_sg U63242 ( .A(n57366), .B(n61680), .X(n61681) );
  nor_x1_sg U63243 ( .A(n57350), .B(n61675), .X(n61676) );
  nor_x1_sg U63244 ( .A(n57350), .B(n61670), .X(n61671) );
  nor_x1_sg U63245 ( .A(n57350), .B(n61665), .X(n61666) );
  nor_x1_sg U63246 ( .A(n57350), .B(n61660), .X(n61661) );
  nor_x1_sg U63247 ( .A(n57350), .B(n61655), .X(n61656) );
  nor_x1_sg U63248 ( .A(n57350), .B(n61650), .X(n61651) );
  nor_x1_sg U63249 ( .A(n57350), .B(n61645), .X(n61646) );
  nor_x1_sg U63250 ( .A(n57350), .B(n61640), .X(n61641) );
  nor_x1_sg U63251 ( .A(n57350), .B(n61635), .X(n61636) );
  nor_x1_sg U63252 ( .A(n57351), .B(n61630), .X(n61631) );
  nor_x1_sg U63253 ( .A(n57351), .B(n61625), .X(n61626) );
  nor_x1_sg U63254 ( .A(n57351), .B(n61620), .X(n61621) );
  nor_x1_sg U63255 ( .A(n57351), .B(n61615), .X(n61616) );
  nor_x1_sg U63256 ( .A(n57351), .B(n61610), .X(n61611) );
  nor_x1_sg U63257 ( .A(n57351), .B(n61605), .X(n61606) );
  nor_x1_sg U63258 ( .A(n57351), .B(n61600), .X(n61601) );
  nor_x1_sg U63259 ( .A(n57351), .B(n61595), .X(n61596) );
  nor_x1_sg U63260 ( .A(n57351), .B(n61590), .X(n61591) );
  nor_x1_sg U63261 ( .A(n57388), .B(n61585), .X(n61586) );
  nor_x1_sg U63262 ( .A(n57352), .B(n61580), .X(n61581) );
  nor_x1_sg U63263 ( .A(n57368), .B(n61575), .X(n61576) );
  nor_x1_sg U63264 ( .A(n57365), .B(n61570), .X(n61571) );
  nor_x1_sg U63265 ( .A(n57359), .B(n61565), .X(n61566) );
  nor_x1_sg U63266 ( .A(n57360), .B(n61560), .X(n61561) );
  nor_x1_sg U63267 ( .A(n57357), .B(n61555), .X(n61556) );
  nor_x1_sg U63268 ( .A(n57358), .B(n61550), .X(n61551) );
  nor_x1_sg U63269 ( .A(n57350), .B(n61545), .X(n61546) );
  nor_x1_sg U63270 ( .A(n57352), .B(n61540), .X(n61541) );
  nor_x1_sg U63271 ( .A(n57352), .B(n61535), .X(n61536) );
  nor_x1_sg U63272 ( .A(n57352), .B(n61530), .X(n61531) );
  nor_x1_sg U63273 ( .A(n57352), .B(n61525), .X(n61526) );
  nor_x1_sg U63274 ( .A(n57352), .B(n61520), .X(n61521) );
  nor_x1_sg U63275 ( .A(n57352), .B(n61515), .X(n61516) );
  nor_x1_sg U63276 ( .A(n57352), .B(n61510), .X(n61511) );
  nor_x1_sg U63277 ( .A(n57352), .B(n61505), .X(n61506) );
  nor_x1_sg U63278 ( .A(n57352), .B(n61500), .X(n61501) );
  nor_x1_sg U63279 ( .A(n57353), .B(n61495), .X(n61496) );
  nor_x1_sg U63280 ( .A(n57353), .B(n61490), .X(n61491) );
  nor_x1_sg U63281 ( .A(n57353), .B(n61485), .X(n61486) );
  nor_x1_sg U63282 ( .A(n57353), .B(n61480), .X(n61481) );
  nor_x1_sg U63283 ( .A(n57353), .B(n61475), .X(n61476) );
  nor_x1_sg U63284 ( .A(n57353), .B(n61470), .X(n61471) );
  nor_x1_sg U63285 ( .A(n57353), .B(n61465), .X(n61466) );
  nor_x1_sg U63286 ( .A(n57353), .B(n61460), .X(n61461) );
  nor_x1_sg U63287 ( .A(n57353), .B(n61455), .X(n61456) );
  nor_x1_sg U63288 ( .A(n57354), .B(n61450), .X(n61451) );
  nor_x1_sg U63289 ( .A(n57354), .B(n61445), .X(n61446) );
  nor_x1_sg U63290 ( .A(n57354), .B(n61440), .X(n61441) );
  nor_x1_sg U63291 ( .A(n57354), .B(n61435), .X(n61436) );
  nor_x1_sg U63292 ( .A(n57354), .B(n61430), .X(n61431) );
  nor_x1_sg U63293 ( .A(n57354), .B(n61425), .X(n61426) );
  nor_x1_sg U63294 ( .A(n57354), .B(n61420), .X(n61421) );
  nor_x1_sg U63295 ( .A(n57354), .B(n61415), .X(n61416) );
  nor_x1_sg U63296 ( .A(n57354), .B(n61410), .X(n61411) );
  nor_x1_sg U63297 ( .A(n57355), .B(n61405), .X(n61406) );
  nor_x1_sg U63298 ( .A(n57355), .B(n61400), .X(n61401) );
  nor_x1_sg U63299 ( .A(n57355), .B(n61395), .X(n61396) );
  nor_x1_sg U63300 ( .A(n57355), .B(n61390), .X(n61391) );
  nor_x1_sg U63301 ( .A(n57355), .B(n61385), .X(n61386) );
  nor_x1_sg U63302 ( .A(n57355), .B(n61380), .X(n61381) );
  nor_x1_sg U63303 ( .A(n57355), .B(n61375), .X(n61376) );
  nor_x1_sg U63304 ( .A(n57355), .B(n61370), .X(n61371) );
  nor_x1_sg U63305 ( .A(n57355), .B(n61365), .X(n61366) );
  nor_x1_sg U63306 ( .A(n57356), .B(n61360), .X(n61361) );
  nor_x1_sg U63307 ( .A(n57356), .B(n61355), .X(n61356) );
  nor_x1_sg U63308 ( .A(n57356), .B(n61350), .X(n61351) );
  nor_x1_sg U63309 ( .A(n57356), .B(n61345), .X(n61346) );
  nor_x1_sg U63310 ( .A(n57356), .B(n61340), .X(n61341) );
  nor_x1_sg U63311 ( .A(n57356), .B(n61335), .X(n61336) );
  nor_x1_sg U63312 ( .A(n57356), .B(n61330), .X(n61331) );
  nor_x1_sg U63313 ( .A(n57356), .B(n61325), .X(n61326) );
  nor_x1_sg U63314 ( .A(n57356), .B(n61320), .X(n61321) );
  nor_x1_sg U63315 ( .A(n57357), .B(n61315), .X(n61316) );
  nor_x1_sg U63316 ( .A(n57357), .B(n61310), .X(n61311) );
  nor_x1_sg U63317 ( .A(n57357), .B(n61305), .X(n61306) );
  nor_x1_sg U63318 ( .A(n57357), .B(n61300), .X(n61301) );
  nor_x1_sg U63319 ( .A(n57357), .B(n61295), .X(n61296) );
  nor_x1_sg U63320 ( .A(n57357), .B(n61290), .X(n61291) );
  nor_x1_sg U63321 ( .A(n57357), .B(n61285), .X(n61286) );
  nor_x1_sg U63322 ( .A(n57357), .B(n61280), .X(n61281) );
  nor_x1_sg U63323 ( .A(n57357), .B(n61275), .X(n61276) );
  nor_x1_sg U63324 ( .A(n57358), .B(n61270), .X(n61271) );
  nor_x1_sg U63325 ( .A(n57358), .B(n61265), .X(n61266) );
  nor_x1_sg U63326 ( .A(n57358), .B(n61260), .X(n61261) );
  nor_x1_sg U63327 ( .A(n57358), .B(n61255), .X(n61256) );
  nor_x1_sg U63328 ( .A(n57358), .B(n61250), .X(n61251) );
  nor_x1_sg U63329 ( .A(n57358), .B(n61245), .X(n61246) );
  nor_x1_sg U63330 ( .A(n57358), .B(n61240), .X(n61241) );
  nor_x1_sg U63331 ( .A(n57358), .B(n61235), .X(n61236) );
  nor_x1_sg U63332 ( .A(n57358), .B(n61230), .X(n61231) );
  nor_x1_sg U63333 ( .A(n57359), .B(n61225), .X(n61226) );
  nor_x1_sg U63334 ( .A(n57359), .B(n61220), .X(n61221) );
  nor_x1_sg U63335 ( .A(n57359), .B(n61215), .X(n61216) );
  nor_x1_sg U63336 ( .A(n57359), .B(n61210), .X(n61211) );
  nor_x1_sg U63337 ( .A(n57359), .B(n61205), .X(n61206) );
  nor_x1_sg U63338 ( .A(n57359), .B(n61200), .X(n61201) );
  nor_x1_sg U63339 ( .A(n57359), .B(n61195), .X(n61196) );
  nor_x1_sg U63340 ( .A(n57359), .B(n61190), .X(n61191) );
  nor_x1_sg U63341 ( .A(n57359), .B(n61185), .X(n61186) );
  nor_x1_sg U63342 ( .A(n57360), .B(n61180), .X(n61181) );
  nor_x1_sg U63343 ( .A(n57360), .B(n61175), .X(n61176) );
  nor_x1_sg U63344 ( .A(n57360), .B(n61170), .X(n61171) );
  nor_x1_sg U63345 ( .A(n57360), .B(n61165), .X(n61166) );
  nor_x1_sg U63346 ( .A(n57360), .B(n61160), .X(n61161) );
  nor_x1_sg U63347 ( .A(n57360), .B(n61155), .X(n61156) );
  nor_x1_sg U63348 ( .A(n57360), .B(n61150), .X(n61151) );
  nor_x1_sg U63349 ( .A(n57360), .B(n61145), .X(n61146) );
  nor_x1_sg U63350 ( .A(n57360), .B(n61140), .X(n61141) );
  nor_x1_sg U63351 ( .A(n57361), .B(n61135), .X(n61136) );
  nor_x1_sg U63352 ( .A(n57361), .B(n61130), .X(n61131) );
  nor_x1_sg U63353 ( .A(n57361), .B(n61125), .X(n61126) );
  nor_x1_sg U63354 ( .A(n57361), .B(n61120), .X(n61121) );
  nor_x1_sg U63355 ( .A(n57361), .B(n61115), .X(n61116) );
  nor_x1_sg U63356 ( .A(n57361), .B(n61110), .X(n61111) );
  nor_x1_sg U63357 ( .A(n57361), .B(n61105), .X(n61106) );
  nor_x1_sg U63358 ( .A(n57361), .B(n61100), .X(n61101) );
  nor_x1_sg U63359 ( .A(n57361), .B(n61095), .X(n61096) );
  nor_x1_sg U63360 ( .A(n57362), .B(n61090), .X(n61091) );
  nor_x1_sg U63361 ( .A(n57362), .B(n61085), .X(n61086) );
  nor_x1_sg U63362 ( .A(n57362), .B(n61080), .X(n61081) );
  nor_x1_sg U63363 ( .A(n57362), .B(n61075), .X(n61076) );
  nor_x1_sg U63364 ( .A(n57362), .B(n61070), .X(n61071) );
  nor_x1_sg U63365 ( .A(n57362), .B(n61065), .X(n61066) );
  nor_x1_sg U63366 ( .A(n57362), .B(n61060), .X(n61061) );
  nor_x1_sg U63367 ( .A(n57362), .B(n61055), .X(n61056) );
  nor_x1_sg U63368 ( .A(n57362), .B(n61050), .X(n61051) );
  nor_x1_sg U63369 ( .A(n57363), .B(n61045), .X(n61046) );
  nor_x1_sg U63370 ( .A(n57363), .B(n61040), .X(n61041) );
  nor_x1_sg U63371 ( .A(n57363), .B(n61035), .X(n61036) );
  nor_x1_sg U63372 ( .A(n57363), .B(n61030), .X(n61031) );
  nor_x1_sg U63373 ( .A(n57363), .B(n61025), .X(n61026) );
  nor_x1_sg U63374 ( .A(n57363), .B(n61020), .X(n61021) );
  nor_x1_sg U63375 ( .A(n57363), .B(n61015), .X(n61016) );
  nor_x1_sg U63376 ( .A(n57363), .B(n61010), .X(n61011) );
  nor_x1_sg U63377 ( .A(n57363), .B(n61005), .X(n61006) );
  nor_x1_sg U63378 ( .A(n57364), .B(n61000), .X(n61001) );
  nor_x1_sg U63379 ( .A(n57364), .B(n60995), .X(n60996) );
  nor_x1_sg U63380 ( .A(n57364), .B(n60990), .X(n60991) );
  nor_x1_sg U63381 ( .A(n57364), .B(n60985), .X(n60986) );
  nor_x1_sg U63382 ( .A(n57364), .B(n60980), .X(n60981) );
  nor_x1_sg U63383 ( .A(n57364), .B(n60975), .X(n60976) );
  nor_x1_sg U63384 ( .A(n57364), .B(n60970), .X(n60971) );
  nor_x1_sg U63385 ( .A(n57364), .B(n60965), .X(n60966) );
  nor_x1_sg U63386 ( .A(n57364), .B(n60960), .X(n60961) );
  nor_x1_sg U63387 ( .A(n57365), .B(n60955), .X(n60956) );
  nor_x1_sg U63388 ( .A(n57365), .B(n60950), .X(n60951) );
  nor_x1_sg U63389 ( .A(n57365), .B(n60945), .X(n60946) );
  nor_x1_sg U63390 ( .A(n57365), .B(n60940), .X(n60941) );
  nor_x1_sg U63391 ( .A(n57365), .B(n60935), .X(n60936) );
  nor_x1_sg U63392 ( .A(n57365), .B(n60930), .X(n60931) );
  nor_x1_sg U63393 ( .A(n57365), .B(n60925), .X(n60926) );
  nor_x1_sg U63394 ( .A(n57365), .B(n60920), .X(n60921) );
  nor_x1_sg U63395 ( .A(n57365), .B(n60915), .X(n60916) );
  nor_x1_sg U63396 ( .A(n57366), .B(n60910), .X(n60911) );
  nor_x1_sg U63397 ( .A(n57366), .B(n60905), .X(n60906) );
  nor_x1_sg U63398 ( .A(n57366), .B(n60900), .X(n60901) );
  nor_x1_sg U63399 ( .A(n57366), .B(n60895), .X(n60896) );
  nor_x1_sg U63400 ( .A(n57366), .B(n60890), .X(n60891) );
  nor_x1_sg U63401 ( .A(n57366), .B(n60885), .X(n60886) );
  nor_x1_sg U63402 ( .A(n57366), .B(n60880), .X(n60881) );
  nor_x1_sg U63403 ( .A(n57366), .B(n60875), .X(n60876) );
  nor_x1_sg U63404 ( .A(n57366), .B(n60870), .X(n60871) );
  nor_x1_sg U63405 ( .A(n57367), .B(n60865), .X(n60866) );
  nor_x1_sg U63406 ( .A(n57367), .B(n60860), .X(n60861) );
  nor_x1_sg U63407 ( .A(n57367), .B(n60855), .X(n60856) );
  nor_x1_sg U63408 ( .A(n57367), .B(n60850), .X(n60851) );
  nor_x1_sg U63409 ( .A(n57367), .B(n60845), .X(n60846) );
  nor_x1_sg U63410 ( .A(n57367), .B(n60840), .X(n60841) );
  nor_x1_sg U63411 ( .A(n57367), .B(n60835), .X(n60836) );
  nor_x1_sg U63412 ( .A(n57367), .B(n60830), .X(n60831) );
  nor_x1_sg U63413 ( .A(n57367), .B(n60825), .X(n60826) );
  nor_x1_sg U63414 ( .A(n57368), .B(n60820), .X(n60821) );
  nor_x1_sg U63415 ( .A(n57368), .B(n60815), .X(n60816) );
  nor_x1_sg U63416 ( .A(n57368), .B(n60810), .X(n60811) );
  nor_x1_sg U63417 ( .A(n57368), .B(n60805), .X(n60806) );
  nor_x1_sg U63418 ( .A(n57368), .B(n60800), .X(n60801) );
  nor_x1_sg U63419 ( .A(n57368), .B(n60795), .X(n60796) );
  nor_x1_sg U63420 ( .A(n57368), .B(n60790), .X(n60791) );
  nor_x1_sg U63421 ( .A(n57368), .B(n60785), .X(n60786) );
  nor_x1_sg U63422 ( .A(n57368), .B(n60780), .X(n60781) );
  nor_x1_sg U63423 ( .A(n57390), .B(n60775), .X(n60776) );
  nor_x1_sg U63424 ( .A(n57387), .B(n60770), .X(n60771) );
  nor_x1_sg U63425 ( .A(n57388), .B(n60765), .X(n60766) );
  nor_x1_sg U63426 ( .A(n57359), .B(n60760), .X(n60761) );
  nor_x1_sg U63427 ( .A(n57360), .B(n60755), .X(n60756) );
  nor_x1_sg U63428 ( .A(n57357), .B(n60750), .X(n60751) );
  nor_x1_sg U63429 ( .A(n57358), .B(n60745), .X(n60746) );
  nor_x1_sg U63430 ( .A(n57367), .B(n60740), .X(n60741) );
  nor_x1_sg U63431 ( .A(n57368), .B(n60735), .X(n60736) );
  nor_x1_sg U63432 ( .A(n57387), .B(n60730), .X(n60731) );
  nor_x1_sg U63433 ( .A(n57387), .B(n60725), .X(n60726) );
  nor_x1_sg U63434 ( .A(n57388), .B(n60720), .X(n60721) );
  nor_x1_sg U63435 ( .A(n57376), .B(n60715), .X(n60716) );
  nor_x1_sg U63436 ( .A(n57359), .B(n60710), .X(n60711) );
  nor_x1_sg U63437 ( .A(n57390), .B(n60705), .X(n60706) );
  nor_x1_sg U63438 ( .A(n57378), .B(n60700), .X(n60701) );
  nor_x1_sg U63439 ( .A(n57387), .B(n60695), .X(n60696) );
  nor_x1_sg U63440 ( .A(n57377), .B(n60690), .X(n60691) );
  nor_x1_sg U63441 ( .A(n57376), .B(n60685), .X(n60686) );
  nor_x1_sg U63442 ( .A(n57365), .B(n60680), .X(n60681) );
  nor_x1_sg U63443 ( .A(n57373), .B(n60675), .X(n60676) );
  nor_x1_sg U63444 ( .A(n57351), .B(n60670), .X(n60671) );
  nor_x1_sg U63445 ( .A(n57387), .B(n60665), .X(n60666) );
  nor_x1_sg U63446 ( .A(n61856), .B(n60660), .X(n60661) );
  nor_x1_sg U63447 ( .A(n57388), .B(n60655), .X(n60656) );
  nor_x1_sg U63448 ( .A(n57373), .B(n60650), .X(n60651) );
  nor_x1_sg U63449 ( .A(n57374), .B(n60645), .X(n60646) );
  nor_x1_sg U63450 ( .A(n57374), .B(n60640), .X(n60641) );
  nor_x1_sg U63451 ( .A(n57366), .B(n60635), .X(n60636) );
  nor_x1_sg U63452 ( .A(n57365), .B(n60630), .X(n60631) );
  nor_x1_sg U63453 ( .A(n57366), .B(n60625), .X(n60626) );
  nor_x1_sg U63454 ( .A(n57387), .B(n60620), .X(n60621) );
  nor_x1_sg U63455 ( .A(n57387), .B(n60615), .X(n60616) );
  nor_x1_sg U63456 ( .A(n57388), .B(n60610), .X(n60611) );
  nor_x1_sg U63457 ( .A(n57378), .B(n60605), .X(n60606) );
  nor_x1_sg U63458 ( .A(n57379), .B(n60600), .X(n60601) );
  nor_x1_sg U63459 ( .A(n61856), .B(n60595), .X(n60596) );
  nor_x1_sg U63460 ( .A(n57387), .B(n60590), .X(n60591) );
  nor_x1_sg U63461 ( .A(n57376), .B(n60585), .X(n60586) );
  nor_x1_sg U63462 ( .A(n57367), .B(n60580), .X(n60581) );
  nor_x1_sg U63463 ( .A(n57375), .B(n60575), .X(n60576) );
  nor_x1_sg U63464 ( .A(n57350), .B(n60570), .X(n60571) );
  nor_x1_sg U63465 ( .A(n57366), .B(n60565), .X(n60566) );
  nor_x1_sg U63466 ( .A(n57373), .B(n60560), .X(n60561) );
  nor_x1_sg U63467 ( .A(n57359), .B(n60555), .X(n60556) );
  nor_x1_sg U63468 ( .A(n57374), .B(n60550), .X(n60551) );
  nor_x1_sg U63469 ( .A(n57376), .B(n60545), .X(n60546) );
  nor_x1_sg U63470 ( .A(n57365), .B(n60540), .X(n60541) );
  nor_x1_sg U63471 ( .A(n57381), .B(n60535), .X(n60536) );
  nor_x1_sg U63472 ( .A(n57357), .B(n60530), .X(n60531) );
  nor_x1_sg U63473 ( .A(n57360), .B(n60525), .X(n60526) );
  nor_x1_sg U63474 ( .A(n57388), .B(n60520), .X(n60521) );
  nor_x1_sg U63475 ( .A(n61856), .B(n60515), .X(n60516) );
  nor_x1_sg U63476 ( .A(n57351), .B(n60510), .X(n60511) );
  nor_x1_sg U63477 ( .A(n57390), .B(n60505), .X(n60506) );
  nor_x1_sg U63478 ( .A(n57390), .B(n60500), .X(n60501) );
  nor_x1_sg U63479 ( .A(n57388), .B(n60495), .X(n60496) );
  nor_x1_sg U63480 ( .A(n57390), .B(n60490), .X(n60491) );
  nor_x1_sg U63481 ( .A(n57388), .B(n60485), .X(n60486) );
  nor_x1_sg U63482 ( .A(n57390), .B(n60480), .X(n60481) );
  nor_x1_sg U63483 ( .A(n57387), .B(n60475), .X(n60476) );
  nor_x1_sg U63484 ( .A(n57388), .B(n60470), .X(n60471) );
  nor_x1_sg U63485 ( .A(n57390), .B(n60465), .X(n60466) );
  nor_x1_sg U63486 ( .A(n61856), .B(n60460), .X(n60461) );
  nor_x1_sg U63487 ( .A(n61856), .B(n60455), .X(n60456) );
  nor_x1_sg U63488 ( .A(n57390), .B(n60450), .X(n60451) );
  nor_x1_sg U63489 ( .A(n57376), .B(n60445), .X(n60446) );
  nor_x1_sg U63490 ( .A(n57376), .B(n60440), .X(n60441) );
  nor_x1_sg U63491 ( .A(n57375), .B(n60435), .X(n60436) );
  nor_x1_sg U63492 ( .A(n57352), .B(n60430), .X(n60431) );
  nor_x1_sg U63493 ( .A(n57387), .B(n60425), .X(n60426) );
  nor_x1_sg U63494 ( .A(n61856), .B(n60420), .X(n60421) );
  nor_x1_sg U63495 ( .A(n57374), .B(n60415), .X(n60416) );
  nor_x1_sg U63496 ( .A(n57352), .B(n60410), .X(n60411) );
  nor_x1_sg U63497 ( .A(n57373), .B(n60405), .X(n60406) );
  nor_x1_sg U63498 ( .A(n57377), .B(n60400), .X(n60401) );
  nor_x1_sg U63499 ( .A(n57358), .B(n60395), .X(n60396) );
  nor_x1_sg U63500 ( .A(n57359), .B(n60390), .X(n60391) );
  nor_x1_sg U63501 ( .A(n57360), .B(n60385), .X(n60386) );
  nor_x1_sg U63502 ( .A(n57357), .B(n60380), .X(n60381) );
  nor_x1_sg U63503 ( .A(n57358), .B(n60375), .X(n60376) );
  nor_x1_sg U63504 ( .A(n57352), .B(n60370), .X(n60371) );
  nor_x1_sg U63505 ( .A(n57360), .B(n60365), .X(n60366) );
  nor_x1_sg U63506 ( .A(n57359), .B(n60360), .X(n60361) );
  nor_x1_sg U63507 ( .A(n57367), .B(n60355), .X(n60356) );
  nor_x1_sg U63508 ( .A(n57368), .B(n60350), .X(n60351) );
  nor_x1_sg U63509 ( .A(n57365), .B(n60345), .X(n60346) );
  nor_x1_sg U63510 ( .A(n57366), .B(n60340), .X(n60341) );
  nor_x1_sg U63511 ( .A(n57378), .B(n60335), .X(n60336) );
  nor_x1_sg U63512 ( .A(n57379), .B(n60330), .X(n60331) );
  nor_x1_sg U63513 ( .A(n57379), .B(n60325), .X(n60326) );
  nor_x1_sg U63514 ( .A(n57359), .B(n60320), .X(n60321) );
  nor_x1_sg U63515 ( .A(n57360), .B(n60315), .X(n60316) );
  nor_x1_sg U63516 ( .A(n57377), .B(n60310), .X(n60311) );
  nor_x1_sg U63517 ( .A(n57365), .B(n60305), .X(n60306) );
  nor_x1_sg U63518 ( .A(n57390), .B(n60300), .X(n60301) );
  nor_x1_sg U63519 ( .A(n57375), .B(n60295), .X(n60296) );
  nor_x1_sg U63520 ( .A(n57350), .B(n60290), .X(n60291) );
  nor_x1_sg U63521 ( .A(n57378), .B(n60285), .X(n60286) );
  nor_x1_sg U63522 ( .A(n57373), .B(n60280), .X(n60281) );
  nor_x1_sg U63523 ( .A(n57390), .B(n60275), .X(n60276) );
  nor_x1_sg U63524 ( .A(n57376), .B(n60270), .X(n60271) );
  nor_x1_sg U63525 ( .A(n57377), .B(n60265), .X(n60266) );
  nor_x1_sg U63526 ( .A(n57359), .B(n60260), .X(n60261) );
  nor_x1_sg U63527 ( .A(n57376), .B(n60255), .X(n60256) );
  nor_x1_sg U63528 ( .A(n57377), .B(n60250), .X(n60251) );
  nor_x1_sg U63529 ( .A(n57372), .B(n60245), .X(n60246) );
  nor_x1_sg U63530 ( .A(n57368), .B(n60240), .X(n60241) );
  nor_x1_sg U63531 ( .A(n57388), .B(n60235), .X(n60236) );
  nor_x1_sg U63532 ( .A(n57359), .B(n60230), .X(n60231) );
  nor_x1_sg U63533 ( .A(n57360), .B(n60225), .X(n60226) );
  nor_x1_sg U63534 ( .A(n57357), .B(n60220), .X(n60221) );
  nor_x1_sg U63535 ( .A(n57358), .B(n60215), .X(n60216) );
  nor_x1_sg U63536 ( .A(n57367), .B(n60210), .X(n60211) );
  nor_x1_sg U63537 ( .A(n57368), .B(n60205), .X(n60206) );
  nor_x1_sg U63538 ( .A(n57365), .B(n60200), .X(n60201) );
  nor_x1_sg U63539 ( .A(n57366), .B(n60195), .X(n60196) );
  nor_x1_sg U63540 ( .A(n57367), .B(n60190), .X(n60191) );
  nor_x1_sg U63541 ( .A(n57379), .B(n60185), .X(n60186) );
  nor_x1_sg U63542 ( .A(n57378), .B(n60180), .X(n60181) );
  nor_x1_sg U63543 ( .A(n57379), .B(n60175), .X(n60176) );
  nor_x1_sg U63544 ( .A(n57375), .B(n60170), .X(n60171) );
  nor_x1_sg U63545 ( .A(n57376), .B(n60165), .X(n60166) );
  nor_x1_sg U63546 ( .A(n57387), .B(n60160), .X(n60161) );
  nor_x1_sg U63547 ( .A(n57375), .B(n60155), .X(n60156) );
  nor_x1_sg U63548 ( .A(n57387), .B(n60150), .X(n60151) );
  nor_x1_sg U63549 ( .A(n57366), .B(n60145), .X(n60146) );
  nor_x1_sg U63550 ( .A(n57377), .B(n60140), .X(n60141) );
  nor_x1_sg U63551 ( .A(n57377), .B(n60135), .X(n60136) );
  nor_x1_sg U63552 ( .A(n57357), .B(n60130), .X(n60131) );
  nor_x1_sg U63553 ( .A(n57358), .B(n60125), .X(n60126) );
  nor_x1_sg U63554 ( .A(n57388), .B(n60120), .X(n60121) );
  nor_x1_sg U63555 ( .A(n57375), .B(n60115), .X(n60116) );
  nor_x1_sg U63556 ( .A(n57375), .B(n60110), .X(n60111) );
  nor_x1_sg U63557 ( .A(n57387), .B(n60105), .X(n60106) );
  nor_x1_sg U63558 ( .A(n57374), .B(n60100), .X(n60101) );
  nor_x1_sg U63559 ( .A(n57387), .B(n60095), .X(n60096) );
  nor_x1_sg U63560 ( .A(n57352), .B(n60090), .X(n60091) );
  nor_x1_sg U63561 ( .A(n57378), .B(n60085), .X(n60086) );
  nor_x1_sg U63562 ( .A(n57379), .B(n60080), .X(n60081) );
  nor_x1_sg U63563 ( .A(n57377), .B(n60075), .X(n60076) );
  nor_x1_sg U63564 ( .A(n57377), .B(n60070), .X(n60071) );
  nor_x1_sg U63565 ( .A(n57375), .B(n60065), .X(n60066) );
  nor_x1_sg U63566 ( .A(n57374), .B(n60060), .X(n60061) );
  nor_x1_sg U63567 ( .A(n57366), .B(n60055), .X(n60056) );
  nor_x1_sg U63568 ( .A(n57390), .B(n60050), .X(n60051) );
  nor_x1_sg U63569 ( .A(n57381), .B(n60045), .X(n60046) );
  nor_x1_sg U63570 ( .A(n57373), .B(n60040), .X(n60041) );
  nor_x1_sg U63571 ( .A(n57374), .B(n60035), .X(n60036) );
  nor_x1_sg U63572 ( .A(n57350), .B(n60030), .X(n60031) );
  nor_x1_sg U63573 ( .A(n57350), .B(n60025), .X(n60026) );
  nor_x1_sg U63574 ( .A(n57378), .B(n60020), .X(n60021) );
  nor_x1_sg U63575 ( .A(n57379), .B(n60015), .X(n60016) );
  nor_x1_sg U63576 ( .A(n57357), .B(n60010), .X(n60011) );
  nor_x1_sg U63577 ( .A(n57358), .B(n60005), .X(n60006) );
  nor_x1_sg U63578 ( .A(n57388), .B(n60000), .X(n60001) );
  nor_x1_sg U63579 ( .A(n57373), .B(n59995), .X(n59996) );
  nor_x1_sg U63580 ( .A(n57374), .B(n59990), .X(n59991) );
  nor_x1_sg U63581 ( .A(n57351), .B(n59985), .X(n59986) );
  nor_x1_sg U63582 ( .A(n57373), .B(n59980), .X(n59981) );
  nor_x1_sg U63583 ( .A(n57387), .B(n59975), .X(n59976) );
  nor_x1_sg U63584 ( .A(n57376), .B(n59970), .X(n59971) );
  nor_x1_sg U63585 ( .A(n57368), .B(n59965), .X(n59966) );
  nor_x1_sg U63586 ( .A(n57388), .B(n59960), .X(n59961) );
  nor_x1_sg U63587 ( .A(n57387), .B(n59955), .X(n59956) );
  nor_x1_sg U63588 ( .A(n57351), .B(n59950), .X(n59951) );
  nor_x1_sg U63589 ( .A(n57367), .B(n59945), .X(n59946) );
  nor_x1_sg U63590 ( .A(n57368), .B(n59940), .X(n59941) );
  nor_x1_sg U63591 ( .A(n57387), .B(n59935), .X(n59936) );
  nor_x1_sg U63592 ( .A(n57378), .B(n59930), .X(n59931) );
  nor_x1_sg U63593 ( .A(n57373), .B(n59925), .X(n59926) );
  nor_x1_sg U63594 ( .A(n57357), .B(n59920), .X(n59921) );
  nor_x1_sg U63595 ( .A(n57358), .B(n59915), .X(n59916) );
  nor_x1_sg U63596 ( .A(n57365), .B(n59910), .X(n59911) );
  nor_x1_sg U63597 ( .A(n57375), .B(n59905), .X(n59906) );
  nor_x1_sg U63598 ( .A(n57351), .B(n59900), .X(n59901) );
  nor_x1_sg U63599 ( .A(n57367), .B(n59895), .X(n59896) );
  nor_x1_sg U63600 ( .A(n57368), .B(n59890), .X(n59891) );
  nor_x1_sg U63601 ( .A(n57365), .B(n59885), .X(n59886) );
  nor_x1_sg U63602 ( .A(n57366), .B(n59880), .X(n59881) );
  nor_x1_sg U63603 ( .A(n57359), .B(n59875), .X(n59876) );
  nor_x1_sg U63604 ( .A(n57360), .B(n59870), .X(n59871) );
  nor_x1_sg U63605 ( .A(n57357), .B(n59865), .X(n59866) );
  nor_x1_sg U63606 ( .A(n57358), .B(n59860), .X(n59861) );
  nor_x1_sg U63607 ( .A(n57371), .B(n59855), .X(n59856) );
  nor_x1_sg U63608 ( .A(n57379), .B(n59850), .X(n59851) );
  nor_x1_sg U63609 ( .A(n57379), .B(n59845), .X(n59846) );
  nor_x1_sg U63610 ( .A(n57376), .B(n59840), .X(n59841) );
  nor_x1_sg U63611 ( .A(n57387), .B(n59835), .X(n59836) );
  nor_x1_sg U63612 ( .A(n57379), .B(n59830), .X(n59831) );
  nor_x1_sg U63613 ( .A(n57377), .B(n59825), .X(n59826) );
  nor_x1_sg U63614 ( .A(n57379), .B(n59820), .X(n59821) );
  nor_x1_sg U63615 ( .A(n57375), .B(n59815), .X(n59816) );
  nor_x1_sg U63616 ( .A(n57375), .B(n59810), .X(n59811) );
  nor_x1_sg U63617 ( .A(n57360), .B(n59805), .X(n59806) );
  nor_x1_sg U63618 ( .A(n57367), .B(n59800), .X(n59801) );
  nor_x1_sg U63619 ( .A(n57350), .B(n59795), .X(n59796) );
  nor_x1_sg U63620 ( .A(n57373), .B(n59790), .X(n59791) );
  nor_x1_sg U63621 ( .A(n57376), .B(n59785), .X(n59786) );
  nor_x1_sg U63622 ( .A(n57366), .B(n59780), .X(n59781) );
  nor_x1_sg U63623 ( .A(n57375), .B(n59775), .X(n59776) );
  nor_x1_sg U63624 ( .A(n57352), .B(n59770), .X(n59771) );
  nor_x1_sg U63625 ( .A(n57367), .B(n59765), .X(n59766) );
  nor_x1_sg U63626 ( .A(n57371), .B(n59760), .X(n59761) );
  nor_x1_sg U63627 ( .A(n57371), .B(n59755), .X(n59756) );
  nor_x1_sg U63628 ( .A(n57388), .B(n59750), .X(n59751) );
  nor_x1_sg U63629 ( .A(n57374), .B(n59745), .X(n59746) );
  nor_x1_sg U63630 ( .A(n57374), .B(n59740), .X(n59741) );
  nor_x1_sg U63631 ( .A(n57358), .B(n59735), .X(n59736) );
  nor_x1_sg U63632 ( .A(n57352), .B(n59730), .X(n59731) );
  nor_x1_sg U63633 ( .A(n57374), .B(n59725), .X(n59726) );
  nor_x1_sg U63634 ( .A(n57378), .B(n59720), .X(n59721) );
  nor_x1_sg U63635 ( .A(n57379), .B(n59715), .X(n59716) );
  nor_x1_sg U63636 ( .A(n57377), .B(n59710), .X(n59711) );
  nor_x1_sg U63637 ( .A(n57378), .B(n59705), .X(n59706) );
  nor_x1_sg U63638 ( .A(n57378), .B(n59700), .X(n59701) );
  nor_x1_sg U63639 ( .A(n57369), .B(n59695), .X(n59696) );
  nor_x1_sg U63640 ( .A(n57369), .B(n59690), .X(n59691) );
  nor_x1_sg U63641 ( .A(n57369), .B(n59685), .X(n59686) );
  nor_x1_sg U63642 ( .A(n57369), .B(n59680), .X(n59681) );
  nor_x1_sg U63643 ( .A(n57369), .B(n59675), .X(n59676) );
  nor_x1_sg U63644 ( .A(n57369), .B(n59670), .X(n59671) );
  nor_x1_sg U63645 ( .A(n57369), .B(n59665), .X(n59666) );
  nor_x1_sg U63646 ( .A(n57369), .B(n59660), .X(n59661) );
  nor_x1_sg U63647 ( .A(n57369), .B(n59655), .X(n59656) );
  nor_x1_sg U63648 ( .A(n57370), .B(n59650), .X(n59651) );
  nor_x1_sg U63649 ( .A(n57370), .B(n59645), .X(n59646) );
  nor_x1_sg U63650 ( .A(n57370), .B(n59640), .X(n59641) );
  nor_x1_sg U63651 ( .A(n57370), .B(n59635), .X(n59636) );
  nor_x1_sg U63652 ( .A(n57370), .B(n59630), .X(n59631) );
  nor_x1_sg U63653 ( .A(n57370), .B(n59625), .X(n59626) );
  nor_x1_sg U63654 ( .A(n57370), .B(n59620), .X(n59621) );
  nor_x1_sg U63655 ( .A(n57370), .B(n59615), .X(n59616) );
  nor_x1_sg U63656 ( .A(n57370), .B(n59610), .X(n59611) );
  nor_x1_sg U63657 ( .A(n57371), .B(n59605), .X(n59606) );
  nor_x1_sg U63658 ( .A(n57371), .B(n59600), .X(n59601) );
  nor_x1_sg U63659 ( .A(n57371), .B(n59595), .X(n59596) );
  nor_x1_sg U63660 ( .A(n57371), .B(n59590), .X(n59591) );
  nor_x1_sg U63661 ( .A(n57371), .B(n59585), .X(n59586) );
  nor_x1_sg U63662 ( .A(n57371), .B(n59580), .X(n59581) );
  nor_x1_sg U63663 ( .A(n57371), .B(n59575), .X(n59576) );
  nor_x1_sg U63664 ( .A(n57371), .B(n59570), .X(n59571) );
  nor_x1_sg U63665 ( .A(n57371), .B(n59565), .X(n59566) );
  nor_x1_sg U63666 ( .A(n57372), .B(n59560), .X(n59561) );
  nor_x1_sg U63667 ( .A(n57372), .B(n59555), .X(n59556) );
  nor_x1_sg U63668 ( .A(n57372), .B(n59550), .X(n59551) );
  nor_x1_sg U63669 ( .A(n57372), .B(n59545), .X(n59546) );
  nor_x1_sg U63670 ( .A(n57372), .B(n59540), .X(n59541) );
  nor_x1_sg U63671 ( .A(n57372), .B(n59535), .X(n59536) );
  nor_x1_sg U63672 ( .A(n57372), .B(n59530), .X(n59531) );
  nor_x1_sg U63673 ( .A(n57372), .B(n59525), .X(n59526) );
  nor_x1_sg U63674 ( .A(n57372), .B(n59520), .X(n59521) );
  nor_x1_sg U63675 ( .A(n57350), .B(n59515), .X(n59516) );
  nor_x1_sg U63676 ( .A(n57350), .B(n59510), .X(n59511) );
  nor_x1_sg U63677 ( .A(n57352), .B(n59505), .X(n59506) );
  nor_x1_sg U63678 ( .A(n57350), .B(n59500), .X(n59501) );
  nor_x1_sg U63679 ( .A(n57352), .B(n59495), .X(n59496) );
  nor_x1_sg U63680 ( .A(n57351), .B(n59490), .X(n59491) );
  nor_x1_sg U63681 ( .A(n57350), .B(n59485), .X(n59486) );
  nor_x1_sg U63682 ( .A(n57352), .B(n59480), .X(n59481) );
  nor_x1_sg U63683 ( .A(n57352), .B(n59475), .X(n59476) );
  nor_x1_sg U63684 ( .A(n57351), .B(n59470), .X(n59471) );
  nor_x1_sg U63685 ( .A(n57351), .B(n59465), .X(n59466) );
  nor_x1_sg U63686 ( .A(n57373), .B(n59460), .X(n59461) );
  nor_x1_sg U63687 ( .A(n57390), .B(n59455), .X(n59456) );
  nor_x1_sg U63688 ( .A(n57374), .B(n59450), .X(n59451) );
  nor_x1_sg U63689 ( .A(n57351), .B(n59445), .X(n59446) );
  nor_x1_sg U63690 ( .A(n57351), .B(n59440), .X(n59441) );
  nor_x1_sg U63691 ( .A(n57375), .B(n59435), .X(n59436) );
  nor_x1_sg U63692 ( .A(n57390), .B(n59430), .X(n59431) );
  nor_x1_sg U63693 ( .A(n57373), .B(n59425), .X(n59426) );
  nor_x1_sg U63694 ( .A(n57373), .B(n59420), .X(n59421) );
  nor_x1_sg U63695 ( .A(n57373), .B(n59415), .X(n59416) );
  nor_x1_sg U63696 ( .A(n57373), .B(n59410), .X(n59411) );
  nor_x1_sg U63697 ( .A(n57373), .B(n59405), .X(n59406) );
  nor_x1_sg U63698 ( .A(n57373), .B(n59400), .X(n59401) );
  nor_x1_sg U63699 ( .A(n57373), .B(n59395), .X(n59396) );
  nor_x1_sg U63700 ( .A(n57373), .B(n59390), .X(n59391) );
  nor_x1_sg U63701 ( .A(n57373), .B(n59385), .X(n59386) );
  nor_x1_sg U63702 ( .A(n57374), .B(n59380), .X(n59381) );
  nor_x1_sg U63703 ( .A(n57374), .B(n59375), .X(n59376) );
  nor_x1_sg U63704 ( .A(n57374), .B(n59370), .X(n59371) );
  nor_x1_sg U63705 ( .A(n57374), .B(n59365), .X(n59366) );
  nor_x1_sg U63706 ( .A(n57374), .B(n59360), .X(n59361) );
  nor_x1_sg U63707 ( .A(n57374), .B(n59355), .X(n59356) );
  nor_x1_sg U63708 ( .A(n57374), .B(n59350), .X(n59351) );
  nor_x1_sg U63709 ( .A(n57374), .B(n59345), .X(n59346) );
  nor_x1_sg U63710 ( .A(n57374), .B(n59340), .X(n59341) );
  nor_x1_sg U63711 ( .A(n57357), .B(n59335), .X(n59336) );
  nor_x1_sg U63712 ( .A(n57358), .B(n59330), .X(n59331) );
  nor_x1_sg U63713 ( .A(n57377), .B(n59325), .X(n59326) );
  nor_x1_sg U63714 ( .A(n57360), .B(n59320), .X(n59321) );
  nor_x1_sg U63715 ( .A(n57387), .B(n59315), .X(n59316) );
  nor_x1_sg U63716 ( .A(n57373), .B(n59310), .X(n59311) );
  nor_x1_sg U63717 ( .A(n57374), .B(n59305), .X(n59306) );
  nor_x1_sg U63718 ( .A(n57350), .B(n59300), .X(n59301) );
  nor_x1_sg U63719 ( .A(n57351), .B(n59295), .X(n59296) );
  nor_x1_sg U63720 ( .A(n57360), .B(n59290), .X(n59291) );
  nor_x1_sg U63721 ( .A(n57390), .B(n59285), .X(n59286) );
  nor_x1_sg U63722 ( .A(n57388), .B(n59280), .X(n59281) );
  nor_x1_sg U63723 ( .A(n57375), .B(n59275), .X(n59276) );
  nor_x1_sg U63724 ( .A(n57368), .B(n59270), .X(n59271) );
  nor_x1_sg U63725 ( .A(n57357), .B(n59265), .X(n59266) );
  nor_x1_sg U63726 ( .A(n57390), .B(n59260), .X(n59261) );
  nor_x1_sg U63727 ( .A(n57376), .B(n59255), .X(n59256) );
  nor_x1_sg U63728 ( .A(n57378), .B(n59250), .X(n59251) );
  nor_x1_sg U63729 ( .A(n57390), .B(n59245), .X(n59246) );
  nor_x1_sg U63730 ( .A(n57359), .B(n59240), .X(n59241) );
  nor_x1_sg U63731 ( .A(n57360), .B(n59235), .X(n59236) );
  nor_x1_sg U63732 ( .A(n57357), .B(n59230), .X(n59231) );
  nor_x1_sg U63733 ( .A(n57388), .B(n59225), .X(n59226) );
  nor_x1_sg U63734 ( .A(n57358), .B(n59220), .X(n59221) );
  nor_x1_sg U63735 ( .A(n57374), .B(n59215), .X(n59216) );
  nor_x1_sg U63736 ( .A(n57387), .B(n59210), .X(n59211) );
  nor_x1_sg U63737 ( .A(n57373), .B(n59205), .X(n59206) );
  nor_x1_sg U63738 ( .A(n57375), .B(n59200), .X(n59201) );
  nor_x1_sg U63739 ( .A(n57387), .B(n59195), .X(n59196) );
  nor_x1_sg U63740 ( .A(n57367), .B(n59190), .X(n59191) );
  nor_x1_sg U63741 ( .A(n57367), .B(n59185), .X(n59186) );
  nor_x1_sg U63742 ( .A(n57368), .B(n59180), .X(n59181) );
  nor_x1_sg U63743 ( .A(n57365), .B(n59175), .X(n59176) );
  nor_x1_sg U63744 ( .A(n57366), .B(n59170), .X(n59171) );
  nor_x1_sg U63745 ( .A(n57376), .B(n59165), .X(n59166) );
  nor_x1_sg U63746 ( .A(n57359), .B(n59160), .X(n59161) );
  nor_x1_sg U63747 ( .A(n57375), .B(n59155), .X(n59156) );
  nor_x1_sg U63748 ( .A(n57375), .B(n59150), .X(n59151) );
  nor_x1_sg U63749 ( .A(n57375), .B(n59145), .X(n59146) );
  nor_x1_sg U63750 ( .A(n57375), .B(n59140), .X(n59141) );
  nor_x1_sg U63751 ( .A(n57375), .B(n59135), .X(n59136) );
  nor_x1_sg U63752 ( .A(n57375), .B(n59130), .X(n59131) );
  nor_x1_sg U63753 ( .A(n57375), .B(n59125), .X(n59126) );
  nor_x1_sg U63754 ( .A(n57375), .B(n59120), .X(n59121) );
  nor_x1_sg U63755 ( .A(n57375), .B(n59115), .X(n59116) );
  nor_x1_sg U63756 ( .A(n57352), .B(n59110), .X(n59111) );
  nor_x1_sg U63757 ( .A(n57352), .B(n59105), .X(n59106) );
  nor_x1_sg U63758 ( .A(n57352), .B(n59100), .X(n59101) );
  nor_x1_sg U63759 ( .A(n57351), .B(n59095), .X(n59096) );
  nor_x1_sg U63760 ( .A(n57350), .B(n59090), .X(n59091) );
  nor_x1_sg U63761 ( .A(n57351), .B(n59085), .X(n59086) );
  nor_x1_sg U63762 ( .A(n57387), .B(n59080), .X(n59081) );
  nor_x1_sg U63763 ( .A(n57350), .B(n59075), .X(n59076) );
  nor_x1_sg U63764 ( .A(n57350), .B(n59070), .X(n59071) );
  nor_x1_sg U63765 ( .A(n57376), .B(n59065), .X(n59066) );
  nor_x1_sg U63766 ( .A(n57376), .B(n59060), .X(n59061) );
  nor_x1_sg U63767 ( .A(n57376), .B(n59055), .X(n59056) );
  nor_x1_sg U63768 ( .A(n57376), .B(n59050), .X(n59051) );
  nor_x1_sg U63769 ( .A(n57376), .B(n59045), .X(n59046) );
  nor_x1_sg U63770 ( .A(n57376), .B(n59040), .X(n59041) );
  nor_x1_sg U63771 ( .A(n57376), .B(n59035), .X(n59036) );
  nor_x1_sg U63772 ( .A(n57376), .B(n59030), .X(n59031) );
  nor_x1_sg U63773 ( .A(n57376), .B(n59025), .X(n59026) );
  nor_x1_sg U63774 ( .A(n57368), .B(n59020), .X(n59021) );
  nor_x1_sg U63775 ( .A(n57365), .B(n59015), .X(n59016) );
  nor_x1_sg U63776 ( .A(n57366), .B(n59010), .X(n59011) );
  nor_x1_sg U63777 ( .A(n57373), .B(n59005), .X(n59006) );
  nor_x1_sg U63778 ( .A(n57374), .B(n59000), .X(n59001) );
  nor_x1_sg U63779 ( .A(n57352), .B(n58995), .X(n58996) );
  nor_x1_sg U63780 ( .A(n57373), .B(n58990), .X(n58991) );
  nor_x1_sg U63781 ( .A(n57387), .B(n58985), .X(n58986) );
  nor_x1_sg U63782 ( .A(n57352), .B(n58980), .X(n58981) );
  nor_x1_sg U63783 ( .A(n57377), .B(n58975), .X(n58976) );
  nor_x1_sg U63784 ( .A(n57377), .B(n58970), .X(n58971) );
  nor_x1_sg U63785 ( .A(n57377), .B(n58965), .X(n58966) );
  nor_x1_sg U63786 ( .A(n57377), .B(n58960), .X(n58961) );
  nor_x1_sg U63787 ( .A(n57377), .B(n58955), .X(n58956) );
  nor_x1_sg U63788 ( .A(n57377), .B(n58950), .X(n58951) );
  nor_x1_sg U63789 ( .A(n57377), .B(n58945), .X(n58946) );
  nor_x1_sg U63790 ( .A(n57377), .B(n58940), .X(n58941) );
  nor_x1_sg U63791 ( .A(n57377), .B(n58935), .X(n58936) );
  nor_x1_sg U63792 ( .A(n57378), .B(n58930), .X(n58931) );
  nor_x1_sg U63793 ( .A(n57379), .B(n58925), .X(n58926) );
  nor_x1_sg U63794 ( .A(n57377), .B(n58920), .X(n58921) );
  nor_x1_sg U63795 ( .A(n57376), .B(n58915), .X(n58916) );
  nor_x1_sg U63796 ( .A(n57387), .B(n58910), .X(n58911) );
  nor_x1_sg U63797 ( .A(n57388), .B(n58905), .X(n58906) );
  nor_x1_sg U63798 ( .A(n57359), .B(n58900), .X(n58901) );
  nor_x1_sg U63799 ( .A(n57360), .B(n58895), .X(n58896) );
  nor_x1_sg U63800 ( .A(n57357), .B(n58890), .X(n58891) );
  nor_x1_sg U63801 ( .A(n57378), .B(n58885), .X(n58886) );
  nor_x1_sg U63802 ( .A(n57378), .B(n58880), .X(n58881) );
  nor_x1_sg U63803 ( .A(n57378), .B(n58875), .X(n58876) );
  nor_x1_sg U63804 ( .A(n57378), .B(n58870), .X(n58871) );
  nor_x1_sg U63805 ( .A(n57378), .B(n58865), .X(n58866) );
  nor_x1_sg U63806 ( .A(n57378), .B(n58860), .X(n58861) );
  nor_x1_sg U63807 ( .A(n57378), .B(n58855), .X(n58856) );
  nor_x1_sg U63808 ( .A(n57378), .B(n58850), .X(n58851) );
  nor_x1_sg U63809 ( .A(n57378), .B(n58845), .X(n58846) );
  nor_x1_sg U63810 ( .A(n57379), .B(n58840), .X(n58841) );
  nor_x1_sg U63811 ( .A(n57379), .B(n58835), .X(n58836) );
  nor_x1_sg U63812 ( .A(n57379), .B(n58830), .X(n58831) );
  nor_x1_sg U63813 ( .A(n57379), .B(n58825), .X(n58826) );
  nor_x1_sg U63814 ( .A(n57379), .B(n58820), .X(n58821) );
  nor_x1_sg U63815 ( .A(n57379), .B(n58815), .X(n58816) );
  nor_x1_sg U63816 ( .A(n57379), .B(n58810), .X(n58811) );
  nor_x1_sg U63817 ( .A(n57379), .B(n58805), .X(n58806) );
  nor_x1_sg U63818 ( .A(n57379), .B(n58800), .X(n58801) );
  nor_x1_sg U63819 ( .A(n57380), .B(n58795), .X(n58796) );
  nor_x1_sg U63820 ( .A(n57380), .B(n58790), .X(n58791) );
  nor_x1_sg U63821 ( .A(n57380), .B(n58785), .X(n58786) );
  nor_x1_sg U63822 ( .A(n57380), .B(n58780), .X(n58781) );
  nor_x1_sg U63823 ( .A(n57380), .B(n58775), .X(n58776) );
  nor_x1_sg U63824 ( .A(n57380), .B(n58770), .X(n58771) );
  nor_x1_sg U63825 ( .A(n57380), .B(n58765), .X(n58766) );
  nor_x1_sg U63826 ( .A(n57380), .B(n58760), .X(n58761) );
  nand_x1_sg U63827 ( .A(n53559), .B(n33098), .X(n33107) );
  nand_x1_sg U63828 ( .A(n50971), .B(n33098), .X(n33101) );
  nand_x1_sg U63829 ( .A(n53557), .B(n33098), .X(n33119) );
  nand_x1_sg U63830 ( .A(n50967), .B(n33098), .X(n33125) );
  nand_x1_sg U63831 ( .A(n50953), .B(n32926), .X(n32929) );
  nand_x1_sg U63832 ( .A(n53537), .B(n32926), .X(n32947) );
  nand_x1_sg U63833 ( .A(n53533), .B(n32926), .X(n32953) );
  nand_x1_sg U63834 ( .A(n53523), .B(n32926), .X(n32935) );
  nand_x1_sg U63835 ( .A(n50887), .B(n33613), .X(n33634) );
  nand_x1_sg U63836 ( .A(n53447), .B(n33613), .X(n33640) );
  nand_x1_sg U63837 ( .A(n50877), .B(n33613), .X(n33622) );
  nand_x1_sg U63838 ( .A(n50873), .B(n33613), .X(n33616) );
  nand_x1_sg U63839 ( .A(n50831), .B(n33140), .X(n33149) );
  nand_x1_sg U63840 ( .A(n53419), .B(n33140), .X(n33143) );
  nand_x1_sg U63841 ( .A(n53417), .B(n33140), .X(n33161) );
  nand_x1_sg U63842 ( .A(n53411), .B(n33140), .X(n33167) );
  nand_x1_sg U63843 ( .A(n50787), .B(n32969), .X(n32978) );
  nand_x1_sg U63844 ( .A(n50781), .B(n32969), .X(n32996) );
  nand_x1_sg U63845 ( .A(n53329), .B(n32969), .X(n32972) );
  nand_x1_sg U63846 ( .A(n53327), .B(n32969), .X(n32990) );
  nand_x1_sg U63847 ( .A(n53219), .B(n33443), .X(n33452) );
  nand_x1_sg U63848 ( .A(n50671), .B(n33443), .X(n33446) );
  nand_x1_sg U63849 ( .A(n53217), .B(n33443), .X(n33464) );
  nand_x1_sg U63850 ( .A(n50667), .B(n33443), .X(n33470) );
  nand_x1_sg U63851 ( .A(n50645), .B(n33012), .X(n33039) );
  nand_x1_sg U63852 ( .A(n53185), .B(n33012), .X(n33015) );
  nand_x1_sg U63853 ( .A(n53183), .B(n33012), .X(n33021) );
  nand_x1_sg U63854 ( .A(n53181), .B(n33012), .X(n33033) );
  nand_x1_sg U63855 ( .A(n53127), .B(n33314), .X(n33335) );
  nand_x1_sg U63856 ( .A(n53123), .B(n33314), .X(n33317) );
  nand_x1_sg U63857 ( .A(n53121), .B(n33314), .X(n33341) );
  nand_x1_sg U63858 ( .A(n50597), .B(n33314), .X(n33323) );
  nand_x1_sg U63859 ( .A(n50587), .B(n33356), .X(n33377) );
  nand_x1_sg U63860 ( .A(n53107), .B(n33356), .X(n33383) );
  nand_x1_sg U63861 ( .A(n50577), .B(n33356), .X(n33365) );
  nand_x1_sg U63862 ( .A(n50573), .B(n33356), .X(n33359) );
  nand_x1_sg U63863 ( .A(n50487), .B(n33055), .X(n33064) );
  nand_x1_sg U63864 ( .A(n50481), .B(n33055), .X(n33082) );
  nand_x1_sg U63865 ( .A(n52989), .B(n33055), .X(n33058) );
  nand_x1_sg U63866 ( .A(n52987), .B(n33055), .X(n33076) );
  nand_x1_sg U63867 ( .A(n50975), .B(n57266), .X(n33095) );
  nand_x1_sg U63868 ( .A(n53563), .B(n57266), .X(n33115) );
  nand_x1_sg U63869 ( .A(n53561), .B(n57265), .X(n33117) );
  nand_x1_sg U63870 ( .A(n50973), .B(n57266), .X(n33109) );
  nand_x1_sg U63871 ( .A(n53555), .B(n57265), .X(n33123) );
  nand_x1_sg U63872 ( .A(n53553), .B(n57266), .X(n33127) );
  nand_x1_sg U63873 ( .A(n50965), .B(n57265), .X(n33099) );
  nand_x1_sg U63874 ( .A(n50961), .B(n57265), .X(n33105) );
  nand_x1_sg U63875 ( .A(n53547), .B(n57266), .X(n33133) );
  nand_x1_sg U63876 ( .A(n53545), .B(n57265), .X(n33135) );
  nand_x1_sg U63877 ( .A(n50959), .B(n57282), .X(n32943) );
  nand_x1_sg U63878 ( .A(n53541), .B(n57281), .X(n32927) );
  nand_x1_sg U63879 ( .A(n50955), .B(n57281), .X(n32945) );
  nand_x1_sg U63880 ( .A(n53539), .B(n57282), .X(n32937) );
  nand_x1_sg U63881 ( .A(n50951), .B(n57282), .X(n32923) );
  nand_x1_sg U63882 ( .A(n50949), .B(n57281), .X(n32951) );
  nand_x1_sg U63883 ( .A(n50947), .B(n57282), .X(n32955) );
  nand_x1_sg U63884 ( .A(n53529), .B(n57281), .X(n32933) );
  nand_x1_sg U63885 ( .A(n53525), .B(n57282), .X(n32961) );
  nand_x1_sg U63886 ( .A(n53521), .B(n57281), .X(n32963) );
  nand_x1_sg U63887 ( .A(n50893), .B(n57221), .X(n33630) );
  nand_x1_sg U63888 ( .A(n50889), .B(n57220), .X(n33632) );
  nand_x1_sg U63889 ( .A(n53449), .B(n57221), .X(n33624) );
  nand_x1_sg U63890 ( .A(n50881), .B(n57220), .X(n33638) );
  nand_x1_sg U63891 ( .A(n50879), .B(n57220), .X(n33614) );
  nand_x1_sg U63892 ( .A(n50875), .B(n57221), .X(n33642) );
  nand_x1_sg U63893 ( .A(n53443), .B(n57220), .X(n33620) );
  nand_x1_sg U63894 ( .A(n53441), .B(n57221), .X(n33648) );
  nand_x1_sg U63895 ( .A(n53439), .B(n57221), .X(n33610) );
  nand_x1_sg U63896 ( .A(n53437), .B(n57220), .X(n33650) );
  nand_x1_sg U63897 ( .A(n53427), .B(n57262), .X(n33137) );
  nand_x1_sg U63898 ( .A(n53425), .B(n57262), .X(n33157) );
  nand_x1_sg U63899 ( .A(n53423), .B(n57261), .X(n33159) );
  nand_x1_sg U63900 ( .A(n53421), .B(n57262), .X(n33151) );
  nand_x1_sg U63901 ( .A(n53413), .B(n57261), .X(n33165) );
  nand_x1_sg U63902 ( .A(n53409), .B(n57262), .X(n33169) );
  nand_x1_sg U63903 ( .A(n53407), .B(n57261), .X(n33141) );
  nand_x1_sg U63904 ( .A(n53401), .B(n57261), .X(n33147) );
  nand_x1_sg U63905 ( .A(n53399), .B(n57262), .X(n33175) );
  nand_x1_sg U63906 ( .A(n53397), .B(n57261), .X(n33177) );
  nand_x1_sg U63907 ( .A(n50795), .B(n57277), .X(n32994) );
  nand_x1_sg U63908 ( .A(n50791), .B(n57278), .X(n33004) );
  nand_x1_sg U63909 ( .A(n50789), .B(n57277), .X(n32970) );
  nand_x1_sg U63910 ( .A(n53341), .B(n57278), .X(n32998) );
  nand_x1_sg U63911 ( .A(n50785), .B(n57278), .X(n32966) );
  nand_x1_sg U63912 ( .A(n50783), .B(n57277), .X(n32976) );
  nand_x1_sg U63913 ( .A(n53335), .B(n57277), .X(n33006) );
  nand_x1_sg U63914 ( .A(n53333), .B(n57277), .X(n32988) );
  nand_x1_sg U63915 ( .A(n53331), .B(n57278), .X(n32980) );
  nand_x1_sg U63916 ( .A(n53325), .B(n57278), .X(n32986) );
  nand_x1_sg U63917 ( .A(n50675), .B(n57234), .X(n33440) );
  nand_x1_sg U63918 ( .A(n53223), .B(n57234), .X(n33460) );
  nand_x1_sg U63919 ( .A(n53221), .B(n57233), .X(n33462) );
  nand_x1_sg U63920 ( .A(n50673), .B(n57234), .X(n33454) );
  nand_x1_sg U63921 ( .A(n53215), .B(n57233), .X(n33468) );
  nand_x1_sg U63922 ( .A(n53213), .B(n57234), .X(n33472) );
  nand_x1_sg U63923 ( .A(n50665), .B(n57233), .X(n33444) );
  nand_x1_sg U63924 ( .A(n50661), .B(n57233), .X(n33450) );
  nand_x1_sg U63925 ( .A(n53207), .B(n57234), .X(n33478) );
  nand_x1_sg U63926 ( .A(n53205), .B(n57233), .X(n33480) );
  nand_x1_sg U63927 ( .A(n50659), .B(n57274), .X(n33047) );
  nand_x1_sg U63928 ( .A(n53201), .B(n57273), .X(n33019) );
  nand_x1_sg U63929 ( .A(n50653), .B(n57274), .X(n33041) );
  nand_x1_sg U63930 ( .A(n53197), .B(n57273), .X(n33013) );
  nand_x1_sg U63931 ( .A(n53195), .B(n57274), .X(n33009) );
  nand_x1_sg U63932 ( .A(n50649), .B(n57273), .X(n33037) );
  nand_x1_sg U63933 ( .A(n53193), .B(n57274), .X(n33029) );
  nand_x1_sg U63934 ( .A(n50647), .B(n57273), .X(n33049) );
  nand_x1_sg U63935 ( .A(n53191), .B(n57274), .X(n33023) );
  nand_x1_sg U63936 ( .A(n53189), .B(n57273), .X(n33031) );
  nand_x1_sg U63937 ( .A(n53137), .B(n57245), .X(n33321) );
  nand_x1_sg U63938 ( .A(n53135), .B(n57246), .X(n33331) );
  nand_x1_sg U63939 ( .A(n53133), .B(n57245), .X(n33333) );
  nand_x1_sg U63940 ( .A(n50601), .B(n57246), .X(n33325) );
  nand_x1_sg U63941 ( .A(n53131), .B(n57246), .X(n33311) );
  nand_x1_sg U63942 ( .A(n53129), .B(n57245), .X(n33315) );
  nand_x1_sg U63943 ( .A(n53125), .B(n57245), .X(n33339) );
  nand_x1_sg U63944 ( .A(n53119), .B(n57246), .X(n33343) );
  nand_x1_sg U63945 ( .A(n53113), .B(n57246), .X(n33349) );
  nand_x1_sg U63946 ( .A(n53111), .B(n57245), .X(n33351) );
  nand_x1_sg U63947 ( .A(n50593), .B(n57242), .X(n33373) );
  nand_x1_sg U63948 ( .A(n50589), .B(n57241), .X(n33375) );
  nand_x1_sg U63949 ( .A(n53109), .B(n57242), .X(n33367) );
  nand_x1_sg U63950 ( .A(n50581), .B(n57241), .X(n33381) );
  nand_x1_sg U63951 ( .A(n50579), .B(n57241), .X(n33357) );
  nand_x1_sg U63952 ( .A(n50575), .B(n57242), .X(n33385) );
  nand_x1_sg U63953 ( .A(n53103), .B(n57241), .X(n33363) );
  nand_x1_sg U63954 ( .A(n53101), .B(n57242), .X(n33391) );
  nand_x1_sg U63955 ( .A(n53099), .B(n57242), .X(n33353) );
  nand_x1_sg U63956 ( .A(n53097), .B(n57241), .X(n33393) );
  nand_x1_sg U63957 ( .A(n50495), .B(n57269), .X(n33080) );
  nand_x1_sg U63958 ( .A(n50491), .B(n57270), .X(n33090) );
  nand_x1_sg U63959 ( .A(n50489), .B(n57269), .X(n33056) );
  nand_x1_sg U63960 ( .A(n53001), .B(n57270), .X(n33084) );
  nand_x1_sg U63961 ( .A(n50485), .B(n57270), .X(n33052) );
  nand_x1_sg U63962 ( .A(n50483), .B(n57269), .X(n33062) );
  nand_x1_sg U63963 ( .A(n52995), .B(n57269), .X(n33092) );
  nand_x1_sg U63964 ( .A(n52993), .B(n57269), .X(n33074) );
  nand_x1_sg U63965 ( .A(n52991), .B(n57270), .X(n33066) );
  nand_x1_sg U63966 ( .A(n52985), .B(n57270), .X(n33072) );
  nand_x1_sg U63967 ( .A(n53549), .B(n33098), .X(n33131) );
  nand_x1_sg U63968 ( .A(n50963), .B(n33098), .X(n33113) );
  nand_x1_sg U63969 ( .A(n50945), .B(n32926), .X(n32959) );
  nand_x1_sg U63970 ( .A(n53527), .B(n32926), .X(n32941) );
  nand_x1_sg U63971 ( .A(n50871), .B(n33613), .X(n33646) );
  nand_x1_sg U63972 ( .A(n50869), .B(n33613), .X(n33628) );
  nand_x1_sg U63973 ( .A(n50829), .B(n33140), .X(n33173) );
  nand_x1_sg U63974 ( .A(n53403), .B(n33140), .X(n33155) );
  nand_x1_sg U63975 ( .A(n53347), .B(n32969), .X(n32984) );
  nand_x1_sg U63976 ( .A(n53343), .B(n32969), .X(n33002) );
  nand_x1_sg U63977 ( .A(n53209), .B(n33443), .X(n33476) );
  nand_x1_sg U63978 ( .A(n50663), .B(n33443), .X(n33458) );
  nand_x1_sg U63979 ( .A(n50657), .B(n33012), .X(n33027) );
  nand_x1_sg U63980 ( .A(n53199), .B(n33012), .X(n33045) );
  nand_x1_sg U63981 ( .A(n53115), .B(n33314), .X(n33329) );
  nand_x1_sg U63982 ( .A(n50595), .B(n33314), .X(n33347) );
  nand_x1_sg U63983 ( .A(n50571), .B(n33356), .X(n33389) );
  nand_x1_sg U63984 ( .A(n50569), .B(n33356), .X(n33371) );
  nand_x1_sg U63985 ( .A(n53007), .B(n33055), .X(n33070) );
  nand_x1_sg U63986 ( .A(n53003), .B(n33055), .X(n33088) );
  nand_x1_sg U63987 ( .A(n53567), .B(n57266), .X(n33103) );
  nand_x1_sg U63988 ( .A(n53565), .B(n57265), .X(n33111) );
  nand_x1_sg U63989 ( .A(n50969), .B(n57266), .X(n33121) );
  nand_x1_sg U63990 ( .A(n53551), .B(n57265), .X(n33129) );
  nand_x1_sg U63991 ( .A(n50957), .B(n57281), .X(n32939) );
  nand_x1_sg U63992 ( .A(n53543), .B(n57282), .X(n32931) );
  nand_x1_sg U63993 ( .A(n53535), .B(n57282), .X(n32949) );
  nand_x1_sg U63994 ( .A(n53531), .B(n57281), .X(n32957) );
  nand_x1_sg U63995 ( .A(n50891), .B(n57220), .X(n33626) );
  nand_x1_sg U63996 ( .A(n50885), .B(n57221), .X(n33618) );
  nand_x1_sg U63997 ( .A(n50883), .B(n57221), .X(n33636) );
  nand_x1_sg U63998 ( .A(n53445), .B(n57220), .X(n33644) );
  nand_x1_sg U63999 ( .A(n50835), .B(n57262), .X(n33145) );
  nand_x1_sg U64000 ( .A(n50833), .B(n57261), .X(n33153) );
  nand_x1_sg U64001 ( .A(n53415), .B(n57262), .X(n33163) );
  nand_x1_sg U64002 ( .A(n53405), .B(n57261), .X(n33171) );
  nand_x1_sg U64003 ( .A(n53345), .B(n57278), .X(n32974) );
  nand_x1_sg U64004 ( .A(n50793), .B(n57278), .X(n32992) );
  nand_x1_sg U64005 ( .A(n53339), .B(n57277), .X(n33000) );
  nand_x1_sg U64006 ( .A(n53337), .B(n57277), .X(n32982) );
  nand_x1_sg U64007 ( .A(n53227), .B(n57234), .X(n33448) );
  nand_x1_sg U64008 ( .A(n53225), .B(n57233), .X(n33456) );
  nand_x1_sg U64009 ( .A(n50669), .B(n57234), .X(n33466) );
  nand_x1_sg U64010 ( .A(n53211), .B(n57233), .X(n33474) );
  nand_x1_sg U64011 ( .A(n53203), .B(n57274), .X(n33017) );
  nand_x1_sg U64012 ( .A(n50655), .B(n57274), .X(n33035) );
  nand_x1_sg U64013 ( .A(n50651), .B(n57273), .X(n33025) );
  nand_x1_sg U64014 ( .A(n53187), .B(n57273), .X(n33043) );
  nand_x1_sg U64015 ( .A(n53141), .B(n57246), .X(n33319) );
  nand_x1_sg U64016 ( .A(n53139), .B(n57245), .X(n33327) );
  nand_x1_sg U64017 ( .A(n50599), .B(n57246), .X(n33337) );
  nand_x1_sg U64018 ( .A(n53117), .B(n57245), .X(n33345) );
  nand_x1_sg U64019 ( .A(n50591), .B(n57241), .X(n33369) );
  nand_x1_sg U64020 ( .A(n50585), .B(n57242), .X(n33361) );
  nand_x1_sg U64021 ( .A(n50583), .B(n57242), .X(n33379) );
  nand_x1_sg U64022 ( .A(n53105), .B(n57241), .X(n33387) );
  nand_x1_sg U64023 ( .A(n53005), .B(n57270), .X(n33060) );
  nand_x1_sg U64024 ( .A(n50493), .B(n57270), .X(n33078) );
  nand_x1_sg U64025 ( .A(n52999), .B(n57269), .X(n33086) );
  nand_x1_sg U64026 ( .A(n52997), .B(n57269), .X(n33068) );
  nand_x1_sg U64027 ( .A(n26113), .B(n51019), .X(n26296) );
  nor_x1_sg U64028 ( .A(n57430), .B(n58648), .X(n58649) );
  nor_x1_sg U64029 ( .A(n57079), .B(n32057), .X(n32056) );
  nand_x2_sg U64030 ( .A(n32058), .B(n32059), .X(n32053) );
  nand_x2_sg U64031 ( .A(n58650), .B(n58649), .X(n32054) );
  nor_x1_sg U64032 ( .A(n57087), .B(n51553), .X(n32058) );
  nand_x1_sg U64033 ( .A(n47775), .B(n31968), .X(n31970) );
  nor_x1_sg U64034 ( .A(n31971), .B(n46857), .X(n31969) );
  nand_x1_sg U64035 ( .A(n57097), .B(n31968), .X(n31991) );
  nor_x1_sg U64036 ( .A(n31996), .B(n46885), .X(n31990) );
  nor_x1_sg U64037 ( .A(n31998), .B(n31974), .X(n31997) );
  nand_x2_sg U64038 ( .A(n26291), .B(n26292), .X(n26290) );
  nand_x1_sg U64039 ( .A(n57106), .B(n47585), .X(n26291) );
  nand_x1_sg U64040 ( .A(n57109), .B(n51045), .X(n26292) );
  nor_x1_sg U64041 ( .A(n57442), .B(n58609), .X(n58610) );
  nor_x1_sg U64042 ( .A(n57077), .B(n32500), .X(n32499) );
  nand_x2_sg U64043 ( .A(n32504), .B(n32505), .X(n32496) );
  nand_x2_sg U64044 ( .A(n58611), .B(n58610), .X(n32497) );
  nor_x1_sg U64045 ( .A(n57083), .B(n51551), .X(n32504) );
  nand_x1_sg U64046 ( .A(n47445), .B(n32368), .X(n32367) );
  nor_x1_sg U64047 ( .A(n32369), .B(n32370), .X(n32366) );
  nor_x1_sg U64048 ( .A(n57390), .B(n58660), .X(n58661) );
  nand_x1_sg U64049 ( .A(n51001), .B(n26113), .X(n26331) );
  nand_x1_sg U64050 ( .A(n26091), .B(n51027), .X(n26278) );
  nor_x1_sg U64051 ( .A(n26275), .B(n26276), .X(n26274) );
  nand_x2_sg U64052 ( .A(n26279), .B(n26280), .X(n26275) );
  nand_x2_sg U64053 ( .A(n26277), .B(n26278), .X(n26276) );
  nand_x1_sg U64054 ( .A(n57111), .B(n51025), .X(n26280) );
  nand_x1_sg U64055 ( .A(n47587), .B(n57111), .X(n26334) );
  nand_x1_sg U64056 ( .A(n51047), .B(n57109), .X(n26335) );
  nand_x1_sg U64057 ( .A(n51049), .B(n26121), .X(n26267) );
  nand_x1_sg U64058 ( .A(n51013), .B(n26121), .X(n26301) );
  nand_x1_sg U64059 ( .A(n47597), .B(n26122), .X(n26268) );
  nand_x2_sg U64060 ( .A(n57308), .B(n67530), .X(n26330) );
  nor_x1_sg U64061 ( .A(n67530), .B(n51069), .X(n26326) );
  nand_x1_sg U64062 ( .A(n57286), .B(n53435), .X(n32878) );
  nand_x1_sg U64063 ( .A(n57286), .B(n53433), .X(n32882) );
  nand_x1_sg U64064 ( .A(n57286), .B(n50867), .X(n32884) );
  nand_x1_sg U64065 ( .A(n57286), .B(n50863), .X(n32890) );
  nand_x1_sg U64066 ( .A(n57286), .B(n50861), .X(n32888) );
  nand_x1_sg U64067 ( .A(n57286), .B(n53431), .X(n32892) );
  nand_x1_sg U64068 ( .A(n57286), .B(n50859), .X(n32906) );
  nand_x1_sg U64069 ( .A(n32881), .B(n50855), .X(n32908) );
  nand_x1_sg U64070 ( .A(n57286), .B(n50851), .X(n32910) );
  nand_x1_sg U64071 ( .A(n57286), .B(n50849), .X(n32898) );
  nand_x1_sg U64072 ( .A(n57286), .B(n50845), .X(n32900) );
  nand_x1_sg U64073 ( .A(n57286), .B(n50843), .X(n32902) );
  nand_x1_sg U64074 ( .A(n57286), .B(n50841), .X(n32916) );
  nand_x1_sg U64075 ( .A(n57286), .B(n50837), .X(n32918) );
  nand_x1_sg U64076 ( .A(n57290), .B(n50567), .X(n32836) );
  nand_x1_sg U64077 ( .A(n57290), .B(n53095), .X(n32838) );
  nand_x1_sg U64078 ( .A(n57290), .B(n50563), .X(n32842) );
  nand_x1_sg U64079 ( .A(n32835), .B(n50561), .X(n32844) );
  nand_x1_sg U64080 ( .A(n57290), .B(n50559), .X(n32846) );
  nand_x1_sg U64081 ( .A(n57290), .B(n50555), .X(n32852) );
  nand_x1_sg U64082 ( .A(n57290), .B(n50553), .X(n32862) );
  nand_x1_sg U64083 ( .A(n57290), .B(n50551), .X(n32854) );
  nand_x1_sg U64084 ( .A(n57290), .B(n50549), .X(n32864) );
  nand_x1_sg U64085 ( .A(n57290), .B(n50547), .X(n32856) );
  nand_x1_sg U64086 ( .A(n57290), .B(n50541), .X(n32832) );
  nand_x1_sg U64087 ( .A(n57290), .B(n50539), .X(n32870) );
  nand_x1_sg U64088 ( .A(n57290), .B(n53089), .X(n32860) );
  nand_x1_sg U64089 ( .A(n57290), .B(n50537), .X(n32872) );
  nand_x1_sg U64090 ( .A(n57286), .B(n50865), .X(n32886) );
  nand_x1_sg U64091 ( .A(n57286), .B(n50857), .X(n32894) );
  nand_x1_sg U64092 ( .A(n57286), .B(n50853), .X(n32896) );
  nand_x1_sg U64093 ( .A(n57286), .B(n50847), .X(n32912) );
  nand_x1_sg U64094 ( .A(n57286), .B(n53429), .X(n32914) );
  nand_x1_sg U64095 ( .A(n57286), .B(n50839), .X(n32904) );
  nand_x1_sg U64096 ( .A(n57290), .B(n50565), .X(n32840) );
  nand_x1_sg U64097 ( .A(n57290), .B(n53093), .X(n32850) );
  nand_x1_sg U64098 ( .A(n57290), .B(n50557), .X(n32848) );
  nand_x1_sg U64099 ( .A(n57290), .B(n50545), .X(n32866) );
  nand_x1_sg U64100 ( .A(n57290), .B(n50543), .X(n32858) );
  nand_x1_sg U64101 ( .A(n57290), .B(n53091), .X(n32868) );
  nand_x4_sg U64102 ( .A(n57091), .B(n57308), .X(n26052) );
  nand_x1_sg U64103 ( .A(n47409), .B(n30627), .X(n40227) );
  nand_x1_sg U64104 ( .A(n50561), .B(n57876), .X(n29734) );
  nand_x1_sg U64105 ( .A(n57089), .B(n46207), .X(n29735) );
  nand_x1_sg U64106 ( .A(n50559), .B(n57880), .X(n29732) );
  nand_x1_sg U64107 ( .A(n57087), .B(n57892), .X(n29733) );
  nand_x1_sg U64108 ( .A(n53093), .B(n57878), .X(n29740) );
  nand_x1_sg U64109 ( .A(n51553), .B(n57911), .X(n29741) );
  nand_x1_sg U64110 ( .A(n50553), .B(n57878), .X(n29720) );
  nand_x1_sg U64111 ( .A(n57079), .B(n57896), .X(n29721) );
  nand_x1_sg U64112 ( .A(n50547), .B(n57875), .X(n29758) );
  nand_x1_sg U64113 ( .A(n57071), .B(n57896), .X(n29759) );
  nand_x1_sg U64114 ( .A(n53091), .B(n57876), .X(n29762) );
  nand_x1_sg U64115 ( .A(n51545), .B(n46207), .X(n29763) );
  nand_x1_sg U64116 ( .A(n53089), .B(n57877), .X(n29752) );
  nand_x1_sg U64117 ( .A(n47773), .B(n46207), .X(n29753) );
  nand_x1_sg U64118 ( .A(n53435), .B(n57878), .X(n30256) );
  nand_x1_sg U64119 ( .A(n51543), .B(n46207), .X(n30257) );
  nand_x1_sg U64120 ( .A(n53433), .B(n57876), .X(n30352) );
  nand_x1_sg U64121 ( .A(n47759), .B(n57895), .X(n30353) );
  nand_x1_sg U64122 ( .A(n53431), .B(n57882), .X(n30178) );
  nand_x1_sg U64123 ( .A(n51551), .B(n46207), .X(n30179) );
  nand_x1_sg U64124 ( .A(n50855), .B(n57878), .X(n30430) );
  nand_x1_sg U64125 ( .A(n57077), .B(n57910), .X(n30431) );
  nand_x1_sg U64126 ( .A(n50849), .B(n57876), .X(n30334) );
  nand_x1_sg U64127 ( .A(n57075), .B(n57895), .X(n30335) );
  nand_x1_sg U64128 ( .A(n50839), .B(n46213), .X(n30502) );
  nand_x1_sg U64129 ( .A(n57073), .B(n57891), .X(n30503) );
  nand_x1_sg U64130 ( .A(n47355), .B(n61911), .X(n57953) );
  nand_x2_sg U64131 ( .A(output_taken), .B(n61906), .X(n57954) );
  nand_x1_sg U64132 ( .A(n50593), .B(n46210), .X(n29842) );
  nand_x1_sg U64133 ( .A(n57063), .B(n57902), .X(n29843) );
  nand_x1_sg U64134 ( .A(n50587), .B(n46209), .X(n29846) );
  nand_x1_sg U64135 ( .A(n57067), .B(n57897), .X(n29847) );
  nand_x1_sg U64136 ( .A(n50585), .B(n57875), .X(n29782) );
  nand_x1_sg U64137 ( .A(n57061), .B(n57886), .X(n29783) );
  nand_x1_sg U64138 ( .A(n53109), .B(n46212), .X(n29780) );
  nand_x1_sg U64139 ( .A(n51541), .B(n57887), .X(n29781) );
  nand_x1_sg U64140 ( .A(n50579), .B(n46213), .X(n29770) );
  nand_x1_sg U64141 ( .A(n57059), .B(n57910), .X(n29771) );
  nand_x1_sg U64142 ( .A(n53107), .B(n57877), .X(n29768) );
  nand_x1_sg U64143 ( .A(n51539), .B(n57907), .X(n29769) );
  nand_x1_sg U64144 ( .A(n50573), .B(n46210), .X(n29806) );
  nand_x1_sg U64145 ( .A(n57057), .B(n57898), .X(n29807) );
  nand_x1_sg U64146 ( .A(n53105), .B(n57880), .X(n29804) );
  nand_x1_sg U64147 ( .A(n51537), .B(n57907), .X(n29805) );
  nand_x1_sg U64148 ( .A(n53103), .B(n46209), .X(n29812) );
  nand_x1_sg U64149 ( .A(n47771), .B(n57896), .X(n29813) );
  nand_x1_sg U64150 ( .A(n53101), .B(n57875), .X(n29792) );
  nand_x1_sg U64151 ( .A(n51535), .B(n57895), .X(n29793) );
  nand_x1_sg U64152 ( .A(n53099), .B(n57875), .X(n29800) );
  nand_x1_sg U64153 ( .A(n47769), .B(n57900), .X(n29801) );
  nand_x1_sg U64154 ( .A(n53097), .B(n57880), .X(n29798) );
  nand_x1_sg U64155 ( .A(n47767), .B(n57900), .X(n29799) );
  nand_x1_sg U64156 ( .A(n50893), .B(n57880), .X(n30404) );
  nand_x1_sg U64157 ( .A(n57055), .B(n57887), .X(n30405) );
  nand_x1_sg U64158 ( .A(n50887), .B(n46212), .X(n30408) );
  nand_x1_sg U64159 ( .A(n57065), .B(n57899), .X(n30409) );
  nand_x1_sg U64160 ( .A(n50885), .B(n57875), .X(n30344) );
  nand_x1_sg U64161 ( .A(n57053), .B(n57900), .X(n30345) );
  nand_x1_sg U64162 ( .A(n53449), .B(n57875), .X(n30342) );
  nand_x1_sg U64163 ( .A(n51533), .B(n57896), .X(n30343) );
  nand_x1_sg U64164 ( .A(n50879), .B(n57875), .X(n30332) );
  nand_x1_sg U64165 ( .A(n57051), .B(n57910), .X(n30333) );
  nand_x1_sg U64166 ( .A(n53447), .B(n57880), .X(n30330) );
  nand_x1_sg U64167 ( .A(n51531), .B(n57908), .X(n30331) );
  nand_x1_sg U64168 ( .A(n50873), .B(n57878), .X(n30368) );
  nand_x1_sg U64169 ( .A(n57049), .B(n57900), .X(n30369) );
  nand_x1_sg U64170 ( .A(n53445), .B(n57878), .X(n30366) );
  nand_x1_sg U64171 ( .A(n51529), .B(n57915), .X(n30367) );
  nand_x1_sg U64172 ( .A(n53443), .B(n46213), .X(n30374) );
  nand_x1_sg U64173 ( .A(n47765), .B(n46207), .X(n30375) );
  nand_x1_sg U64174 ( .A(n53441), .B(n57878), .X(n30354) );
  nand_x1_sg U64175 ( .A(n51527), .B(n57907), .X(n30355) );
  nand_x1_sg U64176 ( .A(n53439), .B(n57876), .X(n30362) );
  nand_x1_sg U64177 ( .A(n47763), .B(n57896), .X(n30363) );
  nand_x1_sg U64178 ( .A(n53437), .B(n46213), .X(n30360) );
  nand_x1_sg U64179 ( .A(n47761), .B(n57900), .X(n30361) );
  nand_x1_sg U64180 ( .A(n50447), .B(n57878), .X(n30084) );
  nand_x1_sg U64181 ( .A(n57029), .B(n57898), .X(n30085) );
  nand_x1_sg U64182 ( .A(n50445), .B(n57878), .X(n30082) );
  nand_x1_sg U64183 ( .A(n57043), .B(n57911), .X(n30083) );
  nand_x1_sg U64184 ( .A(n52935), .B(n57880), .X(n30090) );
  nand_x1_sg U64185 ( .A(n51519), .B(n57898), .X(n30091) );
  nand_x1_sg U64186 ( .A(n50443), .B(n57875), .X(n30088) );
  nand_x1_sg U64187 ( .A(n57027), .B(n57899), .X(n30089) );
  nand_x1_sg U64188 ( .A(n52933), .B(n46213), .X(n30072) );
  nand_x1_sg U64189 ( .A(n51505), .B(n57897), .X(n30073) );
  nand_x1_sg U64190 ( .A(n52931), .B(n57878), .X(n30070) );
  nand_x1_sg U64191 ( .A(n47757), .B(n57895), .X(n30071) );
  nand_x1_sg U64192 ( .A(n50441), .B(n57880), .X(n30078) );
  nand_x1_sg U64193 ( .A(n57041), .B(n57900), .X(n30079) );
  nand_x1_sg U64194 ( .A(n52929), .B(n57878), .X(n30076) );
  nand_x1_sg U64195 ( .A(n51517), .B(n57907), .X(n30077) );
  nand_x1_sg U64196 ( .A(n50439), .B(n46209), .X(n29830) );
  nand_x1_sg U64197 ( .A(n57021), .B(n57900), .X(n29831) );
  nand_x1_sg U64198 ( .A(n52927), .B(n46210), .X(n29828) );
  nand_x1_sg U64199 ( .A(n51503), .B(n57908), .X(n29829) );
  nand_x1_sg U64200 ( .A(n50437), .B(n46210), .X(n29836) );
  nand_x1_sg U64201 ( .A(n57039), .B(n57886), .X(n29837) );
  nand_x1_sg U64202 ( .A(n52925), .B(n57880), .X(n29834) );
  nand_x1_sg U64203 ( .A(n51515), .B(n57887), .X(n29835) );
  nand_x1_sg U64204 ( .A(n50435), .B(n46210), .X(n29818) );
  nand_x1_sg U64205 ( .A(n57013), .B(n57899), .X(n29819) );
  nand_x1_sg U64206 ( .A(n52923), .B(n57875), .X(n29816) );
  nand_x1_sg U64207 ( .A(n51491), .B(n57908), .X(n29817) );
  nand_x1_sg U64208 ( .A(n52921), .B(n46209), .X(n29824) );
  nand_x1_sg U64209 ( .A(n47747), .B(n57909), .X(n29825) );
  nand_x1_sg U64210 ( .A(n50433), .B(n46209), .X(n29822) );
  nand_x1_sg U64211 ( .A(n57015), .B(n57909), .X(n29823) );
  nand_x1_sg U64212 ( .A(n52919), .B(n46210), .X(n29854) );
  nand_x1_sg U64213 ( .A(n51493), .B(n57887), .X(n29855) );
  nand_x1_sg U64214 ( .A(n52917), .B(n46209), .X(n29852) );
  nand_x1_sg U64215 ( .A(n51489), .B(n57911), .X(n29853) );
  nand_x1_sg U64216 ( .A(n52915), .B(n57876), .X(n29860) );
  nand_x1_sg U64217 ( .A(n47745), .B(n57898), .X(n29861) );
  nand_x1_sg U64218 ( .A(n52913), .B(n57880), .X(n29858) );
  nand_x1_sg U64219 ( .A(n47743), .B(n57898), .X(n29859) );
  nand_x1_sg U64220 ( .A(n53275), .B(n46210), .X(n29844) );
  nand_x1_sg U64221 ( .A(n51513), .B(n57899), .X(n29845) );
  nand_x1_sg U64222 ( .A(n50739), .B(n46212), .X(n30392) );
  nand_x1_sg U64223 ( .A(n57019), .B(n57911), .X(n30393) );
  nand_x1_sg U64224 ( .A(n53267), .B(n57878), .X(n30390) );
  nand_x1_sg U64225 ( .A(n51499), .B(n57902), .X(n30391) );
  nand_x1_sg U64226 ( .A(n50737), .B(n57875), .X(n30398) );
  nand_x1_sg U64227 ( .A(n57033), .B(n57901), .X(n30399) );
  nand_x1_sg U64228 ( .A(n53265), .B(n57876), .X(n30396) );
  nand_x1_sg U64229 ( .A(n51509), .B(n57898), .X(n30397) );
  nand_x1_sg U64230 ( .A(n50735), .B(n46213), .X(n30380) );
  nand_x1_sg U64231 ( .A(n57017), .B(n57895), .X(n30381) );
  nand_x1_sg U64232 ( .A(n53263), .B(n57877), .X(n30378) );
  nand_x1_sg U64233 ( .A(n51497), .B(n57907), .X(n30379) );
  nand_x1_sg U64234 ( .A(n53261), .B(n57877), .X(n30386) );
  nand_x1_sg U64235 ( .A(n47753), .B(n57902), .X(n30387) );
  nand_x1_sg U64236 ( .A(n50733), .B(n57878), .X(n30384) );
  nand_x1_sg U64237 ( .A(n57031), .B(n57911), .X(n30385) );
  nand_x1_sg U64238 ( .A(n53259), .B(n57878), .X(n30416) );
  nand_x1_sg U64239 ( .A(n51507), .B(n57911), .X(n30417) );
  nand_x1_sg U64240 ( .A(n53257), .B(n57876), .X(n30414) );
  nand_x1_sg U64241 ( .A(n51495), .B(n57886), .X(n30415) );
  nand_x1_sg U64242 ( .A(n53255), .B(n57880), .X(n30422) );
  nand_x1_sg U64243 ( .A(n47751), .B(n57911), .X(n30423) );
  nand_x1_sg U64244 ( .A(n53253), .B(n57876), .X(n30420) );
  nand_x1_sg U64245 ( .A(n47749), .B(n57903), .X(n30421) );
  nand_x1_sg U64246 ( .A(n50591), .B(n46209), .X(n29840) );
  nand_x1_sg U64247 ( .A(n56967), .B(n57900), .X(n29841) );
  nand_x1_sg U64248 ( .A(n50589), .B(n46210), .X(n29848) );
  nand_x1_sg U64249 ( .A(n56965), .B(n57895), .X(n29849) );
  nand_x1_sg U64250 ( .A(n50583), .B(n57880), .X(n29788) );
  nand_x1_sg U64251 ( .A(n56963), .B(n46207), .X(n29789) );
  nand_x1_sg U64252 ( .A(n50581), .B(n46212), .X(n29786) );
  nand_x1_sg U64253 ( .A(n56961), .B(n57907), .X(n29787) );
  nand_x1_sg U64254 ( .A(n50577), .B(n57878), .X(n29776) );
  nand_x1_sg U64255 ( .A(n56959), .B(n57908), .X(n29777) );
  nand_x1_sg U64256 ( .A(n50575), .B(n46212), .X(n29774) );
  nand_x1_sg U64257 ( .A(n56957), .B(n57898), .X(n29775) );
  nand_x1_sg U64258 ( .A(n50571), .B(n57877), .X(n29810) );
  nand_x1_sg U64259 ( .A(n56955), .B(n57886), .X(n29811) );
  nand_x1_sg U64260 ( .A(n50569), .B(n57876), .X(n29794) );
  nand_x1_sg U64261 ( .A(n56953), .B(n57907), .X(n29795) );
  nand_x1_sg U64262 ( .A(n50891), .B(n57878), .X(n30402) );
  nand_x1_sg U64263 ( .A(n56951), .B(n57899), .X(n30403) );
  nand_x1_sg U64264 ( .A(n50889), .B(n46212), .X(n30410) );
  nand_x1_sg U64265 ( .A(n56949), .B(n57898), .X(n30411) );
  nand_x1_sg U64266 ( .A(n50883), .B(n57880), .X(n30350) );
  nand_x1_sg U64267 ( .A(n56947), .B(n57899), .X(n30351) );
  nand_x1_sg U64268 ( .A(n50881), .B(n57877), .X(n30348) );
  nand_x1_sg U64269 ( .A(n56945), .B(n57895), .X(n30349) );
  nand_x1_sg U64270 ( .A(n50877), .B(n57880), .X(n30338) );
  nand_x1_sg U64271 ( .A(n56943), .B(n57896), .X(n30339) );
  nand_x1_sg U64272 ( .A(n50875), .B(n57872), .X(n30336) );
  nand_x1_sg U64273 ( .A(n56941), .B(n57896), .X(n30337) );
  nand_x1_sg U64274 ( .A(n50871), .B(n57875), .X(n30372) );
  nand_x1_sg U64275 ( .A(n56939), .B(n57909), .X(n30373) );
  nand_x1_sg U64276 ( .A(n50869), .B(n57875), .X(n30356) );
  nand_x1_sg U64277 ( .A(n56937), .B(n57910), .X(n30357) );
  nand_x1_sg U64278 ( .A(n50565), .B(n57872), .X(n30552) );
  nand_x1_sg U64279 ( .A(n56995), .B(n57908), .X(n30553) );
  nand_x1_sg U64280 ( .A(n50557), .B(n57877), .X(n29738) );
  nand_x1_sg U64281 ( .A(n57003), .B(n57900), .X(n29739) );
  nand_x1_sg U64282 ( .A(n50555), .B(n57878), .X(n29722) );
  nand_x1_sg U64283 ( .A(n57001), .B(n57896), .X(n29723) );
  nand_x1_sg U64284 ( .A(n50551), .B(n57882), .X(n29728) );
  nand_x1_sg U64285 ( .A(n57011), .B(n57886), .X(n29729) );
  nand_x1_sg U64286 ( .A(n50549), .B(n57877), .X(n29726) );
  nand_x1_sg U64287 ( .A(n57009), .B(n57895), .X(n29727) );
  nand_x1_sg U64288 ( .A(n50545), .B(n57876), .X(n29756) );
  nand_x1_sg U64289 ( .A(n56981), .B(n57908), .X(n29757) );
  nand_x1_sg U64290 ( .A(n50543), .B(n57876), .X(n29764) );
  nand_x1_sg U64291 ( .A(n56979), .B(n46207), .X(n29765) );
  nand_x1_sg U64292 ( .A(n50541), .B(n57877), .X(n29746) );
  nand_x1_sg U64293 ( .A(n56985), .B(n57907), .X(n29747) );
  nand_x1_sg U64294 ( .A(n50539), .B(n57880), .X(n29744) );
  nand_x1_sg U64295 ( .A(n56983), .B(n57908), .X(n29745) );
  nand_x1_sg U64296 ( .A(n50537), .B(n46213), .X(n29750) );
  nand_x1_sg U64297 ( .A(n57045), .B(n46207), .X(n29751) );
  nand_x1_sg U64298 ( .A(n50867), .B(n57880), .X(n30232) );
  nand_x1_sg U64299 ( .A(n56975), .B(n57910), .X(n30233) );
  nand_x1_sg U64300 ( .A(n50865), .B(n57876), .X(n30496) );
  nand_x1_sg U64301 ( .A(n56973), .B(n57891), .X(n30497) );
  nand_x1_sg U64302 ( .A(n50859), .B(n46209), .X(n30166) );
  nand_x1_sg U64303 ( .A(n56977), .B(n57911), .X(n30167) );
  nand_x1_sg U64304 ( .A(n50857), .B(n57878), .X(n30448) );
  nand_x1_sg U64305 ( .A(n56999), .B(n57894), .X(n30449) );
  nand_x1_sg U64306 ( .A(n50853), .B(n46213), .X(n30418) );
  nand_x1_sg U64307 ( .A(n57007), .B(n57901), .X(n30419) );
  nand_x1_sg U64308 ( .A(n50851), .B(n46213), .X(n30412) );
  nand_x1_sg U64309 ( .A(n57005), .B(n57886), .X(n30413) );
  nand_x1_sg U64310 ( .A(n50847), .B(n57878), .X(n30514) );
  nand_x1_sg U64311 ( .A(n56993), .B(n57890), .X(n30515) );
  nand_x1_sg U64312 ( .A(n50845), .B(n46213), .X(n30436) );
  nand_x1_sg U64313 ( .A(n56991), .B(n57897), .X(n30437) );
  nand_x1_sg U64314 ( .A(n50843), .B(n57878), .X(n30478) );
  nand_x1_sg U64315 ( .A(n56989), .B(n57893), .X(n30479) );
  nand_x1_sg U64316 ( .A(n50841), .B(n57877), .X(n30388) );
  nand_x1_sg U64317 ( .A(n56987), .B(n57901), .X(n30389) );
  nand_x1_sg U64318 ( .A(n50837), .B(n46210), .X(n30160) );
  nand_x1_sg U64319 ( .A(n57047), .B(n57910), .X(n30161) );
  nand_x1_sg U64320 ( .A(n53041), .B(n57877), .X(n29684) );
  nand_x1_sg U64321 ( .A(n47647), .B(n57908), .X(n29685) );
  nand_x1_sg U64322 ( .A(n50513), .B(n46213), .X(n29682) );
  nand_x1_sg U64323 ( .A(n56733), .B(n57909), .X(n29683) );
  nand_x1_sg U64324 ( .A(n50511), .B(n57875), .X(n29702) );
  nand_x1_sg U64325 ( .A(n56689), .B(n57887), .X(n29703) );
  nand_x1_sg U64326 ( .A(n50509), .B(n57878), .X(n29700) );
  nand_x1_sg U64327 ( .A(n56843), .B(n57910), .X(n29701) );
  nand_x1_sg U64328 ( .A(n53031), .B(n46212), .X(n29708) );
  nand_x1_sg U64329 ( .A(n51403), .B(n46207), .X(n29709) );
  nand_x1_sg U64330 ( .A(n53029), .B(n46212), .X(n29706) );
  nand_x1_sg U64331 ( .A(n47691), .B(n57898), .X(n29707) );
  nand_x1_sg U64332 ( .A(n50507), .B(n57875), .X(n29690) );
  nand_x1_sg U64333 ( .A(n56703), .B(n57907), .X(n29691) );
  nand_x1_sg U64334 ( .A(n53027), .B(n57880), .X(n29688) );
  nand_x1_sg U64335 ( .A(n51241), .B(n57910), .X(n29689) );
  nand_x1_sg U64336 ( .A(n50505), .B(n57875), .X(n29696) );
  nand_x1_sg U64337 ( .A(n56731), .B(n57887), .X(n29697) );
  nand_x1_sg U64338 ( .A(n53025), .B(n57880), .X(n29694) );
  nand_x1_sg U64339 ( .A(n51269), .B(n57910), .X(n29695) );
  nand_x1_sg U64340 ( .A(n50491), .B(n57873), .X(n30012) );
  nand_x1_sg U64341 ( .A(n56773), .B(n57902), .X(n30013) );
  nand_x1_sg U64342 ( .A(n53003), .B(n57872), .X(n30010) );
  nand_x1_sg U64343 ( .A(n51315), .B(n57904), .X(n30011) );
  nand_x1_sg U64344 ( .A(n50489), .B(n57873), .X(n30018) );
  nand_x1_sg U64345 ( .A(n56821), .B(n57901), .X(n30019) );
  nand_x1_sg U64346 ( .A(n53001), .B(n57873), .X(n30016) );
  nand_x1_sg U64347 ( .A(n51375), .B(n57887), .X(n30017) );
  nand_x1_sg U64348 ( .A(n50487), .B(n57872), .X(n30000) );
  nand_x1_sg U64349 ( .A(n56771), .B(n57900), .X(n30001) );
  nand_x1_sg U64350 ( .A(n52999), .B(n57872), .X(n29998) );
  nand_x1_sg U64351 ( .A(n51313), .B(n57887), .X(n29999) );
  nand_x1_sg U64352 ( .A(n50485), .B(n57872), .X(n30006) );
  nand_x1_sg U64353 ( .A(n56819), .B(n57895), .X(n30007) );
  nand_x1_sg U64354 ( .A(n52997), .B(n57872), .X(n30004) );
  nand_x1_sg U64355 ( .A(n51373), .B(n57896), .X(n30005) );
  nand_x1_sg U64356 ( .A(n50483), .B(n57878), .X(n30036) );
  nand_x1_sg U64357 ( .A(n56683), .B(n57910), .X(n30037) );
  nand_x1_sg U64358 ( .A(n52995), .B(n46213), .X(n30034) );
  nand_x1_sg U64359 ( .A(n51221), .B(n57910), .X(n30035) );
  nand_x1_sg U64360 ( .A(n52993), .B(n57878), .X(n30042) );
  nand_x1_sg U64361 ( .A(n47635), .B(n57908), .X(n30043) );
  nand_x1_sg U64362 ( .A(n50481), .B(n46212), .X(n30040) );
  nand_x1_sg U64363 ( .A(n56725), .B(n57902), .X(n30041) );
  nand_x1_sg U64364 ( .A(n52991), .B(n57873), .X(n30024) );
  nand_x1_sg U64365 ( .A(n51263), .B(n57907), .X(n30025) );
  nand_x1_sg U64366 ( .A(n52989), .B(n57873), .X(n30022) );
  nand_x1_sg U64367 ( .A(n51219), .B(n57886), .X(n30023) );
  nand_x1_sg U64368 ( .A(n52987), .B(n46210), .X(n30030) );
  nand_x1_sg U64369 ( .A(n47633), .B(n57896), .X(n30031) );
  nand_x1_sg U64370 ( .A(n52985), .B(n57873), .X(n30028) );
  nand_x1_sg U64371 ( .A(n47631), .B(n57899), .X(n30029) );
  nand_x1_sg U64372 ( .A(n52983), .B(n57880), .X(n29974) );
  nand_x1_sg U64373 ( .A(n51327), .B(n57910), .X(n29975) );
  nand_x1_sg U64374 ( .A(n52981), .B(n57880), .X(n29972) );
  nand_x1_sg U64375 ( .A(n47703), .B(n57908), .X(n29973) );
  nand_x1_sg U64376 ( .A(n50479), .B(n57876), .X(n29980) );
  nand_x1_sg U64377 ( .A(n56857), .B(n57910), .X(n29981) );
  nand_x1_sg U64378 ( .A(n52979), .B(n57877), .X(n29978) );
  nand_x1_sg U64379 ( .A(n51421), .B(n57896), .X(n29979) );
  nand_x1_sg U64380 ( .A(n50477), .B(n57876), .X(n29962) );
  nand_x1_sg U64381 ( .A(n56769), .B(n57887), .X(n29963) );
  nand_x1_sg U64382 ( .A(n52977), .B(n57877), .X(n29960) );
  nand_x1_sg U64383 ( .A(n51311), .B(n57911), .X(n29961) );
  nand_x1_sg U64384 ( .A(n52975), .B(n57875), .X(n29968) );
  nand_x1_sg U64385 ( .A(n51371), .B(n57907), .X(n29969) );
  nand_x1_sg U64386 ( .A(n50475), .B(n57875), .X(n29966) );
  nand_x1_sg U64387 ( .A(n56817), .B(n57910), .X(n29967) );
  nand_x1_sg U64388 ( .A(n52973), .B(n57877), .X(n29964) );
  nand_x1_sg U64389 ( .A(n51309), .B(n57887), .X(n29965) );
  nand_x1_sg U64390 ( .A(n50473), .B(n46212), .X(n29716) );
  nand_x1_sg U64391 ( .A(n56767), .B(n46207), .X(n29717) );
  nand_x1_sg U64392 ( .A(n52971), .B(n57873), .X(n30014) );
  nand_x1_sg U64393 ( .A(n51369), .B(n57886), .X(n30015) );
  nand_x1_sg U64394 ( .A(n50471), .B(n57872), .X(n30002) );
  nand_x1_sg U64395 ( .A(n56815), .B(n57907), .X(n30003) );
  nand_x1_sg U64396 ( .A(n52969), .B(n57871), .X(n29988) );
  nand_x1_sg U64397 ( .A(n51217), .B(n46207), .X(n29989) );
  nand_x1_sg U64398 ( .A(n50469), .B(n57871), .X(n29986) );
  nand_x1_sg U64399 ( .A(n56681), .B(n57896), .X(n29987) );
  nand_x1_sg U64400 ( .A(n52967), .B(n57872), .X(n29994) );
  nand_x1_sg U64401 ( .A(n47531), .B(n57895), .X(n29995) );
  nand_x1_sg U64402 ( .A(n52965), .B(n57871), .X(n29992) );
  nand_x1_sg U64403 ( .A(n51261), .B(n57900), .X(n29993) );
  nand_x1_sg U64404 ( .A(n50467), .B(n46209), .X(n30108) );
  nand_x1_sg U64405 ( .A(n56723), .B(n57897), .X(n30109) );
  nand_x1_sg U64406 ( .A(n50465), .B(n46210), .X(n30106) );
  nand_x1_sg U64407 ( .A(n56679), .B(n57897), .X(n30107) );
  nand_x1_sg U64408 ( .A(n52963), .B(n46209), .X(n30114) );
  nand_x1_sg U64409 ( .A(n47529), .B(n57910), .X(n30115) );
  nand_x1_sg U64410 ( .A(n52961), .B(n46210), .X(n30112) );
  nand_x1_sg U64411 ( .A(n47527), .B(n57908), .X(n30113) );
  nand_x1_sg U64412 ( .A(n52959), .B(n57880), .X(n30096) );
  nand_x1_sg U64413 ( .A(n51325), .B(n57897), .X(n30097) );
  nand_x1_sg U64414 ( .A(n50463), .B(n57880), .X(n30094) );
  nand_x1_sg U64415 ( .A(n56855), .B(n57886), .X(n30095) );
  nand_x1_sg U64416 ( .A(n52957), .B(n46209), .X(n30102) );
  nand_x1_sg U64417 ( .A(n47555), .B(n57897), .X(n30103) );
  nand_x1_sg U64418 ( .A(n52955), .B(n57875), .X(n30100) );
  nand_x1_sg U64419 ( .A(n51419), .B(n57897), .X(n30101) );
  nand_x1_sg U64420 ( .A(n52953), .B(n46209), .X(n30132) );
  nand_x1_sg U64421 ( .A(n51307), .B(n57900), .X(n30133) );
  nand_x1_sg U64422 ( .A(n50461), .B(n46210), .X(n30130) );
  nand_x1_sg U64423 ( .A(n56765), .B(n57908), .X(n30131) );
  nand_x1_sg U64424 ( .A(n52951), .B(n57873), .X(n30074) );
  nand_x1_sg U64425 ( .A(n51367), .B(n57886), .X(n30075) );
  nand_x1_sg U64426 ( .A(n50459), .B(n46209), .X(n30122) );
  nand_x1_sg U64427 ( .A(n56813), .B(n57909), .X(n30123) );
  nand_x1_sg U64428 ( .A(n52949), .B(n46210), .X(n30120) );
  nand_x1_sg U64429 ( .A(n51305), .B(n57899), .X(n30121) );
  nand_x1_sg U64430 ( .A(n50457), .B(n46210), .X(n30118) );
  nand_x1_sg U64431 ( .A(n56763), .B(n57904), .X(n30119) );
  nand_x1_sg U64432 ( .A(n52947), .B(n46209), .X(n30126) );
  nand_x1_sg U64433 ( .A(n51365), .B(n57897), .X(n30127) );
  nand_x1_sg U64434 ( .A(n50455), .B(n46210), .X(n30124) );
  nand_x1_sg U64435 ( .A(n56811), .B(n57901), .X(n30125) );
  nand_x1_sg U64436 ( .A(n52945), .B(n46209), .X(n30060) );
  nand_x1_sg U64437 ( .A(n51215), .B(n57908), .X(n30061) );
  nand_x1_sg U64438 ( .A(n50453), .B(n46210), .X(n30058) );
  nand_x1_sg U64439 ( .A(n56677), .B(n57907), .X(n30059) );
  nand_x1_sg U64440 ( .A(n52943), .B(n57877), .X(n30066) );
  nand_x1_sg U64441 ( .A(n47525), .B(n57888), .X(n30067) );
  nand_x1_sg U64442 ( .A(n52941), .B(n46209), .X(n30064) );
  nand_x1_sg U64443 ( .A(n51259), .B(n57898), .X(n30065) );
  nand_x1_sg U64444 ( .A(n50451), .B(n46210), .X(n30048) );
  nand_x1_sg U64445 ( .A(n56721), .B(n57888), .X(n30049) );
  nand_x1_sg U64446 ( .A(n50449), .B(n57878), .X(n30046) );
  nand_x1_sg U64447 ( .A(n56675), .B(n57897), .X(n30047) );
  nand_x1_sg U64448 ( .A(n52939), .B(n46209), .X(n30054) );
  nand_x1_sg U64449 ( .A(n47523), .B(n57903), .X(n30055) );
  nand_x1_sg U64450 ( .A(n52937), .B(n46210), .X(n30052) );
  nand_x1_sg U64451 ( .A(n47521), .B(n57910), .X(n30053) );
  nand_x1_sg U64452 ( .A(n50617), .B(n57875), .X(n29866) );
  nand_x1_sg U64453 ( .A(n56849), .B(n57898), .X(n29867) );
  nand_x1_sg U64454 ( .A(n53165), .B(n57877), .X(n29864) );
  nand_x1_sg U64455 ( .A(n51409), .B(n57898), .X(n29865) );
  nand_x1_sg U64456 ( .A(n53163), .B(n57880), .X(n29872) );
  nand_x1_sg U64457 ( .A(n47697), .B(n46207), .X(n29873) );
  nand_x1_sg U64458 ( .A(n50615), .B(n57878), .X(n29870) );
  nand_x1_sg U64459 ( .A(n56867), .B(n57898), .X(n29871) );
  nand_x1_sg U64460 ( .A(n50613), .B(n57878), .X(n29902) );
  nand_x1_sg U64461 ( .A(n56841), .B(n57910), .X(n29903) );
  nand_x1_sg U64462 ( .A(n53161), .B(n46213), .X(n29900) );
  nand_x1_sg U64463 ( .A(n51401), .B(n57908), .X(n29901) );
  nand_x1_sg U64464 ( .A(n50611), .B(n57878), .X(n29908) );
  nand_x1_sg U64465 ( .A(n56789), .B(n46207), .X(n29909) );
  nand_x1_sg U64466 ( .A(n53159), .B(n46210), .X(n29906) );
  nand_x1_sg U64467 ( .A(n51341), .B(n46207), .X(n29907) );
  nand_x1_sg U64468 ( .A(n50609), .B(n57878), .X(n29890) );
  nand_x1_sg U64469 ( .A(n56839), .B(n57909), .X(n29891) );
  nand_x1_sg U64470 ( .A(n53157), .B(n46209), .X(n29888) );
  nand_x1_sg U64471 ( .A(n51399), .B(n46207), .X(n29889) );
  nand_x1_sg U64472 ( .A(n50607), .B(n46212), .X(n29896) );
  nand_x1_sg U64473 ( .A(n56787), .B(n57898), .X(n29897) );
  nand_x1_sg U64474 ( .A(n53155), .B(n57878), .X(n29894) );
  nand_x1_sg U64475 ( .A(n51339), .B(n57911), .X(n29895) );
  nand_x1_sg U64476 ( .A(n53151), .B(n57878), .X(n30316) );
  nand_x1_sg U64477 ( .A(n47689), .B(n57911), .X(n30317) );
  nand_x1_sg U64478 ( .A(n50603), .B(n57870), .X(n30328) );
  nand_x1_sg U64479 ( .A(n56785), .B(n57909), .X(n30329) );
  nand_x1_sg U64480 ( .A(n53149), .B(n57875), .X(n30310) );
  nand_x1_sg U64481 ( .A(n51337), .B(n57904), .X(n30311) );
  nand_x1_sg U64482 ( .A(n53147), .B(n57882), .X(n30298) );
  nand_x1_sg U64483 ( .A(n51395), .B(n57900), .X(n30299) );
  nand_x1_sg U64484 ( .A(n53145), .B(n57880), .X(n30286) );
  nand_x1_sg U64485 ( .A(n47687), .B(n57908), .X(n30287) );
  nand_x1_sg U64486 ( .A(n53143), .B(n57880), .X(n30280) );
  nand_x1_sg U64487 ( .A(n47685), .B(n46207), .X(n30281) );
  nand_x1_sg U64488 ( .A(n50827), .B(n57878), .X(n29970) );
  nand_x1_sg U64489 ( .A(n56671), .B(n57886), .X(n29971) );
  nand_x1_sg U64490 ( .A(n50825), .B(n57878), .X(n29976) );
  nand_x1_sg U64491 ( .A(n56833), .B(n57896), .X(n29977) );
  nand_x1_sg U64492 ( .A(n53395), .B(n57875), .X(n29916) );
  nand_x1_sg U64493 ( .A(n51391), .B(n57909), .X(n29917) );
  nand_x1_sg U64494 ( .A(n53393), .B(n46209), .X(n30128) );
  nand_x1_sg U64495 ( .A(n47681), .B(n46207), .X(n30129) );
  nand_x1_sg U64496 ( .A(n50823), .B(n46212), .X(n30062) );
  nand_x1_sg U64497 ( .A(n56701), .B(n57888), .X(n30063) );
  nand_x1_sg U64498 ( .A(n53391), .B(n46209), .X(n30056) );
  nand_x1_sg U64499 ( .A(n51239), .B(n57903), .X(n30057) );
  nand_x1_sg U64500 ( .A(n50819), .B(n46210), .X(n30092) );
  nand_x1_sg U64501 ( .A(n56669), .B(n57887), .X(n30093) );
  nand_x1_sg U64502 ( .A(n53387), .B(n46209), .X(n30104) );
  nand_x1_sg U64503 ( .A(n51211), .B(n57897), .X(n30105) );
  nand_x1_sg U64504 ( .A(n50817), .B(n46209), .X(n30086) );
  nand_x1_sg U64505 ( .A(n56715), .B(n57887), .X(n30087) );
  nand_x1_sg U64506 ( .A(n53385), .B(n57877), .X(n30080) );
  nand_x1_sg U64507 ( .A(n51253), .B(n57897), .X(n30081) );
  nand_x1_sg U64508 ( .A(n50809), .B(n57875), .X(n29928) );
  nand_x1_sg U64509 ( .A(n56831), .B(n57909), .X(n29929) );
  nand_x1_sg U64510 ( .A(n53371), .B(n57875), .X(n29922) );
  nand_x1_sg U64511 ( .A(n51389), .B(n57898), .X(n29923) );
  nand_x1_sg U64512 ( .A(n50807), .B(n57875), .X(n29934) );
  nand_x1_sg U64513 ( .A(n56699), .B(n57911), .X(n29935) );
  nand_x1_sg U64514 ( .A(n50805), .B(n57875), .X(n29946) );
  nand_x1_sg U64515 ( .A(n56711), .B(n57897), .X(n29947) );
  nand_x1_sg U64516 ( .A(n53365), .B(n57877), .X(n29952) );
  nand_x1_sg U64517 ( .A(n51249), .B(n57911), .X(n29953) );
  nand_x1_sg U64518 ( .A(n53341), .B(n57875), .X(n29808) );
  nand_x1_sg U64519 ( .A(n51359), .B(n57886), .X(n29809) );
  nand_x1_sg U64520 ( .A(n50785), .B(n57878), .X(n29692) );
  nand_x1_sg U64521 ( .A(n56805), .B(n57895), .X(n29693) );
  nand_x1_sg U64522 ( .A(n53337), .B(n57876), .X(n29892) );
  nand_x1_sg U64523 ( .A(n51357), .B(n46207), .X(n29893) );
  nand_x1_sg U64524 ( .A(n53335), .B(n57872), .X(n30008) );
  nand_x1_sg U64525 ( .A(n51293), .B(n57898), .X(n30009) );
  nand_x1_sg U64526 ( .A(n53331), .B(n57875), .X(n29772) );
  nand_x1_sg U64527 ( .A(n51355), .B(n46207), .X(n29773) );
  nand_x1_sg U64528 ( .A(n53329), .B(n57875), .X(n29874) );
  nand_x1_sg U64529 ( .A(n51291), .B(n57915), .X(n29875) );
  nand_x1_sg U64530 ( .A(n53327), .B(n46212), .X(n29886) );
  nand_x1_sg U64531 ( .A(n47655), .B(n46207), .X(n29887) );
  nand_x1_sg U64532 ( .A(n53325), .B(n46212), .X(n29868) );
  nand_x1_sg U64533 ( .A(n47653), .B(n57898), .X(n29869) );
  nand_x1_sg U64534 ( .A(n53323), .B(n57880), .X(n29814) );
  nand_x1_sg U64535 ( .A(n51323), .B(n57899), .X(n29815) );
  nand_x1_sg U64536 ( .A(n53321), .B(n57875), .X(n29826) );
  nand_x1_sg U64537 ( .A(n47699), .B(n57910), .X(n29827) );
  nand_x1_sg U64538 ( .A(n53319), .B(n57878), .X(n29778) );
  nand_x1_sg U64539 ( .A(n51417), .B(n57895), .X(n29779) );
  nand_x1_sg U64540 ( .A(n50777), .B(n46209), .X(n29850) );
  nand_x1_sg U64541 ( .A(n56755), .B(n57896), .X(n29851) );
  nand_x1_sg U64542 ( .A(n53317), .B(n57876), .X(n29862) );
  nand_x1_sg U64543 ( .A(n51289), .B(n57898), .X(n29863) );
  nand_x1_sg U64544 ( .A(n53313), .B(n57871), .X(n29990) );
  nand_x1_sg U64545 ( .A(n51287), .B(n57893), .X(n29991) );
  nand_x1_sg U64546 ( .A(n53311), .B(n46209), .X(n29838) );
  nand_x1_sg U64547 ( .A(n51351), .B(n57908), .X(n29839) );
  nand_x1_sg U64548 ( .A(n50771), .B(n57877), .X(n29832) );
  nand_x1_sg U64549 ( .A(n56799), .B(n57909), .X(n29833) );
  nand_x1_sg U64550 ( .A(n53309), .B(n57875), .X(n29880) );
  nand_x1_sg U64551 ( .A(n51285), .B(n46207), .X(n29881) );
  nand_x1_sg U64552 ( .A(n53307), .B(n57877), .X(n30098) );
  nand_x1_sg U64553 ( .A(n47547), .B(n57897), .X(n30099) );
  nand_x1_sg U64554 ( .A(n53305), .B(n46212), .X(n29796) );
  nand_x1_sg U64555 ( .A(n51349), .B(n57896), .X(n29797) );
  nand_x1_sg U64556 ( .A(n50767), .B(n57875), .X(n29940) );
  nand_x1_sg U64557 ( .A(n56797), .B(n57903), .X(n29941) );
  nand_x1_sg U64558 ( .A(n53299), .B(n57878), .X(n29766) );
  nand_x1_sg U64559 ( .A(n51321), .B(n46207), .X(n29767) );
  nand_x1_sg U64560 ( .A(n50763), .B(n57876), .X(n30068) );
  nand_x1_sg U64561 ( .A(n56851), .B(n57903), .X(n30069) );
  nand_x1_sg U64562 ( .A(n53293), .B(n57872), .X(n29996) );
  nand_x1_sg U64563 ( .A(n51283), .B(n57894), .X(n29997) );
  nand_x1_sg U64564 ( .A(n50761), .B(n57880), .X(n29982) );
  nand_x1_sg U64565 ( .A(n56747), .B(n57895), .X(n29983) );
  nand_x1_sg U64566 ( .A(n53291), .B(n46209), .X(n29984) );
  nand_x1_sg U64567 ( .A(n51347), .B(n57891), .X(n29985) );
  nand_x1_sg U64568 ( .A(n53287), .B(n57873), .X(n30026) );
  nand_x1_sg U64569 ( .A(n51345), .B(n57910), .X(n30027) );
  nand_x1_sg U64570 ( .A(n50755), .B(n57873), .X(n30020) );
  nand_x1_sg U64571 ( .A(n56793), .B(n57900), .X(n30021) );
  nand_x1_sg U64572 ( .A(n53283), .B(n46210), .X(n30110) );
  nand_x1_sg U64573 ( .A(n47541), .B(n57897), .X(n30111) );
  nand_x1_sg U64574 ( .A(n53281), .B(n57877), .X(n30522) );
  nand_x1_sg U64575 ( .A(n51343), .B(n57890), .X(n30523) );
  nand_x1_sg U64576 ( .A(n53279), .B(n46209), .X(n30116) );
  nand_x1_sg U64577 ( .A(n47539), .B(n57911), .X(n30117) );
  nand_x1_sg U64578 ( .A(n53277), .B(n57870), .X(n29958) );
  nand_x1_sg U64579 ( .A(n47537), .B(n57907), .X(n29959) );
  nand_x1_sg U64580 ( .A(n50917), .B(n57876), .X(n30428) );
  nand_x1_sg U64581 ( .A(n56847), .B(n57903), .X(n30429) );
  nand_x1_sg U64582 ( .A(n53505), .B(n57877), .X(n30426) );
  nand_x1_sg U64583 ( .A(n51407), .B(n57904), .X(n30427) );
  nand_x1_sg U64584 ( .A(n53503), .B(n57876), .X(n30434) );
  nand_x1_sg U64585 ( .A(n47695), .B(n57899), .X(n30435) );
  nand_x1_sg U64586 ( .A(n50915), .B(n46212), .X(n30432) );
  nand_x1_sg U64587 ( .A(n56865), .B(n57887), .X(n30433) );
  nand_x1_sg U64588 ( .A(n50913), .B(n57876), .X(n30464) );
  nand_x1_sg U64589 ( .A(n56829), .B(n57893), .X(n30465) );
  nand_x1_sg U64590 ( .A(n53501), .B(n57870), .X(n30462) );
  nand_x1_sg U64591 ( .A(n51387), .B(n57894), .X(n30463) );
  nand_x1_sg U64592 ( .A(n50911), .B(n57876), .X(n30470) );
  nand_x1_sg U64593 ( .A(n56783), .B(n57893), .X(n30471) );
  nand_x1_sg U64594 ( .A(n53499), .B(n46212), .X(n30468) );
  nand_x1_sg U64595 ( .A(n51335), .B(n57893), .X(n30469) );
  nand_x1_sg U64596 ( .A(n50909), .B(n57871), .X(n30452) );
  nand_x1_sg U64597 ( .A(n56827), .B(n57894), .X(n30453) );
  nand_x1_sg U64598 ( .A(n53497), .B(n57878), .X(n30450) );
  nand_x1_sg U64599 ( .A(n51385), .B(n57894), .X(n30451) );
  nand_x1_sg U64600 ( .A(n50907), .B(n46209), .X(n30458) );
  nand_x1_sg U64601 ( .A(n56781), .B(n57894), .X(n30459) );
  nand_x1_sg U64602 ( .A(n53495), .B(n57871), .X(n30456) );
  nand_x1_sg U64603 ( .A(n51333), .B(n57894), .X(n30457) );
  nand_x1_sg U64604 ( .A(n50905), .B(n57877), .X(n30200) );
  nand_x1_sg U64605 ( .A(n56825), .B(n57896), .X(n30201) );
  nand_x1_sg U64606 ( .A(n53493), .B(n57880), .X(n30198) );
  nand_x1_sg U64607 ( .A(n51383), .B(n57896), .X(n30199) );
  nand_x1_sg U64608 ( .A(n53491), .B(n57877), .X(n30206) );
  nand_x1_sg U64609 ( .A(n47677), .B(n57896), .X(n30207) );
  nand_x1_sg U64610 ( .A(n50903), .B(n57875), .X(n30204) );
  nand_x1_sg U64611 ( .A(n56779), .B(n57896), .X(n30205) );
  nand_x1_sg U64612 ( .A(n53489), .B(n57875), .X(n30188) );
  nand_x1_sg U64613 ( .A(n51331), .B(n57909), .X(n30189) );
  nand_x1_sg U64614 ( .A(n53487), .B(n57880), .X(n30186) );
  nand_x1_sg U64615 ( .A(n51381), .B(n57898), .X(n30187) );
  nand_x1_sg U64616 ( .A(n53485), .B(n57876), .X(n30194) );
  nand_x1_sg U64617 ( .A(n47675), .B(n57896), .X(n30195) );
  nand_x1_sg U64618 ( .A(n53483), .B(n57878), .X(n30192) );
  nand_x1_sg U64619 ( .A(n47673), .B(n57896), .X(n30193) );
  nand_x1_sg U64620 ( .A(n53243), .B(n46209), .X(n30154) );
  nand_x1_sg U64621 ( .A(n47435), .B(n57911), .X(n30155) );
  nand_x1_sg U64622 ( .A(n53241), .B(n57878), .X(n30376) );
  nand_x1_sg U64623 ( .A(n47433), .B(n57895), .X(n30377) );
  nand_x1_sg U64624 ( .A(n53239), .B(n46212), .X(n30202) );
  nand_x1_sg U64625 ( .A(n47371), .B(n57896), .X(n30203) );
  nand_x1_sg U64626 ( .A(n50683), .B(n46213), .X(n29760) );
  nand_x1_sg U64627 ( .A(n56925), .B(n46207), .X(n29761) );
  nand_x1_sg U64628 ( .A(n53235), .B(n57880), .X(n29718) );
  nand_x1_sg U64629 ( .A(n47429), .B(n57909), .X(n29719) );
  nand_x1_sg U64630 ( .A(n53233), .B(n46210), .X(n30142) );
  nand_x1_sg U64631 ( .A(n47369), .B(n57898), .X(n30143) );
  nand_x1_sg U64632 ( .A(n50677), .B(n57872), .X(n30534) );
  nand_x1_sg U64633 ( .A(n56923), .B(n57889), .X(n30535) );
  nand_x1_sg U64634 ( .A(n53231), .B(n46213), .X(n29742) );
  nand_x1_sg U64635 ( .A(n47367), .B(n46207), .X(n29743) );
  nand_x1_sg U64636 ( .A(n53229), .B(n57878), .X(n29736) );
  nand_x1_sg U64637 ( .A(n47365), .B(n57900), .X(n29737) );
  nand_x1_sg U64638 ( .A(n50983), .B(n57873), .X(n30544) );
  nand_x1_sg U64639 ( .A(n56919), .B(n57910), .X(n30545) );
  nand_x1_sg U64640 ( .A(n53575), .B(n57877), .X(n30542) );
  nand_x1_sg U64641 ( .A(n47421), .B(n57889), .X(n30543) );
  nand_x1_sg U64642 ( .A(n53573), .B(n57870), .X(n30550) );
  nand_x1_sg U64643 ( .A(n47361), .B(n57908), .X(n30551) );
  nand_x1_sg U64644 ( .A(n50977), .B(n57870), .X(n30530) );
  nand_x1_sg U64645 ( .A(n56917), .B(n57889), .X(n30531) );
  nand_x1_sg U64646 ( .A(n53571), .B(n57871), .X(n30538) );
  nand_x1_sg U64647 ( .A(n47359), .B(n57889), .X(n30539) );
  nand_x1_sg U64648 ( .A(n53569), .B(n57873), .X(n30536) );
  nand_x1_sg U64649 ( .A(n47357), .B(n57889), .X(n30537) );
  nand_x1_sg U64650 ( .A(n53141), .B(n57875), .X(n29926) );
  nand_x1_sg U64651 ( .A(n51439), .B(n57901), .X(n29927) );
  nand_x1_sg U64652 ( .A(n53139), .B(n57875), .X(n29924) );
  nand_x1_sg U64653 ( .A(n51483), .B(n57910), .X(n29925) );
  nand_x1_sg U64654 ( .A(n53137), .B(n46212), .X(n29932) );
  nand_x1_sg U64655 ( .A(n47735), .B(n57908), .X(n29933) );
  nand_x1_sg U64656 ( .A(n53135), .B(n57884), .X(n29930) );
  nand_x1_sg U64657 ( .A(n47571), .B(n57909), .X(n29931) );
  nand_x1_sg U64658 ( .A(n53133), .B(n57878), .X(n29914) );
  nand_x1_sg U64659 ( .A(n51437), .B(n57900), .X(n29915) );
  nand_x1_sg U64660 ( .A(n50601), .B(n57875), .X(n29912) );
  nand_x1_sg U64661 ( .A(n56883), .B(n57910), .X(n29913) );
  nand_x1_sg U64662 ( .A(n53131), .B(n46209), .X(n29920) );
  nand_x1_sg U64663 ( .A(n51451), .B(n57887), .X(n29921) );
  nand_x1_sg U64664 ( .A(n53129), .B(n46210), .X(n29918) );
  nand_x1_sg U64665 ( .A(n47719), .B(n57908), .X(n29919) );
  nand_x1_sg U64666 ( .A(n53127), .B(n57871), .X(n29950) );
  nand_x1_sg U64667 ( .A(n51435), .B(n57904), .X(n29951) );
  nand_x1_sg U64668 ( .A(n50599), .B(n57876), .X(n29948) );
  nand_x1_sg U64669 ( .A(n56881), .B(n57902), .X(n29949) );
  nand_x1_sg U64670 ( .A(n53125), .B(n57870), .X(n29956) );
  nand_x1_sg U64671 ( .A(n51449), .B(n57909), .X(n29957) );
  nand_x1_sg U64672 ( .A(n53123), .B(n57871), .X(n29954) );
  nand_x1_sg U64673 ( .A(n47717), .B(n57900), .X(n29955) );
  nand_x1_sg U64674 ( .A(n53121), .B(n57875), .X(n29938) );
  nand_x1_sg U64675 ( .A(n51433), .B(n57887), .X(n29939) );
  nand_x1_sg U64676 ( .A(n50597), .B(n57878), .X(n29936) );
  nand_x1_sg U64677 ( .A(n56879), .B(n57900), .X(n29937) );
  nand_x1_sg U64678 ( .A(n53119), .B(n46209), .X(n29944) );
  nand_x1_sg U64679 ( .A(n47567), .B(n57910), .X(n29945) );
  nand_x1_sg U64680 ( .A(n53117), .B(n57877), .X(n29942) );
  nand_x1_sg U64681 ( .A(n51447), .B(n57910), .X(n29943) );
  nand_x1_sg U64682 ( .A(n53115), .B(n57878), .X(n29878) );
  nand_x1_sg U64683 ( .A(n47715), .B(n57910), .X(n29879) );
  nand_x1_sg U64684 ( .A(n50595), .B(n57877), .X(n29876) );
  nand_x1_sg U64685 ( .A(n56877), .B(n46207), .X(n29877) );
  nand_x1_sg U64686 ( .A(n53113), .B(n46210), .X(n29884) );
  nand_x1_sg U64687 ( .A(n47565), .B(n57908), .X(n29885) );
  nand_x1_sg U64688 ( .A(n53111), .B(n57876), .X(n29882) );
  nand_x1_sg U64689 ( .A(n47563), .B(n57900), .X(n29883) );
  nand_x1_sg U64690 ( .A(n50659), .B(n57877), .X(n30304) );
  nand_x1_sg U64691 ( .A(n56895), .B(n57887), .X(n30305) );
  nand_x1_sg U64692 ( .A(n53201), .B(n46210), .X(n29820) );
  nand_x1_sg U64693 ( .A(n47739), .B(n57898), .X(n29821) );
  nand_x1_sg U64694 ( .A(n50655), .B(n57878), .X(n29704) );
  nand_x1_sg U64695 ( .A(n56911), .B(n57896), .X(n29705) );
  nand_x1_sg U64696 ( .A(n50653), .B(n46212), .X(n29686) );
  nand_x1_sg U64697 ( .A(n56909), .B(n57900), .X(n29687) );
  nand_x1_sg U64698 ( .A(n53197), .B(n57882), .X(n29680) );
  nand_x1_sg U64699 ( .A(n51479), .B(n57907), .X(n29681) );
  nand_x1_sg U64700 ( .A(n50651), .B(n46210), .X(n29856) );
  nand_x1_sg U64701 ( .A(n56893), .B(n57898), .X(n29857) );
  nand_x1_sg U64702 ( .A(n53427), .B(n57873), .X(n29802) );
  nand_x1_sg U64703 ( .A(n51393), .B(n57895), .X(n29803) );
  nand_x1_sg U64704 ( .A(n53425), .B(n57875), .X(n29790) );
  nand_x1_sg U64705 ( .A(n47683), .B(n57898), .X(n29791) );
  nand_x1_sg U64706 ( .A(n53423), .B(n57877), .X(n30526) );
  nand_x1_sg U64707 ( .A(n51213), .B(n57890), .X(n30527) );
  nand_x1_sg U64708 ( .A(n53421), .B(n57872), .X(n30524) );
  nand_x1_sg U64709 ( .A(n47629), .B(n57890), .X(n30525) );
  nand_x1_sg U64710 ( .A(n50831), .B(n57876), .X(n29714) );
  nand_x1_sg U64711 ( .A(n56719), .B(n57887), .X(n29715) );
  nand_x1_sg U64712 ( .A(n53419), .B(n57878), .X(n29712) );
  nand_x1_sg U64713 ( .A(n51257), .B(n57898), .X(n29713) );
  nand_x1_sg U64714 ( .A(n53403), .B(n46213), .X(n30050) );
  nand_x1_sg U64715 ( .A(n51361), .B(n57888), .X(n30051) );
  nand_x1_sg U64716 ( .A(n53399), .B(n46213), .X(n30038) );
  nand_x1_sg U64717 ( .A(n47659), .B(n57897), .X(n30039) );
  nand_x1_sg U64718 ( .A(n53397), .B(n46209), .X(n30032) );
  nand_x1_sg U64719 ( .A(n47549), .B(n57908), .X(n30033) );
  nand_x1_sg U64720 ( .A(n53481), .B(n57880), .X(n30488) );
  nand_x1_sg U64721 ( .A(n51431), .B(n57892), .X(n30489) );
  nand_x1_sg U64722 ( .A(n53479), .B(n57877), .X(n30486) );
  nand_x1_sg U64723 ( .A(n51473), .B(n57892), .X(n30487) );
  nand_x1_sg U64724 ( .A(n53477), .B(n57875), .X(n30494) );
  nand_x1_sg U64725 ( .A(n47733), .B(n57892), .X(n30495) );
  nand_x1_sg U64726 ( .A(n53475), .B(n57876), .X(n30492) );
  nand_x1_sg U64727 ( .A(n47569), .B(n57892), .X(n30493) );
  nand_x1_sg U64728 ( .A(n53473), .B(n57880), .X(n30476) );
  nand_x1_sg U64729 ( .A(n51429), .B(n57893), .X(n30477) );
  nand_x1_sg U64730 ( .A(n50901), .B(n57880), .X(n30474) );
  nand_x1_sg U64731 ( .A(n56875), .B(n57893), .X(n30475) );
  nand_x1_sg U64732 ( .A(n53471), .B(n57878), .X(n30482) );
  nand_x1_sg U64733 ( .A(n51445), .B(n57892), .X(n30483) );
  nand_x1_sg U64734 ( .A(n53469), .B(n57877), .X(n30480) );
  nand_x1_sg U64735 ( .A(n47713), .B(n57892), .X(n30481) );
  nand_x1_sg U64736 ( .A(n53467), .B(n46213), .X(n30512) );
  nand_x1_sg U64737 ( .A(n51427), .B(n57890), .X(n30513) );
  nand_x1_sg U64738 ( .A(n50899), .B(n57877), .X(n30510) );
  nand_x1_sg U64739 ( .A(n56873), .B(n57891), .X(n30511) );
  nand_x1_sg U64740 ( .A(n53465), .B(n57875), .X(n30518) );
  nand_x1_sg U64741 ( .A(n51443), .B(n57890), .X(n30519) );
  nand_x1_sg U64742 ( .A(n53463), .B(n46212), .X(n30516) );
  nand_x1_sg U64743 ( .A(n47711), .B(n57890), .X(n30517) );
  nand_x1_sg U64744 ( .A(n53461), .B(n57878), .X(n30500) );
  nand_x1_sg U64745 ( .A(n51425), .B(n57891), .X(n30501) );
  nand_x1_sg U64746 ( .A(n50897), .B(n46212), .X(n30498) );
  nand_x1_sg U64747 ( .A(n56871), .B(n57891), .X(n30499) );
  nand_x1_sg U64748 ( .A(n53459), .B(n46212), .X(n30506) );
  nand_x1_sg U64749 ( .A(n47561), .B(n57891), .X(n30507) );
  nand_x1_sg U64750 ( .A(n53457), .B(n57870), .X(n30504) );
  nand_x1_sg U64751 ( .A(n51441), .B(n57891), .X(n30505) );
  nand_x1_sg U64752 ( .A(n53455), .B(n46212), .X(n30440) );
  nand_x1_sg U64753 ( .A(n47709), .B(n57899), .X(n30441) );
  nand_x1_sg U64754 ( .A(n50895), .B(n46212), .X(n30438) );
  nand_x1_sg U64755 ( .A(n56869), .B(n57901), .X(n30439) );
  nand_x1_sg U64756 ( .A(n53453), .B(n57875), .X(n30446) );
  nand_x1_sg U64757 ( .A(n47559), .B(n57908), .X(n30447) );
  nand_x1_sg U64758 ( .A(n53451), .B(n57876), .X(n30444) );
  nand_x1_sg U64759 ( .A(n47557), .B(n57911), .X(n30445) );
  nand_x1_sg U64760 ( .A(n50959), .B(n46210), .X(n30164) );
  nand_x1_sg U64761 ( .A(n56889), .B(n57908), .X(n30165) );
  nand_x1_sg U64762 ( .A(n50957), .B(n46209), .X(n30162) );
  nand_x1_sg U64763 ( .A(n56913), .B(n57887), .X(n30163) );
  nand_x1_sg U64764 ( .A(n53543), .B(n46210), .X(n30170) );
  nand_x1_sg U64765 ( .A(n51485), .B(n57899), .X(n30171) );
  nand_x1_sg U64766 ( .A(n53541), .B(n46209), .X(n30168) );
  nand_x1_sg U64767 ( .A(n47737), .B(n57910), .X(n30169) );
  nand_x1_sg U64768 ( .A(n50955), .B(n57880), .X(n30296) );
  nand_x1_sg U64769 ( .A(n56903), .B(n57886), .X(n30297) );
  nand_x1_sg U64770 ( .A(n53539), .B(n57880), .X(n30294) );
  nand_x1_sg U64771 ( .A(n51471), .B(n57911), .X(n30295) );
  nand_x1_sg U64772 ( .A(n50953), .B(n57873), .X(n30302) );
  nand_x1_sg U64773 ( .A(n56901), .B(n57908), .X(n30303) );
  nand_x1_sg U64774 ( .A(n53537), .B(n57880), .X(n30300) );
  nand_x1_sg U64775 ( .A(n51469), .B(n57897), .X(n30301) );
  nand_x1_sg U64776 ( .A(n50951), .B(n57880), .X(n30284) );
  nand_x1_sg U64777 ( .A(n56887), .B(n57895), .X(n30285) );
  nand_x1_sg U64778 ( .A(n53535), .B(n57880), .X(n30282) );
  nand_x1_sg U64779 ( .A(n51457), .B(n57908), .X(n30283) );
  nand_x1_sg U64780 ( .A(n50949), .B(n57880), .X(n30290) );
  nand_x1_sg U64781 ( .A(n56899), .B(n57887), .X(n30291) );
  nand_x1_sg U64782 ( .A(n53533), .B(n57880), .X(n30288) );
  nand_x1_sg U64783 ( .A(n51467), .B(n57896), .X(n30289) );
  nand_x1_sg U64784 ( .A(n50947), .B(n57878), .X(n30320) );
  nand_x1_sg U64785 ( .A(n56885), .B(n57907), .X(n30321) );
  nand_x1_sg U64786 ( .A(n53531), .B(n57877), .X(n30318) );
  nand_x1_sg U64787 ( .A(n51455), .B(n57898), .X(n30319) );
  nand_x1_sg U64788 ( .A(n53529), .B(n57877), .X(n30326) );
  nand_x1_sg U64789 ( .A(n47725), .B(n57896), .X(n30327) );
  nand_x1_sg U64790 ( .A(n50945), .B(n57880), .X(n30324) );
  nand_x1_sg U64791 ( .A(n56897), .B(n57898), .X(n30325) );
  nand_x1_sg U64792 ( .A(n53527), .B(n57875), .X(n30308) );
  nand_x1_sg U64793 ( .A(n51465), .B(n57908), .X(n30309) );
  nand_x1_sg U64794 ( .A(n53525), .B(n57876), .X(n30306) );
  nand_x1_sg U64795 ( .A(n51453), .B(n57889), .X(n30307) );
  nand_x1_sg U64796 ( .A(n53523), .B(n46213), .X(n30314) );
  nand_x1_sg U64797 ( .A(n47723), .B(n57890), .X(n30315) );
  nand_x1_sg U64798 ( .A(n53521), .B(n57873), .X(n30312) );
  nand_x1_sg U64799 ( .A(n47721), .B(n57888), .X(n30313) );
  nand_x1_sg U64800 ( .A(n50643), .B(n57880), .X(n30406) );
  nand_x1_sg U64801 ( .A(n55083), .B(n57898), .X(n30407) );
  nand_x1_sg U64802 ( .A(n50637), .B(n57878), .X(n30340) );
  nand_x1_sg U64803 ( .A(n55155), .B(n57886), .X(n30341) );
  nand_x1_sg U64804 ( .A(n53179), .B(n46209), .X(n29898) );
  nand_x1_sg U64805 ( .A(n51149), .B(n46207), .X(n29899) );
  nand_x1_sg U64806 ( .A(n50629), .B(n57875), .X(n30268) );
  nand_x1_sg U64807 ( .A(n55081), .B(n57896), .X(n30269) );
  nand_x1_sg U64808 ( .A(n53177), .B(n57872), .X(n30322) );
  nand_x1_sg U64809 ( .A(n51145), .B(n57911), .X(n30323) );
  nand_x1_sg U64810 ( .A(n50623), .B(n57875), .X(n30472) );
  nand_x1_sg U64811 ( .A(n55079), .B(n57893), .X(n30473) );
  nand_x1_sg U64812 ( .A(n53175), .B(n57877), .X(n30442) );
  nand_x1_sg U64813 ( .A(n51143), .B(n57898), .X(n30443) );
  nand_x1_sg U64814 ( .A(n53169), .B(n57877), .X(n30208) );
  nand_x1_sg U64815 ( .A(n47609), .B(n57910), .X(n30209) );
  nand_x1_sg U64816 ( .A(n53167), .B(n57871), .X(n30508) );
  nand_x1_sg U64817 ( .A(n47607), .B(n57891), .X(n30509) );
  nand_x1_sg U64818 ( .A(n50675), .B(n57876), .X(n30358) );
  nand_x1_sg U64819 ( .A(n55251), .B(n57908), .X(n30359) );
  nand_x1_sg U64820 ( .A(n53217), .B(n46213), .X(n29784) );
  nand_x1_sg U64821 ( .A(n51169), .B(n57907), .X(n29785) );
  nand_x1_sg U64822 ( .A(n53215), .B(n46213), .X(n29904) );
  nand_x1_sg U64823 ( .A(n51167), .B(n57909), .X(n29905) );
  nand_x1_sg U64824 ( .A(n53213), .B(n57878), .X(n30044) );
  nand_x1_sg U64825 ( .A(n51165), .B(n57910), .X(n30045) );
  nand_x1_sg U64826 ( .A(n53211), .B(n46212), .X(n29910) );
  nand_x1_sg U64827 ( .A(n47515), .B(n57908), .X(n29911) );
  nand_x1_sg U64828 ( .A(n53209), .B(n46213), .X(n29710) );
  nand_x1_sg U64829 ( .A(n51163), .B(n46207), .X(n29711) );
  nand_x1_sg U64830 ( .A(n50663), .B(n57875), .X(n29754) );
  nand_x1_sg U64831 ( .A(n55235), .B(n57911), .X(n29755) );
  nand_x1_sg U64832 ( .A(n50661), .B(n57882), .X(n29730) );
  nand_x1_sg U64833 ( .A(n55233), .B(n57896), .X(n29731) );
  nand_x1_sg U64834 ( .A(n53207), .B(n57878), .X(n30196) );
  nand_x1_sg U64835 ( .A(n47513), .B(n57896), .X(n30197) );
  nand_x1_sg U64836 ( .A(n53205), .B(n57878), .X(n30382) );
  nand_x1_sg U64837 ( .A(n47511), .B(n57886), .X(n30383) );
  nand_x1_sg U64838 ( .A(n50943), .B(n57876), .X(n30224) );
  nand_x1_sg U64839 ( .A(n55077), .B(n57910), .X(n30225) );
  nand_x1_sg U64840 ( .A(n50937), .B(n46213), .X(n30228) );
  nand_x1_sg U64841 ( .A(n55153), .B(n57908), .X(n30229) );
  nand_x1_sg U64842 ( .A(n50935), .B(n57880), .X(n30212) );
  nand_x1_sg U64843 ( .A(n55085), .B(n57907), .X(n30213) );
  nand_x1_sg U64844 ( .A(n53519), .B(n57880), .X(n30210) );
  nand_x1_sg U64845 ( .A(n51147), .B(n57899), .X(n30211) );
  nand_x1_sg U64846 ( .A(n50929), .B(n46209), .X(n30152) );
  nand_x1_sg U64847 ( .A(n55075), .B(n57895), .X(n30153) );
  nand_x1_sg U64848 ( .A(n53517), .B(n46210), .X(n30150) );
  nand_x1_sg U64849 ( .A(n51139), .B(n57886), .X(n30151) );
  nand_x1_sg U64850 ( .A(n50923), .B(n46209), .X(n30140) );
  nand_x1_sg U64851 ( .A(n55073), .B(n57909), .X(n30141) );
  nand_x1_sg U64852 ( .A(n53515), .B(n46210), .X(n30138) );
  nand_x1_sg U64853 ( .A(n51137), .B(n57887), .X(n30139) );
  nand_x1_sg U64854 ( .A(n53513), .B(n46209), .X(n30146) );
  nand_x1_sg U64855 ( .A(n47605), .B(n57887), .X(n30147) );
  nand_x1_sg U64856 ( .A(n53511), .B(n57878), .X(n30174) );
  nand_x1_sg U64857 ( .A(n51135), .B(n57886), .X(n30175) );
  nand_x1_sg U64858 ( .A(n53509), .B(n46213), .X(n30182) );
  nand_x1_sg U64859 ( .A(n47603), .B(n57896), .X(n30183) );
  nand_x1_sg U64860 ( .A(n53507), .B(n57875), .X(n30180) );
  nand_x1_sg U64861 ( .A(n47601), .B(n57907), .X(n30181) );
  nand_x1_sg U64862 ( .A(n53567), .B(n46212), .X(n30248) );
  nand_x1_sg U64863 ( .A(n47613), .B(n57895), .X(n30249) );
  nand_x1_sg U64864 ( .A(n53565), .B(n57880), .X(n30246) );
  nand_x1_sg U64865 ( .A(n51179), .B(n57895), .X(n30247) );
  nand_x1_sg U64866 ( .A(n50975), .B(n57876), .X(n30254) );
  nand_x1_sg U64867 ( .A(n55249), .B(n57895), .X(n30255) );
  nand_x1_sg U64868 ( .A(n53563), .B(n57877), .X(n30252) );
  nand_x1_sg U64869 ( .A(n47517), .B(n57895), .X(n30253) );
  nand_x1_sg U64870 ( .A(n53561), .B(n57882), .X(n30236) );
  nand_x1_sg U64871 ( .A(n51175), .B(n57908), .X(n30237) );
  nand_x1_sg U64872 ( .A(n50973), .B(n57876), .X(n30234) );
  nand_x1_sg U64873 ( .A(n55245), .B(n57896), .X(n30235) );
  nand_x1_sg U64874 ( .A(n53559), .B(n57876), .X(n30242) );
  nand_x1_sg U64875 ( .A(n51161), .B(n57895), .X(n30243) );
  nand_x1_sg U64876 ( .A(n50971), .B(n57880), .X(n30240) );
  nand_x1_sg U64877 ( .A(n55231), .B(n57895), .X(n30241) );
  nand_x1_sg U64878 ( .A(n53557), .B(n57880), .X(n30272) );
  nand_x1_sg U64879 ( .A(n51159), .B(n57896), .X(n30273) );
  nand_x1_sg U64880 ( .A(n50969), .B(n57875), .X(n30270) );
  nand_x1_sg U64881 ( .A(n55229), .B(n57895), .X(n30271) );
  nand_x1_sg U64882 ( .A(n53555), .B(n57878), .X(n30278) );
  nand_x1_sg U64883 ( .A(n51157), .B(n57911), .X(n30279) );
  nand_x1_sg U64884 ( .A(n50967), .B(n46213), .X(n30276) );
  nand_x1_sg U64885 ( .A(n55227), .B(n57887), .X(n30277) );
  nand_x1_sg U64886 ( .A(n53553), .B(n57875), .X(n30260) );
  nand_x1_sg U64887 ( .A(n51155), .B(n57911), .X(n30261) );
  nand_x1_sg U64888 ( .A(n50965), .B(n57876), .X(n30258) );
  nand_x1_sg U64889 ( .A(n55225), .B(n57886), .X(n30259) );
  nand_x1_sg U64890 ( .A(n53551), .B(n57876), .X(n30266) );
  nand_x1_sg U64891 ( .A(n47509), .B(n57907), .X(n30267) );
  nand_x1_sg U64892 ( .A(n53549), .B(n57877), .X(n30264) );
  nand_x1_sg U64893 ( .A(n51153), .B(n57898), .X(n30265) );
  nand_x1_sg U64894 ( .A(n50431), .B(n46212), .X(n29724) );
  nand_x1_sg U64895 ( .A(n55259), .B(n46207), .X(n29725) );
  nand_x1_sg U64896 ( .A(n50425), .B(n57875), .X(n30220) );
  nand_x1_sg U64897 ( .A(n55283), .B(n57886), .X(n30221) );
  nand_x1_sg U64898 ( .A(n50417), .B(n57878), .X(n30250) );
  nand_x1_sg U64899 ( .A(n55279), .B(n57895), .X(n30251) );
  nand_x1_sg U64900 ( .A(n50415), .B(n57877), .X(n30466) );
  nand_x1_sg U64901 ( .A(n55257), .B(n57893), .X(n30467) );
  nand_x1_sg U64902 ( .A(n50409), .B(n57875), .X(n30490) );
  nand_x1_sg U64903 ( .A(n55277), .B(n57892), .X(n30491) );
  nand_x1_sg U64904 ( .A(n52909), .B(n46213), .X(n30484) );
  nand_x1_sg U64905 ( .A(n51195), .B(n57892), .X(n30485) );
  nand_x1_sg U64906 ( .A(n50401), .B(n57872), .X(n30394) );
  nand_x1_sg U64907 ( .A(n55273), .B(n57886), .X(n30395) );
  nand_x1_sg U64908 ( .A(n52907), .B(n46212), .X(n30370) );
  nand_x1_sg U64909 ( .A(n51189), .B(n57911), .X(n30371) );
  nand_x1_sg U64910 ( .A(n52905), .B(n57876), .X(n30346) );
  nand_x1_sg U64911 ( .A(n51187), .B(n57895), .X(n30347) );
  nand_x1_sg U64912 ( .A(n50731), .B(n57880), .X(n30568) );
  nand_x1_sg U64913 ( .A(n55255), .B(n57888), .X(n30569) );
  nand_x1_sg U64914 ( .A(n50725), .B(n57875), .X(n30572) );
  nand_x1_sg U64915 ( .A(n55271), .B(n57888), .X(n30573) );
  nand_x1_sg U64916 ( .A(n50723), .B(n57871), .X(n30556) );
  nand_x1_sg U64917 ( .A(n55269), .B(n57910), .X(n30557) );
  nand_x1_sg U64918 ( .A(n53251), .B(n57872), .X(n30554) );
  nand_x1_sg U64919 ( .A(n51193), .B(n57908), .X(n30555) );
  nand_x1_sg U64920 ( .A(n50717), .B(n57875), .X(n30262) );
  nand_x1_sg U64921 ( .A(n55267), .B(n57903), .X(n30263) );
  nand_x1_sg U64922 ( .A(n50715), .B(n46210), .X(n30136) );
  nand_x1_sg U64923 ( .A(n55253), .B(n46207), .X(n30137) );
  nand_x1_sg U64924 ( .A(n50709), .B(n57876), .X(n30226) );
  nand_x1_sg U64925 ( .A(n55265), .B(n57895), .X(n30227) );
  nand_x1_sg U64926 ( .A(n50707), .B(n57876), .X(n29748) );
  nand_x1_sg U64927 ( .A(n55263), .B(n57896), .X(n29749) );
  nand_x1_sg U64928 ( .A(n50701), .B(n57870), .X(n30528) );
  nand_x1_sg U64929 ( .A(n55261), .B(n57889), .X(n30529) );
  nand_x1_sg U64930 ( .A(n53247), .B(n46212), .X(n30570) );
  nand_x1_sg U64931 ( .A(n51185), .B(n57888), .X(n30571) );
  nand_x1_sg U64932 ( .A(n53245), .B(n57877), .X(n30400) );
  nand_x1_sg U64933 ( .A(n51183), .B(n57887), .X(n30401) );
  nand_x1_sg U64934 ( .A(n50699), .B(n57882), .X(n30172) );
  nand_x1_sg U64935 ( .A(n55315), .B(n57887), .X(n30173) );
  nand_x1_sg U64936 ( .A(n50697), .B(n46212), .X(n30424) );
  nand_x1_sg U64937 ( .A(n55313), .B(n57902), .X(n30425) );
  nand_x1_sg U64938 ( .A(n50693), .B(n57880), .X(n30190) );
  nand_x1_sg U64939 ( .A(n55307), .B(n57895), .X(n30191) );
  nand_x1_sg U64940 ( .A(n50691), .B(n57877), .X(n30184) );
  nand_x1_sg U64941 ( .A(n55305), .B(n57900), .X(n30185) );
  nand_x1_sg U64942 ( .A(n50685), .B(n57873), .X(n30460) );
  nand_x1_sg U64943 ( .A(n55301), .B(n57894), .X(n30461) );
  nand_x1_sg U64944 ( .A(n50981), .B(n57873), .X(n30548) );
  nand_x1_sg U64945 ( .A(n55287), .B(n57895), .X(n30549) );
  nand_x1_sg U64946 ( .A(n50979), .B(n57871), .X(n30532) );
  nand_x1_sg U64947 ( .A(n55285), .B(n57889), .X(n30533) );
  nand_x1_sg U64948 ( .A(n50641), .B(n46210), .X(n30148) );
  nand_x1_sg U64949 ( .A(n55061), .B(n57907), .X(n30149) );
  nand_x1_sg U64950 ( .A(n50639), .B(n46212), .X(n30364) );
  nand_x1_sg U64951 ( .A(n55059), .B(n57909), .X(n30365) );
  nand_x1_sg U64952 ( .A(n50627), .B(n57878), .X(n29698) );
  nand_x1_sg U64953 ( .A(n55017), .B(n57895), .X(n29699) );
  nand_x1_sg U64954 ( .A(n50625), .B(n57880), .X(n30292) );
  nand_x1_sg U64955 ( .A(n55015), .B(n57895), .X(n30293) );
  nand_x1_sg U64956 ( .A(n50427), .B(n57877), .X(n30214) );
  nand_x1_sg U64957 ( .A(n55055), .B(n57908), .X(n30215) );
  nand_x1_sg U64958 ( .A(n50421), .B(n57877), .X(n30546) );
  nand_x1_sg U64959 ( .A(n55053), .B(n57888), .X(n30547) );
  nand_x1_sg U64960 ( .A(n50419), .B(n57870), .X(n30540) );
  nand_x1_sg U64961 ( .A(n55051), .B(n57889), .X(n30541) );
  nand_x1_sg U64962 ( .A(n50413), .B(n46212), .X(n30244) );
  nand_x1_sg U64963 ( .A(n55049), .B(n57895), .X(n30245) );
  nand_x1_sg U64964 ( .A(n50411), .B(n57877), .X(n30238) );
  nand_x1_sg U64965 ( .A(n55047), .B(n57900), .X(n30239) );
  nand_x1_sg U64966 ( .A(n50405), .B(n57880), .X(n30274) );
  nand_x1_sg U64967 ( .A(n55045), .B(n57896), .X(n30275) );
  nand_x1_sg U64968 ( .A(n50403), .B(n46213), .X(n30454) );
  nand_x1_sg U64969 ( .A(n55043), .B(n57894), .X(n30455) );
  nand_x1_sg U64970 ( .A(n50941), .B(n57880), .X(n30222) );
  nand_x1_sg U64971 ( .A(n55041), .B(n57887), .X(n30223) );
  nand_x1_sg U64972 ( .A(n50939), .B(n57875), .X(n30230) );
  nand_x1_sg U64973 ( .A(n55039), .B(n57907), .X(n30231) );
  nand_x1_sg U64974 ( .A(n50933), .B(n46213), .X(n30218) );
  nand_x1_sg U64975 ( .A(n55009), .B(n57899), .X(n30219) );
  nand_x1_sg U64976 ( .A(n50931), .B(n57877), .X(n30216) );
  nand_x1_sg U64977 ( .A(n55007), .B(n57909), .X(n30217) );
  nand_x1_sg U64978 ( .A(n50927), .B(n46210), .X(n30158) );
  nand_x1_sg U64979 ( .A(n55005), .B(n57896), .X(n30159) );
  nand_x1_sg U64980 ( .A(n50925), .B(n46209), .X(n30156) );
  nand_x1_sg U64981 ( .A(n55003), .B(n57911), .X(n30157) );
  nand_x1_sg U64982 ( .A(n50921), .B(n46210), .X(n30144) );
  nand_x1_sg U64983 ( .A(n55001), .B(n57909), .X(n30145) );
  nand_x1_sg U64984 ( .A(n50919), .B(n46213), .X(n30176) );
  nand_x1_sg U64985 ( .A(n54999), .B(n57909), .X(n30177) );
  nand_x1_sg U64986 ( .A(n50729), .B(n46210), .X(n30566) );
  nand_x1_sg U64987 ( .A(n55037), .B(n57888), .X(n30567) );
  nand_x1_sg U64988 ( .A(n50727), .B(n57878), .X(n30574) );
  nand_x1_sg U64989 ( .A(n55035), .B(n57888), .X(n30575) );
  nand_x1_sg U64990 ( .A(n50721), .B(n57880), .X(n30562) );
  nand_x1_sg U64991 ( .A(n55033), .B(n57888), .X(n30563) );
  nand_x1_sg U64992 ( .A(n50719), .B(n57875), .X(n30560) );
  nand_x1_sg U64993 ( .A(n55031), .B(n57888), .X(n30561) );
  nand_x1_sg U64994 ( .A(n50713), .B(n46213), .X(n30564) );
  nand_x1_sg U64995 ( .A(n55029), .B(n57888), .X(n30565) );
  nand_x1_sg U64996 ( .A(n50711), .B(n46213), .X(n30558) );
  nand_x1_sg U64997 ( .A(n55027), .B(n57910), .X(n30559) );
  nand_x1_sg U64998 ( .A(n50705), .B(n46209), .X(n30134) );
  nand_x1_sg U64999 ( .A(n55025), .B(n57907), .X(n30135) );
  nand_x1_sg U65000 ( .A(n50703), .B(n57877), .X(n30520) );
  nand_x1_sg U65001 ( .A(n55023), .B(n57890), .X(n30521) );
  nand_x1_sg U65002 ( .A(n57644), .B(n50399), .X(n36381) );
  nand_x1_sg U65003 ( .A(n52903), .B(n46201), .X(n36382) );
  nand_x1_sg U65004 ( .A(n57672), .B(n50397), .X(n36389) );
  nand_x1_sg U65005 ( .A(n52901), .B(n46200), .X(n36390) );
  nand_x1_sg U65006 ( .A(n57672), .B(n50395), .X(n36391) );
  nand_x1_sg U65007 ( .A(n52899), .B(n57728), .X(n36392) );
  nand_x1_sg U65008 ( .A(n57675), .B(n50393), .X(n36433) );
  nand_x1_sg U65009 ( .A(n52897), .B(n57761), .X(n36434) );
  nand_x1_sg U65010 ( .A(n57673), .B(n50391), .X(n36435) );
  nand_x1_sg U65011 ( .A(n52895), .B(n57747), .X(n36436) );
  nand_x1_sg U65012 ( .A(n57680), .B(n50389), .X(n36427) );
  nand_x1_sg U65013 ( .A(n52893), .B(n57759), .X(n36428) );
  nand_x1_sg U65014 ( .A(n57717), .B(n50355), .X(n36637) );
  nand_x1_sg U65015 ( .A(n52859), .B(n57766), .X(n36638) );
  nand_x1_sg U65016 ( .A(n57700), .B(n50353), .X(n36639) );
  nand_x1_sg U65017 ( .A(n52857), .B(n57758), .X(n36640) );
  nand_x1_sg U65018 ( .A(n57697), .B(n50351), .X(n36631) );
  nand_x1_sg U65019 ( .A(n52855), .B(n57748), .X(n36632) );
  nand_x1_sg U65020 ( .A(n57698), .B(n50349), .X(n36633) );
  nand_x1_sg U65021 ( .A(n52853), .B(n57760), .X(n36634) );
  nand_x1_sg U65022 ( .A(n57680), .B(n50347), .X(n36661) );
  nand_x1_sg U65023 ( .A(n52851), .B(n57741), .X(n36662) );
  nand_x1_sg U65024 ( .A(n52851), .B(n57720), .X(n36649) );
  nand_x1_sg U65025 ( .A(n49081), .B(n57740), .X(n36650) );
  nand_x1_sg U65026 ( .A(n57682), .B(n50345), .X(n36663) );
  nand_x1_sg U65027 ( .A(n52849), .B(n57735), .X(n36664) );
  nand_x1_sg U65028 ( .A(n52849), .B(n57720), .X(n36651) );
  nand_x1_sg U65029 ( .A(n49083), .B(n57741), .X(n36652) );
  nand_x1_sg U65030 ( .A(n57681), .B(n50343), .X(n36655) );
  nand_x1_sg U65031 ( .A(n52847), .B(n57740), .X(n36656) );
  nand_x1_sg U65032 ( .A(n52847), .B(n57703), .X(n36643) );
  nand_x1_sg U65033 ( .A(n49085), .B(n57742), .X(n36644) );
  nand_x1_sg U65034 ( .A(n57720), .B(n50341), .X(n36657) );
  nand_x1_sg U65035 ( .A(n52845), .B(n57741), .X(n36658) );
  nand_x1_sg U65036 ( .A(n52845), .B(n57695), .X(n36645) );
  nand_x1_sg U65037 ( .A(n49087), .B(n57744), .X(n36646) );
  nand_x1_sg U65038 ( .A(n57681), .B(n50339), .X(n36673) );
  nand_x1_sg U65039 ( .A(n52843), .B(n57736), .X(n36674) );
  nand_x1_sg U65040 ( .A(n52843), .B(n57698), .X(n36613) );
  nand_x1_sg U65041 ( .A(n49089), .B(n46197), .X(n36614) );
  nand_x1_sg U65042 ( .A(n57682), .B(n50337), .X(n36675) );
  nand_x1_sg U65043 ( .A(n52841), .B(n46200), .X(n36676) );
  nand_x1_sg U65044 ( .A(n52841), .B(n57703), .X(n36615) );
  nand_x1_sg U65045 ( .A(n49091), .B(n57743), .X(n36616) );
  nand_x1_sg U65046 ( .A(n57680), .B(n50335), .X(n36667) );
  nand_x1_sg U65047 ( .A(n52839), .B(n57761), .X(n36668) );
  nand_x1_sg U65048 ( .A(n52839), .B(n57682), .X(n36607) );
  nand_x1_sg U65049 ( .A(n49093), .B(n46200), .X(n36608) );
  nand_x1_sg U65050 ( .A(n57634), .B(n50333), .X(n36669) );
  nand_x1_sg U65051 ( .A(n52837), .B(n57760), .X(n36670) );
  nand_x1_sg U65052 ( .A(n52837), .B(n57695), .X(n36609) );
  nand_x1_sg U65053 ( .A(n49095), .B(n46198), .X(n36610) );
  nand_x1_sg U65054 ( .A(n57681), .B(n50331), .X(n36589) );
  nand_x1_sg U65055 ( .A(n52835), .B(n57742), .X(n36590) );
  nand_x1_sg U65056 ( .A(n52835), .B(n57681), .X(n36625) );
  nand_x1_sg U65057 ( .A(n49097), .B(n57744), .X(n36626) );
  nand_x1_sg U65058 ( .A(n57682), .B(n50329), .X(n36591) );
  nand_x1_sg U65059 ( .A(n52833), .B(n57743), .X(n36592) );
  nand_x1_sg U65060 ( .A(n52833), .B(n57682), .X(n36627) );
  nand_x1_sg U65061 ( .A(n49099), .B(n57759), .X(n36628) );
  nand_x1_sg U65062 ( .A(n57680), .B(n50327), .X(n36583) );
  nand_x1_sg U65063 ( .A(n52831), .B(n57742), .X(n36584) );
  nand_x1_sg U65064 ( .A(n52831), .B(n57680), .X(n36619) );
  nand_x1_sg U65065 ( .A(n49101), .B(n57763), .X(n36620) );
  nand_x1_sg U65066 ( .A(n57634), .B(n50325), .X(n36585) );
  nand_x1_sg U65067 ( .A(n52829), .B(n46200), .X(n36586) );
  nand_x1_sg U65068 ( .A(n52829), .B(n57634), .X(n36621) );
  nand_x1_sg U65069 ( .A(n49103), .B(n57764), .X(n36622) );
  nand_x1_sg U65070 ( .A(n57681), .B(n50323), .X(n36601) );
  nand_x1_sg U65071 ( .A(n52827), .B(n46200), .X(n36602) );
  nand_x1_sg U65072 ( .A(n52827), .B(n57704), .X(n36685) );
  nand_x1_sg U65073 ( .A(n49105), .B(n57733), .X(n36686) );
  nand_x1_sg U65074 ( .A(n57715), .B(n50321), .X(n36603) );
  nand_x1_sg U65075 ( .A(n52825), .B(n46197), .X(n36604) );
  nand_x1_sg U65076 ( .A(n52825), .B(n57720), .X(n36687) );
  nand_x1_sg U65077 ( .A(n49107), .B(n57749), .X(n36688) );
  nand_x1_sg U65078 ( .A(n57720), .B(n50319), .X(n36595) );
  nand_x1_sg U65079 ( .A(n52823), .B(n57743), .X(n36596) );
  nand_x1_sg U65080 ( .A(n52823), .B(n57700), .X(n36679) );
  nand_x1_sg U65081 ( .A(n49109), .B(n57736), .X(n36680) );
  nand_x1_sg U65082 ( .A(n57696), .B(n50317), .X(n36597) );
  nand_x1_sg U65083 ( .A(n52821), .B(n57742), .X(n36598) );
  nand_x1_sg U65084 ( .A(n52821), .B(n57709), .X(n36681) );
  nand_x1_sg U65085 ( .A(n49111), .B(n57732), .X(n36682) );
  nand_x1_sg U65086 ( .A(n57716), .B(n50315), .X(n36577) );
  nand_x1_sg U65087 ( .A(n52819), .B(n46197), .X(n36578) );
  nand_x1_sg U65088 ( .A(n52819), .B(n57703), .X(n36697) );
  nand_x1_sg U65089 ( .A(n49113), .B(n46201), .X(n36698) );
  nand_x1_sg U65090 ( .A(n57634), .B(n50313), .X(n36579) );
  nand_x1_sg U65091 ( .A(n52817), .B(n46198), .X(n36580) );
  nand_x1_sg U65092 ( .A(n52817), .B(n57715), .X(n36699) );
  nand_x1_sg U65093 ( .A(n49115), .B(n57749), .X(n36700) );
  nand_x1_sg U65094 ( .A(n57715), .B(n50311), .X(n36571) );
  nand_x1_sg U65095 ( .A(n52815), .B(n46197), .X(n36572) );
  nand_x1_sg U65096 ( .A(n52815), .B(n57701), .X(n36691) );
  nand_x1_sg U65097 ( .A(n49117), .B(n57750), .X(n36692) );
  nand_x1_sg U65098 ( .A(n57720), .B(n50309), .X(n36573) );
  nand_x1_sg U65099 ( .A(n52813), .B(n46198), .X(n36574) );
  nand_x1_sg U65100 ( .A(n52813), .B(n57702), .X(n36693) );
  nand_x1_sg U65101 ( .A(n49119), .B(n57764), .X(n36694) );
  nand_x1_sg U65102 ( .A(n52803), .B(n57700), .X(n36565) );
  nand_x1_sg U65103 ( .A(n48839), .B(n57755), .X(n36566) );
  nand_x1_sg U65104 ( .A(n57698), .B(n50297), .X(n36843) );
  nand_x1_sg U65105 ( .A(n52801), .B(n57724), .X(n36844) );
  nand_x1_sg U65106 ( .A(n52801), .B(n57680), .X(n36567) );
  nand_x1_sg U65107 ( .A(n48841), .B(n46197), .X(n36568) );
  nand_x1_sg U65108 ( .A(n57682), .B(n50295), .X(n36835) );
  nand_x1_sg U65109 ( .A(n52799), .B(n57731), .X(n36836) );
  nand_x1_sg U65110 ( .A(n52799), .B(n57681), .X(n36559) );
  nand_x1_sg U65111 ( .A(n48843), .B(n57756), .X(n36560) );
  nand_x1_sg U65112 ( .A(n57703), .B(n50293), .X(n36837) );
  nand_x1_sg U65113 ( .A(n52797), .B(n57759), .X(n36838) );
  nand_x1_sg U65114 ( .A(n52797), .B(n57682), .X(n36561) );
  nand_x1_sg U65115 ( .A(n48845), .B(n57744), .X(n36562) );
  nand_x1_sg U65116 ( .A(n57701), .B(n50291), .X(n36805) );
  nand_x1_sg U65117 ( .A(n52795), .B(n57765), .X(n36806) );
  nand_x1_sg U65118 ( .A(n52795), .B(n57697), .X(n36553) );
  nand_x1_sg U65119 ( .A(n48847), .B(n57756), .X(n36554) );
  nand_x1_sg U65120 ( .A(n57717), .B(n50289), .X(n36807) );
  nand_x1_sg U65121 ( .A(n52793), .B(n46200), .X(n36808) );
  nand_x1_sg U65122 ( .A(n52793), .B(n57698), .X(n36555) );
  nand_x1_sg U65123 ( .A(n48849), .B(n57755), .X(n36556) );
  nand_x1_sg U65124 ( .A(n57709), .B(n50287), .X(n36799) );
  nand_x1_sg U65125 ( .A(n52791), .B(n57763), .X(n36800) );
  nand_x1_sg U65126 ( .A(n52791), .B(n57709), .X(n36547) );
  nand_x1_sg U65127 ( .A(n48851), .B(n57742), .X(n36548) );
  nand_x1_sg U65128 ( .A(n57708), .B(n50285), .X(n36801) );
  nand_x1_sg U65129 ( .A(n52789), .B(n57764), .X(n36802) );
  nand_x1_sg U65130 ( .A(n52789), .B(n57718), .X(n36549) );
  nand_x1_sg U65131 ( .A(n48853), .B(n57742), .X(n36550) );
  nand_x1_sg U65132 ( .A(n57718), .B(n50283), .X(n36817) );
  nand_x1_sg U65133 ( .A(n52787), .B(n57764), .X(n36818) );
  nand_x1_sg U65134 ( .A(n52787), .B(n57642), .X(n36445) );
  nand_x1_sg U65135 ( .A(n48855), .B(n57772), .X(n36446) );
  nand_x1_sg U65136 ( .A(n57680), .B(n50281), .X(n36819) );
  nand_x1_sg U65137 ( .A(n52785), .B(n57743), .X(n36820) );
  nand_x1_sg U65138 ( .A(n52785), .B(n57642), .X(n36447) );
  nand_x1_sg U65139 ( .A(n48857), .B(n57763), .X(n36448) );
  nand_x1_sg U65140 ( .A(n57717), .B(n50279), .X(n36811) );
  nand_x1_sg U65141 ( .A(n52783), .B(n57725), .X(n36812) );
  nand_x1_sg U65142 ( .A(n52783), .B(n57717), .X(n36439) );
  nand_x1_sg U65143 ( .A(n48859), .B(n57772), .X(n36440) );
  nand_x1_sg U65144 ( .A(n57718), .B(n50277), .X(n36813) );
  nand_x1_sg U65145 ( .A(n52781), .B(n46197), .X(n36814) );
  nand_x1_sg U65146 ( .A(n52781), .B(n57642), .X(n36441) );
  nand_x1_sg U65147 ( .A(n48861), .B(n57726), .X(n36442) );
  nand_x1_sg U65148 ( .A(n57697), .B(n50275), .X(n36877) );
  nand_x1_sg U65149 ( .A(n52779), .B(n57755), .X(n36878) );
  nand_x1_sg U65150 ( .A(n52779), .B(n57642), .X(n36457) );
  nand_x1_sg U65151 ( .A(n48863), .B(n57748), .X(n36458) );
  nand_x1_sg U65152 ( .A(n57698), .B(n50273), .X(n36879) );
  nand_x1_sg U65153 ( .A(n52777), .B(n46198), .X(n36880) );
  nand_x1_sg U65154 ( .A(n52777), .B(n57641), .X(n36459) );
  nand_x1_sg U65155 ( .A(n48865), .B(n46197), .X(n36460) );
  nand_x1_sg U65156 ( .A(n57718), .B(n50271), .X(n36871) );
  nand_x1_sg U65157 ( .A(n52775), .B(n57728), .X(n36872) );
  nand_x1_sg U65158 ( .A(n52775), .B(n57642), .X(n36451) );
  nand_x1_sg U65159 ( .A(n48867), .B(n57727), .X(n36452) );
  nand_x1_sg U65160 ( .A(n57715), .B(n50269), .X(n36873) );
  nand_x1_sg U65161 ( .A(n52773), .B(n57748), .X(n36874) );
  nand_x1_sg U65162 ( .A(n52773), .B(n57642), .X(n36453) );
  nand_x1_sg U65163 ( .A(n48869), .B(n57724), .X(n36454) );
  nand_x1_sg U65164 ( .A(n57717), .B(n50267), .X(n36889) );
  nand_x1_sg U65165 ( .A(n52771), .B(n57739), .X(n36890) );
  nand_x1_sg U65166 ( .A(n52771), .B(n57681), .X(n36829) );
  nand_x1_sg U65167 ( .A(n48871), .B(n57759), .X(n36830) );
  nand_x1_sg U65168 ( .A(n57694), .B(n50265), .X(n36891) );
  nand_x1_sg U65169 ( .A(n52769), .B(n57739), .X(n36892) );
  nand_x1_sg U65170 ( .A(n52769), .B(n57702), .X(n36831) );
  nand_x1_sg U65171 ( .A(n48873), .B(n57775), .X(n36832) );
  nand_x1_sg U65172 ( .A(n57718), .B(n50263), .X(n36883) );
  nand_x1_sg U65173 ( .A(n52767), .B(n46197), .X(n36884) );
  nand_x1_sg U65174 ( .A(n52767), .B(n57634), .X(n36823) );
  nand_x1_sg U65175 ( .A(n48875), .B(n57761), .X(n36824) );
  nand_x1_sg U65176 ( .A(n57720), .B(n50261), .X(n36885) );
  nand_x1_sg U65177 ( .A(n52765), .B(n57728), .X(n36886) );
  nand_x1_sg U65178 ( .A(n52765), .B(n57717), .X(n36825) );
  nand_x1_sg U65179 ( .A(n48877), .B(n57762), .X(n36826) );
  nand_x1_sg U65180 ( .A(n57703), .B(n50259), .X(n36853) );
  nand_x1_sg U65181 ( .A(n52763), .B(n57728), .X(n36854) );
  nand_x1_sg U65182 ( .A(n52763), .B(n57701), .X(n36841) );
  nand_x1_sg U65183 ( .A(n48879), .B(n57763), .X(n36842) );
  nand_x1_sg U65184 ( .A(n57705), .B(n50257), .X(n36723) );
  nand_x1_sg U65185 ( .A(n52761), .B(n57761), .X(n36724) );
  nand_x1_sg U65186 ( .A(n52761), .B(n57699), .X(n36855) );
  nand_x1_sg U65187 ( .A(n48881), .B(n57746), .X(n36856) );
  nand_x1_sg U65188 ( .A(n57715), .B(n50255), .X(n36715) );
  nand_x1_sg U65189 ( .A(n52759), .B(n57770), .X(n36716) );
  nand_x1_sg U65190 ( .A(n52759), .B(n57702), .X(n36847) );
  nand_x1_sg U65191 ( .A(n48883), .B(n57728), .X(n36848) );
  nand_x1_sg U65192 ( .A(n57720), .B(n50253), .X(n36717) );
  nand_x1_sg U65193 ( .A(n52757), .B(n57762), .X(n36718) );
  nand_x1_sg U65194 ( .A(n52757), .B(n57706), .X(n36849) );
  nand_x1_sg U65195 ( .A(n48885), .B(n57766), .X(n36850) );
  nand_x1_sg U65196 ( .A(n57715), .B(n50251), .X(n36781) );
  nand_x1_sg U65197 ( .A(n52755), .B(n57746), .X(n36782) );
  nand_x1_sg U65198 ( .A(n52755), .B(n57700), .X(n36865) );
  nand_x1_sg U65199 ( .A(n48887), .B(n57743), .X(n36866) );
  nand_x1_sg U65200 ( .A(n57634), .B(n50249), .X(n36783) );
  nand_x1_sg U65201 ( .A(n52753), .B(n57759), .X(n36784) );
  nand_x1_sg U65202 ( .A(n52753), .B(n57720), .X(n36867) );
  nand_x1_sg U65203 ( .A(n48889), .B(n57765), .X(n36868) );
  nand_x1_sg U65204 ( .A(n57708), .B(n50247), .X(n36775) );
  nand_x1_sg U65205 ( .A(n52751), .B(n57760), .X(n36776) );
  nand_x1_sg U65206 ( .A(n52751), .B(n57693), .X(n36859) );
  nand_x1_sg U65207 ( .A(n48891), .B(n57743), .X(n36860) );
  nand_x1_sg U65208 ( .A(n57680), .B(n50245), .X(n36777) );
  nand_x1_sg U65209 ( .A(n52749), .B(n57758), .X(n36778) );
  nand_x1_sg U65210 ( .A(n52749), .B(n57694), .X(n36861) );
  nand_x1_sg U65211 ( .A(n48893), .B(n57746), .X(n36862) );
  nand_x1_sg U65212 ( .A(n57709), .B(n50243), .X(n36793) );
  nand_x1_sg U65213 ( .A(n52747), .B(n46201), .X(n36794) );
  nand_x1_sg U65214 ( .A(n52747), .B(n57705), .X(n36733) );
  nand_x1_sg U65215 ( .A(n48895), .B(n57742), .X(n36734) );
  nand_x1_sg U65216 ( .A(n57708), .B(n50241), .X(n36795) );
  nand_x1_sg U65217 ( .A(n52745), .B(n46200), .X(n36796) );
  nand_x1_sg U65218 ( .A(n52745), .B(n57699), .X(n36735) );
  nand_x1_sg U65219 ( .A(n48897), .B(n57747), .X(n36736) );
  nand_x1_sg U65220 ( .A(n57708), .B(n50239), .X(n36787) );
  nand_x1_sg U65221 ( .A(n52743), .B(n57746), .X(n36788) );
  nand_x1_sg U65222 ( .A(n52743), .B(n57708), .X(n36727) );
  nand_x1_sg U65223 ( .A(n48899), .B(n57765), .X(n36728) );
  nand_x1_sg U65224 ( .A(n57709), .B(n50237), .X(n36789) );
  nand_x1_sg U65225 ( .A(n52741), .B(n57759), .X(n36790) );
  nand_x1_sg U65226 ( .A(n52741), .B(n57709), .X(n36729) );
  nand_x1_sg U65227 ( .A(n48901), .B(n57770), .X(n36730) );
  nand_x1_sg U65228 ( .A(n57709), .B(n50235), .X(n36757) );
  nand_x1_sg U65229 ( .A(n52739), .B(n57741), .X(n36758) );
  nand_x1_sg U65230 ( .A(n52739), .B(n57702), .X(n36745) );
  nand_x1_sg U65231 ( .A(n48903), .B(n57741), .X(n36746) );
  nand_x1_sg U65232 ( .A(n57634), .B(n50233), .X(n36759) );
  nand_x1_sg U65233 ( .A(n52737), .B(n57740), .X(n36760) );
  nand_x1_sg U65234 ( .A(n52737), .B(n57706), .X(n36747) );
  nand_x1_sg U65235 ( .A(n48905), .B(n57741), .X(n36748) );
  nand_x1_sg U65236 ( .A(n57707), .B(n50231), .X(n36751) );
  nand_x1_sg U65237 ( .A(n52735), .B(n57741), .X(n36752) );
  nand_x1_sg U65238 ( .A(n52735), .B(n57704), .X(n36739) );
  nand_x1_sg U65239 ( .A(n48907), .B(n57747), .X(n36740) );
  nand_x1_sg U65240 ( .A(n57705), .B(n50229), .X(n36753) );
  nand_x1_sg U65241 ( .A(n52733), .B(n57741), .X(n36754) );
  nand_x1_sg U65242 ( .A(n52733), .B(n57695), .X(n36741) );
  nand_x1_sg U65243 ( .A(n48909), .B(n57759), .X(n36742) );
  nand_x1_sg U65244 ( .A(n57699), .B(n50227), .X(n36769) );
  nand_x1_sg U65245 ( .A(n52731), .B(n57740), .X(n36770) );
  nand_x1_sg U65246 ( .A(n52731), .B(n57682), .X(n36709) );
  nand_x1_sg U65247 ( .A(n48911), .B(n57750), .X(n36710) );
  nand_x1_sg U65248 ( .A(n57700), .B(n50225), .X(n36771) );
  nand_x1_sg U65249 ( .A(n52729), .B(n57740), .X(n36772) );
  nand_x1_sg U65250 ( .A(n52729), .B(n57703), .X(n36711) );
  nand_x1_sg U65251 ( .A(n48913), .B(n57749), .X(n36712) );
  nand_x1_sg U65252 ( .A(n57715), .B(n50223), .X(n36763) );
  nand_x1_sg U65253 ( .A(n52727), .B(n57740), .X(n36764) );
  nand_x1_sg U65254 ( .A(n52727), .B(n57698), .X(n36703) );
  nand_x1_sg U65255 ( .A(n48915), .B(n57750), .X(n36704) );
  nand_x1_sg U65256 ( .A(n57681), .B(n50221), .X(n36765) );
  nand_x1_sg U65257 ( .A(n52725), .B(n57740), .X(n36766) );
  nand_x1_sg U65258 ( .A(n52725), .B(n57701), .X(n36705) );
  nand_x1_sg U65259 ( .A(n48917), .B(n57748), .X(n36706) );
  nand_x1_sg U65260 ( .A(n52723), .B(n57716), .X(n36721) );
  nand_x1_sg U65261 ( .A(n48919), .B(n57762), .X(n36722) );
  nand_x1_sg U65262 ( .A(n57644), .B(n50215), .X(n36369) );
  nand_x1_sg U65263 ( .A(n52719), .B(n57772), .X(n36370) );
  nand_x1_sg U65264 ( .A(n57644), .B(n50213), .X(n36371) );
  nand_x1_sg U65265 ( .A(n52717), .B(n46200), .X(n36372) );
  nand_x1_sg U65266 ( .A(n52689), .B(n57645), .X(n36359) );
  nand_x1_sg U65267 ( .A(n48953), .B(n46198), .X(n36360) );
  nand_x1_sg U65268 ( .A(n52683), .B(n57645), .X(n36367) );
  nand_x1_sg U65269 ( .A(n48959), .B(n57763), .X(n36368) );
  nand_x1_sg U65270 ( .A(n57717), .B(n50171), .X(n36489) );
  nand_x1_sg U65271 ( .A(n52675), .B(n57743), .X(n36490) );
  nand_x1_sg U65272 ( .A(n57715), .B(n50169), .X(n36491) );
  nand_x1_sg U65273 ( .A(n52673), .B(n57743), .X(n36492) );
  nand_x1_sg U65274 ( .A(n57641), .B(n50167), .X(n36483) );
  nand_x1_sg U65275 ( .A(n52671), .B(n57763), .X(n36484) );
  nand_x1_sg U65276 ( .A(n57647), .B(n50165), .X(n36485) );
  nand_x1_sg U65277 ( .A(n52669), .B(n57760), .X(n36486) );
  nand_x1_sg U65278 ( .A(n57699), .B(n50163), .X(n36501) );
  nand_x1_sg U65279 ( .A(n52667), .B(n57743), .X(n36502) );
  nand_x1_sg U65280 ( .A(n57718), .B(n50161), .X(n36503) );
  nand_x1_sg U65281 ( .A(n52665), .B(n46201), .X(n36504) );
  nand_x1_sg U65282 ( .A(n57707), .B(n50159), .X(n36495) );
  nand_x1_sg U65283 ( .A(n52663), .B(n57743), .X(n36496) );
  nand_x1_sg U65284 ( .A(n57682), .B(n50157), .X(n36497) );
  nand_x1_sg U65285 ( .A(n52661), .B(n57743), .X(n36498) );
  nand_x1_sg U65286 ( .A(n57695), .B(n50155), .X(n36477) );
  nand_x1_sg U65287 ( .A(n52659), .B(n57758), .X(n36478) );
  nand_x1_sg U65288 ( .A(n57695), .B(n50153), .X(n36479) );
  nand_x1_sg U65289 ( .A(n52657), .B(n57765), .X(n36480) );
  nand_x1_sg U65290 ( .A(n57641), .B(n50151), .X(n36471) );
  nand_x1_sg U65291 ( .A(n52655), .B(n57743), .X(n36472) );
  nand_x1_sg U65292 ( .A(n57641), .B(n50149), .X(n36473) );
  nand_x1_sg U65293 ( .A(n52653), .B(n57746), .X(n36474) );
  nand_x1_sg U65294 ( .A(n57695), .B(n50147), .X(n36481) );
  nand_x1_sg U65295 ( .A(n52651), .B(n57749), .X(n36482) );
  nand_x1_sg U65296 ( .A(n57641), .B(n50145), .X(n36469) );
  nand_x1_sg U65297 ( .A(n52649), .B(n46201), .X(n36470) );
  nand_x1_sg U65298 ( .A(n57641), .B(n50143), .X(n36475) );
  nand_x1_sg U65299 ( .A(n52647), .B(n57750), .X(n36476) );
  nand_x1_sg U65300 ( .A(n57641), .B(n50141), .X(n36467) );
  nand_x1_sg U65301 ( .A(n52645), .B(n57725), .X(n36468) );
  nand_x1_sg U65302 ( .A(n57720), .B(n50139), .X(n36529) );
  nand_x1_sg U65303 ( .A(n52643), .B(n46201), .X(n36530) );
  nand_x1_sg U65304 ( .A(n57698), .B(n50137), .X(n36511) );
  nand_x1_sg U65305 ( .A(n52641), .B(n46198), .X(n36512) );
  nand_x1_sg U65306 ( .A(n52641), .B(n57708), .X(n36531) );
  nand_x1_sg U65307 ( .A(n49001), .B(n57742), .X(n36532) );
  nand_x1_sg U65308 ( .A(n57672), .B(n50135), .X(n36395) );
  nand_x1_sg U65309 ( .A(n52639), .B(n57762), .X(n36396) );
  nand_x1_sg U65310 ( .A(n52639), .B(n57709), .X(n36523) );
  nand_x1_sg U65311 ( .A(n49003), .B(n46200), .X(n36524) );
  nand_x1_sg U65312 ( .A(n57672), .B(n50133), .X(n36397) );
  nand_x1_sg U65313 ( .A(n52637), .B(n46197), .X(n36398) );
  nand_x1_sg U65314 ( .A(n52637), .B(n57634), .X(n36525) );
  nand_x1_sg U65315 ( .A(n49005), .B(n57743), .X(n36526) );
  nand_x1_sg U65316 ( .A(n57672), .B(n50131), .X(n36393) );
  nand_x1_sg U65317 ( .A(n52635), .B(n57761), .X(n36394) );
  nand_x1_sg U65318 ( .A(n52635), .B(n57720), .X(n36527) );
  nand_x1_sg U65319 ( .A(n49007), .B(n57742), .X(n36528) );
  nand_x1_sg U65320 ( .A(n57644), .B(n50129), .X(n36375) );
  nand_x1_sg U65321 ( .A(n52633), .B(n46201), .X(n36376) );
  nand_x1_sg U65322 ( .A(n52633), .B(n57697), .X(n36507) );
  nand_x1_sg U65323 ( .A(n49009), .B(n57743), .X(n36508) );
  nand_x1_sg U65324 ( .A(n57643), .B(n50127), .X(n36407) );
  nand_x1_sg U65325 ( .A(n52631), .B(n57764), .X(n36408) );
  nand_x1_sg U65326 ( .A(n52631), .B(n57715), .X(n36519) );
  nand_x1_sg U65327 ( .A(n49011), .B(n46201), .X(n36520) );
  nand_x1_sg U65328 ( .A(n57643), .B(n50125), .X(n36409) );
  nand_x1_sg U65329 ( .A(n52629), .B(n57766), .X(n36410) );
  nand_x1_sg U65330 ( .A(n52629), .B(n57716), .X(n36521) );
  nand_x1_sg U65331 ( .A(n49013), .B(n57743), .X(n36522) );
  nand_x1_sg U65332 ( .A(n57672), .B(n50123), .X(n36401) );
  nand_x1_sg U65333 ( .A(n52627), .B(n57754), .X(n36402) );
  nand_x1_sg U65334 ( .A(n52627), .B(n57699), .X(n36499) );
  nand_x1_sg U65335 ( .A(n49015), .B(n57743), .X(n36500) );
  nand_x1_sg U65336 ( .A(n57704), .B(n50121), .X(n36403) );
  nand_x1_sg U65337 ( .A(n52625), .B(n57766), .X(n36404) );
  nand_x1_sg U65338 ( .A(n52625), .B(n57708), .X(n36487) );
  nand_x1_sg U65339 ( .A(n49017), .B(n57743), .X(n36488) );
  nand_x1_sg U65340 ( .A(n57644), .B(n50119), .X(n36383) );
  nand_x1_sg U65341 ( .A(n52623), .B(n46200), .X(n36384) );
  nand_x1_sg U65342 ( .A(n52623), .B(n57681), .X(n36505) );
  nand_x1_sg U65343 ( .A(n49019), .B(n46200), .X(n36506) );
  nand_x1_sg U65344 ( .A(n57644), .B(n50117), .X(n36385) );
  nand_x1_sg U65345 ( .A(n52621), .B(n46201), .X(n36386) );
  nand_x1_sg U65346 ( .A(n52621), .B(n57634), .X(n36493) );
  nand_x1_sg U65347 ( .A(n49021), .B(n57743), .X(n36494) );
  nand_x1_sg U65348 ( .A(n57644), .B(n50115), .X(n36377) );
  nand_x1_sg U65349 ( .A(n52619), .B(n46200), .X(n36378) );
  nand_x1_sg U65350 ( .A(n52619), .B(n57700), .X(n36515) );
  nand_x1_sg U65351 ( .A(n49023), .B(n57742), .X(n36516) );
  nand_x1_sg U65352 ( .A(n57644), .B(n50113), .X(n36379) );
  nand_x1_sg U65353 ( .A(n52617), .B(n57763), .X(n36380) );
  nand_x1_sg U65354 ( .A(n52617), .B(n57709), .X(n36517) );
  nand_x1_sg U65355 ( .A(n49025), .B(n46197), .X(n36518) );
  nand_x1_sg U65356 ( .A(n57672), .B(n50111), .X(n36387) );
  nand_x1_sg U65357 ( .A(n52615), .B(n57772), .X(n36388) );
  nand_x1_sg U65358 ( .A(n52615), .B(n57715), .X(n36509) );
  nand_x1_sg U65359 ( .A(n49027), .B(n57757), .X(n36510) );
  nand_x1_sg U65360 ( .A(n57702), .B(n50109), .X(n37043) );
  nand_x1_sg U65361 ( .A(n52613), .B(n57759), .X(n37044) );
  nand_x1_sg U65362 ( .A(n52613), .B(n57708), .X(n36429) );
  nand_x1_sg U65363 ( .A(n48633), .B(n57762), .X(n36430) );
  nand_x1_sg U65364 ( .A(n57634), .B(n50107), .X(n37055) );
  nand_x1_sg U65365 ( .A(n52611), .B(n57731), .X(n37056) );
  nand_x1_sg U65366 ( .A(n52611), .B(n57641), .X(n36461) );
  nand_x1_sg U65367 ( .A(n48635), .B(n57764), .X(n36462) );
  nand_x1_sg U65368 ( .A(n57697), .B(n50105), .X(n37061) );
  nand_x1_sg U65369 ( .A(n52609), .B(n57731), .X(n37062) );
  nand_x1_sg U65370 ( .A(n52609), .B(n57709), .X(n36425) );
  nand_x1_sg U65371 ( .A(n48637), .B(n57728), .X(n36426) );
  nand_x1_sg U65372 ( .A(n52607), .B(n57641), .X(n36463) );
  nand_x1_sg U65373 ( .A(n48639), .B(n57772), .X(n36464) );
  nand_x1_sg U65374 ( .A(n52605), .B(n57641), .X(n36465) );
  nand_x1_sg U65375 ( .A(n48641), .B(n57763), .X(n36466) );
  nand_x1_sg U65376 ( .A(n52603), .B(n57704), .X(n36399) );
  nand_x1_sg U65377 ( .A(n48643), .B(n57727), .X(n36400) );
  nand_x1_sg U65378 ( .A(n52601), .B(n57643), .X(n36413) );
  nand_x1_sg U65379 ( .A(n48645), .B(n46198), .X(n36414) );
  nand_x1_sg U65380 ( .A(n52599), .B(n57643), .X(n36419) );
  nand_x1_sg U65381 ( .A(n48647), .B(n57772), .X(n36420) );
  nand_x1_sg U65382 ( .A(n52597), .B(n57643), .X(n36411) );
  nand_x1_sg U65383 ( .A(n48649), .B(n46200), .X(n36412) );
  nand_x1_sg U65384 ( .A(n52595), .B(n57643), .X(n36421) );
  nand_x1_sg U65385 ( .A(n48651), .B(n57764), .X(n36422) );
  nand_x1_sg U65386 ( .A(n52593), .B(n57681), .X(n36423) );
  nand_x1_sg U65387 ( .A(n48653), .B(n57757), .X(n36424) );
  nand_x1_sg U65388 ( .A(n52591), .B(n57643), .X(n36415) );
  nand_x1_sg U65389 ( .A(n48655), .B(n57764), .X(n36416) );
  nand_x1_sg U65390 ( .A(n52589), .B(n57643), .X(n36417) );
  nand_x1_sg U65391 ( .A(n48657), .B(n57724), .X(n36418) );
  nand_x1_sg U65392 ( .A(n57700), .B(n50021), .X(n37343) );
  nand_x1_sg U65393 ( .A(n52525), .B(n57726), .X(n37344) );
  nand_x1_sg U65394 ( .A(n57718), .B(n50019), .X(n37355) );
  nand_x1_sg U65395 ( .A(n52523), .B(n57725), .X(n37356) );
  nand_x1_sg U65396 ( .A(n57718), .B(n50017), .X(n37357) );
  nand_x1_sg U65397 ( .A(n52521), .B(n57725), .X(n37358) );
  nand_x1_sg U65398 ( .A(n57717), .B(n50015), .X(n37351) );
  nand_x1_sg U65399 ( .A(n52519), .B(n57725), .X(n37352) );
  nand_x1_sg U65400 ( .A(n57707), .B(n50013), .X(n37353) );
  nand_x1_sg U65401 ( .A(n52517), .B(n57725), .X(n37354) );
  nand_x1_sg U65402 ( .A(n52505), .B(n57708), .X(n37345) );
  nand_x1_sg U65403 ( .A(n48741), .B(n57726), .X(n37346) );
  nand_x1_sg U65404 ( .A(n52501), .B(n57709), .X(n37339) );
  nand_x1_sg U65405 ( .A(n48745), .B(n57726), .X(n37340) );
  nand_x1_sg U65406 ( .A(n52491), .B(n57708), .X(n37347) );
  nand_x1_sg U65407 ( .A(n48755), .B(n57726), .X(n37348) );
  nand_x1_sg U65408 ( .A(n52489), .B(n57705), .X(n37349) );
  nand_x1_sg U65409 ( .A(n48757), .B(n57726), .X(n37350) );
  nand_x1_sg U65410 ( .A(n52487), .B(n57706), .X(n37341) );
  nand_x1_sg U65411 ( .A(n48759), .B(n57726), .X(n37342) );
  nand_x1_sg U65412 ( .A(n57682), .B(n49911), .X(n37227) );
  nand_x1_sg U65413 ( .A(n52415), .B(n57746), .X(n37228) );
  nand_x1_sg U65414 ( .A(n57682), .B(n49909), .X(n37219) );
  nand_x1_sg U65415 ( .A(n52413), .B(n57743), .X(n37220) );
  nand_x1_sg U65416 ( .A(n57682), .B(n49907), .X(n37221) );
  nand_x1_sg U65417 ( .A(n52411), .B(n57765), .X(n37222) );
  nand_x1_sg U65418 ( .A(n57682), .B(n49851), .X(n36755) );
  nand_x1_sg U65419 ( .A(n52355), .B(n57741), .X(n36756) );
  nand_x1_sg U65420 ( .A(n57680), .B(n49849), .X(n36761) );
  nand_x1_sg U65421 ( .A(n52353), .B(n57740), .X(n36762) );
  nand_x1_sg U65422 ( .A(n57709), .B(n49847), .X(n36779) );
  nand_x1_sg U65423 ( .A(n52351), .B(n57761), .X(n36780) );
  nand_x1_sg U65424 ( .A(n57682), .B(n49845), .X(n36767) );
  nand_x1_sg U65425 ( .A(n52349), .B(n57740), .X(n36768) );
  nand_x1_sg U65426 ( .A(n57681), .B(n49843), .X(n36581) );
  nand_x1_sg U65427 ( .A(n52347), .B(n46198), .X(n36582) );
  nand_x1_sg U65428 ( .A(n57715), .B(n49841), .X(n36665) );
  nand_x1_sg U65429 ( .A(n52345), .B(n57758), .X(n36666) );
  nand_x1_sg U65430 ( .A(n57708), .B(n49839), .X(n36671) );
  nand_x1_sg U65431 ( .A(n52343), .B(n57742), .X(n36672) );
  nand_x1_sg U65432 ( .A(n57702), .B(n49837), .X(n36713) );
  nand_x1_sg U65433 ( .A(n52341), .B(n57762), .X(n36714) );
  nand_x1_sg U65434 ( .A(n57707), .B(n49833), .X(n36851) );
  nand_x1_sg U65435 ( .A(n52337), .B(n57757), .X(n36852) );
  nand_x1_sg U65436 ( .A(n57634), .B(n49831), .X(n36863) );
  nand_x1_sg U65437 ( .A(n52335), .B(n57747), .X(n36864) );
  nand_x1_sg U65438 ( .A(n57680), .B(n49829), .X(n36575) );
  nand_x1_sg U65439 ( .A(n52333), .B(n46197), .X(n36576) );
  nand_x1_sg U65440 ( .A(n57634), .B(n49827), .X(n36791) );
  nand_x1_sg U65441 ( .A(n52331), .B(n57760), .X(n36792) );
  nand_x1_sg U65442 ( .A(n57720), .B(n49825), .X(n36551) );
  nand_x1_sg U65443 ( .A(n52329), .B(n57728), .X(n36552) );
  nand_x1_sg U65444 ( .A(n52329), .B(n57681), .X(n36797) );
  nand_x1_sg U65445 ( .A(n48521), .B(n57766), .X(n36798) );
  nand_x1_sg U65446 ( .A(n57704), .B(n49823), .X(n36617) );
  nand_x1_sg U65447 ( .A(n52327), .B(n57772), .X(n36618) );
  nand_x1_sg U65448 ( .A(n57682), .B(n49821), .X(n36605) );
  nand_x1_sg U65449 ( .A(n52325), .B(n57772), .X(n36606) );
  nand_x1_sg U65450 ( .A(n57642), .B(n49819), .X(n36443) );
  nand_x1_sg U65451 ( .A(n52323), .B(n57725), .X(n36444) );
  nand_x1_sg U65452 ( .A(n52323), .B(n57695), .X(n37139) );
  nand_x1_sg U65453 ( .A(n48527), .B(n57743), .X(n37140) );
  nand_x1_sg U65454 ( .A(n57642), .B(n49817), .X(n36449) );
  nand_x1_sg U65455 ( .A(n52321), .B(n46200), .X(n36450) );
  nand_x1_sg U65456 ( .A(n52321), .B(n57696), .X(n37145) );
  nand_x1_sg U65457 ( .A(n48529), .B(n57728), .X(n37146) );
  nand_x1_sg U65458 ( .A(n57642), .B(n49815), .X(n36455) );
  nand_x1_sg U65459 ( .A(n52319), .B(n46201), .X(n36456) );
  nand_x1_sg U65460 ( .A(n52319), .B(n57682), .X(n37157) );
  nand_x1_sg U65461 ( .A(n48531), .B(n57728), .X(n37158) );
  nand_x1_sg U65462 ( .A(n57698), .B(n49813), .X(n36557) );
  nand_x1_sg U65463 ( .A(n52317), .B(n57746), .X(n36558) );
  nand_x1_sg U65464 ( .A(n52317), .B(n57682), .X(n37163) );
  nand_x1_sg U65465 ( .A(n48533), .B(n57766), .X(n37164) );
  nand_x1_sg U65466 ( .A(n57680), .B(n49807), .X(n36569) );
  nand_x1_sg U65467 ( .A(n52311), .B(n46198), .X(n36570) );
  nand_x1_sg U65468 ( .A(n52307), .B(n57681), .X(n36887) );
  nand_x1_sg U65469 ( .A(n48543), .B(n57739), .X(n36888) );
  nand_x1_sg U65470 ( .A(n52305), .B(n57700), .X(n37007) );
  nand_x1_sg U65471 ( .A(n48545), .B(n57733), .X(n37008) );
  nand_x1_sg U65472 ( .A(n57682), .B(n49799), .X(n36647) );
  nand_x1_sg U65473 ( .A(n52303), .B(n57758), .X(n36648) );
  nand_x1_sg U65474 ( .A(n52303), .B(n57693), .X(n37025) );
  nand_x1_sg U65475 ( .A(n48547), .B(n57732), .X(n37026) );
  nand_x1_sg U65476 ( .A(n57705), .B(n49797), .X(n36677) );
  nand_x1_sg U65477 ( .A(n52301), .B(n57760), .X(n36678) );
  nand_x1_sg U65478 ( .A(n52301), .B(n57699), .X(n37013) );
  nand_x1_sg U65479 ( .A(n48549), .B(n57733), .X(n37014) );
  nand_x1_sg U65480 ( .A(n57720), .B(n49795), .X(n36653) );
  nand_x1_sg U65481 ( .A(n52299), .B(n57743), .X(n36654) );
  nand_x1_sg U65482 ( .A(n52299), .B(n57720), .X(n36815) );
  nand_x1_sg U65483 ( .A(n48551), .B(n57758), .X(n36816) );
  nand_x1_sg U65484 ( .A(n57680), .B(n49793), .X(n36659) );
  nand_x1_sg U65485 ( .A(n52297), .B(n57761), .X(n36660) );
  nand_x1_sg U65486 ( .A(n52297), .B(n57708), .X(n36833) );
  nand_x1_sg U65487 ( .A(n48553), .B(n57765), .X(n36834) );
  nand_x1_sg U65488 ( .A(n57706), .B(n49791), .X(n36689) );
  nand_x1_sg U65489 ( .A(n52295), .B(n57748), .X(n36690) );
  nand_x1_sg U65490 ( .A(n52295), .B(n57680), .X(n36869) );
  nand_x1_sg U65491 ( .A(n48555), .B(n57726), .X(n36870) );
  nand_x1_sg U65492 ( .A(n57707), .B(n49789), .X(n36695) );
  nand_x1_sg U65493 ( .A(n52293), .B(n57758), .X(n36696) );
  nand_x1_sg U65494 ( .A(n52293), .B(n57682), .X(n36875) );
  nand_x1_sg U65495 ( .A(n48557), .B(n57746), .X(n36876) );
  nand_x1_sg U65496 ( .A(n57682), .B(n49787), .X(n36587) );
  nand_x1_sg U65497 ( .A(n52291), .B(n46201), .X(n36588) );
  nand_x1_sg U65498 ( .A(n52291), .B(n57716), .X(n36545) );
  nand_x1_sg U65499 ( .A(n48559), .B(n57742), .X(n36546) );
  nand_x1_sg U65500 ( .A(n52289), .B(n57680), .X(n36593) );
  nand_x1_sg U65501 ( .A(n48561), .B(n57743), .X(n36594) );
  nand_x1_sg U65502 ( .A(n52285), .B(n57708), .X(n36629) );
  nand_x1_sg U65503 ( .A(n48565), .B(n46200), .X(n36630) );
  nand_x1_sg U65504 ( .A(n57705), .B(n49779), .X(n37315) );
  nand_x1_sg U65505 ( .A(n52283), .B(n57755), .X(n37316) );
  nand_x1_sg U65506 ( .A(n52283), .B(n57696), .X(n36737) );
  nand_x1_sg U65507 ( .A(n48567), .B(n57762), .X(n36738) );
  nand_x1_sg U65508 ( .A(n57698), .B(n49777), .X(n37321) );
  nand_x1_sg U65509 ( .A(n52281), .B(n57727), .X(n37322) );
  nand_x1_sg U65510 ( .A(n52281), .B(n57693), .X(n36743) );
  nand_x1_sg U65511 ( .A(n48569), .B(n57741), .X(n36744) );
  nand_x1_sg U65512 ( .A(n52279), .B(n57704), .X(n36839) );
  nand_x1_sg U65513 ( .A(n48571), .B(n57747), .X(n36840) );
  nand_x1_sg U65514 ( .A(n52277), .B(n57709), .X(n36821) );
  nand_x1_sg U65515 ( .A(n48573), .B(n57755), .X(n36822) );
  nand_x1_sg U65516 ( .A(n52275), .B(n57706), .X(n36701) );
  nand_x1_sg U65517 ( .A(n48575), .B(n57734), .X(n36702) );
  nand_x1_sg U65518 ( .A(n52273), .B(n57707), .X(n36707) );
  nand_x1_sg U65519 ( .A(n48577), .B(n57737), .X(n36708) );
  nand_x1_sg U65520 ( .A(n52271), .B(n57717), .X(n36719) );
  nand_x1_sg U65521 ( .A(n48579), .B(n57750), .X(n36720) );
  nand_x1_sg U65522 ( .A(n52269), .B(n57718), .X(n36725) );
  nand_x1_sg U65523 ( .A(n48581), .B(n57742), .X(n36726) );
  nand_x1_sg U65524 ( .A(n52267), .B(n57643), .X(n36405) );
  nand_x1_sg U65525 ( .A(n48583), .B(n57764), .X(n36406) );
  nand_x1_sg U65526 ( .A(n52265), .B(n57634), .X(n36431) );
  nand_x1_sg U65527 ( .A(n48585), .B(n57757), .X(n36432) );
  nand_x1_sg U65528 ( .A(n57702), .B(n49745), .X(n37265) );
  nand_x1_sg U65529 ( .A(n52249), .B(n57757), .X(n37266) );
  nand_x1_sg U65530 ( .A(n57703), .B(n49741), .X(n37271) );
  nand_x1_sg U65531 ( .A(n52245), .B(n57773), .X(n37272) );
  nand_x1_sg U65532 ( .A(n57700), .B(n49739), .X(n37303) );
  nand_x1_sg U65533 ( .A(n52243), .B(n57755), .X(n37304) );
  nand_x1_sg U65534 ( .A(n52243), .B(n57682), .X(n37193) );
  nand_x1_sg U65535 ( .A(n48607), .B(n57743), .X(n37194) );
  nand_x1_sg U65536 ( .A(n57702), .B(n49737), .X(n37309) );
  nand_x1_sg U65537 ( .A(n52241), .B(n46201), .X(n37310) );
  nand_x1_sg U65538 ( .A(n52241), .B(n57682), .X(n37199) );
  nand_x1_sg U65539 ( .A(n48609), .B(n57765), .X(n37200) );
  nand_x1_sg U65540 ( .A(n57718), .B(n49735), .X(n36535) );
  nand_x1_sg U65541 ( .A(n52239), .B(n57742), .X(n36536) );
  nand_x1_sg U65542 ( .A(n52239), .B(n57706), .X(n37235) );
  nand_x1_sg U65543 ( .A(n48611), .B(n57746), .X(n37236) );
  nand_x1_sg U65544 ( .A(n57707), .B(n49733), .X(n36537) );
  nand_x1_sg U65545 ( .A(n52237), .B(n57742), .X(n36538) );
  nand_x1_sg U65546 ( .A(n52237), .B(n57697), .X(n37247) );
  nand_x1_sg U65547 ( .A(n48613), .B(n57743), .X(n37248) );
  nand_x1_sg U65548 ( .A(n57682), .B(n49731), .X(n37211) );
  nand_x1_sg U65549 ( .A(n52235), .B(n57764), .X(n37212) );
  nand_x1_sg U65550 ( .A(n52235), .B(n57717), .X(n37109) );
  nand_x1_sg U65551 ( .A(n48615), .B(n57735), .X(n37110) );
  nand_x1_sg U65552 ( .A(n57682), .B(n49729), .X(n37217) );
  nand_x1_sg U65553 ( .A(n52233), .B(n57743), .X(n37218) );
  nand_x1_sg U65554 ( .A(n52233), .B(n57699), .X(n37115) );
  nand_x1_sg U65555 ( .A(n48617), .B(n57729), .X(n37116) );
  nand_x1_sg U65556 ( .A(n57682), .B(n49727), .X(n37223) );
  nand_x1_sg U65557 ( .A(n52231), .B(n57746), .X(n37224) );
  nand_x1_sg U65558 ( .A(n52231), .B(n57703), .X(n37127) );
  nand_x1_sg U65559 ( .A(n48619), .B(n57728), .X(n37128) );
  nand_x1_sg U65560 ( .A(n57707), .B(n49725), .X(n37241) );
  nand_x1_sg U65561 ( .A(n52229), .B(n57765), .X(n37242) );
  nand_x1_sg U65562 ( .A(n52229), .B(n57682), .X(n37205) );
  nand_x1_sg U65563 ( .A(n48621), .B(n57743), .X(n37206) );
  nand_x1_sg U65564 ( .A(n57708), .B(n49723), .X(n37073) );
  nand_x1_sg U65565 ( .A(n52227), .B(n57755), .X(n37074) );
  nand_x1_sg U65566 ( .A(n52227), .B(n57682), .X(n37175) );
  nand_x1_sg U65567 ( .A(n48623), .B(n57728), .X(n37176) );
  nand_x1_sg U65568 ( .A(n57681), .B(n49721), .X(n37079) );
  nand_x1_sg U65569 ( .A(n52225), .B(n57730), .X(n37080) );
  nand_x1_sg U65570 ( .A(n52225), .B(n57682), .X(n37181) );
  nand_x1_sg U65571 ( .A(n48625), .B(n57757), .X(n37182) );
  nand_x1_sg U65572 ( .A(n57715), .B(n49719), .X(n37091) );
  nand_x1_sg U65573 ( .A(n52223), .B(n57730), .X(n37092) );
  nand_x1_sg U65574 ( .A(n52223), .B(n57700), .X(n37291) );
  nand_x1_sg U65575 ( .A(n48627), .B(n57760), .X(n37292) );
  nand_x1_sg U65576 ( .A(n57681), .B(n49717), .X(n37097) );
  nand_x1_sg U65577 ( .A(n52221), .B(n57741), .X(n37098) );
  nand_x1_sg U65578 ( .A(n52221), .B(n57693), .X(n37297) );
  nand_x1_sg U65579 ( .A(n48629), .B(n57748), .X(n37298) );
  nand_x1_sg U65580 ( .A(n57708), .B(n49715), .X(n37037) );
  nand_x1_sg U65581 ( .A(n52219), .B(n57759), .X(n37038) );
  nand_x1_sg U65582 ( .A(n52219), .B(n57695), .X(n37259) );
  nand_x1_sg U65583 ( .A(n48631), .B(n57728), .X(n37260) );
  nand_x1_sg U65584 ( .A(n57703), .B(n49713), .X(n37031) );
  nand_x1_sg U65585 ( .A(n52217), .B(n57759), .X(n37032) );
  nand_x1_sg U65586 ( .A(n57645), .B(n49711), .X(n36361) );
  nand_x1_sg U65587 ( .A(n52215), .B(n46201), .X(n36362) );
  nand_x1_sg U65588 ( .A(n57697), .B(n49709), .X(n37277) );
  nand_x1_sg U65589 ( .A(n52213), .B(n57756), .X(n37278) );
  nand_x1_sg U65590 ( .A(n52199), .B(n57679), .X(n37381) );
  nand_x1_sg U65591 ( .A(n48255), .B(n57724), .X(n37382) );
  nand_x1_sg U65592 ( .A(n57699), .B(n49691), .X(n37311) );
  nand_x1_sg U65593 ( .A(n52195), .B(n57755), .X(n37312) );
  nand_x1_sg U65594 ( .A(n57716), .B(n49689), .X(n37313) );
  nand_x1_sg U65595 ( .A(n52193), .B(n57743), .X(n37314) );
  nand_x1_sg U65596 ( .A(n57695), .B(n49687), .X(n37305) );
  nand_x1_sg U65597 ( .A(n52191), .B(n57755), .X(n37306) );
  nand_x1_sg U65598 ( .A(n57696), .B(n49685), .X(n37307) );
  nand_x1_sg U65599 ( .A(n52189), .B(n57754), .X(n37308) );
  nand_x1_sg U65600 ( .A(n57703), .B(n49683), .X(n37323) );
  nand_x1_sg U65601 ( .A(n52187), .B(n57727), .X(n37324) );
  nand_x1_sg U65602 ( .A(n57707), .B(n49681), .X(n37325) );
  nand_x1_sg U65603 ( .A(n52185), .B(n57727), .X(n37326) );
  nand_x1_sg U65604 ( .A(n57704), .B(n49679), .X(n37317) );
  nand_x1_sg U65605 ( .A(n52183), .B(n57755), .X(n37318) );
  nand_x1_sg U65606 ( .A(n57703), .B(n49677), .X(n37319) );
  nand_x1_sg U65607 ( .A(n52181), .B(n57727), .X(n37320) );
  nand_x1_sg U65608 ( .A(n57705), .B(n49675), .X(n37287) );
  nand_x1_sg U65609 ( .A(n52179), .B(n57766), .X(n37288) );
  nand_x1_sg U65610 ( .A(n57705), .B(n49673), .X(n37289) );
  nand_x1_sg U65611 ( .A(n52177), .B(n57757), .X(n37290) );
  nand_x1_sg U65612 ( .A(n57694), .B(n49671), .X(n37281) );
  nand_x1_sg U65613 ( .A(n52175), .B(n57772), .X(n37282) );
  nand_x1_sg U65614 ( .A(n57695), .B(n49669), .X(n37363) );
  nand_x1_sg U65615 ( .A(n52173), .B(n57725), .X(n37364) );
  nand_x1_sg U65616 ( .A(n52173), .B(n57704), .X(n37283) );
  nand_x1_sg U65617 ( .A(n48281), .B(n57765), .X(n37284) );
  nand_x1_sg U65618 ( .A(n52171), .B(n57693), .X(n37299) );
  nand_x1_sg U65619 ( .A(n48283), .B(n57750), .X(n37300) );
  nand_x1_sg U65620 ( .A(n52169), .B(n57694), .X(n37301) );
  nand_x1_sg U65621 ( .A(n48285), .B(n57762), .X(n37302) );
  nand_x1_sg U65622 ( .A(n52167), .B(n57699), .X(n37293) );
  nand_x1_sg U65623 ( .A(n48287), .B(n57770), .X(n37294) );
  nand_x1_sg U65624 ( .A(n52165), .B(n57700), .X(n37295) );
  nand_x1_sg U65625 ( .A(n48289), .B(n57747), .X(n37296) );
  nand_x1_sg U65626 ( .A(n52163), .B(n57679), .X(n37375) );
  nand_x1_sg U65627 ( .A(n48291), .B(n57724), .X(n37376) );
  nand_x1_sg U65628 ( .A(n52161), .B(n57679), .X(n37377) );
  nand_x1_sg U65629 ( .A(n48293), .B(n57724), .X(n37378) );
  nand_x1_sg U65630 ( .A(n52159), .B(n57696), .X(n37369) );
  nand_x1_sg U65631 ( .A(n48295), .B(n57724), .X(n37370) );
  nand_x1_sg U65632 ( .A(n52157), .B(n57679), .X(n37371) );
  nand_x1_sg U65633 ( .A(n48297), .B(n57724), .X(n37372) );
  nand_x1_sg U65634 ( .A(n52155), .B(n57679), .X(n37373) );
  nand_x1_sg U65635 ( .A(n48299), .B(n57724), .X(n37374) );
  nand_x1_sg U65636 ( .A(n52153), .B(n57679), .X(n37379) );
  nand_x1_sg U65637 ( .A(n48301), .B(n57724), .X(n37380) );
  nand_x1_sg U65638 ( .A(n52151), .B(n57693), .X(n37365) );
  nand_x1_sg U65639 ( .A(n48303), .B(n57725), .X(n37366) );
  nand_x1_sg U65640 ( .A(n52149), .B(n57694), .X(n37367) );
  nand_x1_sg U65641 ( .A(n48305), .B(n57724), .X(n37368) );
  nand_x1_sg U65642 ( .A(n52147), .B(n57707), .X(n37335) );
  nand_x1_sg U65643 ( .A(n48307), .B(n57726), .X(n37336) );
  nand_x1_sg U65644 ( .A(n52145), .B(n57704), .X(n37337) );
  nand_x1_sg U65645 ( .A(n48309), .B(n57726), .X(n37338) );
  nand_x1_sg U65646 ( .A(n52143), .B(n57694), .X(n37329) );
  nand_x1_sg U65647 ( .A(n48311), .B(n57727), .X(n37330) );
  nand_x1_sg U65648 ( .A(n52141), .B(n57701), .X(n37331) );
  nand_x1_sg U65649 ( .A(n48313), .B(n57727), .X(n37332) );
  nand_x1_sg U65650 ( .A(n52139), .B(n57718), .X(n37359) );
  nand_x1_sg U65651 ( .A(n48315), .B(n57725), .X(n37360) );
  nand_x1_sg U65652 ( .A(n52137), .B(n57702), .X(n37333) );
  nand_x1_sg U65653 ( .A(n48317), .B(n57727), .X(n37334) );
  nand_x1_sg U65654 ( .A(n52135), .B(n57717), .X(n37361) );
  nand_x1_sg U65655 ( .A(n48319), .B(n57725), .X(n37362) );
  nand_x1_sg U65656 ( .A(n57699), .B(n49589), .X(n37005) );
  nand_x1_sg U65657 ( .A(n52093), .B(n57733), .X(n37006) );
  nand_x1_sg U65658 ( .A(n57708), .B(n49587), .X(n37069) );
  nand_x1_sg U65659 ( .A(n52091), .B(n57734), .X(n37070) );
  nand_x1_sg U65660 ( .A(n57634), .B(n49585), .X(n37071) );
  nand_x1_sg U65661 ( .A(n52089), .B(n57730), .X(n37072) );
  nand_x1_sg U65662 ( .A(n57681), .B(n49583), .X(n37063) );
  nand_x1_sg U65663 ( .A(n52087), .B(n57731), .X(n37064) );
  nand_x1_sg U65664 ( .A(n57682), .B(n49581), .X(n37065) );
  nand_x1_sg U65665 ( .A(n52085), .B(n57736), .X(n37066) );
  nand_x1_sg U65666 ( .A(n57709), .B(n49579), .X(n37081) );
  nand_x1_sg U65667 ( .A(n52083), .B(n57730), .X(n37082) );
  nand_x1_sg U65668 ( .A(n52083), .B(n57703), .X(n37021) );
  nand_x1_sg U65669 ( .A(n48371), .B(n57732), .X(n37022) );
  nand_x1_sg U65670 ( .A(n57717), .B(n49577), .X(n37083) );
  nand_x1_sg U65671 ( .A(n52081), .B(n57730), .X(n37084) );
  nand_x1_sg U65672 ( .A(n52081), .B(n57697), .X(n37023) );
  nand_x1_sg U65673 ( .A(n48373), .B(n57732), .X(n37024) );
  nand_x1_sg U65674 ( .A(n57720), .B(n49575), .X(n37075) );
  nand_x1_sg U65675 ( .A(n52079), .B(n57739), .X(n37076) );
  nand_x1_sg U65676 ( .A(n52079), .B(n57720), .X(n37015) );
  nand_x1_sg U65677 ( .A(n48375), .B(n57732), .X(n37016) );
  nand_x1_sg U65678 ( .A(n57709), .B(n49573), .X(n37077) );
  nand_x1_sg U65679 ( .A(n52077), .B(n57738), .X(n37078) );
  nand_x1_sg U65680 ( .A(n52077), .B(n57709), .X(n37017) );
  nand_x1_sg U65681 ( .A(n48377), .B(n57732), .X(n37018) );
  nand_x1_sg U65682 ( .A(n57709), .B(n49571), .X(n37045) );
  nand_x1_sg U65683 ( .A(n52075), .B(n57733), .X(n37046) );
  nand_x1_sg U65684 ( .A(n52075), .B(n57720), .X(n37033) );
  nand_x1_sg U65685 ( .A(n48379), .B(n57759), .X(n37034) );
  nand_x1_sg U65686 ( .A(n57716), .B(n49569), .X(n37047) );
  nand_x1_sg U65687 ( .A(n52073), .B(n57731), .X(n37048) );
  nand_x1_sg U65688 ( .A(n52073), .B(n57718), .X(n37035) );
  nand_x1_sg U65689 ( .A(n48381), .B(n57759), .X(n37036) );
  nand_x1_sg U65690 ( .A(n57717), .B(n49567), .X(n37039) );
  nand_x1_sg U65691 ( .A(n52071), .B(n57759), .X(n37040) );
  nand_x1_sg U65692 ( .A(n52071), .B(n57695), .X(n37027) );
  nand_x1_sg U65693 ( .A(n48383), .B(n57732), .X(n37028) );
  nand_x1_sg U65694 ( .A(n57715), .B(n49565), .X(n37041) );
  nand_x1_sg U65695 ( .A(n52069), .B(n57759), .X(n37042) );
  nand_x1_sg U65696 ( .A(n52069), .B(n57696), .X(n37029) );
  nand_x1_sg U65697 ( .A(n48385), .B(n57732), .X(n37030) );
  nand_x1_sg U65698 ( .A(n57680), .B(n49563), .X(n37057) );
  nand_x1_sg U65699 ( .A(n52067), .B(n57731), .X(n37058) );
  nand_x1_sg U65700 ( .A(n52067), .B(n57700), .X(n36997) );
  nand_x1_sg U65701 ( .A(n48387), .B(n57734), .X(n36998) );
  nand_x1_sg U65702 ( .A(n57715), .B(n49561), .X(n37059) );
  nand_x1_sg U65703 ( .A(n52065), .B(n57731), .X(n37060) );
  nand_x1_sg U65704 ( .A(n52065), .B(n57718), .X(n36999) );
  nand_x1_sg U65705 ( .A(n48389), .B(n57733), .X(n37000) );
  nand_x1_sg U65706 ( .A(n57634), .B(n49559), .X(n37051) );
  nand_x1_sg U65707 ( .A(n52063), .B(n57731), .X(n37052) );
  nand_x1_sg U65708 ( .A(n52063), .B(n57703), .X(n36991) );
  nand_x1_sg U65709 ( .A(n48391), .B(n57734), .X(n36992) );
  nand_x1_sg U65710 ( .A(n57697), .B(n49557), .X(n37053) );
  nand_x1_sg U65711 ( .A(n52061), .B(n57731), .X(n37054) );
  nand_x1_sg U65712 ( .A(n52061), .B(n57703), .X(n36993) );
  nand_x1_sg U65713 ( .A(n48393), .B(n57734), .X(n36994) );
  nand_x1_sg U65714 ( .A(n57702), .B(n49555), .X(n36925) );
  nand_x1_sg U65715 ( .A(n52059), .B(n57737), .X(n36926) );
  nand_x1_sg U65716 ( .A(n52059), .B(n57716), .X(n37009) );
  nand_x1_sg U65717 ( .A(n48395), .B(n57733), .X(n37010) );
  nand_x1_sg U65718 ( .A(n57716), .B(n49553), .X(n36927) );
  nand_x1_sg U65719 ( .A(n52057), .B(n57737), .X(n36928) );
  nand_x1_sg U65720 ( .A(n52057), .B(n57681), .X(n37011) );
  nand_x1_sg U65721 ( .A(n48397), .B(n57733), .X(n37012) );
  nand_x1_sg U65722 ( .A(n57702), .B(n49551), .X(n36919) );
  nand_x1_sg U65723 ( .A(n52055), .B(n57737), .X(n36920) );
  nand_x1_sg U65724 ( .A(n52055), .B(n57708), .X(n37003) );
  nand_x1_sg U65725 ( .A(n48399), .B(n57733), .X(n37004) );
  nand_x1_sg U65726 ( .A(n57703), .B(n49549), .X(n36985) );
  nand_x1_sg U65727 ( .A(n52053), .B(n57734), .X(n36986) );
  nand_x1_sg U65728 ( .A(n52053), .B(n57699), .X(n36921) );
  nand_x1_sg U65729 ( .A(n48401), .B(n57737), .X(n36922) );
  nand_x1_sg U65730 ( .A(n57706), .B(n49547), .X(n36987) );
  nand_x1_sg U65731 ( .A(n52051), .B(n57734), .X(n36988) );
  nand_x1_sg U65732 ( .A(n52051), .B(n57695), .X(n36937) );
  nand_x1_sg U65733 ( .A(n48403), .B(n57736), .X(n36938) );
  nand_x1_sg U65734 ( .A(n57716), .B(n49545), .X(n36979) );
  nand_x1_sg U65735 ( .A(n52049), .B(n57761), .X(n36980) );
  nand_x1_sg U65736 ( .A(n52049), .B(n57696), .X(n36939) );
  nand_x1_sg U65737 ( .A(n48405), .B(n57736), .X(n36940) );
  nand_x1_sg U65738 ( .A(n57695), .B(n49543), .X(n36981) );
  nand_x1_sg U65739 ( .A(n52047), .B(n57761), .X(n36982) );
  nand_x1_sg U65740 ( .A(n52047), .B(n57680), .X(n36931) );
  nand_x1_sg U65741 ( .A(n48407), .B(n57737), .X(n36932) );
  nand_x1_sg U65742 ( .A(n57709), .B(n49541), .X(n36949) );
  nand_x1_sg U65743 ( .A(n52045), .B(n57736), .X(n36950) );
  nand_x1_sg U65744 ( .A(n52045), .B(n57708), .X(n36933) );
  nand_x1_sg U65745 ( .A(n48409), .B(n57737), .X(n36934) );
  nand_x1_sg U65746 ( .A(n57708), .B(n49539), .X(n36951) );
  nand_x1_sg U65747 ( .A(n52043), .B(n57735), .X(n36952) );
  nand_x1_sg U65748 ( .A(n52043), .B(n57699), .X(n36901) );
  nand_x1_sg U65749 ( .A(n48411), .B(n57739), .X(n36902) );
  nand_x1_sg U65750 ( .A(n57693), .B(n49537), .X(n36943) );
  nand_x1_sg U65751 ( .A(n52041), .B(n57736), .X(n36944) );
  nand_x1_sg U65752 ( .A(n52041), .B(n57700), .X(n36903) );
  nand_x1_sg U65753 ( .A(n48413), .B(n57738), .X(n36904) );
  nand_x1_sg U65754 ( .A(n57701), .B(n49535), .X(n36945) );
  nand_x1_sg U65755 ( .A(n52039), .B(n57736), .X(n36946) );
  nand_x1_sg U65756 ( .A(n52039), .B(n57698), .X(n36895) );
  nand_x1_sg U65757 ( .A(n48415), .B(n57739), .X(n36896) );
  nand_x1_sg U65758 ( .A(n57701), .B(n49533), .X(n36961) );
  nand_x1_sg U65759 ( .A(n52037), .B(n57735), .X(n36962) );
  nand_x1_sg U65760 ( .A(n52037), .B(n57697), .X(n36897) );
  nand_x1_sg U65761 ( .A(n48417), .B(n57739), .X(n36898) );
  nand_x1_sg U65762 ( .A(n57706), .B(n49531), .X(n36963) );
  nand_x1_sg U65763 ( .A(n52035), .B(n57735), .X(n36964) );
  nand_x1_sg U65764 ( .A(n52035), .B(n57700), .X(n36913) );
  nand_x1_sg U65765 ( .A(n48419), .B(n57738), .X(n36914) );
  nand_x1_sg U65766 ( .A(n57706), .B(n49529), .X(n36955) );
  nand_x1_sg U65767 ( .A(n52033), .B(n57735), .X(n36956) );
  nand_x1_sg U65768 ( .A(n52033), .B(n57698), .X(n36915) );
  nand_x1_sg U65769 ( .A(n48421), .B(n57738), .X(n36916) );
  nand_x1_sg U65770 ( .A(n57708), .B(n49527), .X(n36957) );
  nand_x1_sg U65771 ( .A(n52031), .B(n57735), .X(n36958) );
  nand_x1_sg U65772 ( .A(n52031), .B(n57697), .X(n36907) );
  nand_x1_sg U65773 ( .A(n48423), .B(n57738), .X(n36908) );
  nand_x1_sg U65774 ( .A(n57682), .B(n49525), .X(n37213) );
  nand_x1_sg U65775 ( .A(n52029), .B(n57765), .X(n37214) );
  nand_x1_sg U65776 ( .A(n52029), .B(n57705), .X(n36909) );
  nand_x1_sg U65777 ( .A(n48425), .B(n57738), .X(n36910) );
  nand_x1_sg U65778 ( .A(n57682), .B(n49523), .X(n37215) );
  nand_x1_sg U65779 ( .A(n52027), .B(n57771), .X(n37216) );
  nand_x1_sg U65780 ( .A(n52027), .B(n57707), .X(n36973) );
  nand_x1_sg U65781 ( .A(n48427), .B(n57739), .X(n36974) );
  nand_x1_sg U65782 ( .A(n57682), .B(n49521), .X(n37207) );
  nand_x1_sg U65783 ( .A(n52025), .B(n57761), .X(n37208) );
  nand_x1_sg U65784 ( .A(n52025), .B(n57704), .X(n36975) );
  nand_x1_sg U65785 ( .A(n48429), .B(n57761), .X(n36976) );
  nand_x1_sg U65786 ( .A(n57682), .B(n49519), .X(n37209) );
  nand_x1_sg U65787 ( .A(n52023), .B(n46201), .X(n37210) );
  nand_x1_sg U65788 ( .A(n52023), .B(n57705), .X(n36967) );
  nand_x1_sg U65789 ( .A(n48431), .B(n57761), .X(n36968) );
  nand_x1_sg U65790 ( .A(n57682), .B(n49517), .X(n37225) );
  nand_x1_sg U65791 ( .A(n52021), .B(n57746), .X(n37226) );
  nand_x1_sg U65792 ( .A(n52021), .B(n57696), .X(n36969) );
  nand_x1_sg U65793 ( .A(n48433), .B(n57761), .X(n36970) );
  nand_x1_sg U65794 ( .A(n52019), .B(n57682), .X(n37189) );
  nand_x1_sg U65795 ( .A(n48039), .B(n57728), .X(n37190) );
  nand_x1_sg U65796 ( .A(n57696), .B(n49513), .X(n37251) );
  nand_x1_sg U65797 ( .A(n52017), .B(n57743), .X(n37252) );
  nand_x1_sg U65798 ( .A(n52017), .B(n57682), .X(n37191) );
  nand_x1_sg U65799 ( .A(n48041), .B(n57762), .X(n37192) );
  nand_x1_sg U65800 ( .A(n57706), .B(n49511), .X(n37243) );
  nand_x1_sg U65801 ( .A(n52015), .B(n57743), .X(n37244) );
  nand_x1_sg U65802 ( .A(n52015), .B(n57682), .X(n37183) );
  nand_x1_sg U65803 ( .A(n48043), .B(n57746), .X(n37184) );
  nand_x1_sg U65804 ( .A(n57707), .B(n49509), .X(n37245) );
  nand_x1_sg U65805 ( .A(n52013), .B(n57743), .X(n37246) );
  nand_x1_sg U65806 ( .A(n52013), .B(n57682), .X(n37185) );
  nand_x1_sg U65807 ( .A(n48045), .B(n57742), .X(n37186) );
  nand_x1_sg U65808 ( .A(n57718), .B(n49507), .X(n37117) );
  nand_x1_sg U65809 ( .A(n52011), .B(n57729), .X(n37118) );
  nand_x1_sg U65810 ( .A(n52011), .B(n57682), .X(n37201) );
  nand_x1_sg U65811 ( .A(n48047), .B(n57763), .X(n37202) );
  nand_x1_sg U65812 ( .A(n57681), .B(n49505), .X(n37119) );
  nand_x1_sg U65813 ( .A(n52009), .B(n57729), .X(n37120) );
  nand_x1_sg U65814 ( .A(n52009), .B(n57682), .X(n37203) );
  nand_x1_sg U65815 ( .A(n48049), .B(n57765), .X(n37204) );
  nand_x1_sg U65816 ( .A(n57682), .B(n49503), .X(n37111) );
  nand_x1_sg U65817 ( .A(n52007), .B(n57729), .X(n37112) );
  nand_x1_sg U65818 ( .A(n52007), .B(n57682), .X(n37195) );
  nand_x1_sg U65819 ( .A(n48051), .B(n57743), .X(n37196) );
  nand_x1_sg U65820 ( .A(n57680), .B(n49501), .X(n37113) );
  nand_x1_sg U65821 ( .A(n52005), .B(n57729), .X(n37114) );
  nand_x1_sg U65822 ( .A(n52005), .B(n57682), .X(n37197) );
  nand_x1_sg U65823 ( .A(n48053), .B(n57744), .X(n37198) );
  nand_x1_sg U65824 ( .A(n57705), .B(n49499), .X(n37129) );
  nand_x1_sg U65825 ( .A(n52003), .B(n46201), .X(n37130) );
  nand_x1_sg U65826 ( .A(n52003), .B(n57693), .X(n37261) );
  nand_x1_sg U65827 ( .A(n48055), .B(n57728), .X(n37262) );
  nand_x1_sg U65828 ( .A(n57701), .B(n49497), .X(n37131) );
  nand_x1_sg U65829 ( .A(n52001), .B(n46197), .X(n37132) );
  nand_x1_sg U65830 ( .A(n52001), .B(n57694), .X(n37263) );
  nand_x1_sg U65831 ( .A(n48057), .B(n57728), .X(n37264) );
  nand_x1_sg U65832 ( .A(n57701), .B(n49495), .X(n37123) );
  nand_x1_sg U65833 ( .A(n51999), .B(n57729), .X(n37124) );
  nand_x1_sg U65834 ( .A(n51999), .B(n57717), .X(n37255) );
  nand_x1_sg U65835 ( .A(n48059), .B(n57757), .X(n37256) );
  nand_x1_sg U65836 ( .A(n57708), .B(n49493), .X(n37125) );
  nand_x1_sg U65837 ( .A(n51997), .B(n57729), .X(n37126) );
  nand_x1_sg U65838 ( .A(n51997), .B(n57697), .X(n37257) );
  nand_x1_sg U65839 ( .A(n48061), .B(n57757), .X(n37258) );
  nand_x1_sg U65840 ( .A(n57708), .B(n49491), .X(n37093) );
  nand_x1_sg U65841 ( .A(n51995), .B(n57730), .X(n37094) );
  nand_x1_sg U65842 ( .A(n51995), .B(n57701), .X(n37273) );
  nand_x1_sg U65843 ( .A(n48063), .B(n57746), .X(n37274) );
  nand_x1_sg U65844 ( .A(n57701), .B(n49489), .X(n37095) );
  nand_x1_sg U65845 ( .A(n51993), .B(n57732), .X(n37096) );
  nand_x1_sg U65846 ( .A(n51993), .B(n57698), .X(n37275) );
  nand_x1_sg U65847 ( .A(n48065), .B(n57742), .X(n37276) );
  nand_x1_sg U65848 ( .A(n57634), .B(n49487), .X(n37087) );
  nand_x1_sg U65849 ( .A(n51991), .B(n57730), .X(n37088) );
  nand_x1_sg U65850 ( .A(n51991), .B(n57705), .X(n37267) );
  nand_x1_sg U65851 ( .A(n48067), .B(n57757), .X(n37268) );
  nand_x1_sg U65852 ( .A(n57716), .B(n49485), .X(n37089) );
  nand_x1_sg U65853 ( .A(n51989), .B(n57730), .X(n37090) );
  nand_x1_sg U65854 ( .A(n51989), .B(n57708), .X(n37269) );
  nand_x1_sg U65855 ( .A(n48069), .B(n57728), .X(n37270) );
  nand_x1_sg U65856 ( .A(n57680), .B(n49483), .X(n37105) );
  nand_x1_sg U65857 ( .A(n51987), .B(n57743), .X(n37106) );
  nand_x1_sg U65858 ( .A(n51987), .B(n57708), .X(n37237) );
  nand_x1_sg U65859 ( .A(n48071), .B(n57746), .X(n37238) );
  nand_x1_sg U65860 ( .A(n57682), .B(n49481), .X(n37107) );
  nand_x1_sg U65861 ( .A(n51985), .B(n57772), .X(n37108) );
  nand_x1_sg U65862 ( .A(n51985), .B(n57709), .X(n37239) );
  nand_x1_sg U65863 ( .A(n48073), .B(n57765), .X(n37240) );
  nand_x1_sg U65864 ( .A(n57717), .B(n49479), .X(n37099) );
  nand_x1_sg U65865 ( .A(n51983), .B(n46200), .X(n37100) );
  nand_x1_sg U65866 ( .A(n51983), .B(n57704), .X(n37231) );
  nand_x1_sg U65867 ( .A(n48075), .B(n57746), .X(n37232) );
  nand_x1_sg U65868 ( .A(n57682), .B(n49477), .X(n37101) );
  nand_x1_sg U65869 ( .A(n51981), .B(n46198), .X(n37102) );
  nand_x1_sg U65870 ( .A(n51981), .B(n57704), .X(n37233) );
  nand_x1_sg U65871 ( .A(n48077), .B(n57746), .X(n37234) );
  nand_x1_sg U65872 ( .A(n57682), .B(n49475), .X(n37165) );
  nand_x1_sg U65873 ( .A(n51979), .B(n57746), .X(n37166) );
  nand_x1_sg U65874 ( .A(n51979), .B(n57695), .X(n37249) );
  nand_x1_sg U65875 ( .A(n48079), .B(n57743), .X(n37250) );
  nand_x1_sg U65876 ( .A(n57715), .B(n49473), .X(n36959) );
  nand_x1_sg U65877 ( .A(n51977), .B(n57735), .X(n36960) );
  nand_x1_sg U65878 ( .A(n51977), .B(n57682), .X(n37167) );
  nand_x1_sg U65879 ( .A(n48081), .B(n57766), .X(n37168) );
  nand_x1_sg U65880 ( .A(n51975), .B(n57682), .X(n37159) );
  nand_x1_sg U65881 ( .A(n48083), .B(n57746), .X(n37160) );
  nand_x1_sg U65882 ( .A(n51973), .B(n57682), .X(n37161) );
  nand_x1_sg U65883 ( .A(n48085), .B(n57766), .X(n37162) );
  nand_x1_sg U65884 ( .A(n51971), .B(n57682), .X(n37177) );
  nand_x1_sg U65885 ( .A(n48087), .B(n57766), .X(n37178) );
  nand_x1_sg U65886 ( .A(n57708), .B(n49465), .X(n36953) );
  nand_x1_sg U65887 ( .A(n51969), .B(n57735), .X(n36954) );
  nand_x1_sg U65888 ( .A(n51969), .B(n57682), .X(n37179) );
  nand_x1_sg U65889 ( .A(n48089), .B(n57757), .X(n37180) );
  nand_x1_sg U65890 ( .A(n51967), .B(n57682), .X(n37171) );
  nand_x1_sg U65891 ( .A(n48091), .B(n57746), .X(n37172) );
  nand_x1_sg U65892 ( .A(n51965), .B(n57682), .X(n37173) );
  nand_x1_sg U65893 ( .A(n48093), .B(n57766), .X(n37174) );
  nand_x1_sg U65894 ( .A(n51963), .B(n57693), .X(n37141) );
  nand_x1_sg U65895 ( .A(n48095), .B(n57733), .X(n37142) );
  nand_x1_sg U65896 ( .A(n51961), .B(n57694), .X(n37143) );
  nand_x1_sg U65897 ( .A(n48097), .B(n57728), .X(n37144) );
  nand_x1_sg U65898 ( .A(n51959), .B(n57702), .X(n37135) );
  nand_x1_sg U65899 ( .A(n48099), .B(n57760), .X(n37136) );
  nand_x1_sg U65900 ( .A(n51957), .B(n57706), .X(n37137) );
  nand_x1_sg U65901 ( .A(n48101), .B(n57749), .X(n37138) );
  nand_x1_sg U65902 ( .A(n51955), .B(n57715), .X(n37153) );
  nand_x1_sg U65903 ( .A(n48103), .B(n57728), .X(n37154) );
  nand_x1_sg U65904 ( .A(n51953), .B(n57708), .X(n37155) );
  nand_x1_sg U65905 ( .A(n48105), .B(n57728), .X(n37156) );
  nand_x1_sg U65906 ( .A(n51951), .B(n57680), .X(n37147) );
  nand_x1_sg U65907 ( .A(n48107), .B(n57728), .X(n37148) );
  nand_x1_sg U65908 ( .A(n57703), .B(n49445), .X(n36977) );
  nand_x1_sg U65909 ( .A(n51949), .B(n57737), .X(n36978) );
  nand_x1_sg U65910 ( .A(n51949), .B(n57634), .X(n37149) );
  nand_x1_sg U65911 ( .A(n48109), .B(n57728), .X(n37150) );
  nand_x1_sg U65912 ( .A(n57695), .B(n49425), .X(n36923) );
  nand_x1_sg U65913 ( .A(n51929), .B(n57737), .X(n36924) );
  nand_x1_sg U65914 ( .A(n57694), .B(n49419), .X(n36941) );
  nand_x1_sg U65915 ( .A(n51923), .B(n57736), .X(n36942) );
  nand_x1_sg U65916 ( .A(n57709), .B(n49417), .X(n36947) );
  nand_x1_sg U65917 ( .A(n51921), .B(n57736), .X(n36948) );
  nand_x1_sg U65918 ( .A(n57715), .B(n49379), .X(n36513) );
  nand_x1_sg U65919 ( .A(n51883), .B(n57755), .X(n36514) );
  nand_x1_sg U65920 ( .A(n57644), .B(n49335), .X(n36373) );
  nand_x1_sg U65921 ( .A(n51839), .B(n46197), .X(n36374) );
  nand_x1_sg U65922 ( .A(n57707), .B(n49327), .X(n37133) );
  nand_x1_sg U65923 ( .A(n51831), .B(n57764), .X(n37134) );
  nand_x1_sg U65924 ( .A(n57682), .B(n49323), .X(n37169) );
  nand_x1_sg U65925 ( .A(n51827), .B(n57766), .X(n37170) );
  nand_x1_sg U65926 ( .A(n57696), .B(n49321), .X(n37253) );
  nand_x1_sg U65927 ( .A(n51825), .B(n57743), .X(n37254) );
  nand_x1_sg U65928 ( .A(n57709), .B(n49319), .X(n37151) );
  nand_x1_sg U65929 ( .A(n51823), .B(n57728), .X(n37152) );
  nand_x1_sg U65930 ( .A(n57708), .B(n49317), .X(n36541) );
  nand_x1_sg U65931 ( .A(n51821), .B(n57742), .X(n36542) );
  nand_x1_sg U65932 ( .A(n51821), .B(n57645), .X(n36363) );
  nand_x1_sg U65933 ( .A(n47841), .B(n57772), .X(n36364) );
  nand_x1_sg U65934 ( .A(n57709), .B(n49315), .X(n36809) );
  nand_x1_sg U65935 ( .A(n51819), .B(n57747), .X(n36810) );
  nand_x1_sg U65936 ( .A(n57682), .B(n49313), .X(n36803) );
  nand_x1_sg U65937 ( .A(n51817), .B(n57758), .X(n36804) );
  nand_x1_sg U65938 ( .A(n57715), .B(n49311), .X(n36543) );
  nand_x1_sg U65939 ( .A(n51815), .B(n57742), .X(n36544) );
  nand_x1_sg U65940 ( .A(n57701), .B(n49307), .X(n36899) );
  nand_x1_sg U65941 ( .A(n51811), .B(n57739), .X(n36900) );
  nand_x1_sg U65942 ( .A(n57696), .B(n49305), .X(n36911) );
  nand_x1_sg U65943 ( .A(n51809), .B(n57738), .X(n36912) );
  nand_x1_sg U65944 ( .A(n57702), .B(n49303), .X(n36893) );
  nand_x1_sg U65945 ( .A(n51807), .B(n57739), .X(n36894) );
  nand_x1_sg U65946 ( .A(n57634), .B(n49301), .X(n37085) );
  nand_x1_sg U65947 ( .A(n51805), .B(n57730), .X(n37086) );
  nand_x1_sg U65948 ( .A(n51803), .B(n57682), .X(n37187) );
  nand_x1_sg U65949 ( .A(n47859), .B(n57728), .X(n37188) );
  nand_x1_sg U65950 ( .A(n51801), .B(n57680), .X(n37121) );
  nand_x1_sg U65951 ( .A(n47861), .B(n57729), .X(n37122) );
  nand_x1_sg U65952 ( .A(n57682), .B(n49295), .X(n36539) );
  nand_x1_sg U65953 ( .A(n51799), .B(n57742), .X(n36540) );
  nand_x1_sg U65954 ( .A(n51795), .B(n57699), .X(n37229) );
  nand_x1_sg U65955 ( .A(n47867), .B(n57746), .X(n37230) );
  nand_x1_sg U65956 ( .A(n57645), .B(n49289), .X(n36365) );
  nand_x1_sg U65957 ( .A(n51793), .B(n46200), .X(n36366) );
  nand_x1_sg U65958 ( .A(n51791), .B(n57720), .X(n37103) );
  nand_x1_sg U65959 ( .A(n47871), .B(n57740), .X(n37104) );
  nand_x1_sg U65960 ( .A(n57702), .B(n49281), .X(n37279) );
  nand_x1_sg U65961 ( .A(n51785), .B(n57750), .X(n37280) );
  nand_x1_sg U65962 ( .A(n51785), .B(n57717), .X(n36599) );
  nand_x1_sg U65963 ( .A(n47877), .B(n57772), .X(n36600) );
  nand_x1_sg U65964 ( .A(n57680), .B(n49279), .X(n36881) );
  nand_x1_sg U65965 ( .A(n51783), .B(n46198), .X(n36882) );
  nand_x1_sg U65966 ( .A(n51783), .B(n57694), .X(n37067) );
  nand_x1_sg U65967 ( .A(n47879), .B(n57739), .X(n37068) );
  nand_x1_sg U65968 ( .A(n51781), .B(n57693), .X(n37019) );
  nand_x1_sg U65969 ( .A(n47881), .B(n57732), .X(n37020) );
  nand_x1_sg U65970 ( .A(n51779), .B(n57720), .X(n36929) );
  nand_x1_sg U65971 ( .A(n47883), .B(n57737), .X(n36930) );
  nand_x1_sg U65972 ( .A(n57698), .B(n49273), .X(n37285) );
  nand_x1_sg U65973 ( .A(n51777), .B(n57744), .X(n37286) );
  nand_x1_sg U65974 ( .A(n51777), .B(n57708), .X(n36965) );
  nand_x1_sg U65975 ( .A(n47885), .B(n57735), .X(n36966) );
  nand_x1_sg U65976 ( .A(n57720), .B(n49271), .X(n36533) );
  nand_x1_sg U65977 ( .A(n51775), .B(n57742), .X(n36534) );
  nand_x1_sg U65978 ( .A(n51775), .B(n57705), .X(n36845) );
  nand_x1_sg U65979 ( .A(n47887), .B(n57763), .X(n36846) );
  nand_x1_sg U65980 ( .A(n51771), .B(n57681), .X(n36827) );
  nand_x1_sg U65981 ( .A(n47891), .B(n57765), .X(n36828) );
  nand_x1_sg U65982 ( .A(n51769), .B(n57701), .X(n36563) );
  nand_x1_sg U65983 ( .A(n47893), .B(n57742), .X(n36564) );
  nand_x1_sg U65984 ( .A(n51765), .B(n57634), .X(n36731) );
  nand_x1_sg U65985 ( .A(n47897), .B(n57772), .X(n36732) );
  nand_x1_sg U65986 ( .A(n57701), .B(n51755), .X(n36995) );
  nand_x1_sg U65987 ( .A(n47907), .B(n57734), .X(n36996) );
  nand_x1_sg U65988 ( .A(n51753), .B(n57680), .X(n37001) );
  nand_x1_sg U65989 ( .A(n47909), .B(n57733), .X(n37002) );
  nand_x1_sg U65990 ( .A(n51745), .B(n57706), .X(n37327) );
  nand_x1_sg U65991 ( .A(n47917), .B(n57727), .X(n37328) );
  nand_x1_sg U65992 ( .A(n57693), .B(n49237), .X(n36917) );
  nand_x1_sg U65993 ( .A(n51741), .B(n57738), .X(n36918) );
  nand_x1_sg U65994 ( .A(n57699), .B(n49229), .X(n36935) );
  nand_x1_sg U65995 ( .A(n51733), .B(n57736), .X(n36936) );
  nand_x1_sg U65996 ( .A(n57709), .B(n49221), .X(n36971) );
  nand_x1_sg U65997 ( .A(n51725), .B(n57737), .X(n36972) );
  nand_x1_sg U65998 ( .A(n57700), .B(n49219), .X(n36989) );
  nand_x1_sg U65999 ( .A(n51723), .B(n57734), .X(n36990) );
  nand_x1_sg U66000 ( .A(n57698), .B(n49215), .X(n36983) );
  nand_x1_sg U66001 ( .A(n51719), .B(n57734), .X(n36984) );
  nand_x1_sg U66002 ( .A(n57716), .B(n49213), .X(n37049) );
  nand_x1_sg U66003 ( .A(n51717), .B(n57731), .X(n37050) );
  nand_x1_sg U66004 ( .A(n51703), .B(n57694), .X(n36905) );
  nand_x1_sg U66005 ( .A(n47959), .B(n57738), .X(n36906) );
  nand_x1_sg U66006 ( .A(n57694), .B(n49149), .X(n36749) );
  nand_x1_sg U66007 ( .A(n51653), .B(n57741), .X(n36750) );
  nand_x1_sg U66008 ( .A(n57634), .B(n49147), .X(n36785) );
  nand_x1_sg U66009 ( .A(n51651), .B(n57743), .X(n36786) );
  nand_x1_sg U66010 ( .A(n57681), .B(n49143), .X(n36773) );
  nand_x1_sg U66011 ( .A(n51647), .B(n57740), .X(n36774) );
  nand_x1_sg U66012 ( .A(n57709), .B(n49139), .X(n36857) );
  nand_x1_sg U66013 ( .A(n51643), .B(n57727), .X(n36858) );
  nand_x1_sg U66014 ( .A(n57704), .B(n49137), .X(n36683) );
  nand_x1_sg U66015 ( .A(n51641), .B(n57762), .X(n36684) );
  nand_x1_sg U66016 ( .A(n57702), .B(n49135), .X(n36635) );
  nand_x1_sg U66017 ( .A(n51639), .B(n57761), .X(n36636) );
  nand_x1_sg U66018 ( .A(n57706), .B(n49131), .X(n36437) );
  nand_x1_sg U66019 ( .A(n51635), .B(n57766), .X(n36438) );
  nand_x1_sg U66020 ( .A(n57680), .B(n49129), .X(n36611) );
  nand_x1_sg U66021 ( .A(n51633), .B(n46198), .X(n36612) );
  nand_x1_sg U66022 ( .A(n57709), .B(n49127), .X(n36623) );
  nand_x1_sg U66023 ( .A(n51631), .B(n46198), .X(n36624) );
  nand_x1_sg U66024 ( .A(n57706), .B(n49123), .X(n36641) );
  nand_x1_sg U66025 ( .A(n51627), .B(n57734), .X(n36642) );
  nand_x1_sg U66026 ( .A(n53095), .B(n57870), .X(n30606) );
  nand_x1_sg U66027 ( .A(n51549), .B(n57886), .X(n30607) );
  nand_x1_sg U66028 ( .A(n50747), .B(n57880), .X(n29470) );
  nand_x1_sg U66029 ( .A(n57025), .B(n57888), .X(n29471) );
  nand_x1_sg U66030 ( .A(n53273), .B(n57880), .X(n29464) );
  nand_x1_sg U66031 ( .A(n51501), .B(n57892), .X(n29465) );
  nand_x1_sg U66032 ( .A(n53271), .B(n57876), .X(n29452) );
  nand_x1_sg U66033 ( .A(n47755), .B(n57903), .X(n29453) );
  nand_x1_sg U66034 ( .A(n50741), .B(n57876), .X(n29440) );
  nand_x1_sg U66035 ( .A(n57035), .B(n57903), .X(n29441) );
  nand_x1_sg U66036 ( .A(n53269), .B(n57877), .X(n29428) );
  nand_x1_sg U66037 ( .A(n51511), .B(n57904), .X(n29429) );
  nand_x1_sg U66038 ( .A(n50563), .B(n57870), .X(n30594) );
  nand_x1_sg U66039 ( .A(n56997), .B(n57886), .X(n30595) );
  nand_x1_sg U66040 ( .A(n50527), .B(n57876), .X(n29522) );
  nand_x1_sg U66041 ( .A(n56695), .B(n57901), .X(n29523) );
  nand_x1_sg U66042 ( .A(n50525), .B(n57877), .X(n29520) );
  nand_x1_sg U66043 ( .A(n56845), .B(n57901), .X(n29521) );
  nand_x1_sg U66044 ( .A(n53055), .B(n57878), .X(n29528) );
  nand_x1_sg U66045 ( .A(n51405), .B(n57901), .X(n29529) );
  nand_x1_sg U66046 ( .A(n53053), .B(n57880), .X(n29526) );
  nand_x1_sg U66047 ( .A(n47693), .B(n57901), .X(n29527) );
  nand_x1_sg U66048 ( .A(n50523), .B(n57880), .X(n29558) );
  nand_x1_sg U66049 ( .A(n56705), .B(n57907), .X(n29559) );
  nand_x1_sg U66050 ( .A(n53051), .B(n57878), .X(n29556) );
  nand_x1_sg U66051 ( .A(n51243), .B(n57910), .X(n29557) );
  nand_x1_sg U66052 ( .A(n50521), .B(n57871), .X(n29564) );
  nand_x1_sg U66053 ( .A(n56737), .B(n57908), .X(n29565) );
  nand_x1_sg U66054 ( .A(n53049), .B(n57878), .X(n29562) );
  nand_x1_sg U66055 ( .A(n51275), .B(n57909), .X(n29563) );
  nand_x1_sg U66056 ( .A(n50519), .B(n46213), .X(n29546) );
  nand_x1_sg U66057 ( .A(n56693), .B(n57904), .X(n29547) );
  nand_x1_sg U66058 ( .A(n53047), .B(n57875), .X(n29544) );
  nand_x1_sg U66059 ( .A(n51233), .B(n57895), .X(n29545) );
  nand_x1_sg U66060 ( .A(n50517), .B(n57877), .X(n29552) );
  nand_x1_sg U66061 ( .A(n56735), .B(n46207), .X(n29553) );
  nand_x1_sg U66062 ( .A(n53045), .B(n57878), .X(n29550) );
  nand_x1_sg U66063 ( .A(n51273), .B(n57900), .X(n29551) );
  nand_x1_sg U66064 ( .A(n50515), .B(n57880), .X(n29678) );
  nand_x1_sg U66065 ( .A(n56691), .B(n57907), .X(n29679) );
  nand_x1_sg U66066 ( .A(n53043), .B(n57875), .X(n29676) );
  nand_x1_sg U66067 ( .A(n51231), .B(n57896), .X(n29677) );
  nand_x1_sg U66068 ( .A(n53039), .B(n57875), .X(n29666) );
  nand_x1_sg U66069 ( .A(n51271), .B(n57910), .X(n29667) );
  nand_x1_sg U66070 ( .A(n53037), .B(n46213), .X(n29664) );
  nand_x1_sg U66071 ( .A(n51229), .B(n57911), .X(n29665) );
  nand_x1_sg U66072 ( .A(n53035), .B(n57876), .X(n29672) );
  nand_x1_sg U66073 ( .A(n47645), .B(n46207), .X(n29673) );
  nand_x1_sg U66074 ( .A(n53033), .B(n57877), .X(n29670) );
  nand_x1_sg U66075 ( .A(n47643), .B(n57900), .X(n29671) );
  nand_x1_sg U66076 ( .A(n50503), .B(n57875), .X(n29630) );
  nand_x1_sg U66077 ( .A(n56687), .B(n57899), .X(n29631) );
  nand_x1_sg U66078 ( .A(n53023), .B(n57875), .X(n29628) );
  nand_x1_sg U66079 ( .A(n51227), .B(n57899), .X(n29629) );
  nand_x1_sg U66080 ( .A(n50501), .B(n57878), .X(n29636) );
  nand_x1_sg U66081 ( .A(n56729), .B(n57886), .X(n29637) );
  nand_x1_sg U66082 ( .A(n53021), .B(n57878), .X(n29634) );
  nand_x1_sg U66083 ( .A(n51267), .B(n57911), .X(n29635) );
  nand_x1_sg U66084 ( .A(n50499), .B(n57877), .X(n29618) );
  nand_x1_sg U66085 ( .A(n56685), .B(n57899), .X(n29619) );
  nand_x1_sg U66086 ( .A(n53019), .B(n46213), .X(n29616) );
  nand_x1_sg U66087 ( .A(n51225), .B(n57899), .X(n29617) );
  nand_x1_sg U66088 ( .A(n53017), .B(n57880), .X(n29624) );
  nand_x1_sg U66089 ( .A(n47641), .B(n57899), .X(n29625) );
  nand_x1_sg U66090 ( .A(n50497), .B(n57880), .X(n29622) );
  nand_x1_sg U66091 ( .A(n56727), .B(n57899), .X(n29623) );
  nand_x1_sg U66092 ( .A(n53015), .B(n57880), .X(n29654) );
  nand_x1_sg U66093 ( .A(n51265), .B(n57908), .X(n29655) );
  nand_x1_sg U66094 ( .A(n53013), .B(n57877), .X(n29652) );
  nand_x1_sg U66095 ( .A(n51223), .B(n57909), .X(n29653) );
  nand_x1_sg U66096 ( .A(n53011), .B(n57877), .X(n29660) );
  nand_x1_sg U66097 ( .A(n47639), .B(n57907), .X(n29661) );
  nand_x1_sg U66098 ( .A(n53009), .B(n57876), .X(n29658) );
  nand_x1_sg U66099 ( .A(n47637), .B(n57898), .X(n29659) );
  nand_x1_sg U66100 ( .A(n50495), .B(n57877), .X(n29642) );
  nand_x1_sg U66101 ( .A(n56777), .B(n57901), .X(n29643) );
  nand_x1_sg U66102 ( .A(n53007), .B(n57877), .X(n29640) );
  nand_x1_sg U66103 ( .A(n51413), .B(n57903), .X(n29641) );
  nand_x1_sg U66104 ( .A(n53005), .B(n57880), .X(n29648) );
  nand_x1_sg U66105 ( .A(n47705), .B(n57887), .X(n29649) );
  nand_x1_sg U66106 ( .A(n50493), .B(n57876), .X(n29646) );
  nand_x1_sg U66107 ( .A(n56863), .B(n57911), .X(n29647) );
  nand_x1_sg U66108 ( .A(n50815), .B(n46212), .X(n29504) );
  nand_x1_sg U66109 ( .A(n56667), .B(n57911), .X(n29505) );
  nand_x1_sg U66110 ( .A(n53383), .B(n57878), .X(n29502) );
  nand_x1_sg U66111 ( .A(n51209), .B(n57898), .X(n29503) );
  nand_x1_sg U66112 ( .A(n53381), .B(n57876), .X(n29510) );
  nand_x1_sg U66113 ( .A(n47627), .B(n57911), .X(n29511) );
  nand_x1_sg U66114 ( .A(n50813), .B(n57877), .X(n29508) );
  nand_x1_sg U66115 ( .A(n56713), .B(n57904), .X(n29509) );
  nand_x1_sg U66116 ( .A(n53379), .B(n46213), .X(n29492) );
  nand_x1_sg U66117 ( .A(n51251), .B(n57898), .X(n29493) );
  nand_x1_sg U66118 ( .A(n53377), .B(n57872), .X(n29490) );
  nand_x1_sg U66119 ( .A(n51207), .B(n57899), .X(n29491) );
  nand_x1_sg U66120 ( .A(n53375), .B(n57875), .X(n29498) );
  nand_x1_sg U66121 ( .A(n47625), .B(n57900), .X(n29499) );
  nand_x1_sg U66122 ( .A(n53373), .B(n57877), .X(n29496) );
  nand_x1_sg U66123 ( .A(n47623), .B(n57895), .X(n29497) );
  nand_x1_sg U66124 ( .A(n50811), .B(n57876), .X(n29516) );
  nand_x1_sg U66125 ( .A(n56665), .B(n57911), .X(n29517) );
  nand_x1_sg U66126 ( .A(n53367), .B(n57878), .X(n29514) );
  nand_x1_sg U66127 ( .A(n51237), .B(n57911), .X(n29515) );
  nand_x1_sg U66128 ( .A(n50803), .B(n57880), .X(n29456) );
  nand_x1_sg U66129 ( .A(n56663), .B(n57889), .X(n29457) );
  nand_x1_sg U66130 ( .A(n53363), .B(n57878), .X(n29454) );
  nand_x1_sg U66131 ( .A(n51205), .B(n57903), .X(n29455) );
  nand_x1_sg U66132 ( .A(n50801), .B(n57877), .X(n29462) );
  nand_x1_sg U66133 ( .A(n56709), .B(n57909), .X(n29463) );
  nand_x1_sg U66134 ( .A(n53361), .B(n57880), .X(n29460) );
  nand_x1_sg U66135 ( .A(n51247), .B(n57893), .X(n29461) );
  nand_x1_sg U66136 ( .A(n50799), .B(n57875), .X(n29444) );
  nand_x1_sg U66137 ( .A(n56661), .B(n57903), .X(n29445) );
  nand_x1_sg U66138 ( .A(n53359), .B(n46213), .X(n29442) );
  nand_x1_sg U66139 ( .A(n51203), .B(n57903), .X(n29443) );
  nand_x1_sg U66140 ( .A(n53357), .B(n57880), .X(n29450) );
  nand_x1_sg U66141 ( .A(n47621), .B(n57903), .X(n29451) );
  nand_x1_sg U66142 ( .A(n50797), .B(n57878), .X(n29448) );
  nand_x1_sg U66143 ( .A(n56707), .B(n57903), .X(n29449) );
  nand_x1_sg U66144 ( .A(n53355), .B(n57873), .X(n29480) );
  nand_x1_sg U66145 ( .A(n51245), .B(n57902), .X(n29481) );
  nand_x1_sg U66146 ( .A(n53353), .B(n57878), .X(n29478) );
  nand_x1_sg U66147 ( .A(n51201), .B(n57902), .X(n29479) );
  nand_x1_sg U66148 ( .A(n53351), .B(n57880), .X(n29486) );
  nand_x1_sg U66149 ( .A(n47619), .B(n57902), .X(n29487) );
  nand_x1_sg U66150 ( .A(n53349), .B(n57876), .X(n29484) );
  nand_x1_sg U66151 ( .A(n47617), .B(n57902), .X(n29485) );
  nand_x1_sg U66152 ( .A(n50795), .B(n57875), .X(n29468) );
  nand_x1_sg U66153 ( .A(n56775), .B(n57890), .X(n29469) );
  nand_x1_sg U66154 ( .A(n53347), .B(n57878), .X(n29466) );
  nand_x1_sg U66155 ( .A(n51411), .B(n57891), .X(n29467) );
  nand_x1_sg U66156 ( .A(n53345), .B(n57880), .X(n29474) );
  nand_x1_sg U66157 ( .A(n47701), .B(n57902), .X(n29475) );
  nand_x1_sg U66158 ( .A(n50793), .B(n46212), .X(n29472) );
  nand_x1_sg U66159 ( .A(n56861), .B(n57902), .X(n29473) );
  nand_x1_sg U66160 ( .A(n50791), .B(n57877), .X(n29632) );
  nand_x1_sg U66161 ( .A(n56761), .B(n57898), .X(n29633) );
  nand_x1_sg U66162 ( .A(n53343), .B(n57875), .X(n29608) );
  nand_x1_sg U66163 ( .A(n51297), .B(n57900), .X(n29609) );
  nand_x1_sg U66164 ( .A(n50789), .B(n57876), .X(n29572) );
  nand_x1_sg U66165 ( .A(n56807), .B(n57886), .X(n29573) );
  nand_x1_sg U66166 ( .A(n50779), .B(n57880), .X(n29506) );
  nand_x1_sg U66167 ( .A(n56853), .B(n57911), .X(n29507) );
  nand_x1_sg U66168 ( .A(n53315), .B(n57878), .X(n29560) );
  nand_x1_sg U66169 ( .A(n51353), .B(n57898), .X(n29561) );
  nand_x1_sg U66170 ( .A(n50775), .B(n57880), .X(n29548) );
  nand_x1_sg U66171 ( .A(n56801), .B(n57898), .X(n29549) );
  nand_x1_sg U66172 ( .A(n50765), .B(n46213), .X(n29512) );
  nand_x1_sg U66173 ( .A(n56749), .B(n57911), .X(n29513) );
  nand_x1_sg U66174 ( .A(n53303), .B(n57878), .X(n29500) );
  nand_x1_sg U66175 ( .A(n47545), .B(n57896), .X(n29501) );
  nand_x1_sg U66176 ( .A(n53301), .B(n46212), .X(n29494) );
  nand_x1_sg U66177 ( .A(n47543), .B(n57887), .X(n29495) );
  nand_x1_sg U66178 ( .A(n53297), .B(n57875), .X(n29458) );
  nand_x1_sg U66179 ( .A(n47553), .B(n57894), .X(n29459) );
  nand_x1_sg U66180 ( .A(n50757), .B(n57876), .X(n29434) );
  nand_x1_sg U66181 ( .A(n56745), .B(n57904), .X(n29435) );
  nand_x1_sg U66182 ( .A(n53285), .B(n57877), .X(n29482) );
  nand_x1_sg U66183 ( .A(n51279), .B(n57902), .X(n29483) );
  nand_x1_sg U66184 ( .A(n50753), .B(n57872), .X(n29476) );
  nand_x1_sg U66185 ( .A(n56743), .B(n57902), .X(n29477) );
  nand_x1_sg U66186 ( .A(n53087), .B(n57871), .X(n29582) );
  nand_x1_sg U66187 ( .A(n51329), .B(n57911), .X(n29583) );
  nand_x1_sg U66188 ( .A(n50535), .B(n57877), .X(n29580) );
  nand_x1_sg U66189 ( .A(n56859), .B(n57909), .X(n29581) );
  nand_x1_sg U66190 ( .A(n53085), .B(n57872), .X(n29588) );
  nand_x1_sg U66191 ( .A(n47707), .B(n57895), .X(n29589) );
  nand_x1_sg U66192 ( .A(n53083), .B(n57875), .X(n29586) );
  nand_x1_sg U66193 ( .A(n51423), .B(n57900), .X(n29587) );
  nand_x1_sg U66194 ( .A(n53081), .B(n57877), .X(n29570) );
  nand_x1_sg U66195 ( .A(n51319), .B(n57907), .X(n29571) );
  nand_x1_sg U66196 ( .A(n53079), .B(n57880), .X(n29568) );
  nand_x1_sg U66197 ( .A(n47667), .B(n57900), .X(n29569) );
  nand_x1_sg U66198 ( .A(n50533), .B(n57876), .X(n29576) );
  nand_x1_sg U66199 ( .A(n56823), .B(n57907), .X(n29577) );
  nand_x1_sg U66200 ( .A(n53077), .B(n57878), .X(n29574) );
  nand_x1_sg U66201 ( .A(n51379), .B(n46207), .X(n29575) );
  nand_x1_sg U66202 ( .A(n53075), .B(n57877), .X(n29606) );
  nand_x1_sg U66203 ( .A(n51317), .B(n57900), .X(n29607) );
  nand_x1_sg U66204 ( .A(n53073), .B(n57876), .X(n29604) );
  nand_x1_sg U66205 ( .A(n47665), .B(n57900), .X(n29605) );
  nand_x1_sg U66206 ( .A(n53071), .B(n57875), .X(n29612) );
  nand_x1_sg U66207 ( .A(n51377), .B(n57900), .X(n29613) );
  nand_x1_sg U66208 ( .A(n53069), .B(n57880), .X(n29610) );
  nand_x1_sg U66209 ( .A(n47671), .B(n57900), .X(n29611) );
  nand_x1_sg U66210 ( .A(n53067), .B(n46209), .X(n29594) );
  nand_x1_sg U66211 ( .A(n51235), .B(n46207), .X(n29595) );
  nand_x1_sg U66212 ( .A(n53065), .B(n46210), .X(n29592) );
  nand_x1_sg U66213 ( .A(n47651), .B(n57887), .X(n29593) );
  nand_x1_sg U66214 ( .A(n53063), .B(n57878), .X(n29600) );
  nand_x1_sg U66215 ( .A(n47535), .B(n57900), .X(n29601) );
  nand_x1_sg U66216 ( .A(n50531), .B(n46212), .X(n29598) );
  nand_x1_sg U66217 ( .A(n56739), .B(n57911), .X(n29599) );
  nand_x1_sg U66218 ( .A(n53061), .B(n57875), .X(n29534) );
  nand_x1_sg U66219 ( .A(n51277), .B(n57901), .X(n29535) );
  nand_x1_sg U66220 ( .A(n53059), .B(n57875), .X(n29532) );
  nand_x1_sg U66221 ( .A(n47649), .B(n57901), .X(n29533) );
  nand_x1_sg U66222 ( .A(n50529), .B(n57875), .X(n29540) );
  nand_x1_sg U66223 ( .A(n56697), .B(n57888), .X(n29541) );
  nand_x1_sg U66224 ( .A(n53057), .B(n46213), .X(n29538) );
  nand_x1_sg U66225 ( .A(n47533), .B(n57902), .X(n29539) );
  nand_x1_sg U66226 ( .A(n53203), .B(n57878), .X(n29446) );
  nand_x1_sg U66227 ( .A(n51487), .B(n57903), .X(n29447) );
  nand_x1_sg U66228 ( .A(n53195), .B(n57877), .X(n29638) );
  nand_x1_sg U66229 ( .A(n51463), .B(n57886), .X(n29639) );
  nand_x1_sg U66230 ( .A(n50649), .B(n57877), .X(n29668) );
  nand_x1_sg U66231 ( .A(n56907), .B(n57907), .X(n29669) );
  nand_x1_sg U66232 ( .A(n53193), .B(n57880), .X(n29662) );
  nand_x1_sg U66233 ( .A(n51477), .B(n57911), .X(n29663) );
  nand_x1_sg U66234 ( .A(n50647), .B(n57875), .X(n29626) );
  nand_x1_sg U66235 ( .A(n56891), .B(n57899), .X(n29627) );
  nand_x1_sg U66236 ( .A(n53191), .B(n57875), .X(n29620) );
  nand_x1_sg U66237 ( .A(n51461), .B(n57899), .X(n29621) );
  nand_x1_sg U66238 ( .A(n53189), .B(n46213), .X(n29614) );
  nand_x1_sg U66239 ( .A(n47731), .B(n57900), .X(n29615) );
  nand_x1_sg U66240 ( .A(n50645), .B(n57877), .X(n29602) );
  nand_x1_sg U66241 ( .A(n56905), .B(n57900), .X(n29603) );
  nand_x1_sg U66242 ( .A(n53187), .B(n57878), .X(n29674) );
  nand_x1_sg U66243 ( .A(n51475), .B(n57895), .X(n29675) );
  nand_x1_sg U66244 ( .A(n53185), .B(n57878), .X(n29656) );
  nand_x1_sg U66245 ( .A(n51459), .B(n46207), .X(n29657) );
  nand_x1_sg U66246 ( .A(n53183), .B(n57877), .X(n29650) );
  nand_x1_sg U66247 ( .A(n47729), .B(n57900), .X(n29651) );
  nand_x1_sg U66248 ( .A(n53181), .B(n57875), .X(n29644) );
  nand_x1_sg U66249 ( .A(n47727), .B(n57886), .X(n29645) );
  nand_x1_sg U66250 ( .A(n53417), .B(n57877), .X(n29432) );
  nand_x1_sg U66251 ( .A(n51303), .B(n57904), .X(n29433) );
  nand_x1_sg U66252 ( .A(n53415), .B(n57876), .X(n29430) );
  nand_x1_sg U66253 ( .A(n47663), .B(n57904), .X(n29431) );
  nand_x1_sg U66254 ( .A(n53413), .B(n57880), .X(n29438) );
  nand_x1_sg U66255 ( .A(n51363), .B(n57904), .X(n29439) );
  nand_x1_sg U66256 ( .A(n53411), .B(n57880), .X(n29436) );
  nand_x1_sg U66257 ( .A(n47669), .B(n57904), .X(n29437) );
  nand_x1_sg U66258 ( .A(n53405), .B(n57877), .X(n29426) );
  nand_x1_sg U66259 ( .A(n47551), .B(n57904), .X(n29427) );
  nand_x1_sg U66260 ( .A(n50829), .B(n57877), .X(n29424) );
  nand_x1_sg U66261 ( .A(n56809), .B(n57904), .X(n29425) );
  nand_x1_sg U66262 ( .A(n50635), .B(n57875), .X(n29596) );
  nand_x1_sg U66263 ( .A(n55087), .B(n57910), .X(n29597) );
  nand_x1_sg U66264 ( .A(n53173), .B(n57880), .X(n29584) );
  nand_x1_sg U66265 ( .A(n47611), .B(n57908), .X(n29585) );
  nand_x1_sg U66266 ( .A(n53227), .B(n46212), .X(n29578) );
  nand_x1_sg U66267 ( .A(n51173), .B(n46207), .X(n29579) );
  nand_x1_sg U66268 ( .A(n53225), .B(n57876), .X(n29566) );
  nand_x1_sg U66269 ( .A(n51181), .B(n57911), .X(n29567) );
  nand_x1_sg U66270 ( .A(n53223), .B(n57875), .X(n29518) );
  nand_x1_sg U66271 ( .A(n47519), .B(n57911), .X(n29519) );
  nand_x1_sg U66272 ( .A(n53221), .B(n57880), .X(n29554) );
  nand_x1_sg U66273 ( .A(n51177), .B(n57907), .X(n29555) );
  nand_x1_sg U66274 ( .A(n50673), .B(n57871), .X(n29542) );
  nand_x1_sg U66275 ( .A(n55247), .B(n57886), .X(n29543) );
  nand_x1_sg U66276 ( .A(n53219), .B(n57876), .X(n29524) );
  nand_x1_sg U66277 ( .A(n51171), .B(n57901), .X(n29525) );
  nand_x1_sg U66278 ( .A(n50671), .B(n46213), .X(n29590) );
  nand_x1_sg U66279 ( .A(n55243), .B(n57900), .X(n29591) );
  nand_x1_sg U66280 ( .A(n50667), .B(n57873), .X(n29488) );
  nand_x1_sg U66281 ( .A(n55239), .B(n57886), .X(n29489) );
  nand_x1_sg U66282 ( .A(n53583), .B(n57873), .X(n30580) );
  nand_x1_sg U66283 ( .A(n47427), .B(n57887), .X(n30581) );
  nand_x1_sg U66284 ( .A(n50995), .B(n57877), .X(n30584) );
  nand_x1_sg U66285 ( .A(n56931), .B(n57887), .X(n30585) );
  nand_x1_sg U66286 ( .A(n50989), .B(n57870), .X(n30604) );
  nand_x1_sg U66287 ( .A(n56921), .B(n57886), .X(n30605) );
  nand_x1_sg U66288 ( .A(n53577), .B(n57870), .X(n30602) );
  nand_x1_sg U66289 ( .A(n47423), .B(n57886), .X(n30603) );
  nand_x1_sg U66290 ( .A(n50963), .B(n57872), .X(n30592) );
  nand_x1_sg U66291 ( .A(n55223), .B(n57886), .X(n30593) );
  nand_x1_sg U66292 ( .A(n50961), .B(n57870), .X(n30590) );
  nand_x1_sg U66293 ( .A(n55221), .B(n57887), .X(n30591) );
  nand_x1_sg U66294 ( .A(n53547), .B(n57870), .X(n30598) );
  nand_x1_sg U66295 ( .A(n51151), .B(n57886), .X(n30599) );
  nand_x1_sg U66296 ( .A(n53545), .B(n57870), .X(n30596) );
  nand_x1_sg U66297 ( .A(n47507), .B(n57886), .X(n30597) );
  nand_x1_sg U66298 ( .A(n50423), .B(n57871), .X(n30582) );
  nand_x1_sg U66299 ( .A(n55281), .B(n57887), .X(n30583) );
  nand_x1_sg U66300 ( .A(n52911), .B(n57876), .X(n30576) );
  nand_x1_sg U66301 ( .A(n51197), .B(n57887), .X(n30577) );
  nand_x1_sg U66302 ( .A(n53249), .B(n57870), .X(n30600) );
  nand_x1_sg U66303 ( .A(n51191), .B(n57886), .X(n30601) );
  nand_x1_sg U66304 ( .A(n50679), .B(n57880), .X(n30588) );
  nand_x1_sg U66305 ( .A(n55297), .B(n57887), .X(n30589) );
  nand_x1_sg U66306 ( .A(n50999), .B(n57877), .X(n30578) );
  nand_x1_sg U66307 ( .A(n55311), .B(n57887), .X(n30579) );
  nand_x1_sg U66308 ( .A(n50997), .B(n57876), .X(n30586) );
  nand_x1_sg U66309 ( .A(n55309), .B(n57887), .X(n30587) );
  nand_x1_sg U66310 ( .A(n50633), .B(n57870), .X(n29536) );
  nand_x1_sg U66311 ( .A(n55021), .B(n57887), .X(n29537) );
  nand_x1_sg U66312 ( .A(n50631), .B(n57873), .X(n29530) );
  nand_x1_sg U66313 ( .A(n55019), .B(n57901), .X(n29531) );
  nand_x1_sg U66314 ( .A(n52903), .B(n57717), .X(n38329) );
  nand_x1_sg U66315 ( .A(n49029), .B(n57765), .X(n38330) );
  nand_x1_sg U66316 ( .A(n52901), .B(n57717), .X(n38327) );
  nand_x1_sg U66317 ( .A(n49031), .B(n57766), .X(n38328) );
  nand_x1_sg U66318 ( .A(n52899), .B(n57717), .X(n38319) );
  nand_x1_sg U66319 ( .A(n49033), .B(n57734), .X(n38320) );
  nand_x1_sg U66320 ( .A(n52897), .B(n57717), .X(n38325) );
  nand_x1_sg U66321 ( .A(n49035), .B(n46198), .X(n38326) );
  nand_x1_sg U66322 ( .A(n52895), .B(n57682), .X(n37595) );
  nand_x1_sg U66323 ( .A(n49037), .B(n57759), .X(n37596) );
  nand_x1_sg U66324 ( .A(n52893), .B(n57681), .X(n37597) );
  nand_x1_sg U66325 ( .A(n49039), .B(n57773), .X(n37598) );
  nand_x1_sg U66326 ( .A(n57634), .B(n50387), .X(n37567) );
  nand_x1_sg U66327 ( .A(n52891), .B(n57766), .X(n37568) );
  nand_x1_sg U66328 ( .A(n52891), .B(n57717), .X(n38323) );
  nand_x1_sg U66329 ( .A(n49041), .B(n46197), .X(n38324) );
  nand_x1_sg U66330 ( .A(n57681), .B(n50385), .X(n37549) );
  nand_x1_sg U66331 ( .A(n52889), .B(n57766), .X(n37550) );
  nand_x1_sg U66332 ( .A(n52889), .B(n57717), .X(n38321) );
  nand_x1_sg U66333 ( .A(n49043), .B(n46201), .X(n38322) );
  nand_x1_sg U66334 ( .A(n57634), .B(n50383), .X(n37569) );
  nand_x1_sg U66335 ( .A(n52887), .B(n57744), .X(n37570) );
  nand_x1_sg U66336 ( .A(n52887), .B(n57676), .X(n38331) );
  nand_x1_sg U66337 ( .A(n49045), .B(n46201), .X(n38332) );
  nand_x1_sg U66338 ( .A(n57680), .B(n50381), .X(n37575) );
  nand_x1_sg U66339 ( .A(n52885), .B(n57756), .X(n37576) );
  nand_x1_sg U66340 ( .A(n52885), .B(n57682), .X(n37593) );
  nand_x1_sg U66341 ( .A(n49047), .B(n57747), .X(n37594) );
  nand_x1_sg U66342 ( .A(n57718), .B(n50379), .X(n37577) );
  nand_x1_sg U66343 ( .A(n52883), .B(n46200), .X(n37578) );
  nand_x1_sg U66344 ( .A(n52883), .B(n57681), .X(n37539) );
  nand_x1_sg U66345 ( .A(n49049), .B(n57754), .X(n37540) );
  nand_x1_sg U66346 ( .A(n57682), .B(n50377), .X(n37579) );
  nand_x1_sg U66347 ( .A(n52881), .B(n57742), .X(n37580) );
  nand_x1_sg U66348 ( .A(n52881), .B(n57682), .X(n37541) );
  nand_x1_sg U66349 ( .A(n49051), .B(n57770), .X(n37542) );
  nand_x1_sg U66350 ( .A(n57682), .B(n50375), .X(n37571) );
  nand_x1_sg U66351 ( .A(n52879), .B(n57758), .X(n37572) );
  nand_x1_sg U66352 ( .A(n52879), .B(n57709), .X(n37533) );
  nand_x1_sg U66353 ( .A(n49053), .B(n57760), .X(n37534) );
  nand_x1_sg U66354 ( .A(n57681), .B(n50373), .X(n37573) );
  nand_x1_sg U66355 ( .A(n52877), .B(n57761), .X(n37574) );
  nand_x1_sg U66356 ( .A(n52877), .B(n57708), .X(n37535) );
  nand_x1_sg U66357 ( .A(n49055), .B(n57749), .X(n37536) );
  nand_x1_sg U66358 ( .A(n57681), .B(n50371), .X(n37551) );
  nand_x1_sg U66359 ( .A(n52875), .B(n57758), .X(n37552) );
  nand_x1_sg U66360 ( .A(n52875), .B(n57682), .X(n37529) );
  nand_x1_sg U66361 ( .A(n49057), .B(n57748), .X(n37530) );
  nand_x1_sg U66362 ( .A(n57681), .B(n50369), .X(n37553) );
  nand_x1_sg U66363 ( .A(n52873), .B(n57764), .X(n37554) );
  nand_x1_sg U66364 ( .A(n52873), .B(n57682), .X(n37543) );
  nand_x1_sg U66365 ( .A(n49059), .B(n46201), .X(n37544) );
  nand_x1_sg U66366 ( .A(n57680), .B(n50367), .X(n37545) );
  nand_x1_sg U66367 ( .A(n52871), .B(n57772), .X(n37546) );
  nand_x1_sg U66368 ( .A(n52871), .B(n57717), .X(n37555) );
  nand_x1_sg U66369 ( .A(n49061), .B(n57771), .X(n37556) );
  nand_x1_sg U66370 ( .A(n57708), .B(n50365), .X(n37547) );
  nand_x1_sg U66371 ( .A(n52869), .B(n57749), .X(n37548) );
  nand_x1_sg U66372 ( .A(n52869), .B(n57682), .X(n37561) );
  nand_x1_sg U66373 ( .A(n49063), .B(n57748), .X(n37562) );
  nand_x1_sg U66374 ( .A(n57708), .B(n50363), .X(n37563) );
  nand_x1_sg U66375 ( .A(n52867), .B(n57748), .X(n37564) );
  nand_x1_sg U66376 ( .A(n52867), .B(n57634), .X(n37513) );
  nand_x1_sg U66377 ( .A(n49065), .B(n57775), .X(n37514) );
  nand_x1_sg U66378 ( .A(n57709), .B(n50361), .X(n37565) );
  nand_x1_sg U66379 ( .A(n52865), .B(n57765), .X(n37566) );
  nand_x1_sg U66380 ( .A(n52865), .B(n57720), .X(n37515) );
  nand_x1_sg U66381 ( .A(n49067), .B(n57742), .X(n37516) );
  nand_x1_sg U66382 ( .A(n57709), .B(n50359), .X(n37557) );
  nand_x1_sg U66383 ( .A(n52863), .B(n57743), .X(n37558) );
  nand_x1_sg U66384 ( .A(n52863), .B(n57634), .X(n37507) );
  nand_x1_sg U66385 ( .A(n49069), .B(n57746), .X(n37508) );
  nand_x1_sg U66386 ( .A(n57634), .B(n50357), .X(n37559) );
  nand_x1_sg U66387 ( .A(n52861), .B(n57760), .X(n37560) );
  nand_x1_sg U66388 ( .A(n52861), .B(n57634), .X(n37509) );
  nand_x1_sg U66389 ( .A(n49071), .B(n57726), .X(n37510) );
  nand_x1_sg U66390 ( .A(n52859), .B(n57680), .X(n37525) );
  nand_x1_sg U66391 ( .A(n49073), .B(n57754), .X(n37526) );
  nand_x1_sg U66392 ( .A(n52857), .B(n57709), .X(n37527) );
  nand_x1_sg U66393 ( .A(n49075), .B(n57762), .X(n37528) );
  nand_x1_sg U66394 ( .A(n52855), .B(n57680), .X(n37519) );
  nand_x1_sg U66395 ( .A(n49077), .B(n57755), .X(n37520) );
  nand_x1_sg U66396 ( .A(n52853), .B(n57720), .X(n37521) );
  nand_x1_sg U66397 ( .A(n49079), .B(n57759), .X(n37522) );
  nand_x1_sg U66398 ( .A(n57676), .B(n50307), .X(n38147) );
  nand_x1_sg U66399 ( .A(n52811), .B(n57739), .X(n38148) );
  nand_x1_sg U66400 ( .A(n57708), .B(n50305), .X(n37683) );
  nand_x1_sg U66401 ( .A(n52809), .B(n57765), .X(n37684) );
  nand_x1_sg U66402 ( .A(n57708), .B(n50303), .X(n37681) );
  nand_x1_sg U66403 ( .A(n52807), .B(n57763), .X(n37682) );
  nand_x1_sg U66404 ( .A(n52807), .B(n57717), .X(n38315) );
  nand_x1_sg U66405 ( .A(n48835), .B(n57758), .X(n38316) );
  nand_x1_sg U66406 ( .A(n57708), .B(n50301), .X(n37673) );
  nand_x1_sg U66407 ( .A(n52805), .B(n46200), .X(n37674) );
  nand_x1_sg U66408 ( .A(n52805), .B(n57717), .X(n38313) );
  nand_x1_sg U66409 ( .A(n48837), .B(n57748), .X(n38314) );
  nand_x1_sg U66410 ( .A(n57708), .B(n50299), .X(n37679) );
  nand_x1_sg U66411 ( .A(n52803), .B(n57755), .X(n37680) );
  nand_x1_sg U66412 ( .A(n57678), .B(n50103), .X(n37403) );
  nand_x1_sg U66413 ( .A(n52607), .B(n57759), .X(n37404) );
  nand_x1_sg U66414 ( .A(n57660), .B(n49981), .X(n37999) );
  nand_x1_sg U66415 ( .A(n52485), .B(n57770), .X(n38000) );
  nand_x1_sg U66416 ( .A(n57656), .B(n49979), .X(n38077) );
  nand_x1_sg U66417 ( .A(n52483), .B(n46197), .X(n38078) );
  nand_x1_sg U66418 ( .A(n57656), .B(n49977), .X(n38075) );
  nand_x1_sg U66419 ( .A(n52481), .B(n46200), .X(n38076) );
  nand_x1_sg U66420 ( .A(n57709), .B(n49975), .X(n37711) );
  nand_x1_sg U66421 ( .A(n52479), .B(n57755), .X(n37712) );
  nand_x1_sg U66422 ( .A(n57709), .B(n49973), .X(n37709) );
  nand_x1_sg U66423 ( .A(n52477), .B(n57756), .X(n37710) );
  nand_x1_sg U66424 ( .A(n57709), .B(n49971), .X(n37715) );
  nand_x1_sg U66425 ( .A(n52475), .B(n57757), .X(n37716) );
  nand_x1_sg U66426 ( .A(n57709), .B(n49969), .X(n37713) );
  nand_x1_sg U66427 ( .A(n52473), .B(n57747), .X(n37714) );
  nand_x1_sg U66428 ( .A(n57709), .B(n49967), .X(n37701) );
  nand_x1_sg U66429 ( .A(n52471), .B(n57764), .X(n37702) );
  nand_x1_sg U66430 ( .A(n57682), .B(n49965), .X(n37699) );
  nand_x1_sg U66431 ( .A(n52469), .B(n57749), .X(n37700) );
  nand_x1_sg U66432 ( .A(n57709), .B(n49963), .X(n37707) );
  nand_x1_sg U66433 ( .A(n52467), .B(n57755), .X(n37708) );
  nand_x1_sg U66434 ( .A(n57709), .B(n49961), .X(n37705) );
  nand_x1_sg U66435 ( .A(n52465), .B(n46198), .X(n37706) );
  nand_x1_sg U66436 ( .A(n57708), .B(n49959), .X(n37723) );
  nand_x1_sg U66437 ( .A(n52463), .B(n46201), .X(n37724) );
  nand_x1_sg U66438 ( .A(n57703), .B(n49957), .X(n37721) );
  nand_x1_sg U66439 ( .A(n52461), .B(n57766), .X(n37722) );
  nand_x1_sg U66440 ( .A(n57709), .B(n49955), .X(n37729) );
  nand_x1_sg U66441 ( .A(n52459), .B(n57758), .X(n37730) );
  nand_x1_sg U66442 ( .A(n57699), .B(n49953), .X(n37727) );
  nand_x1_sg U66443 ( .A(n52457), .B(n57775), .X(n37728) );
  nand_x1_sg U66444 ( .A(n57698), .B(n49951), .X(n37725) );
  nand_x1_sg U66445 ( .A(n52455), .B(n57775), .X(n37726) );
  nand_x1_sg U66446 ( .A(n57703), .B(n49949), .X(n37719) );
  nand_x1_sg U66447 ( .A(n52453), .B(n57775), .X(n37720) );
  nand_x1_sg U66448 ( .A(n57701), .B(n49947), .X(n37703) );
  nand_x1_sg U66449 ( .A(n52451), .B(n57747), .X(n37704) );
  nand_x1_sg U66450 ( .A(n52451), .B(n57661), .X(n37997) );
  nand_x1_sg U66451 ( .A(n48795), .B(n57773), .X(n37998) );
  nand_x1_sg U66452 ( .A(n57702), .B(n49945), .X(n37717) );
  nand_x1_sg U66453 ( .A(n52449), .B(n57771), .X(n37718) );
  nand_x1_sg U66454 ( .A(n52449), .B(n57656), .X(n38073) );
  nand_x1_sg U66455 ( .A(n48797), .B(n57750), .X(n38074) );
  nand_x1_sg U66456 ( .A(n57720), .B(n49943), .X(n37627) );
  nand_x1_sg U66457 ( .A(n52447), .B(n57764), .X(n37628) );
  nand_x1_sg U66458 ( .A(n52447), .B(n57660), .X(n38001) );
  nand_x1_sg U66459 ( .A(n48799), .B(n57771), .X(n38002) );
  nand_x1_sg U66460 ( .A(n57676), .B(n49941), .X(n38129) );
  nand_x1_sg U66461 ( .A(n52445), .B(n57729), .X(n38130) );
  nand_x1_sg U66462 ( .A(n52445), .B(n57682), .X(n37657) );
  nand_x1_sg U66463 ( .A(n48801), .B(n57764), .X(n37658) );
  nand_x1_sg U66464 ( .A(n57680), .B(n49939), .X(n37647) );
  nand_x1_sg U66465 ( .A(n52443), .B(n57745), .X(n37648) );
  nand_x1_sg U66466 ( .A(n52443), .B(n57720), .X(n37613) );
  nand_x1_sg U66467 ( .A(n48803), .B(n57749), .X(n37614) );
  nand_x1_sg U66468 ( .A(n57680), .B(n49937), .X(n37645) );
  nand_x1_sg U66469 ( .A(n52441), .B(n57746), .X(n37646) );
  nand_x1_sg U66470 ( .A(n52441), .B(n57667), .X(n37881) );
  nand_x1_sg U66471 ( .A(n48805), .B(n57756), .X(n37882) );
  nand_x1_sg U66472 ( .A(n57708), .B(n49935), .X(n37649) );
  nand_x1_sg U66473 ( .A(n52439), .B(n57760), .X(n37650) );
  nand_x1_sg U66474 ( .A(n52439), .B(n57682), .X(n37653) );
  nand_x1_sg U66475 ( .A(n48807), .B(n57762), .X(n37654) );
  nand_x1_sg U66476 ( .A(n57676), .B(n49933), .X(n38133) );
  nand_x1_sg U66477 ( .A(n52437), .B(n57745), .X(n38134) );
  nand_x1_sg U66478 ( .A(n52437), .B(n57708), .X(n37655) );
  nand_x1_sg U66479 ( .A(n48809), .B(n57742), .X(n37656) );
  nand_x1_sg U66480 ( .A(n57682), .B(n49931), .X(n37651) );
  nand_x1_sg U66481 ( .A(n52435), .B(n57747), .X(n37652) );
  nand_x1_sg U66482 ( .A(n52435), .B(n57673), .X(n38363) );
  nand_x1_sg U66483 ( .A(n48811), .B(n57759), .X(n38364) );
  nand_x1_sg U66484 ( .A(n57676), .B(n49929), .X(n38131) );
  nand_x1_sg U66485 ( .A(n52433), .B(n46197), .X(n38132) );
  nand_x1_sg U66486 ( .A(n52433), .B(n57707), .X(n38357) );
  nand_x1_sg U66487 ( .A(n48813), .B(n57757), .X(n38358) );
  nand_x1_sg U66488 ( .A(n57706), .B(n49927), .X(n38139) );
  nand_x1_sg U66489 ( .A(n52431), .B(n57755), .X(n38140) );
  nand_x1_sg U66490 ( .A(n52431), .B(n57680), .X(n37659) );
  nand_x1_sg U66491 ( .A(n48815), .B(n57743), .X(n37660) );
  nand_x1_sg U66492 ( .A(n57717), .B(n49925), .X(n38299) );
  nand_x1_sg U66493 ( .A(n52429), .B(n57761), .X(n38300) );
  nand_x1_sg U66494 ( .A(n52429), .B(n57681), .X(n37661) );
  nand_x1_sg U66495 ( .A(n48817), .B(n57744), .X(n37662) );
  nand_x1_sg U66496 ( .A(n57707), .B(n49923), .X(n38281) );
  nand_x1_sg U66497 ( .A(n52427), .B(n57730), .X(n38282) );
  nand_x1_sg U66498 ( .A(n52427), .B(n57667), .X(n37891) );
  nand_x1_sg U66499 ( .A(n48819), .B(n46198), .X(n37892) );
  nand_x1_sg U66500 ( .A(n57660), .B(n49921), .X(n38015) );
  nand_x1_sg U66501 ( .A(n52425), .B(n57758), .X(n38016) );
  nand_x1_sg U66502 ( .A(n52425), .B(n57672), .X(n38401) );
  nand_x1_sg U66503 ( .A(n48821), .B(n57754), .X(n38402) );
  nand_x1_sg U66504 ( .A(n57706), .B(n49919), .X(n38145) );
  nand_x1_sg U66505 ( .A(n52423), .B(n46198), .X(n38146) );
  nand_x1_sg U66506 ( .A(n52423), .B(n57680), .X(n38369) );
  nand_x1_sg U66507 ( .A(n48823), .B(n57758), .X(n38370) );
  nand_x1_sg U66508 ( .A(n57717), .B(n49917), .X(n38303) );
  nand_x1_sg U66509 ( .A(n52421), .B(n57756), .X(n38304) );
  nand_x1_sg U66510 ( .A(n52421), .B(n57682), .X(n37663) );
  nand_x1_sg U66511 ( .A(n48825), .B(n57763), .X(n37664) );
  nand_x1_sg U66512 ( .A(n57717), .B(n49915), .X(n38317) );
  nand_x1_sg U66513 ( .A(n52419), .B(n57765), .X(n38318) );
  nand_x1_sg U66514 ( .A(n52419), .B(n57634), .X(n38383) );
  nand_x1_sg U66515 ( .A(n48827), .B(n57764), .X(n38384) );
  nand_x1_sg U66516 ( .A(n57676), .B(n49913), .X(n38149) );
  nand_x1_sg U66517 ( .A(n52417), .B(n57765), .X(n38150) );
  nand_x1_sg U66518 ( .A(n52417), .B(n57680), .X(n37633) );
  nand_x1_sg U66519 ( .A(n48829), .B(n57743), .X(n37634) );
  nand_x1_sg U66520 ( .A(n52415), .B(n57680), .X(n37671) );
  nand_x1_sg U66521 ( .A(n48435), .B(n57743), .X(n37672) );
  nand_x1_sg U66522 ( .A(n52413), .B(n57681), .X(n37669) );
  nand_x1_sg U66523 ( .A(n48437), .B(n46198), .X(n37670) );
  nand_x1_sg U66524 ( .A(n52411), .B(n57708), .X(n37677) );
  nand_x1_sg U66525 ( .A(n48439), .B(n57744), .X(n37678) );
  nand_x1_sg U66526 ( .A(n57705), .B(n49905), .X(n38345) );
  nand_x1_sg U66527 ( .A(n52409), .B(n57766), .X(n38346) );
  nand_x1_sg U66528 ( .A(n52409), .B(n57680), .X(n37675) );
  nand_x1_sg U66529 ( .A(n48441), .B(n57727), .X(n37676) );
  nand_x1_sg U66530 ( .A(n57676), .B(n49903), .X(n38125) );
  nand_x1_sg U66531 ( .A(n52407), .B(n57765), .X(n38126) );
  nand_x1_sg U66532 ( .A(n52407), .B(n57681), .X(n37693) );
  nand_x1_sg U66533 ( .A(n48443), .B(n57750), .X(n37694) );
  nand_x1_sg U66534 ( .A(n57676), .B(n49901), .X(n38115) );
  nand_x1_sg U66535 ( .A(n52405), .B(n57732), .X(n38116) );
  nand_x1_sg U66536 ( .A(n52405), .B(n57709), .X(n37691) );
  nand_x1_sg U66537 ( .A(n48445), .B(n57760), .X(n37692) );
  nand_x1_sg U66538 ( .A(n57670), .B(n49899), .X(n37825) );
  nand_x1_sg U66539 ( .A(n52403), .B(n57759), .X(n37826) );
  nand_x1_sg U66540 ( .A(n52403), .B(n57699), .X(n37697) );
  nand_x1_sg U66541 ( .A(n48447), .B(n57748), .X(n37698) );
  nand_x1_sg U66542 ( .A(n57717), .B(n49897), .X(n38337) );
  nand_x1_sg U66543 ( .A(n52401), .B(n57766), .X(n38338) );
  nand_x1_sg U66544 ( .A(n52401), .B(n57700), .X(n37695) );
  nand_x1_sg U66545 ( .A(n48449), .B(n57761), .X(n37696) );
  nand_x1_sg U66546 ( .A(n57673), .B(n49895), .X(n38225) );
  nand_x1_sg U66547 ( .A(n52399), .B(n57747), .X(n38226) );
  nand_x1_sg U66548 ( .A(n52399), .B(n57634), .X(n37667) );
  nand_x1_sg U66549 ( .A(n48451), .B(n46200), .X(n37668) );
  nand_x1_sg U66550 ( .A(n57704), .B(n49893), .X(n38223) );
  nand_x1_sg U66551 ( .A(n52397), .B(n46197), .X(n38224) );
  nand_x1_sg U66552 ( .A(n52397), .B(n57697), .X(n37685) );
  nand_x1_sg U66553 ( .A(n48453), .B(n57742), .X(n37686) );
  nand_x1_sg U66554 ( .A(n57673), .B(n49891), .X(n38229) );
  nand_x1_sg U66555 ( .A(n52395), .B(n57762), .X(n38230) );
  nand_x1_sg U66556 ( .A(n52395), .B(n57698), .X(n37689) );
  nand_x1_sg U66557 ( .A(n48455), .B(n57762), .X(n37690) );
  nand_x1_sg U66558 ( .A(n57673), .B(n49889), .X(n38227) );
  nand_x1_sg U66559 ( .A(n52393), .B(n46197), .X(n38228) );
  nand_x1_sg U66560 ( .A(n52393), .B(n57716), .X(n37687) );
  nand_x1_sg U66561 ( .A(n48457), .B(n57772), .X(n37688) );
  nand_x1_sg U66562 ( .A(n57672), .B(n49887), .X(n38217) );
  nand_x1_sg U66563 ( .A(n52391), .B(n57756), .X(n38218) );
  nand_x1_sg U66564 ( .A(n52391), .B(n57716), .X(n38393) );
  nand_x1_sg U66565 ( .A(n48459), .B(n57755), .X(n38394) );
  nand_x1_sg U66566 ( .A(n57704), .B(n49885), .X(n38215) );
  nand_x1_sg U66567 ( .A(n52389), .B(n57765), .X(n38216) );
  nand_x1_sg U66568 ( .A(n52389), .B(n57676), .X(n38107) );
  nand_x1_sg U66569 ( .A(n48461), .B(n57733), .X(n38108) );
  nand_x1_sg U66570 ( .A(n57672), .B(n49883), .X(n38221) );
  nand_x1_sg U66571 ( .A(n52387), .B(n57772), .X(n38222) );
  nand_x1_sg U66572 ( .A(n52387), .B(n57707), .X(n37777) );
  nand_x1_sg U66573 ( .A(n48463), .B(n57747), .X(n37778) );
  nand_x1_sg U66574 ( .A(n57704), .B(n49881), .X(n38219) );
  nand_x1_sg U66575 ( .A(n52385), .B(n57749), .X(n38220) );
  nand_x1_sg U66576 ( .A(n52385), .B(n57708), .X(n37665) );
  nand_x1_sg U66577 ( .A(n48465), .B(n57761), .X(n37666) );
  nand_x1_sg U66578 ( .A(n57673), .B(n49879), .X(n38241) );
  nand_x1_sg U66579 ( .A(n52383), .B(n57747), .X(n38242) );
  nand_x1_sg U66580 ( .A(n52383), .B(n57706), .X(n38143) );
  nand_x1_sg U66581 ( .A(n48467), .B(n57743), .X(n38144) );
  nand_x1_sg U66582 ( .A(n57673), .B(n49877), .X(n38239) );
  nand_x1_sg U66583 ( .A(n52381), .B(n57747), .X(n38240) );
  nand_x1_sg U66584 ( .A(n52381), .B(n57717), .X(n38141) );
  nand_x1_sg U66585 ( .A(n48469), .B(n57746), .X(n38142) );
  nand_x1_sg U66586 ( .A(n57672), .B(n49875), .X(n38245) );
  nand_x1_sg U66587 ( .A(n52379), .B(n57747), .X(n38246) );
  nand_x1_sg U66588 ( .A(n52379), .B(n57681), .X(n37601) );
  nand_x1_sg U66589 ( .A(n48471), .B(n57749), .X(n37602) );
  nand_x1_sg U66590 ( .A(n57672), .B(n49873), .X(n38243) );
  nand_x1_sg U66591 ( .A(n52377), .B(n57766), .X(n38244) );
  nand_x1_sg U66592 ( .A(n52377), .B(n57676), .X(n38105) );
  nand_x1_sg U66593 ( .A(n48473), .B(n57762), .X(n38106) );
  nand_x1_sg U66594 ( .A(n57673), .B(n49871), .X(n38233) );
  nand_x1_sg U66595 ( .A(n52375), .B(n57742), .X(n38234) );
  nand_x1_sg U66596 ( .A(n52375), .B(n57676), .X(n38127) );
  nand_x1_sg U66597 ( .A(n48475), .B(n57773), .X(n38128) );
  nand_x1_sg U66598 ( .A(n57673), .B(n49869), .X(n38231) );
  nand_x1_sg U66599 ( .A(n52373), .B(n57744), .X(n38232) );
  nand_x1_sg U66600 ( .A(n52373), .B(n57676), .X(n38123) );
  nand_x1_sg U66601 ( .A(n48477), .B(n57764), .X(n38124) );
  nand_x1_sg U66602 ( .A(n57673), .B(n49867), .X(n38237) );
  nand_x1_sg U66603 ( .A(n52371), .B(n57743), .X(n38238) );
  nand_x1_sg U66604 ( .A(n52371), .B(n57708), .X(n38343) );
  nand_x1_sg U66605 ( .A(n48479), .B(n46201), .X(n38344) );
  nand_x1_sg U66606 ( .A(n57678), .B(n49865), .X(n38269) );
  nand_x1_sg U66607 ( .A(n52369), .B(n57756), .X(n38270) );
  nand_x1_sg U66608 ( .A(n52369), .B(n57673), .X(n38235) );
  nand_x1_sg U66609 ( .A(n48481), .B(n57744), .X(n38236) );
  nand_x1_sg U66610 ( .A(n57678), .B(n49863), .X(n38259) );
  nand_x1_sg U66611 ( .A(n52367), .B(n57754), .X(n38260) );
  nand_x1_sg U66612 ( .A(n52367), .B(n57672), .X(n38193) );
  nand_x1_sg U66613 ( .A(n48483), .B(n57766), .X(n38194) );
  nand_x1_sg U66614 ( .A(n57672), .B(n49861), .X(n38257) );
  nand_x1_sg U66615 ( .A(n52365), .B(n57755), .X(n38258) );
  nand_x1_sg U66616 ( .A(n52365), .B(n57672), .X(n38191) );
  nand_x1_sg U66617 ( .A(n48485), .B(n57766), .X(n38192) );
  nand_x1_sg U66618 ( .A(n57678), .B(n49859), .X(n38263) );
  nand_x1_sg U66619 ( .A(n52363), .B(n57757), .X(n38264) );
  nand_x1_sg U66620 ( .A(n52363), .B(n57672), .X(n38197) );
  nand_x1_sg U66621 ( .A(n48487), .B(n57766), .X(n38198) );
  nand_x1_sg U66622 ( .A(n57678), .B(n49857), .X(n38261) );
  nand_x1_sg U66623 ( .A(n52361), .B(n57754), .X(n38262) );
  nand_x1_sg U66624 ( .A(n52361), .B(n57672), .X(n38195) );
  nand_x1_sg U66625 ( .A(n48489), .B(n57766), .X(n38196) );
  nand_x1_sg U66626 ( .A(n57707), .B(n49855), .X(n38279) );
  nand_x1_sg U66627 ( .A(n52359), .B(n57760), .X(n38280) );
  nand_x1_sg U66628 ( .A(n52359), .B(n57674), .X(n38185) );
  nand_x1_sg U66629 ( .A(n48491), .B(n57742), .X(n38186) );
  nand_x1_sg U66630 ( .A(n57678), .B(n49853), .X(n38277) );
  nand_x1_sg U66631 ( .A(n52357), .B(n57756), .X(n38278) );
  nand_x1_sg U66632 ( .A(n52357), .B(n57674), .X(n38183) );
  nand_x1_sg U66633 ( .A(n48493), .B(n57748), .X(n38184) );
  nand_x1_sg U66634 ( .A(n52355), .B(n57672), .X(n38189) );
  nand_x1_sg U66635 ( .A(n48495), .B(n57770), .X(n38190) );
  nand_x1_sg U66636 ( .A(n52353), .B(n57674), .X(n38187) );
  nand_x1_sg U66637 ( .A(n48497), .B(n46201), .X(n38188) );
  nand_x1_sg U66638 ( .A(n52351), .B(n57695), .X(n38209) );
  nand_x1_sg U66639 ( .A(n48499), .B(n57775), .X(n38210) );
  nand_x1_sg U66640 ( .A(n52349), .B(n57677), .X(n38207) );
  nand_x1_sg U66641 ( .A(n48501), .B(n46201), .X(n38208) );
  nand_x1_sg U66642 ( .A(n52347), .B(n57679), .X(n38213) );
  nand_x1_sg U66643 ( .A(n48503), .B(n57759), .X(n38214) );
  nand_x1_sg U66644 ( .A(n52345), .B(n57674), .X(n38211) );
  nand_x1_sg U66645 ( .A(n48505), .B(n57746), .X(n38212) );
  nand_x1_sg U66646 ( .A(n52343), .B(n57672), .X(n38201) );
  nand_x1_sg U66647 ( .A(n48507), .B(n57761), .X(n38202) );
  nand_x1_sg U66648 ( .A(n52341), .B(n57672), .X(n38199) );
  nand_x1_sg U66649 ( .A(n48509), .B(n57755), .X(n38200) );
  nand_x1_sg U66650 ( .A(n57672), .B(n49835), .X(n38251) );
  nand_x1_sg U66651 ( .A(n52339), .B(n57750), .X(n38252) );
  nand_x1_sg U66652 ( .A(n52339), .B(n57672), .X(n38205) );
  nand_x1_sg U66653 ( .A(n48511), .B(n57762), .X(n38206) );
  nand_x1_sg U66654 ( .A(n52337), .B(n57672), .X(n38203) );
  nand_x1_sg U66655 ( .A(n48513), .B(n57750), .X(n38204) );
  nand_x1_sg U66656 ( .A(n52335), .B(n57678), .X(n38267) );
  nand_x1_sg U66657 ( .A(n48515), .B(n57757), .X(n38268) );
  nand_x1_sg U66658 ( .A(n52333), .B(n57707), .X(n38265) );
  nand_x1_sg U66659 ( .A(n48517), .B(n57749), .X(n38266) );
  nand_x1_sg U66660 ( .A(n52331), .B(n57678), .X(n38271) );
  nand_x1_sg U66661 ( .A(n48519), .B(n57758), .X(n38272) );
  nand_x1_sg U66662 ( .A(n52327), .B(n57672), .X(n38255) );
  nand_x1_sg U66663 ( .A(n48523), .B(n57754), .X(n38256) );
  nand_x1_sg U66664 ( .A(n52325), .B(n57672), .X(n38253) );
  nand_x1_sg U66665 ( .A(n48525), .B(n57755), .X(n38254) );
  nand_x1_sg U66666 ( .A(n57676), .B(n49811), .X(n38121) );
  nand_x1_sg U66667 ( .A(n52315), .B(n57737), .X(n38122) );
  nand_x1_sg U66668 ( .A(n57676), .B(n49809), .X(n38119) );
  nand_x1_sg U66669 ( .A(n52313), .B(n57738), .X(n38120) );
  nand_x1_sg U66670 ( .A(n52311), .B(n57676), .X(n38137) );
  nand_x1_sg U66671 ( .A(n48539), .B(n57728), .X(n38138) );
  nand_x1_sg U66672 ( .A(n57676), .B(n49805), .X(n38111) );
  nand_x1_sg U66673 ( .A(n52309), .B(n57728), .X(n38112) );
  nand_x1_sg U66674 ( .A(n52309), .B(n57706), .X(n38135) );
  nand_x1_sg U66675 ( .A(n48541), .B(n57747), .X(n38136) );
  nand_x1_sg U66676 ( .A(n57676), .B(n49803), .X(n38113) );
  nand_x1_sg U66677 ( .A(n52307), .B(n57755), .X(n38114) );
  nand_x1_sg U66678 ( .A(n57675), .B(n49785), .X(n38155) );
  nand_x1_sg U66679 ( .A(n52289), .B(n57766), .X(n38156) );
  nand_x1_sg U66680 ( .A(n57675), .B(n49783), .X(n38153) );
  nand_x1_sg U66681 ( .A(n52287), .B(n57757), .X(n38154) );
  nand_x1_sg U66682 ( .A(n57676), .B(n49781), .X(n38151) );
  nand_x1_sg U66683 ( .A(n52285), .B(n46200), .X(n38152) );
  nand_x1_sg U66684 ( .A(n57675), .B(n49775), .X(n38169) );
  nand_x1_sg U66685 ( .A(n52279), .B(n57758), .X(n38170) );
  nand_x1_sg U66686 ( .A(n57675), .B(n49773), .X(n38167) );
  nand_x1_sg U66687 ( .A(n52277), .B(n57759), .X(n38168) );
  nand_x1_sg U66688 ( .A(n57674), .B(n49771), .X(n38173) );
  nand_x1_sg U66689 ( .A(n52275), .B(n57756), .X(n38174) );
  nand_x1_sg U66690 ( .A(n57674), .B(n49769), .X(n38171) );
  nand_x1_sg U66691 ( .A(n52273), .B(n57770), .X(n38172) );
  nand_x1_sg U66692 ( .A(n57675), .B(n49767), .X(n38161) );
  nand_x1_sg U66693 ( .A(n52271), .B(n57758), .X(n38162) );
  nand_x1_sg U66694 ( .A(n57675), .B(n49765), .X(n38159) );
  nand_x1_sg U66695 ( .A(n52269), .B(n57765), .X(n38160) );
  nand_x1_sg U66696 ( .A(n57675), .B(n49763), .X(n38165) );
  nand_x1_sg U66697 ( .A(n52267), .B(n57765), .X(n38166) );
  nand_x1_sg U66698 ( .A(n57675), .B(n49761), .X(n38163) );
  nand_x1_sg U66699 ( .A(n52265), .B(n57760), .X(n38164) );
  nand_x1_sg U66700 ( .A(n57717), .B(n49759), .X(n38297) );
  nand_x1_sg U66701 ( .A(n52263), .B(n57757), .X(n38298) );
  nand_x1_sg U66702 ( .A(n52263), .B(n57674), .X(n38179) );
  nand_x1_sg U66703 ( .A(n48587), .B(n57775), .X(n38180) );
  nand_x1_sg U66704 ( .A(n57717), .B(n49757), .X(n38295) );
  nand_x1_sg U66705 ( .A(n52261), .B(n57737), .X(n38296) );
  nand_x1_sg U66706 ( .A(n52261), .B(n57674), .X(n38177) );
  nand_x1_sg U66707 ( .A(n48589), .B(n46198), .X(n38178) );
  nand_x1_sg U66708 ( .A(n52259), .B(n57674), .X(n38181) );
  nand_x1_sg U66709 ( .A(n48591), .B(n57775), .X(n38182) );
  nand_x1_sg U66710 ( .A(n57682), .B(n49747), .X(n37589) );
  nand_x1_sg U66711 ( .A(n52251), .B(n57744), .X(n37590) );
  nand_x1_sg U66712 ( .A(n52251), .B(n57675), .X(n38157) );
  nand_x1_sg U66713 ( .A(n48599), .B(n57745), .X(n38158) );
  nand_x1_sg U66714 ( .A(n52249), .B(n57682), .X(n37591) );
  nand_x1_sg U66715 ( .A(n48601), .B(n57759), .X(n37592) );
  nand_x1_sg U66716 ( .A(n57707), .B(n49743), .X(n38293) );
  nand_x1_sg U66717 ( .A(n52247), .B(n57754), .X(n38294) );
  nand_x1_sg U66718 ( .A(n52247), .B(n57682), .X(n37583) );
  nand_x1_sg U66719 ( .A(n48603), .B(n57761), .X(n37584) );
  nand_x1_sg U66720 ( .A(n52245), .B(n57682), .X(n37585) );
  nand_x1_sg U66721 ( .A(n48605), .B(n57747), .X(n37586) );
  nand_x1_sg U66722 ( .A(n52217), .B(n57679), .X(n37385) );
  nand_x1_sg U66723 ( .A(n48237), .B(n57770), .X(n37386) );
  nand_x1_sg U66724 ( .A(n52215), .B(n57678), .X(n37405) );
  nand_x1_sg U66725 ( .A(n48239), .B(n57729), .X(n37406) );
  nand_x1_sg U66726 ( .A(n52213), .B(n57673), .X(n37411) );
  nand_x1_sg U66727 ( .A(n48241), .B(n57729), .X(n37412) );
  nand_x1_sg U66728 ( .A(n57673), .B(n49707), .X(n37421) );
  nand_x1_sg U66729 ( .A(n52211), .B(n57754), .X(n37422) );
  nand_x1_sg U66730 ( .A(n52211), .B(n57673), .X(n37413) );
  nand_x1_sg U66731 ( .A(n48243), .B(n57762), .X(n37414) );
  nand_x1_sg U66732 ( .A(n57673), .B(n49705), .X(n37423) );
  nand_x1_sg U66733 ( .A(n52209), .B(n57762), .X(n37424) );
  nand_x1_sg U66734 ( .A(n52209), .B(n57673), .X(n37415) );
  nand_x1_sg U66735 ( .A(n48245), .B(n57747), .X(n37416) );
  nand_x1_sg U66736 ( .A(n57678), .B(n49703), .X(n37391) );
  nand_x1_sg U66737 ( .A(n52207), .B(n57762), .X(n37392) );
  nand_x1_sg U66738 ( .A(n52207), .B(n57673), .X(n37407) );
  nand_x1_sg U66739 ( .A(n48247), .B(n57772), .X(n37408) );
  nand_x1_sg U66740 ( .A(n57678), .B(n49701), .X(n37397) );
  nand_x1_sg U66741 ( .A(n52205), .B(n57765), .X(n37398) );
  nand_x1_sg U66742 ( .A(n52205), .B(n57673), .X(n37409) );
  nand_x1_sg U66743 ( .A(n48249), .B(n57771), .X(n37410) );
  nand_x1_sg U66744 ( .A(n57677), .B(n49699), .X(n37425) );
  nand_x1_sg U66745 ( .A(n52203), .B(n57749), .X(n37426) );
  nand_x1_sg U66746 ( .A(n52203), .B(n57679), .X(n37387) );
  nand_x1_sg U66747 ( .A(n48251), .B(n57756), .X(n37388) );
  nand_x1_sg U66748 ( .A(n57673), .B(n49697), .X(n37419) );
  nand_x1_sg U66749 ( .A(n52201), .B(n57762), .X(n37420) );
  nand_x1_sg U66750 ( .A(n52201), .B(n57678), .X(n37389) );
  nand_x1_sg U66751 ( .A(n48253), .B(n57750), .X(n37390) );
  nand_x1_sg U66752 ( .A(n57677), .B(n49695), .X(n37427) );
  nand_x1_sg U66753 ( .A(n52199), .B(n57755), .X(n37428) );
  nand_x1_sg U66754 ( .A(n57677), .B(n49693), .X(n37429) );
  nand_x1_sg U66755 ( .A(n52197), .B(n57770), .X(n37430) );
  nand_x1_sg U66756 ( .A(n52197), .B(n57679), .X(n37383) );
  nand_x1_sg U66757 ( .A(n48257), .B(n46200), .X(n37384) );
  nand_x1_sg U66758 ( .A(n52195), .B(n57678), .X(n37399) );
  nand_x1_sg U66759 ( .A(n48259), .B(n57759), .X(n37400) );
  nand_x1_sg U66760 ( .A(n52193), .B(n57678), .X(n37401) );
  nand_x1_sg U66761 ( .A(n48261), .B(n57762), .X(n37402) );
  nand_x1_sg U66762 ( .A(n52191), .B(n57678), .X(n37393) );
  nand_x1_sg U66763 ( .A(n48263), .B(n57770), .X(n37394) );
  nand_x1_sg U66764 ( .A(n52189), .B(n57678), .X(n37395) );
  nand_x1_sg U66765 ( .A(n48265), .B(n57761), .X(n37396) );
  nand_x1_sg U66766 ( .A(n52187), .B(n57677), .X(n37439) );
  nand_x1_sg U66767 ( .A(n48267), .B(n57743), .X(n37440) );
  nand_x1_sg U66768 ( .A(n52185), .B(n57677), .X(n37441) );
  nand_x1_sg U66769 ( .A(n48269), .B(n57744), .X(n37442) );
  nand_x1_sg U66770 ( .A(n52183), .B(n57677), .X(n37433) );
  nand_x1_sg U66771 ( .A(n48271), .B(n57748), .X(n37434) );
  nand_x1_sg U66772 ( .A(n52181), .B(n57677), .X(n37435) );
  nand_x1_sg U66773 ( .A(n48273), .B(n57744), .X(n37436) );
  nand_x1_sg U66774 ( .A(n52179), .B(n57673), .X(n37417) );
  nand_x1_sg U66775 ( .A(n48275), .B(n57762), .X(n37418) );
  nand_x1_sg U66776 ( .A(n52177), .B(n57677), .X(n37431) );
  nand_x1_sg U66777 ( .A(n48277), .B(n57750), .X(n37432) );
  nand_x1_sg U66778 ( .A(n52175), .B(n57677), .X(n37437) );
  nand_x1_sg U66779 ( .A(n48279), .B(n57762), .X(n37438) );
  nand_x1_sg U66780 ( .A(n57707), .B(n49667), .X(n37463) );
  nand_x1_sg U66781 ( .A(n52171), .B(n57750), .X(n37464) );
  nand_x1_sg U66782 ( .A(n57704), .B(n49665), .X(n37465) );
  nand_x1_sg U66783 ( .A(n52169), .B(n57773), .X(n37466) );
  nand_x1_sg U66784 ( .A(n57705), .B(n49663), .X(n37457) );
  nand_x1_sg U66785 ( .A(n52167), .B(n57724), .X(n37458) );
  nand_x1_sg U66786 ( .A(n57718), .B(n49661), .X(n37459) );
  nand_x1_sg U66787 ( .A(n52165), .B(n57725), .X(n37460) );
  nand_x1_sg U66788 ( .A(n57682), .B(n49659), .X(n37475) );
  nand_x1_sg U66789 ( .A(n52163), .B(n57771), .X(n37476) );
  nand_x1_sg U66790 ( .A(n57680), .B(n49657), .X(n37477) );
  nand_x1_sg U66791 ( .A(n52161), .B(n57736), .X(n37478) );
  nand_x1_sg U66792 ( .A(n57681), .B(n49655), .X(n37469) );
  nand_x1_sg U66793 ( .A(n52159), .B(n57734), .X(n37470) );
  nand_x1_sg U66794 ( .A(n57681), .B(n49653), .X(n37471) );
  nand_x1_sg U66795 ( .A(n52157), .B(n57739), .X(n37472) );
  nand_x1_sg U66796 ( .A(n57697), .B(n49651), .X(n37445) );
  nand_x1_sg U66797 ( .A(n52155), .B(n57765), .X(n37446) );
  nand_x1_sg U66798 ( .A(n57720), .B(n49649), .X(n37447) );
  nand_x1_sg U66799 ( .A(n52153), .B(n57750), .X(n37448) );
  nand_x1_sg U66800 ( .A(n57718), .B(n49643), .X(n37455) );
  nand_x1_sg U66801 ( .A(n52147), .B(n57766), .X(n37456) );
  nand_x1_sg U66802 ( .A(n57706), .B(n49639), .X(n37443) );
  nand_x1_sg U66803 ( .A(n52143), .B(n57759), .X(n37444) );
  nand_x1_sg U66804 ( .A(n57695), .B(n49635), .X(n37501) );
  nand_x1_sg U66805 ( .A(n52139), .B(n57765), .X(n37502) );
  nand_x1_sg U66806 ( .A(n57696), .B(n49633), .X(n37503) );
  nand_x1_sg U66807 ( .A(n52137), .B(n57765), .X(n37504) );
  nand_x1_sg U66808 ( .A(n57693), .B(n49631), .X(n37497) );
  nand_x1_sg U66809 ( .A(n52135), .B(n57746), .X(n37498) );
  nand_x1_sg U66810 ( .A(n52133), .B(n57694), .X(n37499) );
  nand_x1_sg U66811 ( .A(n48321), .B(n57728), .X(n37500) );
  nand_x1_sg U66812 ( .A(n52131), .B(n57708), .X(n37487) );
  nand_x1_sg U66813 ( .A(n48323), .B(n57773), .X(n37488) );
  nand_x1_sg U66814 ( .A(n52129), .B(n57709), .X(n37481) );
  nand_x1_sg U66815 ( .A(n48325), .B(n57747), .X(n37482) );
  nand_x1_sg U66816 ( .A(n52127), .B(n57715), .X(n37493) );
  nand_x1_sg U66817 ( .A(n48327), .B(n57748), .X(n37494) );
  nand_x1_sg U66818 ( .A(n52125), .B(n57703), .X(n37495) );
  nand_x1_sg U66819 ( .A(n48329), .B(n57759), .X(n37496) );
  nand_x1_sg U66820 ( .A(n52123), .B(n57634), .X(n37473) );
  nand_x1_sg U66821 ( .A(n48331), .B(n57730), .X(n37474) );
  nand_x1_sg U66822 ( .A(n52121), .B(n57697), .X(n37461) );
  nand_x1_sg U66823 ( .A(n48333), .B(n57728), .X(n37462) );
  nand_x1_sg U66824 ( .A(n52119), .B(n57716), .X(n37479) );
  nand_x1_sg U66825 ( .A(n48335), .B(n57758), .X(n37480) );
  nand_x1_sg U66826 ( .A(n52117), .B(n57698), .X(n37467) );
  nand_x1_sg U66827 ( .A(n48337), .B(n57738), .X(n37468) );
  nand_x1_sg U66828 ( .A(n52115), .B(n57703), .X(n37489) );
  nand_x1_sg U66829 ( .A(n48339), .B(n57759), .X(n37490) );
  nand_x1_sg U66830 ( .A(n52113), .B(n57701), .X(n37491) );
  nand_x1_sg U66831 ( .A(n48341), .B(n57759), .X(n37492) );
  nand_x1_sg U66832 ( .A(n52111), .B(n57715), .X(n37483) );
  nand_x1_sg U66833 ( .A(n48343), .B(n57757), .X(n37484) );
  nand_x1_sg U66834 ( .A(n52109), .B(n57681), .X(n37485) );
  nand_x1_sg U66835 ( .A(n48345), .B(n57761), .X(n37486) );
  nand_x1_sg U66836 ( .A(n57681), .B(n49515), .X(n37607) );
  nand_x1_sg U66837 ( .A(n52019), .B(n57763), .X(n37608) );
  nand_x1_sg U66838 ( .A(n57708), .B(n49471), .X(n38373) );
  nand_x1_sg U66839 ( .A(n51975), .B(n57759), .X(n38374) );
  nand_x1_sg U66840 ( .A(n57681), .B(n49469), .X(n38371) );
  nand_x1_sg U66841 ( .A(n51973), .B(n57773), .X(n38372) );
  nand_x1_sg U66842 ( .A(n57682), .B(n49467), .X(n38375) );
  nand_x1_sg U66843 ( .A(n51971), .B(n57761), .X(n38376) );
  nand_x1_sg U66844 ( .A(n57678), .B(n49463), .X(n38361) );
  nand_x1_sg U66845 ( .A(n51967), .B(n57771), .X(n38362) );
  nand_x1_sg U66846 ( .A(n57704), .B(n49461), .X(n38359) );
  nand_x1_sg U66847 ( .A(n51965), .B(n57766), .X(n38360) );
  nand_x1_sg U66848 ( .A(n57705), .B(n49459), .X(n38367) );
  nand_x1_sg U66849 ( .A(n51963), .B(n57754), .X(n38368) );
  nand_x1_sg U66850 ( .A(n57701), .B(n49457), .X(n38365) );
  nand_x1_sg U66851 ( .A(n51961), .B(n46198), .X(n38366) );
  nand_x1_sg U66852 ( .A(n57708), .B(n49455), .X(n38387) );
  nand_x1_sg U66853 ( .A(n51959), .B(n57754), .X(n38388) );
  nand_x1_sg U66854 ( .A(n57681), .B(n49453), .X(n38385) );
  nand_x1_sg U66855 ( .A(n51957), .B(n57770), .X(n38386) );
  nand_x1_sg U66856 ( .A(n57682), .B(n49451), .X(n38391) );
  nand_x1_sg U66857 ( .A(n51955), .B(n57772), .X(n38392) );
  nand_x1_sg U66858 ( .A(n57709), .B(n49449), .X(n38389) );
  nand_x1_sg U66859 ( .A(n51953), .B(n57762), .X(n38390) );
  nand_x1_sg U66860 ( .A(n57701), .B(n49447), .X(n38377) );
  nand_x1_sg U66861 ( .A(n51951), .B(n57764), .X(n38378) );
  nand_x1_sg U66862 ( .A(n57702), .B(n49443), .X(n38381) );
  nand_x1_sg U66863 ( .A(n51947), .B(n57764), .X(n38382) );
  nand_x1_sg U66864 ( .A(n51947), .B(n57680), .X(n38405) );
  nand_x1_sg U66865 ( .A(n48111), .B(n57754), .X(n38406) );
  nand_x1_sg U66866 ( .A(n57706), .B(n49441), .X(n38379) );
  nand_x1_sg U66867 ( .A(n51945), .B(n57760), .X(n38380) );
  nand_x1_sg U66868 ( .A(n51945), .B(n57676), .X(n38403) );
  nand_x1_sg U66869 ( .A(n48113), .B(n57770), .X(n38404) );
  nand_x1_sg U66870 ( .A(n57664), .B(n49439), .X(n37931) );
  nand_x1_sg U66871 ( .A(n51943), .B(n57763), .X(n37932) );
  nand_x1_sg U66872 ( .A(n51943), .B(n57704), .X(n38397) );
  nand_x1_sg U66873 ( .A(n48115), .B(n57764), .X(n38398) );
  nand_x1_sg U66874 ( .A(n57665), .B(n49437), .X(n37919) );
  nand_x1_sg U66875 ( .A(n51941), .B(n57766), .X(n37920) );
  nand_x1_sg U66876 ( .A(n51941), .B(n57707), .X(n38395) );
  nand_x1_sg U66877 ( .A(n48117), .B(n57746), .X(n38396) );
  nand_x1_sg U66878 ( .A(n57666), .B(n49435), .X(n37897) );
  nand_x1_sg U66879 ( .A(n51939), .B(n57747), .X(n37898) );
  nand_x1_sg U66880 ( .A(n51939), .B(n57701), .X(n38399) );
  nand_x1_sg U66881 ( .A(n48119), .B(n57756), .X(n38400) );
  nand_x1_sg U66882 ( .A(n57717), .B(n49433), .X(n38309) );
  nand_x1_sg U66883 ( .A(n51937), .B(n46200), .X(n38310) );
  nand_x1_sg U66884 ( .A(n51937), .B(n57667), .X(n37885) );
  nand_x1_sg U66885 ( .A(n48121), .B(n57743), .X(n37886) );
  nand_x1_sg U66886 ( .A(n51935), .B(n57665), .X(n37925) );
  nand_x1_sg U66887 ( .A(n48123), .B(n57766), .X(n37926) );
  nand_x1_sg U66888 ( .A(n57680), .B(n49429), .X(n37799) );
  nand_x1_sg U66889 ( .A(n51933), .B(n46200), .X(n37800) );
  nand_x1_sg U66890 ( .A(n51933), .B(n57709), .X(n38347) );
  nand_x1_sg U66891 ( .A(n48125), .B(n57762), .X(n38348) );
  nand_x1_sg U66892 ( .A(n57678), .B(n49427), .X(n38287) );
  nand_x1_sg U66893 ( .A(n51931), .B(n57755), .X(n38288) );
  nand_x1_sg U66894 ( .A(n51931), .B(n57664), .X(n37941) );
  nand_x1_sg U66895 ( .A(n48127), .B(n57759), .X(n37942) );
  nand_x1_sg U66896 ( .A(n51929), .B(n57663), .X(n37947) );
  nand_x1_sg U66897 ( .A(n48129), .B(n57772), .X(n37948) );
  nand_x1_sg U66898 ( .A(n51927), .B(n57707), .X(n38275) );
  nand_x1_sg U66899 ( .A(n48131), .B(n57755), .X(n38276) );
  nand_x1_sg U66900 ( .A(n57717), .B(n49421), .X(n38311) );
  nand_x1_sg U66901 ( .A(n51925), .B(n57735), .X(n38312) );
  nand_x1_sg U66902 ( .A(n51925), .B(n57678), .X(n38273) );
  nand_x1_sg U66903 ( .A(n48133), .B(n57771), .X(n38274) );
  nand_x1_sg U66904 ( .A(n51923), .B(n57672), .X(n38249) );
  nand_x1_sg U66905 ( .A(n48135), .B(n57765), .X(n38250) );
  nand_x1_sg U66906 ( .A(n51921), .B(n57672), .X(n38247) );
  nand_x1_sg U66907 ( .A(n48137), .B(n57760), .X(n38248) );
  nand_x1_sg U66908 ( .A(n51919), .B(n57717), .X(n38301) );
  nand_x1_sg U66909 ( .A(n48139), .B(n57750), .X(n38302) );
  nand_x1_sg U66910 ( .A(n51917), .B(n57704), .X(n38289) );
  nand_x1_sg U66911 ( .A(n48141), .B(n57770), .X(n38290) );
  nand_x1_sg U66912 ( .A(n57681), .B(n49411), .X(n38341) );
  nand_x1_sg U66913 ( .A(n51915), .B(n57761), .X(n38342) );
  nand_x1_sg U66914 ( .A(n51915), .B(n57707), .X(n38283) );
  nand_x1_sg U66915 ( .A(n48143), .B(n57770), .X(n38284) );
  nand_x1_sg U66916 ( .A(n57717), .B(n49409), .X(n38339) );
  nand_x1_sg U66917 ( .A(n51913), .B(n57762), .X(n38340) );
  nand_x1_sg U66918 ( .A(n51913), .B(n57678), .X(n38291) );
  nand_x1_sg U66919 ( .A(n48145), .B(n57747), .X(n38292) );
  nand_x1_sg U66920 ( .A(n51911), .B(n57668), .X(n37871) );
  nand_x1_sg U66921 ( .A(n48147), .B(n57744), .X(n37872) );
  nand_x1_sg U66922 ( .A(n57720), .B(n49405), .X(n37623) );
  nand_x1_sg U66923 ( .A(n51909), .B(n57744), .X(n37624) );
  nand_x1_sg U66924 ( .A(n51909), .B(n57681), .X(n37603) );
  nand_x1_sg U66925 ( .A(n48149), .B(n57748), .X(n37604) );
  nand_x1_sg U66926 ( .A(n57663), .B(n49403), .X(n37957) );
  nand_x1_sg U66927 ( .A(n51907), .B(n57761), .X(n37958) );
  nand_x1_sg U66928 ( .A(n51907), .B(n57669), .X(n37847) );
  nand_x1_sg U66929 ( .A(n48151), .B(n57759), .X(n37848) );
  nand_x1_sg U66930 ( .A(n57720), .B(n49401), .X(n37625) );
  nand_x1_sg U66931 ( .A(n51905), .B(n57766), .X(n37626) );
  nand_x1_sg U66932 ( .A(n51905), .B(n57671), .X(n37813) );
  nand_x1_sg U66933 ( .A(n48153), .B(n57750), .X(n37814) );
  nand_x1_sg U66934 ( .A(n57680), .B(n49397), .X(n37639) );
  nand_x1_sg U66935 ( .A(n51901), .B(n57766), .X(n37640) );
  nand_x1_sg U66936 ( .A(n51901), .B(n57681), .X(n37605) );
  nand_x1_sg U66937 ( .A(n48157), .B(n57745), .X(n37606) );
  nand_x1_sg U66938 ( .A(n57680), .B(n49395), .X(n37643) );
  nand_x1_sg U66939 ( .A(n51899), .B(n57756), .X(n37644) );
  nand_x1_sg U66940 ( .A(n57702), .B(n49393), .X(n38349) );
  nand_x1_sg U66941 ( .A(n51897), .B(n57756), .X(n38350) );
  nand_x1_sg U66942 ( .A(n51897), .B(n57680), .X(n37641) );
  nand_x1_sg U66943 ( .A(n48161), .B(n57744), .X(n37642) );
  nand_x1_sg U66944 ( .A(n57670), .B(n49391), .X(n37829) );
  nand_x1_sg U66945 ( .A(n51895), .B(n57761), .X(n37830) );
  nand_x1_sg U66946 ( .A(n51895), .B(n57680), .X(n37631) );
  nand_x1_sg U66947 ( .A(n48163), .B(n57761), .X(n37632) );
  nand_x1_sg U66948 ( .A(n57670), .B(n49389), .X(n37827) );
  nand_x1_sg U66949 ( .A(n51893), .B(n57764), .X(n37828) );
  nand_x1_sg U66950 ( .A(n51893), .B(n57720), .X(n37629) );
  nand_x1_sg U66951 ( .A(n48165), .B(n57760), .X(n37630) );
  nand_x1_sg U66952 ( .A(n57670), .B(n49387), .X(n37833) );
  nand_x1_sg U66953 ( .A(n51891), .B(n57772), .X(n37834) );
  nand_x1_sg U66954 ( .A(n51891), .B(n57680), .X(n37637) );
  nand_x1_sg U66955 ( .A(n48167), .B(n57758), .X(n37638) );
  nand_x1_sg U66956 ( .A(n57670), .B(n49385), .X(n37831) );
  nand_x1_sg U66957 ( .A(n51889), .B(n57764), .X(n37832) );
  nand_x1_sg U66958 ( .A(n51889), .B(n57680), .X(n37635) );
  nand_x1_sg U66959 ( .A(n48169), .B(n57770), .X(n37636) );
  nand_x1_sg U66960 ( .A(n57670), .B(n49383), .X(n37821) );
  nand_x1_sg U66961 ( .A(n51887), .B(n57750), .X(n37822) );
  nand_x1_sg U66962 ( .A(n51887), .B(n57720), .X(n37617) );
  nand_x1_sg U66963 ( .A(n48171), .B(n57775), .X(n37618) );
  nand_x1_sg U66964 ( .A(n57671), .B(n49381), .X(n37819) );
  nand_x1_sg U66965 ( .A(n51885), .B(n46200), .X(n37820) );
  nand_x1_sg U66966 ( .A(n51885), .B(n57720), .X(n37615) );
  nand_x1_sg U66967 ( .A(n48173), .B(n57761), .X(n37616) );
  nand_x1_sg U66968 ( .A(n51883), .B(n57720), .X(n37621) );
  nand_x1_sg U66969 ( .A(n48175), .B(n57749), .X(n37622) );
  nand_x1_sg U66970 ( .A(n57670), .B(n49377), .X(n37823) );
  nand_x1_sg U66971 ( .A(n51881), .B(n46197), .X(n37824) );
  nand_x1_sg U66972 ( .A(n51881), .B(n57720), .X(n37619) );
  nand_x1_sg U66973 ( .A(n48177), .B(n57750), .X(n37620) );
  nand_x1_sg U66974 ( .A(n51879), .B(n57700), .X(n37753) );
  nand_x1_sg U66975 ( .A(n48179), .B(n57775), .X(n37754) );
  nand_x1_sg U66976 ( .A(n51877), .B(n57704), .X(n38285) );
  nand_x1_sg U66977 ( .A(n48181), .B(n57758), .X(n38286) );
  nand_x1_sg U66978 ( .A(n57669), .B(n49371), .X(n37845) );
  nand_x1_sg U66979 ( .A(n51875), .B(n57735), .X(n37846) );
  nand_x1_sg U66980 ( .A(n51875), .B(n57682), .X(n38355) );
  nand_x1_sg U66981 ( .A(n48183), .B(n57757), .X(n38356) );
  nand_x1_sg U66982 ( .A(n57669), .B(n49369), .X(n37843) );
  nand_x1_sg U66983 ( .A(n51873), .B(n57748), .X(n37844) );
  nand_x1_sg U66984 ( .A(n51873), .B(n57704), .X(n38353) );
  nand_x1_sg U66985 ( .A(n48185), .B(n57765), .X(n38354) );
  nand_x1_sg U66986 ( .A(n57670), .B(n49367), .X(n37837) );
  nand_x1_sg U66987 ( .A(n51871), .B(n57744), .X(n37838) );
  nand_x1_sg U66988 ( .A(n51871), .B(n57661), .X(n37985) );
  nand_x1_sg U66989 ( .A(n48187), .B(n57764), .X(n37986) );
  nand_x1_sg U66990 ( .A(n57670), .B(n49365), .X(n37835) );
  nand_x1_sg U66991 ( .A(n51869), .B(n57743), .X(n37836) );
  nand_x1_sg U66992 ( .A(n51869), .B(n57661), .X(n37983) );
  nand_x1_sg U66993 ( .A(n48189), .B(n57770), .X(n37984) );
  nand_x1_sg U66994 ( .A(n57669), .B(n49363), .X(n37841) );
  nand_x1_sg U66995 ( .A(n51867), .B(n57740), .X(n37842) );
  nand_x1_sg U66996 ( .A(n51867), .B(n57717), .X(n38335) );
  nand_x1_sg U66997 ( .A(n48191), .B(n57761), .X(n38336) );
  nand_x1_sg U66998 ( .A(n57669), .B(n49361), .X(n37839) );
  nand_x1_sg U66999 ( .A(n51865), .B(n57743), .X(n37840) );
  nand_x1_sg U67000 ( .A(n51865), .B(n57672), .X(n38333) );
  nand_x1_sg U67001 ( .A(n48193), .B(n57736), .X(n38334) );
  nand_x1_sg U67002 ( .A(n57634), .B(n49359), .X(n37793) );
  nand_x1_sg U67003 ( .A(n51863), .B(n57757), .X(n37794) );
  nand_x1_sg U67004 ( .A(n51863), .B(n57681), .X(n37611) );
  nand_x1_sg U67005 ( .A(n48195), .B(n57750), .X(n37612) );
  nand_x1_sg U67006 ( .A(n57703), .B(n49357), .X(n37791) );
  nand_x1_sg U67007 ( .A(n51861), .B(n57766), .X(n37792) );
  nand_x1_sg U67008 ( .A(n51861), .B(n57681), .X(n37609) );
  nand_x1_sg U67009 ( .A(n48197), .B(n57743), .X(n37610) );
  nand_x1_sg U67010 ( .A(n57682), .B(n49355), .X(n37797) );
  nand_x1_sg U67011 ( .A(n51859), .B(n57747), .X(n37798) );
  nand_x1_sg U67012 ( .A(n51859), .B(n57676), .X(n38351) );
  nand_x1_sg U67013 ( .A(n48199), .B(n57760), .X(n38352) );
  nand_x1_sg U67014 ( .A(n57668), .B(n49353), .X(n37863) );
  nand_x1_sg U67015 ( .A(n51857), .B(n57744), .X(n37864) );
  nand_x1_sg U67016 ( .A(n51857), .B(n57701), .X(n37795) );
  nand_x1_sg U67017 ( .A(n48201), .B(n57763), .X(n37796) );
  nand_x1_sg U67018 ( .A(n57668), .B(n49351), .X(n37869) );
  nand_x1_sg U67019 ( .A(n51855), .B(n57763), .X(n37870) );
  nand_x1_sg U67020 ( .A(n51855), .B(n57702), .X(n37785) );
  nand_x1_sg U67021 ( .A(n48203), .B(n57748), .X(n37786) );
  nand_x1_sg U67022 ( .A(n57668), .B(n49349), .X(n37867) );
  nand_x1_sg U67023 ( .A(n51853), .B(n57766), .X(n37868) );
  nand_x1_sg U67024 ( .A(n51853), .B(n57703), .X(n37783) );
  nand_x1_sg U67025 ( .A(n48205), .B(n57773), .X(n37784) );
  nand_x1_sg U67026 ( .A(n57667), .B(n49347), .X(n37889) );
  nand_x1_sg U67027 ( .A(n51851), .B(n57743), .X(n37890) );
  nand_x1_sg U67028 ( .A(n51851), .B(n57706), .X(n37789) );
  nand_x1_sg U67029 ( .A(n48207), .B(n57765), .X(n37790) );
  nand_x1_sg U67030 ( .A(n57667), .B(n49345), .X(n37887) );
  nand_x1_sg U67031 ( .A(n51849), .B(n57743), .X(n37888) );
  nand_x1_sg U67032 ( .A(n51849), .B(n57707), .X(n37787) );
  nand_x1_sg U67033 ( .A(n48209), .B(n57766), .X(n37788) );
  nand_x1_sg U67034 ( .A(n51847), .B(n57671), .X(n37811) );
  nand_x1_sg U67035 ( .A(n48211), .B(n57749), .X(n37812) );
  nand_x1_sg U67036 ( .A(n51845), .B(n57671), .X(n37809) );
  nand_x1_sg U67037 ( .A(n48213), .B(n57770), .X(n37810) );
  nand_x1_sg U67038 ( .A(n51843), .B(n57671), .X(n37817) );
  nand_x1_sg U67039 ( .A(n48215), .B(n46200), .X(n37818) );
  nand_x1_sg U67040 ( .A(n57667), .B(n49337), .X(n37883) );
  nand_x1_sg U67041 ( .A(n51841), .B(n57742), .X(n37884) );
  nand_x1_sg U67042 ( .A(n51841), .B(n57671), .X(n37815) );
  nand_x1_sg U67043 ( .A(n48217), .B(n57766), .X(n37816) );
  nand_x1_sg U67044 ( .A(n51839), .B(n57671), .X(n37803) );
  nand_x1_sg U67045 ( .A(n48219), .B(n57773), .X(n37804) );
  nand_x1_sg U67046 ( .A(n57682), .B(n49333), .X(n37581) );
  nand_x1_sg U67047 ( .A(n51837), .B(n57749), .X(n37582) );
  nand_x1_sg U67048 ( .A(n51837), .B(n57704), .X(n37801) );
  nand_x1_sg U67049 ( .A(n48221), .B(n57770), .X(n37802) );
  nand_x1_sg U67050 ( .A(n51835), .B(n57671), .X(n37807) );
  nand_x1_sg U67051 ( .A(n48223), .B(n57747), .X(n37808) );
  nand_x1_sg U67052 ( .A(n57682), .B(n49329), .X(n37587) );
  nand_x1_sg U67053 ( .A(n51833), .B(n57750), .X(n37588) );
  nand_x1_sg U67054 ( .A(n51833), .B(n57671), .X(n37805) );
  nand_x1_sg U67055 ( .A(n48225), .B(n57771), .X(n37806) );
  nand_x1_sg U67056 ( .A(n51831), .B(n57667), .X(n37875) );
  nand_x1_sg U67057 ( .A(n48227), .B(n57749), .X(n37876) );
  nand_x1_sg U67058 ( .A(n57669), .B(n49325), .X(n37849) );
  nand_x1_sg U67059 ( .A(n51829), .B(n57743), .X(n37850) );
  nand_x1_sg U67060 ( .A(n51829), .B(n57668), .X(n37873) );
  nand_x1_sg U67061 ( .A(n48229), .B(n57750), .X(n37874) );
  nand_x1_sg U67062 ( .A(n51827), .B(n57667), .X(n37879) );
  nand_x1_sg U67063 ( .A(n48231), .B(n57742), .X(n37880) );
  nand_x1_sg U67064 ( .A(n51825), .B(n57667), .X(n37877) );
  nand_x1_sg U67065 ( .A(n48233), .B(n57764), .X(n37878) );
  nand_x1_sg U67066 ( .A(n51823), .B(n57668), .X(n37865) );
  nand_x1_sg U67067 ( .A(n48235), .B(n57748), .X(n37866) );
  nand_x1_sg U67068 ( .A(n51819), .B(n57668), .X(n37861) );
  nand_x1_sg U67069 ( .A(n47843), .B(n57744), .X(n37862) );
  nand_x1_sg U67070 ( .A(n51817), .B(n57668), .X(n37859) );
  nand_x1_sg U67071 ( .A(n47845), .B(n57758), .X(n37860) );
  nand_x1_sg U67072 ( .A(n51815), .B(n57669), .X(n37853) );
  nand_x1_sg U67073 ( .A(n47847), .B(n57740), .X(n37854) );
  nand_x1_sg U67074 ( .A(n57709), .B(n49309), .X(n37735) );
  nand_x1_sg U67075 ( .A(n51813), .B(n57754), .X(n37736) );
  nand_x1_sg U67076 ( .A(n51813), .B(n57669), .X(n37851) );
  nand_x1_sg U67077 ( .A(n47849), .B(n57741), .X(n37852) );
  nand_x1_sg U67078 ( .A(n51811), .B(n57668), .X(n37857) );
  nand_x1_sg U67079 ( .A(n47851), .B(n57765), .X(n37858) );
  nand_x1_sg U67080 ( .A(n51809), .B(n57669), .X(n37855) );
  nand_x1_sg U67081 ( .A(n47853), .B(n57761), .X(n37856) );
  nand_x1_sg U67082 ( .A(n51807), .B(n57697), .X(n37749) );
  nand_x1_sg U67083 ( .A(n47855), .B(n57763), .X(n37750) );
  nand_x1_sg U67084 ( .A(n51805), .B(n57698), .X(n37747) );
  nand_x1_sg U67085 ( .A(n47857), .B(n46198), .X(n37748) );
  nand_x1_sg U67086 ( .A(n57681), .B(n49299), .X(n37733) );
  nand_x1_sg U67087 ( .A(n51803), .B(n57775), .X(n37734) );
  nand_x1_sg U67088 ( .A(n57709), .B(n49297), .X(n37731) );
  nand_x1_sg U67089 ( .A(n51801), .B(n57775), .X(n37732) );
  nand_x1_sg U67090 ( .A(n51799), .B(n57681), .X(n37743) );
  nand_x1_sg U67091 ( .A(n47863), .B(n57750), .X(n37744) );
  nand_x1_sg U67092 ( .A(n57708), .B(n49293), .X(n37739) );
  nand_x1_sg U67093 ( .A(n51797), .B(n57756), .X(n37740) );
  nand_x1_sg U67094 ( .A(n51797), .B(n57680), .X(n37741) );
  nand_x1_sg U67095 ( .A(n47865), .B(n57773), .X(n37742) );
  nand_x1_sg U67096 ( .A(n51793), .B(n57634), .X(n37745) );
  nand_x1_sg U67097 ( .A(n47869), .B(n57763), .X(n37746) );
  nand_x1_sg U67098 ( .A(n57699), .B(n49283), .X(n37737) );
  nand_x1_sg U67099 ( .A(n51787), .B(n57759), .X(n37738) );
  nand_x1_sg U67100 ( .A(n51787), .B(n57700), .X(n37751) );
  nand_x1_sg U67101 ( .A(n47875), .B(n57771), .X(n37752) );
  nand_x1_sg U67102 ( .A(n57697), .B(n49277), .X(n37755) );
  nand_x1_sg U67103 ( .A(n51781), .B(n46197), .X(n37756) );
  nand_x1_sg U67104 ( .A(n57680), .B(n49269), .X(n37769) );
  nand_x1_sg U67105 ( .A(n51773), .B(n57760), .X(n37770) );
  nand_x1_sg U67106 ( .A(n57705), .B(n49267), .X(n37773) );
  nand_x1_sg U67107 ( .A(n51771), .B(n57755), .X(n37774) );
  nand_x1_sg U67108 ( .A(n57703), .B(n49265), .X(n37771) );
  nand_x1_sg U67109 ( .A(n51769), .B(n57754), .X(n37772) );
  nand_x1_sg U67110 ( .A(n57681), .B(n49263), .X(n37763) );
  nand_x1_sg U67111 ( .A(n51767), .B(n57764), .X(n37764) );
  nand_x1_sg U67112 ( .A(n57704), .B(n49261), .X(n37761) );
  nand_x1_sg U67113 ( .A(n51765), .B(n57748), .X(n37762) );
  nand_x1_sg U67114 ( .A(n57703), .B(n49259), .X(n37767) );
  nand_x1_sg U67115 ( .A(n51763), .B(n57758), .X(n37768) );
  nand_x1_sg U67116 ( .A(n51763), .B(n57634), .X(n37781) );
  nand_x1_sg U67117 ( .A(n47899), .B(n57759), .X(n37782) );
  nand_x1_sg U67118 ( .A(n57702), .B(n49257), .X(n37765) );
  nand_x1_sg U67119 ( .A(n51761), .B(n57763), .X(n37766) );
  nand_x1_sg U67120 ( .A(n51761), .B(n57703), .X(n37779) );
  nand_x1_sg U67121 ( .A(n47901), .B(n46200), .X(n37780) );
  nand_x1_sg U67122 ( .A(n57658), .B(n49255), .X(n38037) );
  nand_x1_sg U67123 ( .A(n51759), .B(n57762), .X(n38038) );
  nand_x1_sg U67124 ( .A(n57658), .B(n49253), .X(n38035) );
  nand_x1_sg U67125 ( .A(n51757), .B(n57771), .X(n38036) );
  nand_x1_sg U67126 ( .A(n51757), .B(n57715), .X(n37775) );
  nand_x1_sg U67127 ( .A(n47905), .B(n57764), .X(n37776) );
  nand_x1_sg U67128 ( .A(n57658), .B(n49249), .X(n38041) );
  nand_x1_sg U67129 ( .A(n51753), .B(n57748), .X(n38042) );
  nand_x1_sg U67130 ( .A(n57659), .B(n49247), .X(n38025) );
  nand_x1_sg U67131 ( .A(n51751), .B(n57764), .X(n38026) );
  nand_x1_sg U67132 ( .A(n57659), .B(n49245), .X(n38023) );
  nand_x1_sg U67133 ( .A(n51749), .B(n57756), .X(n38024) );
  nand_x1_sg U67134 ( .A(n51749), .B(n57705), .X(n37759) );
  nand_x1_sg U67135 ( .A(n47913), .B(n57726), .X(n37760) );
  nand_x1_sg U67136 ( .A(n57659), .B(n49243), .X(n38031) );
  nand_x1_sg U67137 ( .A(n51747), .B(n57749), .X(n38032) );
  nand_x1_sg U67138 ( .A(n57659), .B(n49241), .X(n38029) );
  nand_x1_sg U67139 ( .A(n51745), .B(n57750), .X(n38030) );
  nand_x1_sg U67140 ( .A(n57658), .B(n49239), .X(n38047) );
  nand_x1_sg U67141 ( .A(n51743), .B(n57762), .X(n38048) );
  nand_x1_sg U67142 ( .A(n51743), .B(n57681), .X(n37757) );
  nand_x1_sg U67143 ( .A(n47919), .B(n57764), .X(n37758) );
  nand_x1_sg U67144 ( .A(n51741), .B(n57658), .X(n38045) );
  nand_x1_sg U67145 ( .A(n47921), .B(n57770), .X(n38046) );
  nand_x1_sg U67146 ( .A(n57660), .B(n49235), .X(n38013) );
  nand_x1_sg U67147 ( .A(n51739), .B(n57772), .X(n38014) );
  nand_x1_sg U67148 ( .A(n51739), .B(n57657), .X(n38053) );
  nand_x1_sg U67149 ( .A(n47923), .B(n46200), .X(n38054) );
  nand_x1_sg U67150 ( .A(n57660), .B(n49233), .X(n38011) );
  nand_x1_sg U67151 ( .A(n51737), .B(n57773), .X(n38012) );
  nand_x1_sg U67152 ( .A(n51737), .B(n57658), .X(n38051) );
  nand_x1_sg U67153 ( .A(n47925), .B(n57772), .X(n38052) );
  nand_x1_sg U67154 ( .A(n57706), .B(n49231), .X(n38095) );
  nand_x1_sg U67155 ( .A(n51735), .B(n57731), .X(n38096) );
  nand_x1_sg U67156 ( .A(n51735), .B(n57658), .X(n38043) );
  nand_x1_sg U67157 ( .A(n47927), .B(n57772), .X(n38044) );
  nand_x1_sg U67158 ( .A(n51733), .B(n57659), .X(n38033) );
  nand_x1_sg U67159 ( .A(n47929), .B(n57746), .X(n38034) );
  nand_x1_sg U67160 ( .A(n57717), .B(n49227), .X(n38089) );
  nand_x1_sg U67161 ( .A(n51731), .B(n57733), .X(n38090) );
  nand_x1_sg U67162 ( .A(n51731), .B(n57659), .X(n38027) );
  nand_x1_sg U67163 ( .A(n47931), .B(n57748), .X(n38028) );
  nand_x1_sg U67164 ( .A(n57676), .B(n49225), .X(n38093) );
  nand_x1_sg U67165 ( .A(n51729), .B(n57757), .X(n38094) );
  nand_x1_sg U67166 ( .A(n51729), .B(n57658), .X(n38039) );
  nand_x1_sg U67167 ( .A(n47933), .B(n46201), .X(n38040) );
  nand_x1_sg U67168 ( .A(n57706), .B(n49223), .X(n38087) );
  nand_x1_sg U67169 ( .A(n51727), .B(n57746), .X(n38088) );
  nand_x1_sg U67170 ( .A(n51727), .B(n57660), .X(n38007) );
  nand_x1_sg U67171 ( .A(n47935), .B(n46197), .X(n38008) );
  nand_x1_sg U67172 ( .A(n51725), .B(n57660), .X(n38005) );
  nand_x1_sg U67173 ( .A(n47937), .B(n57763), .X(n38006) );
  nand_x1_sg U67174 ( .A(n51723), .B(n57660), .X(n38003) );
  nand_x1_sg U67175 ( .A(n47939), .B(n57744), .X(n38004) );
  nand_x1_sg U67176 ( .A(n57717), .B(n49217), .X(n38091) );
  nand_x1_sg U67177 ( .A(n51721), .B(n57726), .X(n38092) );
  nand_x1_sg U67178 ( .A(n51721), .B(n57681), .X(n37599) );
  nand_x1_sg U67179 ( .A(n47941), .B(n57746), .X(n37600) );
  nand_x1_sg U67180 ( .A(n51719), .B(n57661), .X(n37991) );
  nand_x1_sg U67181 ( .A(n47943), .B(n57756), .X(n37992) );
  nand_x1_sg U67182 ( .A(n51717), .B(n57661), .X(n37989) );
  nand_x1_sg U67183 ( .A(n47945), .B(n57775), .X(n37990) );
  nand_x1_sg U67184 ( .A(n57676), .B(n49211), .X(n38103) );
  nand_x1_sg U67185 ( .A(n51715), .B(n57763), .X(n38104) );
  nand_x1_sg U67186 ( .A(n51715), .B(n57661), .X(n37995) );
  nand_x1_sg U67187 ( .A(n47947), .B(n57760), .X(n37996) );
  nand_x1_sg U67188 ( .A(n57676), .B(n49209), .X(n38101) );
  nand_x1_sg U67189 ( .A(n51713), .B(n57727), .X(n38102) );
  nand_x1_sg U67190 ( .A(n51713), .B(n57661), .X(n37993) );
  nand_x1_sg U67191 ( .A(n47949), .B(n57771), .X(n37994) );
  nand_x1_sg U67192 ( .A(n57676), .B(n49207), .X(n38085) );
  nand_x1_sg U67193 ( .A(n51711), .B(n46201), .X(n38086) );
  nand_x1_sg U67194 ( .A(n51711), .B(n57659), .X(n38021) );
  nand_x1_sg U67195 ( .A(n47951), .B(n57763), .X(n38022) );
  nand_x1_sg U67196 ( .A(n57676), .B(n49205), .X(n38099) );
  nand_x1_sg U67197 ( .A(n51709), .B(n57724), .X(n38100) );
  nand_x1_sg U67198 ( .A(n51709), .B(n57659), .X(n38019) );
  nand_x1_sg U67199 ( .A(n47953), .B(n46201), .X(n38020) );
  nand_x1_sg U67200 ( .A(n57706), .B(n49203), .X(n38097) );
  nand_x1_sg U67201 ( .A(n51707), .B(n57725), .X(n38098) );
  nand_x1_sg U67202 ( .A(n51707), .B(n57660), .X(n38009) );
  nand_x1_sg U67203 ( .A(n47955), .B(n57764), .X(n38010) );
  nand_x1_sg U67204 ( .A(n57665), .B(n49201), .X(n38083) );
  nand_x1_sg U67205 ( .A(n51705), .B(n57771), .X(n38084) );
  nand_x1_sg U67206 ( .A(n51705), .B(n57659), .X(n38017) );
  nand_x1_sg U67207 ( .A(n47957), .B(n46198), .X(n38018) );
  nand_x1_sg U67208 ( .A(n57657), .B(n49199), .X(n38061) );
  nand_x1_sg U67209 ( .A(n51703), .B(n57765), .X(n38062) );
  nand_x1_sg U67210 ( .A(n57665), .B(n49197), .X(n37921) );
  nand_x1_sg U67211 ( .A(n51701), .B(n46201), .X(n37922) );
  nand_x1_sg U67212 ( .A(n51701), .B(n57657), .X(n38059) );
  nand_x1_sg U67213 ( .A(n47961), .B(n57766), .X(n38060) );
  nand_x1_sg U67214 ( .A(n57664), .B(n49195), .X(n37929) );
  nand_x1_sg U67215 ( .A(n51699), .B(n46197), .X(n37930) );
  nand_x1_sg U67216 ( .A(n51699), .B(n57657), .X(n38067) );
  nand_x1_sg U67217 ( .A(n47963), .B(n57747), .X(n38068) );
  nand_x1_sg U67218 ( .A(n57664), .B(n49193), .X(n37927) );
  nand_x1_sg U67219 ( .A(n51697), .B(n57762), .X(n37928) );
  nand_x1_sg U67220 ( .A(n51697), .B(n57657), .X(n38065) );
  nand_x1_sg U67221 ( .A(n47965), .B(n57747), .X(n38066) );
  nand_x1_sg U67222 ( .A(n57663), .B(n49191), .X(n37951) );
  nand_x1_sg U67223 ( .A(n51695), .B(n57749), .X(n37952) );
  nand_x1_sg U67224 ( .A(n51695), .B(n57657), .X(n38057) );
  nand_x1_sg U67225 ( .A(n47967), .B(n57750), .X(n38058) );
  nand_x1_sg U67226 ( .A(n57663), .B(n49189), .X(n37949) );
  nand_x1_sg U67227 ( .A(n51693), .B(n57762), .X(n37950) );
  nand_x1_sg U67228 ( .A(n51693), .B(n57657), .X(n38063) );
  nand_x1_sg U67229 ( .A(n47969), .B(n57759), .X(n38064) );
  nand_x1_sg U67230 ( .A(n51691), .B(n57658), .X(n38049) );
  nand_x1_sg U67231 ( .A(n47971), .B(n57764), .X(n38050) );
  nand_x1_sg U67232 ( .A(n57663), .B(n49185), .X(n37953) );
  nand_x1_sg U67233 ( .A(n51689), .B(n57750), .X(n37954) );
  nand_x1_sg U67234 ( .A(n51689), .B(n57657), .X(n38055) );
  nand_x1_sg U67235 ( .A(n47973), .B(n57770), .X(n38056) );
  nand_x1_sg U67236 ( .A(n57664), .B(n49183), .X(n37939) );
  nand_x1_sg U67237 ( .A(n51687), .B(n57764), .X(n37940) );
  nand_x1_sg U67238 ( .A(n51687), .B(n57656), .X(n38081) );
  nand_x1_sg U67239 ( .A(n47975), .B(n57771), .X(n38082) );
  nand_x1_sg U67240 ( .A(n57664), .B(n49181), .X(n37937) );
  nand_x1_sg U67241 ( .A(n51685), .B(n46198), .X(n37938) );
  nand_x1_sg U67242 ( .A(n51685), .B(n57656), .X(n38079) );
  nand_x1_sg U67243 ( .A(n47977), .B(n57762), .X(n38080) );
  nand_x1_sg U67244 ( .A(n57663), .B(n49179), .X(n37945) );
  nand_x1_sg U67245 ( .A(n51683), .B(n57749), .X(n37946) );
  nand_x1_sg U67246 ( .A(n51683), .B(n57681), .X(n37523) );
  nand_x1_sg U67247 ( .A(n47979), .B(n57744), .X(n37524) );
  nand_x1_sg U67248 ( .A(n57664), .B(n49177), .X(n37943) );
  nand_x1_sg U67249 ( .A(n51681), .B(n57771), .X(n37944) );
  nand_x1_sg U67250 ( .A(n51681), .B(n57708), .X(n37537) );
  nand_x1_sg U67251 ( .A(n47981), .B(n57773), .X(n37538) );
  nand_x1_sg U67252 ( .A(n57666), .B(n49175), .X(n37901) );
  nand_x1_sg U67253 ( .A(n51679), .B(n57761), .X(n37902) );
  nand_x1_sg U67254 ( .A(n51679), .B(n57657), .X(n38069) );
  nand_x1_sg U67255 ( .A(n47983), .B(n57772), .X(n38070) );
  nand_x1_sg U67256 ( .A(n57666), .B(n49173), .X(n37899) );
  nand_x1_sg U67257 ( .A(n51677), .B(n57746), .X(n37900) );
  nand_x1_sg U67258 ( .A(n51677), .B(n57680), .X(n37531) );
  nand_x1_sg U67259 ( .A(n47985), .B(n57744), .X(n37532) );
  nand_x1_sg U67260 ( .A(n57720), .B(n49171), .X(n37451) );
  nand_x1_sg U67261 ( .A(n51675), .B(n57735), .X(n37452) );
  nand_x1_sg U67262 ( .A(n51675), .B(n57656), .X(n38071) );
  nand_x1_sg U67263 ( .A(n47987), .B(n57764), .X(n38072) );
  nand_x1_sg U67264 ( .A(n57703), .B(n49169), .X(n37453) );
  nand_x1_sg U67265 ( .A(n51673), .B(n57765), .X(n37454) );
  nand_x1_sg U67266 ( .A(n51673), .B(n57702), .X(n37505) );
  nand_x1_sg U67267 ( .A(n47989), .B(n57757), .X(n37506) );
  nand_x1_sg U67268 ( .A(n51671), .B(n57720), .X(n37511) );
  nand_x1_sg U67269 ( .A(n47991), .B(n57747), .X(n37512) );
  nand_x1_sg U67270 ( .A(n51669), .B(n57709), .X(n37517) );
  nand_x1_sg U67271 ( .A(n47993), .B(n57772), .X(n37518) );
  nand_x1_sg U67272 ( .A(n57666), .B(n49163), .X(n37895) );
  nand_x1_sg U67273 ( .A(n51667), .B(n57756), .X(n37896) );
  nand_x1_sg U67274 ( .A(n51667), .B(n57664), .X(n37935) );
  nand_x1_sg U67275 ( .A(n47995), .B(n57765), .X(n37936) );
  nand_x1_sg U67276 ( .A(n57666), .B(n49161), .X(n37893) );
  nand_x1_sg U67277 ( .A(n51665), .B(n57763), .X(n37894) );
  nand_x1_sg U67278 ( .A(n51665), .B(n57664), .X(n37933) );
  nand_x1_sg U67279 ( .A(n47997), .B(n57763), .X(n37934) );
  nand_x1_sg U67280 ( .A(n57665), .B(n49159), .X(n37913) );
  nand_x1_sg U67281 ( .A(n51663), .B(n57744), .X(n37914) );
  nand_x1_sg U67282 ( .A(n51663), .B(n57665), .X(n37923) );
  nand_x1_sg U67283 ( .A(n47999), .B(n57757), .X(n37924) );
  nand_x1_sg U67284 ( .A(n57662), .B(n49157), .X(n37977) );
  nand_x1_sg U67285 ( .A(n51661), .B(n57758), .X(n37978) );
  nand_x1_sg U67286 ( .A(n51661), .B(n57665), .X(n37911) );
  nand_x1_sg U67287 ( .A(n48001), .B(n57754), .X(n37912) );
  nand_x1_sg U67288 ( .A(n57634), .B(n49155), .X(n37449) );
  nand_x1_sg U67289 ( .A(n51659), .B(n57748), .X(n37450) );
  nand_x1_sg U67290 ( .A(n51659), .B(n57665), .X(n37917) );
  nand_x1_sg U67291 ( .A(n48003), .B(n57755), .X(n37918) );
  nand_x1_sg U67292 ( .A(n57661), .B(n49153), .X(n37981) );
  nand_x1_sg U67293 ( .A(n51657), .B(n57766), .X(n37982) );
  nand_x1_sg U67294 ( .A(n51657), .B(n57665), .X(n37915) );
  nand_x1_sg U67295 ( .A(n48005), .B(n57745), .X(n37916) );
  nand_x1_sg U67296 ( .A(n57662), .B(n49151), .X(n37979) );
  nand_x1_sg U67297 ( .A(n51655), .B(n57760), .X(n37980) );
  nand_x1_sg U67298 ( .A(n51655), .B(n57666), .X(n37905) );
  nand_x1_sg U67299 ( .A(n48007), .B(n57757), .X(n37906) );
  nand_x1_sg U67300 ( .A(n51653), .B(n57666), .X(n37903) );
  nand_x1_sg U67301 ( .A(n48009), .B(n46197), .X(n37904) );
  nand_x1_sg U67302 ( .A(n51651), .B(n57666), .X(n37909) );
  nand_x1_sg U67303 ( .A(n48011), .B(n57760), .X(n37910) );
  nand_x1_sg U67304 ( .A(n57663), .B(n49145), .X(n37959) );
  nand_x1_sg U67305 ( .A(n51649), .B(n57773), .X(n37960) );
  nand_x1_sg U67306 ( .A(n51649), .B(n57666), .X(n37907) );
  nand_x1_sg U67307 ( .A(n48013), .B(n57748), .X(n37908) );
  nand_x1_sg U67308 ( .A(n51647), .B(n57662), .X(n37971) );
  nand_x1_sg U67309 ( .A(n48015), .B(n57761), .X(n37972) );
  nand_x1_sg U67310 ( .A(n57663), .B(n49141), .X(n37955) );
  nand_x1_sg U67311 ( .A(n51645), .B(n57764), .X(n37956) );
  nand_x1_sg U67312 ( .A(n51645), .B(n57662), .X(n37969) );
  nand_x1_sg U67313 ( .A(n48017), .B(n57761), .X(n37970) );
  nand_x1_sg U67314 ( .A(n51643), .B(n57662), .X(n37975) );
  nand_x1_sg U67315 ( .A(n48019), .B(n57773), .X(n37976) );
  nand_x1_sg U67316 ( .A(n51641), .B(n57662), .X(n37973) );
  nand_x1_sg U67317 ( .A(n48021), .B(n57761), .X(n37974) );
  nand_x1_sg U67318 ( .A(n51639), .B(n57662), .X(n37963) );
  nand_x1_sg U67319 ( .A(n48023), .B(n57757), .X(n37964) );
  nand_x1_sg U67320 ( .A(n57676), .B(n49133), .X(n38117) );
  nand_x1_sg U67321 ( .A(n51637), .B(n57762), .X(n38118) );
  nand_x1_sg U67322 ( .A(n51637), .B(n57663), .X(n37961) );
  nand_x1_sg U67323 ( .A(n48025), .B(n46201), .X(n37962) );
  nand_x1_sg U67324 ( .A(n51635), .B(n57662), .X(n37967) );
  nand_x1_sg U67325 ( .A(n48027), .B(n57747), .X(n37968) );
  nand_x1_sg U67326 ( .A(n51633), .B(n57662), .X(n37965) );
  nand_x1_sg U67327 ( .A(n48029), .B(n57770), .X(n37966) );
  nand_x1_sg U67328 ( .A(n51631), .B(n57717), .X(n38307) );
  nand_x1_sg U67329 ( .A(n48031), .B(n57759), .X(n38308) );
  nand_x1_sg U67330 ( .A(n57676), .B(n49125), .X(n38109) );
  nand_x1_sg U67331 ( .A(n51629), .B(n57763), .X(n38110) );
  nand_x1_sg U67332 ( .A(n51629), .B(n57717), .X(n38305) );
  nand_x1_sg U67333 ( .A(n48033), .B(n57761), .X(n38306) );
  nand_x1_sg U67334 ( .A(n51627), .B(n57661), .X(n37987) );
  nand_x1_sg U67335 ( .A(n48035), .B(n57763), .X(n37988) );
  nand_x1_sg U67336 ( .A(n57674), .B(n49121), .X(n38175) );
  nand_x1_sg U67337 ( .A(n51625), .B(n57742), .X(n38176) );
  nand_x1_sg U67338 ( .A(n52811), .B(n57700), .X(n36039) );
  nand_x1_sg U67339 ( .A(n48831), .B(n57742), .X(n36040) );
  nand_x1_sg U67340 ( .A(n52809), .B(n57709), .X(n36041) );
  nand_x1_sg U67341 ( .A(n48833), .B(n57744), .X(n36042) );
  nand_x1_sg U67342 ( .A(n57652), .B(n50219), .X(n36241) );
  nand_x1_sg U67343 ( .A(n52723), .B(n57770), .X(n36242) );
  nand_x1_sg U67344 ( .A(n57646), .B(n50217), .X(n36349) );
  nand_x1_sg U67345 ( .A(n52721), .B(n57770), .X(n36350) );
  nand_x1_sg U67346 ( .A(n52721), .B(n57653), .X(n36223) );
  nand_x1_sg U67347 ( .A(n48921), .B(n57761), .X(n36224) );
  nand_x1_sg U67348 ( .A(n52719), .B(n57652), .X(n36243) );
  nand_x1_sg U67349 ( .A(n48923), .B(n57773), .X(n36244) );
  nand_x1_sg U67350 ( .A(n52717), .B(n57651), .X(n36249) );
  nand_x1_sg U67351 ( .A(n48925), .B(n57759), .X(n36250) );
  nand_x1_sg U67352 ( .A(n57650), .B(n50211), .X(n36263) );
  nand_x1_sg U67353 ( .A(n52715), .B(n57772), .X(n36264) );
  nand_x1_sg U67354 ( .A(n52715), .B(n57651), .X(n36251) );
  nand_x1_sg U67355 ( .A(n48927), .B(n57760), .X(n36252) );
  nand_x1_sg U67356 ( .A(n57650), .B(n50209), .X(n36265) );
  nand_x1_sg U67357 ( .A(n52713), .B(n57765), .X(n36266) );
  nand_x1_sg U67358 ( .A(n52713), .B(n57651), .X(n36253) );
  nand_x1_sg U67359 ( .A(n48929), .B(n57775), .X(n36254) );
  nand_x1_sg U67360 ( .A(n57652), .B(n50207), .X(n36229) );
  nand_x1_sg U67361 ( .A(n52711), .B(n57762), .X(n36230) );
  nand_x1_sg U67362 ( .A(n52711), .B(n57651), .X(n36245) );
  nand_x1_sg U67363 ( .A(n48931), .B(n57762), .X(n36246) );
  nand_x1_sg U67364 ( .A(n57652), .B(n50205), .X(n36235) );
  nand_x1_sg U67365 ( .A(n52709), .B(n57760), .X(n36236) );
  nand_x1_sg U67366 ( .A(n52709), .B(n57651), .X(n36247) );
  nand_x1_sg U67367 ( .A(n48933), .B(n57765), .X(n36248) );
  nand_x1_sg U67368 ( .A(n57646), .B(n50203), .X(n36343) );
  nand_x1_sg U67369 ( .A(n52707), .B(n57773), .X(n36344) );
  nand_x1_sg U67370 ( .A(n52707), .B(n57653), .X(n36225) );
  nand_x1_sg U67371 ( .A(n48935), .B(n57757), .X(n36226) );
  nand_x1_sg U67372 ( .A(n57651), .B(n50201), .X(n36261) );
  nand_x1_sg U67373 ( .A(n52705), .B(n57749), .X(n36262) );
  nand_x1_sg U67374 ( .A(n52705), .B(n57652), .X(n36227) );
  nand_x1_sg U67375 ( .A(n48937), .B(n57758), .X(n36228) );
  nand_x1_sg U67376 ( .A(n57646), .B(n50199), .X(n36345) );
  nand_x1_sg U67377 ( .A(n52703), .B(n57770), .X(n36346) );
  nand_x1_sg U67378 ( .A(n52703), .B(n57653), .X(n36219) );
  nand_x1_sg U67379 ( .A(n48939), .B(n46197), .X(n36220) );
  nand_x1_sg U67380 ( .A(n57646), .B(n50197), .X(n36347) );
  nand_x1_sg U67381 ( .A(n52701), .B(n57773), .X(n36348) );
  nand_x1_sg U67382 ( .A(n52701), .B(n57653), .X(n36221) );
  nand_x1_sg U67383 ( .A(n48941), .B(n57763), .X(n36222) );
  nand_x1_sg U67384 ( .A(n57705), .B(n50195), .X(n36167) );
  nand_x1_sg U67385 ( .A(n52699), .B(n46198), .X(n36168) );
  nand_x1_sg U67386 ( .A(n52699), .B(n57652), .X(n36237) );
  nand_x1_sg U67387 ( .A(n48943), .B(n57758), .X(n36238) );
  nand_x1_sg U67388 ( .A(n57655), .B(n50193), .X(n36173) );
  nand_x1_sg U67389 ( .A(n52697), .B(n57749), .X(n36174) );
  nand_x1_sg U67390 ( .A(n52697), .B(n57652), .X(n36239) );
  nand_x1_sg U67391 ( .A(n48945), .B(n57771), .X(n36240) );
  nand_x1_sg U67392 ( .A(n57634), .B(n50191), .X(n36157) );
  nand_x1_sg U67393 ( .A(n52695), .B(n57770), .X(n36158) );
  nand_x1_sg U67394 ( .A(n52695), .B(n57652), .X(n36231) );
  nand_x1_sg U67395 ( .A(n48947), .B(n57771), .X(n36232) );
  nand_x1_sg U67396 ( .A(n57634), .B(n50189), .X(n36159) );
  nand_x1_sg U67397 ( .A(n52693), .B(n57775), .X(n36160) );
  nand_x1_sg U67398 ( .A(n52693), .B(n57652), .X(n36233) );
  nand_x1_sg U67399 ( .A(n48949), .B(n57775), .X(n36234) );
  nand_x1_sg U67400 ( .A(n57634), .B(n50187), .X(n36151) );
  nand_x1_sg U67401 ( .A(n52691), .B(n57761), .X(n36152) );
  nand_x1_sg U67402 ( .A(n52691), .B(n57645), .X(n36357) );
  nand_x1_sg U67403 ( .A(n48951), .B(n46197), .X(n36358) );
  nand_x1_sg U67404 ( .A(n57634), .B(n50185), .X(n36153) );
  nand_x1_sg U67405 ( .A(n52689), .B(n57763), .X(n36154) );
  nand_x1_sg U67406 ( .A(n57634), .B(n50183), .X(n36149) );
  nand_x1_sg U67407 ( .A(n52687), .B(n57766), .X(n36150) );
  nand_x1_sg U67408 ( .A(n52687), .B(n57645), .X(n36351) );
  nand_x1_sg U67409 ( .A(n48955), .B(n57759), .X(n36352) );
  nand_x1_sg U67410 ( .A(n57634), .B(n50181), .X(n36155) );
  nand_x1_sg U67411 ( .A(n52685), .B(n57764), .X(n36156) );
  nand_x1_sg U67412 ( .A(n52685), .B(n57645), .X(n36353) );
  nand_x1_sg U67413 ( .A(n48957), .B(n57775), .X(n36354) );
  nand_x1_sg U67414 ( .A(n57718), .B(n50179), .X(n36163) );
  nand_x1_sg U67415 ( .A(n52683), .B(n57770), .X(n36164) );
  nand_x1_sg U67416 ( .A(n57655), .B(n50177), .X(n36179) );
  nand_x1_sg U67417 ( .A(n52681), .B(n57764), .X(n36180) );
  nand_x1_sg U67418 ( .A(n52681), .B(n57717), .X(n36165) );
  nand_x1_sg U67419 ( .A(n48961), .B(n57758), .X(n36166) );
  nand_x1_sg U67420 ( .A(n57654), .B(n50175), .X(n36199) );
  nand_x1_sg U67421 ( .A(n52679), .B(n57743), .X(n36200) );
  nand_x1_sg U67422 ( .A(n52679), .B(n57634), .X(n36161) );
  nand_x1_sg U67423 ( .A(n48963), .B(n46197), .X(n36162) );
  nand_x1_sg U67424 ( .A(n57654), .B(n50173), .X(n36201) );
  nand_x1_sg U67425 ( .A(n52677), .B(n57748), .X(n36202) );
  nand_x1_sg U67426 ( .A(n52677), .B(n57717), .X(n36117) );
  nand_x1_sg U67427 ( .A(n48965), .B(n57764), .X(n36118) );
  nand_x1_sg U67428 ( .A(n52675), .B(n57655), .X(n36175) );
  nand_x1_sg U67429 ( .A(n48967), .B(n57748), .X(n36176) );
  nand_x1_sg U67430 ( .A(n52673), .B(n57655), .X(n36177) );
  nand_x1_sg U67431 ( .A(n48969), .B(n57763), .X(n36178) );
  nand_x1_sg U67432 ( .A(n52671), .B(n57656), .X(n36169) );
  nand_x1_sg U67433 ( .A(n48971), .B(n57747), .X(n36170) );
  nand_x1_sg U67434 ( .A(n52669), .B(n57656), .X(n36171) );
  nand_x1_sg U67435 ( .A(n48973), .B(n57775), .X(n36172) );
  nand_x1_sg U67436 ( .A(n52667), .B(n57653), .X(n36213) );
  nand_x1_sg U67437 ( .A(n48975), .B(n57761), .X(n36214) );
  nand_x1_sg U67438 ( .A(n52665), .B(n57653), .X(n36215) );
  nand_x1_sg U67439 ( .A(n48977), .B(n57764), .X(n36216) );
  nand_x1_sg U67440 ( .A(n52663), .B(n57654), .X(n36207) );
  nand_x1_sg U67441 ( .A(n48979), .B(n46201), .X(n36208) );
  nand_x1_sg U67442 ( .A(n52661), .B(n57653), .X(n36209) );
  nand_x1_sg U67443 ( .A(n48981), .B(n57764), .X(n36210) );
  nand_x1_sg U67444 ( .A(n52659), .B(n57653), .X(n36211) );
  nand_x1_sg U67445 ( .A(n48983), .B(n57749), .X(n36212) );
  nand_x1_sg U67446 ( .A(n52657), .B(n57653), .X(n36217) );
  nand_x1_sg U67447 ( .A(n48985), .B(n57772), .X(n36218) );
  nand_x1_sg U67448 ( .A(n52655), .B(n57654), .X(n36203) );
  nand_x1_sg U67449 ( .A(n48987), .B(n57760), .X(n36204) );
  nand_x1_sg U67450 ( .A(n52653), .B(n57654), .X(n36205) );
  nand_x1_sg U67451 ( .A(n48989), .B(n57762), .X(n36206) );
  nand_x1_sg U67452 ( .A(n52651), .B(n57655), .X(n36187) );
  nand_x1_sg U67453 ( .A(n48991), .B(n57765), .X(n36188) );
  nand_x1_sg U67454 ( .A(n52649), .B(n57655), .X(n36189) );
  nand_x1_sg U67455 ( .A(n48993), .B(n57762), .X(n36190) );
  nand_x1_sg U67456 ( .A(n52647), .B(n57655), .X(n36181) );
  nand_x1_sg U67457 ( .A(n48995), .B(n57750), .X(n36182) );
  nand_x1_sg U67458 ( .A(n52645), .B(n57655), .X(n36183) );
  nand_x1_sg U67459 ( .A(n48997), .B(n57765), .X(n36184) );
  nand_x1_sg U67460 ( .A(n52643), .B(n57654), .X(n36197) );
  nand_x1_sg U67461 ( .A(n48999), .B(n46201), .X(n36198) );
  nand_x1_sg U67462 ( .A(n57635), .B(n50101), .X(n35965) );
  nand_x1_sg U67463 ( .A(n52605), .B(n57747), .X(n35966) );
  nand_x1_sg U67464 ( .A(n57720), .B(n50099), .X(n35973) );
  nand_x1_sg U67465 ( .A(n52603), .B(n57747), .X(n35974) );
  nand_x1_sg U67466 ( .A(n57635), .B(n50097), .X(n35961) );
  nand_x1_sg U67467 ( .A(n52601), .B(n57747), .X(n35962) );
  nand_x1_sg U67468 ( .A(n57715), .B(n50095), .X(n35967) );
  nand_x1_sg U67469 ( .A(n52599), .B(n57747), .X(n35968) );
  nand_x1_sg U67470 ( .A(n57635), .B(n50093), .X(n35959) );
  nand_x1_sg U67471 ( .A(n52597), .B(n57747), .X(n35960) );
  nand_x1_sg U67472 ( .A(n57698), .B(n50091), .X(n36021) );
  nand_x1_sg U67473 ( .A(n52595), .B(n57756), .X(n36022) );
  nand_x1_sg U67474 ( .A(n57700), .B(n50089), .X(n36023) );
  nand_x1_sg U67475 ( .A(n52593), .B(n57749), .X(n36024) );
  nand_x1_sg U67476 ( .A(n57706), .B(n50087), .X(n36015) );
  nand_x1_sg U67477 ( .A(n52591), .B(n57756), .X(n36016) );
  nand_x1_sg U67478 ( .A(n57707), .B(n50085), .X(n36017) );
  nand_x1_sg U67479 ( .A(n52589), .B(n57756), .X(n36018) );
  nand_x1_sg U67480 ( .A(n57704), .B(n50083), .X(n36013) );
  nand_x1_sg U67481 ( .A(n52587), .B(n57756), .X(n36014) );
  nand_x1_sg U67482 ( .A(n52587), .B(n57706), .X(n35981) );
  nand_x1_sg U67483 ( .A(n48659), .B(n57746), .X(n35982) );
  nand_x1_sg U67484 ( .A(n57699), .B(n50081), .X(n36005) );
  nand_x1_sg U67485 ( .A(n52585), .B(n57745), .X(n36006) );
  nand_x1_sg U67486 ( .A(n52585), .B(n57717), .X(n35983) );
  nand_x1_sg U67487 ( .A(n48661), .B(n57746), .X(n35984) );
  nand_x1_sg U67488 ( .A(n57696), .B(n50079), .X(n36011) );
  nand_x1_sg U67489 ( .A(n52583), .B(n57756), .X(n36012) );
  nand_x1_sg U67490 ( .A(n52583), .B(n57682), .X(n35975) );
  nand_x1_sg U67491 ( .A(n48663), .B(n57746), .X(n35976) );
  nand_x1_sg U67492 ( .A(n57703), .B(n50077), .X(n35999) );
  nand_x1_sg U67493 ( .A(n52581), .B(n57745), .X(n36000) );
  nand_x1_sg U67494 ( .A(n52581), .B(n57697), .X(n35977) );
  nand_x1_sg U67495 ( .A(n48665), .B(n57746), .X(n35978) );
  nand_x1_sg U67496 ( .A(n57702), .B(n50075), .X(n35991) );
  nand_x1_sg U67497 ( .A(n52579), .B(n57745), .X(n35992) );
  nand_x1_sg U67498 ( .A(n52579), .B(n57634), .X(n35993) );
  nand_x1_sg U67499 ( .A(n48667), .B(n57745), .X(n35994) );
  nand_x1_sg U67500 ( .A(n57681), .B(n50073), .X(n35979) );
  nand_x1_sg U67501 ( .A(n52577), .B(n57746), .X(n35980) );
  nand_x1_sg U67502 ( .A(n52577), .B(n57701), .X(n35995) );
  nand_x1_sg U67503 ( .A(n48669), .B(n57745), .X(n35996) );
  nand_x1_sg U67504 ( .A(n57716), .B(n50071), .X(n35997) );
  nand_x1_sg U67505 ( .A(n52575), .B(n57745), .X(n35998) );
  nand_x1_sg U67506 ( .A(n52575), .B(n57705), .X(n35987) );
  nand_x1_sg U67507 ( .A(n48671), .B(n57746), .X(n35988) );
  nand_x1_sg U67508 ( .A(n57693), .B(n50069), .X(n35985) );
  nand_x1_sg U67509 ( .A(n52573), .B(n57746), .X(n35986) );
  nand_x1_sg U67510 ( .A(n52573), .B(n57709), .X(n35989) );
  nand_x1_sg U67511 ( .A(n48673), .B(n57746), .X(n35990) );
  nand_x1_sg U67512 ( .A(n57718), .B(n50067), .X(n36007) );
  nand_x1_sg U67513 ( .A(n52571), .B(n57756), .X(n36008) );
  nand_x1_sg U67514 ( .A(n52571), .B(n57700), .X(n35969) );
  nand_x1_sg U67515 ( .A(n48675), .B(n57747), .X(n35970) );
  nand_x1_sg U67516 ( .A(n57700), .B(n50065), .X(n36009) );
  nand_x1_sg U67517 ( .A(n52569), .B(n57756), .X(n36010) );
  nand_x1_sg U67518 ( .A(n52569), .B(n57697), .X(n35971) );
  nand_x1_sg U67519 ( .A(n48677), .B(n57747), .X(n35972) );
  nand_x1_sg U67520 ( .A(n57703), .B(n50063), .X(n36001) );
  nand_x1_sg U67521 ( .A(n52567), .B(n57745), .X(n36002) );
  nand_x1_sg U67522 ( .A(n52567), .B(n57635), .X(n35963) );
  nand_x1_sg U67523 ( .A(n48679), .B(n57747), .X(n35964) );
  nand_x1_sg U67524 ( .A(n57636), .B(n50061), .X(n35939) );
  nand_x1_sg U67525 ( .A(n52565), .B(n57749), .X(n35940) );
  nand_x1_sg U67526 ( .A(n52565), .B(n57708), .X(n36003) );
  nand_x1_sg U67527 ( .A(n48681), .B(n57745), .X(n36004) );
  nand_x1_sg U67528 ( .A(n57635), .B(n50059), .X(n35953) );
  nand_x1_sg U67529 ( .A(n52563), .B(n57750), .X(n35954) );
  nand_x1_sg U67530 ( .A(n52563), .B(n57638), .X(n35905) );
  nand_x1_sg U67531 ( .A(n48683), .B(n57744), .X(n35906) );
  nand_x1_sg U67532 ( .A(n57636), .B(n50057), .X(n35935) );
  nand_x1_sg U67533 ( .A(n52561), .B(n57760), .X(n35936) );
  nand_x1_sg U67534 ( .A(n52561), .B(n57638), .X(n35907) );
  nand_x1_sg U67535 ( .A(n48685), .B(n57750), .X(n35908) );
  nand_x1_sg U67536 ( .A(n57635), .B(n50055), .X(n35955) );
  nand_x1_sg U67537 ( .A(n52559), .B(n57748), .X(n35956) );
  nand_x1_sg U67538 ( .A(n52559), .B(n57638), .X(n35903) );
  nand_x1_sg U67539 ( .A(n48687), .B(n57748), .X(n35904) );
  nand_x1_sg U67540 ( .A(n57635), .B(n50053), .X(n35957) );
  nand_x1_sg U67541 ( .A(n52557), .B(n57742), .X(n35958) );
  nand_x1_sg U67542 ( .A(n52557), .B(n57639), .X(n35891) );
  nand_x1_sg U67543 ( .A(n48689), .B(n57748), .X(n35892) );
  nand_x1_sg U67544 ( .A(n57638), .B(n50051), .X(n35909) );
  nand_x1_sg U67545 ( .A(n52555), .B(n57749), .X(n35910) );
  nand_x1_sg U67546 ( .A(n52555), .B(n57637), .X(n35917) );
  nand_x1_sg U67547 ( .A(n48691), .B(n57773), .X(n35918) );
  nand_x1_sg U67548 ( .A(n57637), .B(n50049), .X(n35923) );
  nand_x1_sg U67549 ( .A(n52553), .B(n57770), .X(n35924) );
  nand_x1_sg U67550 ( .A(n52553), .B(n57637), .X(n35919) );
  nand_x1_sg U67551 ( .A(n48693), .B(n46198), .X(n35920) );
  nand_x1_sg U67552 ( .A(n57637), .B(n50047), .X(n35929) );
  nand_x1_sg U67553 ( .A(n52551), .B(n57771), .X(n35930) );
  nand_x1_sg U67554 ( .A(n52551), .B(n57638), .X(n35911) );
  nand_x1_sg U67555 ( .A(n48695), .B(n57773), .X(n35912) );
  nand_x1_sg U67556 ( .A(n57637), .B(n50045), .X(n35921) );
  nand_x1_sg U67557 ( .A(n52549), .B(n57762), .X(n35922) );
  nand_x1_sg U67558 ( .A(n52549), .B(n57637), .X(n35913) );
  nand_x1_sg U67559 ( .A(n48697), .B(n57749), .X(n35914) );
  nand_x1_sg U67560 ( .A(n57636), .B(n50043), .X(n35931) );
  nand_x1_sg U67561 ( .A(n52547), .B(n46198), .X(n35932) );
  nand_x1_sg U67562 ( .A(n52547), .B(n57639), .X(n35893) );
  nand_x1_sg U67563 ( .A(n48699), .B(n57748), .X(n35894) );
  nand_x1_sg U67564 ( .A(n57636), .B(n50041), .X(n35933) );
  nand_x1_sg U67565 ( .A(n52545), .B(n46198), .X(n35934) );
  nand_x1_sg U67566 ( .A(n52545), .B(n57638), .X(n35895) );
  nand_x1_sg U67567 ( .A(n48701), .B(n57747), .X(n35896) );
  nand_x1_sg U67568 ( .A(n57637), .B(n50039), .X(n35925) );
  nand_x1_sg U67569 ( .A(n52543), .B(n57749), .X(n35926) );
  nand_x1_sg U67570 ( .A(n52543), .B(n57639), .X(n35887) );
  nand_x1_sg U67571 ( .A(n48703), .B(n57748), .X(n35888) );
  nand_x1_sg U67572 ( .A(n57637), .B(n50037), .X(n35927) );
  nand_x1_sg U67573 ( .A(n52541), .B(n57770), .X(n35928) );
  nand_x1_sg U67574 ( .A(n52541), .B(n57639), .X(n35889) );
  nand_x1_sg U67575 ( .A(n48705), .B(n57748), .X(n35890) );
  nand_x1_sg U67576 ( .A(n57634), .B(n50035), .X(n36145) );
  nand_x1_sg U67577 ( .A(n52539), .B(n57770), .X(n36146) );
  nand_x1_sg U67578 ( .A(n52539), .B(n57638), .X(n35897) );
  nand_x1_sg U67579 ( .A(n48707), .B(n57764), .X(n35898) );
  nand_x1_sg U67580 ( .A(n57634), .B(n50033), .X(n36147) );
  nand_x1_sg U67581 ( .A(n52537), .B(n57759), .X(n36148) );
  nand_x1_sg U67582 ( .A(n52537), .B(n57639), .X(n35885) );
  nand_x1_sg U67583 ( .A(n48709), .B(n57748), .X(n35886) );
  nand_x1_sg U67584 ( .A(n57715), .B(n50031), .X(n36139) );
  nand_x1_sg U67585 ( .A(n52535), .B(n46197), .X(n36140) );
  nand_x1_sg U67586 ( .A(n52535), .B(n57638), .X(n35899) );
  nand_x1_sg U67587 ( .A(n48711), .B(n57765), .X(n35900) );
  nand_x1_sg U67588 ( .A(n57716), .B(n50029), .X(n36141) );
  nand_x1_sg U67589 ( .A(n52533), .B(n57770), .X(n36142) );
  nand_x1_sg U67590 ( .A(n52533), .B(n57638), .X(n35901) );
  nand_x1_sg U67591 ( .A(n48713), .B(n57746), .X(n35902) );
  nand_x1_sg U67592 ( .A(n57715), .B(n50027), .X(n36101) );
  nand_x1_sg U67593 ( .A(n52531), .B(n57743), .X(n36102) );
  nand_x1_sg U67594 ( .A(n52531), .B(n57636), .X(n35943) );
  nand_x1_sg U67595 ( .A(n48715), .B(n57771), .X(n35944) );
  nand_x1_sg U67596 ( .A(n57720), .B(n50025), .X(n36137) );
  nand_x1_sg U67597 ( .A(n52529), .B(n57770), .X(n36138) );
  nand_x1_sg U67598 ( .A(n52529), .B(n57636), .X(n35945) );
  nand_x1_sg U67599 ( .A(n48717), .B(n57748), .X(n35946) );
  nand_x1_sg U67600 ( .A(n57709), .B(n50023), .X(n36143) );
  nand_x1_sg U67601 ( .A(n52527), .B(n46198), .X(n36144) );
  nand_x1_sg U67602 ( .A(n52527), .B(n57636), .X(n35937) );
  nand_x1_sg U67603 ( .A(n48719), .B(n57750), .X(n35938) );
  nand_x1_sg U67604 ( .A(n52525), .B(n57717), .X(n36135) );
  nand_x1_sg U67605 ( .A(n48721), .B(n57762), .X(n36136) );
  nand_x1_sg U67606 ( .A(n52523), .B(n57718), .X(n36111) );
  nand_x1_sg U67607 ( .A(n48723), .B(n57748), .X(n36112) );
  nand_x1_sg U67608 ( .A(n52521), .B(n57634), .X(n36113) );
  nand_x1_sg U67609 ( .A(n48725), .B(n57770), .X(n36114) );
  nand_x1_sg U67610 ( .A(n52519), .B(n57699), .X(n36105) );
  nand_x1_sg U67611 ( .A(n48727), .B(n57747), .X(n36106) );
  nand_x1_sg U67612 ( .A(n52517), .B(n57698), .X(n36107) );
  nand_x1_sg U67613 ( .A(n48729), .B(n57749), .X(n36108) );
  nand_x1_sg U67614 ( .A(n57715), .B(n50011), .X(n36059) );
  nand_x1_sg U67615 ( .A(n52515), .B(n57744), .X(n36060) );
  nand_x1_sg U67616 ( .A(n52515), .B(n57715), .X(n36131) );
  nand_x1_sg U67617 ( .A(n48731), .B(n57749), .X(n36132) );
  nand_x1_sg U67618 ( .A(n57715), .B(n50009), .X(n36061) );
  nand_x1_sg U67619 ( .A(n52513), .B(n57742), .X(n36062) );
  nand_x1_sg U67620 ( .A(n52513), .B(n57716), .X(n36133) );
  nand_x1_sg U67621 ( .A(n48733), .B(n57750), .X(n36134) );
  nand_x1_sg U67622 ( .A(n57697), .B(n50007), .X(n36053) );
  nand_x1_sg U67623 ( .A(n52511), .B(n57742), .X(n36054) );
  nand_x1_sg U67624 ( .A(n52511), .B(n57682), .X(n36129) );
  nand_x1_sg U67625 ( .A(n48735), .B(n57757), .X(n36130) );
  nand_x1_sg U67626 ( .A(n57715), .B(n50005), .X(n36055) );
  nand_x1_sg U67627 ( .A(n52509), .B(n57744), .X(n36056) );
  nand_x1_sg U67628 ( .A(n52509), .B(n57701), .X(n36103) );
  nand_x1_sg U67629 ( .A(n48737), .B(n57750), .X(n36104) );
  nand_x1_sg U67630 ( .A(n57715), .B(n50003), .X(n36063) );
  nand_x1_sg U67631 ( .A(n52507), .B(n57742), .X(n36064) );
  nand_x1_sg U67632 ( .A(n52507), .B(n57639), .X(n35883) );
  nand_x1_sg U67633 ( .A(n48739), .B(n57748), .X(n35884) );
  nand_x1_sg U67634 ( .A(n57707), .B(n50001), .X(n36051) );
  nand_x1_sg U67635 ( .A(n52505), .B(n57744), .X(n36052) );
  nand_x1_sg U67636 ( .A(n57716), .B(n49999), .X(n36057) );
  nand_x1_sg U67637 ( .A(n52503), .B(n57744), .X(n36058) );
  nand_x1_sg U67638 ( .A(n52503), .B(n57715), .X(n36115) );
  nand_x1_sg U67639 ( .A(n48743), .B(n57748), .X(n36116) );
  nand_x1_sg U67640 ( .A(n57718), .B(n49997), .X(n36049) );
  nand_x1_sg U67641 ( .A(n52501), .B(n57742), .X(n36050) );
  nand_x1_sg U67642 ( .A(n57697), .B(n49995), .X(n36033) );
  nand_x1_sg U67643 ( .A(n52499), .B(n57743), .X(n36034) );
  nand_x1_sg U67644 ( .A(n52499), .B(n57717), .X(n36125) );
  nand_x1_sg U67645 ( .A(n48747), .B(n57772), .X(n36126) );
  nand_x1_sg U67646 ( .A(n57698), .B(n49993), .X(n36035) );
  nand_x1_sg U67647 ( .A(n52497), .B(n57766), .X(n36036) );
  nand_x1_sg U67648 ( .A(n52497), .B(n57682), .X(n36127) );
  nand_x1_sg U67649 ( .A(n48749), .B(n57764), .X(n36128) );
  nand_x1_sg U67650 ( .A(n57716), .B(n49991), .X(n36027) );
  nand_x1_sg U67651 ( .A(n52495), .B(n57742), .X(n36028) );
  nand_x1_sg U67652 ( .A(n52495), .B(n57634), .X(n36119) );
  nand_x1_sg U67653 ( .A(n48751), .B(n46200), .X(n36120) );
  nand_x1_sg U67654 ( .A(n57699), .B(n49989), .X(n36029) );
  nand_x1_sg U67655 ( .A(n52493), .B(n57744), .X(n36030) );
  nand_x1_sg U67656 ( .A(n52493), .B(n57716), .X(n36121) );
  nand_x1_sg U67657 ( .A(n48753), .B(n57748), .X(n36122) );
  nand_x1_sg U67658 ( .A(n57717), .B(n49987), .X(n36043) );
  nand_x1_sg U67659 ( .A(n52491), .B(n57744), .X(n36044) );
  nand_x1_sg U67660 ( .A(n57706), .B(n49985), .X(n36025) );
  nand_x1_sg U67661 ( .A(n52489), .B(n57743), .X(n36026) );
  nand_x1_sg U67662 ( .A(n57680), .B(n49983), .X(n36045) );
  nand_x1_sg U67663 ( .A(n52487), .B(n57742), .X(n36046) );
  nand_x1_sg U67664 ( .A(n52485), .B(n57704), .X(n36047) );
  nand_x1_sg U67665 ( .A(n48761), .B(n57744), .X(n36048) );
  nand_x1_sg U67666 ( .A(n52483), .B(n57717), .X(n36087) );
  nand_x1_sg U67667 ( .A(n48763), .B(n57743), .X(n36088) );
  nand_x1_sg U67668 ( .A(n52481), .B(n57695), .X(n36069) );
  nand_x1_sg U67669 ( .A(n48765), .B(n57742), .X(n36070) );
  nand_x1_sg U67670 ( .A(n52479), .B(n57720), .X(n36089) );
  nand_x1_sg U67671 ( .A(n48767), .B(n57743), .X(n36090) );
  nand_x1_sg U67672 ( .A(n52477), .B(n57716), .X(n36095) );
  nand_x1_sg U67673 ( .A(n48769), .B(n57743), .X(n36096) );
  nand_x1_sg U67674 ( .A(n52475), .B(n57697), .X(n36097) );
  nand_x1_sg U67675 ( .A(n48771), .B(n57743), .X(n36098) );
  nand_x1_sg U67676 ( .A(n52473), .B(n57718), .X(n36099) );
  nand_x1_sg U67677 ( .A(n48773), .B(n57743), .X(n36100) );
  nand_x1_sg U67678 ( .A(n52471), .B(n57634), .X(n36091) );
  nand_x1_sg U67679 ( .A(n48775), .B(n57743), .X(n36092) );
  nand_x1_sg U67680 ( .A(n52469), .B(n57699), .X(n36093) );
  nand_x1_sg U67681 ( .A(n48777), .B(n57743), .X(n36094) );
  nand_x1_sg U67682 ( .A(n52467), .B(n57696), .X(n36071) );
  nand_x1_sg U67683 ( .A(n48779), .B(n57744), .X(n36072) );
  nand_x1_sg U67684 ( .A(n52465), .B(n57709), .X(n36073) );
  nand_x1_sg U67685 ( .A(n48781), .B(n57744), .X(n36074) );
  nand_x1_sg U67686 ( .A(n52463), .B(n57693), .X(n36065) );
  nand_x1_sg U67687 ( .A(n48783), .B(n57744), .X(n36066) );
  nand_x1_sg U67688 ( .A(n52461), .B(n57694), .X(n36067) );
  nand_x1_sg U67689 ( .A(n48785), .B(n57742), .X(n36068) );
  nand_x1_sg U67690 ( .A(n52459), .B(n57699), .X(n36083) );
  nand_x1_sg U67691 ( .A(n48787), .B(n57744), .X(n36084) );
  nand_x1_sg U67692 ( .A(n52457), .B(n57718), .X(n36085) );
  nand_x1_sg U67693 ( .A(n48789), .B(n57744), .X(n36086) );
  nand_x1_sg U67694 ( .A(n52455), .B(n57716), .X(n36077) );
  nand_x1_sg U67695 ( .A(n48791), .B(n57744), .X(n36078) );
  nand_x1_sg U67696 ( .A(n52453), .B(n57708), .X(n36079) );
  nand_x1_sg U67697 ( .A(n48793), .B(n57744), .X(n36080) );
  nand_x1_sg U67698 ( .A(n52315), .B(n57640), .X(n35859) );
  nand_x1_sg U67699 ( .A(n48535), .B(n57750), .X(n35860) );
  nand_x1_sg U67700 ( .A(n52313), .B(n57640), .X(n35861) );
  nand_x1_sg U67701 ( .A(n48537), .B(n57750), .X(n35862) );
  nand_x1_sg U67702 ( .A(n57634), .B(n49801), .X(n36037) );
  nand_x1_sg U67703 ( .A(n52305), .B(n57746), .X(n36038) );
  nand_x1_sg U67704 ( .A(n52287), .B(n57640), .X(n35873) );
  nand_x1_sg U67705 ( .A(n48563), .B(n57749), .X(n35874) );
  nand_x1_sg U67706 ( .A(n57695), .B(n49755), .X(n35855) );
  nand_x1_sg U67707 ( .A(n52259), .B(n57750), .X(n35856) );
  nand_x1_sg U67708 ( .A(n57695), .B(n49753), .X(n35857) );
  nand_x1_sg U67709 ( .A(n52257), .B(n57750), .X(n35858) );
  nand_x1_sg U67710 ( .A(n52257), .B(n57650), .X(n36267) );
  nand_x1_sg U67711 ( .A(n48593), .B(n57775), .X(n36268) );
  nand_x1_sg U67712 ( .A(n57682), .B(n49751), .X(n35849) );
  nand_x1_sg U67713 ( .A(n52255), .B(n57750), .X(n35850) );
  nand_x1_sg U67714 ( .A(n52255), .B(n57640), .X(n35867) );
  nand_x1_sg U67715 ( .A(n48595), .B(n57749), .X(n35868) );
  nand_x1_sg U67716 ( .A(n57639), .B(n49749), .X(n35851) );
  nand_x1_sg U67717 ( .A(n52253), .B(n57750), .X(n35852) );
  nand_x1_sg U67718 ( .A(n52253), .B(n57640), .X(n35869) );
  nand_x1_sg U67719 ( .A(n48597), .B(n57749), .X(n35870) );
  nand_x1_sg U67720 ( .A(n57646), .B(n49647), .X(n36333) );
  nand_x1_sg U67721 ( .A(n52151), .B(n57759), .X(n36334) );
  nand_x1_sg U67722 ( .A(n57646), .B(n49645), .X(n36335) );
  nand_x1_sg U67723 ( .A(n52149), .B(n57758), .X(n36336) );
  nand_x1_sg U67724 ( .A(n57647), .B(n49641), .X(n36331) );
  nand_x1_sg U67725 ( .A(n52145), .B(n57759), .X(n36332) );
  nand_x1_sg U67726 ( .A(n57647), .B(n49637), .X(n36325) );
  nand_x1_sg U67727 ( .A(n52141), .B(n57758), .X(n36326) );
  nand_x1_sg U67728 ( .A(n57649), .B(n49629), .X(n36297) );
  nand_x1_sg U67729 ( .A(n52133), .B(n57763), .X(n36298) );
  nand_x1_sg U67730 ( .A(n57650), .B(n49627), .X(n36277) );
  nand_x1_sg U67731 ( .A(n52131), .B(n46198), .X(n36278) );
  nand_x1_sg U67732 ( .A(n57650), .B(n49625), .X(n36279) );
  nand_x1_sg U67733 ( .A(n52129), .B(n57772), .X(n36280) );
  nand_x1_sg U67734 ( .A(n57650), .B(n49623), .X(n36271) );
  nand_x1_sg U67735 ( .A(n52127), .B(n57762), .X(n36272) );
  nand_x1_sg U67736 ( .A(n57650), .B(n49621), .X(n36273) );
  nand_x1_sg U67737 ( .A(n52125), .B(n46197), .X(n36274) );
  nand_x1_sg U67738 ( .A(n57649), .B(n49619), .X(n36281) );
  nand_x1_sg U67739 ( .A(n52123), .B(n57758), .X(n36282) );
  nand_x1_sg U67740 ( .A(n57650), .B(n49617), .X(n36275) );
  nand_x1_sg U67741 ( .A(n52121), .B(n57771), .X(n36276) );
  nand_x1_sg U67742 ( .A(n57649), .B(n49615), .X(n36283) );
  nand_x1_sg U67743 ( .A(n52119), .B(n57747), .X(n36284) );
  nand_x1_sg U67744 ( .A(n57649), .B(n49613), .X(n36285) );
  nand_x1_sg U67745 ( .A(n52117), .B(n57765), .X(n36286) );
  nand_x1_sg U67746 ( .A(n57647), .B(n49611), .X(n36327) );
  nand_x1_sg U67747 ( .A(n52115), .B(n57775), .X(n36328) );
  nand_x1_sg U67748 ( .A(n57647), .B(n49609), .X(n36329) );
  nand_x1_sg U67749 ( .A(n52113), .B(n46197), .X(n36330) );
  nand_x1_sg U67750 ( .A(n57647), .B(n49607), .X(n36321) );
  nand_x1_sg U67751 ( .A(n52111), .B(n57759), .X(n36322) );
  nand_x1_sg U67752 ( .A(n57647), .B(n49605), .X(n36323) );
  nand_x1_sg U67753 ( .A(n52109), .B(n57758), .X(n36324) );
  nand_x1_sg U67754 ( .A(n57646), .B(n49603), .X(n36337) );
  nand_x1_sg U67755 ( .A(n52107), .B(n57770), .X(n36338) );
  nand_x1_sg U67756 ( .A(n52107), .B(n57649), .X(n36289) );
  nand_x1_sg U67757 ( .A(n48347), .B(n57770), .X(n36290) );
  nand_x1_sg U67758 ( .A(n57647), .B(n49601), .X(n36319) );
  nand_x1_sg U67759 ( .A(n52105), .B(n57760), .X(n36320) );
  nand_x1_sg U67760 ( .A(n52105), .B(n57649), .X(n36291) );
  nand_x1_sg U67761 ( .A(n48349), .B(n57758), .X(n36292) );
  nand_x1_sg U67762 ( .A(n57646), .B(n49599), .X(n36339) );
  nand_x1_sg U67763 ( .A(n52103), .B(n57773), .X(n36340) );
  nand_x1_sg U67764 ( .A(n52103), .B(n57649), .X(n36287) );
  nand_x1_sg U67765 ( .A(n48351), .B(n57747), .X(n36288) );
  nand_x1_sg U67766 ( .A(n57646), .B(n49597), .X(n36341) );
  nand_x1_sg U67767 ( .A(n52101), .B(n57764), .X(n36342) );
  nand_x1_sg U67768 ( .A(n52101), .B(n57650), .X(n36269) );
  nand_x1_sg U67769 ( .A(n48353), .B(n57772), .X(n36270) );
  nand_x1_sg U67770 ( .A(n57648), .B(n49595), .X(n36305) );
  nand_x1_sg U67771 ( .A(n52099), .B(n57761), .X(n36306) );
  nand_x1_sg U67772 ( .A(n52099), .B(n57648), .X(n36301) );
  nand_x1_sg U67773 ( .A(n48355), .B(n57766), .X(n36302) );
  nand_x1_sg U67774 ( .A(n57649), .B(n49593), .X(n36293) );
  nand_x1_sg U67775 ( .A(n52097), .B(n57748), .X(n36294) );
  nand_x1_sg U67776 ( .A(n52097), .B(n57648), .X(n36303) );
  nand_x1_sg U67777 ( .A(n48357), .B(n57760), .X(n36304) );
  nand_x1_sg U67778 ( .A(n57648), .B(n49591), .X(n36307) );
  nand_x1_sg U67779 ( .A(n52095), .B(n57762), .X(n36308) );
  nand_x1_sg U67780 ( .A(n52095), .B(n57649), .X(n36295) );
  nand_x1_sg U67781 ( .A(n48359), .B(n57758), .X(n36296) );
  nand_x1_sg U67782 ( .A(n52093), .B(n57648), .X(n36313) );
  nand_x1_sg U67783 ( .A(n48361), .B(n57761), .X(n36314) );
  nand_x1_sg U67784 ( .A(n52091), .B(n57648), .X(n36315) );
  nand_x1_sg U67785 ( .A(n48363), .B(n57760), .X(n36316) );
  nand_x1_sg U67786 ( .A(n52089), .B(n57647), .X(n36317) );
  nand_x1_sg U67787 ( .A(n48365), .B(n57761), .X(n36318) );
  nand_x1_sg U67788 ( .A(n52087), .B(n57648), .X(n36309) );
  nand_x1_sg U67789 ( .A(n48367), .B(n57775), .X(n36310) );
  nand_x1_sg U67790 ( .A(n52085), .B(n57648), .X(n36311) );
  nand_x1_sg U67791 ( .A(n48369), .B(n57760), .X(n36312) );
  nand_x1_sg U67792 ( .A(n57636), .B(n49431), .X(n35941) );
  nand_x1_sg U67793 ( .A(n51935), .B(n57746), .X(n35942) );
  nand_x1_sg U67794 ( .A(n57637), .B(n49423), .X(n35915) );
  nand_x1_sg U67795 ( .A(n51927), .B(n57775), .X(n35916) );
  nand_x1_sg U67796 ( .A(n57707), .B(n49415), .X(n36019) );
  nand_x1_sg U67797 ( .A(n51919), .B(n57756), .X(n36020) );
  nand_x1_sg U67798 ( .A(n57718), .B(n49413), .X(n36109) );
  nand_x1_sg U67799 ( .A(n51917), .B(n57775), .X(n36110) );
  nand_x1_sg U67800 ( .A(n57680), .B(n49407), .X(n36075) );
  nand_x1_sg U67801 ( .A(n51911), .B(n57744), .X(n36076) );
  nand_x1_sg U67802 ( .A(n57698), .B(n49399), .X(n36081) );
  nand_x1_sg U67803 ( .A(n51903), .B(n57744), .X(n36082) );
  nand_x1_sg U67804 ( .A(n51903), .B(n57634), .X(n36123) );
  nand_x1_sg U67805 ( .A(n48155), .B(n46201), .X(n36124) );
  nand_x1_sg U67806 ( .A(n51899), .B(n57704), .X(n36031) );
  nand_x1_sg U67807 ( .A(n48159), .B(n57765), .X(n36032) );
  nand_x1_sg U67808 ( .A(n57645), .B(n49375), .X(n36355) );
  nand_x1_sg U67809 ( .A(n51879), .B(n46198), .X(n36356) );
  nand_x1_sg U67810 ( .A(n57655), .B(n49373), .X(n36185) );
  nand_x1_sg U67811 ( .A(n51877), .B(n57762), .X(n36186) );
  nand_x1_sg U67812 ( .A(n57654), .B(n49343), .X(n36195) );
  nand_x1_sg U67813 ( .A(n51847), .B(n57749), .X(n36196) );
  nand_x1_sg U67814 ( .A(n57640), .B(n49341), .X(n35863) );
  nand_x1_sg U67815 ( .A(n51845), .B(n57749), .X(n35864) );
  nand_x1_sg U67816 ( .A(n57654), .B(n49339), .X(n36191) );
  nand_x1_sg U67817 ( .A(n51843), .B(n57749), .X(n36192) );
  nand_x1_sg U67818 ( .A(n57654), .B(n49331), .X(n36193) );
  nand_x1_sg U67819 ( .A(n51835), .B(n57759), .X(n36194) );
  nand_x1_sg U67820 ( .A(n57635), .B(n49291), .X(n35951) );
  nand_x1_sg U67821 ( .A(n51795), .B(n57755), .X(n35952) );
  nand_x1_sg U67822 ( .A(n57635), .B(n49287), .X(n35949) );
  nand_x1_sg U67823 ( .A(n51791), .B(n57765), .X(n35950) );
  nand_x1_sg U67824 ( .A(n57636), .B(n49285), .X(n35947) );
  nand_x1_sg U67825 ( .A(n51789), .B(n57766), .X(n35948) );
  nand_x1_sg U67826 ( .A(n51789), .B(n57640), .X(n35865) );
  nand_x1_sg U67827 ( .A(n47873), .B(n57749), .X(n35866) );
  nand_x1_sg U67828 ( .A(n57639), .B(n49275), .X(n35877) );
  nand_x1_sg U67829 ( .A(n51779), .B(n57749), .X(n35878) );
  nand_x1_sg U67830 ( .A(n51773), .B(n57640), .X(n35875) );
  nand_x1_sg U67831 ( .A(n47889), .B(n57749), .X(n35876) );
  nand_x1_sg U67832 ( .A(n51767), .B(n57640), .X(n35871) );
  nand_x1_sg U67833 ( .A(n47895), .B(n57749), .X(n35872) );
  nand_x1_sg U67834 ( .A(n51759), .B(n57639), .X(n35879) );
  nand_x1_sg U67835 ( .A(n47903), .B(n57748), .X(n35880) );
  nand_x1_sg U67836 ( .A(n57656), .B(n49251), .X(n35845) );
  nand_x1_sg U67837 ( .A(n51755), .B(n57750), .X(n35846) );
  nand_x1_sg U67838 ( .A(n51751), .B(n57639), .X(n35881) );
  nand_x1_sg U67839 ( .A(n47911), .B(n57748), .X(n35882) );
  nand_x1_sg U67840 ( .A(n51747), .B(n57640), .X(n35853) );
  nand_x1_sg U67841 ( .A(n47915), .B(n57750), .X(n35854) );
  nand_x1_sg U67842 ( .A(n57648), .B(n49187), .X(n36299) );
  nand_x1_sg U67843 ( .A(n51691), .B(n46197), .X(n36300) );
  nand_x1_sg U67844 ( .A(n57651), .B(n49167), .X(n36257) );
  nand_x1_sg U67845 ( .A(n51671), .B(n57750), .X(n36258) );
  nand_x1_sg U67846 ( .A(n57651), .B(n49165), .X(n36259) );
  nand_x1_sg U67847 ( .A(n51669), .B(n57748), .X(n36260) );
  nand_x1_sg U67848 ( .A(n51625), .B(n57651), .X(n36255) );
  nand_x1_sg U67849 ( .A(n48037), .B(n57749), .X(n36256) );
  nand_x1_sg U67850 ( .A(n50567), .B(n57871), .X(n30618) );
  nand_x1_sg U67851 ( .A(n57081), .B(n57907), .X(n30619) );
  nand_x1_sg U67852 ( .A(n50863), .B(n57875), .X(n29368) );
  nand_x1_sg U67853 ( .A(n57085), .B(n57910), .X(n29369) );
  nand_x1_sg U67854 ( .A(n50861), .B(n57877), .X(n29370) );
  nand_x1_sg U67855 ( .A(n57083), .B(n57910), .X(n29371) );
  nand_x1_sg U67856 ( .A(n53429), .B(n57877), .X(n29360) );
  nand_x1_sg U67857 ( .A(n51547), .B(n57909), .X(n29361) );
  nand_x1_sg U67858 ( .A(n50745), .B(n57877), .X(n29416) );
  nand_x1_sg U67859 ( .A(n57037), .B(n57886), .X(n29417) );
  nand_x1_sg U67860 ( .A(n50743), .B(n57878), .X(n29404) );
  nand_x1_sg U67861 ( .A(n57023), .B(n57898), .X(n29405) );
  nand_x1_sg U67862 ( .A(n50605), .B(n46212), .X(n29382) );
  nand_x1_sg U67863 ( .A(n56837), .B(n57907), .X(n29383) );
  nand_x1_sg U67864 ( .A(n53153), .B(n57875), .X(n29386) );
  nand_x1_sg U67865 ( .A(n51397), .B(n57909), .X(n29387) );
  nand_x1_sg U67866 ( .A(n50821), .B(n57878), .X(n29394) );
  nand_x1_sg U67867 ( .A(n56717), .B(n57895), .X(n29395) );
  nand_x1_sg U67868 ( .A(n53389), .B(n57876), .X(n29392) );
  nand_x1_sg U67869 ( .A(n51255), .B(n57886), .X(n29393) );
  nand_x1_sg U67870 ( .A(n53369), .B(n57875), .X(n29412) );
  nand_x1_sg U67871 ( .A(n47679), .B(n57904), .X(n29413) );
  nand_x1_sg U67872 ( .A(n50787), .B(n57880), .X(n29398) );
  nand_x1_sg U67873 ( .A(n56759), .B(n57887), .X(n29399) );
  nand_x1_sg U67874 ( .A(n53339), .B(n57877), .X(n29396) );
  nand_x1_sg U67875 ( .A(n51295), .B(n57910), .X(n29397) );
  nand_x1_sg U67876 ( .A(n53333), .B(n46209), .X(n29378) );
  nand_x1_sg U67877 ( .A(n47657), .B(n57899), .X(n29379) );
  nand_x1_sg U67878 ( .A(n50781), .B(n57875), .X(n29422) );
  nand_x1_sg U67879 ( .A(n56803), .B(n57909), .X(n29423) );
  nand_x1_sg U67880 ( .A(n50773), .B(n57870), .X(n29388) );
  nand_x1_sg U67881 ( .A(n56753), .B(n57899), .X(n29389) );
  nand_x1_sg U67882 ( .A(n50769), .B(n57880), .X(n29402) );
  nand_x1_sg U67883 ( .A(n56751), .B(n57898), .X(n29403) );
  nand_x1_sg U67884 ( .A(n53295), .B(n57878), .X(n29410) );
  nand_x1_sg U67885 ( .A(n51415), .B(n57908), .X(n29411) );
  nand_x1_sg U67886 ( .A(n50759), .B(n57875), .X(n29408) );
  nand_x1_sg U67887 ( .A(n56795), .B(n57886), .X(n29409) );
  nand_x1_sg U67888 ( .A(n53289), .B(n57876), .X(n29390) );
  nand_x1_sg U67889 ( .A(n51281), .B(n57896), .X(n29391) );
  nand_x1_sg U67890 ( .A(n50749), .B(n57878), .X(n29380) );
  nand_x1_sg U67891 ( .A(n56741), .B(n57900), .X(n29381) );
  nand_x1_sg U67892 ( .A(n53581), .B(n57871), .X(n30616) );
  nand_x1_sg U67893 ( .A(n47425), .B(n57907), .X(n30617) );
  nand_x1_sg U67894 ( .A(n53579), .B(n57871), .X(n30614) );
  nand_x1_sg U67895 ( .A(n47363), .B(n57898), .X(n30615) );
  nand_x1_sg U67896 ( .A(n50657), .B(n57877), .X(n29406) );
  nand_x1_sg U67897 ( .A(n56915), .B(n57887), .X(n29407) );
  nand_x1_sg U67898 ( .A(n53199), .B(n57877), .X(n29384) );
  nand_x1_sg U67899 ( .A(n51481), .B(n57907), .X(n29385) );
  nand_x1_sg U67900 ( .A(n50835), .B(n57872), .X(n29414) );
  nand_x1_sg U67901 ( .A(n56673), .B(n57898), .X(n29415) );
  nand_x1_sg U67902 ( .A(n53409), .B(n57880), .X(n29420) );
  nand_x1_sg U67903 ( .A(n51301), .B(n57910), .X(n29421) );
  nand_x1_sg U67904 ( .A(n53407), .B(n46212), .X(n29418) );
  nand_x1_sg U67905 ( .A(n47661), .B(n57886), .X(n29419) );
  nand_x1_sg U67906 ( .A(n53171), .B(n57877), .X(n29364) );
  nand_x1_sg U67907 ( .A(n51141), .B(n57908), .X(n29365) );
  nand_x1_sg U67908 ( .A(n50669), .B(n57875), .X(n29400) );
  nand_x1_sg U67909 ( .A(n55241), .B(n57896), .X(n29401) );
  nand_x1_sg U67910 ( .A(n50665), .B(n46212), .X(n29376) );
  nand_x1_sg U67911 ( .A(n55237), .B(n57900), .X(n29377) );
  nand_x1_sg U67912 ( .A(n50407), .B(n57878), .X(n29374) );
  nand_x1_sg U67913 ( .A(n55275), .B(n57909), .X(n29375) );
  nand_x1_sg U67914 ( .A(n50687), .B(n46210), .X(n29372) );
  nand_x1_sg U67915 ( .A(n55303), .B(n57907), .X(n29373) );
  nand_x1_sg U67916 ( .A(n50681), .B(n57871), .X(n30612) );
  nand_x1_sg U67917 ( .A(n55299), .B(n57911), .X(n30613) );
  nand_x1_sg U67918 ( .A(n50993), .B(n46213), .X(n30622) );
  nand_x1_sg U67919 ( .A(n55295), .B(n46207), .X(n30623) );
  nand_x1_sg U67920 ( .A(n50991), .B(n57871), .X(n30620) );
  nand_x1_sg U67921 ( .A(n55293), .B(n57908), .X(n30621) );
  nand_x1_sg U67922 ( .A(n50987), .B(n57870), .X(n30610) );
  nand_x1_sg U67923 ( .A(n55291), .B(n57909), .X(n30611) );
  nand_x1_sg U67924 ( .A(n50985), .B(n57870), .X(n30608) );
  nand_x1_sg U67925 ( .A(n55289), .B(n57908), .X(n30609) );
  nand_x1_sg U67926 ( .A(n50621), .B(n46210), .X(n29366) );
  nand_x1_sg U67927 ( .A(n55013), .B(n57910), .X(n29367) );
  nand_x1_sg U67928 ( .A(n50619), .B(n57877), .X(n29362) );
  nand_x1_sg U67929 ( .A(n55011), .B(n57895), .X(n29363) );
  nand_x1_sg U67930 ( .A(n50783), .B(n57877), .X(n29352) );
  nand_x1_sg U67931 ( .A(n56757), .B(n57909), .X(n29353) );
  nand_x1_sg U67932 ( .A(n50751), .B(n57880), .X(n29348) );
  nand_x1_sg U67933 ( .A(n56791), .B(n57886), .X(n29349) );
  nand_x1_sg U67934 ( .A(n50695), .B(n46210), .X(n29358) );
  nand_x1_sg U67935 ( .A(n56933), .B(n57907), .X(n29359) );
  nand_x1_sg U67936 ( .A(n50689), .B(n46210), .X(n29356) );
  nand_x1_sg U67937 ( .A(n56927), .B(n57907), .X(n29357) );
  nand_x1_sg U67938 ( .A(n53237), .B(n57884), .X(n29354) );
  nand_x1_sg U67939 ( .A(n47431), .B(n57907), .X(n29355) );
  nand_x1_sg U67940 ( .A(n50833), .B(n57878), .X(n29344) );
  nand_x1_sg U67941 ( .A(n56835), .B(n57896), .X(n29345) );
  nand_x1_sg U67942 ( .A(n53401), .B(n57880), .X(n29350) );
  nand_x1_sg U67943 ( .A(n51299), .B(n57907), .X(n29351) );
  nand_x4_sg U67944 ( .A(n40225), .B(n40226), .X(n39839) );
  nor_x1_sg U67945 ( .A(n47437), .B(n47353), .X(n40226) );
  nor_x1_sg U67946 ( .A(n57168), .B(n68270), .X(n40225) );
  nand_x1_sg U67947 ( .A(n50309), .B(n57533), .X(n35387) );
  nand_x1_sg U67948 ( .A(n56595), .B(n57810), .X(n35388) );
  nand_x1_sg U67949 ( .A(n50311), .B(n57552), .X(n35381) );
  nand_x1_sg U67950 ( .A(n56593), .B(n57811), .X(n35382) );
  nand_x1_sg U67951 ( .A(n50313), .B(n57553), .X(n35371) );
  nand_x1_sg U67952 ( .A(n56591), .B(n57811), .X(n35372) );
  nand_x1_sg U67953 ( .A(n50315), .B(n57535), .X(n35365) );
  nand_x1_sg U67954 ( .A(n56589), .B(n57812), .X(n35366) );
  nand_x1_sg U67955 ( .A(n50317), .B(n57533), .X(n35323) );
  nand_x1_sg U67956 ( .A(n56587), .B(n57814), .X(n35324) );
  nand_x1_sg U67957 ( .A(n50321), .B(n57554), .X(n35317) );
  nand_x1_sg U67958 ( .A(n56583), .B(n57815), .X(n35318) );
  nand_x1_sg U67959 ( .A(n50323), .B(n57554), .X(n35311) );
  nand_x1_sg U67960 ( .A(n56581), .B(n57815), .X(n35312) );
  nand_x1_sg U67961 ( .A(n50325), .B(n57536), .X(n35359) );
  nand_x1_sg U67962 ( .A(n56579), .B(n57812), .X(n35360) );
  nand_x1_sg U67963 ( .A(n50327), .B(n57537), .X(n35353) );
  nand_x1_sg U67964 ( .A(n56577), .B(n57812), .X(n35354) );
  nand_x1_sg U67965 ( .A(n50329), .B(n57551), .X(n35337) );
  nand_x1_sg U67966 ( .A(n56575), .B(n57813), .X(n35338) );
  nand_x1_sg U67967 ( .A(n50331), .B(n57550), .X(n35333) );
  nand_x1_sg U67968 ( .A(n56573), .B(n57814), .X(n35334) );
  nand_x1_sg U67969 ( .A(n50333), .B(n57553), .X(n35209) );
  nand_x1_sg U67970 ( .A(n56571), .B(n57809), .X(n35210) );
  nand_x1_sg U67971 ( .A(n50335), .B(n57550), .X(n35197) );
  nand_x1_sg U67972 ( .A(n56569), .B(n57846), .X(n35198) );
  nand_x1_sg U67973 ( .A(n50337), .B(n57550), .X(n35399) );
  nand_x1_sg U67974 ( .A(n56567), .B(n57810), .X(n35400) );
  nand_x1_sg U67975 ( .A(n50339), .B(n57533), .X(n35393) );
  nand_x1_sg U67976 ( .A(n56565), .B(n57810), .X(n35394) );
  nand_x1_sg U67977 ( .A(n50341), .B(n57534), .X(n35283) );
  nand_x1_sg U67978 ( .A(n56563), .B(n57817), .X(n35284) );
  nand_x1_sg U67979 ( .A(n50343), .B(n57552), .X(n35295) );
  nand_x1_sg U67980 ( .A(n56561), .B(n57816), .X(n35296) );
  nand_x1_sg U67981 ( .A(n50345), .B(n57552), .X(n35281) );
  nand_x1_sg U67982 ( .A(n56559), .B(n57817), .X(n35282) );
  nand_x1_sg U67983 ( .A(n50347), .B(n57557), .X(n35275) );
  nand_x1_sg U67984 ( .A(n56557), .B(n57817), .X(n35276) );
  nand_x1_sg U67985 ( .A(n50349), .B(n57539), .X(n34917) );
  nand_x1_sg U67986 ( .A(n56555), .B(n57844), .X(n34918) );
  nand_x1_sg U67987 ( .A(n50351), .B(n57539), .X(n34911) );
  nand_x1_sg U67988 ( .A(n56553), .B(n57825), .X(n34912) );
  nand_x1_sg U67989 ( .A(n50353), .B(n57539), .X(n34905) );
  nand_x1_sg U67990 ( .A(n56551), .B(n57824), .X(n34906) );
  nand_x1_sg U67991 ( .A(n50355), .B(n57540), .X(n34899) );
  nand_x1_sg U67992 ( .A(n56549), .B(n57846), .X(n34900) );
  nand_x1_sg U67993 ( .A(n50357), .B(n57537), .X(n34941) );
  nand_x1_sg U67994 ( .A(n56547), .B(n57840), .X(n34942) );
  nand_x1_sg U67995 ( .A(n50359), .B(n57537), .X(n34953) );
  nand_x1_sg U67996 ( .A(n56545), .B(n57842), .X(n34954) );
  nand_x1_sg U67997 ( .A(n50361), .B(n57538), .X(n34935) );
  nand_x1_sg U67998 ( .A(n56543), .B(n57821), .X(n34936) );
  nand_x1_sg U67999 ( .A(n50363), .B(n57538), .X(n34929) );
  nand_x1_sg U68000 ( .A(n56541), .B(n57836), .X(n34930) );
  nand_x1_sg U68001 ( .A(n50365), .B(n57537), .X(n34985) );
  nand_x1_sg U68002 ( .A(n56539), .B(n46204), .X(n34986) );
  nand_x1_sg U68003 ( .A(n50367), .B(n57536), .X(n34979) );
  nand_x1_sg U68004 ( .A(n56537), .B(n57846), .X(n34980) );
  nand_x1_sg U68005 ( .A(n50369), .B(n57533), .X(n34973) );
  nand_x1_sg U68006 ( .A(n56535), .B(n57844), .X(n34974) );
  nand_x1_sg U68007 ( .A(n50371), .B(n57554), .X(n34969) );
  nand_x1_sg U68008 ( .A(n56533), .B(n57845), .X(n34970) );
  nand_x1_sg U68009 ( .A(n50373), .B(n57541), .X(n34881) );
  nand_x1_sg U68010 ( .A(n56531), .B(n57821), .X(n34882) );
  nand_x1_sg U68011 ( .A(n50375), .B(n57550), .X(n34875) );
  nand_x1_sg U68012 ( .A(n56529), .B(n57821), .X(n34876) );
  nand_x1_sg U68013 ( .A(n50377), .B(n57535), .X(n35021) );
  nand_x1_sg U68014 ( .A(n56527), .B(n57822), .X(n35022) );
  nand_x1_sg U68015 ( .A(n50385), .B(n57552), .X(n34863) );
  nand_x1_sg U68016 ( .A(n56519), .B(n57844), .X(n34864) );
  nand_x1_sg U68017 ( .A(n50387), .B(n57541), .X(n34857) );
  nand_x1_sg U68018 ( .A(n56517), .B(n57821), .X(n34858) );
  nand_x1_sg U68019 ( .A(n50389), .B(n57553), .X(n34821) );
  nand_x1_sg U68020 ( .A(n56515), .B(n57824), .X(n34822) );
  nand_x1_sg U68021 ( .A(n50391), .B(n57557), .X(n34815) );
  nand_x1_sg U68022 ( .A(n56513), .B(n57824), .X(n34816) );
  nand_x1_sg U68023 ( .A(n50393), .B(n57541), .X(n34809) );
  nand_x1_sg U68024 ( .A(n56511), .B(n57824), .X(n34810) );
  nand_x1_sg U68025 ( .A(n50395), .B(n57541), .X(n34803) );
  nand_x1_sg U68026 ( .A(n56509), .B(n57846), .X(n34804) );
  nand_x1_sg U68027 ( .A(n50397), .B(n57536), .X(n35027) );
  nand_x1_sg U68028 ( .A(n56507), .B(n57824), .X(n35028) );
  nand_x1_sg U68029 ( .A(n50115), .B(n57534), .X(n34827) );
  nand_x1_sg U68030 ( .A(n56499), .B(n57823), .X(n34828) );
  nand_x1_sg U68031 ( .A(n50117), .B(n57541), .X(n34839) );
  nand_x1_sg U68032 ( .A(n56497), .B(n57823), .X(n34840) );
  nand_x1_sg U68033 ( .A(n50123), .B(n57534), .X(n35139) );
  nand_x1_sg U68034 ( .A(n56491), .B(n57799), .X(n35140) );
  nand_x1_sg U68035 ( .A(n50125), .B(n57554), .X(n35133) );
  nand_x1_sg U68036 ( .A(n56489), .B(n57844), .X(n35134) );
  nand_x1_sg U68037 ( .A(n50127), .B(n57533), .X(n35127) );
  nand_x1_sg U68038 ( .A(n56487), .B(n57800), .X(n35128) );
  nand_x1_sg U68039 ( .A(n50129), .B(n57534), .X(n35121) );
  nand_x1_sg U68040 ( .A(n56485), .B(n57796), .X(n35122) );
  nand_x1_sg U68041 ( .A(n50131), .B(n57537), .X(n35163) );
  nand_x1_sg U68042 ( .A(n56483), .B(n57845), .X(n35164) );
  nand_x1_sg U68043 ( .A(n50133), .B(n57551), .X(n35175) );
  nand_x1_sg U68044 ( .A(n56481), .B(n57844), .X(n35176) );
  nand_x1_sg U68045 ( .A(n50135), .B(n57550), .X(n35157) );
  nand_x1_sg U68046 ( .A(n56479), .B(n57850), .X(n35158) );
  nand_x1_sg U68047 ( .A(n50137), .B(n57553), .X(n35151) );
  nand_x1_sg U68048 ( .A(n56477), .B(n57827), .X(n35152) );
  nand_x1_sg U68049 ( .A(n50139), .B(n57551), .X(n35233) );
  nand_x1_sg U68050 ( .A(n56475), .B(n57820), .X(n35234) );
  nand_x1_sg U68051 ( .A(n50143), .B(n57550), .X(n35229) );
  nand_x1_sg U68052 ( .A(n56471), .B(n57820), .X(n35230) );
  nand_x1_sg U68053 ( .A(n50145), .B(n57558), .X(n35225) );
  nand_x1_sg U68054 ( .A(n56469), .B(n57820), .X(n35226) );
  nand_x1_sg U68055 ( .A(n50147), .B(n57554), .X(n35269) );
  nand_x1_sg U68056 ( .A(n56467), .B(n57818), .X(n35270) );
  nand_x1_sg U68057 ( .A(n50149), .B(n57550), .X(n35257) );
  nand_x1_sg U68058 ( .A(n56465), .B(n57818), .X(n35258) );
  nand_x1_sg U68059 ( .A(n50151), .B(n57553), .X(n35219) );
  nand_x1_sg U68060 ( .A(n56463), .B(n57806), .X(n35220) );
  nand_x1_sg U68061 ( .A(n50153), .B(n57554), .X(n35203) );
  nand_x1_sg U68062 ( .A(n56461), .B(n57839), .X(n35204) );
  nand_x1_sg U68063 ( .A(n50155), .B(n57554), .X(n35115) );
  nand_x1_sg U68064 ( .A(n56459), .B(n57827), .X(n35116) );
  nand_x1_sg U68065 ( .A(n50159), .B(n57533), .X(n35109) );
  nand_x1_sg U68066 ( .A(n56455), .B(n57824), .X(n35110) );
  nand_x1_sg U68067 ( .A(n50161), .B(n57554), .X(n35103) );
  nand_x1_sg U68068 ( .A(n56453), .B(n57845), .X(n35104) );
  nand_x1_sg U68069 ( .A(n50163), .B(n57537), .X(n35015) );
  nand_x1_sg U68070 ( .A(n56451), .B(n57826), .X(n35016) );
  nand_x1_sg U68071 ( .A(n50165), .B(n57535), .X(n35009) );
  nand_x1_sg U68072 ( .A(n56449), .B(n57849), .X(n35010) );
  nand_x1_sg U68073 ( .A(n50167), .B(n57536), .X(n34997) );
  nand_x1_sg U68074 ( .A(n56447), .B(n57846), .X(n34998) );
  nand_x1_sg U68075 ( .A(n50169), .B(n57537), .X(n34991) );
  nand_x1_sg U68076 ( .A(n56445), .B(n57836), .X(n34992) );
  nand_x1_sg U68077 ( .A(n50171), .B(n57550), .X(n35049) );
  nand_x1_sg U68078 ( .A(n56443), .B(n57824), .X(n35050) );
  nand_x1_sg U68079 ( .A(n50173), .B(n57551), .X(n35045) );
  nand_x1_sg U68080 ( .A(n56441), .B(n57824), .X(n35046) );
  nand_x1_sg U68081 ( .A(n50175), .B(n57533), .X(n35039) );
  nand_x1_sg U68082 ( .A(n56439), .B(n57850), .X(n35040) );
  nand_x1_sg U68083 ( .A(n50177), .B(n57551), .X(n35033) );
  nand_x1_sg U68084 ( .A(n56437), .B(n46204), .X(n35034) );
  nand_x1_sg U68085 ( .A(n50179), .B(n57554), .X(n35073) );
  nand_x1_sg U68086 ( .A(n56435), .B(n57795), .X(n35074) );
  nand_x1_sg U68087 ( .A(n50181), .B(n57553), .X(n35085) );
  nand_x1_sg U68088 ( .A(n56433), .B(n46204), .X(n35086) );
  nand_x1_sg U68089 ( .A(n50183), .B(n57551), .X(n35067) );
  nand_x1_sg U68090 ( .A(n56431), .B(n57836), .X(n35068) );
  nand_x1_sg U68091 ( .A(n50185), .B(n57550), .X(n35061) );
  nand_x1_sg U68092 ( .A(n56429), .B(n57813), .X(n35062) );
  nand_x1_sg U68093 ( .A(n50271), .B(n57554), .X(n34699) );
  nand_x1_sg U68094 ( .A(n56343), .B(n57823), .X(n34700) );
  nand_x1_sg U68095 ( .A(n50273), .B(n57533), .X(n34697) );
  nand_x1_sg U68096 ( .A(n56341), .B(n57822), .X(n34698) );
  nand_x1_sg U68097 ( .A(n49939), .B(n57536), .X(n35487) );
  nand_x1_sg U68098 ( .A(n56279), .B(n57839), .X(n35488) );
  nand_x1_sg U68099 ( .A(n49941), .B(n57550), .X(n35485) );
  nand_x1_sg U68100 ( .A(n56277), .B(n57795), .X(n35486) );
  nand_x1_sg U68101 ( .A(n49947), .B(n57533), .X(n35499) );
  nand_x1_sg U68102 ( .A(n56271), .B(n57804), .X(n35500) );
  nand_x1_sg U68103 ( .A(n49949), .B(n57552), .X(n35497) );
  nand_x1_sg U68104 ( .A(n56269), .B(n57804), .X(n35498) );
  nand_x1_sg U68105 ( .A(n49951), .B(n57553), .X(n35505) );
  nand_x1_sg U68106 ( .A(n56267), .B(n57804), .X(n35506) );
  nand_x1_sg U68107 ( .A(n49953), .B(n57534), .X(n35503) );
  nand_x1_sg U68108 ( .A(n56265), .B(n57804), .X(n35504) );
  nand_x1_sg U68109 ( .A(n49959), .B(n57553), .X(n35247) );
  nand_x1_sg U68110 ( .A(n56259), .B(n57819), .X(n35248) );
  nand_x1_sg U68111 ( .A(n49961), .B(n57550), .X(n35237) );
  nand_x1_sg U68112 ( .A(n56257), .B(n57820), .X(n35238) );
  nand_x1_sg U68113 ( .A(n49963), .B(n57554), .X(n35213) );
  nand_x1_sg U68114 ( .A(n56255), .B(n57807), .X(n35214) );
  nand_x1_sg U68115 ( .A(n49965), .B(n57554), .X(n35417) );
  nand_x1_sg U68116 ( .A(n56253), .B(n57808), .X(n35418) );
  nand_x1_sg U68117 ( .A(n49971), .B(n57558), .X(n35263) );
  nand_x1_sg U68118 ( .A(n56247), .B(n57818), .X(n35264) );
  nand_x1_sg U68119 ( .A(n50047), .B(n57534), .X(n35047) );
  nand_x1_sg U68120 ( .A(n56171), .B(n46204), .X(n35048) );
  nand_x1_sg U68121 ( .A(n50051), .B(n57551), .X(n35053) );
  nand_x1_sg U68122 ( .A(n56167), .B(n57810), .X(n35054) );
  nand_x1_sg U68123 ( .A(n50053), .B(n57552), .X(n35051) );
  nand_x1_sg U68124 ( .A(n56165), .B(n57811), .X(n35052) );
  nand_x1_sg U68125 ( .A(n50055), .B(n57554), .X(n35037) );
  nand_x1_sg U68126 ( .A(n56163), .B(n57850), .X(n35038) );
  nand_x1_sg U68127 ( .A(n50057), .B(n57538), .X(n35035) );
  nand_x1_sg U68128 ( .A(n56161), .B(n46204), .X(n35036) );
  nand_x1_sg U68129 ( .A(n50059), .B(n57551), .X(n35043) );
  nand_x1_sg U68130 ( .A(n56159), .B(n57824), .X(n35044) );
  nand_x1_sg U68131 ( .A(n50061), .B(n57550), .X(n35041) );
  nand_x1_sg U68132 ( .A(n56157), .B(n57825), .X(n35042) );
  nand_x1_sg U68133 ( .A(n50063), .B(n57534), .X(n35071) );
  nand_x1_sg U68134 ( .A(n56155), .B(n57836), .X(n35072) );
  nand_x1_sg U68135 ( .A(n50065), .B(n57552), .X(n35069) );
  nand_x1_sg U68136 ( .A(n56153), .B(n57819), .X(n35070) );
  nand_x1_sg U68137 ( .A(n50067), .B(n57534), .X(n35077) );
  nand_x1_sg U68138 ( .A(n56151), .B(n57836), .X(n35078) );
  nand_x1_sg U68139 ( .A(n50069), .B(n57553), .X(n35075) );
  nand_x1_sg U68140 ( .A(n56149), .B(n57827), .X(n35076) );
  nand_x1_sg U68141 ( .A(n50071), .B(n57553), .X(n35059) );
  nand_x1_sg U68142 ( .A(n56147), .B(n57815), .X(n35060) );
  nand_x1_sg U68143 ( .A(n50073), .B(n57550), .X(n35057) );
  nand_x1_sg U68144 ( .A(n56145), .B(n57816), .X(n35058) );
  nand_x1_sg U68145 ( .A(n50075), .B(n57550), .X(n35065) );
  nand_x1_sg U68146 ( .A(n56143), .B(n57826), .X(n35066) );
  nand_x1_sg U68147 ( .A(n50077), .B(n57551), .X(n35063) );
  nand_x1_sg U68148 ( .A(n56141), .B(n57820), .X(n35064) );
  nand_x1_sg U68149 ( .A(n50079), .B(n57552), .X(n35001) );
  nand_x1_sg U68150 ( .A(n56139), .B(n57850), .X(n35002) );
  nand_x1_sg U68151 ( .A(n50081), .B(n57553), .X(n34999) );
  nand_x1_sg U68152 ( .A(n56137), .B(n57844), .X(n35000) );
  nand_x1_sg U68153 ( .A(n50083), .B(n57534), .X(n35007) );
  nand_x1_sg U68154 ( .A(n56135), .B(n57849), .X(n35008) );
  nand_x1_sg U68155 ( .A(n50085), .B(n57534), .X(n35005) );
  nand_x1_sg U68156 ( .A(n56133), .B(n57846), .X(n35006) );
  nand_x1_sg U68157 ( .A(n50087), .B(n57538), .X(n34989) );
  nand_x1_sg U68158 ( .A(n56131), .B(n57845), .X(n34990) );
  nand_x1_sg U68159 ( .A(n50089), .B(n57554), .X(n34987) );
  nand_x1_sg U68160 ( .A(n56129), .B(n46204), .X(n34988) );
  nand_x1_sg U68161 ( .A(n50091), .B(n57533), .X(n34995) );
  nand_x1_sg U68162 ( .A(n56127), .B(n46204), .X(n34996) );
  nand_x1_sg U68163 ( .A(n50093), .B(n57533), .X(n34993) );
  nand_x1_sg U68164 ( .A(n56125), .B(n57850), .X(n34994) );
  nand_x1_sg U68165 ( .A(n50095), .B(n57538), .X(n35025) );
  nand_x1_sg U68166 ( .A(n56123), .B(n57846), .X(n35026) );
  nand_x1_sg U68167 ( .A(n50097), .B(n57535), .X(n35023) );
  nand_x1_sg U68168 ( .A(n56121), .B(n57821), .X(n35024) );
  nand_x1_sg U68169 ( .A(n50099), .B(n57552), .X(n35031) );
  nand_x1_sg U68170 ( .A(n56119), .B(n57825), .X(n35032) );
  nand_x1_sg U68171 ( .A(n50101), .B(n57553), .X(n35029) );
  nand_x1_sg U68172 ( .A(n56117), .B(n57825), .X(n35030) );
  nand_x1_sg U68173 ( .A(n50103), .B(n57551), .X(n35013) );
  nand_x1_sg U68174 ( .A(n56115), .B(n57824), .X(n35014) );
  nand_x1_sg U68175 ( .A(n50105), .B(n57551), .X(n35011) );
  nand_x1_sg U68176 ( .A(n56113), .B(n57824), .X(n35012) );
  nand_x1_sg U68177 ( .A(n50107), .B(n57533), .X(n35019) );
  nand_x1_sg U68178 ( .A(n56111), .B(n57803), .X(n35020) );
  nand_x1_sg U68179 ( .A(n50109), .B(n57558), .X(n35017) );
  nand_x1_sg U68180 ( .A(n56109), .B(n57804), .X(n35018) );
  nand_x1_sg U68181 ( .A(n49715), .B(n57551), .X(n35143) );
  nand_x1_sg U68182 ( .A(n56107), .B(n57818), .X(n35144) );
  nand_x1_sg U68183 ( .A(n49717), .B(n57550), .X(n35141) );
  nand_x1_sg U68184 ( .A(n56105), .B(n57845), .X(n35142) );
  nand_x1_sg U68185 ( .A(n49719), .B(n57551), .X(n35149) );
  nand_x1_sg U68186 ( .A(n56103), .B(n57826), .X(n35150) );
  nand_x1_sg U68187 ( .A(n49721), .B(n57551), .X(n35147) );
  nand_x1_sg U68188 ( .A(n56101), .B(n57836), .X(n35148) );
  nand_x1_sg U68189 ( .A(n49723), .B(n57558), .X(n35131) );
  nand_x1_sg U68190 ( .A(n56099), .B(n57798), .X(n35132) );
  nand_x1_sg U68191 ( .A(n49725), .B(n57553), .X(n35129) );
  nand_x1_sg U68192 ( .A(n56097), .B(n57795), .X(n35130) );
  nand_x1_sg U68193 ( .A(n49727), .B(n57550), .X(n35137) );
  nand_x1_sg U68194 ( .A(n56095), .B(n57797), .X(n35138) );
  nand_x1_sg U68195 ( .A(n49729), .B(n57534), .X(n35135) );
  nand_x1_sg U68196 ( .A(n56093), .B(n57843), .X(n35136) );
  nand_x1_sg U68197 ( .A(n49731), .B(n57558), .X(n35167) );
  nand_x1_sg U68198 ( .A(n56091), .B(n57850), .X(n35168) );
  nand_x1_sg U68199 ( .A(n49733), .B(n57552), .X(n35165) );
  nand_x1_sg U68200 ( .A(n56089), .B(n57838), .X(n35166) );
  nand_x1_sg U68201 ( .A(n49735), .B(n57553), .X(n35173) );
  nand_x1_sg U68202 ( .A(n56087), .B(n57839), .X(n35174) );
  nand_x1_sg U68203 ( .A(n49737), .B(n57558), .X(n35171) );
  nand_x1_sg U68204 ( .A(n56085), .B(n57837), .X(n35172) );
  nand_x1_sg U68205 ( .A(n49739), .B(n57554), .X(n35155) );
  nand_x1_sg U68206 ( .A(n56083), .B(n57849), .X(n35156) );
  nand_x1_sg U68207 ( .A(n49741), .B(n57551), .X(n35153) );
  nand_x1_sg U68208 ( .A(n56081), .B(n57827), .X(n35154) );
  nand_x1_sg U68209 ( .A(n49743), .B(n57552), .X(n35161) );
  nand_x1_sg U68210 ( .A(n56079), .B(n57838), .X(n35162) );
  nand_x1_sg U68211 ( .A(n49745), .B(n57533), .X(n35159) );
  nand_x1_sg U68212 ( .A(n56077), .B(n57850), .X(n35160) );
  nand_x1_sg U68213 ( .A(n49747), .B(n57534), .X(n35095) );
  nand_x1_sg U68214 ( .A(n56075), .B(n57817), .X(n35096) );
  nand_x1_sg U68215 ( .A(n49749), .B(n57558), .X(n35093) );
  nand_x1_sg U68216 ( .A(n56073), .B(n57814), .X(n35094) );
  nand_x1_sg U68217 ( .A(n49751), .B(n57558), .X(n35101) );
  nand_x1_sg U68218 ( .A(n56071), .B(n57836), .X(n35102) );
  nand_x1_sg U68219 ( .A(n49753), .B(n57550), .X(n35099) );
  nand_x1_sg U68220 ( .A(n56069), .B(n57846), .X(n35100) );
  nand_x1_sg U68221 ( .A(n49755), .B(n57553), .X(n35083) );
  nand_x1_sg U68222 ( .A(n56067), .B(n57808), .X(n35084) );
  nand_x1_sg U68223 ( .A(n49757), .B(n57550), .X(n35081) );
  nand_x1_sg U68224 ( .A(n56065), .B(n57809), .X(n35082) );
  nand_x1_sg U68225 ( .A(n49759), .B(n57534), .X(n35089) );
  nand_x1_sg U68226 ( .A(n56063), .B(n57806), .X(n35090) );
  nand_x1_sg U68227 ( .A(n49761), .B(n57534), .X(n35087) );
  nand_x1_sg U68228 ( .A(n56061), .B(n57807), .X(n35088) );
  nand_x1_sg U68229 ( .A(n49763), .B(n57534), .X(n35119) );
  nand_x1_sg U68230 ( .A(n56059), .B(n57844), .X(n35120) );
  nand_x1_sg U68231 ( .A(n49765), .B(n57550), .X(n35117) );
  nand_x1_sg U68232 ( .A(n56057), .B(n57801), .X(n35118) );
  nand_x1_sg U68233 ( .A(n49767), .B(n57533), .X(n35125) );
  nand_x1_sg U68234 ( .A(n56055), .B(n57839), .X(n35126) );
  nand_x1_sg U68235 ( .A(n49769), .B(n57534), .X(n35123) );
  nand_x1_sg U68236 ( .A(n56053), .B(n57805), .X(n35124) );
  nand_x1_sg U68237 ( .A(n49771), .B(n57551), .X(n35107) );
  nand_x1_sg U68238 ( .A(n56051), .B(n57846), .X(n35108) );
  nand_x1_sg U68239 ( .A(n49773), .B(n57552), .X(n35105) );
  nand_x1_sg U68240 ( .A(n56049), .B(n57824), .X(n35106) );
  nand_x1_sg U68241 ( .A(n49775), .B(n57553), .X(n35113) );
  nand_x1_sg U68242 ( .A(n56047), .B(n57802), .X(n35114) );
  nand_x1_sg U68243 ( .A(n49777), .B(n57533), .X(n35111) );
  nand_x1_sg U68244 ( .A(n56045), .B(n57827), .X(n35112) );
  nand_x1_sg U68245 ( .A(n49779), .B(n57552), .X(n34861) );
  nand_x1_sg U68246 ( .A(n56043), .B(n57825), .X(n34862) );
  nand_x1_sg U68247 ( .A(n49781), .B(n57541), .X(n34859) );
  nand_x1_sg U68248 ( .A(n56041), .B(n57844), .X(n34860) );
  nand_x1_sg U68249 ( .A(n49783), .B(n57552), .X(n34867) );
  nand_x1_sg U68250 ( .A(n56039), .B(n57821), .X(n34868) );
  nand_x1_sg U68251 ( .A(n49785), .B(n57552), .X(n34865) );
  nand_x1_sg U68252 ( .A(n56037), .B(n57837), .X(n34866) );
  nand_x1_sg U68253 ( .A(n49787), .B(n57541), .X(n34849) );
  nand_x1_sg U68254 ( .A(n56035), .B(n57822), .X(n34850) );
  nand_x1_sg U68255 ( .A(n49789), .B(n57541), .X(n34847) );
  nand_x1_sg U68256 ( .A(n56033), .B(n57822), .X(n34848) );
  nand_x1_sg U68257 ( .A(n49791), .B(n57552), .X(n34855) );
  nand_x1_sg U68258 ( .A(n56031), .B(n57822), .X(n34856) );
  nand_x1_sg U68259 ( .A(n49793), .B(n57541), .X(n34853) );
  nand_x1_sg U68260 ( .A(n56029), .B(n57822), .X(n34854) );
  nand_x1_sg U68261 ( .A(n49795), .B(n57540), .X(n34885) );
  nand_x1_sg U68262 ( .A(n56027), .B(n57821), .X(n34886) );
  nand_x1_sg U68263 ( .A(n49797), .B(n57538), .X(n34883) );
  nand_x1_sg U68264 ( .A(n56025), .B(n57821), .X(n34884) );
  nand_x1_sg U68265 ( .A(n49799), .B(n57540), .X(n34891) );
  nand_x1_sg U68266 ( .A(n56023), .B(n57824), .X(n34892) );
  nand_x1_sg U68267 ( .A(n49801), .B(n57540), .X(n34889) );
  nand_x1_sg U68268 ( .A(n56021), .B(n57844), .X(n34890) );
  nand_x1_sg U68269 ( .A(n49803), .B(n57541), .X(n34873) );
  nand_x1_sg U68270 ( .A(n56019), .B(n57821), .X(n34874) );
  nand_x1_sg U68271 ( .A(n49805), .B(n57553), .X(n34871) );
  nand_x1_sg U68272 ( .A(n56017), .B(n57838), .X(n34872) );
  nand_x1_sg U68273 ( .A(n49807), .B(n57554), .X(n34879) );
  nand_x1_sg U68274 ( .A(n56015), .B(n57821), .X(n34880) );
  nand_x1_sg U68275 ( .A(n49809), .B(n57550), .X(n34877) );
  nand_x1_sg U68276 ( .A(n56013), .B(n57821), .X(n34878) );
  nand_x1_sg U68277 ( .A(n49811), .B(n57533), .X(n34813) );
  nand_x1_sg U68278 ( .A(n56011), .B(n57825), .X(n34814) );
  nand_x1_sg U68279 ( .A(n49813), .B(n57541), .X(n34811) );
  nand_x1_sg U68280 ( .A(n56009), .B(n57823), .X(n34812) );
  nand_x1_sg U68281 ( .A(n49815), .B(n57537), .X(n34819) );
  nand_x1_sg U68282 ( .A(n56007), .B(n57824), .X(n34820) );
  nand_x1_sg U68283 ( .A(n49817), .B(n57536), .X(n34817) );
  nand_x1_sg U68284 ( .A(n56005), .B(n57824), .X(n34818) );
  nand_x1_sg U68285 ( .A(n49819), .B(n57541), .X(n34801) );
  nand_x1_sg U68286 ( .A(n56003), .B(n57846), .X(n34802) );
  nand_x1_sg U68287 ( .A(n49821), .B(n57541), .X(n34799) );
  nand_x1_sg U68288 ( .A(n56001), .B(n57846), .X(n34800) );
  nand_x1_sg U68289 ( .A(n49823), .B(n57541), .X(n34807) );
  nand_x1_sg U68290 ( .A(n55999), .B(n57846), .X(n34808) );
  nand_x1_sg U68291 ( .A(n49825), .B(n57552), .X(n34805) );
  nand_x1_sg U68292 ( .A(n55997), .B(n57845), .X(n34806) );
  nand_x1_sg U68293 ( .A(n49827), .B(n57541), .X(n34837) );
  nand_x1_sg U68294 ( .A(n55995), .B(n57823), .X(n34838) );
  nand_x1_sg U68295 ( .A(n49829), .B(n57541), .X(n34835) );
  nand_x1_sg U68296 ( .A(n55993), .B(n57823), .X(n34836) );
  nand_x1_sg U68297 ( .A(n49831), .B(n57541), .X(n34843) );
  nand_x1_sg U68298 ( .A(n55991), .B(n57822), .X(n34844) );
  nand_x1_sg U68299 ( .A(n49833), .B(n57541), .X(n34841) );
  nand_x1_sg U68300 ( .A(n55989), .B(n57822), .X(n34842) );
  nand_x1_sg U68301 ( .A(n49835), .B(n57535), .X(n34825) );
  nand_x1_sg U68302 ( .A(n55987), .B(n57823), .X(n34826) );
  nand_x1_sg U68303 ( .A(n49837), .B(n57538), .X(n34823) );
  nand_x1_sg U68304 ( .A(n55985), .B(n57844), .X(n34824) );
  nand_x1_sg U68305 ( .A(n49839), .B(n57541), .X(n34831) );
  nand_x1_sg U68306 ( .A(n55983), .B(n57823), .X(n34832) );
  nand_x1_sg U68307 ( .A(n49841), .B(n57552), .X(n34829) );
  nand_x1_sg U68308 ( .A(n55981), .B(n57823), .X(n34830) );
  nand_x1_sg U68309 ( .A(n49843), .B(n57536), .X(n34957) );
  nand_x1_sg U68310 ( .A(n55979), .B(n57824), .X(n34958) );
  nand_x1_sg U68311 ( .A(n49845), .B(n57537), .X(n34955) );
  nand_x1_sg U68312 ( .A(n55977), .B(n57824), .X(n34956) );
  nand_x1_sg U68313 ( .A(n49847), .B(n57536), .X(n34963) );
  nand_x1_sg U68314 ( .A(n55975), .B(n57850), .X(n34964) );
  nand_x1_sg U68315 ( .A(n49849), .B(n57536), .X(n34961) );
  nand_x1_sg U68316 ( .A(n55973), .B(n57824), .X(n34962) );
  nand_x1_sg U68317 ( .A(n49851), .B(n57537), .X(n34945) );
  nand_x1_sg U68318 ( .A(n55971), .B(n57841), .X(n34946) );
  nand_x1_sg U68319 ( .A(n49853), .B(n57537), .X(n34943) );
  nand_x1_sg U68320 ( .A(n55969), .B(n57842), .X(n34944) );
  nand_x1_sg U68321 ( .A(n49855), .B(n57537), .X(n34951) );
  nand_x1_sg U68322 ( .A(n55967), .B(n57850), .X(n34952) );
  nand_x1_sg U68323 ( .A(n49857), .B(n57537), .X(n34949) );
  nand_x1_sg U68324 ( .A(n55965), .B(n57844), .X(n34950) );
  nand_x1_sg U68325 ( .A(n49859), .B(n57534), .X(n34977) );
  nand_x1_sg U68326 ( .A(n55963), .B(n46204), .X(n34978) );
  nand_x1_sg U68327 ( .A(n49861), .B(n57558), .X(n34975) );
  nand_x1_sg U68328 ( .A(n55961), .B(n46204), .X(n34976) );
  nand_x1_sg U68329 ( .A(n49863), .B(n57551), .X(n34983) );
  nand_x1_sg U68330 ( .A(n55959), .B(n57843), .X(n34984) );
  nand_x1_sg U68331 ( .A(n49865), .B(n57554), .X(n34981) );
  nand_x1_sg U68332 ( .A(n55957), .B(n57840), .X(n34982) );
  nand_x1_sg U68333 ( .A(n49867), .B(n57541), .X(n34967) );
  nand_x1_sg U68334 ( .A(n55955), .B(n57846), .X(n34968) );
  nand_x1_sg U68335 ( .A(n49871), .B(n57551), .X(n34971) );
  nand_x1_sg U68336 ( .A(n55951), .B(n57841), .X(n34972) );
  nand_x1_sg U68337 ( .A(n49875), .B(n57539), .X(n34909) );
  nand_x1_sg U68338 ( .A(n55947), .B(n57846), .X(n34910) );
  nand_x1_sg U68339 ( .A(n49877), .B(n57539), .X(n34907) );
  nand_x1_sg U68340 ( .A(n55945), .B(n57844), .X(n34908) );
  nand_x1_sg U68341 ( .A(n49879), .B(n57539), .X(n34915) );
  nand_x1_sg U68342 ( .A(n55943), .B(n57822), .X(n34916) );
  nand_x1_sg U68343 ( .A(n49881), .B(n57539), .X(n34913) );
  nand_x1_sg U68344 ( .A(n55941), .B(n57823), .X(n34914) );
  nand_x1_sg U68345 ( .A(n49883), .B(n57540), .X(n34897) );
  nand_x1_sg U68346 ( .A(n55939), .B(n57844), .X(n34898) );
  nand_x1_sg U68347 ( .A(n49885), .B(n57540), .X(n34895) );
  nand_x1_sg U68348 ( .A(n55937), .B(n57821), .X(n34896) );
  nand_x1_sg U68349 ( .A(n49887), .B(n57539), .X(n34903) );
  nand_x1_sg U68350 ( .A(n55935), .B(n57844), .X(n34904) );
  nand_x1_sg U68351 ( .A(n49889), .B(n57540), .X(n34901) );
  nand_x1_sg U68352 ( .A(n55933), .B(n57822), .X(n34902) );
  nand_x1_sg U68353 ( .A(n49891), .B(n57538), .X(n34933) );
  nand_x1_sg U68354 ( .A(n55931), .B(n57845), .X(n34934) );
  nand_x1_sg U68355 ( .A(n49893), .B(n57538), .X(n34931) );
  nand_x1_sg U68356 ( .A(n55929), .B(n57825), .X(n34932) );
  nand_x1_sg U68357 ( .A(n49895), .B(n57537), .X(n34939) );
  nand_x1_sg U68358 ( .A(n55927), .B(n57825), .X(n34940) );
  nand_x1_sg U68359 ( .A(n49897), .B(n57538), .X(n34937) );
  nand_x1_sg U68360 ( .A(n55925), .B(n57844), .X(n34938) );
  nand_x1_sg U68361 ( .A(n49899), .B(n57538), .X(n34921) );
  nand_x1_sg U68362 ( .A(n55923), .B(n57825), .X(n34922) );
  nand_x1_sg U68363 ( .A(n49901), .B(n57539), .X(n34919) );
  nand_x1_sg U68364 ( .A(n55921), .B(n57821), .X(n34920) );
  nand_x1_sg U68365 ( .A(n49903), .B(n57538), .X(n34927) );
  nand_x1_sg U68366 ( .A(n55919), .B(n57823), .X(n34928) );
  nand_x1_sg U68367 ( .A(n49905), .B(n57538), .X(n34925) );
  nand_x1_sg U68368 ( .A(n55917), .B(n57844), .X(n34926) );
  nand_x1_sg U68369 ( .A(n49907), .B(n57558), .X(n35403) );
  nand_x1_sg U68370 ( .A(n55915), .B(n57809), .X(n35404) );
  nand_x1_sg U68371 ( .A(n49909), .B(n57534), .X(n35401) );
  nand_x1_sg U68372 ( .A(n55913), .B(n57809), .X(n35402) );
  nand_x1_sg U68373 ( .A(n49911), .B(n57554), .X(n35409) );
  nand_x1_sg U68374 ( .A(n55911), .B(n57809), .X(n35410) );
  nand_x1_sg U68375 ( .A(n49517), .B(n57537), .X(n35407) );
  nand_x1_sg U68376 ( .A(n55909), .B(n57809), .X(n35408) );
  nand_x1_sg U68377 ( .A(n49519), .B(n57534), .X(n35391) );
  nand_x1_sg U68378 ( .A(n55907), .B(n57810), .X(n35392) );
  nand_x1_sg U68379 ( .A(n49521), .B(n57550), .X(n35389) );
  nand_x1_sg U68380 ( .A(n55905), .B(n57810), .X(n35390) );
  nand_x1_sg U68381 ( .A(n49523), .B(n57535), .X(n35397) );
  nand_x1_sg U68382 ( .A(n55903), .B(n57810), .X(n35398) );
  nand_x1_sg U68383 ( .A(n49525), .B(n57536), .X(n35395) );
  nand_x1_sg U68384 ( .A(n55901), .B(n57810), .X(n35396) );
  nand_x1_sg U68385 ( .A(n49527), .B(n57551), .X(n35427) );
  nand_x1_sg U68386 ( .A(n55899), .B(n57808), .X(n35428) );
  nand_x1_sg U68387 ( .A(n49529), .B(n57534), .X(n35425) );
  nand_x1_sg U68388 ( .A(n55897), .B(n57808), .X(n35426) );
  nand_x1_sg U68389 ( .A(n49531), .B(n57535), .X(n35433) );
  nand_x1_sg U68390 ( .A(n55895), .B(n57807), .X(n35434) );
  nand_x1_sg U68391 ( .A(n49533), .B(n57550), .X(n35431) );
  nand_x1_sg U68392 ( .A(n55893), .B(n57808), .X(n35432) );
  nand_x1_sg U68393 ( .A(n49535), .B(n57538), .X(n35415) );
  nand_x1_sg U68394 ( .A(n55891), .B(n57809), .X(n35416) );
  nand_x1_sg U68395 ( .A(n49537), .B(n57534), .X(n35413) );
  nand_x1_sg U68396 ( .A(n55889), .B(n57809), .X(n35414) );
  nand_x1_sg U68397 ( .A(n49539), .B(n57533), .X(n35421) );
  nand_x1_sg U68398 ( .A(n55887), .B(n57808), .X(n35422) );
  nand_x1_sg U68399 ( .A(n49541), .B(n57554), .X(n35419) );
  nand_x1_sg U68400 ( .A(n55885), .B(n57808), .X(n35420) );
  nand_x1_sg U68401 ( .A(n49543), .B(n57538), .X(n35357) );
  nand_x1_sg U68402 ( .A(n55883), .B(n57812), .X(n35358) );
  nand_x1_sg U68403 ( .A(n49545), .B(n57535), .X(n35355) );
  nand_x1_sg U68404 ( .A(n55881), .B(n57812), .X(n35356) );
  nand_x1_sg U68405 ( .A(n49547), .B(n57536), .X(n35363) );
  nand_x1_sg U68406 ( .A(n55879), .B(n57812), .X(n35364) );
  nand_x1_sg U68407 ( .A(n49549), .B(n57537), .X(n35361) );
  nand_x1_sg U68408 ( .A(n55877), .B(n57812), .X(n35362) );
  nand_x1_sg U68409 ( .A(n49551), .B(n57550), .X(n35345) );
  nand_x1_sg U68410 ( .A(n55875), .B(n57813), .X(n35346) );
  nand_x1_sg U68411 ( .A(n49553), .B(n57554), .X(n35343) );
  nand_x1_sg U68412 ( .A(n55873), .B(n57813), .X(n35344) );
  nand_x1_sg U68413 ( .A(n49555), .B(n57538), .X(n35351) );
  nand_x1_sg U68414 ( .A(n55871), .B(n57813), .X(n35352) );
  nand_x1_sg U68415 ( .A(n49557), .B(n57534), .X(n35349) );
  nand_x1_sg U68416 ( .A(n55869), .B(n57813), .X(n35350) );
  nand_x1_sg U68417 ( .A(n49559), .B(n57533), .X(n35379) );
  nand_x1_sg U68418 ( .A(n55867), .B(n57811), .X(n35380) );
  nand_x1_sg U68419 ( .A(n49561), .B(n57551), .X(n35377) );
  nand_x1_sg U68420 ( .A(n55865), .B(n57811), .X(n35378) );
  nand_x1_sg U68421 ( .A(n49563), .B(n57551), .X(n35385) );
  nand_x1_sg U68422 ( .A(n55863), .B(n57810), .X(n35386) );
  nand_x1_sg U68423 ( .A(n49565), .B(n57533), .X(n35383) );
  nand_x1_sg U68424 ( .A(n55861), .B(n57811), .X(n35384) );
  nand_x1_sg U68425 ( .A(n49567), .B(n57534), .X(n35369) );
  nand_x1_sg U68426 ( .A(n55859), .B(n57811), .X(n35370) );
  nand_x1_sg U68427 ( .A(n49569), .B(n57554), .X(n35367) );
  nand_x1_sg U68428 ( .A(n55857), .B(n57812), .X(n35368) );
  nand_x1_sg U68429 ( .A(n49571), .B(n57550), .X(n35375) );
  nand_x1_sg U68430 ( .A(n55855), .B(n57811), .X(n35376) );
  nand_x1_sg U68431 ( .A(n49573), .B(n57550), .X(n35373) );
  nand_x1_sg U68432 ( .A(n55853), .B(n57811), .X(n35374) );
  nand_x1_sg U68433 ( .A(n49575), .B(n57553), .X(n35461) );
  nand_x1_sg U68434 ( .A(n55851), .B(n57806), .X(n35462) );
  nand_x1_sg U68435 ( .A(n49577), .B(n57534), .X(n35459) );
  nand_x1_sg U68436 ( .A(n55849), .B(n57806), .X(n35460) );
  nand_x1_sg U68437 ( .A(n49579), .B(n57537), .X(n35439) );
  nand_x1_sg U68438 ( .A(n55847), .B(n57807), .X(n35440) );
  nand_x1_sg U68439 ( .A(n49581), .B(n57534), .X(n35467) );
  nand_x1_sg U68440 ( .A(n55845), .B(n57805), .X(n35468) );
  nand_x1_sg U68441 ( .A(n49583), .B(n57533), .X(n35465) );
  nand_x1_sg U68442 ( .A(n55843), .B(n57805), .X(n35466) );
  nand_x1_sg U68443 ( .A(n49585), .B(n57534), .X(n35463) );
  nand_x1_sg U68444 ( .A(n55841), .B(n57806), .X(n35464) );
  nand_x1_sg U68445 ( .A(n49587), .B(n57535), .X(n35471) );
  nand_x1_sg U68446 ( .A(n55839), .B(n57805), .X(n35472) );
  nand_x1_sg U68447 ( .A(n49589), .B(n57536), .X(n35469) );
  nand_x1_sg U68448 ( .A(n55837), .B(n57805), .X(n35470) );
  nand_x1_sg U68449 ( .A(n49591), .B(n57550), .X(n35493) );
  nand_x1_sg U68450 ( .A(n55835), .B(n57839), .X(n35494) );
  nand_x1_sg U68451 ( .A(n49593), .B(n57550), .X(n35491) );
  nand_x1_sg U68452 ( .A(n55833), .B(n57795), .X(n35492) );
  nand_x1_sg U68453 ( .A(n49595), .B(n57537), .X(n35473) );
  nand_x1_sg U68454 ( .A(n55831), .B(n57805), .X(n35474) );
  nand_x1_sg U68455 ( .A(n49597), .B(n57554), .X(n35489) );
  nand_x1_sg U68456 ( .A(n55829), .B(n57839), .X(n35490) );
  nand_x1_sg U68457 ( .A(n49599), .B(n57558), .X(n35477) );
  nand_x1_sg U68458 ( .A(n55827), .B(n57805), .X(n35478) );
  nand_x1_sg U68459 ( .A(n49601), .B(n57538), .X(n35475) );
  nand_x1_sg U68460 ( .A(n55825), .B(n57805), .X(n35476) );
  nand_x1_sg U68461 ( .A(n49603), .B(n57550), .X(n35481) );
  nand_x1_sg U68462 ( .A(n55823), .B(n57795), .X(n35482) );
  nand_x1_sg U68463 ( .A(n49605), .B(n57533), .X(n35479) );
  nand_x1_sg U68464 ( .A(n55821), .B(n57805), .X(n35480) );
  nand_x1_sg U68465 ( .A(n49607), .B(n57550), .X(n35429) );
  nand_x1_sg U68466 ( .A(n55819), .B(n57808), .X(n35430) );
  nand_x1_sg U68467 ( .A(n49609), .B(n57551), .X(n35437) );
  nand_x1_sg U68468 ( .A(n55817), .B(n57807), .X(n35438) );
  nand_x1_sg U68469 ( .A(n49611), .B(n57533), .X(n35445) );
  nand_x1_sg U68470 ( .A(n55815), .B(n57807), .X(n35446) );
  nand_x1_sg U68471 ( .A(n49613), .B(n57533), .X(n35443) );
  nand_x1_sg U68472 ( .A(n55813), .B(n57807), .X(n35444) );
  nand_x1_sg U68473 ( .A(n49615), .B(n57533), .X(n35423) );
  nand_x1_sg U68474 ( .A(n55811), .B(n57808), .X(n35424) );
  nand_x1_sg U68475 ( .A(n49623), .B(n57551), .X(n35435) );
  nand_x1_sg U68476 ( .A(n55803), .B(n57807), .X(n35436) );
  nand_x1_sg U68477 ( .A(n49625), .B(n57558), .X(n35453) );
  nand_x1_sg U68478 ( .A(n55801), .B(n57806), .X(n35454) );
  nand_x1_sg U68479 ( .A(n49627), .B(n57534), .X(n35457) );
  nand_x1_sg U68480 ( .A(n55799), .B(n57806), .X(n35458) );
  nand_x1_sg U68481 ( .A(n49629), .B(n57554), .X(n35455) );
  nand_x1_sg U68482 ( .A(n55797), .B(n57806), .X(n35456) );
  nand_x1_sg U68483 ( .A(n49631), .B(n57534), .X(n35451) );
  nand_x1_sg U68484 ( .A(n55795), .B(n57806), .X(n35452) );
  nand_x1_sg U68485 ( .A(n49633), .B(n57551), .X(n35449) );
  nand_x1_sg U68486 ( .A(n55793), .B(n57806), .X(n35450) );
  nand_x1_sg U68487 ( .A(n49635), .B(n57537), .X(n35441) );
  nand_x1_sg U68488 ( .A(n55791), .B(n57807), .X(n35442) );
  nand_x1_sg U68489 ( .A(n49637), .B(n57538), .X(n35447) );
  nand_x1_sg U68490 ( .A(n55789), .B(n57807), .X(n35448) );
  nand_x1_sg U68491 ( .A(n49639), .B(n57558), .X(n35231) );
  nand_x1_sg U68492 ( .A(n55787), .B(n57820), .X(n35232) );
  nand_x1_sg U68493 ( .A(n49645), .B(n57554), .X(n35235) );
  nand_x1_sg U68494 ( .A(n55781), .B(n57820), .X(n35236) );
  nand_x1_sg U68495 ( .A(n49647), .B(n57554), .X(n35223) );
  nand_x1_sg U68496 ( .A(n55779), .B(n57808), .X(n35224) );
  nand_x1_sg U68497 ( .A(n49649), .B(n57552), .X(n35221) );
  nand_x1_sg U68498 ( .A(n55777), .B(n57814), .X(n35222) );
  nand_x1_sg U68499 ( .A(n49651), .B(n57558), .X(n35227) );
  nand_x1_sg U68500 ( .A(n55775), .B(n57820), .X(n35228) );
  nand_x1_sg U68501 ( .A(n49655), .B(n57534), .X(n35249) );
  nand_x1_sg U68502 ( .A(n55771), .B(n57819), .X(n35250) );
  nand_x1_sg U68503 ( .A(n49659), .B(n57534), .X(n35255) );
  nand_x1_sg U68504 ( .A(n55767), .B(n57819), .X(n35256) );
  nand_x1_sg U68505 ( .A(n49661), .B(n57551), .X(n35253) );
  nand_x1_sg U68506 ( .A(n55765), .B(n57819), .X(n35254) );
  nand_x1_sg U68507 ( .A(n49663), .B(n57534), .X(n35239) );
  nand_x1_sg U68508 ( .A(n55763), .B(n57820), .X(n35240) );
  nand_x1_sg U68509 ( .A(n49667), .B(n57557), .X(n35245) );
  nand_x1_sg U68510 ( .A(n55759), .B(n57819), .X(n35246) );
  nand_x1_sg U68511 ( .A(n49669), .B(n57557), .X(n35243) );
  nand_x1_sg U68512 ( .A(n55757), .B(n57819), .X(n35244) );
  nand_x1_sg U68513 ( .A(n49671), .B(n57551), .X(n35189) );
  nand_x1_sg U68514 ( .A(n55755), .B(n57824), .X(n35190) );
  nand_x1_sg U68515 ( .A(n49675), .B(n57558), .X(n35195) );
  nand_x1_sg U68516 ( .A(n55751), .B(n57837), .X(n35196) );
  nand_x1_sg U68517 ( .A(n49677), .B(n57533), .X(n35193) );
  nand_x1_sg U68518 ( .A(n55749), .B(n57838), .X(n35194) );
  nand_x1_sg U68519 ( .A(n49679), .B(n57550), .X(n35179) );
  nand_x1_sg U68520 ( .A(n55747), .B(n57850), .X(n35180) );
  nand_x1_sg U68521 ( .A(n49681), .B(n57557), .X(n35177) );
  nand_x1_sg U68522 ( .A(n55745), .B(n57844), .X(n35178) );
  nand_x1_sg U68523 ( .A(n49683), .B(n57552), .X(n35185) );
  nand_x1_sg U68524 ( .A(n55743), .B(n57850), .X(n35186) );
  nand_x1_sg U68525 ( .A(n49685), .B(n57551), .X(n35183) );
  nand_x1_sg U68526 ( .A(n55741), .B(n57845), .X(n35184) );
  nand_x1_sg U68527 ( .A(n49689), .B(n57552), .X(n35211) );
  nand_x1_sg U68528 ( .A(n55737), .B(n57815), .X(n35212) );
  nand_x1_sg U68529 ( .A(n49691), .B(n57558), .X(n35217) );
  nand_x1_sg U68530 ( .A(n55735), .B(n57816), .X(n35218) );
  nand_x1_sg U68531 ( .A(n49693), .B(n57534), .X(n35215) );
  nand_x1_sg U68532 ( .A(n55733), .B(n57817), .X(n35216) );
  nand_x1_sg U68533 ( .A(n49695), .B(n57534), .X(n35201) );
  nand_x1_sg U68534 ( .A(n55731), .B(n57826), .X(n35202) );
  nand_x1_sg U68535 ( .A(n49697), .B(n57551), .X(n35199) );
  nand_x1_sg U68536 ( .A(n55729), .B(n57846), .X(n35200) );
  nand_x1_sg U68537 ( .A(n49699), .B(n57550), .X(n35207) );
  nand_x1_sg U68538 ( .A(n55727), .B(n57845), .X(n35208) );
  nand_x1_sg U68539 ( .A(n49701), .B(n57533), .X(n35205) );
  nand_x1_sg U68540 ( .A(n55725), .B(n57845), .X(n35206) );
  nand_x1_sg U68541 ( .A(n49703), .B(n57559), .X(n35315) );
  nand_x1_sg U68542 ( .A(n55723), .B(n57815), .X(n35316) );
  nand_x1_sg U68543 ( .A(n49705), .B(n57554), .X(n35313) );
  nand_x1_sg U68544 ( .A(n55721), .B(n57815), .X(n35314) );
  nand_x1_sg U68545 ( .A(n49707), .B(n57554), .X(n35321) );
  nand_x1_sg U68546 ( .A(n55719), .B(n57814), .X(n35322) );
  nand_x1_sg U68547 ( .A(n49709), .B(n57533), .X(n35319) );
  nand_x1_sg U68548 ( .A(n55717), .B(n57815), .X(n35320) );
  nand_x1_sg U68549 ( .A(n49711), .B(n57554), .X(n35305) );
  nand_x1_sg U68550 ( .A(n55715), .B(n57815), .X(n35306) );
  nand_x1_sg U68551 ( .A(n49713), .B(n57558), .X(n35303) );
  nand_x1_sg U68552 ( .A(n55713), .B(n57816), .X(n35304) );
  nand_x1_sg U68553 ( .A(n49319), .B(n57557), .X(n35309) );
  nand_x1_sg U68554 ( .A(n55711), .B(n57815), .X(n35310) );
  nand_x1_sg U68555 ( .A(n49323), .B(n57554), .X(n35335) );
  nand_x1_sg U68556 ( .A(n55707), .B(n57814), .X(n35336) );
  nand_x1_sg U68557 ( .A(n49327), .B(n57551), .X(n35339) );
  nand_x1_sg U68558 ( .A(n55703), .B(n57813), .X(n35340) );
  nand_x1_sg U68559 ( .A(n49331), .B(n57534), .X(n35325) );
  nand_x1_sg U68560 ( .A(n55699), .B(n57814), .X(n35326) );
  nand_x1_sg U68561 ( .A(n49335), .B(n57554), .X(n35331) );
  nand_x1_sg U68562 ( .A(n55695), .B(n57814), .X(n35332) );
  nand_x1_sg U68563 ( .A(n49337), .B(n57558), .X(n35329) );
  nand_x1_sg U68564 ( .A(n55693), .B(n57814), .X(n35330) );
  nand_x1_sg U68565 ( .A(n49339), .B(n57534), .X(n35273) );
  nand_x1_sg U68566 ( .A(n55691), .B(n57817), .X(n35274) );
  nand_x1_sg U68567 ( .A(n49341), .B(n57551), .X(n35271) );
  nand_x1_sg U68568 ( .A(n55689), .B(n57818), .X(n35272) );
  nand_x1_sg U68569 ( .A(n49343), .B(n57550), .X(n35279) );
  nand_x1_sg U68570 ( .A(n55687), .B(n57817), .X(n35280) );
  nand_x1_sg U68571 ( .A(n49345), .B(n57551), .X(n35277) );
  nand_x1_sg U68572 ( .A(n55685), .B(n57817), .X(n35278) );
  nand_x1_sg U68573 ( .A(n49347), .B(n57535), .X(n35261) );
  nand_x1_sg U68574 ( .A(n55683), .B(n57818), .X(n35262) );
  nand_x1_sg U68575 ( .A(n49349), .B(n57558), .X(n35259) );
  nand_x1_sg U68576 ( .A(n55681), .B(n57818), .X(n35260) );
  nand_x1_sg U68577 ( .A(n49351), .B(n57557), .X(n35267) );
  nand_x1_sg U68578 ( .A(n55679), .B(n57818), .X(n35268) );
  nand_x1_sg U68579 ( .A(n49353), .B(n57554), .X(n35265) );
  nand_x1_sg U68580 ( .A(n55677), .B(n57818), .X(n35266) );
  nand_x1_sg U68581 ( .A(n49355), .B(n57553), .X(n35293) );
  nand_x1_sg U68582 ( .A(n55675), .B(n57816), .X(n35294) );
  nand_x1_sg U68583 ( .A(n49357), .B(n57537), .X(n35291) );
  nand_x1_sg U68584 ( .A(n55673), .B(n57816), .X(n35292) );
  nand_x1_sg U68585 ( .A(n49359), .B(n57536), .X(n35299) );
  nand_x1_sg U68586 ( .A(n55671), .B(n57816), .X(n35300) );
  nand_x1_sg U68587 ( .A(n49361), .B(n57538), .X(n35297) );
  nand_x1_sg U68588 ( .A(n55669), .B(n57816), .X(n35298) );
  nand_x1_sg U68589 ( .A(n49367), .B(n57551), .X(n35287) );
  nand_x1_sg U68590 ( .A(n55663), .B(n57817), .X(n35288) );
  nand_x1_sg U68591 ( .A(n49369), .B(n57550), .X(n35285) );
  nand_x1_sg U68592 ( .A(n55661), .B(n57817), .X(n35286) );
  nand_x1_sg U68593 ( .A(n49371), .B(n57545), .X(n34707) );
  nand_x1_sg U68594 ( .A(n55659), .B(n57846), .X(n34708) );
  nand_x1_sg U68595 ( .A(n49373), .B(n57552), .X(n34701) );
  nand_x1_sg U68596 ( .A(n55657), .B(n57824), .X(n34702) );
  nand_x1_sg U68597 ( .A(n49377), .B(n57545), .X(n34713) );
  nand_x1_sg U68598 ( .A(n55653), .B(n57821), .X(n34714) );
  nand_x1_sg U68599 ( .A(n49379), .B(n57544), .X(n34725) );
  nand_x1_sg U68600 ( .A(n55651), .B(n57825), .X(n34726) );
  nand_x1_sg U68601 ( .A(n49381), .B(n57545), .X(n34719) );
  nand_x1_sg U68602 ( .A(n55649), .B(n57825), .X(n34720) );
  nand_x1_sg U68603 ( .A(n49435), .B(n57554), .X(n35509) );
  nand_x1_sg U68604 ( .A(n55595), .B(n57804), .X(n35510) );
  nand_x1_sg U68605 ( .A(n49437), .B(n57540), .X(n34887) );
  nand_x1_sg U68606 ( .A(n55593), .B(n57821), .X(n34888) );
  nand_x1_sg U68607 ( .A(n49439), .B(n57551), .X(n34869) );
  nand_x1_sg U68608 ( .A(n55591), .B(n57839), .X(n34870) );
  nand_x1_sg U68609 ( .A(n49441), .B(n57551), .X(n35405) );
  nand_x1_sg U68610 ( .A(n55589), .B(n57809), .X(n35406) );
  nand_x1_sg U68611 ( .A(n49443), .B(n57550), .X(n35341) );
  nand_x1_sg U68612 ( .A(n55587), .B(n57813), .X(n35342) );
  nand_x1_sg U68613 ( .A(n49445), .B(n57534), .X(n35507) );
  nand_x1_sg U68614 ( .A(n55585), .B(n57804), .X(n35508) );
  nand_x1_sg U68615 ( .A(n49451), .B(n57550), .X(n35181) );
  nand_x1_sg U68616 ( .A(n55579), .B(n46204), .X(n35182) );
  nand_x1_sg U68617 ( .A(n49455), .B(n57533), .X(n35307) );
  nand_x1_sg U68618 ( .A(n55575), .B(n57815), .X(n35308) );
  nand_x1_sg U68619 ( .A(n49457), .B(n57533), .X(n35097) );
  nand_x1_sg U68620 ( .A(n55573), .B(n57824), .X(n35098) );
  nand_x1_sg U68621 ( .A(n49459), .B(n57533), .X(n35301) );
  nand_x1_sg U68622 ( .A(n55571), .B(n57816), .X(n35302) );
  nand_x1_sg U68623 ( .A(n49461), .B(n57533), .X(n35289) );
  nand_x1_sg U68624 ( .A(n55569), .B(n57816), .X(n35290) );
  nand_x1_sg U68625 ( .A(n49463), .B(n57558), .X(n35327) );
  nand_x1_sg U68626 ( .A(n55567), .B(n57814), .X(n35328) );
  nand_x1_sg U68627 ( .A(n49465), .B(n57554), .X(n35347) );
  nand_x1_sg U68628 ( .A(n55565), .B(n57813), .X(n35348) );
  nand_x1_sg U68629 ( .A(n49495), .B(n57550), .X(n35003) );
  nand_x1_sg U68630 ( .A(n55535), .B(n46204), .X(n35004) );
  nand_x1_sg U68631 ( .A(n49499), .B(n57551), .X(n35169) );
  nand_x1_sg U68632 ( .A(n55531), .B(n57826), .X(n35170) );
  nand_x1_sg U68633 ( .A(n49501), .B(n57553), .X(n35091) );
  nand_x1_sg U68634 ( .A(n55529), .B(n57812), .X(n35092) );
  nand_x1_sg U68635 ( .A(n49503), .B(n57552), .X(n35055) );
  nand_x1_sg U68636 ( .A(n55527), .B(n57843), .X(n35056) );
  nand_x1_sg U68637 ( .A(n49505), .B(n57551), .X(n35079) );
  nand_x1_sg U68638 ( .A(n55525), .B(n57822), .X(n35080) );
  nand_x1_sg U68639 ( .A(n49507), .B(n57535), .X(n35191) );
  nand_x1_sg U68640 ( .A(n55523), .B(n57845), .X(n35192) );
  nand_x1_sg U68641 ( .A(n49513), .B(n57536), .X(n35187) );
  nand_x1_sg U68642 ( .A(n55517), .B(n57846), .X(n35188) );
  nand_x1_sg U68643 ( .A(n49125), .B(n57536), .X(n35251) );
  nand_x1_sg U68644 ( .A(n55509), .B(n57819), .X(n35252) );
  nand_x1_sg U68645 ( .A(n49129), .B(n57558), .X(n35501) );
  nand_x1_sg U68646 ( .A(n55505), .B(n57804), .X(n35502) );
  nand_x1_sg U68647 ( .A(n49133), .B(n57536), .X(n34965) );
  nand_x1_sg U68648 ( .A(n55501), .B(n57844), .X(n34966) );
  nand_x1_sg U68649 ( .A(n49135), .B(n57543), .X(n34755) );
  nand_x1_sg U68650 ( .A(n55499), .B(n57844), .X(n34756) );
  nand_x1_sg U68651 ( .A(n49137), .B(n57543), .X(n34749) );
  nand_x1_sg U68652 ( .A(n55497), .B(n57825), .X(n34750) );
  nand_x1_sg U68653 ( .A(n49139), .B(n57543), .X(n34743) );
  nand_x1_sg U68654 ( .A(n55495), .B(n57825), .X(n34744) );
  nand_x1_sg U68655 ( .A(n49141), .B(n57544), .X(n34737) );
  nand_x1_sg U68656 ( .A(n55493), .B(n57825), .X(n34738) );
  nand_x1_sg U68657 ( .A(n49143), .B(n57541), .X(n34779) );
  nand_x1_sg U68658 ( .A(n55491), .B(n57824), .X(n34780) );
  nand_x1_sg U68659 ( .A(n49145), .B(n57541), .X(n34791) );
  nand_x1_sg U68660 ( .A(n55489), .B(n57824), .X(n34792) );
  nand_x1_sg U68661 ( .A(n49147), .B(n57542), .X(n34773) );
  nand_x1_sg U68662 ( .A(n55487), .B(n57844), .X(n34774) );
  nand_x1_sg U68663 ( .A(n49149), .B(n57542), .X(n34767) );
  nand_x1_sg U68664 ( .A(n55485), .B(n57845), .X(n34768) );
  nand_x1_sg U68665 ( .A(n49151), .B(n57541), .X(n34845) );
  nand_x1_sg U68666 ( .A(n55483), .B(n57822), .X(n34846) );
  nand_x1_sg U68667 ( .A(n49153), .B(n57557), .X(n35241) );
  nand_x1_sg U68668 ( .A(n55481), .B(n57819), .X(n35242) );
  nand_x1_sg U68669 ( .A(n49155), .B(n57541), .X(n34833) );
  nand_x1_sg U68670 ( .A(n55479), .B(n57823), .X(n34834) );
  nand_x1_sg U68671 ( .A(n49157), .B(n57552), .X(n34851) );
  nand_x1_sg U68672 ( .A(n55477), .B(n57822), .X(n34852) );
  nand_x1_sg U68673 ( .A(n49159), .B(n57536), .X(n34959) );
  nand_x1_sg U68674 ( .A(n55475), .B(n46204), .X(n34960) );
  nand_x1_sg U68675 ( .A(n49161), .B(n57540), .X(n34893) );
  nand_x1_sg U68676 ( .A(n55473), .B(n57823), .X(n34894) );
  nand_x1_sg U68677 ( .A(n49163), .B(n57538), .X(n34923) );
  nand_x1_sg U68678 ( .A(n55471), .B(n57846), .X(n34924) );
  nand_x1_sg U68679 ( .A(n49165), .B(n57537), .X(n34947) );
  nand_x1_sg U68680 ( .A(n55469), .B(n57822), .X(n34948) );
  nand_x1_sg U68681 ( .A(n49173), .B(n57550), .X(n35483) );
  nand_x1_sg U68682 ( .A(n55461), .B(n57839), .X(n35484) );
  nand_x1_sg U68683 ( .A(n49199), .B(n57550), .X(n35411) );
  nand_x1_sg U68684 ( .A(n55435), .B(n57809), .X(n35412) );
  nand_x1_sg U68685 ( .A(n49215), .B(n57534), .X(n35495) );
  nand_x1_sg U68686 ( .A(n55419), .B(n57795), .X(n35496) );
  nand_x1_sg U68687 ( .A(n49231), .B(n57542), .X(n34765) );
  nand_x1_sg U68688 ( .A(n55403), .B(n57846), .X(n34766) );
  nand_x1_sg U68689 ( .A(n49233), .B(n57542), .X(n34763) );
  nand_x1_sg U68690 ( .A(n55401), .B(n57824), .X(n34764) );
  nand_x1_sg U68691 ( .A(n49235), .B(n57542), .X(n34771) );
  nand_x1_sg U68692 ( .A(n55399), .B(n57844), .X(n34772) );
  nand_x1_sg U68693 ( .A(n49237), .B(n57542), .X(n34769) );
  nand_x1_sg U68694 ( .A(n55397), .B(n57845), .X(n34770) );
  nand_x1_sg U68695 ( .A(n49239), .B(n57543), .X(n34753) );
  nand_x1_sg U68696 ( .A(n55395), .B(n57844), .X(n34754) );
  nand_x1_sg U68697 ( .A(n49241), .B(n57543), .X(n34751) );
  nand_x1_sg U68698 ( .A(n55393), .B(n57825), .X(n34752) );
  nand_x1_sg U68699 ( .A(n49243), .B(n57543), .X(n34759) );
  nand_x1_sg U68700 ( .A(n55391), .B(n57844), .X(n34760) );
  nand_x1_sg U68701 ( .A(n49245), .B(n57543), .X(n34757) );
  nand_x1_sg U68702 ( .A(n55389), .B(n57825), .X(n34758) );
  nand_x1_sg U68703 ( .A(n49247), .B(n57541), .X(n34789) );
  nand_x1_sg U68704 ( .A(n55387), .B(n57824), .X(n34790) );
  nand_x1_sg U68705 ( .A(n49249), .B(n57541), .X(n34787) );
  nand_x1_sg U68706 ( .A(n55385), .B(n57824), .X(n34788) );
  nand_x1_sg U68707 ( .A(n49251), .B(n57541), .X(n34795) );
  nand_x1_sg U68708 ( .A(n55383), .B(n57824), .X(n34796) );
  nand_x1_sg U68709 ( .A(n49253), .B(n57541), .X(n34793) );
  nand_x1_sg U68710 ( .A(n55381), .B(n57823), .X(n34794) );
  nand_x1_sg U68711 ( .A(n49255), .B(n57542), .X(n34777) );
  nand_x1_sg U68712 ( .A(n55379), .B(n57824), .X(n34778) );
  nand_x1_sg U68713 ( .A(n49257), .B(n57542), .X(n34775) );
  nand_x1_sg U68714 ( .A(n55377), .B(n57846), .X(n34776) );
  nand_x1_sg U68715 ( .A(n49259), .B(n57541), .X(n34783) );
  nand_x1_sg U68716 ( .A(n55375), .B(n57824), .X(n34784) );
  nand_x1_sg U68717 ( .A(n49261), .B(n57541), .X(n34781) );
  nand_x1_sg U68718 ( .A(n55373), .B(n57824), .X(n34782) );
  nand_x1_sg U68719 ( .A(n49263), .B(n57545), .X(n34717) );
  nand_x1_sg U68720 ( .A(n55371), .B(n57825), .X(n34718) );
  nand_x1_sg U68721 ( .A(n49265), .B(n57545), .X(n34715) );
  nand_x1_sg U68722 ( .A(n55369), .B(n57846), .X(n34716) );
  nand_x1_sg U68723 ( .A(n49267), .B(n57545), .X(n34723) );
  nand_x1_sg U68724 ( .A(n55367), .B(n57825), .X(n34724) );
  nand_x1_sg U68725 ( .A(n49269), .B(n57545), .X(n34721) );
  nand_x1_sg U68726 ( .A(n55365), .B(n57824), .X(n34722) );
  nand_x1_sg U68727 ( .A(n49271), .B(n57553), .X(n34705) );
  nand_x1_sg U68728 ( .A(n55363), .B(n57846), .X(n34706) );
  nand_x1_sg U68729 ( .A(n49273), .B(n57554), .X(n34703) );
  nand_x1_sg U68730 ( .A(n55361), .B(n57823), .X(n34704) );
  nand_x1_sg U68731 ( .A(n49275), .B(n57545), .X(n34711) );
  nand_x1_sg U68732 ( .A(n55359), .B(n57822), .X(n34712) );
  nand_x1_sg U68733 ( .A(n49277), .B(n57545), .X(n34709) );
  nand_x1_sg U68734 ( .A(n55357), .B(n57821), .X(n34710) );
  nand_x1_sg U68735 ( .A(n49279), .B(n57544), .X(n34741) );
  nand_x1_sg U68736 ( .A(n55355), .B(n57825), .X(n34742) );
  nand_x1_sg U68737 ( .A(n49281), .B(n57544), .X(n34739) );
  nand_x1_sg U68738 ( .A(n55353), .B(n57825), .X(n34740) );
  nand_x1_sg U68739 ( .A(n49283), .B(n57543), .X(n34747) );
  nand_x1_sg U68740 ( .A(n55351), .B(n57844), .X(n34748) );
  nand_x1_sg U68741 ( .A(n49285), .B(n57543), .X(n34745) );
  nand_x1_sg U68742 ( .A(n55349), .B(n57825), .X(n34746) );
  nand_x1_sg U68743 ( .A(n49287), .B(n57544), .X(n34729) );
  nand_x1_sg U68744 ( .A(n55347), .B(n57825), .X(n34730) );
  nand_x1_sg U68745 ( .A(n49289), .B(n57544), .X(n34727) );
  nand_x1_sg U68746 ( .A(n55345), .B(n57824), .X(n34728) );
  nand_x1_sg U68747 ( .A(n49291), .B(n57544), .X(n34735) );
  nand_x1_sg U68748 ( .A(n55343), .B(n57825), .X(n34736) );
  nand_x1_sg U68749 ( .A(n49293), .B(n57544), .X(n34733) );
  nand_x1_sg U68750 ( .A(n55341), .B(n57825), .X(n34734) );
  nand_x1_sg U68751 ( .A(n49299), .B(n57552), .X(n34797) );
  nand_x1_sg U68752 ( .A(n55335), .B(n57821), .X(n34798) );
  nand_x1_sg U68753 ( .A(n49303), .B(n57550), .X(n35145) );
  nand_x1_sg U68754 ( .A(n55331), .B(n57827), .X(n35146) );
  nand_x1_sg U68755 ( .A(n49311), .B(n57542), .X(n34761) );
  nand_x1_sg U68756 ( .A(n55323), .B(n57824), .X(n34762) );
  nand_x1_sg U68757 ( .A(n49313), .B(n57541), .X(n34785) );
  nand_x1_sg U68758 ( .A(n55321), .B(n57824), .X(n34786) );
  nand_x1_sg U68759 ( .A(n49315), .B(n57544), .X(n34731) );
  nand_x1_sg U68760 ( .A(n55319), .B(n57825), .X(n34732) );
  nand_x1_sg U68761 ( .A(n47337), .B(n57804), .X(n39840) );
  nand_x1_sg U68762 ( .A(n47595), .B(n57796), .X(n40180) );
  nand_x1_sg U68763 ( .A(n53633), .B(n57796), .X(n40175) );
  nand_x1_sg U68764 ( .A(n53631), .B(n57796), .X(n40170) );
  nand_x1_sg U68765 ( .A(n53629), .B(n57796), .X(n40165) );
  nand_x1_sg U68766 ( .A(n47503), .B(n57796), .X(n40160) );
  nand_x1_sg U68767 ( .A(n53627), .B(n57796), .X(n40150) );
  nand_x1_sg U68768 ( .A(n53647), .B(n57796), .X(n40145) );
  nand_x1_sg U68769 ( .A(n47347), .B(n57839), .X(n40140) );
  nand_x1_sg U68770 ( .A(n51039), .B(n57826), .X(n40135) );
  nand_x1_sg U68771 ( .A(n53625), .B(n57795), .X(n40130) );
  nand_x1_sg U68772 ( .A(n53623), .B(n57824), .X(n40125) );
  nand_x1_sg U68773 ( .A(n47405), .B(n57846), .X(n40120) );
  nand_x1_sg U68774 ( .A(n47581), .B(n57796), .X(n40115) );
  nand_x1_sg U68775 ( .A(n51037), .B(n57804), .X(n40110) );
  nand_x1_sg U68776 ( .A(n53621), .B(n57805), .X(n40105) );
  nand_x1_sg U68777 ( .A(n47593), .B(n57797), .X(n40100) );
  nand_x1_sg U68778 ( .A(n53619), .B(n57797), .X(n40095) );
  nand_x1_sg U68779 ( .A(n53617), .B(n57797), .X(n40090) );
  nand_x1_sg U68780 ( .A(n53615), .B(n57797), .X(n40085) );
  nand_x1_sg U68781 ( .A(n47501), .B(n57797), .X(n40080) );
  nand_x1_sg U68782 ( .A(n53613), .B(n57797), .X(n40070) );
  nand_x1_sg U68783 ( .A(n53645), .B(n57797), .X(n40065) );
  nand_x1_sg U68784 ( .A(n47345), .B(n57843), .X(n40060) );
  nand_x1_sg U68785 ( .A(n51035), .B(n57820), .X(n40055) );
  nand_x1_sg U68786 ( .A(n53611), .B(n57843), .X(n40050) );
  nand_x1_sg U68787 ( .A(n53609), .B(n57797), .X(n40045) );
  nand_x1_sg U68788 ( .A(n47403), .B(n57843), .X(n40040) );
  nand_x1_sg U68789 ( .A(n47579), .B(n57843), .X(n40035) );
  nand_x1_sg U68790 ( .A(n51033), .B(n57843), .X(n40030) );
  nand_x1_sg U68791 ( .A(n53607), .B(n57798), .X(n40025) );
  nand_x1_sg U68792 ( .A(n47591), .B(n57798), .X(n40020) );
  nand_x1_sg U68793 ( .A(n53605), .B(n57798), .X(n40015) );
  nand_x1_sg U68794 ( .A(n53603), .B(n57798), .X(n40010) );
  nand_x1_sg U68795 ( .A(n53601), .B(n57798), .X(n40005) );
  nand_x1_sg U68796 ( .A(n47499), .B(n57798), .X(n40000) );
  nand_x1_sg U68797 ( .A(n53599), .B(n57798), .X(n39990) );
  nand_x1_sg U68798 ( .A(n53643), .B(n57798), .X(n39985) );
  nand_x1_sg U68799 ( .A(n47343), .B(n57825), .X(n39980) );
  nand_x1_sg U68800 ( .A(n51031), .B(n57826), .X(n39975) );
  nand_x1_sg U68801 ( .A(n53597), .B(n57844), .X(n39970) );
  nand_x1_sg U68802 ( .A(n53595), .B(n57824), .X(n39965) );
  nand_x1_sg U68803 ( .A(n47401), .B(n57820), .X(n39960) );
  nand_x1_sg U68804 ( .A(n47577), .B(n57839), .X(n39955) );
  nand_x1_sg U68805 ( .A(n51029), .B(n57846), .X(n39950) );
  nand_x1_sg U68806 ( .A(n53593), .B(n57827), .X(n39945) );
  nand_x1_sg U68807 ( .A(n47589), .B(n57799), .X(n39940) );
  nand_x1_sg U68808 ( .A(n53591), .B(n57799), .X(n39935) );
  nand_x1_sg U68809 ( .A(n53589), .B(n57799), .X(n39930) );
  nand_x1_sg U68810 ( .A(n53587), .B(n57799), .X(n39925) );
  nand_x1_sg U68811 ( .A(n47497), .B(n57799), .X(n39920) );
  nand_x1_sg U68812 ( .A(n53585), .B(n57799), .X(n39910) );
  nand_x1_sg U68813 ( .A(n53641), .B(n57799), .X(n39905) );
  nand_x1_sg U68814 ( .A(n55069), .B(n57796), .X(n40155) );
  nand_x1_sg U68815 ( .A(n55067), .B(n57797), .X(n40075) );
  nand_x1_sg U68816 ( .A(n55065), .B(n57798), .X(n39995) );
  nand_x1_sg U68817 ( .A(n55063), .B(n57799), .X(n39915) );
  nand_x1_sg U68818 ( .A(n50429), .B(n57875), .X(n29346) );
  nand_x1_sg U68819 ( .A(n55057), .B(n57895), .X(n29347) );
  nand_x1_sg U68820 ( .A(o_mask[31]), .B(n57554), .X(n39903) );
  nand_x1_sg U68821 ( .A(n57800), .B(n47341), .X(n39904) );
  nand_x1_sg U68822 ( .A(o_mask[30]), .B(n57533), .X(n39901) );
  nand_x1_sg U68823 ( .A(n57800), .B(n51049), .X(n39902) );
  nand_x1_sg U68824 ( .A(o_mask[29]), .B(n57534), .X(n39899) );
  nand_x1_sg U68825 ( .A(n57800), .B(n51027), .X(n39900) );
  nand_x1_sg U68826 ( .A(o_mask[28]), .B(n57551), .X(n39897) );
  nand_x1_sg U68827 ( .A(n57800), .B(n51025), .X(n39898) );
  nand_x1_sg U68828 ( .A(o_mask[27]), .B(n57538), .X(n39895) );
  nand_x1_sg U68829 ( .A(n57800), .B(n47399), .X(n39896) );
  nand_x1_sg U68830 ( .A(o_mask[26]), .B(n57554), .X(n39893) );
  nand_x1_sg U68831 ( .A(n57800), .B(n47597), .X(n39894) );
  nand_x1_sg U68832 ( .A(o_mask[25]), .B(n57533), .X(n39891) );
  nand_x1_sg U68833 ( .A(n57800), .B(n51023), .X(n39892) );
  nand_x1_sg U68834 ( .A(o_mask[24]), .B(n57536), .X(n39889) );
  nand_x1_sg U68835 ( .A(n57800), .B(n51021), .X(n39890) );
  nand_x1_sg U68836 ( .A(o_mask[23]), .B(n57537), .X(n39887) );
  nand_x1_sg U68837 ( .A(n57801), .B(n51051), .X(n39888) );
  nand_x1_sg U68838 ( .A(o_mask[22]), .B(n57538), .X(n39885) );
  nand_x1_sg U68839 ( .A(n57801), .B(n51019), .X(n39886) );
  nand_x1_sg U68840 ( .A(o_mask[21]), .B(n57533), .X(n39883) );
  nand_x1_sg U68841 ( .A(n57801), .B(n51045), .X(n39884) );
  nand_x1_sg U68842 ( .A(o_mask[20]), .B(n57554), .X(n39881) );
  nand_x1_sg U68843 ( .A(n57801), .B(n51017), .X(n39882) );
  nand_x1_sg U68844 ( .A(o_mask[19]), .B(n57551), .X(n39879) );
  nand_x1_sg U68845 ( .A(n57801), .B(n47599), .X(n39880) );
  nand_x1_sg U68846 ( .A(o_mask[18]), .B(n57550), .X(n39877) );
  nand_x1_sg U68847 ( .A(n57801), .B(n51059), .X(n39878) );
  nand_x1_sg U68848 ( .A(o_mask[17]), .B(n57551), .X(n39875) );
  nand_x1_sg U68849 ( .A(n57801), .B(n47585), .X(n39876) );
  nand_x1_sg U68850 ( .A(o_mask[16]), .B(n57533), .X(n39873) );
  nand_x1_sg U68851 ( .A(n57801), .B(n51015), .X(n39874) );
  nand_x1_sg U68852 ( .A(o_mask[15]), .B(n57550), .X(n39871) );
  nand_x1_sg U68853 ( .A(n57802), .B(n47339), .X(n39872) );
  nand_x1_sg U68854 ( .A(o_mask[14]), .B(n57552), .X(n39869) );
  nand_x1_sg U68855 ( .A(n57802), .B(n51013), .X(n39870) );
  nand_x1_sg U68856 ( .A(o_mask[13]), .B(n57553), .X(n39867) );
  nand_x1_sg U68857 ( .A(n57802), .B(n51011), .X(n39868) );
  nand_x1_sg U68858 ( .A(o_mask[12]), .B(n57534), .X(n39865) );
  nand_x1_sg U68859 ( .A(n57802), .B(n51009), .X(n39866) );
  nand_x1_sg U68860 ( .A(o_mask[11]), .B(n57534), .X(n39863) );
  nand_x1_sg U68861 ( .A(n57802), .B(n47397), .X(n39864) );
  nand_x1_sg U68862 ( .A(o_mask[10]), .B(n57533), .X(n39861) );
  nand_x1_sg U68863 ( .A(n57802), .B(n47575), .X(n39862) );
  nand_x1_sg U68864 ( .A(o_mask[9]), .B(n57535), .X(n39859) );
  nand_x1_sg U68865 ( .A(n57802), .B(n51007), .X(n39860) );
  nand_x1_sg U68866 ( .A(o_mask[8]), .B(n57533), .X(n39857) );
  nand_x1_sg U68867 ( .A(n57802), .B(n51005), .X(n39858) );
  nand_x1_sg U68868 ( .A(o_mask[7]), .B(n57550), .X(n39855) );
  nand_x1_sg U68869 ( .A(n57803), .B(n51003), .X(n39856) );
  nand_x1_sg U68870 ( .A(o_mask[6]), .B(n57551), .X(n39853) );
  nand_x1_sg U68871 ( .A(n57803), .B(n51001), .X(n39854) );
  nand_x1_sg U68872 ( .A(o_mask[5]), .B(n57558), .X(n39851) );
  nand_x1_sg U68873 ( .A(n57803), .B(n51047), .X(n39852) );
  nand_x1_sg U68874 ( .A(o_mask[4]), .B(n57536), .X(n39849) );
  nand_x1_sg U68875 ( .A(n57803), .B(n47587), .X(n39850) );
  nand_x1_sg U68876 ( .A(o_mask[3]), .B(n57537), .X(n39847) );
  nand_x1_sg U68877 ( .A(n57803), .B(n51063), .X(n39848) );
  nand_x1_sg U68878 ( .A(o_mask[2]), .B(n57538), .X(n39845) );
  nand_x1_sg U68879 ( .A(n57803), .B(n51061), .X(n39846) );
  nand_x1_sg U68880 ( .A(o_mask[1]), .B(n57533), .X(n39843) );
  nand_x1_sg U68881 ( .A(n51069), .B(n57803), .X(n39844) );
  nand_x1_sg U68882 ( .A(o_mask[0]), .B(n57535), .X(n39841) );
  nand_x1_sg U68883 ( .A(n51067), .B(n57803), .X(n39842) );
  nand_x1_sg U68884 ( .A(n47349), .B(n57795), .X(n40221) );
  nand_x1_sg U68885 ( .A(n51043), .B(n57795), .X(n40215) );
  nand_x1_sg U68886 ( .A(n53639), .B(n57795), .X(n40210) );
  nand_x1_sg U68887 ( .A(n53637), .B(n57795), .X(n40205) );
  nand_x1_sg U68888 ( .A(n47407), .B(n57795), .X(n40200) );
  nand_x1_sg U68889 ( .A(n47583), .B(n57795), .X(n40195) );
  nand_x1_sg U68890 ( .A(n51041), .B(n57795), .X(n40190) );
  nand_x1_sg U68891 ( .A(n53635), .B(n57795), .X(n40185) );
  nand_x1_sg U68892 ( .A(n50319), .B(n57554), .X(n34391) );
  nand_x1_sg U68893 ( .A(n56585), .B(n57827), .X(n34392) );
  nand_x1_sg U68894 ( .A(n50379), .B(n57534), .X(n34337) );
  nand_x1_sg U68895 ( .A(n56525), .B(n46204), .X(n34338) );
  nand_x1_sg U68896 ( .A(n50381), .B(n57533), .X(n34355) );
  nand_x1_sg U68897 ( .A(n56523), .B(n57826), .X(n34356) );
  nand_x1_sg U68898 ( .A(n50383), .B(n57533), .X(n34353) );
  nand_x1_sg U68899 ( .A(n56521), .B(n57827), .X(n34354) );
  nand_x1_sg U68900 ( .A(n50399), .B(n57533), .X(n34357) );
  nand_x1_sg U68901 ( .A(n56505), .B(n57827), .X(n34358) );
  nand_x1_sg U68902 ( .A(n50111), .B(n57533), .X(n34335) );
  nand_x1_sg U68903 ( .A(n56503), .B(n57839), .X(n34336) );
  nand_x1_sg U68904 ( .A(n50113), .B(n57533), .X(n34349) );
  nand_x1_sg U68905 ( .A(n56501), .B(n57826), .X(n34350) );
  nand_x1_sg U68906 ( .A(n50119), .B(n57534), .X(n34575) );
  nand_x1_sg U68907 ( .A(n56495), .B(n57846), .X(n34576) );
  nand_x1_sg U68908 ( .A(n50121), .B(n57551), .X(n34393) );
  nand_x1_sg U68909 ( .A(n56493), .B(n57839), .X(n34394) );
  nand_x1_sg U68910 ( .A(n50141), .B(n57554), .X(n34379) );
  nand_x1_sg U68911 ( .A(n56473), .B(n57826), .X(n34380) );
  nand_x1_sg U68912 ( .A(n50157), .B(n57558), .X(n34367) );
  nand_x1_sg U68913 ( .A(n56457), .B(n57826), .X(n34368) );
  nand_x1_sg U68914 ( .A(n50187), .B(n57554), .X(n34579) );
  nand_x1_sg U68915 ( .A(n56427), .B(n57836), .X(n34580) );
  nand_x1_sg U68916 ( .A(n50189), .B(n57558), .X(n34577) );
  nand_x1_sg U68917 ( .A(n56425), .B(n57845), .X(n34578) );
  nand_x1_sg U68918 ( .A(n50191), .B(n57554), .X(n34585) );
  nand_x1_sg U68919 ( .A(n56423), .B(n57836), .X(n34586) );
  nand_x1_sg U68920 ( .A(n50193), .B(n57535), .X(n34583) );
  nand_x1_sg U68921 ( .A(n56421), .B(n57838), .X(n34584) );
  nand_x1_sg U68922 ( .A(n50195), .B(n57553), .X(n34567) );
  nand_x1_sg U68923 ( .A(n56419), .B(n57845), .X(n34568) );
  nand_x1_sg U68924 ( .A(n50197), .B(n57554), .X(n34565) );
  nand_x1_sg U68925 ( .A(n56417), .B(n57824), .X(n34566) );
  nand_x1_sg U68926 ( .A(n50199), .B(n57554), .X(n34573) );
  nand_x1_sg U68927 ( .A(n56415), .B(n57850), .X(n34574) );
  nand_x1_sg U68928 ( .A(n50201), .B(n57558), .X(n34571) );
  nand_x1_sg U68929 ( .A(n56413), .B(n57824), .X(n34572) );
  nand_x1_sg U68930 ( .A(n50203), .B(n57554), .X(n34603) );
  nand_x1_sg U68931 ( .A(n56411), .B(n57838), .X(n34604) );
  nand_x1_sg U68932 ( .A(n50205), .B(n57554), .X(n34601) );
  nand_x1_sg U68933 ( .A(n56409), .B(n57839), .X(n34602) );
  nand_x1_sg U68934 ( .A(n50207), .B(n57554), .X(n34609) );
  nand_x1_sg U68935 ( .A(n56407), .B(n57849), .X(n34610) );
  nand_x1_sg U68936 ( .A(n50209), .B(n57559), .X(n34607) );
  nand_x1_sg U68937 ( .A(n56405), .B(n57827), .X(n34608) );
  nand_x1_sg U68938 ( .A(n50211), .B(n57536), .X(n34591) );
  nand_x1_sg U68939 ( .A(n56403), .B(n57850), .X(n34592) );
  nand_x1_sg U68940 ( .A(n50213), .B(n57537), .X(n34589) );
  nand_x1_sg U68941 ( .A(n56401), .B(n57843), .X(n34590) );
  nand_x1_sg U68942 ( .A(n50215), .B(n57538), .X(n34597) );
  nand_x1_sg U68943 ( .A(n56399), .B(n57840), .X(n34598) );
  nand_x1_sg U68944 ( .A(n50217), .B(n57537), .X(n34595) );
  nand_x1_sg U68945 ( .A(n56397), .B(n57841), .X(n34596) );
  nand_x1_sg U68946 ( .A(n50219), .B(n57550), .X(n34531) );
  nand_x1_sg U68947 ( .A(n56395), .B(n57840), .X(n34532) );
  nand_x1_sg U68948 ( .A(n50221), .B(n57558), .X(n34529) );
  nand_x1_sg U68949 ( .A(n56393), .B(n57844), .X(n34530) );
  nand_x1_sg U68950 ( .A(n50223), .B(n57550), .X(n34537) );
  nand_x1_sg U68951 ( .A(n56391), .B(n57850), .X(n34538) );
  nand_x1_sg U68952 ( .A(n50225), .B(n57550), .X(n34535) );
  nand_x1_sg U68953 ( .A(n56389), .B(n57846), .X(n34536) );
  nand_x1_sg U68954 ( .A(n50227), .B(n57550), .X(n34519) );
  nand_x1_sg U68955 ( .A(n56387), .B(n57839), .X(n34520) );
  nand_x1_sg U68956 ( .A(n50229), .B(n57550), .X(n34517) );
  nand_x1_sg U68957 ( .A(n56385), .B(n57849), .X(n34518) );
  nand_x1_sg U68958 ( .A(n50231), .B(n57550), .X(n34525) );
  nand_x1_sg U68959 ( .A(n56383), .B(n57849), .X(n34526) );
  nand_x1_sg U68960 ( .A(n50233), .B(n57551), .X(n34523) );
  nand_x1_sg U68961 ( .A(n56381), .B(n57836), .X(n34524) );
  nand_x1_sg U68962 ( .A(n50235), .B(n57537), .X(n34555) );
  nand_x1_sg U68963 ( .A(n56379), .B(n57845), .X(n34556) );
  nand_x1_sg U68964 ( .A(n50237), .B(n57538), .X(n34553) );
  nand_x1_sg U68965 ( .A(n56377), .B(n57846), .X(n34554) );
  nand_x1_sg U68966 ( .A(n50239), .B(n57534), .X(n34561) );
  nand_x1_sg U68967 ( .A(n56375), .B(n57824), .X(n34562) );
  nand_x1_sg U68968 ( .A(n50241), .B(n57533), .X(n34559) );
  nand_x1_sg U68969 ( .A(n56373), .B(n57846), .X(n34560) );
  nand_x1_sg U68970 ( .A(n50243), .B(n57550), .X(n34543) );
  nand_x1_sg U68971 ( .A(n56371), .B(n34232), .X(n34544) );
  nand_x1_sg U68972 ( .A(n50245), .B(n57551), .X(n34541) );
  nand_x1_sg U68973 ( .A(n56369), .B(n57836), .X(n34542) );
  nand_x1_sg U68974 ( .A(n50247), .B(n57533), .X(n34549) );
  nand_x1_sg U68975 ( .A(n56367), .B(n57843), .X(n34550) );
  nand_x1_sg U68976 ( .A(n50249), .B(n57550), .X(n34547) );
  nand_x1_sg U68977 ( .A(n56365), .B(n57840), .X(n34548) );
  nand_x1_sg U68978 ( .A(n50251), .B(n57535), .X(n34671) );
  nand_x1_sg U68979 ( .A(n56363), .B(n57839), .X(n34672) );
  nand_x1_sg U68980 ( .A(n50253), .B(n57546), .X(n34669) );
  nand_x1_sg U68981 ( .A(n56361), .B(n57827), .X(n34670) );
  nand_x1_sg U68982 ( .A(n50255), .B(n57536), .X(n34677) );
  nand_x1_sg U68983 ( .A(n56359), .B(n46204), .X(n34678) );
  nand_x1_sg U68984 ( .A(n50257), .B(n57537), .X(n34675) );
  nand_x1_sg U68985 ( .A(n56357), .B(n46204), .X(n34676) );
  nand_x1_sg U68986 ( .A(n50259), .B(n57546), .X(n34659) );
  nand_x1_sg U68987 ( .A(n56355), .B(n46204), .X(n34660) );
  nand_x1_sg U68988 ( .A(n50261), .B(n57546), .X(n34657) );
  nand_x1_sg U68989 ( .A(n56353), .B(n57849), .X(n34658) );
  nand_x1_sg U68990 ( .A(n50263), .B(n57546), .X(n34665) );
  nand_x1_sg U68991 ( .A(n56351), .B(n57837), .X(n34666) );
  nand_x1_sg U68992 ( .A(n50265), .B(n57546), .X(n34663) );
  nand_x1_sg U68993 ( .A(n56349), .B(n46204), .X(n34664) );
  nand_x1_sg U68994 ( .A(n50267), .B(n57551), .X(n34693) );
  nand_x1_sg U68995 ( .A(n56347), .B(n57846), .X(n34694) );
  nand_x1_sg U68996 ( .A(n50269), .B(n57557), .X(n34691) );
  nand_x1_sg U68997 ( .A(n56345), .B(n57846), .X(n34692) );
  nand_x1_sg U68998 ( .A(n50275), .B(n57554), .X(n34683) );
  nand_x1_sg U68999 ( .A(n56339), .B(n57827), .X(n34684) );
  nand_x1_sg U69000 ( .A(n50277), .B(n57557), .X(n34681) );
  nand_x1_sg U69001 ( .A(n56337), .B(n57839), .X(n34682) );
  nand_x1_sg U69002 ( .A(n50279), .B(n57534), .X(n34689) );
  nand_x1_sg U69003 ( .A(n56335), .B(n57844), .X(n34690) );
  nand_x1_sg U69004 ( .A(n50281), .B(n57551), .X(n34687) );
  nand_x1_sg U69005 ( .A(n56333), .B(n57845), .X(n34688) );
  nand_x1_sg U69006 ( .A(n50283), .B(n57558), .X(n34625) );
  nand_x1_sg U69007 ( .A(n56331), .B(n46204), .X(n34626) );
  nand_x1_sg U69008 ( .A(n50285), .B(n57534), .X(n34623) );
  nand_x1_sg U69009 ( .A(n56329), .B(n57843), .X(n34624) );
  nand_x1_sg U69010 ( .A(n50287), .B(n57533), .X(n34631) );
  nand_x1_sg U69011 ( .A(n56327), .B(n57840), .X(n34632) );
  nand_x1_sg U69012 ( .A(n50289), .B(n57550), .X(n34629) );
  nand_x1_sg U69013 ( .A(n56325), .B(n57841), .X(n34630) );
  nand_x1_sg U69014 ( .A(n50291), .B(n57558), .X(n34613) );
  nand_x1_sg U69015 ( .A(n56323), .B(n57839), .X(n34614) );
  nand_x1_sg U69016 ( .A(n50293), .B(n57558), .X(n34611) );
  nand_x1_sg U69017 ( .A(n56321), .B(n57826), .X(n34612) );
  nand_x1_sg U69018 ( .A(n50295), .B(n57533), .X(n34619) );
  nand_x1_sg U69019 ( .A(n56319), .B(n57842), .X(n34620) );
  nand_x1_sg U69020 ( .A(n50297), .B(n57534), .X(n34617) );
  nand_x1_sg U69021 ( .A(n56317), .B(n57826), .X(n34618) );
  nand_x1_sg U69022 ( .A(n50299), .B(n57547), .X(n34649) );
  nand_x1_sg U69023 ( .A(n56315), .B(n57838), .X(n34650) );
  nand_x1_sg U69024 ( .A(n50301), .B(n57547), .X(n34647) );
  nand_x1_sg U69025 ( .A(n56313), .B(n57837), .X(n34648) );
  nand_x1_sg U69026 ( .A(n50303), .B(n57546), .X(n34655) );
  nand_x1_sg U69027 ( .A(n56311), .B(n57843), .X(n34656) );
  nand_x1_sg U69028 ( .A(n50305), .B(n57546), .X(n34653) );
  nand_x1_sg U69029 ( .A(n56309), .B(n57840), .X(n34654) );
  nand_x1_sg U69030 ( .A(n50307), .B(n57547), .X(n34637) );
  nand_x1_sg U69031 ( .A(n56307), .B(n57849), .X(n34638) );
  nand_x1_sg U69032 ( .A(n49913), .B(n57547), .X(n34635) );
  nand_x1_sg U69033 ( .A(n56305), .B(n57849), .X(n34636) );
  nand_x1_sg U69034 ( .A(n49915), .B(n57547), .X(n34643) );
  nand_x1_sg U69035 ( .A(n56303), .B(n57843), .X(n34644) );
  nand_x1_sg U69036 ( .A(n49917), .B(n57547), .X(n34641) );
  nand_x1_sg U69037 ( .A(n56301), .B(n57840), .X(n34642) );
  nand_x1_sg U69038 ( .A(n49919), .B(n57533), .X(n34303) );
  nand_x1_sg U69039 ( .A(n56299), .B(n57827), .X(n34304) );
  nand_x1_sg U69040 ( .A(n49921), .B(n57533), .X(n34301) );
  nand_x1_sg U69041 ( .A(n56297), .B(n57836), .X(n34302) );
  nand_x1_sg U69042 ( .A(n49923), .B(n57534), .X(n34309) );
  nand_x1_sg U69043 ( .A(n56295), .B(n57842), .X(n34310) );
  nand_x1_sg U69044 ( .A(n49925), .B(n57534), .X(n34307) );
  nand_x1_sg U69045 ( .A(n56293), .B(n57837), .X(n34308) );
  nand_x1_sg U69046 ( .A(n49927), .B(n57551), .X(n34291) );
  nand_x1_sg U69047 ( .A(n56291), .B(n57845), .X(n34292) );
  nand_x1_sg U69048 ( .A(n49929), .B(n57551), .X(n34289) );
  nand_x1_sg U69049 ( .A(n56289), .B(n57844), .X(n34290) );
  nand_x1_sg U69050 ( .A(n49931), .B(n57554), .X(n34297) );
  nand_x1_sg U69051 ( .A(n56287), .B(n57849), .X(n34298) );
  nand_x1_sg U69052 ( .A(n49933), .B(n57534), .X(n34295) );
  nand_x1_sg U69053 ( .A(n56285), .B(n57838), .X(n34296) );
  nand_x1_sg U69054 ( .A(n49935), .B(n57558), .X(n34333) );
  nand_x1_sg U69055 ( .A(n56283), .B(n57843), .X(n34334) );
  nand_x1_sg U69056 ( .A(n49937), .B(n57551), .X(n34331) );
  nand_x1_sg U69057 ( .A(n56281), .B(n57840), .X(n34332) );
  nand_x1_sg U69058 ( .A(n49943), .B(n57533), .X(n34387) );
  nand_x1_sg U69059 ( .A(n56275), .B(n46204), .X(n34388) );
  nand_x1_sg U69060 ( .A(n49945), .B(n57550), .X(n34385) );
  nand_x1_sg U69061 ( .A(n56273), .B(n57845), .X(n34386) );
  nand_x1_sg U69062 ( .A(n49955), .B(n57534), .X(n34401) );
  nand_x1_sg U69063 ( .A(n56263), .B(n57837), .X(n34402) );
  nand_x1_sg U69064 ( .A(n49957), .B(n57550), .X(n34399) );
  nand_x1_sg U69065 ( .A(n56261), .B(n57850), .X(n34400) );
  nand_x1_sg U69066 ( .A(n49967), .B(n57554), .X(n34375) );
  nand_x1_sg U69067 ( .A(n56251), .B(n57826), .X(n34376) );
  nand_x1_sg U69068 ( .A(n49969), .B(n57551), .X(n34373) );
  nand_x1_sg U69069 ( .A(n56249), .B(n57826), .X(n34374) );
  nand_x1_sg U69070 ( .A(n49973), .B(n57558), .X(n34397) );
  nand_x1_sg U69071 ( .A(n56245), .B(n57846), .X(n34398) );
  nand_x1_sg U69072 ( .A(n49975), .B(n57532), .X(n34411) );
  nand_x1_sg U69073 ( .A(n56243), .B(n57838), .X(n34412) );
  nand_x1_sg U69074 ( .A(n49977), .B(n57532), .X(n34409) );
  nand_x1_sg U69075 ( .A(n56241), .B(n57845), .X(n34410) );
  nand_x1_sg U69076 ( .A(n49979), .B(n57532), .X(n34417) );
  nand_x1_sg U69077 ( .A(n56239), .B(n57844), .X(n34418) );
  nand_x1_sg U69078 ( .A(n49981), .B(n57532), .X(n34415) );
  nand_x1_sg U69079 ( .A(n56237), .B(n57849), .X(n34416) );
  nand_x1_sg U69080 ( .A(n49983), .B(n57551), .X(n34483) );
  nand_x1_sg U69081 ( .A(n56235), .B(n57850), .X(n34484) );
  nand_x1_sg U69082 ( .A(n49985), .B(n57550), .X(n34481) );
  nand_x1_sg U69083 ( .A(n56233), .B(n57838), .X(n34482) );
  nand_x1_sg U69084 ( .A(n49987), .B(n57550), .X(n34489) );
  nand_x1_sg U69085 ( .A(n56231), .B(n57850), .X(n34490) );
  nand_x1_sg U69086 ( .A(n49989), .B(n57551), .X(n34487) );
  nand_x1_sg U69087 ( .A(n56229), .B(n57839), .X(n34488) );
  nand_x1_sg U69088 ( .A(n49991), .B(n57530), .X(n34471) );
  nand_x1_sg U69089 ( .A(n56227), .B(n57850), .X(n34472) );
  nand_x1_sg U69090 ( .A(n49993), .B(n57530), .X(n34469) );
  nand_x1_sg U69091 ( .A(n56225), .B(n57842), .X(n34470) );
  nand_x1_sg U69092 ( .A(n49995), .B(n57550), .X(n34477) );
  nand_x1_sg U69093 ( .A(n56223), .B(n57827), .X(n34478) );
  nand_x1_sg U69094 ( .A(n49997), .B(n57551), .X(n34475) );
  nand_x1_sg U69095 ( .A(n56221), .B(n57850), .X(n34476) );
  nand_x1_sg U69096 ( .A(n49999), .B(n57538), .X(n34507) );
  nand_x1_sg U69097 ( .A(n56219), .B(n57838), .X(n34508) );
  nand_x1_sg U69098 ( .A(n50001), .B(n57551), .X(n34505) );
  nand_x1_sg U69099 ( .A(n56217), .B(n46204), .X(n34506) );
  nand_x1_sg U69100 ( .A(n50003), .B(n57554), .X(n34513) );
  nand_x1_sg U69101 ( .A(n56215), .B(n57846), .X(n34514) );
  nand_x1_sg U69102 ( .A(n50005), .B(n57550), .X(n34511) );
  nand_x1_sg U69103 ( .A(n56213), .B(n57837), .X(n34512) );
  nand_x1_sg U69104 ( .A(n50007), .B(n57558), .X(n34495) );
  nand_x1_sg U69105 ( .A(n56211), .B(n57850), .X(n34496) );
  nand_x1_sg U69106 ( .A(n50009), .B(n57550), .X(n34493) );
  nand_x1_sg U69107 ( .A(n56209), .B(n57836), .X(n34494) );
  nand_x1_sg U69108 ( .A(n50011), .B(n57551), .X(n34501) );
  nand_x1_sg U69109 ( .A(n56207), .B(n46204), .X(n34502) );
  nand_x1_sg U69110 ( .A(n50013), .B(n57554), .X(n34499) );
  nand_x1_sg U69111 ( .A(n56205), .B(n57838), .X(n34500) );
  nand_x1_sg U69112 ( .A(n50015), .B(n57534), .X(n34435) );
  nand_x1_sg U69113 ( .A(n56203), .B(n57837), .X(n34436) );
  nand_x1_sg U69114 ( .A(n50017), .B(n57533), .X(n34433) );
  nand_x1_sg U69115 ( .A(n56201), .B(n57838), .X(n34434) );
  nand_x1_sg U69116 ( .A(n50019), .B(n57531), .X(n34441) );
  nand_x1_sg U69117 ( .A(n56199), .B(n57844), .X(n34442) );
  nand_x1_sg U69118 ( .A(n50021), .B(n57531), .X(n34439) );
  nand_x1_sg U69119 ( .A(n56197), .B(n57839), .X(n34440) );
  nand_x1_sg U69120 ( .A(n50023), .B(n57534), .X(n34423) );
  nand_x1_sg U69121 ( .A(n56195), .B(n46204), .X(n34424) );
  nand_x1_sg U69122 ( .A(n50025), .B(n57533), .X(n34421) );
  nand_x1_sg U69123 ( .A(n56193), .B(n46204), .X(n34422) );
  nand_x1_sg U69124 ( .A(n50027), .B(n57535), .X(n34429) );
  nand_x1_sg U69125 ( .A(n56191), .B(n57849), .X(n34430) );
  nand_x1_sg U69126 ( .A(n50029), .B(n57536), .X(n34427) );
  nand_x1_sg U69127 ( .A(n56189), .B(n57844), .X(n34428) );
  nand_x1_sg U69128 ( .A(n50031), .B(n57530), .X(n34459) );
  nand_x1_sg U69129 ( .A(n56187), .B(n57836), .X(n34460) );
  nand_x1_sg U69130 ( .A(n50033), .B(n57530), .X(n34457) );
  nand_x1_sg U69131 ( .A(n56185), .B(n57845), .X(n34458) );
  nand_x1_sg U69132 ( .A(n50035), .B(n57530), .X(n34465) );
  nand_x1_sg U69133 ( .A(n56183), .B(n57843), .X(n34466) );
  nand_x1_sg U69134 ( .A(n50037), .B(n57530), .X(n34463) );
  nand_x1_sg U69135 ( .A(n56181), .B(n57842), .X(n34464) );
  nand_x1_sg U69136 ( .A(n50039), .B(n57531), .X(n34447) );
  nand_x1_sg U69137 ( .A(n56179), .B(n57845), .X(n34448) );
  nand_x1_sg U69138 ( .A(n50041), .B(n57531), .X(n34445) );
  nand_x1_sg U69139 ( .A(n56177), .B(n57842), .X(n34446) );
  nand_x1_sg U69140 ( .A(n50043), .B(n57531), .X(n34453) );
  nand_x1_sg U69141 ( .A(n56175), .B(n57840), .X(n34454) );
  nand_x1_sg U69142 ( .A(n50045), .B(n57531), .X(n34451) );
  nand_x1_sg U69143 ( .A(n56173), .B(n57841), .X(n34452) );
  nand_x1_sg U69144 ( .A(n49617), .B(n57533), .X(n34363) );
  nand_x1_sg U69145 ( .A(n55809), .B(n57826), .X(n34364) );
  nand_x1_sg U69146 ( .A(n49619), .B(n57533), .X(n34361) );
  nand_x1_sg U69147 ( .A(n55807), .B(n57826), .X(n34362) );
  nand_x1_sg U69148 ( .A(n49621), .B(n57533), .X(n34359) );
  nand_x1_sg U69149 ( .A(n55805), .B(n57826), .X(n34360) );
  nand_x1_sg U69150 ( .A(n49653), .B(n57536), .X(n34259) );
  nand_x1_sg U69151 ( .A(n55773), .B(n57843), .X(n34260) );
  nand_x1_sg U69152 ( .A(n49657), .B(n57535), .X(n34255) );
  nand_x1_sg U69153 ( .A(n55769), .B(n57837), .X(n34256) );
  nand_x1_sg U69154 ( .A(n49665), .B(n57535), .X(n34257) );
  nand_x1_sg U69155 ( .A(n55761), .B(n57845), .X(n34258) );
  nand_x1_sg U69156 ( .A(n49673), .B(n57535), .X(n34251) );
  nand_x1_sg U69157 ( .A(n55753), .B(n57845), .X(n34252) );
  nand_x1_sg U69158 ( .A(n49321), .B(n57535), .X(n34249) );
  nand_x1_sg U69159 ( .A(n55709), .B(n57849), .X(n34250) );
  nand_x1_sg U69160 ( .A(n49325), .B(n57535), .X(n34253) );
  nand_x1_sg U69161 ( .A(n55705), .B(n57826), .X(n34254) );
  nand_x1_sg U69162 ( .A(n49363), .B(n57550), .X(n34269) );
  nand_x1_sg U69163 ( .A(n55667), .B(n57843), .X(n34270) );
  nand_x1_sg U69164 ( .A(n49365), .B(n57534), .X(n34267) );
  nand_x1_sg U69165 ( .A(n55665), .B(n57826), .X(n34268) );
  nand_x1_sg U69166 ( .A(n49375), .B(n57533), .X(n34271) );
  nand_x1_sg U69167 ( .A(n55655), .B(n57827), .X(n34272) );
  nand_x1_sg U69168 ( .A(n49383), .B(n57535), .X(n34581) );
  nand_x1_sg U69169 ( .A(n55647), .B(n57839), .X(n34582) );
  nand_x1_sg U69170 ( .A(n49385), .B(n57550), .X(n34605) );
  nand_x1_sg U69171 ( .A(n55645), .B(n46204), .X(n34606) );
  nand_x1_sg U69172 ( .A(n49387), .B(n57552), .X(n34569) );
  nand_x1_sg U69173 ( .A(n55643), .B(n57837), .X(n34570) );
  nand_x1_sg U69174 ( .A(n49389), .B(n57554), .X(n34563) );
  nand_x1_sg U69175 ( .A(n55641), .B(n57839), .X(n34564) );
  nand_x1_sg U69176 ( .A(n49391), .B(n57533), .X(n34557) );
  nand_x1_sg U69177 ( .A(n55639), .B(n57841), .X(n34558) );
  nand_x1_sg U69178 ( .A(n49393), .B(n57534), .X(n34551) );
  nand_x1_sg U69179 ( .A(n55637), .B(n57841), .X(n34552) );
  nand_x1_sg U69180 ( .A(n49395), .B(n57532), .X(n34599) );
  nand_x1_sg U69181 ( .A(n55635), .B(n57842), .X(n34600) );
  nand_x1_sg U69182 ( .A(n49397), .B(n57551), .X(n34615) );
  nand_x1_sg U69183 ( .A(n55633), .B(n46204), .X(n34616) );
  nand_x1_sg U69184 ( .A(n49399), .B(n57533), .X(n34593) );
  nand_x1_sg U69185 ( .A(n55631), .B(n57850), .X(n34594) );
  nand_x1_sg U69186 ( .A(n49401), .B(n57533), .X(n34587) );
  nand_x1_sg U69187 ( .A(n55629), .B(n57837), .X(n34588) );
  nand_x1_sg U69188 ( .A(n49403), .B(n57554), .X(n34341) );
  nand_x1_sg U69189 ( .A(n55627), .B(n57841), .X(n34342) );
  nand_x1_sg U69190 ( .A(n49405), .B(n57550), .X(n34343) );
  nand_x1_sg U69191 ( .A(n55625), .B(n57850), .X(n34344) );
  nand_x1_sg U69192 ( .A(n49407), .B(n57550), .X(n34533) );
  nand_x1_sg U69193 ( .A(n55623), .B(n57843), .X(n34534) );
  nand_x1_sg U69194 ( .A(n49409), .B(n57558), .X(n34527) );
  nand_x1_sg U69195 ( .A(n55621), .B(n57840), .X(n34528) );
  nand_x1_sg U69196 ( .A(n49411), .B(n57551), .X(n34479) );
  nand_x1_sg U69197 ( .A(n55619), .B(n57846), .X(n34480) );
  nand_x1_sg U69198 ( .A(n49413), .B(n57533), .X(n34345) );
  nand_x1_sg U69199 ( .A(n55617), .B(n57827), .X(n34346) );
  nand_x1_sg U69200 ( .A(n49415), .B(n57550), .X(n34485) );
  nand_x1_sg U69201 ( .A(n55615), .B(n57844), .X(n34486) );
  nand_x1_sg U69202 ( .A(n49417), .B(n57530), .X(n34461) );
  nand_x1_sg U69203 ( .A(n55613), .B(n57840), .X(n34462) );
  nand_x1_sg U69204 ( .A(n49419), .B(n57534), .X(n34497) );
  nand_x1_sg U69205 ( .A(n55611), .B(n57839), .X(n34498) );
  nand_x1_sg U69206 ( .A(n49421), .B(n57550), .X(n34515) );
  nand_x1_sg U69207 ( .A(n55609), .B(n57844), .X(n34516) );
  nand_x1_sg U69208 ( .A(n49423), .B(n57538), .X(n34545) );
  nand_x1_sg U69209 ( .A(n55607), .B(n57850), .X(n34546) );
  nand_x1_sg U69210 ( .A(n49425), .B(n57534), .X(n34521) );
  nand_x1_sg U69211 ( .A(n55605), .B(n57841), .X(n34522) );
  nand_x1_sg U69212 ( .A(n49427), .B(n57533), .X(n34503) );
  nand_x1_sg U69213 ( .A(n55603), .B(n57837), .X(n34504) );
  nand_x1_sg U69214 ( .A(n49429), .B(n57533), .X(n34509) );
  nand_x1_sg U69215 ( .A(n55601), .B(n57836), .X(n34510) );
  nand_x1_sg U69216 ( .A(n49431), .B(n57550), .X(n34539) );
  nand_x1_sg U69217 ( .A(n55599), .B(n57838), .X(n34540) );
  nand_x1_sg U69218 ( .A(n49433), .B(n57558), .X(n34491) );
  nand_x1_sg U69219 ( .A(n55597), .B(n57849), .X(n34492) );
  nand_x1_sg U69220 ( .A(n49447), .B(n57554), .X(n34673) );
  nand_x1_sg U69221 ( .A(n55583), .B(n57838), .X(n34674) );
  nand_x1_sg U69222 ( .A(n49449), .B(n57533), .X(n34695) );
  nand_x1_sg U69223 ( .A(n55581), .B(n57846), .X(n34696) );
  nand_x1_sg U69224 ( .A(n49453), .B(n57554), .X(n34389) );
  nand_x1_sg U69225 ( .A(n55577), .B(n34232), .X(n34390) );
  nand_x1_sg U69226 ( .A(n49467), .B(n57554), .X(n34621) );
  nand_x1_sg U69227 ( .A(n55563), .B(n57844), .X(n34622) );
  nand_x1_sg U69228 ( .A(n49469), .B(n57546), .X(n34667) );
  nand_x1_sg U69229 ( .A(n55561), .B(n57839), .X(n34668) );
  nand_x1_sg U69230 ( .A(n49471), .B(n57547), .X(n34645) );
  nand_x1_sg U69231 ( .A(n55559), .B(n57841), .X(n34646) );
  nand_x1_sg U69232 ( .A(n49473), .B(n57558), .X(n34627) );
  nand_x1_sg U69233 ( .A(n55557), .B(n57846), .X(n34628) );
  nand_x1_sg U69234 ( .A(n49475), .B(n57546), .X(n34661) );
  nand_x1_sg U69235 ( .A(n55555), .B(n57841), .X(n34662) );
  nand_x1_sg U69236 ( .A(n49479), .B(n57547), .X(n34639) );
  nand_x1_sg U69237 ( .A(n55551), .B(n57842), .X(n34640) );
  nand_x1_sg U69238 ( .A(n49481), .B(n57534), .X(n34633) );
  nand_x1_sg U69239 ( .A(n55549), .B(n46204), .X(n34634) );
  nand_x1_sg U69240 ( .A(n49483), .B(n57535), .X(n34263) );
  nand_x1_sg U69241 ( .A(n55547), .B(n57842), .X(n34264) );
  nand_x1_sg U69242 ( .A(n49485), .B(n57536), .X(n34261) );
  nand_x1_sg U69243 ( .A(n55545), .B(n57844), .X(n34262) );
  nand_x1_sg U69244 ( .A(n49487), .B(n57557), .X(n34685) );
  nand_x1_sg U69245 ( .A(n55543), .B(n57824), .X(n34686) );
  nand_x1_sg U69246 ( .A(n49489), .B(n57534), .X(n34679) );
  nand_x1_sg U69247 ( .A(n55541), .B(n57849), .X(n34680) );
  nand_x1_sg U69248 ( .A(n49491), .B(n57547), .X(n34651) );
  nand_x1_sg U69249 ( .A(n55539), .B(n57842), .X(n34652) );
  nand_x1_sg U69250 ( .A(n49493), .B(n57537), .X(n34265) );
  nand_x1_sg U69251 ( .A(n55537), .B(n57837), .X(n34266) );
  nand_x1_sg U69252 ( .A(n49497), .B(n57533), .X(n34369) );
  nand_x1_sg U69253 ( .A(n55533), .B(n57826), .X(n34370) );
  nand_x1_sg U69254 ( .A(n49509), .B(n57551), .X(n34277) );
  nand_x1_sg U69255 ( .A(n55521), .B(n57842), .X(n34278) );
  nand_x1_sg U69256 ( .A(n49511), .B(n57558), .X(n34381) );
  nand_x1_sg U69257 ( .A(n55519), .B(n57849), .X(n34382) );
  nand_x1_sg U69258 ( .A(n49515), .B(n57532), .X(n34413) );
  nand_x1_sg U69259 ( .A(n55515), .B(n46204), .X(n34414) );
  nand_x1_sg U69260 ( .A(n49121), .B(n57550), .X(n34283) );
  nand_x1_sg U69261 ( .A(n55513), .B(n57844), .X(n34284) );
  nand_x1_sg U69262 ( .A(n49123), .B(n57532), .X(n34407) );
  nand_x1_sg U69263 ( .A(n55511), .B(n57844), .X(n34408) );
  nand_x1_sg U69264 ( .A(n49127), .B(n57533), .X(n34285) );
  nand_x1_sg U69265 ( .A(n55507), .B(n57844), .X(n34286) );
  nand_x1_sg U69266 ( .A(n49131), .B(n57554), .X(n34281) );
  nand_x1_sg U69267 ( .A(n55503), .B(n57846), .X(n34282) );
  nand_x1_sg U69268 ( .A(n49167), .B(n57537), .X(n34425) );
  nand_x1_sg U69269 ( .A(n55467), .B(n57845), .X(n34426) );
  nand_x1_sg U69270 ( .A(n49169), .B(n57534), .X(n34321) );
  nand_x1_sg U69271 ( .A(n55465), .B(n57827), .X(n34322) );
  nand_x1_sg U69272 ( .A(n49171), .B(n57538), .X(n34419) );
  nand_x1_sg U69273 ( .A(n55463), .B(n46204), .X(n34420) );
  nand_x1_sg U69274 ( .A(n49175), .B(n57534), .X(n34317) );
  nand_x1_sg U69275 ( .A(n55459), .B(n57827), .X(n34318) );
  nand_x1_sg U69276 ( .A(n49177), .B(n57534), .X(n34319) );
  nand_x1_sg U69277 ( .A(n55457), .B(n57827), .X(n34320) );
  nand_x1_sg U69278 ( .A(n49179), .B(n57531), .X(n34443) );
  nand_x1_sg U69279 ( .A(n55455), .B(n57836), .X(n34444) );
  nand_x1_sg U69280 ( .A(n49181), .B(n57531), .X(n34437) );
  nand_x1_sg U69281 ( .A(n55453), .B(n57838), .X(n34438) );
  nand_x1_sg U69282 ( .A(n49183), .B(n57534), .X(n34323) );
  nand_x1_sg U69283 ( .A(n55451), .B(n57827), .X(n34324) );
  nand_x1_sg U69284 ( .A(n49185), .B(n57534), .X(n34325) );
  nand_x1_sg U69285 ( .A(n55449), .B(n57827), .X(n34326) );
  nand_x1_sg U69286 ( .A(n49187), .B(n57554), .X(n34473) );
  nand_x1_sg U69287 ( .A(n55447), .B(n57844), .X(n34474) );
  nand_x1_sg U69288 ( .A(n49189), .B(n57530), .X(n34467) );
  nand_x1_sg U69289 ( .A(n55445), .B(n57841), .X(n34468) );
  nand_x1_sg U69290 ( .A(n49191), .B(n57531), .X(n34449) );
  nand_x1_sg U69291 ( .A(n55443), .B(n57846), .X(n34450) );
  nand_x1_sg U69292 ( .A(n49193), .B(n57534), .X(n34327) );
  nand_x1_sg U69293 ( .A(n55441), .B(n57827), .X(n34328) );
  nand_x1_sg U69294 ( .A(n49195), .B(n57530), .X(n34455) );
  nand_x1_sg U69295 ( .A(n55439), .B(n57837), .X(n34456) );
  nand_x1_sg U69296 ( .A(n49197), .B(n57561), .X(n34431) );
  nand_x1_sg U69297 ( .A(n55437), .B(n57826), .X(n34432) );
  nand_x1_sg U69298 ( .A(n49201), .B(n57550), .X(n34311) );
  nand_x1_sg U69299 ( .A(n55433), .B(n57826), .X(n34312) );
  nand_x1_sg U69300 ( .A(n49203), .B(n57534), .X(n34329) );
  nand_x1_sg U69301 ( .A(n55431), .B(n57846), .X(n34330) );
  nand_x1_sg U69302 ( .A(n49205), .B(n57534), .X(n34313) );
  nand_x1_sg U69303 ( .A(n55429), .B(n57827), .X(n34314) );
  nand_x1_sg U69304 ( .A(n49207), .B(n57532), .X(n34403) );
  nand_x1_sg U69305 ( .A(n55427), .B(n57845), .X(n34404) );
  nand_x1_sg U69306 ( .A(n49209), .B(n57534), .X(n34315) );
  nand_x1_sg U69307 ( .A(n55425), .B(n57827), .X(n34316) );
  nand_x1_sg U69308 ( .A(n49211), .B(n57551), .X(n34395) );
  nand_x1_sg U69309 ( .A(n55423), .B(n57839), .X(n34396) );
  nand_x1_sg U69310 ( .A(n49213), .B(n57550), .X(n34377) );
  nand_x1_sg U69311 ( .A(n55421), .B(n57837), .X(n34378) );
  nand_x1_sg U69312 ( .A(n49217), .B(n57535), .X(n34293) );
  nand_x1_sg U69313 ( .A(n55417), .B(n57843), .X(n34294) );
  nand_x1_sg U69314 ( .A(n49219), .B(n57558), .X(n34299) );
  nand_x1_sg U69315 ( .A(n55415), .B(n57837), .X(n34300) );
  nand_x1_sg U69316 ( .A(n49221), .B(n57554), .X(n34371) );
  nand_x1_sg U69317 ( .A(n55413), .B(n57826), .X(n34372) );
  nand_x1_sg U69318 ( .A(n49223), .B(n57534), .X(n34383) );
  nand_x1_sg U69319 ( .A(n55411), .B(n57836), .X(n34384) );
  nand_x1_sg U69320 ( .A(n49225), .B(n57551), .X(n34305) );
  nand_x1_sg U69321 ( .A(n55409), .B(n57826), .X(n34306) );
  nand_x1_sg U69322 ( .A(n49227), .B(n57550), .X(n34287) );
  nand_x1_sg U69323 ( .A(n55407), .B(n57846), .X(n34288) );
  nand_x1_sg U69324 ( .A(n49229), .B(n57532), .X(n34405) );
  nand_x1_sg U69325 ( .A(n55405), .B(n57838), .X(n34406) );
  nand_x1_sg U69326 ( .A(n49295), .B(n57534), .X(n34347) );
  nand_x1_sg U69327 ( .A(n55339), .B(n57838), .X(n34348) );
  nand_x1_sg U69328 ( .A(n49297), .B(n57538), .X(n34273) );
  nand_x1_sg U69329 ( .A(n55337), .B(n57850), .X(n34274) );
  nand_x1_sg U69330 ( .A(n49301), .B(n57533), .X(n34339) );
  nand_x1_sg U69331 ( .A(n55333), .B(n46204), .X(n34340) );
  nand_x1_sg U69332 ( .A(n49305), .B(n57552), .X(n34275) );
  nand_x1_sg U69333 ( .A(n55329), .B(n57837), .X(n34276) );
  nand_x1_sg U69334 ( .A(n49307), .B(n57533), .X(n34365) );
  nand_x1_sg U69335 ( .A(n55327), .B(n57826), .X(n34366) );
  nand_x1_sg U69336 ( .A(n49309), .B(n57533), .X(n34279) );
  nand_x1_sg U69337 ( .A(n55325), .B(n57836), .X(n34280) );
  nand_x1_sg U69338 ( .A(n49317), .B(n57533), .X(n34351) );
  nand_x1_sg U69339 ( .A(n55317), .B(n57839), .X(n34352) );
  nand_x1_sg U69340 ( .A(n50049), .B(n57536), .X(n34233) );
  nand_x1_sg U69341 ( .A(n56169), .B(n57838), .X(n34234) );
  nand_x1_sg U69342 ( .A(n49869), .B(n57536), .X(n34237) );
  nand_x1_sg U69343 ( .A(n55953), .B(n57846), .X(n34238) );
  nand_x1_sg U69344 ( .A(n49873), .B(n57535), .X(n34241) );
  nand_x1_sg U69345 ( .A(n55949), .B(n57827), .X(n34242) );
  nand_x1_sg U69346 ( .A(n49641), .B(n57535), .X(n34245) );
  nand_x1_sg U69347 ( .A(n55785), .B(n57839), .X(n34246) );
  nand_x1_sg U69348 ( .A(n49687), .B(n57536), .X(n34235) );
  nand_x1_sg U69349 ( .A(n55739), .B(n57795), .X(n34236) );
  nand_x1_sg U69350 ( .A(n49329), .B(n57535), .X(n34243) );
  nand_x1_sg U69351 ( .A(n55701), .B(n57844), .X(n34244) );
  nand_x1_sg U69352 ( .A(n49333), .B(n57535), .X(n34247) );
  nand_x1_sg U69353 ( .A(n55697), .B(n57836), .X(n34248) );
  nand_x1_sg U69354 ( .A(n49477), .B(n57536), .X(n34239) );
  nand_x1_sg U69355 ( .A(n55553), .B(n57837), .X(n34240) );
  nand_x1_sg U69356 ( .A(n47409), .B(n57911), .X(n29326) );
  nand_x1_sg U69357 ( .A(n49643), .B(n57551), .X(n34230) );
  nand_x1_sg U69358 ( .A(n55783), .B(n46204), .X(n34231) );
  nand_x4_sg U69359 ( .A(n38411), .B(n39835), .X(n38415) );
  nor_x1_sg U69360 ( .A(state[0]), .B(state[1]), .X(n39836) );
  nand_x1_sg U69361 ( .A(n57522), .B(n49103), .X(n38743) );
  nand_x1_sg U69362 ( .A(n57519), .B(n49097), .X(n38735) );
  nand_x1_sg U69363 ( .A(n57522), .B(n49095), .X(n39193) );
  nand_x1_sg U69364 ( .A(n57523), .B(n49093), .X(n38737) );
  nand_x1_sg U69365 ( .A(n57522), .B(n49091), .X(n39199) );
  nand_x1_sg U69366 ( .A(n57527), .B(n49089), .X(n39205) );
  nand_x1_sg U69367 ( .A(n57520), .B(n49087), .X(n39211) );
  nand_x1_sg U69368 ( .A(n57523), .B(n49083), .X(n38745) );
  nand_x1_sg U69369 ( .A(n57519), .B(n49081), .X(n38747) );
  nand_x1_sg U69370 ( .A(n57526), .B(n49079), .X(n38739) );
  nand_x1_sg U69371 ( .A(n57519), .B(n49077), .X(n38741) );
  nand_x1_sg U69372 ( .A(n57520), .B(n48867), .X(n39129) );
  nand_x1_sg U69373 ( .A(n57520), .B(n48865), .X(n39131) );
  nand_x1_sg U69374 ( .A(n57524), .B(n48863), .X(n39123) );
  nand_x1_sg U69375 ( .A(n57522), .B(n48861), .X(n39125) );
  nand_x1_sg U69376 ( .A(n57520), .B(n48859), .X(n39141) );
  nand_x1_sg U69377 ( .A(n57520), .B(n48857), .X(n39143) );
  nand_x1_sg U69378 ( .A(n57520), .B(n48855), .X(n39135) );
  nand_x1_sg U69379 ( .A(n57520), .B(n48853), .X(n39137) );
  nand_x1_sg U69380 ( .A(n57524), .B(n48851), .X(n39105) );
  nand_x1_sg U69381 ( .A(n57524), .B(n48849), .X(n39107) );
  nand_x1_sg U69382 ( .A(n57524), .B(n48847), .X(n39099) );
  nand_x1_sg U69383 ( .A(n57522), .B(n48845), .X(n39101) );
  nand_x1_sg U69384 ( .A(n57524), .B(n48843), .X(n39117) );
  nand_x1_sg U69385 ( .A(n57521), .B(n48841), .X(n39119) );
  nand_x1_sg U69386 ( .A(n57519), .B(n48839), .X(n39111) );
  nand_x1_sg U69387 ( .A(n57525), .B(n48837), .X(n39113) );
  nand_x1_sg U69388 ( .A(n57527), .B(n48835), .X(n39177) );
  nand_x1_sg U69389 ( .A(n57520), .B(n48833), .X(n39179) );
  nand_x1_sg U69390 ( .A(n57523), .B(n48831), .X(n39171) );
  nand_x1_sg U69391 ( .A(n57525), .B(n48829), .X(n39173) );
  nand_x1_sg U69392 ( .A(n57521), .B(n48827), .X(n39189) );
  nand_x1_sg U69393 ( .A(n57523), .B(n48825), .X(n39191) );
  nand_x1_sg U69394 ( .A(n57521), .B(n48823), .X(n39183) );
  nand_x1_sg U69395 ( .A(n57523), .B(n48821), .X(n39185) );
  nand_x1_sg U69396 ( .A(n57521), .B(n48819), .X(n39153) );
  nand_x1_sg U69397 ( .A(n57523), .B(n48817), .X(n39155) );
  nand_x1_sg U69398 ( .A(n57525), .B(n48815), .X(n39147) );
  nand_x1_sg U69399 ( .A(n57519), .B(n48813), .X(n39149) );
  nand_x1_sg U69400 ( .A(n57525), .B(n48811), .X(n39165) );
  nand_x1_sg U69401 ( .A(n57520), .B(n48809), .X(n39167) );
  nand_x1_sg U69402 ( .A(n57524), .B(n48807), .X(n39159) );
  nand_x1_sg U69403 ( .A(n57525), .B(n48805), .X(n39161) );
  nand_x1_sg U69404 ( .A(n57522), .B(n48803), .X(n38943) );
  nand_x1_sg U69405 ( .A(n57522), .B(n48801), .X(n38945) );
  nand_x1_sg U69406 ( .A(n57522), .B(n48799), .X(n38937) );
  nand_x1_sg U69407 ( .A(n57522), .B(n48797), .X(n38939) );
  nand_x1_sg U69408 ( .A(n57521), .B(n48795), .X(n39035) );
  nand_x1_sg U69409 ( .A(n57521), .B(n48793), .X(n38891) );
  nand_x1_sg U69410 ( .A(n57520), .B(n48789), .X(n38689) );
  nand_x1_sg U69411 ( .A(n57526), .B(n48771), .X(n39081) );
  nand_x1_sg U69412 ( .A(n57524), .B(n48769), .X(n39083) );
  nand_x1_sg U69413 ( .A(n57521), .B(n48767), .X(n39075) );
  nand_x1_sg U69414 ( .A(n57524), .B(n48765), .X(n39077) );
  nand_x1_sg U69415 ( .A(n57520), .B(n48763), .X(n39093) );
  nand_x1_sg U69416 ( .A(n57524), .B(n48761), .X(n39095) );
  nand_x1_sg U69417 ( .A(n57519), .B(n48759), .X(n39087) );
  nand_x1_sg U69418 ( .A(n57519), .B(n48757), .X(n39089) );
  nand_x1_sg U69419 ( .A(n57520), .B(n48755), .X(n38917) );
  nand_x1_sg U69420 ( .A(n57521), .B(n48753), .X(n38979) );
  nand_x1_sg U69421 ( .A(n57522), .B(n48751), .X(n39053) );
  nand_x1_sg U69422 ( .A(n57519), .B(n48749), .X(n38985) );
  nand_x1_sg U69423 ( .A(n57522), .B(n48747), .X(n38931) );
  nand_x1_sg U69424 ( .A(n57522), .B(n48745), .X(n38933) );
  nand_x1_sg U69425 ( .A(n57526), .B(n48743), .X(n38925) );
  nand_x1_sg U69426 ( .A(n57523), .B(n48741), .X(n38927) );
  nand_x1_sg U69427 ( .A(n57521), .B(n48675), .X(n39225) );
  nand_x1_sg U69428 ( .A(n57527), .B(n48673), .X(n39227) );
  nand_x1_sg U69429 ( .A(n57519), .B(n48671), .X(n39219) );
  nand_x1_sg U69430 ( .A(n57527), .B(n48669), .X(n39221) );
  nand_x1_sg U69431 ( .A(n57520), .B(n48667), .X(n39237) );
  nand_x1_sg U69432 ( .A(n57520), .B(n48665), .X(n39239) );
  nand_x1_sg U69433 ( .A(n57519), .B(n48663), .X(n39231) );
  nand_x1_sg U69434 ( .A(n57526), .B(n48661), .X(n39233) );
  nand_x1_sg U69435 ( .A(n57521), .B(n48659), .X(n39201) );
  nand_x1_sg U69436 ( .A(n57520), .B(n48657), .X(n39203) );
  nand_x1_sg U69437 ( .A(n57526), .B(n48655), .X(n39195) );
  nand_x1_sg U69438 ( .A(n57523), .B(n48653), .X(n39197) );
  nand_x1_sg U69439 ( .A(n57519), .B(n48651), .X(n39213) );
  nand_x1_sg U69440 ( .A(n57522), .B(n48649), .X(n39215) );
  nand_x1_sg U69441 ( .A(n57521), .B(n48647), .X(n39207) );
  nand_x1_sg U69442 ( .A(n57522), .B(n48645), .X(n39209) );
  nand_x1_sg U69443 ( .A(n57520), .B(n48627), .X(n39249) );
  nand_x1_sg U69444 ( .A(n57520), .B(n48625), .X(n39251) );
  nand_x1_sg U69445 ( .A(n57520), .B(n48623), .X(n39243) );
  nand_x1_sg U69446 ( .A(n57520), .B(n48621), .X(n39245) );
  nand_x1_sg U69447 ( .A(n57520), .B(n48615), .X(n39255) );
  nand_x1_sg U69448 ( .A(n57520), .B(n48613), .X(n39257) );
  nand_x1_sg U69449 ( .A(n57520), .B(n48543), .X(n39241) );
  nand_x1_sg U69450 ( .A(n57520), .B(n48541), .X(n39259) );
  nand_x1_sg U69451 ( .A(n57521), .B(n48483), .X(n38695) );
  nand_x1_sg U69452 ( .A(n57524), .B(n48475), .X(n38705) );
  nand_x1_sg U69453 ( .A(n57524), .B(n48473), .X(n38707) );
  nand_x1_sg U69454 ( .A(n57521), .B(n48471), .X(n38699) );
  nand_x1_sg U69455 ( .A(n57526), .B(n48469), .X(n38701) );
  nand_x1_sg U69456 ( .A(n57523), .B(n48459), .X(n38691) );
  nand_x1_sg U69457 ( .A(n57526), .B(n48457), .X(n38693) );
  nand_x1_sg U69458 ( .A(n57526), .B(n48455), .X(n38685) );
  nand_x1_sg U69459 ( .A(n57525), .B(n48453), .X(n38687) );
  nand_x1_sg U69460 ( .A(n57520), .B(n48441), .X(n38709) );
  nand_x1_sg U69461 ( .A(n57526), .B(n48439), .X(n38727) );
  nand_x1_sg U69462 ( .A(n57526), .B(n48435), .X(n38717) );
  nand_x1_sg U69463 ( .A(n57519), .B(n48433), .X(n38703) );
  nand_x1_sg U69464 ( .A(n57526), .B(n48431), .X(n38719) );
  nand_x1_sg U69465 ( .A(n57526), .B(n48429), .X(n38721) );
  nand_x1_sg U69466 ( .A(n57521), .B(n48427), .X(n38713) );
  nand_x1_sg U69467 ( .A(n57519), .B(n48425), .X(n38715) );
  nand_x1_sg U69468 ( .A(n57523), .B(n48423), .X(n38711) );
  nand_x1_sg U69469 ( .A(n57525), .B(n48421), .X(n38697) );
  nand_x1_sg U69470 ( .A(n57519), .B(n48355), .X(n39187) );
  nand_x1_sg U69471 ( .A(n57520), .B(n48329), .X(n39253) );
  nand_x1_sg U69472 ( .A(n57522), .B(n48289), .X(n38935) );
  nand_x1_sg U69473 ( .A(n57519), .B(n48285), .X(n39109) );
  nand_x1_sg U69474 ( .A(n57521), .B(n48283), .X(n39115) );
  nand_x1_sg U69475 ( .A(n57520), .B(n48281), .X(n39133) );
  nand_x1_sg U69476 ( .A(n57520), .B(n48277), .X(n39139) );
  nand_x1_sg U69477 ( .A(n57525), .B(n48259), .X(n39151) );
  nand_x1_sg U69478 ( .A(n57523), .B(n48257), .X(n39157) );
  nand_x1_sg U69479 ( .A(n57519), .B(n48253), .X(n39175) );
  nand_x1_sg U69480 ( .A(n57525), .B(n48251), .X(n39145) );
  nand_x1_sg U69481 ( .A(n57526), .B(n48249), .X(n39169) );
  nand_x1_sg U69482 ( .A(n57521), .B(n48247), .X(n39163) );
  nand_x1_sg U69483 ( .A(n57524), .B(n48245), .X(n39181) );
  nand_x1_sg U69484 ( .A(n57525), .B(n48241), .X(n39071) );
  nand_x1_sg U69485 ( .A(n57523), .B(n48239), .X(n39085) );
  nand_x1_sg U69486 ( .A(n57519), .B(n48237), .X(n39091) );
  nand_x1_sg U69487 ( .A(n57524), .B(n48235), .X(n39073) );
  nand_x1_sg U69488 ( .A(n57522), .B(n48233), .X(n38941) );
  nand_x1_sg U69489 ( .A(n57523), .B(n48231), .X(n39103) );
  nand_x1_sg U69490 ( .A(n57520), .B(n48229), .X(n39079) );
  nand_x1_sg U69491 ( .A(n57520), .B(n48227), .X(n39127) );
  nand_x1_sg U69492 ( .A(n57526), .B(n48225), .X(n39217) );
  nand_x1_sg U69493 ( .A(n57521), .B(n48223), .X(n39223) );
  nand_x1_sg U69494 ( .A(n57526), .B(n48221), .X(n39229) );
  nand_x1_sg U69495 ( .A(n57526), .B(n48217), .X(n38839) );
  nand_x1_sg U69496 ( .A(n57522), .B(n48215), .X(n38929) );
  nand_x1_sg U69497 ( .A(n57524), .B(n48213), .X(n39097) );
  nand_x1_sg U69498 ( .A(n57523), .B(n48211), .X(n38827) );
  nand_x1_sg U69499 ( .A(n57524), .B(n48209), .X(n38833) );
  nand_x1_sg U69500 ( .A(n57522), .B(n48207), .X(n39059) );
  nand_x1_sg U69501 ( .A(n57519), .B(n48205), .X(n38877) );
  nand_x1_sg U69502 ( .A(n57519), .B(n48203), .X(n38803) );
  nand_x1_sg U69503 ( .A(n57523), .B(n48201), .X(n38809) );
  nand_x1_sg U69504 ( .A(n57525), .B(n48199), .X(n38815) );
  nand_x1_sg U69505 ( .A(n57524), .B(n48197), .X(n38821) );
  nand_x1_sg U69506 ( .A(n57520), .B(n48183), .X(n39235) );
  nand_x1_sg U69507 ( .A(n57524), .B(n48175), .X(n39121) );
  nand_x1_sg U69508 ( .A(n57525), .B(n48173), .X(n38923) );
  nand_x1_sg U69509 ( .A(n57520), .B(n48139), .X(n39247) );
  nand_x1_sg U69510 ( .A(n57525), .B(n48131), .X(n38779) );
  nand_x1_sg U69511 ( .A(n57520), .B(n48129), .X(n38785) );
  nand_x1_sg U69512 ( .A(n57526), .B(n48123), .X(n38755) );
  nand_x1_sg U69513 ( .A(n57520), .B(n48121), .X(n38761) );
  nand_x1_sg U69514 ( .A(n57522), .B(n48119), .X(n38767) );
  nand_x1_sg U69515 ( .A(n57527), .B(n48117), .X(n38773) );
  nand_x1_sg U69516 ( .A(n57525), .B(n48111), .X(n38749) );
  nand_x1_sg U69517 ( .A(n57525), .B(n48107), .X(n38791) );
  nand_x1_sg U69518 ( .A(n57522), .B(n48105), .X(n38797) );
  nand_x1_sg U69519 ( .A(n57521), .B(n48099), .X(n38867) );
  nand_x1_sg U69520 ( .A(n57519), .B(n48097), .X(n38869) );
  nand_x1_sg U69521 ( .A(n57522), .B(n48095), .X(n38861) );
  nand_x1_sg U69522 ( .A(n57522), .B(n48093), .X(n38863) );
  nand_x1_sg U69523 ( .A(n57521), .B(n48091), .X(n38879) );
  nand_x1_sg U69524 ( .A(n57520), .B(n48089), .X(n38881) );
  nand_x1_sg U69525 ( .A(n57526), .B(n48087), .X(n38873) );
  nand_x1_sg U69526 ( .A(n57522), .B(n48085), .X(n38875) );
  nand_x1_sg U69527 ( .A(n57527), .B(n48083), .X(n38855) );
  nand_x1_sg U69528 ( .A(n57523), .B(n48081), .X(n38857) );
  nand_x1_sg U69529 ( .A(n57525), .B(n48079), .X(n38849) );
  nand_x1_sg U69530 ( .A(n57526), .B(n48077), .X(n38851) );
  nand_x1_sg U69531 ( .A(n57524), .B(n48075), .X(n38729) );
  nand_x1_sg U69532 ( .A(n57521), .B(n48073), .X(n38853) );
  nand_x1_sg U69533 ( .A(n57520), .B(n48071), .X(n38845) );
  nand_x1_sg U69534 ( .A(n57521), .B(n48069), .X(n38847) );
  nand_x1_sg U69535 ( .A(n57523), .B(n48067), .X(n38907) );
  nand_x1_sg U69536 ( .A(n57524), .B(n48065), .X(n38909) );
  nand_x1_sg U69537 ( .A(n57520), .B(n48063), .X(n38901) );
  nand_x1_sg U69538 ( .A(n57523), .B(n48061), .X(n38903) );
  nand_x1_sg U69539 ( .A(n57523), .B(n48059), .X(n38905) );
  nand_x1_sg U69540 ( .A(n57523), .B(n48057), .X(n38885) );
  nand_x1_sg U69541 ( .A(n57522), .B(n48055), .X(n38897) );
  nand_x1_sg U69542 ( .A(n57519), .B(n48053), .X(n38899) );
  nand_x1_sg U69543 ( .A(n57519), .B(n48051), .X(n38871) );
  nand_x1_sg U69544 ( .A(n57519), .B(n48049), .X(n38859) );
  nand_x1_sg U69545 ( .A(n57522), .B(n48047), .X(n38883) );
  nand_x1_sg U69546 ( .A(n57527), .B(n48045), .X(n38865) );
  nand_x1_sg U69547 ( .A(n57522), .B(n48043), .X(n38893) );
  nand_x1_sg U69548 ( .A(n57525), .B(n48041), .X(n38895) );
  nand_x1_sg U69549 ( .A(n57521), .B(n48039), .X(n38887) );
  nand_x1_sg U69550 ( .A(n57519), .B(n48037), .X(n38889) );
  nand_x1_sg U69551 ( .A(n57520), .B(n48035), .X(n38781) );
  nand_x1_sg U69552 ( .A(n57522), .B(n48033), .X(n38783) );
  nand_x1_sg U69553 ( .A(n57519), .B(n48031), .X(n38775) );
  nand_x1_sg U69554 ( .A(n57524), .B(n48029), .X(n38777) );
  nand_x1_sg U69555 ( .A(n57522), .B(n48027), .X(n38793) );
  nand_x1_sg U69556 ( .A(n57521), .B(n48025), .X(n38795) );
  nand_x1_sg U69557 ( .A(n57525), .B(n48023), .X(n38787) );
  nand_x1_sg U69558 ( .A(n57525), .B(n48021), .X(n38789) );
  nand_x1_sg U69559 ( .A(n57522), .B(n48019), .X(n38757) );
  nand_x1_sg U69560 ( .A(n57523), .B(n48017), .X(n38759) );
  nand_x1_sg U69561 ( .A(n57526), .B(n48015), .X(n38751) );
  nand_x1_sg U69562 ( .A(n57521), .B(n48013), .X(n38753) );
  nand_x1_sg U69563 ( .A(n57523), .B(n48011), .X(n38769) );
  nand_x1_sg U69564 ( .A(n57521), .B(n48009), .X(n38771) );
  nand_x1_sg U69565 ( .A(n57524), .B(n48007), .X(n38763) );
  nand_x1_sg U69566 ( .A(n57523), .B(n48005), .X(n38765) );
  nand_x1_sg U69567 ( .A(n57522), .B(n48003), .X(n38829) );
  nand_x1_sg U69568 ( .A(n57523), .B(n48001), .X(n38831) );
  nand_x1_sg U69569 ( .A(n57524), .B(n47999), .X(n38823) );
  nand_x1_sg U69570 ( .A(n57524), .B(n47997), .X(n38825) );
  nand_x1_sg U69571 ( .A(n57519), .B(n47995), .X(n38841) );
  nand_x1_sg U69572 ( .A(n57522), .B(n47993), .X(n38843) );
  nand_x1_sg U69573 ( .A(n57526), .B(n47991), .X(n38835) );
  nand_x1_sg U69574 ( .A(n57526), .B(n47989), .X(n38837) );
  nand_x1_sg U69575 ( .A(n57520), .B(n47987), .X(n38805) );
  nand_x1_sg U69576 ( .A(n57520), .B(n47985), .X(n38807) );
  nand_x1_sg U69577 ( .A(n57527), .B(n47983), .X(n38799) );
  nand_x1_sg U69578 ( .A(n57519), .B(n47981), .X(n38801) );
  nand_x1_sg U69579 ( .A(n57522), .B(n47979), .X(n38817) );
  nand_x1_sg U69580 ( .A(n57520), .B(n47977), .X(n38819) );
  nand_x1_sg U69581 ( .A(n57521), .B(n47975), .X(n38811) );
  nand_x1_sg U69582 ( .A(n57521), .B(n47973), .X(n38813) );
  nand_x1_sg U69583 ( .A(n57523), .B(n47971), .X(n39037) );
  nand_x1_sg U69584 ( .A(n57520), .B(n47969), .X(n39039) );
  nand_x1_sg U69585 ( .A(n57527), .B(n47967), .X(n39031) );
  nand_x1_sg U69586 ( .A(n57519), .B(n47965), .X(n39033) );
  nand_x1_sg U69587 ( .A(n57521), .B(n47963), .X(n39015) );
  nand_x1_sg U69588 ( .A(n57524), .B(n47961), .X(n39029) );
  nand_x1_sg U69589 ( .A(n57526), .B(n47959), .X(n39017) );
  nand_x1_sg U69590 ( .A(n57527), .B(n47957), .X(n39019) );
  nand_x1_sg U69591 ( .A(n57525), .B(n47955), .X(n39011) );
  nand_x1_sg U69592 ( .A(n57525), .B(n47953), .X(n39013) );
  nand_x1_sg U69593 ( .A(n57527), .B(n47951), .X(n39007) );
  nand_x1_sg U69594 ( .A(n57523), .B(n47949), .X(n39009) );
  nand_x1_sg U69595 ( .A(n57527), .B(n47947), .X(n39023) );
  nand_x1_sg U69596 ( .A(n57524), .B(n47945), .X(n39025) );
  nand_x1_sg U69597 ( .A(n57527), .B(n47943), .X(n39005) );
  nand_x1_sg U69598 ( .A(n57522), .B(n47941), .X(n39021) );
  nand_x1_sg U69599 ( .A(n57519), .B(n47939), .X(n39069) );
  nand_x1_sg U69600 ( .A(n57527), .B(n47937), .X(n39027) );
  nand_x1_sg U69601 ( .A(n57523), .B(n47935), .X(n39041) );
  nand_x1_sg U69602 ( .A(n57525), .B(n47933), .X(n39047) );
  nand_x1_sg U69603 ( .A(n57519), .B(n47931), .X(n38723) );
  nand_x1_sg U69604 ( .A(n57519), .B(n47929), .X(n38725) );
  nand_x1_sg U69605 ( .A(n57524), .B(n47927), .X(n39065) );
  nand_x1_sg U69606 ( .A(n57526), .B(n47925), .X(n39067) );
  nand_x1_sg U69607 ( .A(n57522), .B(n47923), .X(n39049) );
  nand_x1_sg U69608 ( .A(n57525), .B(n47921), .X(n39051) );
  nand_x1_sg U69609 ( .A(n57526), .B(n47919), .X(n39043) );
  nand_x1_sg U69610 ( .A(n57519), .B(n47917), .X(n39045) );
  nand_x1_sg U69611 ( .A(n57520), .B(n47915), .X(n39061) );
  nand_x1_sg U69612 ( .A(n57522), .B(n47913), .X(n39063) );
  nand_x1_sg U69613 ( .A(n57525), .B(n47911), .X(n39055) );
  nand_x1_sg U69614 ( .A(n57526), .B(n47909), .X(n39057) );
  nand_x1_sg U69615 ( .A(n57526), .B(n47907), .X(n38963) );
  nand_x1_sg U69616 ( .A(n57521), .B(n47905), .X(n38965) );
  nand_x1_sg U69617 ( .A(n57523), .B(n47903), .X(n38957) );
  nand_x1_sg U69618 ( .A(n57524), .B(n47901), .X(n38959) );
  nand_x1_sg U69619 ( .A(n57521), .B(n47899), .X(n38967) );
  nand_x1_sg U69620 ( .A(n57519), .B(n47897), .X(n38955) );
  nand_x1_sg U69621 ( .A(n57521), .B(n47895), .X(n38961) );
  nand_x1_sg U69622 ( .A(n57520), .B(n47893), .X(n38953) );
  nand_x1_sg U69623 ( .A(n57526), .B(n47891), .X(n38919) );
  nand_x1_sg U69624 ( .A(n57523), .B(n47889), .X(n38921) );
  nand_x1_sg U69625 ( .A(n57522), .B(n47887), .X(n38913) );
  nand_x1_sg U69626 ( .A(n57522), .B(n47885), .X(n38915) );
  nand_x1_sg U69627 ( .A(n57522), .B(n47883), .X(n38947) );
  nand_x1_sg U69628 ( .A(n57527), .B(n47881), .X(n38911) );
  nand_x1_sg U69629 ( .A(n57526), .B(n47879), .X(n38949) );
  nand_x1_sg U69630 ( .A(n57527), .B(n47877), .X(n38951) );
  nand_x1_sg U69631 ( .A(n57521), .B(n47875), .X(n38973) );
  nand_x1_sg U69632 ( .A(n57524), .B(n47873), .X(n38991) );
  nand_x1_sg U69633 ( .A(n57527), .B(n47871), .X(n38993) );
  nand_x1_sg U69634 ( .A(n57519), .B(n47869), .X(n38999) );
  nand_x1_sg U69635 ( .A(n57524), .B(n47867), .X(n39001) );
  nand_x1_sg U69636 ( .A(n57527), .B(n47865), .X(n39003) );
  nand_x1_sg U69637 ( .A(n57523), .B(n47863), .X(n38995) );
  nand_x1_sg U69638 ( .A(n57523), .B(n47861), .X(n38997) );
  nand_x1_sg U69639 ( .A(n57521), .B(n47859), .X(n38975) );
  nand_x1_sg U69640 ( .A(n57521), .B(n47857), .X(n38977) );
  nand_x1_sg U69641 ( .A(n57521), .B(n47855), .X(n38969) );
  nand_x1_sg U69642 ( .A(n57521), .B(n47853), .X(n38971) );
  nand_x1_sg U69643 ( .A(n57521), .B(n47851), .X(n38987) );
  nand_x1_sg U69644 ( .A(n57519), .B(n47849), .X(n38989) );
  nand_x1_sg U69645 ( .A(n57521), .B(n47847), .X(n38981) );
  nand_x1_sg U69646 ( .A(n57522), .B(n47845), .X(n38983) );
  nand_x1_sg U69647 ( .A(n57521), .B(n47843), .X(n38731) );
  nand_x1_sg U69648 ( .A(n57524), .B(n47841), .X(n38733) );
  nand_x1_sg U69649 ( .A(n57519), .B(n47791), .X(n39810) );
  nand_x1_sg U69650 ( .A(n57519), .B(n47789), .X(n39812) );
  nand_x1_sg U69651 ( .A(n57519), .B(n47787), .X(n39814) );
  nand_x1_sg U69652 ( .A(n57519), .B(n47785), .X(n39816) );
  nand_x1_sg U69653 ( .A(n57519), .B(n47783), .X(n39818) );
  nand_x1_sg U69654 ( .A(n57527), .B(n47781), .X(n39820) );
  nand_x1_sg U69655 ( .A(n57527), .B(n47779), .X(n39822) );
  nand_x1_sg U69656 ( .A(n57520), .B(n47777), .X(n39824) );
  nand_x1_sg U69657 ( .A(n57522), .B(n51567), .X(n39826) );
  nand_x1_sg U69658 ( .A(n57526), .B(n49119), .X(n38647) );
  nand_x1_sg U69659 ( .A(n57519), .B(n49109), .X(n38641) );
  nand_x1_sg U69660 ( .A(n57520), .B(n48791), .X(n38635) );
  nand_x1_sg U69661 ( .A(n57525), .B(n48787), .X(n38649) );
  nand_x1_sg U69662 ( .A(n57520), .B(n48785), .X(n38651) );
  nand_x1_sg U69663 ( .A(n57526), .B(n48783), .X(n38643) );
  nand_x1_sg U69664 ( .A(n57521), .B(n48781), .X(n38645) );
  nand_x1_sg U69665 ( .A(n57523), .B(n48779), .X(n38661) );
  nand_x1_sg U69666 ( .A(n57519), .B(n48777), .X(n38663) );
  nand_x1_sg U69667 ( .A(n57525), .B(n48775), .X(n38655) );
  nand_x1_sg U69668 ( .A(n57520), .B(n48773), .X(n38657) );
  nand_x1_sg U69669 ( .A(n57523), .B(n48611), .X(n38541) );
  nand_x1_sg U69670 ( .A(n57523), .B(n48609), .X(n38543) );
  nand_x1_sg U69671 ( .A(n57523), .B(n48607), .X(n38535) );
  nand_x1_sg U69672 ( .A(n57523), .B(n48605), .X(n38537) );
  nand_x1_sg U69673 ( .A(n57523), .B(n48603), .X(n38539) );
  nand_x1_sg U69674 ( .A(n57521), .B(n48601), .X(n38519) );
  nand_x1_sg U69675 ( .A(n57519), .B(n48599), .X(n38531) );
  nand_x1_sg U69676 ( .A(n57523), .B(n48597), .X(n38533) );
  nand_x1_sg U69677 ( .A(n57519), .B(n48595), .X(n38505) );
  nand_x1_sg U69678 ( .A(n57525), .B(n48593), .X(n38511) );
  nand_x1_sg U69679 ( .A(n57526), .B(n48591), .X(n38517) );
  nand_x1_sg U69680 ( .A(n57522), .B(n48589), .X(n38503) );
  nand_x1_sg U69681 ( .A(n57522), .B(n48587), .X(n38527) );
  nand_x1_sg U69682 ( .A(n57525), .B(n48585), .X(n38529) );
  nand_x1_sg U69683 ( .A(n57520), .B(n48583), .X(n38521) );
  nand_x1_sg U69684 ( .A(n57523), .B(n48581), .X(n38523) );
  nand_x1_sg U69685 ( .A(n57522), .B(n48579), .X(n38569) );
  nand_x1_sg U69686 ( .A(n57522), .B(n48577), .X(n38571) );
  nand_x1_sg U69687 ( .A(n57522), .B(n48575), .X(n38563) );
  nand_x1_sg U69688 ( .A(n57522), .B(n48573), .X(n38565) );
  nand_x1_sg U69689 ( .A(n57522), .B(n48571), .X(n38579) );
  nand_x1_sg U69690 ( .A(n57522), .B(n48569), .X(n38573) );
  nand_x1_sg U69691 ( .A(n57520), .B(n48567), .X(n38561) );
  nand_x1_sg U69692 ( .A(n57521), .B(n48565), .X(n38559) );
  nand_x1_sg U69693 ( .A(n57519), .B(n48563), .X(n38555) );
  nand_x1_sg U69694 ( .A(n57524), .B(n48561), .X(n38557) );
  nand_x1_sg U69695 ( .A(n57523), .B(n48559), .X(n38549) );
  nand_x1_sg U69696 ( .A(n57522), .B(n48557), .X(n38551) );
  nand_x1_sg U69697 ( .A(n57523), .B(n48555), .X(n38567) );
  nand_x1_sg U69698 ( .A(n57523), .B(n48553), .X(n38547) );
  nand_x1_sg U69699 ( .A(n57523), .B(n48551), .X(n38553) );
  nand_x1_sg U69700 ( .A(n57523), .B(n48549), .X(n38545) );
  nand_x1_sg U69701 ( .A(n57521), .B(n48531), .X(n38483) );
  nand_x1_sg U69702 ( .A(n57519), .B(n48529), .X(n38467) );
  nand_x1_sg U69703 ( .A(n57524), .B(n48525), .X(n38461) );
  nand_x1_sg U69704 ( .A(n57525), .B(n48523), .X(n38469) );
  nand_x1_sg U69705 ( .A(n57526), .B(n48519), .X(n38463) );
  nand_x1_sg U69706 ( .A(n57521), .B(n48517), .X(n38465) );
  nand_x1_sg U69707 ( .A(n57519), .B(n48515), .X(n38475) );
  nand_x1_sg U69708 ( .A(n57524), .B(n48513), .X(n38477) );
  nand_x1_sg U69709 ( .A(n57522), .B(n48511), .X(n38473) );
  nand_x1_sg U69710 ( .A(n57519), .B(n48509), .X(n38485) );
  nand_x1_sg U69711 ( .A(n57523), .B(n48507), .X(n38513) );
  nand_x1_sg U69712 ( .A(n57522), .B(n48505), .X(n38515) );
  nand_x1_sg U69713 ( .A(n57527), .B(n48503), .X(n38507) );
  nand_x1_sg U69714 ( .A(n57526), .B(n48501), .X(n38509) );
  nand_x1_sg U69715 ( .A(n57521), .B(n48499), .X(n38493) );
  nand_x1_sg U69716 ( .A(n57522), .B(n48497), .X(n38495) );
  nand_x1_sg U69717 ( .A(n57522), .B(n48495), .X(n38487) );
  nand_x1_sg U69718 ( .A(n57523), .B(n48493), .X(n38489) );
  nand_x1_sg U69719 ( .A(n57527), .B(n48491), .X(n38497) );
  nand_x1_sg U69720 ( .A(n57521), .B(n48487), .X(n38499) );
  nand_x1_sg U69721 ( .A(n57527), .B(n48485), .X(n38501) );
  nand_x1_sg U69722 ( .A(n57524), .B(n48481), .X(n38671) );
  nand_x1_sg U69723 ( .A(n57525), .B(n48479), .X(n38677) );
  nand_x1_sg U69724 ( .A(n57520), .B(n48477), .X(n38683) );
  nand_x1_sg U69725 ( .A(n57521), .B(n48467), .X(n38679) );
  nand_x1_sg U69726 ( .A(n57522), .B(n48465), .X(n38681) );
  nand_x1_sg U69727 ( .A(n57522), .B(n48463), .X(n38673) );
  nand_x1_sg U69728 ( .A(n57520), .B(n48461), .X(n38675) );
  nand_x1_sg U69729 ( .A(n57524), .B(n48451), .X(n38525) );
  nand_x1_sg U69730 ( .A(n57523), .B(n48449), .X(n38491) );
  nand_x1_sg U69731 ( .A(n57524), .B(n48447), .X(n38449) );
  nand_x1_sg U69732 ( .A(n57524), .B(n48445), .X(n38451) );
  nand_x1_sg U69733 ( .A(n57523), .B(n48443), .X(n38591) );
  nand_x1_sg U69734 ( .A(n57524), .B(n48437), .X(n38447) );
  nand_x1_sg U69735 ( .A(n57523), .B(n48419), .X(n38597) );
  nand_x1_sg U69736 ( .A(n57522), .B(n48417), .X(n38585) );
  nand_x1_sg U69737 ( .A(n57526), .B(n48415), .X(n38599) );
  nand_x1_sg U69738 ( .A(n57523), .B(n48413), .X(n38605) );
  nand_x1_sg U69739 ( .A(n57523), .B(n48411), .X(n38607) );
  nand_x1_sg U69740 ( .A(n57523), .B(n48409), .X(n38609) );
  nand_x1_sg U69741 ( .A(n57521), .B(n48407), .X(n38601) );
  nand_x1_sg U69742 ( .A(n57525), .B(n48405), .X(n38603) );
  nand_x1_sg U69743 ( .A(n57526), .B(n48403), .X(n38581) );
  nand_x1_sg U69744 ( .A(n57526), .B(n48401), .X(n38583) );
  nand_x1_sg U69745 ( .A(n57525), .B(n48399), .X(n38575) );
  nand_x1_sg U69746 ( .A(n57520), .B(n48397), .X(n38577) );
  nand_x1_sg U69747 ( .A(n57520), .B(n48395), .X(n38593) );
  nand_x1_sg U69748 ( .A(n57521), .B(n48393), .X(n38595) );
  nand_x1_sg U69749 ( .A(n57519), .B(n48391), .X(n38587) );
  nand_x1_sg U69750 ( .A(n57524), .B(n48389), .X(n38589) );
  nand_x1_sg U69751 ( .A(n57525), .B(n48387), .X(n38637) );
  nand_x1_sg U69752 ( .A(n57523), .B(n48385), .X(n38639) );
  nand_x1_sg U69753 ( .A(n57526), .B(n48383), .X(n38631) );
  nand_x1_sg U69754 ( .A(n57520), .B(n48381), .X(n38633) );
  nand_x1_sg U69755 ( .A(n57524), .B(n48379), .X(n38665) );
  nand_x1_sg U69756 ( .A(n57525), .B(n48377), .X(n38629) );
  nand_x1_sg U69757 ( .A(n57526), .B(n48375), .X(n38667) );
  nand_x1_sg U69758 ( .A(n57522), .B(n48373), .X(n38669) );
  nand_x1_sg U69759 ( .A(n57526), .B(n48371), .X(n38619) );
  nand_x1_sg U69760 ( .A(n57523), .B(n48369), .X(n38621) );
  nand_x1_sg U69761 ( .A(n57526), .B(n48367), .X(n38613) );
  nand_x1_sg U69762 ( .A(n57519), .B(n48365), .X(n38615) );
  nand_x1_sg U69763 ( .A(n57520), .B(n48363), .X(n38623) );
  nand_x1_sg U69764 ( .A(n57523), .B(n48361), .X(n38611) );
  nand_x1_sg U69765 ( .A(n57526), .B(n48359), .X(n38625) );
  nand_x1_sg U69766 ( .A(n57522), .B(n48357), .X(n38627) );
  nand_x1_sg U69767 ( .A(n57524), .B(n48351), .X(n38443) );
  nand_x1_sg U69768 ( .A(n57524), .B(n48343), .X(n38441) );
  nand_x1_sg U69769 ( .A(n57522), .B(n48341), .X(n38439) );
  nand_x1_sg U69770 ( .A(n57519), .B(n48335), .X(n38435) );
  nand_x1_sg U69771 ( .A(n57521), .B(n48333), .X(n38433) );
  nand_x1_sg U69772 ( .A(n57519), .B(n48327), .X(n38437) );
  nand_x1_sg U69773 ( .A(n57524), .B(n48303), .X(n38459) );
  nand_x1_sg U69774 ( .A(n57525), .B(n48273), .X(n38653) );
  nand_x1_sg U69775 ( .A(n57525), .B(n48265), .X(n38659) );
  nand_x1_sg U69776 ( .A(n57525), .B(n48243), .X(n38617) );
  nand_x1_sg U69777 ( .A(n57523), .B(n48219), .X(n38471) );
  nand_x1_sg U69778 ( .A(n57521), .B(n48187), .X(n38479) );
  nand_x1_sg U69779 ( .A(n57519), .B(n48185), .X(n38481) );
  nand_x1_sg U69780 ( .A(n57524), .B(n48127), .X(n38457) );
  nand_x1_sg U69781 ( .A(n57524), .B(n48125), .X(n38445) );
  nand_x1_sg U69782 ( .A(n57524), .B(n48103), .X(n38453) );
  nand_x1_sg U69783 ( .A(n57524), .B(n48101), .X(n38455) );
  nand_x1_sg U69784 ( .A(n57527), .B(n49117), .X(n39631) );
  nand_x1_sg U69785 ( .A(n57526), .B(n49115), .X(n39559) );
  nand_x1_sg U69786 ( .A(n57524), .B(n49113), .X(n39529) );
  nand_x1_sg U69787 ( .A(n57526), .B(n49111), .X(n39271) );
  nand_x1_sg U69788 ( .A(n57519), .B(n49107), .X(n39385) );
  nand_x1_sg U69789 ( .A(n57525), .B(n49105), .X(n39391) );
  nand_x1_sg U69790 ( .A(n57525), .B(n49101), .X(n39397) );
  nand_x1_sg U69791 ( .A(n57521), .B(n49099), .X(n39403) );
  nand_x1_sg U69792 ( .A(n57520), .B(n49085), .X(n39265) );
  nand_x1_sg U69793 ( .A(n57521), .B(n49075), .X(n39393) );
  nand_x1_sg U69794 ( .A(n57524), .B(n49073), .X(n39395) );
  nand_x1_sg U69795 ( .A(n57524), .B(n49071), .X(n39387) );
  nand_x1_sg U69796 ( .A(n57519), .B(n49069), .X(n39389) );
  nand_x1_sg U69797 ( .A(n57521), .B(n49067), .X(n39405) );
  nand_x1_sg U69798 ( .A(n57525), .B(n49065), .X(n39407) );
  nand_x1_sg U69799 ( .A(n57525), .B(n49063), .X(n39399) );
  nand_x1_sg U69800 ( .A(n57520), .B(n49061), .X(n39401) );
  nand_x1_sg U69801 ( .A(n57527), .B(n49059), .X(n39441) );
  nand_x1_sg U69802 ( .A(n57522), .B(n49057), .X(n39443) );
  nand_x1_sg U69803 ( .A(n57522), .B(n49055), .X(n39435) );
  nand_x1_sg U69804 ( .A(n57521), .B(n49053), .X(n39437) );
  nand_x1_sg U69805 ( .A(n57525), .B(n49051), .X(n39453) );
  nand_x1_sg U69806 ( .A(n57524), .B(n49049), .X(n39455) );
  nand_x1_sg U69807 ( .A(n57523), .B(n49047), .X(n39447) );
  nand_x1_sg U69808 ( .A(n57519), .B(n49045), .X(n39449) );
  nand_x1_sg U69809 ( .A(n57525), .B(n49043), .X(n39417) );
  nand_x1_sg U69810 ( .A(n57526), .B(n49041), .X(n39419) );
  nand_x1_sg U69811 ( .A(n57525), .B(n49039), .X(n39411) );
  nand_x1_sg U69812 ( .A(n57524), .B(n49037), .X(n39413) );
  nand_x1_sg U69813 ( .A(n57522), .B(n49035), .X(n39429) );
  nand_x1_sg U69814 ( .A(n57521), .B(n49033), .X(n39431) );
  nand_x1_sg U69815 ( .A(n57525), .B(n49031), .X(n39423) );
  nand_x1_sg U69816 ( .A(n57521), .B(n49029), .X(n39425) );
  nand_x1_sg U69817 ( .A(n57525), .B(n49027), .X(n39489) );
  nand_x1_sg U69818 ( .A(n57526), .B(n49025), .X(n39491) );
  nand_x1_sg U69819 ( .A(n57520), .B(n49023), .X(n39483) );
  nand_x1_sg U69820 ( .A(n57525), .B(n49021), .X(n39485) );
  nand_x1_sg U69821 ( .A(n57519), .B(n49019), .X(n39501) );
  nand_x1_sg U69822 ( .A(n57526), .B(n49017), .X(n39503) );
  nand_x1_sg U69823 ( .A(n57519), .B(n49015), .X(n39495) );
  nand_x1_sg U69824 ( .A(n57520), .B(n49013), .X(n39497) );
  nand_x1_sg U69825 ( .A(n57527), .B(n49011), .X(n39465) );
  nand_x1_sg U69826 ( .A(n57525), .B(n49009), .X(n39467) );
  nand_x1_sg U69827 ( .A(n57526), .B(n49007), .X(n39459) );
  nand_x1_sg U69828 ( .A(n57525), .B(n49005), .X(n39461) );
  nand_x1_sg U69829 ( .A(n57520), .B(n49003), .X(n39477) );
  nand_x1_sg U69830 ( .A(n57520), .B(n49001), .X(n39479) );
  nand_x1_sg U69831 ( .A(n57526), .B(n48999), .X(n39471) );
  nand_x1_sg U69832 ( .A(n57521), .B(n48997), .X(n39473) );
  nand_x1_sg U69833 ( .A(n57527), .B(n48995), .X(n39633) );
  nand_x1_sg U69834 ( .A(n57527), .B(n48993), .X(n39635) );
  nand_x1_sg U69835 ( .A(n57524), .B(n48991), .X(n39627) );
  nand_x1_sg U69836 ( .A(n57525), .B(n48989), .X(n39629) );
  nand_x1_sg U69837 ( .A(n57529), .B(n48987), .X(n39645) );
  nand_x1_sg U69838 ( .A(n57523), .B(n48985), .X(n39647) );
  nand_x1_sg U69839 ( .A(n57522), .B(n48983), .X(n39639) );
  nand_x1_sg U69840 ( .A(n57527), .B(n48981), .X(n39641) );
  nand_x1_sg U69841 ( .A(n57524), .B(n48979), .X(n39609) );
  nand_x1_sg U69842 ( .A(n57520), .B(n48977), .X(n39611) );
  nand_x1_sg U69843 ( .A(n57521), .B(n48975), .X(n39603) );
  nand_x1_sg U69844 ( .A(n57524), .B(n48973), .X(n39605) );
  nand_x1_sg U69845 ( .A(n57526), .B(n48971), .X(n39621) );
  nand_x1_sg U69846 ( .A(n57523), .B(n48969), .X(n39623) );
  nand_x1_sg U69847 ( .A(n57525), .B(n48967), .X(n39615) );
  nand_x1_sg U69848 ( .A(n57527), .B(n48965), .X(n39617) );
  nand_x1_sg U69849 ( .A(n57527), .B(n48963), .X(n39681) );
  nand_x1_sg U69850 ( .A(n57523), .B(n48961), .X(n39683) );
  nand_x1_sg U69851 ( .A(n57527), .B(n48959), .X(n39675) );
  nand_x1_sg U69852 ( .A(n57527), .B(n48957), .X(n39677) );
  nand_x1_sg U69853 ( .A(n57527), .B(n48955), .X(n39693) );
  nand_x1_sg U69854 ( .A(n57527), .B(n48953), .X(n39695) );
  nand_x1_sg U69855 ( .A(n57521), .B(n48951), .X(n39687) );
  nand_x1_sg U69856 ( .A(n57523), .B(n48949), .X(n39689) );
  nand_x1_sg U69857 ( .A(n57521), .B(n48947), .X(n39657) );
  nand_x1_sg U69858 ( .A(n57519), .B(n48945), .X(n39659) );
  nand_x1_sg U69859 ( .A(n57524), .B(n48943), .X(n39651) );
  nand_x1_sg U69860 ( .A(n57521), .B(n48941), .X(n39653) );
  nand_x1_sg U69861 ( .A(n57524), .B(n48939), .X(n39669) );
  nand_x1_sg U69862 ( .A(n57520), .B(n48937), .X(n39671) );
  nand_x1_sg U69863 ( .A(n57525), .B(n48935), .X(n39663) );
  nand_x1_sg U69864 ( .A(n57524), .B(n48933), .X(n39665) );
  nand_x1_sg U69865 ( .A(n57526), .B(n48931), .X(n39537) );
  nand_x1_sg U69866 ( .A(n57521), .B(n48929), .X(n39539) );
  nand_x1_sg U69867 ( .A(n57526), .B(n48927), .X(n39531) );
  nand_x1_sg U69868 ( .A(n57525), .B(n48925), .X(n39533) );
  nand_x1_sg U69869 ( .A(n57520), .B(n48923), .X(n39549) );
  nand_x1_sg U69870 ( .A(n57527), .B(n48921), .X(n39551) );
  nand_x1_sg U69871 ( .A(n57524), .B(n48919), .X(n39543) );
  nand_x1_sg U69872 ( .A(n57523), .B(n48917), .X(n39545) );
  nand_x1_sg U69873 ( .A(n57519), .B(n48915), .X(n39513) );
  nand_x1_sg U69874 ( .A(n57524), .B(n48913), .X(n39515) );
  nand_x1_sg U69875 ( .A(n57524), .B(n48911), .X(n39507) );
  nand_x1_sg U69876 ( .A(n57525), .B(n48909), .X(n39509) );
  nand_x1_sg U69877 ( .A(n57522), .B(n48907), .X(n39525) );
  nand_x1_sg U69878 ( .A(n57526), .B(n48905), .X(n39527) );
  nand_x1_sg U69879 ( .A(n57523), .B(n48903), .X(n39519) );
  nand_x1_sg U69880 ( .A(n57520), .B(n48901), .X(n39521) );
  nand_x1_sg U69881 ( .A(n57521), .B(n48899), .X(n39585) );
  nand_x1_sg U69882 ( .A(n57524), .B(n48897), .X(n39587) );
  nand_x1_sg U69883 ( .A(n57523), .B(n48895), .X(n39579) );
  nand_x1_sg U69884 ( .A(n57519), .B(n48893), .X(n39581) );
  nand_x1_sg U69885 ( .A(n57526), .B(n48891), .X(n39597) );
  nand_x1_sg U69886 ( .A(n57526), .B(n48889), .X(n39599) );
  nand_x1_sg U69887 ( .A(n57524), .B(n48887), .X(n39591) );
  nand_x1_sg U69888 ( .A(n57521), .B(n48885), .X(n39593) );
  nand_x1_sg U69889 ( .A(n57522), .B(n48883), .X(n39561) );
  nand_x1_sg U69890 ( .A(n57524), .B(n48881), .X(n39563) );
  nand_x1_sg U69891 ( .A(n57521), .B(n48879), .X(n39555) );
  nand_x1_sg U69892 ( .A(n57521), .B(n48877), .X(n39557) );
  nand_x1_sg U69893 ( .A(n57525), .B(n48875), .X(n39573) );
  nand_x1_sg U69894 ( .A(n57522), .B(n48873), .X(n39575) );
  nand_x1_sg U69895 ( .A(n57519), .B(n48871), .X(n39567) );
  nand_x1_sg U69896 ( .A(n57526), .B(n48869), .X(n39569) );
  nand_x1_sg U69897 ( .A(n57526), .B(n48739), .X(n39321) );
  nand_x1_sg U69898 ( .A(n57521), .B(n48737), .X(n39323) );
  nand_x1_sg U69899 ( .A(n57527), .B(n48735), .X(n39315) );
  nand_x1_sg U69900 ( .A(n57526), .B(n48733), .X(n39317) );
  nand_x1_sg U69901 ( .A(n57527), .B(n48731), .X(n39333) );
  nand_x1_sg U69902 ( .A(n57520), .B(n48729), .X(n39335) );
  nand_x1_sg U69903 ( .A(n57525), .B(n48727), .X(n39327) );
  nand_x1_sg U69904 ( .A(n57526), .B(n48725), .X(n39329) );
  nand_x1_sg U69905 ( .A(n57522), .B(n48723), .X(n39297) );
  nand_x1_sg U69906 ( .A(n57523), .B(n48721), .X(n39299) );
  nand_x1_sg U69907 ( .A(n57522), .B(n48719), .X(n39291) );
  nand_x1_sg U69908 ( .A(n57523), .B(n48717), .X(n39293) );
  nand_x1_sg U69909 ( .A(n57521), .B(n48715), .X(n39309) );
  nand_x1_sg U69910 ( .A(n57524), .B(n48713), .X(n39311) );
  nand_x1_sg U69911 ( .A(n57526), .B(n48711), .X(n39303) );
  nand_x1_sg U69912 ( .A(n57527), .B(n48709), .X(n39305) );
  nand_x1_sg U69913 ( .A(n57524), .B(n48707), .X(n39369) );
  nand_x1_sg U69914 ( .A(n57519), .B(n48705), .X(n39371) );
  nand_x1_sg U69915 ( .A(n57525), .B(n48703), .X(n39363) );
  nand_x1_sg U69916 ( .A(n57521), .B(n48701), .X(n39365) );
  nand_x1_sg U69917 ( .A(n57521), .B(n48699), .X(n39381) );
  nand_x1_sg U69918 ( .A(n57522), .B(n48697), .X(n39383) );
  nand_x1_sg U69919 ( .A(n57526), .B(n48695), .X(n39375) );
  nand_x1_sg U69920 ( .A(n57525), .B(n48693), .X(n39377) );
  nand_x1_sg U69921 ( .A(n57519), .B(n48691), .X(n39345) );
  nand_x1_sg U69922 ( .A(n57526), .B(n48689), .X(n39347) );
  nand_x1_sg U69923 ( .A(n57527), .B(n48687), .X(n39339) );
  nand_x1_sg U69924 ( .A(n57525), .B(n48685), .X(n39341) );
  nand_x1_sg U69925 ( .A(n57526), .B(n48683), .X(n39357) );
  nand_x1_sg U69926 ( .A(n57526), .B(n48681), .X(n39359) );
  nand_x1_sg U69927 ( .A(n57523), .B(n48679), .X(n39351) );
  nand_x1_sg U69928 ( .A(n57526), .B(n48677), .X(n39353) );
  nand_x1_sg U69929 ( .A(n57525), .B(n48643), .X(n39273) );
  nand_x1_sg U69930 ( .A(n57527), .B(n48641), .X(n39275) );
  nand_x1_sg U69931 ( .A(n57520), .B(n48639), .X(n39267) );
  nand_x1_sg U69932 ( .A(n57520), .B(n48637), .X(n39269) );
  nand_x1_sg U69933 ( .A(n57526), .B(n48635), .X(n39285) );
  nand_x1_sg U69934 ( .A(n57523), .B(n48633), .X(n39287) );
  nand_x1_sg U69935 ( .A(n57523), .B(n48631), .X(n39279) );
  nand_x1_sg U69936 ( .A(n57525), .B(n48629), .X(n39281) );
  nand_x1_sg U69937 ( .A(n57520), .B(n48619), .X(n39261) );
  nand_x1_sg U69938 ( .A(n57520), .B(n48617), .X(n39263) );
  nand_x1_sg U69939 ( .A(n57527), .B(n48547), .X(n39673) );
  nand_x1_sg U69940 ( .A(n57519), .B(n48545), .X(n39679) );
  nand_x1_sg U69941 ( .A(n57521), .B(n48539), .X(n39601) );
  nand_x1_sg U69942 ( .A(n57525), .B(n48537), .X(n39691) );
  nand_x1_sg U69943 ( .A(n57521), .B(n48535), .X(n39685) );
  nand_x1_sg U69944 ( .A(n57525), .B(n48533), .X(n39325) );
  nand_x1_sg U69945 ( .A(n57525), .B(n48527), .X(n39577) );
  nand_x1_sg U69946 ( .A(n57521), .B(n48521), .X(n39331) );
  nand_x1_sg U69947 ( .A(n57526), .B(n48489), .X(n39355) );
  nand_x1_sg U69948 ( .A(n57522), .B(n48353), .X(n39319) );
  nand_x1_sg U69949 ( .A(n57526), .B(n48349), .X(n39313) );
  nand_x1_sg U69950 ( .A(n57525), .B(n48347), .X(n39373) );
  nand_x1_sg U69951 ( .A(n57525), .B(n48345), .X(n39409) );
  nand_x1_sg U69952 ( .A(n57527), .B(n48339), .X(n39301) );
  nand_x1_sg U69953 ( .A(n57526), .B(n48337), .X(n39307) );
  nand_x1_sg U69954 ( .A(n57522), .B(n48331), .X(n39295) );
  nand_x1_sg U69955 ( .A(n57527), .B(n48325), .X(n39289) );
  nand_x1_sg U69956 ( .A(n57526), .B(n48323), .X(n39439) );
  nand_x1_sg U69957 ( .A(n57523), .B(n48321), .X(n39445) );
  nand_x1_sg U69958 ( .A(n57523), .B(n48319), .X(n39493) );
  nand_x1_sg U69959 ( .A(n57520), .B(n48317), .X(n39499) );
  nand_x1_sg U69960 ( .A(n57523), .B(n48315), .X(n39451) );
  nand_x1_sg U69961 ( .A(n57521), .B(n48313), .X(n39433) );
  nand_x1_sg U69962 ( .A(n57520), .B(n48311), .X(n39505) );
  nand_x1_sg U69963 ( .A(n57527), .B(n48309), .X(n39481) );
  nand_x1_sg U69964 ( .A(n57522), .B(n48307), .X(n39343) );
  nand_x1_sg U69965 ( .A(n57524), .B(n48305), .X(n39415) );
  nand_x1_sg U69966 ( .A(n57527), .B(n48301), .X(n39337) );
  nand_x1_sg U69967 ( .A(n57526), .B(n48299), .X(n39517) );
  nand_x1_sg U69968 ( .A(n57525), .B(n48297), .X(n39523) );
  nand_x1_sg U69969 ( .A(n57525), .B(n48295), .X(n39511) );
  nand_x1_sg U69970 ( .A(n57524), .B(n48293), .X(n39421) );
  nand_x1_sg U69971 ( .A(n57526), .B(n48275), .X(n39643) );
  nand_x1_sg U69972 ( .A(n57526), .B(n48267), .X(n39637) );
  nand_x1_sg U69973 ( .A(n57526), .B(n48261), .X(n39625) );
  nand_x1_sg U69974 ( .A(n57523), .B(n48195), .X(n39361) );
  nand_x1_sg U69975 ( .A(n57524), .B(n48193), .X(n39367) );
  nand_x1_sg U69976 ( .A(n57520), .B(n48191), .X(n39379) );
  nand_x1_sg U69977 ( .A(n57519), .B(n48189), .X(n39457) );
  nand_x1_sg U69978 ( .A(n57526), .B(n48181), .X(n39349) );
  nand_x1_sg U69979 ( .A(n57519), .B(n48177), .X(n39547) );
  nand_x1_sg U69980 ( .A(n57519), .B(n48171), .X(n39463) );
  nand_x1_sg U69981 ( .A(n57524), .B(n48169), .X(n39469) );
  nand_x1_sg U69982 ( .A(n57519), .B(n48167), .X(n39475) );
  nand_x1_sg U69983 ( .A(n57524), .B(n48165), .X(n39541) );
  nand_x1_sg U69984 ( .A(n57522), .B(n48163), .X(n39649) );
  nand_x1_sg U69985 ( .A(n57527), .B(n48161), .X(n39655) );
  nand_x1_sg U69986 ( .A(n57525), .B(n48159), .X(n39661) );
  nand_x1_sg U69987 ( .A(n57526), .B(n48157), .X(n39667) );
  nand_x1_sg U69988 ( .A(n57523), .B(n48155), .X(n39583) );
  nand_x1_sg U69989 ( .A(n57524), .B(n48153), .X(n39589) );
  nand_x1_sg U69990 ( .A(n57520), .B(n48151), .X(n39607) );
  nand_x1_sg U69991 ( .A(n57520), .B(n48149), .X(n39613) );
  nand_x1_sg U69992 ( .A(n57524), .B(n48147), .X(n39535) );
  nand_x1_sg U69993 ( .A(n57524), .B(n48145), .X(n39553) );
  nand_x1_sg U69994 ( .A(n57527), .B(n48143), .X(n39565) );
  nand_x1_sg U69995 ( .A(n57520), .B(n48141), .X(n39571) );
  nand_x1_sg U69996 ( .A(n57527), .B(n48137), .X(n39277) );
  nand_x1_sg U69997 ( .A(n57522), .B(n48135), .X(n39427) );
  nand_x1_sg U69998 ( .A(n57525), .B(n48133), .X(n39487) );
  nand_x1_sg U69999 ( .A(n57525), .B(n48115), .X(n39619) );
  nand_x1_sg U70000 ( .A(n57524), .B(n48113), .X(n39595) );
  nand_x1_sg U70001 ( .A(n57523), .B(n48109), .X(n39283) );
  nand_x1_sg U70002 ( .A(n57519), .B(n47839), .X(n39706) );
  nand_x1_sg U70003 ( .A(n57524), .B(n51623), .X(n39708) );
  nand_x1_sg U70004 ( .A(n57524), .B(n51621), .X(n39710) );
  nand_x1_sg U70005 ( .A(n57521), .B(n51619), .X(n39712) );
  nand_x1_sg U70006 ( .A(n57519), .B(n47837), .X(n39714) );
  nand_x1_sg U70007 ( .A(n57525), .B(n47835), .X(n39716) );
  nand_x1_sg U70008 ( .A(n57523), .B(n51617), .X(n39718) );
  nand_x1_sg U70009 ( .A(n57519), .B(n51615), .X(n39720) );
  nand_x1_sg U70010 ( .A(n57521), .B(n51613), .X(n39722) );
  nand_x1_sg U70011 ( .A(n57523), .B(n51611), .X(n39724) );
  nand_x1_sg U70012 ( .A(n57527), .B(n51609), .X(n39726) );
  nand_x1_sg U70013 ( .A(n57524), .B(n51607), .X(n39728) );
  nand_x1_sg U70014 ( .A(n57525), .B(n51605), .X(n39730) );
  nand_x1_sg U70015 ( .A(n57523), .B(n51603), .X(n39732) );
  nand_x1_sg U70016 ( .A(n57527), .B(n51601), .X(n39734) );
  nand_x1_sg U70017 ( .A(n57527), .B(n51599), .X(n39736) );
  nand_x1_sg U70018 ( .A(n57520), .B(n51597), .X(n39738) );
  nand_x1_sg U70019 ( .A(n57526), .B(n47833), .X(n39740) );
  nand_x1_sg U70020 ( .A(n57525), .B(n51595), .X(n39742) );
  nand_x1_sg U70021 ( .A(n57525), .B(n51593), .X(n39744) );
  nand_x1_sg U70022 ( .A(n57527), .B(n51591), .X(n39746) );
  nand_x1_sg U70023 ( .A(n57522), .B(n51589), .X(n39748) );
  nand_x1_sg U70024 ( .A(n57524), .B(n51587), .X(n39750) );
  nand_x1_sg U70025 ( .A(n57520), .B(n51585), .X(n39752) );
  nand_x1_sg U70026 ( .A(n57522), .B(n51583), .X(n39754) );
  nand_x1_sg U70027 ( .A(n57527), .B(n51581), .X(n39756) );
  nand_x1_sg U70028 ( .A(n57527), .B(n51579), .X(n39758) );
  nand_x1_sg U70029 ( .A(n57523), .B(n51577), .X(n39760) );
  nand_x1_sg U70030 ( .A(n57520), .B(n47831), .X(n39762) );
  nand_x1_sg U70031 ( .A(n57519), .B(n47829), .X(n39764) );
  nand_x1_sg U70032 ( .A(n57521), .B(n47827), .X(n39766) );
  nand_x1_sg U70033 ( .A(n57522), .B(n47825), .X(n39768) );
  nand_x1_sg U70034 ( .A(n57522), .B(n51575), .X(n39770) );
  nand_x1_sg U70035 ( .A(n57525), .B(n47823), .X(n39772) );
  nand_x1_sg U70036 ( .A(n57526), .B(n47821), .X(n39774) );
  nand_x1_sg U70037 ( .A(n57525), .B(n47819), .X(n39776) );
  nand_x1_sg U70038 ( .A(n57525), .B(n51573), .X(n39778) );
  nand_x1_sg U70039 ( .A(n57525), .B(n51571), .X(n39780) );
  nand_x1_sg U70040 ( .A(n57527), .B(n47817), .X(n39782) );
  nand_x1_sg U70041 ( .A(n57526), .B(n47815), .X(n39784) );
  nand_x1_sg U70042 ( .A(n57519), .B(n47813), .X(n39786) );
  nand_x1_sg U70043 ( .A(n57524), .B(n47811), .X(n39788) );
  nand_x1_sg U70044 ( .A(n57523), .B(n47809), .X(n39790) );
  nand_x1_sg U70045 ( .A(n57521), .B(n47807), .X(n39792) );
  nand_x1_sg U70046 ( .A(n57520), .B(n47805), .X(n39794) );
  nand_x1_sg U70047 ( .A(n57525), .B(n47803), .X(n39796) );
  nand_x1_sg U70048 ( .A(n57522), .B(n47801), .X(n39798) );
  nand_x1_sg U70049 ( .A(n57526), .B(n47799), .X(n39800) );
  nand_x1_sg U70050 ( .A(n57519), .B(n47797), .X(n39802) );
  nand_x1_sg U70051 ( .A(n57519), .B(n51569), .X(n39804) );
  nand_x1_sg U70052 ( .A(n57519), .B(n47795), .X(n39806) );
  nand_x1_sg U70053 ( .A(n57519), .B(n47793), .X(n39808) );
  nand_x1_sg U70054 ( .A(n57521), .B(n48291), .X(n38431) );
  nand_x1_sg U70055 ( .A(n57523), .B(n48287), .X(n38427) );
  nand_x1_sg U70056 ( .A(n57524), .B(n48279), .X(n38429) );
  nand_x1_sg U70057 ( .A(n57522), .B(n48271), .X(n38423) );
  nand_x1_sg U70058 ( .A(n57519), .B(n48269), .X(n38421) );
  nand_x1_sg U70059 ( .A(n57527), .B(n48263), .X(n38425) );
  nand_x1_sg U70060 ( .A(n57519), .B(n48255), .X(n38419) );
  nand_x1_sg U70061 ( .A(n57526), .B(n48179), .X(n38417) );
  nand_x1_sg U70062 ( .A(n57519), .B(n51565), .X(n39828) );
  nand_x1_sg U70063 ( .A(n57527), .B(n51563), .X(n39830) );
  nand_x1_sg U70064 ( .A(n57527), .B(n51561), .X(n39832) );
  nand_x1_sg U70065 ( .A(input_taken), .B(n57527), .X(n39834) );
  nand_x1_sg U70066 ( .A(n68240), .B(n51133), .X(n35534) );
  nand_x1_sg U70067 ( .A(o_mask[31]), .B(n57790), .X(n35533) );
  nand_x1_sg U70068 ( .A(n68241), .B(n51131), .X(n35527) );
  nand_x1_sg U70069 ( .A(o_mask[30]), .B(n57791), .X(n35526) );
  nand_x1_sg U70070 ( .A(n68237), .B(n51129), .X(n35520) );
  nand_x1_sg U70071 ( .A(o_mask[29]), .B(n57791), .X(n35519) );
  nand_x1_sg U70072 ( .A(n68238), .B(n51127), .X(n35512) );
  nand_x1_sg U70073 ( .A(o_mask[28]), .B(n57791), .X(n35511) );
  nand_x1_sg U70074 ( .A(n68251), .B(n51113), .X(n35642) );
  nand_x1_sg U70075 ( .A(o_mask[25]), .B(n57788), .X(n35641) );
  nand_x1_sg U70076 ( .A(n68252), .B(n51111), .X(n35636) );
  nand_x1_sg U70077 ( .A(o_mask[24]), .B(n57788), .X(n35635) );
  nand_x1_sg U70078 ( .A(n68234), .B(n51125), .X(n35587) );
  nand_x1_sg U70079 ( .A(o_mask[17]), .B(n57789), .X(n35586) );
  nand_x1_sg U70080 ( .A(n68250), .B(n51095), .X(n35648) );
  nand_x1_sg U70081 ( .A(o_mask[15]), .B(n57788), .X(n35647) );
  nand_x1_sg U70082 ( .A(n68254), .B(n51093), .X(n35624) );
  nand_x1_sg U70083 ( .A(o_mask[14]), .B(n57789), .X(n35623) );
  nand_x1_sg U70084 ( .A(n68258), .B(n51091), .X(n35600) );
  nand_x1_sg U70085 ( .A(o_mask[13]), .B(n57790), .X(n35599) );
  nand_x1_sg U70086 ( .A(n68259), .B(n51089), .X(n35594) );
  nand_x1_sg U70087 ( .A(o_mask[12]), .B(n57791), .X(n35593) );
  nand_x1_sg U70088 ( .A(n68257), .B(n51087), .X(n35606) );
  nand_x1_sg U70089 ( .A(o_mask[11]), .B(n57791), .X(n35605) );
  nand_x1_sg U70090 ( .A(n68256), .B(n51085), .X(n35612) );
  nand_x1_sg U70091 ( .A(o_mask[10]), .B(n57788), .X(n35611) );
  nand_x1_sg U70092 ( .A(n68253), .B(n51083), .X(n35630) );
  nand_x1_sg U70093 ( .A(o_mask[9]), .B(n57789), .X(n35629) );
  nand_x1_sg U70094 ( .A(n68255), .B(n51081), .X(n35618) );
  nand_x1_sg U70095 ( .A(o_mask[8]), .B(n57789), .X(n35617) );
  nand_x1_sg U70096 ( .A(n68260), .B(n51079), .X(n35581) );
  nand_x1_sg U70097 ( .A(o_mask[7]), .B(n57791), .X(n35580) );
  nand_x1_sg U70098 ( .A(n68261), .B(n51077), .X(n35575) );
  nand_x1_sg U70099 ( .A(o_mask[6]), .B(n57788), .X(n35574) );
  nand_x1_sg U70100 ( .A(n68245), .B(n51123), .X(n35556) );
  nand_x1_sg U70101 ( .A(o_mask[5]), .B(n57789), .X(n35555) );
  nand_x1_sg U70102 ( .A(n68246), .B(n51121), .X(n35548) );
  nand_x1_sg U70103 ( .A(o_mask[4]), .B(n57790), .X(n35547) );
  nand_x1_sg U70104 ( .A(n68263), .B(n51075), .X(n35563) );
  nand_x1_sg U70105 ( .A(o_mask[3]), .B(n57790), .X(n35562) );
  nand_x1_sg U70106 ( .A(n68262), .B(n51073), .X(n35569) );
  nand_x1_sg U70107 ( .A(o_mask[2]), .B(n57789), .X(n35568) );
  nand_x1_sg U70108 ( .A(n68249), .B(n51119), .X(n35541) );
  nand_x1_sg U70109 ( .A(o_mask[0]), .B(n57790), .X(n35540) );
  nand_x1_sg U70110 ( .A(n51133), .B(n57786), .X(n35584) );
  nand_x1_sg U70111 ( .A(n55151), .B(n57788), .X(n35585) );
  nand_x1_sg U70112 ( .A(n51131), .B(n57786), .X(n35582) );
  nand_x1_sg U70113 ( .A(n55149), .B(n57789), .X(n35583) );
  nand_x1_sg U70114 ( .A(n51129), .B(n57786), .X(n35591) );
  nand_x1_sg U70115 ( .A(n55147), .B(n57789), .X(n35592) );
  nand_x1_sg U70116 ( .A(n51127), .B(n57786), .X(n35589) );
  nand_x1_sg U70117 ( .A(n55145), .B(n57790), .X(n35590) );
  nand_x1_sg U70118 ( .A(n55219), .B(n57791), .X(n35573) );
  nand_x1_sg U70119 ( .A(n55217), .B(n57788), .X(n35571) );
  nand_x1_sg U70120 ( .A(n55215), .B(n57791), .X(n35579) );
  nand_x1_sg U70121 ( .A(n55213), .B(n57788), .X(n35577) );
  nand_x1_sg U70122 ( .A(n55211), .B(n57788), .X(n35610) );
  nand_x1_sg U70123 ( .A(n55209), .B(n57789), .X(n35608) );
  nand_x1_sg U70124 ( .A(n55207), .B(n57789), .X(n35616) );
  nand_x1_sg U70125 ( .A(n55205), .B(n57789), .X(n35614) );
  nand_x1_sg U70126 ( .A(n55203), .B(n57790), .X(n35598) );
  nand_x1_sg U70127 ( .A(n55201), .B(n57791), .X(n35596) );
  nand_x1_sg U70128 ( .A(n51125), .B(n57786), .X(n35603) );
  nand_x1_sg U70129 ( .A(n55143), .B(n57789), .X(n35604) );
  nand_x1_sg U70130 ( .A(n55199), .B(n57789), .X(n35602) );
  nand_x1_sg U70131 ( .A(n55197), .B(n57790), .X(n35532) );
  nand_x1_sg U70132 ( .A(n55195), .B(n57791), .X(n35530) );
  nand_x1_sg U70133 ( .A(n55193), .B(n57790), .X(n35539) );
  nand_x1_sg U70134 ( .A(n55191), .B(n57790), .X(n35537) );
  nand_x1_sg U70135 ( .A(n55189), .B(n57791), .X(n35518) );
  nand_x1_sg U70136 ( .A(n55187), .B(n57791), .X(n35516) );
  nand_x1_sg U70137 ( .A(n55185), .B(n57791), .X(n35525) );
  nand_x1_sg U70138 ( .A(n55183), .B(n57791), .X(n35523) );
  nand_x1_sg U70139 ( .A(n55181), .B(n57790), .X(n35561) );
  nand_x1_sg U70140 ( .A(n55179), .B(n57791), .X(n35559) );
  nand_x1_sg U70141 ( .A(n51123), .B(n57786), .X(n35566) );
  nand_x1_sg U70142 ( .A(n55141), .B(n57790), .X(n35567) );
  nand_x1_sg U70143 ( .A(n51121), .B(n57786), .X(n35564) );
  nand_x1_sg U70144 ( .A(n55139), .B(n57791), .X(n35565) );
  nand_x1_sg U70145 ( .A(n55177), .B(n57790), .X(n35546) );
  nand_x1_sg U70146 ( .A(n55175), .B(n57790), .X(n35544) );
  nand_x1_sg U70147 ( .A(n55173), .B(n57788), .X(n35554) );
  nand_x1_sg U70148 ( .A(n51119), .B(n57786), .X(n35550) );
  nand_x1_sg U70149 ( .A(n55137), .B(n57791), .X(n35551) );
  nand_x1_sg U70150 ( .A(n51095), .B(n57786), .X(n35633) );
  nand_x1_sg U70151 ( .A(n55113), .B(n57788), .X(n35634) );
  nand_x1_sg U70152 ( .A(n51093), .B(n57786), .X(n35631) );
  nand_x1_sg U70153 ( .A(n55111), .B(n57789), .X(n35632) );
  nand_x1_sg U70154 ( .A(n51091), .B(n57786), .X(n35639) );
  nand_x1_sg U70155 ( .A(n55109), .B(n57788), .X(n35640) );
  nand_x1_sg U70156 ( .A(n51089), .B(n57786), .X(n35637) );
  nand_x1_sg U70157 ( .A(n55107), .B(n57788), .X(n35638) );
  nand_x1_sg U70158 ( .A(n51087), .B(n57786), .X(n35621) );
  nand_x1_sg U70159 ( .A(n55105), .B(n57789), .X(n35622) );
  nand_x1_sg U70160 ( .A(n51085), .B(n57786), .X(n35619) );
  nand_x1_sg U70161 ( .A(n55103), .B(n57789), .X(n35620) );
  nand_x1_sg U70162 ( .A(n51083), .B(n57786), .X(n35627) );
  nand_x1_sg U70163 ( .A(n55101), .B(n57789), .X(n35628) );
  nand_x1_sg U70164 ( .A(n51081), .B(n57786), .X(n35625) );
  nand_x1_sg U70165 ( .A(n55099), .B(n57789), .X(n35626) );
  nand_x1_sg U70166 ( .A(n51075), .B(n57786), .X(n35645) );
  nand_x1_sg U70167 ( .A(n55093), .B(n57788), .X(n35646) );
  nand_x1_sg U70168 ( .A(n51073), .B(n57786), .X(n35643) );
  nand_x1_sg U70169 ( .A(n55091), .B(n57788), .X(n35644) );
  nand_x1_sg U70170 ( .A(n68232), .B(n51117), .X(n35700) );
  nand_x1_sg U70171 ( .A(o_mask[27]), .B(n57790), .X(n35699) );
  nand_x1_sg U70172 ( .A(n68233), .B(n51115), .X(n35694) );
  nand_x1_sg U70173 ( .A(o_mask[26]), .B(n57791), .X(n35693) );
  nand_x1_sg U70174 ( .A(n68239), .B(n51109), .X(n35679) );
  nand_x1_sg U70175 ( .A(o_mask[23]), .B(n57793), .X(n35678) );
  nand_x1_sg U70176 ( .A(n68242), .B(n51107), .X(n35675) );
  nand_x1_sg U70177 ( .A(o_mask[22]), .B(n57788), .X(n35674) );
  nand_x1_sg U70178 ( .A(n68247), .B(n51105), .X(n35659) );
  nand_x1_sg U70179 ( .A(o_mask[21]), .B(n57788), .X(n35658) );
  nand_x1_sg U70180 ( .A(n68248), .B(n51103), .X(n35653) );
  nand_x1_sg U70181 ( .A(o_mask[20]), .B(n57789), .X(n35652) );
  nand_x1_sg U70182 ( .A(n68244), .B(n51101), .X(n35663) );
  nand_x1_sg U70183 ( .A(o_mask[19]), .B(n57790), .X(n35662) );
  nand_x1_sg U70184 ( .A(n68243), .B(n51099), .X(n35669) );
  nand_x1_sg U70185 ( .A(o_mask[18]), .B(n57788), .X(n35668) );
  nand_x1_sg U70186 ( .A(n68236), .B(n51097), .X(n35683) );
  nand_x1_sg U70187 ( .A(o_mask[16]), .B(n57789), .X(n35682) );
  nand_x1_sg U70188 ( .A(n68235), .B(n51071), .X(n35689) );
  nand_x1_sg U70189 ( .A(o_mask[1]), .B(n57790), .X(n35688) );
  nand_x1_sg U70190 ( .A(n55171), .B(n57790), .X(n35677) );
  nand_x1_sg U70191 ( .A(n55169), .B(n57791), .X(n35676) );
  nand_x1_sg U70192 ( .A(n55167), .B(n57791), .X(n35681) );
  nand_x1_sg U70193 ( .A(n55165), .B(n57790), .X(n35680) );
  nand_x1_sg U70194 ( .A(n51117), .B(n57786), .X(n35666) );
  nand_x1_sg U70195 ( .A(n55135), .B(n57791), .X(n35667) );
  nand_x1_sg U70196 ( .A(n51115), .B(n57786), .X(n35664) );
  nand_x1_sg U70197 ( .A(n55133), .B(n57788), .X(n35665) );
  nand_x1_sg U70198 ( .A(n51113), .B(n57786), .X(n35672) );
  nand_x1_sg U70199 ( .A(n55131), .B(n57788), .X(n35673) );
  nand_x1_sg U70200 ( .A(n51111), .B(n57786), .X(n35670) );
  nand_x1_sg U70201 ( .A(n55129), .B(n57790), .X(n35671) );
  nand_x1_sg U70202 ( .A(n51109), .B(n57786), .X(n35697) );
  nand_x1_sg U70203 ( .A(n55127), .B(n57790), .X(n35698) );
  nand_x1_sg U70204 ( .A(n51107), .B(n57786), .X(n35695) );
  nand_x1_sg U70205 ( .A(n55125), .B(n57791), .X(n35696) );
  nand_x1_sg U70206 ( .A(n51105), .B(n57786), .X(n35703) );
  nand_x1_sg U70207 ( .A(n55123), .B(n57791), .X(n35704) );
  nand_x1_sg U70208 ( .A(n51103), .B(n57786), .X(n35701) );
  nand_x1_sg U70209 ( .A(n55121), .B(n57789), .X(n35702) );
  nand_x1_sg U70210 ( .A(n51101), .B(n57786), .X(n35686) );
  nand_x1_sg U70211 ( .A(n55119), .B(n57788), .X(n35687) );
  nand_x1_sg U70212 ( .A(n51099), .B(n57786), .X(n35684) );
  nand_x1_sg U70213 ( .A(n55117), .B(n57789), .X(n35685) );
  nand_x1_sg U70214 ( .A(n55163), .B(n57789), .X(n35692) );
  nand_x1_sg U70215 ( .A(n51097), .B(n57786), .X(n35690) );
  nand_x1_sg U70216 ( .A(n55115), .B(n57790), .X(n35691) );
  nand_x1_sg U70217 ( .A(n51079), .B(n57786), .X(n35656) );
  nand_x1_sg U70218 ( .A(n55097), .B(n57788), .X(n35657) );
  nand_x1_sg U70219 ( .A(n51077), .B(n57786), .X(n35654) );
  nand_x1_sg U70220 ( .A(n55095), .B(n57791), .X(n35655) );
  nand_x1_sg U70221 ( .A(n55161), .B(n57789), .X(n35661) );
  nand_x1_sg U70222 ( .A(n55159), .B(n57790), .X(n35660) );
  nand_x1_sg U70223 ( .A(n51071), .B(n57786), .X(n35650) );
  nand_x1_sg U70224 ( .A(n55089), .B(n57790), .X(n35651) );
  nand_x1_sg U70225 ( .A(n55157), .B(n57788), .X(n35649) );
  nand_x1_sg U70226 ( .A(n61907), .B(n61905), .X(n32484) );
  nand_x1_sg U70227 ( .A(n68372), .B(n47337), .X(n35841) );
  nor_x1_sg U70228 ( .A(n57065), .B(n32560), .X(n32559) );
  nand_x2_sg U70229 ( .A(n32547), .B(n32548), .X(n32546) );
  nor_x1_sg U70230 ( .A(n47763), .B(n57055), .X(n32547) );
  nor_x1_sg U70231 ( .A(n51527), .B(n32549), .X(n32548) );
  nand_x2_sg U70232 ( .A(n32550), .B(n32551), .X(n32545) );
  nor_x1_sg U70233 ( .A(n51529), .B(n47765), .X(n32550) );
  nor_x1_sg U70234 ( .A(n57049), .B(n32552), .X(n32551) );
  nand_x2_sg U70235 ( .A(n32555), .B(n32556), .X(n32554) );
  nor_x1_sg U70236 ( .A(n51531), .B(n47761), .X(n32555) );
  nor_x1_sg U70237 ( .A(n57051), .B(n32557), .X(n32556) );
  nor_x1_sg U70238 ( .A(n57067), .B(n32115), .X(n32114) );
  nand_x2_sg U70239 ( .A(n32102), .B(n32103), .X(n32101) );
  nor_x1_sg U70240 ( .A(n47769), .B(n57063), .X(n32102) );
  nor_x1_sg U70241 ( .A(n51535), .B(n32104), .X(n32103) );
  nand_x2_sg U70242 ( .A(n32105), .B(n32106), .X(n32100) );
  nor_x1_sg U70243 ( .A(n51537), .B(n47771), .X(n32105) );
  nor_x1_sg U70244 ( .A(n57057), .B(n32107), .X(n32106) );
  nand_x2_sg U70245 ( .A(n32110), .B(n32111), .X(n32109) );
  nor_x1_sg U70246 ( .A(n51539), .B(n47767), .X(n32110) );
  nor_x1_sg U70247 ( .A(n57059), .B(n32112), .X(n32111) );
  nor_x1_sg U70248 ( .A(n51493), .B(n57015), .X(n32283) );
  nor_x1_sg U70249 ( .A(n51515), .B(n57039), .X(n32286) );
  nor_x1_sg U70250 ( .A(n51517), .B(n57041), .X(n32291) );
  nor_x1_sg U70251 ( .A(n51519), .B(n57043), .X(n32294) );
  nor_x1_sg U70252 ( .A(n51507), .B(n57031), .X(n32728) );
  nor_x1_sg U70253 ( .A(n51509), .B(n57033), .X(n32731) );
  nor_x1_sg U70254 ( .A(n51511), .B(n57035), .X(n32736) );
  nor_x1_sg U70255 ( .A(n51513), .B(n57037), .X(n32739) );
  nand_x2_sg U70256 ( .A(n32281), .B(n32282), .X(n32280) );
  nor_x1_sg U70257 ( .A(n47745), .B(n57029), .X(n32281) );
  nor_x1_sg U70258 ( .A(n51489), .B(n68537), .X(n32282) );
  nand_x2_sg U70259 ( .A(n32284), .B(n32285), .X(n32279) );
  nor_x1_sg U70260 ( .A(n51491), .B(n47747), .X(n32284) );
  nor_x1_sg U70261 ( .A(n57013), .B(n68538), .X(n32285) );
  nand_x2_sg U70262 ( .A(n32289), .B(n32290), .X(n32288) );
  nor_x1_sg U70263 ( .A(n51503), .B(n47743), .X(n32289) );
  nor_x1_sg U70264 ( .A(n57021), .B(n68539), .X(n32290) );
  nand_x2_sg U70265 ( .A(n32292), .B(n32293), .X(n32287) );
  nor_x1_sg U70266 ( .A(n51505), .B(n47757), .X(n32292) );
  nor_x1_sg U70267 ( .A(n57027), .B(n68540), .X(n32293) );
  nand_x2_sg U70268 ( .A(n32726), .B(n32727), .X(n32725) );
  nor_x1_sg U70269 ( .A(n47751), .B(n57025), .X(n32726) );
  nor_x1_sg U70270 ( .A(n51495), .B(n68444), .X(n32727) );
  nand_x2_sg U70271 ( .A(n32729), .B(n32730), .X(n32724) );
  nor_x1_sg U70272 ( .A(n51497), .B(n47753), .X(n32729) );
  nor_x1_sg U70273 ( .A(n57017), .B(n68445), .X(n32730) );
  nand_x2_sg U70274 ( .A(n32734), .B(n32735), .X(n32733) );
  nor_x1_sg U70275 ( .A(n51499), .B(n47749), .X(n32734) );
  nor_x1_sg U70276 ( .A(n57019), .B(n68446), .X(n32735) );
  nand_x2_sg U70277 ( .A(n32737), .B(n32738), .X(n32732) );
  nor_x1_sg U70278 ( .A(n51501), .B(n47755), .X(n32737) );
  nor_x1_sg U70279 ( .A(n57023), .B(n68447), .X(n32738) );
  nand_x1_sg U70280 ( .A(n57069), .B(n57294), .X(n32801) );
  nand_x1_sg U70281 ( .A(n56971), .B(n57294), .X(n32815) );
  nand_x1_sg U70282 ( .A(n51523), .B(n57294), .X(n32826) );
  nand_x1_sg U70283 ( .A(n47441), .B(n57294), .X(n32822) );
  nand_x1_sg U70284 ( .A(n51561), .B(n57780), .X(n35796) );
  nand_x1_sg U70285 ( .A(n57782), .B(n51133), .X(n35797) );
  nand_x1_sg U70286 ( .A(n51563), .B(n57780), .X(n35810) );
  nand_x1_sg U70287 ( .A(n57782), .B(n51131), .X(n35811) );
  nand_x1_sg U70288 ( .A(n51565), .B(n57780), .X(n35802) );
  nand_x1_sg U70289 ( .A(n57782), .B(n51129), .X(n35803) );
  nand_x1_sg U70290 ( .A(n51567), .B(n57780), .X(n35794) );
  nand_x1_sg U70291 ( .A(n57782), .B(n51127), .X(n35795) );
  nand_x1_sg U70292 ( .A(n51569), .B(n57780), .X(n35784) );
  nand_x1_sg U70293 ( .A(n57784), .B(n51125), .X(n35785) );
  nand_x1_sg U70294 ( .A(n51571), .B(n57780), .X(n35812) );
  nand_x1_sg U70295 ( .A(n57782), .B(n51123), .X(n35813) );
  nand_x1_sg U70296 ( .A(n51573), .B(n57780), .X(n35814) );
  nand_x1_sg U70297 ( .A(n57782), .B(n51121), .X(n35815) );
  nand_x1_sg U70298 ( .A(n51575), .B(n57780), .X(n35728) );
  nand_x1_sg U70299 ( .A(n57784), .B(n51119), .X(n35729) );
  nand_x1_sg U70300 ( .A(n51577), .B(n57780), .X(n35744) );
  nand_x1_sg U70301 ( .A(n57782), .B(n51117), .X(n35745) );
  nand_x1_sg U70302 ( .A(n51579), .B(n57780), .X(n35746) );
  nand_x1_sg U70303 ( .A(n57782), .B(n51115), .X(n35747) );
  nand_x1_sg U70304 ( .A(n51581), .B(n57780), .X(n35738) );
  nand_x1_sg U70305 ( .A(n57782), .B(n51113), .X(n35739) );
  nand_x1_sg U70306 ( .A(n51583), .B(n57780), .X(n35740) );
  nand_x1_sg U70307 ( .A(n57782), .B(n51111), .X(n35741) );
  nand_x1_sg U70308 ( .A(n51585), .B(n57779), .X(n35718) );
  nand_x1_sg U70309 ( .A(n35708), .B(n51109), .X(n35719) );
  nand_x1_sg U70310 ( .A(n51587), .B(n57779), .X(n35720) );
  nand_x1_sg U70311 ( .A(n35708), .B(n51107), .X(n35721) );
  nand_x1_sg U70312 ( .A(n51589), .B(n57779), .X(n35712) );
  nand_x1_sg U70313 ( .A(n35708), .B(n51105), .X(n35713) );
  nand_x1_sg U70314 ( .A(n51591), .B(n57779), .X(n35714) );
  nand_x1_sg U70315 ( .A(n57782), .B(n51103), .X(n35715) );
  nand_x1_sg U70316 ( .A(n51593), .B(n57780), .X(n35730) );
  nand_x1_sg U70317 ( .A(n57782), .B(n51101), .X(n35731) );
  nand_x1_sg U70318 ( .A(n51595), .B(n57780), .X(n35732) );
  nand_x1_sg U70319 ( .A(n57782), .B(n51099), .X(n35733) );
  nand_x1_sg U70320 ( .A(n51597), .B(n57780), .X(n35726) );
  nand_x1_sg U70321 ( .A(n57782), .B(n51097), .X(n35727) );
  nand_x1_sg U70322 ( .A(n51599), .B(n57780), .X(n35748) );
  nand_x1_sg U70323 ( .A(n57782), .B(n51095), .X(n35749) );
  nand_x1_sg U70324 ( .A(n51601), .B(n57780), .X(n35754) );
  nand_x1_sg U70325 ( .A(n57782), .B(n51093), .X(n35755) );
  nand_x1_sg U70326 ( .A(n51603), .B(n57780), .X(n35774) );
  nand_x1_sg U70327 ( .A(n57782), .B(n51091), .X(n35775) );
  nand_x1_sg U70328 ( .A(n51605), .B(n57780), .X(n35766) );
  nand_x1_sg U70329 ( .A(n57782), .B(n51089), .X(n35767) );
  nand_x1_sg U70330 ( .A(n51607), .B(n57780), .X(n35776) );
  nand_x1_sg U70331 ( .A(n57782), .B(n51087), .X(n35777) );
  nand_x1_sg U70332 ( .A(n51609), .B(n57780), .X(n35778) );
  nand_x1_sg U70333 ( .A(n57782), .B(n51085), .X(n35779) );
  nand_x1_sg U70334 ( .A(n51611), .B(n57780), .X(n35770) );
  nand_x1_sg U70335 ( .A(n57782), .B(n51083), .X(n35771) );
  nand_x1_sg U70336 ( .A(n51613), .B(n57780), .X(n35772) );
  nand_x1_sg U70337 ( .A(n57782), .B(n51081), .X(n35773) );
  nand_x1_sg U70338 ( .A(n51615), .B(n57780), .X(n35756) );
  nand_x1_sg U70339 ( .A(n57782), .B(n51079), .X(n35757) );
  nand_x1_sg U70340 ( .A(n51617), .B(n57780), .X(n35758) );
  nand_x1_sg U70341 ( .A(n57782), .B(n51077), .X(n35759) );
  nand_x1_sg U70342 ( .A(n51619), .B(n57780), .X(n35706) );
  nand_x1_sg U70343 ( .A(n57782), .B(n51075), .X(n35707) );
  nand_x1_sg U70344 ( .A(n51621), .B(n57780), .X(n35760) );
  nand_x1_sg U70345 ( .A(n57782), .B(n51073), .X(n35761) );
  nand_x1_sg U70346 ( .A(n51623), .B(n57780), .X(n35762) );
  nand_x1_sg U70347 ( .A(n57782), .B(n51071), .X(n35763) );
  nand_x1_sg U70348 ( .A(n47373), .B(n57294), .X(n32830) );
  nand_x1_sg U70349 ( .A(n56935), .B(n57294), .X(n32811) );
  nand_x1_sg U70350 ( .A(n47777), .B(n57780), .X(n35804) );
  nand_x1_sg U70351 ( .A(n57782), .B(n53711), .X(n35805) );
  nand_x1_sg U70352 ( .A(n47779), .B(n57780), .X(n35806) );
  nand_x1_sg U70353 ( .A(n57782), .B(n53709), .X(n35807) );
  nand_x1_sg U70354 ( .A(n47781), .B(n57780), .X(n35798) );
  nand_x1_sg U70355 ( .A(n57782), .B(n53707), .X(n35799) );
  nand_x1_sg U70356 ( .A(n47783), .B(n57780), .X(n35800) );
  nand_x1_sg U70357 ( .A(n57782), .B(n53705), .X(n35801) );
  nand_x1_sg U70358 ( .A(n47785), .B(n57780), .X(n35782) );
  nand_x1_sg U70359 ( .A(n57782), .B(n53703), .X(n35783) );
  nand_x1_sg U70360 ( .A(n47787), .B(n57780), .X(n35816) );
  nand_x1_sg U70361 ( .A(n57782), .B(n53701), .X(n35817) );
  nand_x1_sg U70362 ( .A(n47789), .B(n57780), .X(n35788) );
  nand_x1_sg U70363 ( .A(n57782), .B(n53699), .X(n35789) );
  nand_x1_sg U70364 ( .A(n47791), .B(n57780), .X(n35780) );
  nand_x1_sg U70365 ( .A(n57782), .B(n53697), .X(n35781) );
  nand_x1_sg U70366 ( .A(n47793), .B(n57780), .X(n35790) );
  nand_x1_sg U70367 ( .A(n57782), .B(n53695), .X(n35791) );
  nand_x1_sg U70368 ( .A(n47795), .B(n57780), .X(n35792) );
  nand_x1_sg U70369 ( .A(n57782), .B(n53693), .X(n35793) );
  nand_x1_sg U70370 ( .A(n47797), .B(n57780), .X(n35786) );
  nand_x1_sg U70371 ( .A(n57782), .B(n53691), .X(n35787) );
  nand_x1_sg U70372 ( .A(n47799), .B(n57780), .X(n35824) );
  nand_x1_sg U70373 ( .A(n57782), .B(n53689), .X(n35825) );
  nand_x1_sg U70374 ( .A(n47801), .B(n57780), .X(n35808) );
  nand_x1_sg U70375 ( .A(n57782), .B(n53687), .X(n35809) );
  nand_x1_sg U70376 ( .A(n47803), .B(n57780), .X(n35830) );
  nand_x1_sg U70377 ( .A(n57782), .B(n53685), .X(n35831) );
  nand_x1_sg U70378 ( .A(n47805), .B(n57780), .X(n35822) );
  nand_x1_sg U70379 ( .A(n57782), .B(n53683), .X(n35823) );
  nand_x1_sg U70380 ( .A(n47807), .B(n57780), .X(n35832) );
  nand_x1_sg U70381 ( .A(n57782), .B(n53681), .X(n35833) );
  nand_x1_sg U70382 ( .A(n47809), .B(n57779), .X(n35834) );
  nand_x1_sg U70383 ( .A(n57782), .B(n53679), .X(n35835) );
  nand_x1_sg U70384 ( .A(n47811), .B(n57780), .X(n35826) );
  nand_x1_sg U70385 ( .A(n57782), .B(n53677), .X(n35827) );
  nand_x1_sg U70386 ( .A(n47813), .B(n57780), .X(n35828) );
  nand_x1_sg U70387 ( .A(n57782), .B(n53675), .X(n35829) );
  nand_x1_sg U70388 ( .A(n47815), .B(n57780), .X(n35818) );
  nand_x1_sg U70389 ( .A(n57782), .B(n53673), .X(n35819) );
  nand_x1_sg U70390 ( .A(n47817), .B(n57780), .X(n35820) );
  nand_x1_sg U70391 ( .A(n57782), .B(n53671), .X(n35821) );
  nand_x1_sg U70392 ( .A(n47819), .B(n57779), .X(n35710) );
  nand_x1_sg U70393 ( .A(n57782), .B(n53669), .X(n35711) );
  nand_x1_sg U70394 ( .A(n47821), .B(n57779), .X(n35716) );
  nand_x1_sg U70395 ( .A(n57782), .B(n53667), .X(n35717) );
  nand_x1_sg U70396 ( .A(n47823), .B(n57780), .X(n35722) );
  nand_x1_sg U70397 ( .A(n57782), .B(n53665), .X(n35723) );
  nand_x1_sg U70398 ( .A(n47825), .B(n57780), .X(n35736) );
  nand_x1_sg U70399 ( .A(n57782), .B(n53663), .X(n35737) );
  nand_x1_sg U70400 ( .A(n47827), .B(n57780), .X(n35768) );
  nand_x1_sg U70401 ( .A(n57782), .B(n53661), .X(n35769) );
  nand_x1_sg U70402 ( .A(n47829), .B(n57780), .X(n35742) );
  nand_x1_sg U70403 ( .A(n57782), .B(n53659), .X(n35743) );
  nand_x1_sg U70404 ( .A(n47831), .B(n57780), .X(n35734) );
  nand_x1_sg U70405 ( .A(n57782), .B(n53657), .X(n35735) );
  nand_x1_sg U70406 ( .A(n47833), .B(n57780), .X(n35724) );
  nand_x1_sg U70407 ( .A(n57782), .B(n53655), .X(n35725) );
  nand_x1_sg U70408 ( .A(n47835), .B(n57780), .X(n35750) );
  nand_x1_sg U70409 ( .A(n57782), .B(n53653), .X(n35751) );
  nand_x1_sg U70410 ( .A(n47837), .B(n57780), .X(n35752) );
  nand_x1_sg U70411 ( .A(n57782), .B(n53651), .X(n35753) );
  nand_x1_sg U70412 ( .A(n47839), .B(n57780), .X(n35764) );
  nand_x1_sg U70413 ( .A(n57782), .B(n53649), .X(n35765) );
  nor_x1_sg U70414 ( .A(n56865), .B(n68437), .X(n32597) );
  nor_x1_sg U70415 ( .A(n47695), .B(n51407), .X(n32598) );
  nor_x1_sg U70416 ( .A(n51331), .B(n56779), .X(n32587) );
  nor_x1_sg U70417 ( .A(n51333), .B(n56781), .X(n32590) );
  nor_x1_sg U70418 ( .A(n51335), .B(n56783), .X(n32595) );
  nand_x2_sg U70419 ( .A(n32585), .B(n32586), .X(n32584) );
  nor_x1_sg U70420 ( .A(n47675), .B(n56847), .X(n32585) );
  nor_x1_sg U70421 ( .A(n51381), .B(n68434), .X(n32586) );
  nand_x2_sg U70422 ( .A(n32588), .B(n32589), .X(n32583) );
  nor_x1_sg U70423 ( .A(n51383), .B(n47677), .X(n32588) );
  nor_x1_sg U70424 ( .A(n56825), .B(n68435), .X(n32589) );
  nand_x2_sg U70425 ( .A(n32593), .B(n32594), .X(n32592) );
  nor_x1_sg U70426 ( .A(n51385), .B(n47673), .X(n32593) );
  nor_x1_sg U70427 ( .A(n56827), .B(n68436), .X(n32594) );
  nor_x1_sg U70428 ( .A(n57053), .B(n51533), .X(n32558) );
  nor_x1_sg U70429 ( .A(n56867), .B(n68528), .X(n32152) );
  nor_x1_sg U70430 ( .A(n47697), .B(n51409), .X(n32153) );
  nor_x1_sg U70431 ( .A(n51337), .B(n56785), .X(n32142) );
  nor_x1_sg U70432 ( .A(n51339), .B(n56787), .X(n32145) );
  nor_x1_sg U70433 ( .A(n51341), .B(n56789), .X(n32150) );
  nand_x1_sg U70434 ( .A(n57091), .B(n32802), .X(n32828) );
  nand_x1_sg U70435 ( .A(n51525), .B(n57294), .X(n32813) );
  nand_x2_sg U70436 ( .A(n32140), .B(n32141), .X(n32139) );
  nor_x1_sg U70437 ( .A(n47687), .B(n56849), .X(n32140) );
  nor_x1_sg U70438 ( .A(n51395), .B(n68525), .X(n32141) );
  nand_x2_sg U70439 ( .A(n32143), .B(n32144), .X(n32138) );
  nor_x1_sg U70440 ( .A(n51397), .B(n47689), .X(n32143) );
  nor_x1_sg U70441 ( .A(n56837), .B(n68526), .X(n32144) );
  nand_x2_sg U70442 ( .A(n32148), .B(n32149), .X(n32147) );
  nor_x1_sg U70443 ( .A(n51399), .B(n47685), .X(n32148) );
  nor_x1_sg U70444 ( .A(n56839), .B(n68527), .X(n32149) );
  nor_x1_sg U70445 ( .A(n57061), .B(n51541), .X(n32113) );
  nand_x1_sg U70446 ( .A(n47443), .B(n57294), .X(n32824) );
  nand_x1_sg U70447 ( .A(n56969), .B(n57294), .X(n32817) );
  nand_x1_sg U70448 ( .A(n47375), .B(n57294), .X(n32805) );
  nor_x1_sg U70449 ( .A(n56861), .B(n68462), .X(n32719) );
  nor_x1_sg U70450 ( .A(n47701), .B(n51411), .X(n32720) );
  nor_x1_sg U70451 ( .A(n47569), .B(n68441), .X(n32577) );
  nor_x1_sg U70452 ( .A(n47733), .B(n51473), .X(n32578) );
  nor_x1_sg U70453 ( .A(n51355), .B(n56803), .X(n32709) );
  nor_x1_sg U70454 ( .A(n51357), .B(n56805), .X(n32712) );
  nor_x1_sg U70455 ( .A(n51359), .B(n56807), .X(n32717) );
  nor_x1_sg U70456 ( .A(n51475), .B(n56905), .X(n32181) );
  nor_x1_sg U70457 ( .A(n51477), .B(n56907), .X(n32184) );
  nor_x1_sg U70458 ( .A(n51479), .B(n56909), .X(n32189) );
  nor_x1_sg U70459 ( .A(n51465), .B(n56897), .X(n32626) );
  nor_x1_sg U70460 ( .A(n51467), .B(n56899), .X(n32629) );
  nor_x1_sg U70461 ( .A(n51469), .B(n56901), .X(n32634) );
  nor_x1_sg U70462 ( .A(n47739), .B(n68513), .X(n32191) );
  nor_x1_sg U70463 ( .A(n51487), .B(n56915), .X(n32192) );
  nor_x1_sg U70464 ( .A(n47737), .B(n68424), .X(n32636) );
  nor_x1_sg U70465 ( .A(n51485), .B(n56913), .X(n32637) );
  nor_x1_sg U70466 ( .A(n47715), .B(n51447), .X(n32122) );
  nor_x1_sg U70467 ( .A(n47717), .B(n51449), .X(n32125) );
  nor_x1_sg U70468 ( .A(n47719), .B(n51451), .X(n32130) );
  nor_x1_sg U70469 ( .A(n47709), .B(n51441), .X(n32567) );
  nor_x1_sg U70470 ( .A(n47711), .B(n51443), .X(n32570) );
  nor_x1_sg U70471 ( .A(n47713), .B(n51445), .X(n32575) );
  nor_x1_sg U70472 ( .A(n47571), .B(n68533), .X(n32132) );
  nor_x1_sg U70473 ( .A(n47735), .B(n51483), .X(n32133) );
  nand_x2_sg U70474 ( .A(n32707), .B(n32708), .X(n32706) );
  nor_x1_sg U70475 ( .A(n47655), .B(n56775), .X(n32707) );
  nor_x1_sg U70476 ( .A(n51291), .B(n68459), .X(n32708) );
  nand_x2_sg U70477 ( .A(n32710), .B(n32711), .X(n32705) );
  nor_x1_sg U70478 ( .A(n51293), .B(n47657), .X(n32710) );
  nor_x1_sg U70479 ( .A(n56757), .B(n68460), .X(n32711) );
  nand_x2_sg U70480 ( .A(n32715), .B(n32716), .X(n32714) );
  nor_x1_sg U70481 ( .A(n51295), .B(n47653), .X(n32715) );
  nor_x1_sg U70482 ( .A(n56759), .B(n68461), .X(n32716) );
  nand_x2_sg U70483 ( .A(n32179), .B(n32180), .X(n32178) );
  nor_x1_sg U70484 ( .A(n47729), .B(n56895), .X(n32179) );
  nor_x1_sg U70485 ( .A(n51459), .B(n68510), .X(n32180) );
  nand_x2_sg U70486 ( .A(n32182), .B(n32183), .X(n32177) );
  nor_x1_sg U70487 ( .A(n51461), .B(n47731), .X(n32182) );
  nor_x1_sg U70488 ( .A(n56891), .B(n68511), .X(n32183) );
  nand_x2_sg U70489 ( .A(n32187), .B(n32188), .X(n32186) );
  nor_x1_sg U70490 ( .A(n51463), .B(n47727), .X(n32187) );
  nor_x1_sg U70491 ( .A(n56893), .B(n68512), .X(n32188) );
  nand_x2_sg U70492 ( .A(n32624), .B(n32625), .X(n32623) );
  nor_x1_sg U70493 ( .A(n47723), .B(n56889), .X(n32624) );
  nor_x1_sg U70494 ( .A(n51453), .B(n68421), .X(n32625) );
  nand_x2_sg U70495 ( .A(n32627), .B(n32628), .X(n32622) );
  nor_x1_sg U70496 ( .A(n51455), .B(n47725), .X(n32627) );
  nor_x1_sg U70497 ( .A(n56885), .B(n68422), .X(n32628) );
  nand_x2_sg U70498 ( .A(n32632), .B(n32633), .X(n32631) );
  nor_x1_sg U70499 ( .A(n51457), .B(n47721), .X(n32632) );
  nor_x1_sg U70500 ( .A(n56887), .B(n68423), .X(n32633) );
  nand_x2_sg U70501 ( .A(n32120), .B(n32121), .X(n32119) );
  nor_x1_sg U70502 ( .A(n47565), .B(n51439), .X(n32120) );
  nor_x1_sg U70503 ( .A(n56877), .B(n68530), .X(n32121) );
  nand_x2_sg U70504 ( .A(n32123), .B(n32124), .X(n32118) );
  nor_x1_sg U70505 ( .A(n56879), .B(n47567), .X(n32123) );
  nor_x1_sg U70506 ( .A(n51433), .B(n68531), .X(n32124) );
  nand_x2_sg U70507 ( .A(n32128), .B(n32129), .X(n32127) );
  nor_x1_sg U70508 ( .A(n56881), .B(n47563), .X(n32128) );
  nor_x1_sg U70509 ( .A(n51435), .B(n68532), .X(n32129) );
  nand_x2_sg U70510 ( .A(n32565), .B(n32566), .X(n32564) );
  nor_x1_sg U70511 ( .A(n47559), .B(n51431), .X(n32565) );
  nor_x1_sg U70512 ( .A(n56869), .B(n68438), .X(n32566) );
  nand_x2_sg U70513 ( .A(n32568), .B(n32569), .X(n32563) );
  nor_x1_sg U70514 ( .A(n56871), .B(n47561), .X(n32568) );
  nor_x1_sg U70515 ( .A(n51425), .B(n68439), .X(n32569) );
  nand_x2_sg U70516 ( .A(n32573), .B(n32574), .X(n32572) );
  nor_x1_sg U70517 ( .A(n56873), .B(n47557), .X(n32573) );
  nor_x1_sg U70518 ( .A(n51427), .B(n68440), .X(n32574) );
  nor_x1_sg U70519 ( .A(n56863), .B(n68555), .X(n32274) );
  nor_x1_sg U70520 ( .A(n47705), .B(n51413), .X(n32275) );
  nor_x1_sg U70521 ( .A(n51263), .B(n56725), .X(n32264) );
  nor_x1_sg U70522 ( .A(n51373), .B(n56819), .X(n32267) );
  nor_x1_sg U70523 ( .A(n51375), .B(n56821), .X(n32272) );
  nand_x2_sg U70524 ( .A(n32262), .B(n32263), .X(n32261) );
  nor_x1_sg U70525 ( .A(n47633), .B(n56777), .X(n32262) );
  nor_x1_sg U70526 ( .A(n51219), .B(n68552), .X(n32263) );
  nand_x2_sg U70527 ( .A(n32265), .B(n32266), .X(n32260) );
  nor_x1_sg U70528 ( .A(n51221), .B(n47635), .X(n32265) );
  nor_x1_sg U70529 ( .A(n56683), .B(n68553), .X(n32266) );
  nand_x2_sg U70530 ( .A(n32270), .B(n32271), .X(n32269) );
  nor_x1_sg U70531 ( .A(n51313), .B(n47631), .X(n32270) );
  nor_x1_sg U70532 ( .A(n56771), .B(n68554), .X(n32271) );
  nor_x1_sg U70533 ( .A(n47681), .B(n68471), .X(n32683) );
  nor_x1_sg U70534 ( .A(n51391), .B(n56833), .X(n32684) );
  nor_x1_sg U70535 ( .A(n51251), .B(n56713), .X(n32673) );
  nor_x1_sg U70536 ( .A(n51253), .B(n56715), .X(n32676) );
  nor_x1_sg U70537 ( .A(n51255), .B(n56717), .X(n32681) );
  nand_x2_sg U70538 ( .A(n32671), .B(n32672), .X(n32670) );
  nor_x1_sg U70539 ( .A(n47625), .B(n56671), .X(n32671) );
  nor_x1_sg U70540 ( .A(n51207), .B(n68468), .X(n32672) );
  nand_x2_sg U70541 ( .A(n32674), .B(n32675), .X(n32669) );
  nor_x1_sg U70542 ( .A(n51209), .B(n47627), .X(n32674) );
  nor_x1_sg U70543 ( .A(n56667), .B(n68469), .X(n32675) );
  nand_x2_sg U70544 ( .A(n32679), .B(n32680), .X(n32678) );
  nor_x1_sg U70545 ( .A(n51211), .B(n47623), .X(n32679) );
  nor_x1_sg U70546 ( .A(n56669), .B(n68470), .X(n32680) );
  nor_x1_sg U70547 ( .A(n47693), .B(n68564), .X(n32238) );
  nor_x1_sg U70548 ( .A(n51405), .B(n56845), .X(n32239) );
  nor_x1_sg U70549 ( .A(n51271), .B(n56733), .X(n32228) );
  nor_x1_sg U70550 ( .A(n51273), .B(n56735), .X(n32231) );
  nor_x1_sg U70551 ( .A(n51275), .B(n56737), .X(n32236) );
  nand_x2_sg U70552 ( .A(n32226), .B(n32227), .X(n32225) );
  nor_x1_sg U70553 ( .A(n47645), .B(n56695), .X(n32226) );
  nor_x1_sg U70554 ( .A(n51229), .B(n68561), .X(n32227) );
  nand_x2_sg U70555 ( .A(n32229), .B(n32230), .X(n32224) );
  nor_x1_sg U70556 ( .A(n51231), .B(n47647), .X(n32229) );
  nor_x1_sg U70557 ( .A(n56691), .B(n68562), .X(n32230) );
  nand_x2_sg U70558 ( .A(n32234), .B(n32235), .X(n32233) );
  nor_x1_sg U70559 ( .A(n51233), .B(n47643), .X(n32234) );
  nor_x1_sg U70560 ( .A(n56693), .B(n68563), .X(n32235) );
  nor_x1_sg U70561 ( .A(n47683), .B(n68476), .X(n32701) );
  nor_x1_sg U70562 ( .A(n51393), .B(n56835), .X(n32702) );
  nor_x1_sg U70563 ( .A(n51361), .B(n56809), .X(n32691) );
  nor_x1_sg U70564 ( .A(n47669), .B(n51363), .X(n32694) );
  nor_x1_sg U70565 ( .A(n51257), .B(n56719), .X(n32699) );
  nand_x2_sg U70566 ( .A(n32689), .B(n32690), .X(n32688) );
  nor_x1_sg U70567 ( .A(n47659), .B(n56673), .X(n32689) );
  nor_x1_sg U70568 ( .A(n51299), .B(n68473), .X(n32690) );
  nand_x2_sg U70569 ( .A(n32692), .B(n32693), .X(n32687) );
  nor_x1_sg U70570 ( .A(n47661), .B(n47551), .X(n32692) );
  nor_x1_sg U70571 ( .A(n51301), .B(n68474), .X(n32693) );
  nand_x2_sg U70572 ( .A(n32697), .B(n32698), .X(n32696) );
  nor_x1_sg U70573 ( .A(n47663), .B(n47549), .X(n32697) );
  nor_x1_sg U70574 ( .A(n51303), .B(n68475), .X(n32698) );
  nor_x1_sg U70575 ( .A(n51277), .B(n56739), .X(n32246) );
  nor_x1_sg U70576 ( .A(n47671), .B(n51377), .X(n32249) );
  nor_x1_sg U70577 ( .A(n51379), .B(n56823), .X(n32254) );
  nor_x1_sg U70578 ( .A(n51423), .B(n68569), .X(n32256) );
  nor_x1_sg U70579 ( .A(n47707), .B(n56859), .X(n32257) );
  nand_x1_sg U70580 ( .A(n47299), .B(n38411), .X(n38408) );
  nand_x1_sg U70581 ( .A(n57522), .B(state[1]), .X(n38409) );
  nand_x2_sg U70582 ( .A(n32244), .B(n32245), .X(n32243) );
  nor_x1_sg U70583 ( .A(n56697), .B(n51329), .X(n32244) );
  nor_x1_sg U70584 ( .A(n47649), .B(n68566), .X(n32245) );
  nand_x2_sg U70585 ( .A(n32247), .B(n32248), .X(n32242) );
  nor_x1_sg U70586 ( .A(n47651), .B(n47535), .X(n32247) );
  nor_x1_sg U70587 ( .A(n51235), .B(n68567), .X(n32248) );
  nand_x2_sg U70588 ( .A(n32252), .B(n32253), .X(n32251) );
  nor_x1_sg U70589 ( .A(n47665), .B(n47533), .X(n32252) );
  nor_x1_sg U70590 ( .A(n51317), .B(n68568), .X(n32253) );
  nor_x1_sg U70591 ( .A(n47691), .B(n68560), .X(n32332) );
  nor_x1_sg U70592 ( .A(n51403), .B(n56843), .X(n32333) );
  nor_x1_sg U70593 ( .A(n47679), .B(n68467), .X(n32777) );
  nor_x1_sg U70594 ( .A(n51389), .B(n56831), .X(n32778) );
  nor_x1_sg U70595 ( .A(n51265), .B(n56727), .X(n32322) );
  nor_x1_sg U70596 ( .A(n51267), .B(n56729), .X(n32325) );
  nor_x1_sg U70597 ( .A(n51269), .B(n56731), .X(n32330) );
  nor_x1_sg U70598 ( .A(n51245), .B(n56707), .X(n32767) );
  nor_x1_sg U70599 ( .A(n51247), .B(n56709), .X(n32770) );
  nor_x1_sg U70600 ( .A(n51249), .B(n56711), .X(n32775) );
  nand_x2_sg U70601 ( .A(n32320), .B(n32321), .X(n32319) );
  nor_x1_sg U70602 ( .A(n47639), .B(n56689), .X(n32320) );
  nor_x1_sg U70603 ( .A(n51223), .B(n68557), .X(n32321) );
  nand_x2_sg U70604 ( .A(n32323), .B(n32324), .X(n32318) );
  nor_x1_sg U70605 ( .A(n51225), .B(n47641), .X(n32323) );
  nor_x1_sg U70606 ( .A(n56685), .B(n68558), .X(n32324) );
  nand_x2_sg U70607 ( .A(n32328), .B(n32329), .X(n32327) );
  nor_x1_sg U70608 ( .A(n51227), .B(n47637), .X(n32328) );
  nor_x1_sg U70609 ( .A(n56687), .B(n68559), .X(n32329) );
  nand_x2_sg U70610 ( .A(n32765), .B(n32766), .X(n32764) );
  nor_x1_sg U70611 ( .A(n47619), .B(n56665), .X(n32765) );
  nor_x1_sg U70612 ( .A(n51201), .B(n68464), .X(n32766) );
  nand_x2_sg U70613 ( .A(n32768), .B(n32769), .X(n32763) );
  nor_x1_sg U70614 ( .A(n51203), .B(n47621), .X(n32768) );
  nor_x1_sg U70615 ( .A(n56661), .B(n68465), .X(n32769) );
  nand_x2_sg U70616 ( .A(n32773), .B(n32774), .X(n32772) );
  nor_x1_sg U70617 ( .A(n51205), .B(n47617), .X(n32773) );
  nor_x1_sg U70618 ( .A(n56663), .B(n68466), .X(n32774) );
  nor_x1_sg U70619 ( .A(n47351), .B(n47439), .X(n39705) );
  nor_x1_sg U70620 ( .A(n56829), .B(n51387), .X(n32596) );
  nor_x1_sg U70621 ( .A(n56841), .B(n51401), .X(n32151) );
  nor_x1_sg U70622 ( .A(n56761), .B(n51297), .X(n32718) );
  nor_x1_sg U70623 ( .A(n56911), .B(n51481), .X(n32190) );
  nor_x1_sg U70624 ( .A(n56903), .B(n51471), .X(n32635) );
  nor_x1_sg U70625 ( .A(n51437), .B(n56883), .X(n32131) );
  nor_x1_sg U70626 ( .A(n51429), .B(n56875), .X(n32576) );
  nor_x1_sg U70627 ( .A(n51419), .B(n68545), .X(n32314) );
  nor_x1_sg U70628 ( .A(n47555), .B(n56855), .X(n32315) );
  nor_x1_sg U70629 ( .A(n56773), .B(n51315), .X(n32273) );
  nor_x1_sg U70630 ( .A(n51415), .B(n68452), .X(n32759) );
  nor_x1_sg U70631 ( .A(n47553), .B(n56851), .X(n32760) );
  nor_x1_sg U70632 ( .A(n56721), .B(n51259), .X(n32304) );
  nor_x1_sg U70633 ( .A(n56811), .B(n51365), .X(n32307) );
  nor_x1_sg U70634 ( .A(n56813), .B(n51367), .X(n32312) );
  nor_x1_sg U70635 ( .A(n56791), .B(n51343), .X(n32749) );
  nor_x1_sg U70636 ( .A(n56793), .B(n51345), .X(n32752) );
  nor_x1_sg U70637 ( .A(n56795), .B(n51347), .X(n32757) );
  nand_x2_sg U70638 ( .A(n32302), .B(n32303), .X(n32301) );
  nor_x1_sg U70639 ( .A(n47523), .B(n51325), .X(n32302) );
  nor_x1_sg U70640 ( .A(n56675), .B(n68542), .X(n32303) );
  nand_x2_sg U70641 ( .A(n32305), .B(n32306), .X(n32300) );
  nor_x1_sg U70642 ( .A(n56677), .B(n47525), .X(n32305) );
  nor_x1_sg U70643 ( .A(n51215), .B(n68543), .X(n32306) );
  nand_x2_sg U70644 ( .A(n32310), .B(n32311), .X(n32309) );
  nor_x1_sg U70645 ( .A(n56763), .B(n47521), .X(n32310) );
  nor_x1_sg U70646 ( .A(n51305), .B(n68544), .X(n32311) );
  nand_x2_sg U70647 ( .A(n32747), .B(n32748), .X(n32746) );
  nor_x1_sg U70648 ( .A(n47539), .B(n51321), .X(n32747) );
  nor_x1_sg U70649 ( .A(n56741), .B(n68449), .X(n32748) );
  nand_x2_sg U70650 ( .A(n32750), .B(n32751), .X(n32745) );
  nor_x1_sg U70651 ( .A(n56743), .B(n47541), .X(n32750) );
  nor_x1_sg U70652 ( .A(n51279), .B(n68450), .X(n32751) );
  nand_x2_sg U70653 ( .A(n32755), .B(n32756), .X(n32754) );
  nor_x1_sg U70654 ( .A(n56745), .B(n47537), .X(n32755) );
  nor_x1_sg U70655 ( .A(n51281), .B(n68451), .X(n32756) );
  nor_x1_sg U70656 ( .A(n55155), .B(n32171), .X(n32170) );
  nor_x1_sg U70657 ( .A(n55153), .B(n32616), .X(n32615) );
  nand_x2_sg U70658 ( .A(n32158), .B(n32159), .X(n32157) );
  nor_x1_sg U70659 ( .A(n47609), .B(n55083), .X(n32158) );
  nor_x1_sg U70660 ( .A(n51141), .B(n32160), .X(n32159) );
  nand_x2_sg U70661 ( .A(n32161), .B(n32162), .X(n32156) );
  nor_x1_sg U70662 ( .A(n51143), .B(n47611), .X(n32161) );
  nor_x1_sg U70663 ( .A(n55079), .B(n32163), .X(n32162) );
  nand_x2_sg U70664 ( .A(n32166), .B(n32167), .X(n32165) );
  nor_x1_sg U70665 ( .A(n51145), .B(n47607), .X(n32166) );
  nor_x1_sg U70666 ( .A(n55081), .B(n32168), .X(n32167) );
  nand_x2_sg U70667 ( .A(n32603), .B(n32604), .X(n32602) );
  nor_x1_sg U70668 ( .A(n47603), .B(n55077), .X(n32603) );
  nor_x1_sg U70669 ( .A(n51135), .B(n32605), .X(n32604) );
  nand_x2_sg U70670 ( .A(n32606), .B(n32607), .X(n32601) );
  nor_x1_sg U70671 ( .A(n51137), .B(n47605), .X(n32606) );
  nor_x1_sg U70672 ( .A(n55073), .B(n32608), .X(n32607) );
  nand_x2_sg U70673 ( .A(n32611), .B(n32612), .X(n32610) );
  nor_x1_sg U70674 ( .A(n51139), .B(n47601), .X(n32611) );
  nor_x1_sg U70675 ( .A(n55075), .B(n32613), .X(n32612) );
  nor_x1_sg U70676 ( .A(n56705), .B(n51243), .X(n32237) );
  nor_x1_sg U70677 ( .A(n56701), .B(n51239), .X(n32682) );
  nor_x1_sg U70678 ( .A(n51213), .B(n47629), .X(n32700) );
  nand_x1_sg U70679 ( .A(n47352), .B(n51065), .X(n34229) );
  nor_x1_sg U70680 ( .A(n51319), .B(n47667), .X(n32255) );
  nand_x1_sg U70681 ( .A(n32820), .B(n47437), .X(n34224) );
  nor_x1_sg U70682 ( .A(n47318), .B(n32820), .X(n34226) );
  nor_x1_sg U70683 ( .A(n51421), .B(n68550), .X(n32351) );
  nor_x1_sg U70684 ( .A(n56857), .B(n47703), .X(n32352) );
  nor_x1_sg U70685 ( .A(n51417), .B(n68457), .X(n32796) );
  nor_x1_sg U70686 ( .A(n56853), .B(n47699), .X(n32797) );
  nor_x1_sg U70687 ( .A(n56723), .B(n51261), .X(n32341) );
  nor_x1_sg U70688 ( .A(n56815), .B(n51369), .X(n32344) );
  nor_x1_sg U70689 ( .A(n56817), .B(n51371), .X(n32349) );
  nor_x1_sg U70690 ( .A(n56797), .B(n51349), .X(n32786) );
  nor_x1_sg U70691 ( .A(n56799), .B(n51351), .X(n32789) );
  nor_x1_sg U70692 ( .A(n56801), .B(n51353), .X(n32794) );
  nand_x2_sg U70693 ( .A(n32339), .B(n32340), .X(n32338) );
  nor_x1_sg U70694 ( .A(n47529), .B(n51327), .X(n32339) );
  nor_x1_sg U70695 ( .A(n56679), .B(n68547), .X(n32340) );
  nand_x2_sg U70696 ( .A(n32342), .B(n32343), .X(n32337) );
  nor_x1_sg U70697 ( .A(n56681), .B(n47531), .X(n32342) );
  nor_x1_sg U70698 ( .A(n51217), .B(n68548), .X(n32343) );
  nand_x2_sg U70699 ( .A(n32347), .B(n32348), .X(n32346) );
  nor_x1_sg U70700 ( .A(n56767), .B(n47527), .X(n32347) );
  nor_x1_sg U70701 ( .A(n51309), .B(n68549), .X(n32348) );
  nand_x2_sg U70702 ( .A(n32784), .B(n32785), .X(n32783) );
  nor_x1_sg U70703 ( .A(n47545), .B(n51323), .X(n32784) );
  nor_x1_sg U70704 ( .A(n56749), .B(n68454), .X(n32785) );
  nand_x2_sg U70705 ( .A(n32787), .B(n32788), .X(n32782) );
  nor_x1_sg U70706 ( .A(n56751), .B(n47547), .X(n32787) );
  nor_x1_sg U70707 ( .A(n51285), .B(n68455), .X(n32788) );
  nand_x2_sg U70708 ( .A(n32792), .B(n32793), .X(n32791) );
  nor_x1_sg U70709 ( .A(n56753), .B(n47543), .X(n32792) );
  nor_x1_sg U70710 ( .A(n51287), .B(n68456), .X(n32793) );
  nor_x1_sg U70711 ( .A(n56933), .B(n32210), .X(n32209) );
  nor_x1_sg U70712 ( .A(n56931), .B(n32655), .X(n32654) );
  nand_x2_sg U70713 ( .A(n32197), .B(n32198), .X(n32196) );
  nor_x1_sg U70714 ( .A(n47367), .B(n47435), .X(n32197) );
  nor_x1_sg U70715 ( .A(n56923), .B(n32199), .X(n32198) );
  nand_x2_sg U70716 ( .A(n32200), .B(n32201), .X(n32195) );
  nor_x1_sg U70717 ( .A(n47429), .B(n47369), .X(n32200) );
  nor_x1_sg U70718 ( .A(n56925), .B(n32202), .X(n32201) );
  nand_x2_sg U70719 ( .A(n32205), .B(n32206), .X(n32204) );
  nor_x1_sg U70720 ( .A(n47431), .B(n47365), .X(n32205) );
  nor_x1_sg U70721 ( .A(n56927), .B(n32207), .X(n32206) );
  nand_x2_sg U70722 ( .A(n32642), .B(n32643), .X(n32641) );
  nor_x1_sg U70723 ( .A(n47359), .B(n47427), .X(n32642) );
  nor_x1_sg U70724 ( .A(n56917), .B(n32644), .X(n32643) );
  nand_x2_sg U70725 ( .A(n32645), .B(n32646), .X(n32640) );
  nor_x1_sg U70726 ( .A(n47421), .B(n47361), .X(n32645) );
  nor_x1_sg U70727 ( .A(n56919), .B(n32647), .X(n32646) );
  nand_x2_sg U70728 ( .A(n32650), .B(n32651), .X(n32649) );
  nor_x1_sg U70729 ( .A(n47423), .B(n47357), .X(n32650) );
  nor_x1_sg U70730 ( .A(n56921), .B(n32652), .X(n32651) );
  nor_x1_sg U70731 ( .A(n56703), .B(n51241), .X(n32331) );
  nor_x1_sg U70732 ( .A(n56699), .B(n51237), .X(n32776) );
  nor_x1_sg U70733 ( .A(n55085), .B(n51147), .X(n32614) );
  nor_x1_sg U70734 ( .A(n55087), .B(n51149), .X(n32169) );
  nand_x1_sg U70735 ( .A(n47411), .B(n57170), .X(n32819) );
  nand_x1_sg U70736 ( .A(n32820), .B(n47353), .X(n32818) );
  nor_x1_sg U70737 ( .A(n47433), .B(n47371), .X(n32208) );
  nor_x1_sg U70738 ( .A(n47425), .B(n47363), .X(n32653) );
  nor_x1_sg U70739 ( .A(n51307), .B(n56765), .X(n32313) );
  nor_x1_sg U70740 ( .A(n51283), .B(n56747), .X(n32758) );
  nor_x1_sg U70741 ( .A(n56769), .B(n51311), .X(n32350) );
  nor_x1_sg U70742 ( .A(n56755), .B(n51289), .X(n32795) );
  nor_x1_sg U70743 ( .A(n57089), .B(n32060), .X(n32059) );
  nand_x2_sg U70744 ( .A(n32046), .B(n32047), .X(n32045) );
  nor_x1_sg U70745 ( .A(n57081), .B(n51549), .X(n32046) );
  nor_x1_sg U70746 ( .A(n47773), .B(n32048), .X(n32047) );
  nand_x2_sg U70747 ( .A(n32049), .B(n32050), .X(n32044) );
  nor_x1_sg U70748 ( .A(n51545), .B(n32052), .X(n32049) );
  nor_x1_sg U70749 ( .A(n57071), .B(n32051), .X(n32050) );
  nor_x1_sg U70750 ( .A(n57085), .B(n32506), .X(n32505) );
  nand_x2_sg U70751 ( .A(n32489), .B(n32490), .X(n32488) );
  nor_x1_sg U70752 ( .A(n51543), .B(n47759), .X(n32489) );
  nor_x1_sg U70753 ( .A(n57073), .B(n32491), .X(n32490) );
  nand_x2_sg U70754 ( .A(n32492), .B(n32493), .X(n32487) );
  nor_x1_sg U70755 ( .A(n51547), .B(n32495), .X(n32492) );
  nor_x1_sg U70756 ( .A(n57075), .B(n32494), .X(n32493) );
  nor_x1_sg U70757 ( .A(n47519), .B(n68508), .X(n32018) );
  nor_x1_sg U70758 ( .A(n55251), .B(n51181), .X(n32019) );
  nor_x1_sg U70759 ( .A(n47517), .B(n68419), .X(n32460) );
  nor_x1_sg U70760 ( .A(n55249), .B(n51179), .X(n32461) );
  nor_x1_sg U70761 ( .A(n55235), .B(n51163), .X(n32008) );
  nor_x1_sg U70762 ( .A(n55239), .B(n51167), .X(n32011) );
  nor_x1_sg U70763 ( .A(n55243), .B(n51171), .X(n32016) );
  nor_x1_sg U70764 ( .A(n55223), .B(n51153), .X(n32450) );
  nor_x1_sg U70765 ( .A(n55227), .B(n51157), .X(n32453) );
  nor_x1_sg U70766 ( .A(n55231), .B(n51161), .X(n32458) );
  nand_x2_sg U70767 ( .A(n32006), .B(n32007), .X(n32005) );
  nor_x1_sg U70768 ( .A(n47513), .B(n51173), .X(n32006) );
  nor_x1_sg U70769 ( .A(n55233), .B(n68505), .X(n32007) );
  nand_x2_sg U70770 ( .A(n32009), .B(n32010), .X(n32004) );
  nor_x1_sg U70771 ( .A(n55237), .B(n47515), .X(n32009) );
  nor_x1_sg U70772 ( .A(n51165), .B(n68506), .X(n32010) );
  nand_x2_sg U70773 ( .A(n32014), .B(n32015), .X(n32013) );
  nor_x1_sg U70774 ( .A(n55241), .B(n47511), .X(n32014) );
  nor_x1_sg U70775 ( .A(n51169), .B(n68507), .X(n32015) );
  nand_x2_sg U70776 ( .A(n32448), .B(n32449), .X(n32447) );
  nor_x1_sg U70777 ( .A(n51151), .B(n47613), .X(n32448) );
  nor_x1_sg U70778 ( .A(n55221), .B(n68416), .X(n32449) );
  nand_x2_sg U70779 ( .A(n32451), .B(n32452), .X(n32446) );
  nor_x1_sg U70780 ( .A(n55225), .B(n47509), .X(n32451) );
  nor_x1_sg U70781 ( .A(n51155), .B(n68417), .X(n32452) );
  nand_x2_sg U70782 ( .A(n32456), .B(n32457), .X(n32455) );
  nor_x1_sg U70783 ( .A(n55229), .B(n47507), .X(n32456) );
  nor_x1_sg U70784 ( .A(n51159), .B(n68418), .X(n32457) );
  nor_x1_sg U70785 ( .A(n55261), .B(n32469), .X(n32468) );
  nor_x1_sg U70786 ( .A(n55265), .B(n32472), .X(n32471) );
  nor_x1_sg U70787 ( .A(n55267), .B(n32477), .X(n32476) );
  nor_x1_sg U70788 ( .A(n55271), .B(n32480), .X(n32479) );
  nand_x2_sg U70789 ( .A(n32470), .B(n32471), .X(n32465) );
  nand_x2_sg U70790 ( .A(n32467), .B(n32468), .X(n32466) );
  nor_x1_sg U70791 ( .A(n55263), .B(n51191), .X(n32470) );
  nand_x2_sg U70792 ( .A(n32478), .B(n32479), .X(n32473) );
  nand_x2_sg U70793 ( .A(n32475), .B(n32476), .X(n32474) );
  nor_x1_sg U70794 ( .A(n55269), .B(n51193), .X(n32478) );
  nor_x1_sg U70795 ( .A(n55273), .B(n32027), .X(n32026) );
  nor_x1_sg U70796 ( .A(n55277), .B(n32030), .X(n32029) );
  nor_x1_sg U70797 ( .A(n55279), .B(n32035), .X(n32034) );
  nor_x1_sg U70798 ( .A(n55283), .B(n32038), .X(n32037) );
  nand_x2_sg U70799 ( .A(n32028), .B(n32029), .X(n32023) );
  nand_x2_sg U70800 ( .A(n32025), .B(n32026), .X(n32024) );
  nor_x1_sg U70801 ( .A(n55275), .B(n51195), .X(n32028) );
  nand_x2_sg U70802 ( .A(n32036), .B(n32037), .X(n32031) );
  nand_x2_sg U70803 ( .A(n32033), .B(n32034), .X(n32032) );
  nor_x1_sg U70804 ( .A(n55281), .B(n51197), .X(n32036) );
  nand_x1_sg U70805 ( .A(n39699), .B(n56929), .X(n39698) );
  nand_x1_sg U70806 ( .A(n51199), .B(n39700), .X(n39697) );
  nor_x1_sg U70807 ( .A(n51199), .B(n68370), .X(n39699) );
  nor_x1_sg U70808 ( .A(n51189), .B(n55259), .X(n32025) );
  nor_x1_sg U70809 ( .A(n55257), .B(n51187), .X(n32033) );
  nor_x1_sg U70810 ( .A(n51185), .B(n55255), .X(n32467) );
  nor_x1_sg U70811 ( .A(n55253), .B(n51183), .X(n32475) );
  nor_x1_sg U70812 ( .A(n51177), .B(n55247), .X(n32017) );
  nor_x1_sg U70813 ( .A(n51175), .B(n55245), .X(n32459) );
  nor_x1_sg U70814 ( .A(n51199), .B(n56929), .X(n35843) );
  nor_x1_sg U70815 ( .A(n35836), .B(n35705), .X(n44270) );
  nand_x2_sg U70816 ( .A(n35844), .B(n56928), .X(n39701) );
  nand_x1_sg U70817 ( .A(n39704), .B(n56929), .X(n39703) );
  nor_x1_sg U70818 ( .A(n35844), .B(n68269), .X(n39704) );
  nor_x1_sg U70819 ( .A(n68368), .B(n55151), .X(n40224) );
  nor_x1_sg U70820 ( .A(n68367), .B(n55149), .X(n40219) );
  nor_x1_sg U70821 ( .A(n68366), .B(n55147), .X(n40214) );
  nor_x1_sg U70822 ( .A(n68365), .B(n55145), .X(n40209) );
  nor_x1_sg U70823 ( .A(n68364), .B(n55219), .X(n40204) );
  nor_x1_sg U70824 ( .A(n68363), .B(n55217), .X(n40199) );
  nor_x1_sg U70825 ( .A(n68362), .B(n55215), .X(n40194) );
  nor_x1_sg U70826 ( .A(n68361), .B(n55213), .X(n40189) );
  nor_x1_sg U70827 ( .A(n68360), .B(n55211), .X(n40184) );
  nor_x1_sg U70828 ( .A(n68359), .B(n55209), .X(n40179) );
  nor_x1_sg U70829 ( .A(n68358), .B(n55207), .X(n40174) );
  nor_x1_sg U70830 ( .A(n68357), .B(n55205), .X(n40169) );
  nor_x1_sg U70831 ( .A(n68356), .B(n55203), .X(n40164) );
  nor_x1_sg U70832 ( .A(n68355), .B(n55201), .X(n40159) );
  nor_x1_sg U70833 ( .A(n68354), .B(n55143), .X(n40154) );
  nor_x1_sg U70834 ( .A(n68353), .B(n55199), .X(n40149) );
  nor_x1_sg U70835 ( .A(n68352), .B(n55197), .X(n40144) );
  nor_x1_sg U70836 ( .A(n68351), .B(n55195), .X(n40139) );
  nor_x1_sg U70837 ( .A(n68350), .B(n55193), .X(n40134) );
  nor_x1_sg U70838 ( .A(n68349), .B(n55191), .X(n40129) );
  nor_x1_sg U70839 ( .A(n68348), .B(n55189), .X(n40124) );
  nor_x1_sg U70840 ( .A(n68347), .B(n55187), .X(n40119) );
  nor_x1_sg U70841 ( .A(n68346), .B(n55185), .X(n40114) );
  nor_x1_sg U70842 ( .A(n68345), .B(n55183), .X(n40109) );
  nor_x1_sg U70843 ( .A(n68344), .B(n55181), .X(n40104) );
  nor_x1_sg U70844 ( .A(n68343), .B(n55179), .X(n40099) );
  nor_x1_sg U70845 ( .A(n68342), .B(n55141), .X(n40094) );
  nor_x1_sg U70846 ( .A(n68341), .B(n55139), .X(n40089) );
  nor_x1_sg U70847 ( .A(n68340), .B(n55177), .X(n40084) );
  nor_x1_sg U70848 ( .A(n68339), .B(n55175), .X(n40079) );
  nor_x1_sg U70849 ( .A(n68338), .B(n55173), .X(n40074) );
  nor_x1_sg U70850 ( .A(n68337), .B(n55137), .X(n40069) );
  nor_x1_sg U70851 ( .A(n68368), .B(n55171), .X(n40064) );
  nor_x1_sg U70852 ( .A(n68367), .B(n55169), .X(n40059) );
  nor_x1_sg U70853 ( .A(n68366), .B(n55167), .X(n40054) );
  nor_x1_sg U70854 ( .A(n68365), .B(n55165), .X(n40049) );
  nor_x1_sg U70855 ( .A(n68364), .B(n55135), .X(n40044) );
  nor_x1_sg U70856 ( .A(n68363), .B(n55133), .X(n40039) );
  nor_x1_sg U70857 ( .A(n68362), .B(n55131), .X(n40034) );
  nor_x1_sg U70858 ( .A(n68361), .B(n55129), .X(n40029) );
  nor_x1_sg U70859 ( .A(n68360), .B(n55127), .X(n40024) );
  nor_x1_sg U70860 ( .A(n68359), .B(n55125), .X(n40019) );
  nor_x1_sg U70861 ( .A(n68358), .B(n55123), .X(n40014) );
  nor_x1_sg U70862 ( .A(n68357), .B(n55121), .X(n40009) );
  nor_x1_sg U70863 ( .A(n68356), .B(n55119), .X(n40004) );
  nor_x1_sg U70864 ( .A(n68355), .B(n55117), .X(n39999) );
  nor_x1_sg U70865 ( .A(n68354), .B(n55163), .X(n39994) );
  nor_x1_sg U70866 ( .A(n68353), .B(n55115), .X(n39989) );
  nor_x1_sg U70867 ( .A(n68352), .B(n55113), .X(n39984) );
  nor_x1_sg U70868 ( .A(n68351), .B(n55111), .X(n39979) );
  nor_x1_sg U70869 ( .A(n68350), .B(n55109), .X(n39974) );
  nor_x1_sg U70870 ( .A(n68349), .B(n55107), .X(n39969) );
  nor_x1_sg U70871 ( .A(n68348), .B(n55105), .X(n39964) );
  nor_x1_sg U70872 ( .A(n68347), .B(n55103), .X(n39959) );
  nor_x1_sg U70873 ( .A(n68346), .B(n55101), .X(n39954) );
  nor_x1_sg U70874 ( .A(n68345), .B(n55099), .X(n39949) );
  nor_x1_sg U70875 ( .A(n68344), .B(n55097), .X(n39944) );
  nor_x1_sg U70876 ( .A(n68343), .B(n55095), .X(n39939) );
  nor_x1_sg U70877 ( .A(n68342), .B(n55161), .X(n39934) );
  nor_x1_sg U70878 ( .A(n68341), .B(n55159), .X(n39929) );
  nor_x1_sg U70879 ( .A(n68340), .B(n55093), .X(n39924) );
  nor_x1_sg U70880 ( .A(n68339), .B(n55091), .X(n39919) );
  nor_x1_sg U70881 ( .A(n68338), .B(n55089), .X(n39914) );
  nor_x1_sg U70882 ( .A(n68337), .B(n55157), .X(n39909) );
  nand_x1_sg U70883 ( .A(n55151), .B(n68368), .X(n40223) );
  nand_x1_sg U70884 ( .A(n55149), .B(n68367), .X(n40218) );
  nand_x1_sg U70885 ( .A(n55147), .B(n68366), .X(n40213) );
  nand_x1_sg U70886 ( .A(n55145), .B(n68365), .X(n40208) );
  nand_x1_sg U70887 ( .A(n55219), .B(n68364), .X(n40203) );
  nand_x1_sg U70888 ( .A(n55217), .B(n68363), .X(n40198) );
  nand_x1_sg U70889 ( .A(n55215), .B(n68362), .X(n40193) );
  nand_x1_sg U70890 ( .A(n55213), .B(n68361), .X(n40188) );
  nand_x1_sg U70891 ( .A(n55211), .B(n68360), .X(n40183) );
  nand_x1_sg U70892 ( .A(n55209), .B(n68359), .X(n40178) );
  nand_x1_sg U70893 ( .A(n55207), .B(n68358), .X(n40173) );
  nand_x1_sg U70894 ( .A(n55205), .B(n68357), .X(n40168) );
  nand_x1_sg U70895 ( .A(n55203), .B(n68356), .X(n40163) );
  nand_x1_sg U70896 ( .A(n55201), .B(n68355), .X(n40158) );
  nand_x1_sg U70897 ( .A(n55143), .B(n68354), .X(n40153) );
  nand_x1_sg U70898 ( .A(n55199), .B(n68353), .X(n40148) );
  nand_x1_sg U70899 ( .A(n55197), .B(n68352), .X(n40143) );
  nand_x1_sg U70900 ( .A(n55195), .B(n68351), .X(n40138) );
  nand_x1_sg U70901 ( .A(n55193), .B(n68350), .X(n40133) );
  nand_x1_sg U70902 ( .A(n55191), .B(n68349), .X(n40128) );
  nand_x1_sg U70903 ( .A(n55189), .B(n68348), .X(n40123) );
  nand_x1_sg U70904 ( .A(n55187), .B(n68347), .X(n40118) );
  nand_x1_sg U70905 ( .A(n55185), .B(n68346), .X(n40113) );
  nand_x1_sg U70906 ( .A(n55183), .B(n68345), .X(n40108) );
  nand_x1_sg U70907 ( .A(n55181), .B(n68344), .X(n40103) );
  nand_x1_sg U70908 ( .A(n55179), .B(n68343), .X(n40098) );
  nand_x1_sg U70909 ( .A(n55141), .B(n68342), .X(n40093) );
  nand_x1_sg U70910 ( .A(n55139), .B(n68341), .X(n40088) );
  nand_x1_sg U70911 ( .A(n55177), .B(n68340), .X(n40083) );
  nand_x1_sg U70912 ( .A(n55175), .B(n68339), .X(n40078) );
  nand_x1_sg U70913 ( .A(n55173), .B(n68338), .X(n40073) );
  nand_x1_sg U70914 ( .A(n55137), .B(n68337), .X(n40068) );
  nand_x1_sg U70915 ( .A(n55171), .B(n68368), .X(n40063) );
  nand_x1_sg U70916 ( .A(n55169), .B(n68367), .X(n40058) );
  nand_x1_sg U70917 ( .A(n55167), .B(n68366), .X(n40053) );
  nand_x1_sg U70918 ( .A(n55165), .B(n68365), .X(n40048) );
  nand_x1_sg U70919 ( .A(n55135), .B(n68364), .X(n40043) );
  nand_x1_sg U70920 ( .A(n55133), .B(n68363), .X(n40038) );
  nand_x1_sg U70921 ( .A(n55131), .B(n68362), .X(n40033) );
  nand_x1_sg U70922 ( .A(n55129), .B(n68361), .X(n40028) );
  nand_x1_sg U70923 ( .A(n55127), .B(n68360), .X(n40023) );
  nand_x1_sg U70924 ( .A(n55125), .B(n68359), .X(n40018) );
  nand_x1_sg U70925 ( .A(n55123), .B(n68358), .X(n40013) );
  nand_x1_sg U70926 ( .A(n55121), .B(n68357), .X(n40008) );
  nand_x1_sg U70927 ( .A(n55119), .B(n68356), .X(n40003) );
  nand_x1_sg U70928 ( .A(n55117), .B(n68355), .X(n39998) );
  nand_x1_sg U70929 ( .A(n55163), .B(n68354), .X(n39993) );
  nand_x1_sg U70930 ( .A(n55115), .B(n68353), .X(n39988) );
  nand_x1_sg U70931 ( .A(n55113), .B(n68352), .X(n39983) );
  nand_x1_sg U70932 ( .A(n55111), .B(n68351), .X(n39978) );
  nand_x1_sg U70933 ( .A(n55109), .B(n68350), .X(n39973) );
  nand_x1_sg U70934 ( .A(n55107), .B(n68349), .X(n39968) );
  nand_x1_sg U70935 ( .A(n55105), .B(n68348), .X(n39963) );
  nand_x1_sg U70936 ( .A(n55103), .B(n68347), .X(n39958) );
  nand_x1_sg U70937 ( .A(n55101), .B(n68346), .X(n39953) );
  nand_x1_sg U70938 ( .A(n55099), .B(n68345), .X(n39948) );
  nand_x1_sg U70939 ( .A(n55097), .B(n68344), .X(n39943) );
  nand_x1_sg U70940 ( .A(n55095), .B(n68343), .X(n39938) );
  nand_x1_sg U70941 ( .A(n55161), .B(n68342), .X(n39933) );
  nand_x1_sg U70942 ( .A(n55159), .B(n68341), .X(n39928) );
  nand_x1_sg U70943 ( .A(n55093), .B(n68340), .X(n39923) );
  nand_x1_sg U70944 ( .A(n55091), .B(n68339), .X(n39918) );
  nand_x1_sg U70945 ( .A(n55089), .B(n68338), .X(n39913) );
  nand_x1_sg U70946 ( .A(n55157), .B(n68337), .X(n39908) );
  nand_x1_sg U70947 ( .A(n22698), .B(n22471), .X(n22697) );
  nand_x1_sg U70948 ( .A(n57862), .B(n68573), .X(n22696) );
  nor_x1_sg U70949 ( .A(n57091), .B(n57113), .X(\filter_0/n8272 ) );
  nor_x1_sg U70950 ( .A(n57073), .B(n22395), .X(\shifter_0/n12760 ) );
  nor_x1_sg U70951 ( .A(n51547), .B(n22395), .X(\shifter_0/n12748 ) );
  nor_x1_sg U70952 ( .A(n57075), .B(n22395), .X(\shifter_0/n12736 ) );
  nor_x1_sg U70953 ( .A(n57077), .B(n22395), .X(\shifter_0/n12724 ) );
  nor_x1_sg U70954 ( .A(n51551), .B(n22395), .X(\shifter_0/n12712 ) );
  nor_x1_sg U70955 ( .A(n57083), .B(n22395), .X(\shifter_0/n12708 ) );
  nor_x1_sg U70956 ( .A(n57085), .B(n22395), .X(\shifter_0/n12704 ) );
  nor_x1_sg U70957 ( .A(n47759), .B(n22395), .X(\shifter_0/n12692 ) );
  nor_x1_sg U70958 ( .A(n51543), .B(n22395), .X(\shifter_0/n12688 ) );
  nor_x1_sg U70959 ( .A(n47773), .B(n26003), .X(\shifter_0/n10280 ) );
  nor_x1_sg U70960 ( .A(n51545), .B(n26003), .X(\shifter_0/n10268 ) );
  nor_x1_sg U70961 ( .A(n57071), .B(n26003), .X(\shifter_0/n10256 ) );
  nor_x1_sg U70962 ( .A(n57079), .B(n26003), .X(\shifter_0/n10244 ) );
  nor_x1_sg U70963 ( .A(n51553), .B(n26003), .X(\shifter_0/n10232 ) );
  nor_x1_sg U70964 ( .A(n57087), .B(n26003), .X(\shifter_0/n10228 ) );
  nor_x1_sg U70965 ( .A(n57089), .B(n26003), .X(\shifter_0/n10224 ) );
  nor_x1_sg U70966 ( .A(n51549), .B(n26003), .X(\shifter_0/n10212 ) );
  nor_x1_sg U70967 ( .A(n57081), .B(n26003), .X(\shifter_0/n10208 ) );
  nand_x1_sg U70968 ( .A(n26043), .B(n47343), .X(n26152) );
  nand_x1_sg U70969 ( .A(n26043), .B(n47345), .X(n26115) );
  nand_x1_sg U70970 ( .A(n26043), .B(n47347), .X(n26244) );
  nand_x1_sg U70971 ( .A(n26043), .B(n47349), .X(n26210) );
  nand_x1_sg U70972 ( .A(n47637), .B(n57453), .X(n24808) );
  nand_x1_sg U70973 ( .A(n47643), .B(n57450), .X(n24807) );
  nand_x1_sg U70974 ( .A(n47639), .B(n57453), .X(n24844) );
  nand_x1_sg U70975 ( .A(n47645), .B(n57450), .X(n24843) );
  nand_x1_sg U70976 ( .A(n51223), .B(n57453), .X(n24874) );
  nand_x1_sg U70977 ( .A(n51229), .B(n57450), .X(n24873) );
  nand_x1_sg U70978 ( .A(n51265), .B(n57453), .X(n24904) );
  nand_x1_sg U70979 ( .A(n51271), .B(n57450), .X(n24903) );
  nand_x1_sg U70980 ( .A(n56727), .B(n57453), .X(n24934) );
  nand_x1_sg U70981 ( .A(n56733), .B(n57450), .X(n24933) );
  nand_x1_sg U70982 ( .A(n47641), .B(n57453), .X(n24964) );
  nand_x1_sg U70983 ( .A(n47647), .B(n57450), .X(n24963) );
  nand_x1_sg U70984 ( .A(n51225), .B(n57453), .X(n24994) );
  nand_x1_sg U70985 ( .A(n51231), .B(n57450), .X(n24993) );
  nand_x1_sg U70986 ( .A(n56685), .B(n57453), .X(n25024) );
  nand_x1_sg U70987 ( .A(n56691), .B(n57450), .X(n25023) );
  nand_x1_sg U70988 ( .A(n51267), .B(n57453), .X(n25054) );
  nand_x1_sg U70989 ( .A(n51273), .B(n57450), .X(n25053) );
  nand_x1_sg U70990 ( .A(n56729), .B(n57453), .X(n25084) );
  nand_x1_sg U70991 ( .A(n56735), .B(n57450), .X(n25083) );
  nand_x1_sg U70992 ( .A(n51227), .B(n57453), .X(n25114) );
  nand_x1_sg U70993 ( .A(n51233), .B(n57450), .X(n25113) );
  nand_x1_sg U70994 ( .A(n56687), .B(n57453), .X(n25144) );
  nand_x1_sg U70995 ( .A(n56693), .B(n57450), .X(n25143) );
  nand_x1_sg U70996 ( .A(n51269), .B(n57453), .X(n25174) );
  nand_x1_sg U70997 ( .A(n51275), .B(n57450), .X(n25173) );
  nand_x1_sg U70998 ( .A(n56731), .B(n57451), .X(n25204) );
  nand_x1_sg U70999 ( .A(n56737), .B(n57450), .X(n25203) );
  nand_x1_sg U71000 ( .A(n51241), .B(n57451), .X(n25234) );
  nand_x1_sg U71001 ( .A(n51243), .B(n57450), .X(n25233) );
  nand_x1_sg U71002 ( .A(n56703), .B(n57453), .X(n25264) );
  nand_x1_sg U71003 ( .A(n56705), .B(n57450), .X(n25263) );
  nand_x1_sg U71004 ( .A(n47691), .B(n57453), .X(n25294) );
  nand_x1_sg U71005 ( .A(n47693), .B(n57450), .X(n25293) );
  nand_x1_sg U71006 ( .A(n51403), .B(n57453), .X(n25324) );
  nand_x1_sg U71007 ( .A(n51405), .B(n57450), .X(n25323) );
  nand_x1_sg U71008 ( .A(n56843), .B(n57453), .X(n25354) );
  nand_x1_sg U71009 ( .A(n56845), .B(n57450), .X(n25353) );
  nand_x1_sg U71010 ( .A(n56689), .B(n57453), .X(n25385) );
  nand_x1_sg U71011 ( .A(n56695), .B(n57450), .X(n25384) );
  nand_x1_sg U71012 ( .A(n47617), .B(n57453), .X(n25416) );
  nand_x1_sg U71013 ( .A(n47623), .B(n57450), .X(n25415) );
  nand_x1_sg U71014 ( .A(n47619), .B(n57453), .X(n25446) );
  nand_x1_sg U71015 ( .A(n47625), .B(n57450), .X(n25445) );
  nand_x1_sg U71016 ( .A(n51201), .B(n57453), .X(n25476) );
  nand_x1_sg U71017 ( .A(n51207), .B(n57450), .X(n25475) );
  nand_x1_sg U71018 ( .A(n51245), .B(n57452), .X(n25506) );
  nand_x1_sg U71019 ( .A(n51251), .B(n57450), .X(n25505) );
  nand_x1_sg U71020 ( .A(n56707), .B(n57452), .X(n25536) );
  nand_x1_sg U71021 ( .A(n56713), .B(n57450), .X(n25535) );
  nand_x1_sg U71022 ( .A(n47621), .B(n57453), .X(n25566) );
  nand_x1_sg U71023 ( .A(n47627), .B(n57450), .X(n25565) );
  nand_x1_sg U71024 ( .A(n51203), .B(n57453), .X(n25596) );
  nand_x1_sg U71025 ( .A(n51209), .B(n57450), .X(n25595) );
  nand_x1_sg U71026 ( .A(n56661), .B(n57453), .X(n25626) );
  nand_x1_sg U71027 ( .A(n56667), .B(n57450), .X(n25625) );
  nand_x1_sg U71028 ( .A(n51247), .B(n57453), .X(n25656) );
  nand_x1_sg U71029 ( .A(n51253), .B(n57450), .X(n25655) );
  nand_x1_sg U71030 ( .A(n56709), .B(n57453), .X(n25686) );
  nand_x1_sg U71031 ( .A(n56715), .B(n57450), .X(n25685) );
  nand_x1_sg U71032 ( .A(n51205), .B(n57453), .X(n25716) );
  nand_x1_sg U71033 ( .A(n51211), .B(n57450), .X(n25715) );
  nand_x1_sg U71034 ( .A(n56663), .B(n57453), .X(n25746) );
  nand_x1_sg U71035 ( .A(n56669), .B(n57450), .X(n25745) );
  nand_x1_sg U71036 ( .A(n51249), .B(n57453), .X(n25776) );
  nand_x1_sg U71037 ( .A(n51255), .B(n57450), .X(n25775) );
  nand_x1_sg U71038 ( .A(n56711), .B(n57453), .X(n25806) );
  nand_x1_sg U71039 ( .A(n56717), .B(n57450), .X(n25805) );
  nand_x1_sg U71040 ( .A(n51237), .B(n57453), .X(n25836) );
  nand_x1_sg U71041 ( .A(n51239), .B(n57450), .X(n25835) );
  nand_x1_sg U71042 ( .A(n56699), .B(n57453), .X(n25866) );
  nand_x1_sg U71043 ( .A(n56701), .B(n57450), .X(n25865) );
  nand_x1_sg U71044 ( .A(n47679), .B(n57453), .X(n25896) );
  nand_x1_sg U71045 ( .A(n47681), .B(n57450), .X(n25895) );
  nand_x1_sg U71046 ( .A(n51389), .B(n57453), .X(n25926) );
  nand_x1_sg U71047 ( .A(n51391), .B(n57450), .X(n25925) );
  nand_x1_sg U71048 ( .A(n56831), .B(n57453), .X(n25956) );
  nand_x1_sg U71049 ( .A(n56833), .B(n57450), .X(n25955) );
  nand_x1_sg U71050 ( .A(n56665), .B(n57453), .X(n25987) );
  nand_x1_sg U71051 ( .A(n56671), .B(n57450), .X(n25986) );
  nand_x1_sg U71052 ( .A(n47365), .B(n57857), .X(n24828) );
  nand_x1_sg U71053 ( .A(n47367), .B(n57857), .X(n24859) );
  nand_x1_sg U71054 ( .A(n56923), .B(n57857), .X(n24889) );
  nand_x1_sg U71055 ( .A(n47369), .B(n57857), .X(n24979) );
  nand_x1_sg U71056 ( .A(n47429), .B(n57857), .X(n25009) );
  nand_x1_sg U71057 ( .A(n56925), .B(n57857), .X(n25039) );
  nand_x1_sg U71058 ( .A(n47431), .B(n57857), .X(n25129) );
  nand_x1_sg U71059 ( .A(n56927), .B(n57857), .X(n25159) );
  nand_x1_sg U71060 ( .A(n47371), .B(n57857), .X(n25249) );
  nand_x1_sg U71061 ( .A(n47433), .B(n57857), .X(n25279) );
  nand_x1_sg U71062 ( .A(n56933), .B(n57857), .X(n25309) );
  nand_x1_sg U71063 ( .A(n47435), .B(n57857), .X(n25400) );
  nand_x1_sg U71064 ( .A(n47357), .B(n57857), .X(n25431) );
  nand_x1_sg U71065 ( .A(n47359), .B(n57857), .X(n25461) );
  nand_x1_sg U71066 ( .A(n56917), .B(n57857), .X(n25491) );
  nand_x1_sg U71067 ( .A(n47361), .B(n57857), .X(n25581) );
  nand_x1_sg U71068 ( .A(n47421), .B(n57857), .X(n25611) );
  nand_x1_sg U71069 ( .A(n56919), .B(n57857), .X(n25641) );
  nand_x1_sg U71070 ( .A(n47423), .B(n57857), .X(n25731) );
  nand_x1_sg U71071 ( .A(n56921), .B(n57857), .X(n25761) );
  nand_x1_sg U71072 ( .A(n47363), .B(n57857), .X(n25851) );
  nand_x1_sg U71073 ( .A(n47425), .B(n57857), .X(n25881) );
  nand_x1_sg U71074 ( .A(n56931), .B(n57101), .X(n25911) );
  nand_x1_sg U71075 ( .A(n47427), .B(n57857), .X(n26002) );
  nor_x1_sg U71076 ( .A(n57047), .B(n22395), .X(\shifter_0/n10204 ) );
  nor_x1_sg U71077 ( .A(n56987), .B(n22395), .X(\shifter_0/n12756 ) );
  nor_x1_sg U71078 ( .A(n56989), .B(n22395), .X(\shifter_0/n12752 ) );
  nor_x1_sg U71079 ( .A(n56991), .B(n22395), .X(\shifter_0/n12744 ) );
  nor_x1_sg U71080 ( .A(n56993), .B(n22395), .X(\shifter_0/n12740 ) );
  nor_x1_sg U71081 ( .A(n57005), .B(n22395), .X(\shifter_0/n12732 ) );
  nor_x1_sg U71082 ( .A(n57007), .B(n22395), .X(\shifter_0/n12728 ) );
  nor_x1_sg U71083 ( .A(n56999), .B(n22395), .X(\shifter_0/n12720 ) );
  nor_x1_sg U71084 ( .A(n56977), .B(n22395), .X(\shifter_0/n12716 ) );
  nor_x1_sg U71085 ( .A(n56973), .B(n22395), .X(\shifter_0/n12700 ) );
  nor_x1_sg U71086 ( .A(n56975), .B(n22395), .X(\shifter_0/n12696 ) );
  nor_x1_sg U71087 ( .A(n57045), .B(n26003), .X(\shifter_0/n10284 ) );
  nor_x1_sg U71088 ( .A(n56983), .B(n26003), .X(\shifter_0/n10276 ) );
  nor_x1_sg U71089 ( .A(n56985), .B(n26003), .X(\shifter_0/n10272 ) );
  nor_x1_sg U71090 ( .A(n56979), .B(n26003), .X(\shifter_0/n10264 ) );
  nor_x1_sg U71091 ( .A(n56981), .B(n26003), .X(\shifter_0/n10260 ) );
  nor_x1_sg U71092 ( .A(n57009), .B(n26003), .X(\shifter_0/n10252 ) );
  nor_x1_sg U71093 ( .A(n57011), .B(n26003), .X(\shifter_0/n10248 ) );
  nor_x1_sg U71094 ( .A(n57001), .B(n26003), .X(\shifter_0/n10240 ) );
  nor_x1_sg U71095 ( .A(n57003), .B(n26003), .X(\shifter_0/n10236 ) );
  nor_x1_sg U71096 ( .A(n56997), .B(n26003), .X(\shifter_0/n10220 ) );
  nor_x1_sg U71097 ( .A(n56995), .B(n26003), .X(\shifter_0/n10216 ) );
  nand_x1_sg U71098 ( .A(n47401), .B(n26117), .X(n26153) );
  nand_x1_sg U71099 ( .A(n47403), .B(n26117), .X(n26116) );
  nand_x1_sg U71100 ( .A(n47405), .B(n26117), .X(n26245) );
  nand_x1_sg U71101 ( .A(n47407), .B(n26117), .X(n26211) );
  nand_x1_sg U71102 ( .A(n47607), .B(n57328), .X(n58330) );
  nand_x1_sg U71103 ( .A(n47609), .B(n57328), .X(n58325) );
  nand_x1_sg U71104 ( .A(n51141), .B(n57328), .X(n58320) );
  nand_x1_sg U71105 ( .A(n47611), .B(n57328), .X(n58305) );
  nand_x1_sg U71106 ( .A(n51143), .B(n57328), .X(n58300) );
  nand_x1_sg U71107 ( .A(n55079), .B(n57328), .X(n58295) );
  nand_x1_sg U71108 ( .A(n51145), .B(n57328), .X(n58280) );
  nand_x1_sg U71109 ( .A(n55081), .B(n57328), .X(n58275) );
  nand_x1_sg U71110 ( .A(n51149), .B(n57328), .X(n58260) );
  nand_x1_sg U71111 ( .A(n55087), .B(n57328), .X(n58255) );
  nand_x1_sg U71112 ( .A(n55155), .B(n57328), .X(n58250) );
  nand_x1_sg U71113 ( .A(n55083), .B(n57328), .X(n58235) );
  nand_x1_sg U71114 ( .A(n47601), .B(n57328), .X(n58230) );
  nand_x1_sg U71115 ( .A(n47603), .B(n57328), .X(n58225) );
  nand_x1_sg U71116 ( .A(n51135), .B(n57328), .X(n58220) );
  nand_x1_sg U71117 ( .A(n47605), .B(n57328), .X(n58205) );
  nand_x1_sg U71118 ( .A(n51137), .B(n57328), .X(n58200) );
  nand_x1_sg U71119 ( .A(n55073), .B(n57328), .X(n58195) );
  nand_x1_sg U71120 ( .A(n51139), .B(n57328), .X(n58180) );
  nand_x1_sg U71121 ( .A(n55075), .B(n57326), .X(n58175) );
  nand_x1_sg U71122 ( .A(n51147), .B(n57327), .X(n58160) );
  nand_x1_sg U71123 ( .A(n55085), .B(n57328), .X(n58155) );
  nand_x1_sg U71124 ( .A(n55153), .B(n57328), .X(n58150) );
  nand_x1_sg U71125 ( .A(n55077), .B(n57328), .X(n58135) );
  nor_x1_sg U71126 ( .A(n24479), .B(n57949), .X(n58130) );
  nor_x1_sg U71127 ( .A(n24591), .B(n57949), .X(n58128) );
  nor_x1_sg U71128 ( .A(n55317), .B(n26249), .X(\filter_0/n8235 ) );
  nor_x1_sg U71129 ( .A(n55319), .B(n26249), .X(\filter_0/n10843 ) );
  nor_x1_sg U71130 ( .A(n55321), .B(n26249), .X(\filter_0/n10839 ) );
  nor_x1_sg U71131 ( .A(n55323), .B(n26249), .X(\filter_0/n10835 ) );
  nor_x1_sg U71132 ( .A(n55325), .B(n26249), .X(\filter_0/n10831 ) );
  nor_x1_sg U71133 ( .A(n55327), .B(n26249), .X(\filter_0/n10827 ) );
  nor_x1_sg U71134 ( .A(n55329), .B(n26249), .X(\filter_0/n10823 ) );
  nor_x1_sg U71135 ( .A(n55331), .B(n26249), .X(\filter_0/n10819 ) );
  nor_x1_sg U71136 ( .A(n55333), .B(n26249), .X(\filter_0/n10815 ) );
  nor_x1_sg U71137 ( .A(n55335), .B(n26249), .X(\filter_0/n10811 ) );
  nor_x1_sg U71138 ( .A(n55337), .B(n26249), .X(\filter_0/n10807 ) );
  nor_x1_sg U71139 ( .A(n55339), .B(n26249), .X(\filter_0/n10803 ) );
  nor_x1_sg U71140 ( .A(n55341), .B(n26249), .X(\filter_0/n10799 ) );
  nor_x1_sg U71141 ( .A(n55343), .B(n26249), .X(\filter_0/n10795 ) );
  nor_x1_sg U71142 ( .A(n55345), .B(n26249), .X(\filter_0/n10791 ) );
  nor_x1_sg U71143 ( .A(n55347), .B(n26249), .X(\filter_0/n10787 ) );
  nor_x1_sg U71144 ( .A(n55349), .B(n26249), .X(\filter_0/n10783 ) );
  nor_x1_sg U71145 ( .A(n55351), .B(n26249), .X(\filter_0/n10779 ) );
  nor_x1_sg U71146 ( .A(n55353), .B(n26249), .X(\filter_0/n10775 ) );
  nor_x1_sg U71147 ( .A(n55355), .B(n26249), .X(\filter_0/n10771 ) );
  nor_x1_sg U71148 ( .A(n55357), .B(n26250), .X(\filter_0/n10767 ) );
  nor_x1_sg U71149 ( .A(n55359), .B(n26250), .X(\filter_0/n10763 ) );
  nor_x1_sg U71150 ( .A(n55361), .B(n26250), .X(\filter_0/n10759 ) );
  nor_x1_sg U71151 ( .A(n55363), .B(n26250), .X(\filter_0/n10755 ) );
  nor_x1_sg U71152 ( .A(n55365), .B(n26250), .X(\filter_0/n10751 ) );
  nor_x1_sg U71153 ( .A(n55367), .B(n26250), .X(\filter_0/n10747 ) );
  nor_x1_sg U71154 ( .A(n55369), .B(n26250), .X(\filter_0/n10743 ) );
  nor_x1_sg U71155 ( .A(n55371), .B(n26250), .X(\filter_0/n10739 ) );
  nor_x1_sg U71156 ( .A(n55373), .B(n26250), .X(\filter_0/n10735 ) );
  nor_x1_sg U71157 ( .A(n55375), .B(n26250), .X(\filter_0/n10731 ) );
  nor_x1_sg U71158 ( .A(n55377), .B(n26250), .X(\filter_0/n10727 ) );
  nor_x1_sg U71159 ( .A(n55379), .B(n26250), .X(\filter_0/n10723 ) );
  nor_x1_sg U71160 ( .A(n55381), .B(n26250), .X(\filter_0/n10719 ) );
  nor_x1_sg U71161 ( .A(n55383), .B(n26250), .X(\filter_0/n10715 ) );
  nor_x1_sg U71162 ( .A(n55385), .B(n26250), .X(\filter_0/n10711 ) );
  nor_x1_sg U71163 ( .A(n55387), .B(n26250), .X(\filter_0/n10707 ) );
  nor_x1_sg U71164 ( .A(n55389), .B(n26250), .X(\filter_0/n10703 ) );
  nor_x1_sg U71165 ( .A(n55391), .B(n26250), .X(\filter_0/n10699 ) );
  nor_x1_sg U71166 ( .A(n55393), .B(n26250), .X(\filter_0/n10695 ) );
  nor_x1_sg U71167 ( .A(n55395), .B(n26250), .X(\filter_0/n10691 ) );
  nor_x1_sg U71168 ( .A(n55397), .B(n26251), .X(\filter_0/n10687 ) );
  nor_x1_sg U71169 ( .A(n55399), .B(n26251), .X(\filter_0/n10683 ) );
  nor_x1_sg U71170 ( .A(n55401), .B(n26251), .X(\filter_0/n10679 ) );
  nor_x1_sg U71171 ( .A(n55403), .B(n26251), .X(\filter_0/n10675 ) );
  nor_x1_sg U71172 ( .A(n55405), .B(n26251), .X(\filter_0/n10671 ) );
  nor_x1_sg U71173 ( .A(n55407), .B(n26251), .X(\filter_0/n10667 ) );
  nor_x1_sg U71174 ( .A(n55409), .B(n26251), .X(\filter_0/n10663 ) );
  nor_x1_sg U71175 ( .A(n55411), .B(n26251), .X(\filter_0/n10659 ) );
  nor_x1_sg U71176 ( .A(n55413), .B(n26251), .X(\filter_0/n10655 ) );
  nor_x1_sg U71177 ( .A(n55415), .B(n26251), .X(\filter_0/n10651 ) );
  nor_x1_sg U71178 ( .A(n55417), .B(n26251), .X(\filter_0/n10647 ) );
  nor_x1_sg U71179 ( .A(n55419), .B(n26251), .X(\filter_0/n10643 ) );
  nor_x1_sg U71180 ( .A(n55421), .B(n26251), .X(\filter_0/n10639 ) );
  nor_x1_sg U71181 ( .A(n55423), .B(n26251), .X(\filter_0/n10635 ) );
  nor_x1_sg U71182 ( .A(n55425), .B(n26251), .X(\filter_0/n10631 ) );
  nor_x1_sg U71183 ( .A(n55427), .B(n26251), .X(\filter_0/n10627 ) );
  nor_x1_sg U71184 ( .A(n55429), .B(n26251), .X(\filter_0/n10623 ) );
  nor_x1_sg U71185 ( .A(n55431), .B(n26251), .X(\filter_0/n10619 ) );
  nor_x1_sg U71186 ( .A(n55433), .B(n26251), .X(\filter_0/n10615 ) );
  nor_x1_sg U71187 ( .A(n55435), .B(n26251), .X(\filter_0/n10611 ) );
  nor_x1_sg U71188 ( .A(n55437), .B(n26252), .X(\filter_0/n10607 ) );
  nor_x1_sg U71189 ( .A(n55439), .B(n26252), .X(\filter_0/n10603 ) );
  nor_x1_sg U71190 ( .A(n55441), .B(n26252), .X(\filter_0/n10599 ) );
  nor_x1_sg U71191 ( .A(n55443), .B(n26252), .X(\filter_0/n10595 ) );
  nor_x1_sg U71192 ( .A(n55445), .B(n26252), .X(\filter_0/n10591 ) );
  nor_x1_sg U71193 ( .A(n55447), .B(n26252), .X(\filter_0/n10587 ) );
  nor_x1_sg U71194 ( .A(n55449), .B(n26252), .X(\filter_0/n10583 ) );
  nor_x1_sg U71195 ( .A(n55451), .B(n26252), .X(\filter_0/n10579 ) );
  nor_x1_sg U71196 ( .A(n55453), .B(n26252), .X(\filter_0/n10575 ) );
  nor_x1_sg U71197 ( .A(n55455), .B(n26252), .X(\filter_0/n10571 ) );
  nor_x1_sg U71198 ( .A(n55457), .B(n26252), .X(\filter_0/n10567 ) );
  nor_x1_sg U71199 ( .A(n55459), .B(n26252), .X(\filter_0/n10563 ) );
  nor_x1_sg U71200 ( .A(n55461), .B(n26252), .X(\filter_0/n10559 ) );
  nor_x1_sg U71201 ( .A(n55463), .B(n26252), .X(\filter_0/n10555 ) );
  nor_x1_sg U71202 ( .A(n55465), .B(n26252), .X(\filter_0/n10551 ) );
  nor_x1_sg U71203 ( .A(n55467), .B(n26252), .X(\filter_0/n10547 ) );
  nor_x1_sg U71204 ( .A(n55469), .B(n26252), .X(\filter_0/n10543 ) );
  nor_x1_sg U71205 ( .A(n55471), .B(n26252), .X(\filter_0/n10539 ) );
  nor_x1_sg U71206 ( .A(n55473), .B(n26252), .X(\filter_0/n10535 ) );
  nor_x1_sg U71207 ( .A(n55475), .B(n26252), .X(\filter_0/n10531 ) );
  nor_x1_sg U71208 ( .A(n55477), .B(n26253), .X(\filter_0/n10527 ) );
  nor_x1_sg U71209 ( .A(n55479), .B(n26253), .X(\filter_0/n10523 ) );
  nor_x1_sg U71210 ( .A(n55481), .B(n26253), .X(\filter_0/n10519 ) );
  nor_x1_sg U71211 ( .A(n55483), .B(n26253), .X(\filter_0/n10515 ) );
  nor_x1_sg U71212 ( .A(n55485), .B(n26253), .X(\filter_0/n10511 ) );
  nor_x1_sg U71213 ( .A(n55487), .B(n26253), .X(\filter_0/n10507 ) );
  nor_x1_sg U71214 ( .A(n55489), .B(n26253), .X(\filter_0/n10503 ) );
  nor_x1_sg U71215 ( .A(n55491), .B(n26253), .X(\filter_0/n10499 ) );
  nor_x1_sg U71216 ( .A(n55493), .B(n26253), .X(\filter_0/n10495 ) );
  nor_x1_sg U71217 ( .A(n55495), .B(n26253), .X(\filter_0/n10491 ) );
  nor_x1_sg U71218 ( .A(n55497), .B(n26253), .X(\filter_0/n10487 ) );
  nor_x1_sg U71219 ( .A(n55499), .B(n26253), .X(\filter_0/n10483 ) );
  nor_x1_sg U71220 ( .A(n55501), .B(n26253), .X(\filter_0/n10479 ) );
  nor_x1_sg U71221 ( .A(n55503), .B(n26253), .X(\filter_0/n10475 ) );
  nor_x1_sg U71222 ( .A(n55505), .B(n26253), .X(\filter_0/n10471 ) );
  nor_x1_sg U71223 ( .A(n55507), .B(n26253), .X(\filter_0/n10467 ) );
  nor_x1_sg U71224 ( .A(n55509), .B(n26253), .X(\filter_0/n10463 ) );
  nor_x1_sg U71225 ( .A(n55511), .B(n26253), .X(\filter_0/n10459 ) );
  nor_x1_sg U71226 ( .A(n55513), .B(n26253), .X(\filter_0/n10455 ) );
  nor_x1_sg U71227 ( .A(n55515), .B(n26253), .X(\filter_0/n10451 ) );
  nor_x1_sg U71228 ( .A(n55517), .B(n26254), .X(\filter_0/n10447 ) );
  nor_x1_sg U71229 ( .A(n55519), .B(n26254), .X(\filter_0/n10443 ) );
  nor_x1_sg U71230 ( .A(n55521), .B(n26254), .X(\filter_0/n10439 ) );
  nor_x1_sg U71231 ( .A(n55523), .B(n26254), .X(\filter_0/n10435 ) );
  nor_x1_sg U71232 ( .A(n55525), .B(n26254), .X(\filter_0/n10431 ) );
  nor_x1_sg U71233 ( .A(n55527), .B(n26254), .X(\filter_0/n10427 ) );
  nor_x1_sg U71234 ( .A(n55529), .B(n26254), .X(\filter_0/n10423 ) );
  nor_x1_sg U71235 ( .A(n55531), .B(n26254), .X(\filter_0/n10419 ) );
  nor_x1_sg U71236 ( .A(n55533), .B(n26254), .X(\filter_0/n10415 ) );
  nor_x1_sg U71237 ( .A(n55535), .B(n26254), .X(\filter_0/n10411 ) );
  nor_x1_sg U71238 ( .A(n55537), .B(n26254), .X(\filter_0/n10407 ) );
  nor_x1_sg U71239 ( .A(n55539), .B(n26254), .X(\filter_0/n10403 ) );
  nor_x1_sg U71240 ( .A(n55541), .B(n26254), .X(\filter_0/n10399 ) );
  nor_x1_sg U71241 ( .A(n55543), .B(n26254), .X(\filter_0/n10395 ) );
  nor_x1_sg U71242 ( .A(n55545), .B(n26254), .X(\filter_0/n10391 ) );
  nor_x1_sg U71243 ( .A(n55547), .B(n26254), .X(\filter_0/n10387 ) );
  nor_x1_sg U71244 ( .A(n55549), .B(n26254), .X(\filter_0/n10383 ) );
  nor_x1_sg U71245 ( .A(n55551), .B(n26254), .X(\filter_0/n10379 ) );
  nor_x1_sg U71246 ( .A(n55553), .B(n26254), .X(\filter_0/n10375 ) );
  nor_x1_sg U71247 ( .A(n55555), .B(n26254), .X(\filter_0/n10371 ) );
  nor_x1_sg U71248 ( .A(n55557), .B(n26255), .X(\filter_0/n10367 ) );
  nor_x1_sg U71249 ( .A(n55559), .B(n26255), .X(\filter_0/n10363 ) );
  nor_x1_sg U71250 ( .A(n55561), .B(n26255), .X(\filter_0/n10359 ) );
  nor_x1_sg U71251 ( .A(n55563), .B(n26255), .X(\filter_0/n10355 ) );
  nor_x1_sg U71252 ( .A(n55565), .B(n26255), .X(\filter_0/n10351 ) );
  nor_x1_sg U71253 ( .A(n55567), .B(n26255), .X(\filter_0/n10347 ) );
  nor_x1_sg U71254 ( .A(n55569), .B(n26255), .X(\filter_0/n10343 ) );
  nor_x1_sg U71255 ( .A(n55571), .B(n26255), .X(\filter_0/n10339 ) );
  nor_x1_sg U71256 ( .A(n55573), .B(n26255), .X(\filter_0/n10335 ) );
  nor_x1_sg U71257 ( .A(n55575), .B(n26255), .X(\filter_0/n10331 ) );
  nor_x1_sg U71258 ( .A(n55577), .B(n26255), .X(\filter_0/n10327 ) );
  nor_x1_sg U71259 ( .A(n55579), .B(n26255), .X(\filter_0/n10323 ) );
  nor_x1_sg U71260 ( .A(n55581), .B(n26255), .X(\filter_0/n10319 ) );
  nor_x1_sg U71261 ( .A(n55583), .B(n26255), .X(\filter_0/n10315 ) );
  nor_x1_sg U71262 ( .A(n55585), .B(n26255), .X(\filter_0/n10311 ) );
  nor_x1_sg U71263 ( .A(n55587), .B(n26255), .X(\filter_0/n10307 ) );
  nor_x1_sg U71264 ( .A(n55589), .B(n26255), .X(\filter_0/n10303 ) );
  nor_x1_sg U71265 ( .A(n55591), .B(n26255), .X(\filter_0/n10299 ) );
  nor_x1_sg U71266 ( .A(n55593), .B(n26255), .X(\filter_0/n10295 ) );
  nor_x1_sg U71267 ( .A(n55595), .B(n26255), .X(\filter_0/n10291 ) );
  nor_x1_sg U71268 ( .A(n55597), .B(n26256), .X(\filter_0/n10287 ) );
  nor_x1_sg U71269 ( .A(n55599), .B(n26256), .X(\filter_0/n10283 ) );
  nor_x1_sg U71270 ( .A(n55601), .B(n26256), .X(\filter_0/n10279 ) );
  nor_x1_sg U71271 ( .A(n55603), .B(n26256), .X(\filter_0/n10275 ) );
  nor_x1_sg U71272 ( .A(n55605), .B(n26256), .X(\filter_0/n10271 ) );
  nor_x1_sg U71273 ( .A(n55607), .B(n26256), .X(\filter_0/n10267 ) );
  nor_x1_sg U71274 ( .A(n55609), .B(n26256), .X(\filter_0/n10263 ) );
  nor_x1_sg U71275 ( .A(n55611), .B(n26256), .X(\filter_0/n10259 ) );
  nor_x1_sg U71276 ( .A(n55613), .B(n26256), .X(\filter_0/n10255 ) );
  nor_x1_sg U71277 ( .A(n55615), .B(n26256), .X(\filter_0/n10251 ) );
  nor_x1_sg U71278 ( .A(n55617), .B(n26256), .X(\filter_0/n10247 ) );
  nor_x1_sg U71279 ( .A(n55619), .B(n26256), .X(\filter_0/n10243 ) );
  nor_x1_sg U71280 ( .A(n55621), .B(n26256), .X(\filter_0/n10239 ) );
  nor_x1_sg U71281 ( .A(n55623), .B(n26256), .X(\filter_0/n10235 ) );
  nor_x1_sg U71282 ( .A(n55625), .B(n26256), .X(\filter_0/n10231 ) );
  nor_x1_sg U71283 ( .A(n55627), .B(n26256), .X(\filter_0/n10227 ) );
  nor_x1_sg U71284 ( .A(n55629), .B(n26256), .X(\filter_0/n10223 ) );
  nor_x1_sg U71285 ( .A(n55631), .B(n26256), .X(\filter_0/n10219 ) );
  nor_x1_sg U71286 ( .A(n55633), .B(n26256), .X(\filter_0/n10215 ) );
  nor_x1_sg U71287 ( .A(n55635), .B(n26256), .X(\filter_0/n10211 ) );
  nor_x1_sg U71288 ( .A(n55637), .B(n26257), .X(\filter_0/n10207 ) );
  nor_x1_sg U71289 ( .A(n55639), .B(n26257), .X(\filter_0/n10203 ) );
  nor_x1_sg U71290 ( .A(n55641), .B(n26257), .X(\filter_0/n10199 ) );
  nor_x1_sg U71291 ( .A(n55643), .B(n26257), .X(\filter_0/n10195 ) );
  nor_x1_sg U71292 ( .A(n55645), .B(n26257), .X(\filter_0/n10191 ) );
  nor_x1_sg U71293 ( .A(n55647), .B(n26257), .X(\filter_0/n10187 ) );
  nor_x1_sg U71294 ( .A(n55649), .B(n26257), .X(\filter_0/n10183 ) );
  nor_x1_sg U71295 ( .A(n55651), .B(n26257), .X(\filter_0/n10179 ) );
  nor_x1_sg U71296 ( .A(n55653), .B(n26257), .X(\filter_0/n10175 ) );
  nor_x1_sg U71297 ( .A(n55655), .B(n26257), .X(\filter_0/n10171 ) );
  nor_x1_sg U71298 ( .A(n55657), .B(n26257), .X(\filter_0/n10167 ) );
  nor_x1_sg U71299 ( .A(n55659), .B(n26257), .X(\filter_0/n10163 ) );
  nor_x1_sg U71300 ( .A(n55661), .B(n26257), .X(\filter_0/n10159 ) );
  nor_x1_sg U71301 ( .A(n55663), .B(n26257), .X(\filter_0/n10155 ) );
  nor_x1_sg U71302 ( .A(n55665), .B(n26257), .X(\filter_0/n10151 ) );
  nor_x1_sg U71303 ( .A(n55667), .B(n26257), .X(\filter_0/n10147 ) );
  nor_x1_sg U71304 ( .A(n55669), .B(n26257), .X(\filter_0/n10143 ) );
  nor_x1_sg U71305 ( .A(n55671), .B(n26257), .X(\filter_0/n10139 ) );
  nor_x1_sg U71306 ( .A(n55673), .B(n26257), .X(\filter_0/n10135 ) );
  nor_x1_sg U71307 ( .A(n55675), .B(n26257), .X(\filter_0/n10131 ) );
  nor_x1_sg U71308 ( .A(n55677), .B(n26259), .X(\filter_0/n10127 ) );
  nor_x1_sg U71309 ( .A(n55679), .B(n26259), .X(\filter_0/n10123 ) );
  nor_x1_sg U71310 ( .A(n55681), .B(n26259), .X(\filter_0/n10119 ) );
  nor_x1_sg U71311 ( .A(n55683), .B(n26259), .X(\filter_0/n10115 ) );
  nor_x1_sg U71312 ( .A(n55685), .B(n26259), .X(\filter_0/n10111 ) );
  nor_x1_sg U71313 ( .A(n55687), .B(n26259), .X(\filter_0/n10107 ) );
  nor_x1_sg U71314 ( .A(n55689), .B(n26259), .X(\filter_0/n10103 ) );
  nor_x1_sg U71315 ( .A(n55691), .B(n26259), .X(\filter_0/n10099 ) );
  nor_x1_sg U71316 ( .A(n55693), .B(n26259), .X(\filter_0/n10095 ) );
  nor_x1_sg U71317 ( .A(n55695), .B(n26259), .X(\filter_0/n10091 ) );
  nor_x1_sg U71318 ( .A(n55697), .B(n26259), .X(\filter_0/n10087 ) );
  nor_x1_sg U71319 ( .A(n55699), .B(n26259), .X(\filter_0/n10083 ) );
  nor_x1_sg U71320 ( .A(n55701), .B(n26259), .X(\filter_0/n10079 ) );
  nor_x1_sg U71321 ( .A(n55703), .B(n26259), .X(\filter_0/n10075 ) );
  nor_x1_sg U71322 ( .A(n55705), .B(n26259), .X(\filter_0/n10071 ) );
  nor_x1_sg U71323 ( .A(n55707), .B(n26259), .X(\filter_0/n10067 ) );
  nor_x1_sg U71324 ( .A(n55709), .B(n26259), .X(\filter_0/n10063 ) );
  nor_x1_sg U71325 ( .A(n55711), .B(n26259), .X(\filter_0/n10059 ) );
  nor_x1_sg U71326 ( .A(n55713), .B(n26259), .X(\filter_0/n10055 ) );
  nor_x1_sg U71327 ( .A(n55715), .B(n26259), .X(\filter_0/n10051 ) );
  nor_x1_sg U71328 ( .A(n55717), .B(n26006), .X(\filter_0/n10047 ) );
  nor_x1_sg U71329 ( .A(n55719), .B(n26006), .X(\filter_0/n10043 ) );
  nor_x1_sg U71330 ( .A(n55721), .B(n26006), .X(\filter_0/n10039 ) );
  nor_x1_sg U71331 ( .A(n55723), .B(n26006), .X(\filter_0/n10035 ) );
  nor_x1_sg U71332 ( .A(n55725), .B(n26006), .X(\filter_0/n10031 ) );
  nor_x1_sg U71333 ( .A(n55727), .B(n26006), .X(\filter_0/n10027 ) );
  nor_x1_sg U71334 ( .A(n55729), .B(n26006), .X(\filter_0/n10023 ) );
  nor_x1_sg U71335 ( .A(n55731), .B(n26006), .X(\filter_0/n10019 ) );
  nor_x1_sg U71336 ( .A(n55733), .B(n26006), .X(\filter_0/n10015 ) );
  nor_x1_sg U71337 ( .A(n55735), .B(n26006), .X(\filter_0/n10011 ) );
  nor_x1_sg U71338 ( .A(n55737), .B(n26006), .X(\filter_0/n10007 ) );
  nor_x1_sg U71339 ( .A(n55739), .B(n26006), .X(\filter_0/n10003 ) );
  nor_x1_sg U71340 ( .A(n55741), .B(n26006), .X(\filter_0/n9999 ) );
  nor_x1_sg U71341 ( .A(n55743), .B(n26006), .X(\filter_0/n9995 ) );
  nor_x1_sg U71342 ( .A(n55745), .B(n26006), .X(\filter_0/n9991 ) );
  nor_x1_sg U71343 ( .A(n55747), .B(n26006), .X(\filter_0/n9987 ) );
  nor_x1_sg U71344 ( .A(n55749), .B(n26006), .X(\filter_0/n9983 ) );
  nor_x1_sg U71345 ( .A(n55751), .B(n26006), .X(\filter_0/n9979 ) );
  nor_x1_sg U71346 ( .A(n55753), .B(n26006), .X(\filter_0/n9975 ) );
  nor_x1_sg U71347 ( .A(n55755), .B(n26006), .X(\filter_0/n9971 ) );
  nor_x1_sg U71348 ( .A(n55757), .B(n26007), .X(\filter_0/n9967 ) );
  nor_x1_sg U71349 ( .A(n55759), .B(n26007), .X(\filter_0/n9963 ) );
  nor_x1_sg U71350 ( .A(n55761), .B(n26007), .X(\filter_0/n9959 ) );
  nor_x1_sg U71351 ( .A(n55763), .B(n26007), .X(\filter_0/n9955 ) );
  nor_x1_sg U71352 ( .A(n55765), .B(n26007), .X(\filter_0/n9951 ) );
  nor_x1_sg U71353 ( .A(n55767), .B(n26007), .X(\filter_0/n9947 ) );
  nor_x1_sg U71354 ( .A(n55769), .B(n26007), .X(\filter_0/n9943 ) );
  nor_x1_sg U71355 ( .A(n55771), .B(n26007), .X(\filter_0/n9939 ) );
  nor_x1_sg U71356 ( .A(n55773), .B(n26007), .X(\filter_0/n9935 ) );
  nor_x1_sg U71357 ( .A(n55775), .B(n26007), .X(\filter_0/n9931 ) );
  nor_x1_sg U71358 ( .A(n55777), .B(n26007), .X(\filter_0/n9927 ) );
  nor_x1_sg U71359 ( .A(n55779), .B(n26007), .X(\filter_0/n9923 ) );
  nor_x1_sg U71360 ( .A(n55781), .B(n26007), .X(\filter_0/n9919 ) );
  nor_x1_sg U71361 ( .A(n55783), .B(n26007), .X(\filter_0/n9915 ) );
  nor_x1_sg U71362 ( .A(n55785), .B(n26007), .X(\filter_0/n9911 ) );
  nor_x1_sg U71363 ( .A(n55787), .B(n26007), .X(\filter_0/n9907 ) );
  nor_x1_sg U71364 ( .A(n55789), .B(n26007), .X(\filter_0/n9903 ) );
  nor_x1_sg U71365 ( .A(n55791), .B(n26007), .X(\filter_0/n9899 ) );
  nor_x1_sg U71366 ( .A(n55793), .B(n26007), .X(\filter_0/n9895 ) );
  nor_x1_sg U71367 ( .A(n55795), .B(n26007), .X(\filter_0/n9891 ) );
  nor_x1_sg U71368 ( .A(n55797), .B(n26009), .X(\filter_0/n9887 ) );
  nor_x1_sg U71369 ( .A(n55799), .B(n26009), .X(\filter_0/n9883 ) );
  nor_x1_sg U71370 ( .A(n55801), .B(n26009), .X(\filter_0/n9879 ) );
  nor_x1_sg U71371 ( .A(n55803), .B(n26009), .X(\filter_0/n9875 ) );
  nor_x1_sg U71372 ( .A(n55805), .B(n26009), .X(\filter_0/n9871 ) );
  nor_x1_sg U71373 ( .A(n55807), .B(n26009), .X(\filter_0/n9867 ) );
  nor_x1_sg U71374 ( .A(n55809), .B(n26009), .X(\filter_0/n9863 ) );
  nor_x1_sg U71375 ( .A(n55811), .B(n26009), .X(\filter_0/n9859 ) );
  nor_x1_sg U71376 ( .A(n55813), .B(n26009), .X(\filter_0/n9855 ) );
  nor_x1_sg U71377 ( .A(n55815), .B(n26009), .X(\filter_0/n9851 ) );
  nor_x1_sg U71378 ( .A(n55817), .B(n26009), .X(\filter_0/n9847 ) );
  nor_x1_sg U71379 ( .A(n55819), .B(n26009), .X(\filter_0/n9843 ) );
  nor_x1_sg U71380 ( .A(n55821), .B(n26009), .X(\filter_0/n9839 ) );
  nor_x1_sg U71381 ( .A(n55823), .B(n26009), .X(\filter_0/n9835 ) );
  nor_x1_sg U71382 ( .A(n55825), .B(n26009), .X(\filter_0/n9831 ) );
  nor_x1_sg U71383 ( .A(n55827), .B(n26009), .X(\filter_0/n9827 ) );
  nor_x1_sg U71384 ( .A(n55829), .B(n26009), .X(\filter_0/n9823 ) );
  nor_x1_sg U71385 ( .A(n55831), .B(n26009), .X(\filter_0/n9819 ) );
  nor_x1_sg U71386 ( .A(n55833), .B(n26009), .X(\filter_0/n9815 ) );
  nor_x1_sg U71387 ( .A(n55835), .B(n26009), .X(\filter_0/n9811 ) );
  nor_x1_sg U71388 ( .A(n55837), .B(n26011), .X(\filter_0/n9807 ) );
  nor_x1_sg U71389 ( .A(n55839), .B(n26011), .X(\filter_0/n9803 ) );
  nor_x1_sg U71390 ( .A(n55841), .B(n26011), .X(\filter_0/n9799 ) );
  nor_x1_sg U71391 ( .A(n55843), .B(n26011), .X(\filter_0/n9795 ) );
  nor_x1_sg U71392 ( .A(n55845), .B(n26011), .X(\filter_0/n9791 ) );
  nor_x1_sg U71393 ( .A(n55847), .B(n26011), .X(\filter_0/n9787 ) );
  nor_x1_sg U71394 ( .A(n55849), .B(n26011), .X(\filter_0/n9783 ) );
  nor_x1_sg U71395 ( .A(n55851), .B(n26011), .X(\filter_0/n9779 ) );
  nor_x1_sg U71396 ( .A(n55853), .B(n26011), .X(\filter_0/n9775 ) );
  nor_x1_sg U71397 ( .A(n55855), .B(n26011), .X(\filter_0/n9771 ) );
  nor_x1_sg U71398 ( .A(n55857), .B(n26011), .X(\filter_0/n9767 ) );
  nor_x1_sg U71399 ( .A(n55859), .B(n26011), .X(\filter_0/n9763 ) );
  nor_x1_sg U71400 ( .A(n55861), .B(n26011), .X(\filter_0/n9759 ) );
  nor_x1_sg U71401 ( .A(n55863), .B(n26011), .X(\filter_0/n9755 ) );
  nor_x1_sg U71402 ( .A(n55865), .B(n26011), .X(\filter_0/n9751 ) );
  nor_x1_sg U71403 ( .A(n55867), .B(n26011), .X(\filter_0/n9747 ) );
  nor_x1_sg U71404 ( .A(n55869), .B(n26011), .X(\filter_0/n9743 ) );
  nor_x1_sg U71405 ( .A(n55871), .B(n26011), .X(\filter_0/n9739 ) );
  nor_x1_sg U71406 ( .A(n55873), .B(n26011), .X(\filter_0/n9735 ) );
  nor_x1_sg U71407 ( .A(n55875), .B(n26011), .X(\filter_0/n9731 ) );
  nor_x1_sg U71408 ( .A(n55877), .B(n26013), .X(\filter_0/n9727 ) );
  nor_x1_sg U71409 ( .A(n55879), .B(n26013), .X(\filter_0/n9723 ) );
  nor_x1_sg U71410 ( .A(n55881), .B(n26013), .X(\filter_0/n9719 ) );
  nor_x1_sg U71411 ( .A(n55883), .B(n26013), .X(\filter_0/n9715 ) );
  nor_x1_sg U71412 ( .A(n55885), .B(n26013), .X(\filter_0/n9711 ) );
  nor_x1_sg U71413 ( .A(n55887), .B(n26013), .X(\filter_0/n9707 ) );
  nor_x1_sg U71414 ( .A(n55889), .B(n26013), .X(\filter_0/n9703 ) );
  nor_x1_sg U71415 ( .A(n55891), .B(n26013), .X(\filter_0/n9699 ) );
  nor_x1_sg U71416 ( .A(n55893), .B(n26013), .X(\filter_0/n9695 ) );
  nor_x1_sg U71417 ( .A(n55895), .B(n26013), .X(\filter_0/n9691 ) );
  nor_x1_sg U71418 ( .A(n55897), .B(n26013), .X(\filter_0/n9687 ) );
  nor_x1_sg U71419 ( .A(n55899), .B(n26013), .X(\filter_0/n9683 ) );
  nor_x1_sg U71420 ( .A(n55901), .B(n26013), .X(\filter_0/n9679 ) );
  nor_x1_sg U71421 ( .A(n55903), .B(n26013), .X(\filter_0/n9675 ) );
  nor_x1_sg U71422 ( .A(n55905), .B(n26013), .X(\filter_0/n9671 ) );
  nor_x1_sg U71423 ( .A(n55907), .B(n26013), .X(\filter_0/n9667 ) );
  nor_x1_sg U71424 ( .A(n55909), .B(n26013), .X(\filter_0/n9663 ) );
  nor_x1_sg U71425 ( .A(n55911), .B(n26013), .X(\filter_0/n9659 ) );
  nor_x1_sg U71426 ( .A(n55913), .B(n26013), .X(\filter_0/n9655 ) );
  nor_x1_sg U71427 ( .A(n55915), .B(n26013), .X(\filter_0/n9651 ) );
  nor_x1_sg U71428 ( .A(n55917), .B(n26015), .X(\filter_0/n9647 ) );
  nor_x1_sg U71429 ( .A(n55919), .B(n26015), .X(\filter_0/n9643 ) );
  nor_x1_sg U71430 ( .A(n55921), .B(n26015), .X(\filter_0/n9639 ) );
  nor_x1_sg U71431 ( .A(n55923), .B(n26015), .X(\filter_0/n9635 ) );
  nor_x1_sg U71432 ( .A(n55925), .B(n26015), .X(\filter_0/n9631 ) );
  nor_x1_sg U71433 ( .A(n55927), .B(n26015), .X(\filter_0/n9627 ) );
  nor_x1_sg U71434 ( .A(n55929), .B(n26015), .X(\filter_0/n9623 ) );
  nor_x1_sg U71435 ( .A(n55931), .B(n26015), .X(\filter_0/n9619 ) );
  nor_x1_sg U71436 ( .A(n55933), .B(n26015), .X(\filter_0/n9615 ) );
  nor_x1_sg U71437 ( .A(n55935), .B(n26015), .X(\filter_0/n9611 ) );
  nor_x1_sg U71438 ( .A(n55937), .B(n26015), .X(\filter_0/n9607 ) );
  nor_x1_sg U71439 ( .A(n55939), .B(n26015), .X(\filter_0/n9603 ) );
  nor_x1_sg U71440 ( .A(n55941), .B(n26015), .X(\filter_0/n9599 ) );
  nor_x1_sg U71441 ( .A(n55943), .B(n26015), .X(\filter_0/n9595 ) );
  nor_x1_sg U71442 ( .A(n55945), .B(n26015), .X(\filter_0/n9591 ) );
  nor_x1_sg U71443 ( .A(n55947), .B(n26015), .X(\filter_0/n9587 ) );
  nor_x1_sg U71444 ( .A(n55949), .B(n26015), .X(\filter_0/n9583 ) );
  nor_x1_sg U71445 ( .A(n55951), .B(n26015), .X(\filter_0/n9579 ) );
  nor_x1_sg U71446 ( .A(n55953), .B(n26015), .X(\filter_0/n9575 ) );
  nor_x1_sg U71447 ( .A(n55955), .B(n26015), .X(\filter_0/n9571 ) );
  nor_x1_sg U71448 ( .A(n55957), .B(n26016), .X(\filter_0/n9567 ) );
  nor_x1_sg U71449 ( .A(n55959), .B(n26016), .X(\filter_0/n9563 ) );
  nor_x1_sg U71450 ( .A(n55961), .B(n26016), .X(\filter_0/n9559 ) );
  nor_x1_sg U71451 ( .A(n55963), .B(n26016), .X(\filter_0/n9555 ) );
  nor_x1_sg U71452 ( .A(n55965), .B(n26016), .X(\filter_0/n9551 ) );
  nor_x1_sg U71453 ( .A(n55967), .B(n26016), .X(\filter_0/n9547 ) );
  nor_x1_sg U71454 ( .A(n55969), .B(n26016), .X(\filter_0/n9543 ) );
  nor_x1_sg U71455 ( .A(n55971), .B(n26016), .X(\filter_0/n9539 ) );
  nor_x1_sg U71456 ( .A(n55973), .B(n26016), .X(\filter_0/n9535 ) );
  nor_x1_sg U71457 ( .A(n55975), .B(n26016), .X(\filter_0/n9531 ) );
  nor_x1_sg U71458 ( .A(n55977), .B(n26016), .X(\filter_0/n9527 ) );
  nor_x1_sg U71459 ( .A(n55979), .B(n26016), .X(\filter_0/n9523 ) );
  nor_x1_sg U71460 ( .A(n55981), .B(n26016), .X(\filter_0/n9519 ) );
  nor_x1_sg U71461 ( .A(n55983), .B(n26016), .X(\filter_0/n9515 ) );
  nor_x1_sg U71462 ( .A(n55985), .B(n26016), .X(\filter_0/n9511 ) );
  nor_x1_sg U71463 ( .A(n55987), .B(n26016), .X(\filter_0/n9507 ) );
  nor_x1_sg U71464 ( .A(n55989), .B(n26016), .X(\filter_0/n9503 ) );
  nor_x1_sg U71465 ( .A(n55991), .B(n26016), .X(\filter_0/n9499 ) );
  nor_x1_sg U71466 ( .A(n55993), .B(n26016), .X(\filter_0/n9495 ) );
  nor_x1_sg U71467 ( .A(n55995), .B(n26016), .X(\filter_0/n9491 ) );
  nor_x1_sg U71468 ( .A(n55997), .B(n26018), .X(\filter_0/n9487 ) );
  nor_x1_sg U71469 ( .A(n55999), .B(n26018), .X(\filter_0/n9483 ) );
  nor_x1_sg U71470 ( .A(n56001), .B(n26018), .X(\filter_0/n9479 ) );
  nor_x1_sg U71471 ( .A(n56003), .B(n26018), .X(\filter_0/n9475 ) );
  nor_x1_sg U71472 ( .A(n56005), .B(n26018), .X(\filter_0/n9471 ) );
  nor_x1_sg U71473 ( .A(n56007), .B(n26018), .X(\filter_0/n9467 ) );
  nor_x1_sg U71474 ( .A(n56009), .B(n26018), .X(\filter_0/n9463 ) );
  nor_x1_sg U71475 ( .A(n56011), .B(n26018), .X(\filter_0/n9459 ) );
  nor_x1_sg U71476 ( .A(n56013), .B(n26018), .X(\filter_0/n9455 ) );
  nor_x1_sg U71477 ( .A(n56015), .B(n26018), .X(\filter_0/n9451 ) );
  nor_x1_sg U71478 ( .A(n56017), .B(n26018), .X(\filter_0/n9447 ) );
  nor_x1_sg U71479 ( .A(n56019), .B(n26018), .X(\filter_0/n9443 ) );
  nor_x1_sg U71480 ( .A(n56021), .B(n26018), .X(\filter_0/n9439 ) );
  nor_x1_sg U71481 ( .A(n56023), .B(n26018), .X(\filter_0/n9435 ) );
  nor_x1_sg U71482 ( .A(n56025), .B(n26018), .X(\filter_0/n9431 ) );
  nor_x1_sg U71483 ( .A(n56027), .B(n26018), .X(\filter_0/n9427 ) );
  nor_x1_sg U71484 ( .A(n56029), .B(n26018), .X(\filter_0/n9423 ) );
  nor_x1_sg U71485 ( .A(n56031), .B(n26018), .X(\filter_0/n9419 ) );
  nor_x1_sg U71486 ( .A(n56033), .B(n26018), .X(\filter_0/n9415 ) );
  nor_x1_sg U71487 ( .A(n56035), .B(n26018), .X(\filter_0/n9411 ) );
  nor_x1_sg U71488 ( .A(n56037), .B(n26020), .X(\filter_0/n9407 ) );
  nor_x1_sg U71489 ( .A(n56039), .B(n26020), .X(\filter_0/n9403 ) );
  nor_x1_sg U71490 ( .A(n56041), .B(n26020), .X(\filter_0/n9399 ) );
  nor_x1_sg U71491 ( .A(n56043), .B(n26020), .X(\filter_0/n9395 ) );
  nor_x1_sg U71492 ( .A(n56045), .B(n26020), .X(\filter_0/n9391 ) );
  nor_x1_sg U71493 ( .A(n56047), .B(n26020), .X(\filter_0/n9387 ) );
  nor_x1_sg U71494 ( .A(n56049), .B(n26020), .X(\filter_0/n9383 ) );
  nor_x1_sg U71495 ( .A(n56051), .B(n26020), .X(\filter_0/n9379 ) );
  nor_x1_sg U71496 ( .A(n56053), .B(n26020), .X(\filter_0/n9375 ) );
  nor_x1_sg U71497 ( .A(n56055), .B(n26020), .X(\filter_0/n9371 ) );
  nor_x1_sg U71498 ( .A(n56057), .B(n26020), .X(\filter_0/n9367 ) );
  nor_x1_sg U71499 ( .A(n56059), .B(n26020), .X(\filter_0/n9363 ) );
  nor_x1_sg U71500 ( .A(n56061), .B(n26020), .X(\filter_0/n9359 ) );
  nor_x1_sg U71501 ( .A(n56063), .B(n26020), .X(\filter_0/n9355 ) );
  nor_x1_sg U71502 ( .A(n56065), .B(n26020), .X(\filter_0/n9351 ) );
  nor_x1_sg U71503 ( .A(n56067), .B(n26020), .X(\filter_0/n9347 ) );
  nor_x1_sg U71504 ( .A(n56069), .B(n26020), .X(\filter_0/n9343 ) );
  nor_x1_sg U71505 ( .A(n56071), .B(n26020), .X(\filter_0/n9339 ) );
  nor_x1_sg U71506 ( .A(n56073), .B(n26020), .X(\filter_0/n9335 ) );
  nor_x1_sg U71507 ( .A(n56075), .B(n26020), .X(\filter_0/n9331 ) );
  nor_x1_sg U71508 ( .A(n56077), .B(n26022), .X(\filter_0/n9327 ) );
  nor_x1_sg U71509 ( .A(n56079), .B(n26022), .X(\filter_0/n9323 ) );
  nor_x1_sg U71510 ( .A(n56081), .B(n26022), .X(\filter_0/n9319 ) );
  nor_x1_sg U71511 ( .A(n56083), .B(n26022), .X(\filter_0/n9315 ) );
  nor_x1_sg U71512 ( .A(n56085), .B(n26022), .X(\filter_0/n9311 ) );
  nor_x1_sg U71513 ( .A(n56087), .B(n26022), .X(\filter_0/n9307 ) );
  nor_x1_sg U71514 ( .A(n56089), .B(n26022), .X(\filter_0/n9303 ) );
  nor_x1_sg U71515 ( .A(n56091), .B(n26022), .X(\filter_0/n9299 ) );
  nor_x1_sg U71516 ( .A(n56093), .B(n26022), .X(\filter_0/n9295 ) );
  nor_x1_sg U71517 ( .A(n56095), .B(n26022), .X(\filter_0/n9291 ) );
  nor_x1_sg U71518 ( .A(n56097), .B(n26022), .X(\filter_0/n9287 ) );
  nor_x1_sg U71519 ( .A(n56099), .B(n26022), .X(\filter_0/n9283 ) );
  nor_x1_sg U71520 ( .A(n56101), .B(n26022), .X(\filter_0/n9279 ) );
  nor_x1_sg U71521 ( .A(n56103), .B(n26022), .X(\filter_0/n9275 ) );
  nor_x1_sg U71522 ( .A(n56105), .B(n26022), .X(\filter_0/n9271 ) );
  nor_x1_sg U71523 ( .A(n56107), .B(n26022), .X(\filter_0/n9267 ) );
  nor_x1_sg U71524 ( .A(n56109), .B(n26022), .X(\filter_0/n9263 ) );
  nor_x1_sg U71525 ( .A(n56111), .B(n26022), .X(\filter_0/n9259 ) );
  nor_x1_sg U71526 ( .A(n56113), .B(n26022), .X(\filter_0/n9255 ) );
  nor_x1_sg U71527 ( .A(n56115), .B(n26022), .X(\filter_0/n9251 ) );
  nor_x1_sg U71528 ( .A(n56117), .B(n26024), .X(\filter_0/n9247 ) );
  nor_x1_sg U71529 ( .A(n56119), .B(n26024), .X(\filter_0/n9243 ) );
  nor_x1_sg U71530 ( .A(n56121), .B(n26024), .X(\filter_0/n9239 ) );
  nor_x1_sg U71531 ( .A(n56123), .B(n26024), .X(\filter_0/n9235 ) );
  nor_x1_sg U71532 ( .A(n56125), .B(n26024), .X(\filter_0/n9231 ) );
  nor_x1_sg U71533 ( .A(n56127), .B(n26024), .X(\filter_0/n9227 ) );
  nor_x1_sg U71534 ( .A(n56129), .B(n26024), .X(\filter_0/n9223 ) );
  nor_x1_sg U71535 ( .A(n56131), .B(n26024), .X(\filter_0/n9219 ) );
  nor_x1_sg U71536 ( .A(n56133), .B(n26024), .X(\filter_0/n9215 ) );
  nor_x1_sg U71537 ( .A(n56135), .B(n26024), .X(\filter_0/n9211 ) );
  nor_x1_sg U71538 ( .A(n56137), .B(n26024), .X(\filter_0/n9207 ) );
  nor_x1_sg U71539 ( .A(n56139), .B(n26024), .X(\filter_0/n9203 ) );
  nor_x1_sg U71540 ( .A(n56141), .B(n26024), .X(\filter_0/n9199 ) );
  nor_x1_sg U71541 ( .A(n56143), .B(n26024), .X(\filter_0/n9195 ) );
  nor_x1_sg U71542 ( .A(n56145), .B(n26024), .X(\filter_0/n9191 ) );
  nor_x1_sg U71543 ( .A(n56147), .B(n26024), .X(\filter_0/n9187 ) );
  nor_x1_sg U71544 ( .A(n56149), .B(n26024), .X(\filter_0/n9183 ) );
  nor_x1_sg U71545 ( .A(n56151), .B(n26024), .X(\filter_0/n9179 ) );
  nor_x1_sg U71546 ( .A(n56153), .B(n26024), .X(\filter_0/n9175 ) );
  nor_x1_sg U71547 ( .A(n56155), .B(n26024), .X(\filter_0/n9171 ) );
  nor_x1_sg U71548 ( .A(n56157), .B(n26025), .X(\filter_0/n9167 ) );
  nor_x1_sg U71549 ( .A(n56159), .B(n26025), .X(\filter_0/n9163 ) );
  nor_x1_sg U71550 ( .A(n56161), .B(n26025), .X(\filter_0/n9159 ) );
  nor_x1_sg U71551 ( .A(n56163), .B(n26025), .X(\filter_0/n9155 ) );
  nor_x1_sg U71552 ( .A(n56165), .B(n26025), .X(\filter_0/n9151 ) );
  nor_x1_sg U71553 ( .A(n56167), .B(n26025), .X(\filter_0/n9147 ) );
  nor_x1_sg U71554 ( .A(n56169), .B(n26025), .X(\filter_0/n9143 ) );
  nor_x1_sg U71555 ( .A(n56171), .B(n26025), .X(\filter_0/n9139 ) );
  nor_x1_sg U71556 ( .A(n56173), .B(n26025), .X(\filter_0/n9135 ) );
  nor_x1_sg U71557 ( .A(n56175), .B(n26025), .X(\filter_0/n9131 ) );
  nor_x1_sg U71558 ( .A(n56177), .B(n26025), .X(\filter_0/n9127 ) );
  nor_x1_sg U71559 ( .A(n56179), .B(n26025), .X(\filter_0/n9123 ) );
  nor_x1_sg U71560 ( .A(n56181), .B(n26025), .X(\filter_0/n9119 ) );
  nor_x1_sg U71561 ( .A(n56183), .B(n26025), .X(\filter_0/n9115 ) );
  nor_x1_sg U71562 ( .A(n56185), .B(n26025), .X(\filter_0/n9111 ) );
  nor_x1_sg U71563 ( .A(n56187), .B(n26025), .X(\filter_0/n9107 ) );
  nor_x1_sg U71564 ( .A(n56189), .B(n26025), .X(\filter_0/n9103 ) );
  nor_x1_sg U71565 ( .A(n56191), .B(n26025), .X(\filter_0/n9099 ) );
  nor_x1_sg U71566 ( .A(n56193), .B(n26025), .X(\filter_0/n9095 ) );
  nor_x1_sg U71567 ( .A(n56195), .B(n26025), .X(\filter_0/n9091 ) );
  nor_x1_sg U71568 ( .A(n56197), .B(n26026), .X(\filter_0/n9087 ) );
  nor_x1_sg U71569 ( .A(n56199), .B(n26026), .X(\filter_0/n9083 ) );
  nor_x1_sg U71570 ( .A(n56201), .B(n26026), .X(\filter_0/n9079 ) );
  nor_x1_sg U71571 ( .A(n56203), .B(n26026), .X(\filter_0/n9075 ) );
  nor_x1_sg U71572 ( .A(n56205), .B(n26026), .X(\filter_0/n9071 ) );
  nor_x1_sg U71573 ( .A(n56207), .B(n26026), .X(\filter_0/n9067 ) );
  nor_x1_sg U71574 ( .A(n56209), .B(n26026), .X(\filter_0/n9063 ) );
  nor_x1_sg U71575 ( .A(n56211), .B(n26026), .X(\filter_0/n9059 ) );
  nor_x1_sg U71576 ( .A(n56213), .B(n26026), .X(\filter_0/n9055 ) );
  nor_x1_sg U71577 ( .A(n56215), .B(n26026), .X(\filter_0/n9051 ) );
  nor_x1_sg U71578 ( .A(n56217), .B(n26026), .X(\filter_0/n9047 ) );
  nor_x1_sg U71579 ( .A(n56219), .B(n26026), .X(\filter_0/n9043 ) );
  nor_x1_sg U71580 ( .A(n56221), .B(n26026), .X(\filter_0/n9039 ) );
  nor_x1_sg U71581 ( .A(n56223), .B(n26026), .X(\filter_0/n9035 ) );
  nor_x1_sg U71582 ( .A(n56225), .B(n26026), .X(\filter_0/n9031 ) );
  nor_x1_sg U71583 ( .A(n56227), .B(n26026), .X(\filter_0/n9027 ) );
  nor_x1_sg U71584 ( .A(n56229), .B(n26026), .X(\filter_0/n9023 ) );
  nor_x1_sg U71585 ( .A(n56231), .B(n26026), .X(\filter_0/n9019 ) );
  nor_x1_sg U71586 ( .A(n56233), .B(n26026), .X(\filter_0/n9015 ) );
  nor_x1_sg U71587 ( .A(n56235), .B(n26026), .X(\filter_0/n9011 ) );
  nor_x1_sg U71588 ( .A(n56237), .B(n26027), .X(\filter_0/n9007 ) );
  nor_x1_sg U71589 ( .A(n56239), .B(n26027), .X(\filter_0/n9003 ) );
  nor_x1_sg U71590 ( .A(n56241), .B(n26027), .X(\filter_0/n8999 ) );
  nor_x1_sg U71591 ( .A(n56243), .B(n26027), .X(\filter_0/n8995 ) );
  nor_x1_sg U71592 ( .A(n56245), .B(n26027), .X(\filter_0/n8991 ) );
  nor_x1_sg U71593 ( .A(n56247), .B(n26027), .X(\filter_0/n8987 ) );
  nor_x1_sg U71594 ( .A(n56249), .B(n26027), .X(\filter_0/n8983 ) );
  nor_x1_sg U71595 ( .A(n56251), .B(n26027), .X(\filter_0/n8979 ) );
  nor_x1_sg U71596 ( .A(n56253), .B(n26027), .X(\filter_0/n8975 ) );
  nor_x1_sg U71597 ( .A(n56255), .B(n26027), .X(\filter_0/n8971 ) );
  nor_x1_sg U71598 ( .A(n56257), .B(n26027), .X(\filter_0/n8967 ) );
  nor_x1_sg U71599 ( .A(n56259), .B(n26027), .X(\filter_0/n8963 ) );
  nor_x1_sg U71600 ( .A(n56261), .B(n26027), .X(\filter_0/n8959 ) );
  nor_x1_sg U71601 ( .A(n56263), .B(n26027), .X(\filter_0/n8955 ) );
  nor_x1_sg U71602 ( .A(n56265), .B(n26027), .X(\filter_0/n8951 ) );
  nor_x1_sg U71603 ( .A(n56267), .B(n26027), .X(\filter_0/n8947 ) );
  nor_x1_sg U71604 ( .A(n56269), .B(n26027), .X(\filter_0/n8943 ) );
  nor_x1_sg U71605 ( .A(n56271), .B(n26027), .X(\filter_0/n8939 ) );
  nor_x1_sg U71606 ( .A(n56273), .B(n26027), .X(\filter_0/n8935 ) );
  nor_x1_sg U71607 ( .A(n56275), .B(n26027), .X(\filter_0/n8931 ) );
  nor_x1_sg U71608 ( .A(n56277), .B(n26028), .X(\filter_0/n8927 ) );
  nor_x1_sg U71609 ( .A(n56279), .B(n26028), .X(\filter_0/n8923 ) );
  nor_x1_sg U71610 ( .A(n56281), .B(n26028), .X(\filter_0/n8919 ) );
  nor_x1_sg U71611 ( .A(n56283), .B(n26028), .X(\filter_0/n8915 ) );
  nor_x1_sg U71612 ( .A(n56285), .B(n26028), .X(\filter_0/n8911 ) );
  nor_x1_sg U71613 ( .A(n56287), .B(n26028), .X(\filter_0/n8907 ) );
  nor_x1_sg U71614 ( .A(n56289), .B(n26028), .X(\filter_0/n8903 ) );
  nor_x1_sg U71615 ( .A(n56291), .B(n26028), .X(\filter_0/n8899 ) );
  nor_x1_sg U71616 ( .A(n56293), .B(n26028), .X(\filter_0/n8895 ) );
  nor_x1_sg U71617 ( .A(n56295), .B(n26028), .X(\filter_0/n8891 ) );
  nor_x1_sg U71618 ( .A(n56297), .B(n26028), .X(\filter_0/n8887 ) );
  nor_x1_sg U71619 ( .A(n56299), .B(n26028), .X(\filter_0/n8883 ) );
  nor_x1_sg U71620 ( .A(n56301), .B(n26028), .X(\filter_0/n8879 ) );
  nor_x1_sg U71621 ( .A(n56303), .B(n26028), .X(\filter_0/n8875 ) );
  nor_x1_sg U71622 ( .A(n56305), .B(n26028), .X(\filter_0/n8871 ) );
  nor_x1_sg U71623 ( .A(n56307), .B(n26028), .X(\filter_0/n8867 ) );
  nor_x1_sg U71624 ( .A(n56309), .B(n26028), .X(\filter_0/n8863 ) );
  nor_x1_sg U71625 ( .A(n56311), .B(n26028), .X(\filter_0/n8859 ) );
  nor_x1_sg U71626 ( .A(n56313), .B(n26028), .X(\filter_0/n8855 ) );
  nor_x1_sg U71627 ( .A(n56315), .B(n26028), .X(\filter_0/n8851 ) );
  nor_x1_sg U71628 ( .A(n56317), .B(n26029), .X(\filter_0/n8847 ) );
  nor_x1_sg U71629 ( .A(n56319), .B(n26029), .X(\filter_0/n8843 ) );
  nor_x1_sg U71630 ( .A(n56321), .B(n26029), .X(\filter_0/n8839 ) );
  nor_x1_sg U71631 ( .A(n56323), .B(n26029), .X(\filter_0/n8835 ) );
  nor_x1_sg U71632 ( .A(n56325), .B(n26029), .X(\filter_0/n8831 ) );
  nor_x1_sg U71633 ( .A(n56327), .B(n26029), .X(\filter_0/n8827 ) );
  nor_x1_sg U71634 ( .A(n56329), .B(n26029), .X(\filter_0/n8823 ) );
  nor_x1_sg U71635 ( .A(n56331), .B(n26029), .X(\filter_0/n8819 ) );
  nor_x1_sg U71636 ( .A(n56333), .B(n26029), .X(\filter_0/n8815 ) );
  nor_x1_sg U71637 ( .A(n56335), .B(n26029), .X(\filter_0/n8811 ) );
  nor_x1_sg U71638 ( .A(n56337), .B(n26029), .X(\filter_0/n8807 ) );
  nor_x1_sg U71639 ( .A(n56339), .B(n26029), .X(\filter_0/n8803 ) );
  nor_x1_sg U71640 ( .A(n56341), .B(n26029), .X(\filter_0/n8799 ) );
  nor_x1_sg U71641 ( .A(n56343), .B(n26029), .X(\filter_0/n8795 ) );
  nor_x1_sg U71642 ( .A(n56345), .B(n26029), .X(\filter_0/n8791 ) );
  nor_x1_sg U71643 ( .A(n56347), .B(n26029), .X(\filter_0/n8787 ) );
  nor_x1_sg U71644 ( .A(n56349), .B(n26029), .X(\filter_0/n8783 ) );
  nor_x1_sg U71645 ( .A(n56351), .B(n26029), .X(\filter_0/n8779 ) );
  nor_x1_sg U71646 ( .A(n56353), .B(n26029), .X(\filter_0/n8775 ) );
  nor_x1_sg U71647 ( .A(n56355), .B(n26029), .X(\filter_0/n8771 ) );
  nor_x1_sg U71648 ( .A(n56357), .B(n26030), .X(\filter_0/n8767 ) );
  nor_x1_sg U71649 ( .A(n56359), .B(n26030), .X(\filter_0/n8763 ) );
  nor_x1_sg U71650 ( .A(n56361), .B(n26030), .X(\filter_0/n8759 ) );
  nor_x1_sg U71651 ( .A(n56363), .B(n26030), .X(\filter_0/n8755 ) );
  nor_x1_sg U71652 ( .A(n56365), .B(n26030), .X(\filter_0/n8751 ) );
  nor_x1_sg U71653 ( .A(n56367), .B(n26030), .X(\filter_0/n8747 ) );
  nor_x1_sg U71654 ( .A(n56369), .B(n26030), .X(\filter_0/n8743 ) );
  nor_x1_sg U71655 ( .A(n56371), .B(n26030), .X(\filter_0/n8739 ) );
  nor_x1_sg U71656 ( .A(n56373), .B(n26030), .X(\filter_0/n8735 ) );
  nor_x1_sg U71657 ( .A(n56375), .B(n26030), .X(\filter_0/n8731 ) );
  nor_x1_sg U71658 ( .A(n56377), .B(n26030), .X(\filter_0/n8727 ) );
  nor_x1_sg U71659 ( .A(n56379), .B(n26030), .X(\filter_0/n8723 ) );
  nor_x1_sg U71660 ( .A(n56381), .B(n26030), .X(\filter_0/n8719 ) );
  nor_x1_sg U71661 ( .A(n56383), .B(n26030), .X(\filter_0/n8715 ) );
  nor_x1_sg U71662 ( .A(n56385), .B(n26030), .X(\filter_0/n8711 ) );
  nor_x1_sg U71663 ( .A(n56387), .B(n26030), .X(\filter_0/n8707 ) );
  nor_x1_sg U71664 ( .A(n56389), .B(n26030), .X(\filter_0/n8703 ) );
  nor_x1_sg U71665 ( .A(n56391), .B(n26030), .X(\filter_0/n8699 ) );
  nor_x1_sg U71666 ( .A(n56393), .B(n26030), .X(\filter_0/n8695 ) );
  nor_x1_sg U71667 ( .A(n56395), .B(n26030), .X(\filter_0/n8691 ) );
  nor_x1_sg U71668 ( .A(n56397), .B(n26031), .X(\filter_0/n8687 ) );
  nor_x1_sg U71669 ( .A(n56399), .B(n26031), .X(\filter_0/n8683 ) );
  nor_x1_sg U71670 ( .A(n56401), .B(n26031), .X(\filter_0/n8679 ) );
  nor_x1_sg U71671 ( .A(n56403), .B(n26031), .X(\filter_0/n8675 ) );
  nor_x1_sg U71672 ( .A(n56405), .B(n26031), .X(\filter_0/n8671 ) );
  nor_x1_sg U71673 ( .A(n56407), .B(n26031), .X(\filter_0/n8667 ) );
  nor_x1_sg U71674 ( .A(n56409), .B(n26031), .X(\filter_0/n8663 ) );
  nor_x1_sg U71675 ( .A(n56411), .B(n26031), .X(\filter_0/n8659 ) );
  nor_x1_sg U71676 ( .A(n56413), .B(n26031), .X(\filter_0/n8655 ) );
  nor_x1_sg U71677 ( .A(n56415), .B(n26031), .X(\filter_0/n8651 ) );
  nor_x1_sg U71678 ( .A(n56417), .B(n26031), .X(\filter_0/n8647 ) );
  nor_x1_sg U71679 ( .A(n56419), .B(n26031), .X(\filter_0/n8643 ) );
  nor_x1_sg U71680 ( .A(n56421), .B(n26031), .X(\filter_0/n8639 ) );
  nor_x1_sg U71681 ( .A(n56423), .B(n26031), .X(\filter_0/n8635 ) );
  nor_x1_sg U71682 ( .A(n56425), .B(n26031), .X(\filter_0/n8631 ) );
  nor_x1_sg U71683 ( .A(n56427), .B(n26031), .X(\filter_0/n8627 ) );
  nor_x1_sg U71684 ( .A(n56429), .B(n26031), .X(\filter_0/n8623 ) );
  nor_x1_sg U71685 ( .A(n56431), .B(n26031), .X(\filter_0/n8619 ) );
  nor_x1_sg U71686 ( .A(n56433), .B(n26031), .X(\filter_0/n8615 ) );
  nor_x1_sg U71687 ( .A(n56435), .B(n26031), .X(\filter_0/n8611 ) );
  nor_x1_sg U71688 ( .A(n56437), .B(n26032), .X(\filter_0/n8607 ) );
  nor_x1_sg U71689 ( .A(n56439), .B(n26032), .X(\filter_0/n8603 ) );
  nor_x1_sg U71690 ( .A(n56441), .B(n26032), .X(\filter_0/n8599 ) );
  nor_x1_sg U71691 ( .A(n56443), .B(n26032), .X(\filter_0/n8595 ) );
  nor_x1_sg U71692 ( .A(n56445), .B(n26032), .X(\filter_0/n8591 ) );
  nor_x1_sg U71693 ( .A(n56447), .B(n26032), .X(\filter_0/n8587 ) );
  nor_x1_sg U71694 ( .A(n56449), .B(n26032), .X(\filter_0/n8583 ) );
  nor_x1_sg U71695 ( .A(n56451), .B(n26032), .X(\filter_0/n8579 ) );
  nor_x1_sg U71696 ( .A(n56453), .B(n26032), .X(\filter_0/n8575 ) );
  nor_x1_sg U71697 ( .A(n56455), .B(n26032), .X(\filter_0/n8571 ) );
  nor_x1_sg U71698 ( .A(n56457), .B(n26032), .X(\filter_0/n8567 ) );
  nor_x1_sg U71699 ( .A(n56459), .B(n26032), .X(\filter_0/n8563 ) );
  nor_x1_sg U71700 ( .A(n56461), .B(n26032), .X(\filter_0/n8559 ) );
  nor_x1_sg U71701 ( .A(n56463), .B(n26032), .X(\filter_0/n8555 ) );
  nor_x1_sg U71702 ( .A(n56465), .B(n26032), .X(\filter_0/n8551 ) );
  nor_x1_sg U71703 ( .A(n56467), .B(n26032), .X(\filter_0/n8547 ) );
  nor_x1_sg U71704 ( .A(n56469), .B(n26032), .X(\filter_0/n8543 ) );
  nor_x1_sg U71705 ( .A(n56471), .B(n26032), .X(\filter_0/n8539 ) );
  nor_x1_sg U71706 ( .A(n56473), .B(n26032), .X(\filter_0/n8535 ) );
  nor_x1_sg U71707 ( .A(n56475), .B(n26032), .X(\filter_0/n8531 ) );
  nor_x1_sg U71708 ( .A(n56477), .B(n26035), .X(\filter_0/n8527 ) );
  nor_x1_sg U71709 ( .A(n56479), .B(n26035), .X(\filter_0/n8523 ) );
  nor_x1_sg U71710 ( .A(n56481), .B(n26035), .X(\filter_0/n8519 ) );
  nor_x1_sg U71711 ( .A(n56483), .B(n26035), .X(\filter_0/n8515 ) );
  nor_x1_sg U71712 ( .A(n56485), .B(n26035), .X(\filter_0/n8511 ) );
  nor_x1_sg U71713 ( .A(n56487), .B(n26035), .X(\filter_0/n8507 ) );
  nor_x1_sg U71714 ( .A(n56489), .B(n26035), .X(\filter_0/n8503 ) );
  nor_x1_sg U71715 ( .A(n56491), .B(n26035), .X(\filter_0/n8499 ) );
  nor_x1_sg U71716 ( .A(n56493), .B(n26035), .X(\filter_0/n8495 ) );
  nor_x1_sg U71717 ( .A(n56495), .B(n26035), .X(\filter_0/n8491 ) );
  nor_x1_sg U71718 ( .A(n56497), .B(n26035), .X(\filter_0/n8487 ) );
  nor_x1_sg U71719 ( .A(n56499), .B(n26035), .X(\filter_0/n8483 ) );
  nor_x1_sg U71720 ( .A(n56501), .B(n26035), .X(\filter_0/n8479 ) );
  nor_x1_sg U71721 ( .A(n56503), .B(n26035), .X(\filter_0/n8475 ) );
  nor_x1_sg U71722 ( .A(n56505), .B(n26035), .X(\filter_0/n8471 ) );
  nor_x1_sg U71723 ( .A(n56507), .B(n26035), .X(\filter_0/n8467 ) );
  nor_x1_sg U71724 ( .A(n56509), .B(n26035), .X(\filter_0/n8463 ) );
  nor_x1_sg U71725 ( .A(n56511), .B(n26035), .X(\filter_0/n8459 ) );
  nor_x1_sg U71726 ( .A(n56513), .B(n26035), .X(\filter_0/n8455 ) );
  nor_x1_sg U71727 ( .A(n56515), .B(n26035), .X(\filter_0/n8451 ) );
  nor_x1_sg U71728 ( .A(n56517), .B(n26037), .X(\filter_0/n8447 ) );
  nor_x1_sg U71729 ( .A(n56519), .B(n26037), .X(\filter_0/n8443 ) );
  nor_x1_sg U71730 ( .A(n56521), .B(n26037), .X(\filter_0/n8439 ) );
  nor_x1_sg U71731 ( .A(n56523), .B(n26037), .X(\filter_0/n8435 ) );
  nor_x1_sg U71732 ( .A(n56525), .B(n26037), .X(\filter_0/n8431 ) );
  nor_x1_sg U71733 ( .A(n56527), .B(n26037), .X(\filter_0/n8427 ) );
  nor_x1_sg U71734 ( .A(n56529), .B(n26037), .X(\filter_0/n8423 ) );
  nor_x1_sg U71735 ( .A(n56531), .B(n26037), .X(\filter_0/n8419 ) );
  nor_x1_sg U71736 ( .A(n56533), .B(n26037), .X(\filter_0/n8415 ) );
  nor_x1_sg U71737 ( .A(n56535), .B(n26037), .X(\filter_0/n8411 ) );
  nor_x1_sg U71738 ( .A(n56537), .B(n26037), .X(\filter_0/n8407 ) );
  nor_x1_sg U71739 ( .A(n56539), .B(n26037), .X(\filter_0/n8403 ) );
  nor_x1_sg U71740 ( .A(n56541), .B(n26037), .X(\filter_0/n8399 ) );
  nor_x1_sg U71741 ( .A(n56543), .B(n26037), .X(\filter_0/n8395 ) );
  nor_x1_sg U71742 ( .A(n56545), .B(n26037), .X(\filter_0/n8391 ) );
  nor_x1_sg U71743 ( .A(n56547), .B(n26037), .X(\filter_0/n8387 ) );
  nor_x1_sg U71744 ( .A(n56549), .B(n26037), .X(\filter_0/n8383 ) );
  nor_x1_sg U71745 ( .A(n56551), .B(n26037), .X(\filter_0/n8379 ) );
  nor_x1_sg U71746 ( .A(n56553), .B(n26037), .X(\filter_0/n8375 ) );
  nor_x1_sg U71747 ( .A(n56555), .B(n26037), .X(\filter_0/n8371 ) );
  nor_x1_sg U71748 ( .A(n56557), .B(n26038), .X(\filter_0/n8367 ) );
  nor_x1_sg U71749 ( .A(n56559), .B(n26038), .X(\filter_0/n8363 ) );
  nor_x1_sg U71750 ( .A(n56561), .B(n26038), .X(\filter_0/n8359 ) );
  nor_x1_sg U71751 ( .A(n56563), .B(n26038), .X(\filter_0/n8355 ) );
  nor_x1_sg U71752 ( .A(n56565), .B(n26038), .X(\filter_0/n8351 ) );
  nor_x1_sg U71753 ( .A(n56567), .B(n26038), .X(\filter_0/n8347 ) );
  nor_x1_sg U71754 ( .A(n56569), .B(n26038), .X(\filter_0/n8343 ) );
  nor_x1_sg U71755 ( .A(n56571), .B(n26038), .X(\filter_0/n8339 ) );
  nor_x1_sg U71756 ( .A(n56573), .B(n26038), .X(\filter_0/n8335 ) );
  nor_x1_sg U71757 ( .A(n56575), .B(n26038), .X(\filter_0/n8331 ) );
  nor_x1_sg U71758 ( .A(n56577), .B(n26038), .X(\filter_0/n8327 ) );
  nor_x1_sg U71759 ( .A(n56579), .B(n26038), .X(\filter_0/n8323 ) );
  nor_x1_sg U71760 ( .A(n56581), .B(n26038), .X(\filter_0/n8319 ) );
  nor_x1_sg U71761 ( .A(n56583), .B(n26038), .X(\filter_0/n8315 ) );
  nor_x1_sg U71762 ( .A(n56585), .B(n26038), .X(\filter_0/n8311 ) );
  nor_x1_sg U71763 ( .A(n56587), .B(n26038), .X(\filter_0/n8307 ) );
  nor_x1_sg U71764 ( .A(n56589), .B(n26038), .X(\filter_0/n8303 ) );
  nor_x1_sg U71765 ( .A(n56591), .B(n26038), .X(\filter_0/n8299 ) );
  nor_x1_sg U71766 ( .A(n56593), .B(n26038), .X(\filter_0/n8295 ) );
  nor_x1_sg U71767 ( .A(n56595), .B(n26038), .X(\filter_0/n8291 ) );
  nand_x4_sg U71768 ( .A(n26041), .B(n26042), .X(n26040) );
  nand_x1_sg U71769 ( .A(n26043), .B(n68373), .X(n26041) );
  nand_x1_sg U71770 ( .A(n57069), .B(n68374), .X(n26042) );
  nand_x4_sg U71771 ( .A(n26074), .B(n26075), .X(n26073) );
  nand_x1_sg U71772 ( .A(n56969), .B(n67576), .X(n26075) );
  nand_x1_sg U71773 ( .A(n26076), .B(n51523), .X(n26074) );
  nor_x1_sg U71774 ( .A(n47417), .B(n67575), .X(n26076) );
  nand_x4_sg U71775 ( .A(n26170), .B(n26171), .X(n26169) );
  nand_x1_sg U71776 ( .A(n56971), .B(n67582), .X(n26171) );
  nand_x1_sg U71777 ( .A(n26172), .B(n51525), .X(n26170) );
  nor_x1_sg U71778 ( .A(n47416), .B(n67581), .X(n26172) );
  nand_x4_sg U71779 ( .A(n26058), .B(n26059), .X(n26056) );
  nand_x1_sg U71780 ( .A(n67575), .B(n68380), .X(n26058) );
  nand_x1_sg U71781 ( .A(n51523), .B(n26060), .X(n26059) );
  nand_x4_sg U71782 ( .A(n26175), .B(n26176), .X(n26173) );
  nand_x1_sg U71783 ( .A(n67581), .B(n68386), .X(n26175) );
  nand_x1_sg U71784 ( .A(n51525), .B(n26177), .X(n26176) );
  nand_x4_sg U71785 ( .A(n23423), .B(n23424), .X(n23420) );
  nand_x1_sg U71786 ( .A(n47563), .B(n57320), .X(n23424) );
  nand_x1_sg U71787 ( .A(n47767), .B(n57318), .X(n23423) );
  nand_x4_sg U71788 ( .A(n23431), .B(n23432), .X(n23429) );
  nand_x1_sg U71789 ( .A(n47565), .B(n57320), .X(n23432) );
  nand_x1_sg U71790 ( .A(n47769), .B(n57318), .X(n23431) );
  nand_x4_sg U71791 ( .A(n23437), .B(n23438), .X(n23435) );
  nand_x1_sg U71792 ( .A(n56877), .B(n57320), .X(n23438) );
  nand_x1_sg U71793 ( .A(n51535), .B(n57318), .X(n23437) );
  nand_x4_sg U71794 ( .A(n23455), .B(n23456), .X(n23453) );
  nand_x1_sg U71795 ( .A(n47567), .B(n57320), .X(n23456) );
  nand_x1_sg U71796 ( .A(n47771), .B(n57318), .X(n23455) );
  nand_x4_sg U71797 ( .A(n23461), .B(n23462), .X(n23459) );
  nand_x1_sg U71798 ( .A(n56879), .B(n57320), .X(n23462) );
  nand_x1_sg U71799 ( .A(n51537), .B(n57318), .X(n23461) );
  nand_x4_sg U71800 ( .A(n23467), .B(n23468), .X(n23465) );
  nand_x1_sg U71801 ( .A(n51433), .B(n57320), .X(n23468) );
  nand_x1_sg U71802 ( .A(n57057), .B(n57318), .X(n23467) );
  nand_x4_sg U71803 ( .A(n23485), .B(n23486), .X(n23483) );
  nand_x1_sg U71804 ( .A(n56881), .B(n57320), .X(n23486) );
  nand_x1_sg U71805 ( .A(n51539), .B(n57318), .X(n23485) );
  nand_x4_sg U71806 ( .A(n23491), .B(n23492), .X(n23489) );
  nand_x1_sg U71807 ( .A(n51435), .B(n57320), .X(n23492) );
  nand_x1_sg U71808 ( .A(n57059), .B(n57318), .X(n23491) );
  nand_x4_sg U71809 ( .A(n23509), .B(n23510), .X(n23507) );
  nand_x1_sg U71810 ( .A(n56883), .B(n57320), .X(n23510) );
  nand_x1_sg U71811 ( .A(n51541), .B(n57318), .X(n23509) );
  nand_x4_sg U71812 ( .A(n23515), .B(n23516), .X(n23513) );
  nand_x1_sg U71813 ( .A(n51437), .B(n57320), .X(n23516) );
  nand_x1_sg U71814 ( .A(n57061), .B(n57318), .X(n23515) );
  nand_x4_sg U71815 ( .A(n23521), .B(n23522), .X(n23519) );
  nand_x1_sg U71816 ( .A(n47571), .B(n57320), .X(n23522) );
  nand_x1_sg U71817 ( .A(n57067), .B(n57318), .X(n23521) );
  nand_x4_sg U71818 ( .A(n23550), .B(n23551), .X(n23537) );
  nand_x1_sg U71819 ( .A(n51439), .B(n57320), .X(n23551) );
  nand_x1_sg U71820 ( .A(n57063), .B(n57318), .X(n23550) );
  nand_x4_sg U71821 ( .A(n23557), .B(n23558), .X(n23554) );
  nand_x1_sg U71822 ( .A(n47557), .B(n57320), .X(n23558) );
  nand_x1_sg U71823 ( .A(n47761), .B(n57318), .X(n23557) );
  nand_x4_sg U71824 ( .A(n23563), .B(n23564), .X(n23561) );
  nand_x1_sg U71825 ( .A(n47559), .B(n57320), .X(n23564) );
  nand_x1_sg U71826 ( .A(n47763), .B(n57318), .X(n23563) );
  nand_x4_sg U71827 ( .A(n23569), .B(n23570), .X(n23567) );
  nand_x1_sg U71828 ( .A(n56869), .B(n57320), .X(n23570) );
  nand_x1_sg U71829 ( .A(n51527), .B(n57318), .X(n23569) );
  nand_x4_sg U71830 ( .A(n23587), .B(n23588), .X(n23585) );
  nand_x1_sg U71831 ( .A(n47561), .B(n57320), .X(n23588) );
  nand_x1_sg U71832 ( .A(n47765), .B(n57318), .X(n23587) );
  nand_x4_sg U71833 ( .A(n23593), .B(n23594), .X(n23591) );
  nand_x1_sg U71834 ( .A(n56871), .B(n57320), .X(n23594) );
  nand_x1_sg U71835 ( .A(n51529), .B(n57318), .X(n23593) );
  nand_x4_sg U71836 ( .A(n23599), .B(n23600), .X(n23597) );
  nand_x1_sg U71837 ( .A(n51425), .B(n57320), .X(n23600) );
  nand_x1_sg U71838 ( .A(n57049), .B(n57318), .X(n23599) );
  nand_x4_sg U71839 ( .A(n23617), .B(n23618), .X(n23615) );
  nand_x1_sg U71840 ( .A(n56873), .B(n57320), .X(n23618) );
  nand_x1_sg U71841 ( .A(n51531), .B(n57318), .X(n23617) );
  nand_x4_sg U71842 ( .A(n23623), .B(n23624), .X(n23621) );
  nand_x1_sg U71843 ( .A(n51427), .B(n57320), .X(n23624) );
  nand_x1_sg U71844 ( .A(n57051), .B(n57318), .X(n23623) );
  nand_x4_sg U71845 ( .A(n23641), .B(n23642), .X(n23639) );
  nand_x1_sg U71846 ( .A(n56875), .B(n58388), .X(n23642) );
  nand_x1_sg U71847 ( .A(n51533), .B(n58387), .X(n23641) );
  nand_x4_sg U71848 ( .A(n23647), .B(n23648), .X(n23645) );
  nand_x1_sg U71849 ( .A(n51429), .B(n57320), .X(n23648) );
  nand_x1_sg U71850 ( .A(n57053), .B(n57318), .X(n23647) );
  nand_x4_sg U71851 ( .A(n23653), .B(n23654), .X(n23651) );
  nand_x1_sg U71852 ( .A(n47569), .B(n57320), .X(n23654) );
  nand_x1_sg U71853 ( .A(n57065), .B(n57318), .X(n23653) );
  nand_x4_sg U71854 ( .A(n23681), .B(n23682), .X(n23669) );
  nand_x1_sg U71855 ( .A(n51431), .B(n57320), .X(n23682) );
  nand_x1_sg U71856 ( .A(n57055), .B(n57318), .X(n23681) );
  nand_x1_sg U71857 ( .A(n57109), .B(n53589), .X(n26147) );
  nand_x1_sg U71858 ( .A(n57106), .B(n53585), .X(n26146) );
  nand_x1_sg U71859 ( .A(n57111), .B(n53587), .X(n26149) );
  nand_x1_sg U71860 ( .A(n57109), .B(n53603), .X(n26108) );
  nand_x1_sg U71861 ( .A(n57106), .B(n53599), .X(n26107) );
  nand_x1_sg U71862 ( .A(n57111), .B(n53601), .X(n26110) );
  nand_x1_sg U71863 ( .A(n57109), .B(n53617), .X(n26239) );
  nand_x1_sg U71864 ( .A(n57106), .B(n53613), .X(n26238) );
  nand_x1_sg U71865 ( .A(n57111), .B(n53615), .X(n26241) );
  nand_x1_sg U71866 ( .A(n57109), .B(n53631), .X(n26205) );
  nand_x1_sg U71867 ( .A(n57106), .B(n53627), .X(n26204) );
  nand_x1_sg U71868 ( .A(n57111), .B(n53629), .X(n26207) );
  nand_x4_sg U71869 ( .A(n26070), .B(n26071), .X(n26069) );
  nand_x1_sg U71870 ( .A(n26066), .B(n67528), .X(n26070) );
  nand_x1_sg U71871 ( .A(n47441), .B(n67576), .X(n26071) );
  nand_x4_sg U71872 ( .A(n26166), .B(n26167), .X(n26165) );
  nand_x1_sg U71873 ( .A(n26162), .B(n67525), .X(n26166) );
  nand_x1_sg U71874 ( .A(n47443), .B(n67582), .X(n26167) );
  nand_x1_sg U71875 ( .A(n26113), .B(n53591), .X(n26151) );
  nand_x1_sg U71876 ( .A(n26113), .B(n53605), .X(n26112) );
  nand_x1_sg U71877 ( .A(n26113), .B(n53619), .X(n26243) );
  nand_x1_sg U71878 ( .A(n26113), .B(n53633), .X(n26209) );
  nand_x1_sg U71879 ( .A(n47563), .B(n57949), .X(n58328) );
  nand_x1_sg U71880 ( .A(n47767), .B(n57929), .X(n58329) );
  nand_x1_sg U71881 ( .A(n47565), .B(n57949), .X(n58323) );
  nand_x1_sg U71882 ( .A(n47769), .B(n57929), .X(n58324) );
  nand_x1_sg U71883 ( .A(n56877), .B(n57949), .X(n58318) );
  nand_x1_sg U71884 ( .A(n51535), .B(n57930), .X(n58319) );
  nand_x1_sg U71885 ( .A(n47567), .B(n57949), .X(n58303) );
  nand_x1_sg U71886 ( .A(n47771), .B(n57951), .X(n58304) );
  nand_x1_sg U71887 ( .A(n56879), .B(n57949), .X(n58298) );
  nand_x1_sg U71888 ( .A(n51537), .B(n57926), .X(n58299) );
  nand_x1_sg U71889 ( .A(n51433), .B(n57949), .X(n58293) );
  nand_x1_sg U71890 ( .A(n57057), .B(n57951), .X(n58294) );
  nand_x1_sg U71891 ( .A(n56881), .B(n57949), .X(n58278) );
  nand_x1_sg U71892 ( .A(n51539), .B(n57931), .X(n58279) );
  nand_x1_sg U71893 ( .A(n51435), .B(n57949), .X(n58273) );
  nand_x1_sg U71894 ( .A(n57059), .B(n57932), .X(n58274) );
  nand_x1_sg U71895 ( .A(n56883), .B(n57949), .X(n58258) );
  nand_x1_sg U71896 ( .A(n51541), .B(n57940), .X(n58259) );
  nand_x1_sg U71897 ( .A(n51437), .B(n57949), .X(n58253) );
  nand_x1_sg U71898 ( .A(n57061), .B(n57933), .X(n58254) );
  nand_x1_sg U71899 ( .A(n47571), .B(n57949), .X(n58248) );
  nand_x1_sg U71900 ( .A(n57067), .B(n57933), .X(n58249) );
  nand_x1_sg U71901 ( .A(n51439), .B(n57949), .X(n58233) );
  nand_x1_sg U71902 ( .A(n57063), .B(n57934), .X(n58234) );
  nand_x1_sg U71903 ( .A(n47557), .B(n57949), .X(n58228) );
  nand_x1_sg U71904 ( .A(n47761), .B(n57934), .X(n58229) );
  nand_x1_sg U71905 ( .A(n47559), .B(n57949), .X(n58223) );
  nand_x1_sg U71906 ( .A(n47763), .B(n57935), .X(n58224) );
  nand_x1_sg U71907 ( .A(n56869), .B(n57949), .X(n58218) );
  nand_x1_sg U71908 ( .A(n51527), .B(n57935), .X(n58219) );
  nand_x1_sg U71909 ( .A(n47561), .B(n57949), .X(n58203) );
  nand_x1_sg U71910 ( .A(n47765), .B(n57936), .X(n58204) );
  nand_x1_sg U71911 ( .A(n56871), .B(n57949), .X(n58198) );
  nand_x1_sg U71912 ( .A(n51529), .B(n57936), .X(n58199) );
  nand_x1_sg U71913 ( .A(n51425), .B(n57949), .X(n58193) );
  nand_x1_sg U71914 ( .A(n57049), .B(n57937), .X(n58194) );
  nand_x1_sg U71915 ( .A(n56873), .B(n57949), .X(n58178) );
  nand_x1_sg U71916 ( .A(n51531), .B(n57938), .X(n58179) );
  nand_x1_sg U71917 ( .A(n51427), .B(n57949), .X(n58173) );
  nand_x1_sg U71918 ( .A(n57051), .B(n57938), .X(n58174) );
  nand_x1_sg U71919 ( .A(n56875), .B(n57949), .X(n58158) );
  nand_x1_sg U71920 ( .A(n51533), .B(n57939), .X(n58159) );
  nand_x1_sg U71921 ( .A(n51429), .B(n57949), .X(n58153) );
  nand_x1_sg U71922 ( .A(n57053), .B(n57939), .X(n58154) );
  nand_x1_sg U71923 ( .A(n47569), .B(n57949), .X(n58148) );
  nand_x1_sg U71924 ( .A(n57065), .B(n57940), .X(n58149) );
  nand_x1_sg U71925 ( .A(n51431), .B(n57949), .X(n58133) );
  nand_x1_sg U71926 ( .A(n57055), .B(n57941), .X(n58134) );
  nand_x1_sg U71927 ( .A(n47685), .B(n57349), .X(n24822) );
  nand_x1_sg U71928 ( .A(n47687), .B(n57348), .X(n24853) );
  nand_x1_sg U71929 ( .A(n51395), .B(n57348), .X(n24883) );
  nand_x1_sg U71930 ( .A(n51337), .B(n57348), .X(n24913) );
  nand_x1_sg U71931 ( .A(n56785), .B(n57348), .X(n24943) );
  nand_x1_sg U71932 ( .A(n47689), .B(n57349), .X(n24973) );
  nand_x1_sg U71933 ( .A(n51397), .B(n57349), .X(n25003) );
  nand_x1_sg U71934 ( .A(n56837), .B(n57348), .X(n25033) );
  nand_x1_sg U71935 ( .A(n51339), .B(n57348), .X(n25063) );
  nand_x1_sg U71936 ( .A(n56787), .B(n57349), .X(n25093) );
  nand_x1_sg U71937 ( .A(n51399), .B(n57348), .X(n25123) );
  nand_x1_sg U71938 ( .A(n56839), .B(n57349), .X(n25153) );
  nand_x1_sg U71939 ( .A(n51341), .B(n57348), .X(n25183) );
  nand_x1_sg U71940 ( .A(n56789), .B(n57349), .X(n25213) );
  nand_x1_sg U71941 ( .A(n51401), .B(n57348), .X(n25243) );
  nand_x1_sg U71942 ( .A(n56841), .B(n57349), .X(n25273) );
  nand_x1_sg U71943 ( .A(n56867), .B(n57348), .X(n25303) );
  nand_x1_sg U71944 ( .A(n47697), .B(n57348), .X(n25333) );
  nand_x1_sg U71945 ( .A(n51409), .B(n57349), .X(n25363) );
  nand_x1_sg U71946 ( .A(n56849), .B(n57349), .X(n25394) );
  nand_x1_sg U71947 ( .A(n47673), .B(n57348), .X(n25425) );
  nand_x1_sg U71948 ( .A(n47675), .B(n57349), .X(n25455) );
  nand_x1_sg U71949 ( .A(n51381), .B(n57348), .X(n25485) );
  nand_x1_sg U71950 ( .A(n51331), .B(n57349), .X(n25515) );
  nand_x1_sg U71951 ( .A(n56779), .B(n57348), .X(n25545) );
  nand_x1_sg U71952 ( .A(n47677), .B(n57348), .X(n25575) );
  nand_x1_sg U71953 ( .A(n51383), .B(n57348), .X(n25605) );
  nand_x1_sg U71954 ( .A(n56825), .B(n57348), .X(n25635) );
  nand_x1_sg U71955 ( .A(n51333), .B(n57349), .X(n25665) );
  nand_x1_sg U71956 ( .A(n56781), .B(n57348), .X(n25695) );
  nand_x1_sg U71957 ( .A(n51385), .B(n57348), .X(n25725) );
  nand_x1_sg U71958 ( .A(n56827), .B(n57348), .X(n25755) );
  nand_x1_sg U71959 ( .A(n51335), .B(n57349), .X(n25785) );
  nand_x1_sg U71960 ( .A(n56783), .B(n57348), .X(n25815) );
  nand_x1_sg U71961 ( .A(n51387), .B(n57348), .X(n25845) );
  nand_x1_sg U71962 ( .A(n56829), .B(n57348), .X(n25875) );
  nand_x1_sg U71963 ( .A(n56865), .B(n57348), .X(n25905) );
  nand_x1_sg U71964 ( .A(n47695), .B(n57348), .X(n25935) );
  nand_x1_sg U71965 ( .A(n51407), .B(n57348), .X(n25965) );
  nand_x1_sg U71966 ( .A(n56847), .B(n57348), .X(n25996) );
  nand_x4_sg U71967 ( .A(n23443), .B(n23444), .X(n23441) );
  nand_x1_sg U71968 ( .A(n47715), .B(n57320), .X(n23444) );
  nand_x1_sg U71969 ( .A(n56953), .B(n57318), .X(n23443) );
  nand_x4_sg U71970 ( .A(n23449), .B(n23450), .X(n23447) );
  nand_x1_sg U71971 ( .A(n51447), .B(n57320), .X(n23450) );
  nand_x1_sg U71972 ( .A(n56955), .B(n57318), .X(n23449) );
  nand_x4_sg U71973 ( .A(n23473), .B(n23474), .X(n23471) );
  nand_x1_sg U71974 ( .A(n47717), .B(n57320), .X(n23474) );
  nand_x1_sg U71975 ( .A(n56957), .B(n57318), .X(n23473) );
  nand_x4_sg U71976 ( .A(n23479), .B(n23480), .X(n23477) );
  nand_x1_sg U71977 ( .A(n51449), .B(n57320), .X(n23480) );
  nand_x1_sg U71978 ( .A(n56959), .B(n57318), .X(n23479) );
  nand_x4_sg U71979 ( .A(n23497), .B(n23498), .X(n23495) );
  nand_x1_sg U71980 ( .A(n47719), .B(n57320), .X(n23498) );
  nand_x1_sg U71981 ( .A(n56961), .B(n57318), .X(n23497) );
  nand_x4_sg U71982 ( .A(n23503), .B(n23504), .X(n23501) );
  nand_x1_sg U71983 ( .A(n51451), .B(n57320), .X(n23504) );
  nand_x1_sg U71984 ( .A(n56963), .B(n57318), .X(n23503) );
  nand_x4_sg U71985 ( .A(n23527), .B(n23528), .X(n23525) );
  nand_x1_sg U71986 ( .A(n47735), .B(n57320), .X(n23528) );
  nand_x1_sg U71987 ( .A(n56965), .B(n57318), .X(n23527) );
  nand_x4_sg U71988 ( .A(n23533), .B(n23534), .X(n23531) );
  nand_x1_sg U71989 ( .A(n51483), .B(n57320), .X(n23534) );
  nand_x1_sg U71990 ( .A(n56967), .B(n57318), .X(n23533) );
  nand_x4_sg U71991 ( .A(n23575), .B(n23576), .X(n23573) );
  nand_x1_sg U71992 ( .A(n47709), .B(n57320), .X(n23576) );
  nand_x1_sg U71993 ( .A(n56937), .B(n57318), .X(n23575) );
  nand_x4_sg U71994 ( .A(n23581), .B(n23582), .X(n23579) );
  nand_x1_sg U71995 ( .A(n51441), .B(n57320), .X(n23582) );
  nand_x1_sg U71996 ( .A(n56939), .B(n57318), .X(n23581) );
  nand_x4_sg U71997 ( .A(n23605), .B(n23606), .X(n23603) );
  nand_x1_sg U71998 ( .A(n47711), .B(n57320), .X(n23606) );
  nand_x1_sg U71999 ( .A(n56941), .B(n57318), .X(n23605) );
  nand_x4_sg U72000 ( .A(n23611), .B(n23612), .X(n23609) );
  nand_x1_sg U72001 ( .A(n51443), .B(n57320), .X(n23612) );
  nand_x1_sg U72002 ( .A(n56943), .B(n57318), .X(n23611) );
  nand_x4_sg U72003 ( .A(n23629), .B(n23630), .X(n23627) );
  nand_x1_sg U72004 ( .A(n47713), .B(n57320), .X(n23630) );
  nand_x1_sg U72005 ( .A(n56945), .B(n57318), .X(n23629) );
  nand_x4_sg U72006 ( .A(n23635), .B(n23636), .X(n23633) );
  nand_x1_sg U72007 ( .A(n51445), .B(n57320), .X(n23636) );
  nand_x1_sg U72008 ( .A(n56947), .B(n57318), .X(n23635) );
  nand_x4_sg U72009 ( .A(n23659), .B(n23660), .X(n23657) );
  nand_x1_sg U72010 ( .A(n47733), .B(n57320), .X(n23660) );
  nand_x1_sg U72011 ( .A(n56949), .B(n57318), .X(n23659) );
  nand_x4_sg U72012 ( .A(n23665), .B(n23666), .X(n23663) );
  nand_x1_sg U72013 ( .A(n51473), .B(n57320), .X(n23666) );
  nand_x1_sg U72014 ( .A(n56951), .B(n57318), .X(n23665) );
  nand_x4_sg U72015 ( .A(n23687), .B(n23688), .X(n23684) );
  nand_x1_sg U72016 ( .A(n47685), .B(n57316), .X(n23688) );
  nand_x4_sg U72017 ( .A(n23694), .B(n23695), .X(n23692) );
  nand_x1_sg U72018 ( .A(n47687), .B(n57316), .X(n23695) );
  nand_x4_sg U72019 ( .A(n23700), .B(n23701), .X(n23698) );
  nand_x1_sg U72020 ( .A(n51395), .B(n57316), .X(n23701) );
  nand_x4_sg U72021 ( .A(n23706), .B(n23707), .X(n23704) );
  nand_x1_sg U72022 ( .A(n51337), .B(n57316), .X(n23707) );
  nand_x4_sg U72023 ( .A(n23712), .B(n23713), .X(n23710) );
  nand_x1_sg U72024 ( .A(n56785), .B(n57316), .X(n23713) );
  nand_x4_sg U72025 ( .A(n23718), .B(n23719), .X(n23716) );
  nand_x1_sg U72026 ( .A(n47689), .B(n57316), .X(n23719) );
  nand_x4_sg U72027 ( .A(n23724), .B(n23725), .X(n23722) );
  nand_x1_sg U72028 ( .A(n51397), .B(n57316), .X(n23725) );
  nand_x4_sg U72029 ( .A(n23730), .B(n23731), .X(n23728) );
  nand_x1_sg U72030 ( .A(n56837), .B(n57316), .X(n23731) );
  nand_x4_sg U72031 ( .A(n23736), .B(n23737), .X(n23734) );
  nand_x1_sg U72032 ( .A(n51339), .B(n57316), .X(n23737) );
  nand_x4_sg U72033 ( .A(n23742), .B(n23743), .X(n23740) );
  nand_x1_sg U72034 ( .A(n56787), .B(n57316), .X(n23743) );
  nand_x4_sg U72035 ( .A(n23748), .B(n23749), .X(n23746) );
  nand_x1_sg U72036 ( .A(n51399), .B(n57316), .X(n23749) );
  nand_x4_sg U72037 ( .A(n23754), .B(n23755), .X(n23752) );
  nand_x1_sg U72038 ( .A(n56839), .B(n57316), .X(n23755) );
  nand_x4_sg U72039 ( .A(n23760), .B(n23761), .X(n23758) );
  nand_x1_sg U72040 ( .A(n51341), .B(n57316), .X(n23761) );
  nand_x4_sg U72041 ( .A(n23766), .B(n23767), .X(n23764) );
  nand_x1_sg U72042 ( .A(n56789), .B(n57316), .X(n23767) );
  nand_x4_sg U72043 ( .A(n23772), .B(n23773), .X(n23770) );
  nand_x1_sg U72044 ( .A(n51401), .B(n57316), .X(n23773) );
  nand_x4_sg U72045 ( .A(n23778), .B(n23779), .X(n23776) );
  nand_x1_sg U72046 ( .A(n56841), .B(n57316), .X(n23779) );
  nand_x4_sg U72047 ( .A(n23784), .B(n23785), .X(n23782) );
  nand_x1_sg U72048 ( .A(n56867), .B(n57316), .X(n23785) );
  nand_x4_sg U72049 ( .A(n23790), .B(n23791), .X(n23788) );
  nand_x1_sg U72050 ( .A(n47697), .B(n57316), .X(n23791) );
  nand_x4_sg U72051 ( .A(n23796), .B(n23797), .X(n23794) );
  nand_x1_sg U72052 ( .A(n51409), .B(n57316), .X(n23797) );
  nand_x4_sg U72053 ( .A(n23810), .B(n23811), .X(n23800) );
  nand_x1_sg U72054 ( .A(n56849), .B(n57316), .X(n23811) );
  nand_x4_sg U72055 ( .A(n23817), .B(n23818), .X(n23814) );
  nand_x1_sg U72056 ( .A(n47673), .B(n57316), .X(n23818) );
  nand_x4_sg U72057 ( .A(n23823), .B(n23824), .X(n23821) );
  nand_x1_sg U72058 ( .A(n47675), .B(n57316), .X(n23824) );
  nand_x4_sg U72059 ( .A(n23829), .B(n23830), .X(n23827) );
  nand_x1_sg U72060 ( .A(n51381), .B(n57316), .X(n23830) );
  nand_x4_sg U72061 ( .A(n23835), .B(n23836), .X(n23833) );
  nand_x1_sg U72062 ( .A(n51331), .B(n57316), .X(n23836) );
  nand_x4_sg U72063 ( .A(n23841), .B(n23842), .X(n23839) );
  nand_x1_sg U72064 ( .A(n56779), .B(n57316), .X(n23842) );
  nand_x4_sg U72065 ( .A(n23847), .B(n23848), .X(n23845) );
  nand_x1_sg U72066 ( .A(n47677), .B(n57316), .X(n23848) );
  nand_x4_sg U72067 ( .A(n23853), .B(n23854), .X(n23851) );
  nand_x1_sg U72068 ( .A(n51383), .B(n57316), .X(n23854) );
  nand_x4_sg U72069 ( .A(n23859), .B(n23860), .X(n23857) );
  nand_x1_sg U72070 ( .A(n56825), .B(n57316), .X(n23860) );
  nand_x4_sg U72071 ( .A(n23865), .B(n23866), .X(n23863) );
  nand_x1_sg U72072 ( .A(n51333), .B(n57316), .X(n23866) );
  nand_x4_sg U72073 ( .A(n23871), .B(n23872), .X(n23869) );
  nand_x1_sg U72074 ( .A(n56781), .B(n57316), .X(n23872) );
  nand_x4_sg U72075 ( .A(n23877), .B(n23878), .X(n23875) );
  nand_x1_sg U72076 ( .A(n51385), .B(n57316), .X(n23878) );
  nand_x4_sg U72077 ( .A(n23883), .B(n23884), .X(n23881) );
  nand_x1_sg U72078 ( .A(n56827), .B(n57316), .X(n23884) );
  nand_x4_sg U72079 ( .A(n23889), .B(n23890), .X(n23887) );
  nand_x1_sg U72080 ( .A(n51335), .B(n58376), .X(n23890) );
  nand_x4_sg U72081 ( .A(n23895), .B(n23896), .X(n23893) );
  nand_x1_sg U72082 ( .A(n56783), .B(n57316), .X(n23896) );
  nand_x4_sg U72083 ( .A(n23901), .B(n23902), .X(n23899) );
  nand_x1_sg U72084 ( .A(n51387), .B(n57316), .X(n23902) );
  nand_x4_sg U72085 ( .A(n23907), .B(n23908), .X(n23905) );
  nand_x1_sg U72086 ( .A(n56829), .B(n57316), .X(n23908) );
  nand_x4_sg U72087 ( .A(n23913), .B(n23914), .X(n23911) );
  nand_x1_sg U72088 ( .A(n56865), .B(n57316), .X(n23914) );
  nand_x4_sg U72089 ( .A(n23919), .B(n23920), .X(n23917) );
  nand_x1_sg U72090 ( .A(n47695), .B(n57316), .X(n23920) );
  nand_x4_sg U72091 ( .A(n23925), .B(n23926), .X(n23923) );
  nand_x1_sg U72092 ( .A(n51407), .B(n57316), .X(n23926) );
  nand_x4_sg U72093 ( .A(n23939), .B(n23940), .X(n23929) );
  nand_x1_sg U72094 ( .A(n56847), .B(n57316), .X(n23940) );
  nand_x4_sg U72095 ( .A(n67161), .B(n22752), .X(n22598) );
  nand_x1_sg U72096 ( .A(n47527), .B(n57864), .X(n22752) );
  nand_x4_sg U72097 ( .A(n67160), .B(n22766), .X(n22599) );
  nand_x1_sg U72098 ( .A(n47529), .B(n57864), .X(n22766) );
  nand_x4_sg U72099 ( .A(n67159), .B(n22777), .X(n22600) );
  nand_x1_sg U72100 ( .A(n56679), .B(n57864), .X(n22777) );
  nand_x4_sg U72101 ( .A(n67158), .B(n22788), .X(n22601) );
  nand_x1_sg U72102 ( .A(n56723), .B(n57864), .X(n22788) );
  nand_x4_sg U72103 ( .A(n67157), .B(n22799), .X(n22602) );
  nand_x1_sg U72104 ( .A(n51261), .B(n57864), .X(n22799) );
  nand_x4_sg U72105 ( .A(n67156), .B(n22810), .X(n22603) );
  nand_x1_sg U72106 ( .A(n47531), .B(n57864), .X(n22810) );
  nand_x4_sg U72107 ( .A(n67155), .B(n22821), .X(n22604) );
  nand_x1_sg U72108 ( .A(n56681), .B(n57864), .X(n22821) );
  nand_x4_sg U72109 ( .A(n67154), .B(n22832), .X(n22605) );
  nand_x1_sg U72110 ( .A(n51217), .B(n57864), .X(n22832) );
  nand_x4_sg U72111 ( .A(n67153), .B(n22843), .X(n22606) );
  nand_x1_sg U72112 ( .A(n56815), .B(n57864), .X(n22843) );
  nand_x4_sg U72113 ( .A(n67152), .B(n22854), .X(n22607) );
  nand_x1_sg U72114 ( .A(n51369), .B(n57864), .X(n22854) );
  nand_x4_sg U72115 ( .A(n67151), .B(n22865), .X(n22608) );
  nand_x1_sg U72116 ( .A(n56767), .B(n57864), .X(n22865) );
  nand_x4_sg U72117 ( .A(n67150), .B(n22876), .X(n22609) );
  nand_x1_sg U72118 ( .A(n51309), .B(n57864), .X(n22876) );
  nand_x4_sg U72119 ( .A(n67149), .B(n22887), .X(n22610) );
  nand_x1_sg U72120 ( .A(n56817), .B(n57864), .X(n22887) );
  nand_x4_sg U72121 ( .A(n67148), .B(n22898), .X(n22611) );
  nand_x1_sg U72122 ( .A(n51371), .B(n57864), .X(n22898) );
  nand_x4_sg U72123 ( .A(n67147), .B(n22909), .X(n22612) );
  nand_x1_sg U72124 ( .A(n51311), .B(n57864), .X(n22909) );
  nand_x4_sg U72125 ( .A(n67146), .B(n22920), .X(n22613) );
  nand_x1_sg U72126 ( .A(n56769), .B(n57864), .X(n22920) );
  nand_x4_sg U72127 ( .A(n67145), .B(n22931), .X(n22614) );
  nand_x1_sg U72128 ( .A(n51421), .B(n57864), .X(n22931) );
  nand_x4_sg U72129 ( .A(n67144), .B(n22942), .X(n22615) );
  nand_x1_sg U72130 ( .A(n56857), .B(n57864), .X(n22942) );
  nand_x4_sg U72131 ( .A(n67143), .B(n22953), .X(n22616) );
  nand_x1_sg U72132 ( .A(n47703), .B(n57864), .X(n22953) );
  nand_x4_sg U72133 ( .A(n67142), .B(n22964), .X(n22617) );
  nand_x1_sg U72134 ( .A(n51327), .B(n57864), .X(n22964) );
  nand_x4_sg U72135 ( .A(n67374), .B(n22980), .X(n22625) );
  nand_x1_sg U72136 ( .A(n47543), .B(n57864), .X(n22980) );
  nand_x4_sg U72137 ( .A(n67373), .B(n22993), .X(n22626) );
  nand_x1_sg U72138 ( .A(n47545), .B(n57864), .X(n22993) );
  nand_x4_sg U72139 ( .A(n67372), .B(n23004), .X(n22627) );
  nand_x1_sg U72140 ( .A(n56749), .B(n57864), .X(n23004) );
  nand_x4_sg U72141 ( .A(n67371), .B(n23015), .X(n22628) );
  nand_x1_sg U72142 ( .A(n56797), .B(n57864), .X(n23015) );
  nand_x4_sg U72143 ( .A(n67370), .B(n23026), .X(n22629) );
  nand_x1_sg U72144 ( .A(n51349), .B(n57864), .X(n23026) );
  nand_x4_sg U72145 ( .A(n67369), .B(n23037), .X(n22630) );
  nand_x1_sg U72146 ( .A(n47547), .B(n57864), .X(n23037) );
  nand_x4_sg U72147 ( .A(n67368), .B(n23048), .X(n22631) );
  nand_x1_sg U72148 ( .A(n56751), .B(n57864), .X(n23048) );
  nand_x4_sg U72149 ( .A(n67367), .B(n23059), .X(n22632) );
  nand_x1_sg U72150 ( .A(n51285), .B(n57864), .X(n23059) );
  nand_x4_sg U72151 ( .A(n67366), .B(n23070), .X(n22633) );
  nand_x1_sg U72152 ( .A(n56799), .B(n57864), .X(n23070) );
  nand_x4_sg U72153 ( .A(n67365), .B(n23081), .X(n22634) );
  nand_x1_sg U72154 ( .A(n51351), .B(n57864), .X(n23081) );
  nand_x4_sg U72155 ( .A(n67364), .B(n23092), .X(n22635) );
  nand_x1_sg U72156 ( .A(n56753), .B(n57864), .X(n23092) );
  nand_x4_sg U72157 ( .A(n67363), .B(n23103), .X(n22636) );
  nand_x1_sg U72158 ( .A(n51287), .B(n57864), .X(n23103) );
  nand_x4_sg U72159 ( .A(n67362), .B(n23114), .X(n22637) );
  nand_x1_sg U72160 ( .A(n56801), .B(n57864), .X(n23114) );
  nand_x4_sg U72161 ( .A(n67361), .B(n23125), .X(n22638) );
  nand_x1_sg U72162 ( .A(n51353), .B(n57864), .X(n23125) );
  nand_x4_sg U72163 ( .A(n67360), .B(n23136), .X(n22639) );
  nand_x1_sg U72164 ( .A(n51289), .B(n57864), .X(n23136) );
  nand_x4_sg U72165 ( .A(n67359), .B(n23147), .X(n22640) );
  nand_x1_sg U72166 ( .A(n56755), .B(n57864), .X(n23147) );
  nand_x4_sg U72167 ( .A(n67358), .B(n23158), .X(n22641) );
  nand_x1_sg U72168 ( .A(n51417), .B(n57864), .X(n23158) );
  nand_x4_sg U72169 ( .A(n67357), .B(n23169), .X(n22642) );
  nand_x1_sg U72170 ( .A(n56853), .B(n57864), .X(n23169) );
  nand_x4_sg U72171 ( .A(n67356), .B(n23180), .X(n22643) );
  nand_x1_sg U72172 ( .A(n47699), .B(n57864), .X(n23180) );
  nand_x4_sg U72173 ( .A(n67355), .B(n23191), .X(n22644) );
  nand_x1_sg U72174 ( .A(n51323), .B(n57864), .X(n23191) );
  nand_x4_sg U72175 ( .A(n67141), .B(n22753), .X(n22547) );
  nand_x1_sg U72176 ( .A(n47631), .B(n57345), .X(n22753) );
  nand_x4_sg U72177 ( .A(n67140), .B(n22767), .X(n22548) );
  nand_x1_sg U72178 ( .A(n47633), .B(n57345), .X(n22767) );
  nand_x4_sg U72179 ( .A(n67139), .B(n22778), .X(n22549) );
  nand_x1_sg U72180 ( .A(n51219), .B(n57345), .X(n22778) );
  nand_x4_sg U72181 ( .A(n67138), .B(n22789), .X(n22550) );
  nand_x1_sg U72182 ( .A(n51263), .B(n57345), .X(n22789) );
  nand_x4_sg U72183 ( .A(n67137), .B(n22800), .X(n22551) );
  nand_x1_sg U72184 ( .A(n56725), .B(n57345), .X(n22800) );
  nand_x4_sg U72185 ( .A(n67136), .B(n22811), .X(n22552) );
  nand_x1_sg U72186 ( .A(n47635), .B(n57345), .X(n22811) );
  nand_x4_sg U72187 ( .A(n67135), .B(n22822), .X(n22553) );
  nand_x1_sg U72188 ( .A(n51221), .B(n57345), .X(n22822) );
  nand_x4_sg U72189 ( .A(n67134), .B(n22833), .X(n22554) );
  nand_x1_sg U72190 ( .A(n56683), .B(n57345), .X(n22833) );
  nand_x4_sg U72191 ( .A(n67133), .B(n22844), .X(n22555) );
  nand_x1_sg U72192 ( .A(n51373), .B(n57345), .X(n22844) );
  nand_x4_sg U72193 ( .A(n67132), .B(n22855), .X(n22556) );
  nand_x1_sg U72194 ( .A(n56819), .B(n57345), .X(n22855) );
  nand_x4_sg U72195 ( .A(n67131), .B(n22866), .X(n22557) );
  nand_x1_sg U72196 ( .A(n51313), .B(n57345), .X(n22866) );
  nand_x4_sg U72197 ( .A(n67130), .B(n22877), .X(n22558) );
  nand_x1_sg U72198 ( .A(n56771), .B(n57345), .X(n22877) );
  nand_x4_sg U72199 ( .A(n67129), .B(n22888), .X(n22559) );
  nand_x1_sg U72200 ( .A(n51375), .B(n57345), .X(n22888) );
  nand_x4_sg U72201 ( .A(n67128), .B(n22899), .X(n22560) );
  nand_x1_sg U72202 ( .A(n56821), .B(n57345), .X(n22899) );
  nand_x4_sg U72203 ( .A(n67127), .B(n22910), .X(n22561) );
  nand_x1_sg U72204 ( .A(n51315), .B(n57345), .X(n22910) );
  nand_x4_sg U72205 ( .A(n67126), .B(n22921), .X(n22562) );
  nand_x1_sg U72206 ( .A(n56773), .B(n57345), .X(n22921) );
  nand_x4_sg U72207 ( .A(n67125), .B(n22932), .X(n22563) );
  nand_x1_sg U72208 ( .A(n56863), .B(n57345), .X(n22932) );
  nand_x4_sg U72209 ( .A(n67124), .B(n22943), .X(n22564) );
  nand_x1_sg U72210 ( .A(n47705), .B(n57345), .X(n22943) );
  nand_x4_sg U72211 ( .A(n67123), .B(n22954), .X(n22565) );
  nand_x1_sg U72212 ( .A(n51413), .B(n57345), .X(n22954) );
  nand_x4_sg U72213 ( .A(n67122), .B(n22965), .X(n22566) );
  nand_x1_sg U72214 ( .A(n56777), .B(n57345), .X(n22965) );
  nand_x4_sg U72215 ( .A(n67354), .B(n22981), .X(n22573) );
  nand_x1_sg U72216 ( .A(n47653), .B(n57345), .X(n22981) );
  nand_x4_sg U72217 ( .A(n67353), .B(n22994), .X(n22574) );
  nand_x1_sg U72218 ( .A(n47655), .B(n57345), .X(n22994) );
  nand_x4_sg U72219 ( .A(n67352), .B(n23005), .X(n22575) );
  nand_x1_sg U72220 ( .A(n51291), .B(n57345), .X(n23005) );
  nand_x4_sg U72221 ( .A(n67351), .B(n23016), .X(n22576) );
  nand_x1_sg U72222 ( .A(n51355), .B(n57345), .X(n23016) );
  nand_x4_sg U72223 ( .A(n67350), .B(n23027), .X(n22577) );
  nand_x1_sg U72224 ( .A(n56803), .B(n57345), .X(n23027) );
  nand_x4_sg U72225 ( .A(n67349), .B(n23038), .X(n22578) );
  nand_x1_sg U72226 ( .A(n47657), .B(n57345), .X(n23038) );
  nand_x4_sg U72227 ( .A(n67348), .B(n23049), .X(n22579) );
  nand_x1_sg U72228 ( .A(n51293), .B(n57345), .X(n23049) );
  nand_x4_sg U72229 ( .A(n67347), .B(n23060), .X(n22580) );
  nand_x1_sg U72230 ( .A(n56757), .B(n57345), .X(n23060) );
  nand_x4_sg U72231 ( .A(n67346), .B(n23071), .X(n22581) );
  nand_x1_sg U72232 ( .A(n51357), .B(n57345), .X(n23071) );
  nand_x4_sg U72233 ( .A(n67345), .B(n23082), .X(n22582) );
  nand_x1_sg U72234 ( .A(n56805), .B(n57345), .X(n23082) );
  nand_x4_sg U72235 ( .A(n67344), .B(n23093), .X(n22583) );
  nand_x1_sg U72236 ( .A(n51295), .B(n57345), .X(n23093) );
  nand_x4_sg U72237 ( .A(n67343), .B(n23104), .X(n22584) );
  nand_x1_sg U72238 ( .A(n56759), .B(n57345), .X(n23104) );
  nand_x4_sg U72239 ( .A(n67342), .B(n23115), .X(n22585) );
  nand_x1_sg U72240 ( .A(n51359), .B(n57345), .X(n23115) );
  nand_x4_sg U72241 ( .A(n67341), .B(n23126), .X(n22586) );
  nand_x1_sg U72242 ( .A(n56807), .B(n57345), .X(n23126) );
  nand_x4_sg U72243 ( .A(n67340), .B(n23137), .X(n22587) );
  nand_x1_sg U72244 ( .A(n51297), .B(n57345), .X(n23137) );
  nand_x4_sg U72245 ( .A(n67339), .B(n23148), .X(n22588) );
  nand_x1_sg U72246 ( .A(n56761), .B(n57345), .X(n23148) );
  nand_x4_sg U72247 ( .A(n67338), .B(n23159), .X(n22589) );
  nand_x1_sg U72248 ( .A(n56861), .B(n57345), .X(n23159) );
  nand_x4_sg U72249 ( .A(n67337), .B(n23170), .X(n22590) );
  nand_x1_sg U72250 ( .A(n47701), .B(n57345), .X(n23170) );
  nand_x4_sg U72251 ( .A(n67336), .B(n23181), .X(n22591) );
  nand_x1_sg U72252 ( .A(n51411), .B(n57345), .X(n23181) );
  nand_x4_sg U72253 ( .A(n67335), .B(n23192), .X(n22592) );
  nand_x1_sg U72254 ( .A(n56775), .B(n57345), .X(n23192) );
  nand_x4_sg U72255 ( .A(n67121), .B(n22754), .X(n22499) );
  nand_x1_sg U72256 ( .A(n47637), .B(n57858), .X(n22754) );
  nand_x4_sg U72257 ( .A(n67120), .B(n22768), .X(n22500) );
  nand_x1_sg U72258 ( .A(n47639), .B(n57858), .X(n22768) );
  nand_x4_sg U72259 ( .A(n67119), .B(n22779), .X(n22501) );
  nand_x1_sg U72260 ( .A(n51223), .B(n57858), .X(n22779) );
  nand_x4_sg U72261 ( .A(n67118), .B(n22790), .X(n22502) );
  nand_x1_sg U72262 ( .A(n51265), .B(n57858), .X(n22790) );
  nand_x4_sg U72263 ( .A(n67117), .B(n22801), .X(n22503) );
  nand_x1_sg U72264 ( .A(n56727), .B(n57858), .X(n22801) );
  nand_x4_sg U72265 ( .A(n67116), .B(n22812), .X(n22504) );
  nand_x1_sg U72266 ( .A(n47641), .B(n57858), .X(n22812) );
  nand_x4_sg U72267 ( .A(n67115), .B(n22823), .X(n22505) );
  nand_x1_sg U72268 ( .A(n51225), .B(n57860), .X(n22823) );
  nand_x4_sg U72269 ( .A(n67114), .B(n22834), .X(n22506) );
  nand_x1_sg U72270 ( .A(n56685), .B(n57860), .X(n22834) );
  nand_x4_sg U72271 ( .A(n67113), .B(n22845), .X(n22507) );
  nand_x1_sg U72272 ( .A(n51267), .B(n57860), .X(n22845) );
  nand_x4_sg U72273 ( .A(n67112), .B(n22856), .X(n22508) );
  nand_x1_sg U72274 ( .A(n56729), .B(n57860), .X(n22856) );
  nand_x4_sg U72275 ( .A(n67111), .B(n22867), .X(n22509) );
  nand_x1_sg U72276 ( .A(n51227), .B(n57860), .X(n22867) );
  nand_x4_sg U72277 ( .A(n67110), .B(n22878), .X(n22510) );
  nand_x1_sg U72278 ( .A(n56687), .B(n57860), .X(n22878) );
  nand_x4_sg U72279 ( .A(n67109), .B(n22889), .X(n22511) );
  nand_x1_sg U72280 ( .A(n51269), .B(n57860), .X(n22889) );
  nand_x4_sg U72281 ( .A(n67108), .B(n22900), .X(n22512) );
  nand_x1_sg U72282 ( .A(n56731), .B(n57860), .X(n22900) );
  nand_x4_sg U72283 ( .A(n67107), .B(n22911), .X(n22513) );
  nand_x1_sg U72284 ( .A(n51241), .B(n57860), .X(n22911) );
  nand_x4_sg U72285 ( .A(n67106), .B(n22922), .X(n22514) );
  nand_x1_sg U72286 ( .A(n56703), .B(n57860), .X(n22922) );
  nand_x4_sg U72287 ( .A(n67105), .B(n22933), .X(n22515) );
  nand_x1_sg U72288 ( .A(n47691), .B(n57858), .X(n22933) );
  nand_x4_sg U72289 ( .A(n67104), .B(n22944), .X(n22516) );
  nand_x1_sg U72290 ( .A(n51403), .B(n57860), .X(n22944) );
  nand_x4_sg U72291 ( .A(n67103), .B(n22955), .X(n22517) );
  nand_x1_sg U72292 ( .A(n56843), .B(n57860), .X(n22955) );
  nand_x4_sg U72293 ( .A(n67102), .B(n22966), .X(n22518) );
  nand_x1_sg U72294 ( .A(n56689), .B(n57860), .X(n22966) );
  nand_x4_sg U72295 ( .A(n67334), .B(n22982), .X(n22524) );
  nand_x1_sg U72296 ( .A(n47617), .B(n57860), .X(n22982) );
  nand_x4_sg U72297 ( .A(n67333), .B(n22995), .X(n22525) );
  nand_x1_sg U72298 ( .A(n47619), .B(n57860), .X(n22995) );
  nand_x4_sg U72299 ( .A(n67332), .B(n23006), .X(n22526) );
  nand_x1_sg U72300 ( .A(n51201), .B(n57860), .X(n23006) );
  nand_x4_sg U72301 ( .A(n67331), .B(n23017), .X(n22527) );
  nand_x1_sg U72302 ( .A(n51245), .B(n57860), .X(n23017) );
  nand_x4_sg U72303 ( .A(n67330), .B(n23028), .X(n22528) );
  nand_x1_sg U72304 ( .A(n56707), .B(n57860), .X(n23028) );
  nand_x4_sg U72305 ( .A(n67329), .B(n23039), .X(n22529) );
  nand_x1_sg U72306 ( .A(n47621), .B(n57860), .X(n23039) );
  nand_x4_sg U72307 ( .A(n67328), .B(n23050), .X(n22530) );
  nand_x1_sg U72308 ( .A(n51203), .B(n57860), .X(n23050) );
  nand_x4_sg U72309 ( .A(n67327), .B(n23061), .X(n22531) );
  nand_x1_sg U72310 ( .A(n56661), .B(n57860), .X(n23061) );
  nand_x4_sg U72311 ( .A(n67326), .B(n23072), .X(n22532) );
  nand_x1_sg U72312 ( .A(n51247), .B(n57860), .X(n23072) );
  nand_x4_sg U72313 ( .A(n67325), .B(n23083), .X(n22533) );
  nand_x1_sg U72314 ( .A(n56709), .B(n57860), .X(n23083) );
  nand_x4_sg U72315 ( .A(n67324), .B(n23094), .X(n22534) );
  nand_x1_sg U72316 ( .A(n51205), .B(n29333), .X(n23094) );
  nand_x4_sg U72317 ( .A(n67323), .B(n23105), .X(n22535) );
  nand_x1_sg U72318 ( .A(n56663), .B(n57860), .X(n23105) );
  nand_x4_sg U72319 ( .A(n67322), .B(n23116), .X(n22536) );
  nand_x1_sg U72320 ( .A(n51249), .B(n57860), .X(n23116) );
  nand_x4_sg U72321 ( .A(n67321), .B(n23127), .X(n22537) );
  nand_x1_sg U72322 ( .A(n56711), .B(n57860), .X(n23127) );
  nand_x4_sg U72323 ( .A(n67320), .B(n23138), .X(n22538) );
  nand_x1_sg U72324 ( .A(n51237), .B(n57860), .X(n23138) );
  nand_x4_sg U72325 ( .A(n67319), .B(n23149), .X(n22539) );
  nand_x1_sg U72326 ( .A(n56699), .B(n57860), .X(n23149) );
  nand_x4_sg U72327 ( .A(n67318), .B(n23160), .X(n22540) );
  nand_x1_sg U72328 ( .A(n47679), .B(n57860), .X(n23160) );
  nand_x4_sg U72329 ( .A(n67317), .B(n23171), .X(n22541) );
  nand_x1_sg U72330 ( .A(n51389), .B(n57860), .X(n23171) );
  nand_x4_sg U72331 ( .A(n67316), .B(n23182), .X(n22542) );
  nand_x1_sg U72332 ( .A(n56831), .B(n29333), .X(n23182) );
  nand_x4_sg U72333 ( .A(n67315), .B(n23193), .X(n22543) );
  nand_x1_sg U72334 ( .A(n56665), .B(n57860), .X(n23193) );
  nand_x4_sg U72335 ( .A(n67281), .B(n24606), .X(n24603) );
  nor_x1_sg U72336 ( .A(n58125), .B(n47364), .X(n58126) );
  nand_x4_sg U72337 ( .A(n67280), .B(n24611), .X(n24609) );
  nor_x1_sg U72338 ( .A(n58125), .B(n47366), .X(n58120) );
  nand_x4_sg U72339 ( .A(n67279), .B(n24615), .X(n24613) );
  nor_x1_sg U72340 ( .A(n58125), .B(n56922), .X(n58117) );
  nand_x4_sg U72341 ( .A(n67278), .B(n24619), .X(n24617) );
  nor_x1_sg U72342 ( .A(n58125), .B(n58113), .X(n58114) );
  nand_x4_sg U72343 ( .A(n67277), .B(n24623), .X(n24621) );
  nor_x1_sg U72344 ( .A(n58125), .B(n58109), .X(n58110) );
  nand_x4_sg U72345 ( .A(n67276), .B(n24627), .X(n24625) );
  nor_x1_sg U72346 ( .A(n58125), .B(n47368), .X(n58106) );
  nand_x4_sg U72347 ( .A(n67275), .B(n24631), .X(n24629) );
  nor_x1_sg U72348 ( .A(n58125), .B(n47428), .X(n58103) );
  nand_x4_sg U72349 ( .A(n67274), .B(n24635), .X(n24633) );
  nor_x1_sg U72350 ( .A(n58125), .B(n56924), .X(n58100) );
  nand_x4_sg U72351 ( .A(n67273), .B(n24639), .X(n24637) );
  nor_x1_sg U72352 ( .A(n58125), .B(n58096), .X(n58097) );
  nand_x4_sg U72353 ( .A(n67272), .B(n24643), .X(n24641) );
  nor_x1_sg U72354 ( .A(n58125), .B(n58092), .X(n58093) );
  nand_x4_sg U72355 ( .A(n67271), .B(n24647), .X(n24645) );
  nor_x1_sg U72356 ( .A(n58125), .B(n47430), .X(n58089) );
  nand_x4_sg U72357 ( .A(n67270), .B(n24651), .X(n24649) );
  nor_x1_sg U72358 ( .A(n58125), .B(n56926), .X(n58086) );
  nand_x4_sg U72359 ( .A(n67269), .B(n24655), .X(n24653) );
  nor_x1_sg U72360 ( .A(n58125), .B(n58082), .X(n58083) );
  nand_x4_sg U72361 ( .A(n67268), .B(n24659), .X(n24657) );
  nor_x1_sg U72362 ( .A(n58125), .B(n58078), .X(n58079) );
  nand_x4_sg U72363 ( .A(n67267), .B(n24663), .X(n24661) );
  nor_x1_sg U72364 ( .A(n58125), .B(n47370), .X(n58075) );
  nand_x4_sg U72365 ( .A(n67266), .B(n24667), .X(n24665) );
  nor_x1_sg U72366 ( .A(n58125), .B(n47432), .X(n58072) );
  nand_x4_sg U72367 ( .A(n67265), .B(n24671), .X(n24669) );
  nor_x1_sg U72368 ( .A(n58125), .B(n56932), .X(n58069) );
  nand_x4_sg U72369 ( .A(n67264), .B(n24675), .X(n24673) );
  nor_x1_sg U72370 ( .A(n58125), .B(n58065), .X(n58066) );
  nand_x4_sg U72371 ( .A(n67263), .B(n24679), .X(n24677) );
  nor_x1_sg U72372 ( .A(n58125), .B(n58061), .X(n58062) );
  nand_x4_sg U72373 ( .A(n67262), .B(n24696), .X(n24681) );
  nor_x1_sg U72374 ( .A(n58125), .B(n47434), .X(n58058) );
  nand_x4_sg U72375 ( .A(n67474), .B(n24701), .X(n24698) );
  nor_x1_sg U72376 ( .A(n58125), .B(n47356), .X(n58055) );
  nand_x4_sg U72377 ( .A(n67473), .B(n24705), .X(n24703) );
  nor_x1_sg U72378 ( .A(n58125), .B(n47358), .X(n58050) );
  nand_x4_sg U72379 ( .A(n67472), .B(n24709), .X(n24707) );
  nor_x1_sg U72380 ( .A(n58125), .B(n56916), .X(n58047) );
  nand_x4_sg U72381 ( .A(n67471), .B(n24713), .X(n24711) );
  nor_x1_sg U72382 ( .A(n58125), .B(n58043), .X(n58044) );
  nand_x4_sg U72383 ( .A(n67470), .B(n24717), .X(n24715) );
  nor_x1_sg U72384 ( .A(n58125), .B(n58039), .X(n58040) );
  nand_x4_sg U72385 ( .A(n67469), .B(n24721), .X(n24719) );
  nor_x1_sg U72386 ( .A(n58125), .B(n47360), .X(n58036) );
  nand_x4_sg U72387 ( .A(n67468), .B(n24725), .X(n24723) );
  nor_x1_sg U72388 ( .A(n58125), .B(n47420), .X(n58033) );
  nand_x4_sg U72389 ( .A(n67467), .B(n24729), .X(n24727) );
  nor_x1_sg U72390 ( .A(n58125), .B(n56918), .X(n58030) );
  nand_x4_sg U72391 ( .A(n67466), .B(n24733), .X(n24731) );
  nor_x1_sg U72392 ( .A(n58125), .B(n58026), .X(n58027) );
  nand_x4_sg U72393 ( .A(n67465), .B(n24737), .X(n24735) );
  nor_x1_sg U72394 ( .A(n58125), .B(n58022), .X(n58023) );
  nand_x4_sg U72395 ( .A(n67464), .B(n24741), .X(n24739) );
  nor_x1_sg U72396 ( .A(n58125), .B(n47422), .X(n58019) );
  nand_x4_sg U72397 ( .A(n67463), .B(n24745), .X(n24743) );
  nor_x1_sg U72398 ( .A(n58125), .B(n56920), .X(n58016) );
  nand_x4_sg U72399 ( .A(n67462), .B(n24749), .X(n24747) );
  nor_x1_sg U72400 ( .A(n58125), .B(n58012), .X(n58013) );
  nand_x4_sg U72401 ( .A(n67461), .B(n24753), .X(n24751) );
  nor_x1_sg U72402 ( .A(n58125), .B(n58008), .X(n58009) );
  nand_x4_sg U72403 ( .A(n67460), .B(n24757), .X(n24755) );
  nor_x1_sg U72404 ( .A(n58125), .B(n47362), .X(n58005) );
  nand_x4_sg U72405 ( .A(n67459), .B(n24761), .X(n24759) );
  nor_x1_sg U72406 ( .A(n58125), .B(n47424), .X(n58002) );
  nand_x4_sg U72407 ( .A(n67458), .B(n24765), .X(n24763) );
  nor_x1_sg U72408 ( .A(n58125), .B(n56930), .X(n57999) );
  nand_x4_sg U72409 ( .A(n67457), .B(n24769), .X(n24767) );
  nor_x1_sg U72410 ( .A(n58125), .B(n57995), .X(n57996) );
  nand_x4_sg U72411 ( .A(n67456), .B(n24773), .X(n24771) );
  nor_x1_sg U72412 ( .A(n58125), .B(n57991), .X(n57992) );
  nand_x4_sg U72413 ( .A(n67455), .B(n24789), .X(n24775) );
  nor_x1_sg U72414 ( .A(n58125), .B(n47426), .X(n57988) );
  nand_x4_sg U72415 ( .A(n61862), .B(n22755), .X(n22447) );
  nand_x1_sg U72416 ( .A(n47643), .B(n57463), .X(n22755) );
  nand_x4_sg U72417 ( .A(n61863), .B(n22769), .X(n22448) );
  nand_x1_sg U72418 ( .A(n47645), .B(n57463), .X(n22769) );
  nand_x4_sg U72419 ( .A(n61864), .B(n22780), .X(n22449) );
  nand_x1_sg U72420 ( .A(n51229), .B(n57463), .X(n22780) );
  nand_x4_sg U72421 ( .A(n61865), .B(n22791), .X(n22450) );
  nand_x1_sg U72422 ( .A(n51271), .B(n57463), .X(n22791) );
  nand_x4_sg U72423 ( .A(n61866), .B(n22802), .X(n22451) );
  nand_x1_sg U72424 ( .A(n56733), .B(n57463), .X(n22802) );
  nand_x4_sg U72425 ( .A(n61867), .B(n22813), .X(n22452) );
  nand_x1_sg U72426 ( .A(n47647), .B(n57463), .X(n22813) );
  nand_x4_sg U72427 ( .A(n61868), .B(n22824), .X(n22453) );
  nand_x1_sg U72428 ( .A(n51231), .B(n57463), .X(n22824) );
  nand_x4_sg U72429 ( .A(n61869), .B(n22835), .X(n22454) );
  nand_x1_sg U72430 ( .A(n56691), .B(n57463), .X(n22835) );
  nand_x4_sg U72431 ( .A(n61870), .B(n22846), .X(n22455) );
  nand_x1_sg U72432 ( .A(n51273), .B(n57463), .X(n22846) );
  nand_x4_sg U72433 ( .A(n61871), .B(n22857), .X(n22456) );
  nand_x1_sg U72434 ( .A(n56735), .B(n57463), .X(n22857) );
  nand_x4_sg U72435 ( .A(n61872), .B(n22868), .X(n22457) );
  nand_x1_sg U72436 ( .A(n51233), .B(n57463), .X(n22868) );
  nand_x4_sg U72437 ( .A(n61873), .B(n22879), .X(n22458) );
  nand_x1_sg U72438 ( .A(n56693), .B(n57463), .X(n22879) );
  nand_x4_sg U72439 ( .A(n61874), .B(n22890), .X(n22459) );
  nand_x1_sg U72440 ( .A(n51275), .B(n57463), .X(n22890) );
  nand_x4_sg U72441 ( .A(n61875), .B(n22901), .X(n22460) );
  nand_x1_sg U72442 ( .A(n56737), .B(n57463), .X(n22901) );
  nand_x4_sg U72443 ( .A(n61876), .B(n22912), .X(n22461) );
  nand_x1_sg U72444 ( .A(n51243), .B(n57463), .X(n22912) );
  nand_x4_sg U72445 ( .A(n61877), .B(n22923), .X(n22462) );
  nand_x1_sg U72446 ( .A(n56705), .B(n57463), .X(n22923) );
  nand_x4_sg U72447 ( .A(n61878), .B(n22934), .X(n22463) );
  nand_x1_sg U72448 ( .A(n47693), .B(n57463), .X(n22934) );
  nand_x4_sg U72449 ( .A(n61879), .B(n22945), .X(n22464) );
  nand_x1_sg U72450 ( .A(n51405), .B(n57463), .X(n22945) );
  nand_x4_sg U72451 ( .A(n61880), .B(n22956), .X(n22465) );
  nand_x1_sg U72452 ( .A(n56845), .B(n57463), .X(n22956) );
  nand_x4_sg U72453 ( .A(n61881), .B(n22967), .X(n22466) );
  nand_x1_sg U72454 ( .A(n56695), .B(n57463), .X(n22967) );
  nand_x4_sg U72455 ( .A(n61882), .B(n22983), .X(n22474) );
  nand_x1_sg U72456 ( .A(n47623), .B(n57463), .X(n22983) );
  nand_x4_sg U72457 ( .A(n61883), .B(n22996), .X(n22475) );
  nand_x1_sg U72458 ( .A(n47625), .B(n57463), .X(n22996) );
  nand_x4_sg U72459 ( .A(n61884), .B(n23007), .X(n22476) );
  nand_x1_sg U72460 ( .A(n51207), .B(n57463), .X(n23007) );
  nand_x4_sg U72461 ( .A(n61885), .B(n23018), .X(n22477) );
  nand_x1_sg U72462 ( .A(n51251), .B(n57463), .X(n23018) );
  nand_x4_sg U72463 ( .A(n61886), .B(n23029), .X(n22478) );
  nand_x1_sg U72464 ( .A(n56713), .B(n57463), .X(n23029) );
  nand_x4_sg U72465 ( .A(n61887), .B(n23040), .X(n22479) );
  nand_x1_sg U72466 ( .A(n47627), .B(n57463), .X(n23040) );
  nand_x4_sg U72467 ( .A(n61888), .B(n23051), .X(n22480) );
  nand_x1_sg U72468 ( .A(n51209), .B(n57463), .X(n23051) );
  nand_x4_sg U72469 ( .A(n61889), .B(n23062), .X(n22481) );
  nand_x1_sg U72470 ( .A(n56667), .B(n57463), .X(n23062) );
  nand_x4_sg U72471 ( .A(n61890), .B(n23073), .X(n22482) );
  nand_x1_sg U72472 ( .A(n51253), .B(n57463), .X(n23073) );
  nand_x4_sg U72473 ( .A(n61891), .B(n23084), .X(n22483) );
  nand_x1_sg U72474 ( .A(n56715), .B(n57463), .X(n23084) );
  nand_x4_sg U72475 ( .A(n61892), .B(n23095), .X(n22484) );
  nand_x1_sg U72476 ( .A(n51211), .B(n57463), .X(n23095) );
  nand_x4_sg U72477 ( .A(n61893), .B(n23106), .X(n22485) );
  nand_x1_sg U72478 ( .A(n56669), .B(n57463), .X(n23106) );
  nand_x4_sg U72479 ( .A(n61894), .B(n23117), .X(n22486) );
  nand_x1_sg U72480 ( .A(n51255), .B(n57463), .X(n23117) );
  nand_x4_sg U72481 ( .A(n61895), .B(n23128), .X(n22487) );
  nand_x1_sg U72482 ( .A(n56717), .B(n57463), .X(n23128) );
  nand_x4_sg U72483 ( .A(n61896), .B(n23139), .X(n22488) );
  nand_x1_sg U72484 ( .A(n51239), .B(n57463), .X(n23139) );
  nand_x4_sg U72485 ( .A(n61897), .B(n23150), .X(n22489) );
  nand_x1_sg U72486 ( .A(n56701), .B(n57463), .X(n23150) );
  nand_x4_sg U72487 ( .A(n61898), .B(n23161), .X(n22490) );
  nand_x1_sg U72488 ( .A(n47681), .B(n57463), .X(n23161) );
  nand_x4_sg U72489 ( .A(n61899), .B(n23172), .X(n22491) );
  nand_x1_sg U72490 ( .A(n51391), .B(n57463), .X(n23172) );
  nand_x4_sg U72491 ( .A(n61900), .B(n23183), .X(n22492) );
  nand_x1_sg U72492 ( .A(n56833), .B(n57463), .X(n23183) );
  nand_x4_sg U72493 ( .A(n61901), .B(n23194), .X(n22493) );
  nand_x1_sg U72494 ( .A(n56671), .B(n57463), .X(n23194) );
  nand_x1_sg U72495 ( .A(n47715), .B(n57949), .X(n58313) );
  nand_x1_sg U72496 ( .A(n56953), .B(n57930), .X(n58314) );
  nand_x1_sg U72497 ( .A(n51447), .B(n57949), .X(n58308) );
  nand_x1_sg U72498 ( .A(n56955), .B(n57930), .X(n58309) );
  nand_x1_sg U72499 ( .A(n47717), .B(n57949), .X(n58288) );
  nand_x1_sg U72500 ( .A(n56957), .B(n57931), .X(n58289) );
  nand_x1_sg U72501 ( .A(n51449), .B(n57949), .X(n58283) );
  nand_x1_sg U72502 ( .A(n56959), .B(n57931), .X(n58284) );
  nand_x1_sg U72503 ( .A(n47719), .B(n57949), .X(n58268) );
  nand_x1_sg U72504 ( .A(n56961), .B(n57932), .X(n58269) );
  nand_x1_sg U72505 ( .A(n51451), .B(n57949), .X(n58263) );
  nand_x1_sg U72506 ( .A(n56963), .B(n57932), .X(n58264) );
  nand_x1_sg U72507 ( .A(n47735), .B(n57949), .X(n58243) );
  nand_x1_sg U72508 ( .A(n56965), .B(n57933), .X(n58244) );
  nand_x1_sg U72509 ( .A(n51483), .B(n57949), .X(n58238) );
  nand_x1_sg U72510 ( .A(n56967), .B(n57934), .X(n58239) );
  nand_x1_sg U72511 ( .A(n47709), .B(n57949), .X(n58213) );
  nand_x1_sg U72512 ( .A(n56937), .B(n57935), .X(n58214) );
  nand_x1_sg U72513 ( .A(n51441), .B(n57949), .X(n58208) );
  nand_x1_sg U72514 ( .A(n56939), .B(n57936), .X(n58209) );
  nand_x1_sg U72515 ( .A(n47711), .B(n57949), .X(n58188) );
  nand_x1_sg U72516 ( .A(n56941), .B(n57937), .X(n58189) );
  nand_x1_sg U72517 ( .A(n51443), .B(n57949), .X(n58183) );
  nand_x1_sg U72518 ( .A(n56943), .B(n57937), .X(n58184) );
  nand_x1_sg U72519 ( .A(n47713), .B(n57949), .X(n58168) );
  nand_x1_sg U72520 ( .A(n56945), .B(n57938), .X(n58169) );
  nand_x1_sg U72521 ( .A(n51445), .B(n57949), .X(n58163) );
  nand_x1_sg U72522 ( .A(n56947), .B(n57939), .X(n58164) );
  nand_x1_sg U72523 ( .A(n47733), .B(n57949), .X(n58143) );
  nand_x1_sg U72524 ( .A(n56949), .B(n57940), .X(n58144) );
  nand_x1_sg U72525 ( .A(n51473), .B(n57949), .X(n58138) );
  nand_x1_sg U72526 ( .A(n56951), .B(n57941), .X(n58139) );
  nor_x1_sg U72527 ( .A(n23308), .B(n23309), .X(n23307) );
  nand_x2_sg U72528 ( .A(n24801), .B(n24802), .X(n24796) );
  nand_x1_sg U72529 ( .A(n57501), .B(n47527), .X(n24802) );
  nand_x1_sg U72530 ( .A(n57504), .B(n47743), .X(n24801) );
  nand_x2_sg U72531 ( .A(n24839), .B(n24840), .X(n24835) );
  nand_x1_sg U72532 ( .A(n57499), .B(n47529), .X(n24840) );
  nand_x1_sg U72533 ( .A(n57502), .B(n47745), .X(n24839) );
  nand_x2_sg U72534 ( .A(n24869), .B(n24870), .X(n24865) );
  nand_x1_sg U72535 ( .A(n57499), .B(n56679), .X(n24870) );
  nand_x1_sg U72536 ( .A(n57502), .B(n51489), .X(n24869) );
  nand_x2_sg U72537 ( .A(n24899), .B(n24900), .X(n24895) );
  nand_x1_sg U72538 ( .A(n57499), .B(n56723), .X(n24900) );
  nand_x1_sg U72539 ( .A(n57502), .B(n51493), .X(n24899) );
  nand_x2_sg U72540 ( .A(n24929), .B(n24930), .X(n24925) );
  nand_x1_sg U72541 ( .A(n57499), .B(n51261), .X(n24930) );
  nand_x1_sg U72542 ( .A(n57502), .B(n57015), .X(n24929) );
  nand_x2_sg U72543 ( .A(n24959), .B(n24960), .X(n24955) );
  nand_x1_sg U72544 ( .A(n57499), .B(n47531), .X(n24960) );
  nand_x1_sg U72545 ( .A(n57502), .B(n47747), .X(n24959) );
  nand_x2_sg U72546 ( .A(n24989), .B(n24990), .X(n24985) );
  nand_x1_sg U72547 ( .A(n57499), .B(n56681), .X(n24990) );
  nand_x1_sg U72548 ( .A(n57502), .B(n51491), .X(n24989) );
  nand_x2_sg U72549 ( .A(n25019), .B(n25020), .X(n25015) );
  nand_x1_sg U72550 ( .A(n57499), .B(n51217), .X(n25020) );
  nand_x1_sg U72551 ( .A(n57502), .B(n57013), .X(n25019) );
  nand_x2_sg U72552 ( .A(n25049), .B(n25050), .X(n25045) );
  nand_x1_sg U72553 ( .A(n57499), .B(n56815), .X(n25050) );
  nand_x1_sg U72554 ( .A(n57502), .B(n51515), .X(n25049) );
  nand_x2_sg U72555 ( .A(n25079), .B(n25080), .X(n25075) );
  nand_x1_sg U72556 ( .A(n57499), .B(n51369), .X(n25080) );
  nand_x1_sg U72557 ( .A(n57502), .B(n57039), .X(n25079) );
  nand_x2_sg U72558 ( .A(n25109), .B(n25110), .X(n25105) );
  nand_x1_sg U72559 ( .A(n57499), .B(n56767), .X(n25110) );
  nand_x1_sg U72560 ( .A(n57502), .B(n51503), .X(n25109) );
  nand_x2_sg U72561 ( .A(n25139), .B(n25140), .X(n25135) );
  nand_x1_sg U72562 ( .A(n57499), .B(n51309), .X(n25140) );
  nand_x1_sg U72563 ( .A(n57502), .B(n57021), .X(n25139) );
  nand_x2_sg U72564 ( .A(n25169), .B(n25170), .X(n25165) );
  nand_x1_sg U72565 ( .A(n57499), .B(n56817), .X(n25170) );
  nand_x1_sg U72566 ( .A(n57502), .B(n51517), .X(n25169) );
  nand_x2_sg U72567 ( .A(n25199), .B(n25200), .X(n25195) );
  nand_x1_sg U72568 ( .A(n57499), .B(n51371), .X(n25200) );
  nand_x1_sg U72569 ( .A(n57502), .B(n57041), .X(n25199) );
  nand_x2_sg U72570 ( .A(n25229), .B(n25230), .X(n25225) );
  nand_x1_sg U72571 ( .A(n57499), .B(n51311), .X(n25230) );
  nand_x1_sg U72572 ( .A(n57502), .B(n47757), .X(n25229) );
  nand_x2_sg U72573 ( .A(n25259), .B(n25260), .X(n25255) );
  nand_x1_sg U72574 ( .A(n57499), .B(n56769), .X(n25260) );
  nand_x1_sg U72575 ( .A(n57502), .B(n51505), .X(n25259) );
  nand_x2_sg U72576 ( .A(n25289), .B(n25290), .X(n25285) );
  nand_x1_sg U72577 ( .A(n57499), .B(n51421), .X(n25290) );
  nand_x1_sg U72578 ( .A(n57502), .B(n57027), .X(n25289) );
  nand_x2_sg U72579 ( .A(n25319), .B(n25320), .X(n25315) );
  nand_x1_sg U72580 ( .A(n57499), .B(n56857), .X(n25320) );
  nand_x1_sg U72581 ( .A(n57502), .B(n51519), .X(n25319) );
  nand_x2_sg U72582 ( .A(n25349), .B(n25350), .X(n25345) );
  nand_x1_sg U72583 ( .A(n57499), .B(n47703), .X(n25350) );
  nand_x1_sg U72584 ( .A(n57502), .B(n57043), .X(n25349) );
  nand_x2_sg U72585 ( .A(n25380), .B(n25381), .X(n25376) );
  nand_x1_sg U72586 ( .A(n57499), .B(n51327), .X(n25381) );
  nand_x1_sg U72587 ( .A(n57502), .B(n57029), .X(n25380) );
  nand_x2_sg U72588 ( .A(n25411), .B(n25412), .X(n25407) );
  nand_x1_sg U72589 ( .A(n57499), .B(n47543), .X(n25412) );
  nand_x1_sg U72590 ( .A(n57502), .B(n47749), .X(n25411) );
  nand_x2_sg U72591 ( .A(n25441), .B(n25442), .X(n25437) );
  nand_x1_sg U72592 ( .A(n57499), .B(n47545), .X(n25442) );
  nand_x1_sg U72593 ( .A(n57502), .B(n47751), .X(n25441) );
  nand_x2_sg U72594 ( .A(n25471), .B(n25472), .X(n25467) );
  nand_x1_sg U72595 ( .A(n57499), .B(n56749), .X(n25472) );
  nand_x1_sg U72596 ( .A(n57502), .B(n51495), .X(n25471) );
  nand_x2_sg U72597 ( .A(n25501), .B(n25502), .X(n25497) );
  nand_x1_sg U72598 ( .A(n57499), .B(n56797), .X(n25502) );
  nand_x1_sg U72599 ( .A(n57502), .B(n51507), .X(n25501) );
  nand_x2_sg U72600 ( .A(n25531), .B(n25532), .X(n25527) );
  nand_x1_sg U72601 ( .A(n57499), .B(n51349), .X(n25532) );
  nand_x1_sg U72602 ( .A(n57502), .B(n57031), .X(n25531) );
  nand_x2_sg U72603 ( .A(n25561), .B(n25562), .X(n25557) );
  nand_x1_sg U72604 ( .A(n57499), .B(n47547), .X(n25562) );
  nand_x1_sg U72605 ( .A(n57502), .B(n47753), .X(n25561) );
  nand_x2_sg U72606 ( .A(n25591), .B(n25592), .X(n25587) );
  nand_x1_sg U72607 ( .A(n57499), .B(n56751), .X(n25592) );
  nand_x1_sg U72608 ( .A(n57502), .B(n51497), .X(n25591) );
  nand_x2_sg U72609 ( .A(n25621), .B(n25622), .X(n25617) );
  nand_x1_sg U72610 ( .A(n57499), .B(n51285), .X(n25622) );
  nand_x1_sg U72611 ( .A(n57502), .B(n57017), .X(n25621) );
  nand_x2_sg U72612 ( .A(n25651), .B(n25652), .X(n25647) );
  nand_x1_sg U72613 ( .A(n57499), .B(n56799), .X(n25652) );
  nand_x1_sg U72614 ( .A(n57502), .B(n51509), .X(n25651) );
  nand_x2_sg U72615 ( .A(n25681), .B(n25682), .X(n25677) );
  nand_x1_sg U72616 ( .A(n57499), .B(n51351), .X(n25682) );
  nand_x1_sg U72617 ( .A(n57502), .B(n57033), .X(n25681) );
  nand_x2_sg U72618 ( .A(n25711), .B(n25712), .X(n25707) );
  nand_x1_sg U72619 ( .A(n57499), .B(n56753), .X(n25712) );
  nand_x1_sg U72620 ( .A(n57502), .B(n51499), .X(n25711) );
  nand_x2_sg U72621 ( .A(n25741), .B(n25742), .X(n25737) );
  nand_x1_sg U72622 ( .A(n57499), .B(n51287), .X(n25742) );
  nand_x1_sg U72623 ( .A(n57502), .B(n57019), .X(n25741) );
  nand_x2_sg U72624 ( .A(n25771), .B(n25772), .X(n25767) );
  nand_x1_sg U72625 ( .A(n57499), .B(n56801), .X(n25772) );
  nand_x1_sg U72626 ( .A(n57502), .B(n51511), .X(n25771) );
  nand_x2_sg U72627 ( .A(n25801), .B(n25802), .X(n25797) );
  nand_x1_sg U72628 ( .A(n57499), .B(n51353), .X(n25802) );
  nand_x1_sg U72629 ( .A(n57502), .B(n57035), .X(n25801) );
  nand_x2_sg U72630 ( .A(n25831), .B(n25832), .X(n25827) );
  nand_x1_sg U72631 ( .A(n57499), .B(n51289), .X(n25832) );
  nand_x1_sg U72632 ( .A(n57502), .B(n47755), .X(n25831) );
  nand_x2_sg U72633 ( .A(n25861), .B(n25862), .X(n25857) );
  nand_x1_sg U72634 ( .A(n57499), .B(n56755), .X(n25862) );
  nand_x1_sg U72635 ( .A(n57502), .B(n51501), .X(n25861) );
  nand_x2_sg U72636 ( .A(n25891), .B(n25892), .X(n25887) );
  nand_x1_sg U72637 ( .A(n57499), .B(n51417), .X(n25892) );
  nand_x1_sg U72638 ( .A(n57502), .B(n57023), .X(n25891) );
  nand_x2_sg U72639 ( .A(n25921), .B(n25922), .X(n25917) );
  nand_x1_sg U72640 ( .A(n57499), .B(n56853), .X(n25922) );
  nand_x1_sg U72641 ( .A(n57502), .B(n51513), .X(n25921) );
  nand_x2_sg U72642 ( .A(n25951), .B(n25952), .X(n25947) );
  nand_x1_sg U72643 ( .A(n57499), .B(n47699), .X(n25952) );
  nand_x1_sg U72644 ( .A(n57502), .B(n57037), .X(n25951) );
  nand_x2_sg U72645 ( .A(n25982), .B(n25983), .X(n25978) );
  nand_x1_sg U72646 ( .A(n57499), .B(n51323), .X(n25983) );
  nand_x1_sg U72647 ( .A(n57502), .B(n57025), .X(n25982) );
  nand_x4_sg U72648 ( .A(n24164), .B(n24165), .X(n24161) );
  nand_x1_sg U72649 ( .A(n47727), .B(n57455), .X(n24165) );
  nand_x4_sg U72650 ( .A(n24169), .B(n24170), .X(n24167) );
  nand_x1_sg U72651 ( .A(n47729), .B(n57454), .X(n24170) );
  nand_x4_sg U72652 ( .A(n24174), .B(n24175), .X(n24172) );
  nand_x1_sg U72653 ( .A(n51459), .B(n57455), .X(n24175) );
  nand_x4_sg U72654 ( .A(n24179), .B(n24180), .X(n24177) );
  nand_x1_sg U72655 ( .A(n51475), .B(n57454), .X(n24180) );
  nand_x4_sg U72656 ( .A(n24184), .B(n24185), .X(n24182) );
  nand_x1_sg U72657 ( .A(n56905), .B(n57455), .X(n24185) );
  nand_x4_sg U72658 ( .A(n24189), .B(n24190), .X(n24187) );
  nand_x1_sg U72659 ( .A(n47731), .B(n57454), .X(n24190) );
  nand_x4_sg U72660 ( .A(n24194), .B(n24195), .X(n24192) );
  nand_x1_sg U72661 ( .A(n51461), .B(n57455), .X(n24195) );
  nand_x4_sg U72662 ( .A(n24199), .B(n24200), .X(n24197) );
  nand_x1_sg U72663 ( .A(n56891), .B(n57455), .X(n24200) );
  nand_x4_sg U72664 ( .A(n24204), .B(n24205), .X(n24202) );
  nand_x1_sg U72665 ( .A(n51477), .B(n57454), .X(n24205) );
  nand_x4_sg U72666 ( .A(n24209), .B(n24210), .X(n24207) );
  nand_x1_sg U72667 ( .A(n56907), .B(n57455), .X(n24210) );
  nand_x4_sg U72668 ( .A(n24214), .B(n24215), .X(n24212) );
  nand_x1_sg U72669 ( .A(n51463), .B(n57455), .X(n24215) );
  nand_x4_sg U72670 ( .A(n24219), .B(n24220), .X(n24217) );
  nand_x1_sg U72671 ( .A(n56893), .B(n57454), .X(n24220) );
  nand_x4_sg U72672 ( .A(n24224), .B(n24225), .X(n24222) );
  nand_x1_sg U72673 ( .A(n51479), .B(n57454), .X(n24225) );
  nand_x4_sg U72674 ( .A(n24229), .B(n24230), .X(n24227) );
  nand_x1_sg U72675 ( .A(n56909), .B(n57455), .X(n24230) );
  nand_x4_sg U72676 ( .A(n24234), .B(n24235), .X(n24232) );
  nand_x1_sg U72677 ( .A(n51481), .B(n57454), .X(n24235) );
  nand_x4_sg U72678 ( .A(n24239), .B(n24240), .X(n24237) );
  nand_x1_sg U72679 ( .A(n56911), .B(n57454), .X(n24240) );
  nand_x4_sg U72680 ( .A(n24244), .B(n24245), .X(n24242) );
  nand_x1_sg U72681 ( .A(n47739), .B(n57455), .X(n24245) );
  nand_x4_sg U72682 ( .A(n24249), .B(n24250), .X(n24247) );
  nand_x1_sg U72683 ( .A(n51487), .B(n57454), .X(n24250) );
  nand_x4_sg U72684 ( .A(n24254), .B(n24255), .X(n24252) );
  nand_x1_sg U72685 ( .A(n56915), .B(n57454), .X(n24255) );
  nand_x4_sg U72686 ( .A(n24267), .B(n24268), .X(n24257) );
  nand_x1_sg U72687 ( .A(n56895), .B(n57454), .X(n24268) );
  nand_x4_sg U72688 ( .A(n24273), .B(n24274), .X(n24270) );
  nand_x1_sg U72689 ( .A(n47721), .B(n57454), .X(n24274) );
  nand_x4_sg U72690 ( .A(n24278), .B(n24279), .X(n24276) );
  nand_x1_sg U72691 ( .A(n47723), .B(n57454), .X(n24279) );
  nand_x4_sg U72692 ( .A(n24283), .B(n24284), .X(n24281) );
  nand_x1_sg U72693 ( .A(n51453), .B(n57455), .X(n24284) );
  nand_x4_sg U72694 ( .A(n24288), .B(n24289), .X(n24286) );
  nand_x1_sg U72695 ( .A(n51465), .B(n57455), .X(n24289) );
  nand_x4_sg U72696 ( .A(n24293), .B(n24294), .X(n24291) );
  nand_x1_sg U72697 ( .A(n56897), .B(n57454), .X(n24294) );
  nand_x4_sg U72698 ( .A(n24298), .B(n24299), .X(n24296) );
  nand_x1_sg U72699 ( .A(n47725), .B(n57455), .X(n24299) );
  nand_x4_sg U72700 ( .A(n24303), .B(n24304), .X(n24301) );
  nand_x1_sg U72701 ( .A(n51455), .B(n57454), .X(n24304) );
  nand_x4_sg U72702 ( .A(n24308), .B(n24309), .X(n24306) );
  nand_x1_sg U72703 ( .A(n56885), .B(n57454), .X(n24309) );
  nand_x4_sg U72704 ( .A(n24313), .B(n24314), .X(n24311) );
  nand_x1_sg U72705 ( .A(n51467), .B(n57455), .X(n24314) );
  nand_x4_sg U72706 ( .A(n24318), .B(n24319), .X(n24316) );
  nand_x1_sg U72707 ( .A(n56899), .B(n57454), .X(n24319) );
  nand_x4_sg U72708 ( .A(n24323), .B(n24324), .X(n24321) );
  nand_x1_sg U72709 ( .A(n51457), .B(n57455), .X(n24324) );
  nand_x4_sg U72710 ( .A(n24328), .B(n24329), .X(n24326) );
  nand_x1_sg U72711 ( .A(n56887), .B(n57455), .X(n24329) );
  nand_x4_sg U72712 ( .A(n24333), .B(n24334), .X(n24331) );
  nand_x1_sg U72713 ( .A(n51469), .B(n57455), .X(n24334) );
  nand_x4_sg U72714 ( .A(n24338), .B(n24339), .X(n24336) );
  nand_x1_sg U72715 ( .A(n56901), .B(n57454), .X(n24339) );
  nand_x4_sg U72716 ( .A(n24343), .B(n24344), .X(n24341) );
  nand_x1_sg U72717 ( .A(n51471), .B(n57455), .X(n24344) );
  nand_x4_sg U72718 ( .A(n24348), .B(n24349), .X(n24346) );
  nand_x1_sg U72719 ( .A(n56903), .B(n57454), .X(n24349) );
  nand_x4_sg U72720 ( .A(n24353), .B(n24354), .X(n24351) );
  nand_x1_sg U72721 ( .A(n47737), .B(n57455), .X(n24354) );
  nand_x4_sg U72722 ( .A(n24358), .B(n24359), .X(n24356) );
  nand_x1_sg U72723 ( .A(n51485), .B(n57455), .X(n24359) );
  nand_x4_sg U72724 ( .A(n24363), .B(n24364), .X(n24361) );
  nand_x1_sg U72725 ( .A(n56913), .B(n57454), .X(n24364) );
  nand_x4_sg U72726 ( .A(n24376), .B(n24377), .X(n24366) );
  nand_x1_sg U72727 ( .A(n56889), .B(n57454), .X(n24377) );
  nand_x1_sg U72728 ( .A(n47767), .B(n57464), .X(n23203) );
  nand_x1_sg U72729 ( .A(n47769), .B(n57464), .X(n23210) );
  nand_x1_sg U72730 ( .A(n51535), .B(n57464), .X(n23215) );
  nand_x1_sg U72731 ( .A(n47771), .B(n57464), .X(n23230) );
  nand_x1_sg U72732 ( .A(n51537), .B(n57464), .X(n23235) );
  nand_x1_sg U72733 ( .A(n57057), .B(n57464), .X(n23240) );
  nand_x1_sg U72734 ( .A(n51539), .B(n57464), .X(n23255) );
  nand_x1_sg U72735 ( .A(n57059), .B(n57464), .X(n23260) );
  nand_x1_sg U72736 ( .A(n51541), .B(n57464), .X(n23275) );
  nand_x1_sg U72737 ( .A(n57061), .B(n57464), .X(n23280) );
  nand_x1_sg U72738 ( .A(n57067), .B(n57464), .X(n23285) );
  nand_x1_sg U72739 ( .A(n57063), .B(n57464), .X(n23300) );
  nand_x1_sg U72740 ( .A(n47761), .B(n57472), .X(n23311) );
  nand_x1_sg U72741 ( .A(n47763), .B(n57472), .X(n23318) );
  nand_x1_sg U72742 ( .A(n51527), .B(n57472), .X(n23323) );
  nand_x1_sg U72743 ( .A(n47765), .B(n57472), .X(n23338) );
  nand_x1_sg U72744 ( .A(n51529), .B(n57472), .X(n23343) );
  nand_x1_sg U72745 ( .A(n57049), .B(n57472), .X(n23348) );
  nand_x1_sg U72746 ( .A(n51531), .B(n57472), .X(n23363) );
  nand_x1_sg U72747 ( .A(n57051), .B(n57472), .X(n23368) );
  nand_x1_sg U72748 ( .A(n51533), .B(n57472), .X(n23383) );
  nand_x1_sg U72749 ( .A(n57053), .B(n57472), .X(n23388) );
  nand_x1_sg U72750 ( .A(n57065), .B(n57472), .X(n23393) );
  nand_x1_sg U72751 ( .A(n57055), .B(n57472), .X(n23408) );
  nand_x4_sg U72752 ( .A(n26050), .B(n26051), .X(n26049) );
  nand_x1_sg U72753 ( .A(n56935), .B(n26052), .X(n26050) );
  nor_x1_sg U72754 ( .A(n26078), .B(n26079), .X(n26077) );
  nor_x1_sg U72755 ( .A(n26179), .B(n26180), .X(n26178) );
  nand_x1_sg U72756 ( .A(n47511), .B(n57949), .X(n58123) );
  nand_x1_sg U72757 ( .A(n47727), .B(n57941), .X(n58124) );
  nand_x1_sg U72758 ( .A(n47513), .B(n57949), .X(n58118) );
  nand_x1_sg U72759 ( .A(n47729), .B(n57942), .X(n58119) );
  nand_x1_sg U72760 ( .A(n55233), .B(n57949), .X(n58115) );
  nand_x1_sg U72761 ( .A(n51459), .B(n57942), .X(n58116) );
  nand_x1_sg U72762 ( .A(n55235), .B(n57949), .X(n58111) );
  nand_x1_sg U72763 ( .A(n51475), .B(n57942), .X(n58112) );
  nand_x1_sg U72764 ( .A(n51163), .B(n57949), .X(n58107) );
  nand_x1_sg U72765 ( .A(n56905), .B(n57947), .X(n58108) );
  nand_x1_sg U72766 ( .A(n47515), .B(n57949), .X(n58104) );
  nand_x1_sg U72767 ( .A(n47731), .B(n57947), .X(n58105) );
  nand_x1_sg U72768 ( .A(n55237), .B(n57949), .X(n58101) );
  nand_x1_sg U72769 ( .A(n51461), .B(n57944), .X(n58102) );
  nand_x1_sg U72770 ( .A(n51165), .B(n57949), .X(n58098) );
  nand_x1_sg U72771 ( .A(n56891), .B(n57937), .X(n58099) );
  nand_x1_sg U72772 ( .A(n55239), .B(n57949), .X(n58094) );
  nand_x1_sg U72773 ( .A(n51477), .B(n57938), .X(n58095) );
  nand_x1_sg U72774 ( .A(n51167), .B(n57949), .X(n58090) );
  nand_x1_sg U72775 ( .A(n56907), .B(n57943), .X(n58091) );
  nand_x1_sg U72776 ( .A(n55241), .B(n57949), .X(n58087) );
  nand_x1_sg U72777 ( .A(n51463), .B(n57943), .X(n58088) );
  nand_x1_sg U72778 ( .A(n51169), .B(n57949), .X(n58084) );
  nand_x1_sg U72779 ( .A(n56893), .B(n57943), .X(n58085) );
  nand_x1_sg U72780 ( .A(n55243), .B(n57949), .X(n58080) );
  nand_x1_sg U72781 ( .A(n51479), .B(n57943), .X(n58081) );
  nand_x1_sg U72782 ( .A(n51171), .B(n57949), .X(n58076) );
  nand_x1_sg U72783 ( .A(n56909), .B(n57944), .X(n58077) );
  nand_x1_sg U72784 ( .A(n55247), .B(n57949), .X(n58073) );
  nand_x1_sg U72785 ( .A(n51481), .B(n57944), .X(n58074) );
  nand_x1_sg U72786 ( .A(n51177), .B(n57949), .X(n58070) );
  nand_x1_sg U72787 ( .A(n56911), .B(n57944), .X(n58071) );
  nand_x1_sg U72788 ( .A(n47519), .B(n57949), .X(n58067) );
  nand_x1_sg U72789 ( .A(n47739), .B(n57929), .X(n58068) );
  nand_x1_sg U72790 ( .A(n55251), .B(n57949), .X(n58063) );
  nand_x1_sg U72791 ( .A(n51487), .B(n57951), .X(n58064) );
  nand_x1_sg U72792 ( .A(n51181), .B(n57949), .X(n58059) );
  nand_x1_sg U72793 ( .A(n56915), .B(n57951), .X(n58060) );
  nand_x1_sg U72794 ( .A(n51173), .B(n57949), .X(n58056) );
  nand_x1_sg U72795 ( .A(n56895), .B(n57948), .X(n58057) );
  nand_x1_sg U72796 ( .A(n47507), .B(n57949), .X(n58053) );
  nand_x1_sg U72797 ( .A(n47721), .B(n57951), .X(n58054) );
  nand_x1_sg U72798 ( .A(n51151), .B(n57949), .X(n58048) );
  nand_x1_sg U72799 ( .A(n47723), .B(n57940), .X(n58049) );
  nand_x1_sg U72800 ( .A(n55221), .B(n57949), .X(n58045) );
  nand_x1_sg U72801 ( .A(n51453), .B(n57933), .X(n58046) );
  nand_x1_sg U72802 ( .A(n55223), .B(n57949), .X(n58041) );
  nand_x1_sg U72803 ( .A(n51465), .B(n57934), .X(n58042) );
  nand_x1_sg U72804 ( .A(n51153), .B(n57949), .X(n58037) );
  nand_x1_sg U72805 ( .A(n56897), .B(n57939), .X(n58038) );
  nand_x1_sg U72806 ( .A(n47509), .B(n57949), .X(n58034) );
  nand_x1_sg U72807 ( .A(n47725), .B(n57945), .X(n58035) );
  nand_x1_sg U72808 ( .A(n55225), .B(n57949), .X(n58031) );
  nand_x1_sg U72809 ( .A(n51455), .B(n57945), .X(n58032) );
  nand_x1_sg U72810 ( .A(n51155), .B(n57949), .X(n58028) );
  nand_x1_sg U72811 ( .A(n56885), .B(n57945), .X(n58029) );
  nand_x1_sg U72812 ( .A(n55227), .B(n57949), .X(n58024) );
  nand_x1_sg U72813 ( .A(n51467), .B(n57941), .X(n58025) );
  nand_x1_sg U72814 ( .A(n51157), .B(n57949), .X(n58020) );
  nand_x1_sg U72815 ( .A(n56899), .B(n57942), .X(n58021) );
  nand_x1_sg U72816 ( .A(n55229), .B(n57949), .X(n58017) );
  nand_x1_sg U72817 ( .A(n51457), .B(n57945), .X(n58018) );
  nand_x1_sg U72818 ( .A(n51159), .B(n57949), .X(n58014) );
  nand_x1_sg U72819 ( .A(n56887), .B(n57948), .X(n58015) );
  nand_x1_sg U72820 ( .A(n55231), .B(n57949), .X(n58010) );
  nand_x1_sg U72821 ( .A(n51469), .B(n57948), .X(n58011) );
  nand_x1_sg U72822 ( .A(n51161), .B(n57949), .X(n58006) );
  nand_x1_sg U72823 ( .A(n56901), .B(n57936), .X(n58007) );
  nand_x1_sg U72824 ( .A(n55245), .B(n57949), .X(n58003) );
  nand_x1_sg U72825 ( .A(n51471), .B(n57930), .X(n58004) );
  nand_x1_sg U72826 ( .A(n51175), .B(n57949), .X(n58000) );
  nand_x1_sg U72827 ( .A(n56903), .B(n57951), .X(n58001) );
  nand_x1_sg U72828 ( .A(n47517), .B(n57949), .X(n57997) );
  nand_x1_sg U72829 ( .A(n47737), .B(n57935), .X(n57998) );
  nand_x1_sg U72830 ( .A(n55249), .B(n57949), .X(n57993) );
  nand_x1_sg U72831 ( .A(n51485), .B(n57948), .X(n57994) );
  nand_x1_sg U72832 ( .A(n51179), .B(n57949), .X(n57989) );
  nand_x1_sg U72833 ( .A(n56913), .B(n57931), .X(n57990) );
  nand_x1_sg U72834 ( .A(n47613), .B(n57949), .X(n57985) );
  nand_x1_sg U72835 ( .A(n56889), .B(n57932), .X(n57986) );
  nand_x4_sg U72836 ( .A(n22757), .B(n58580), .X(n22397) );
  nand_x1_sg U72837 ( .A(n47533), .B(n57865), .X(n22757) );
  nor_x1_sg U72838 ( .A(n57331), .B(n58650), .X(n58579) );
  nand_x4_sg U72839 ( .A(n22771), .B(n58578), .X(n22398) );
  nand_x1_sg U72840 ( .A(n56697), .B(n57865), .X(n22771) );
  nor_x1_sg U72841 ( .A(n57332), .B(n58576), .X(n58577) );
  nand_x4_sg U72842 ( .A(n22782), .B(n58575), .X(n22399) );
  nand_x1_sg U72843 ( .A(n47649), .B(n57865), .X(n22782) );
  nor_x1_sg U72844 ( .A(n57333), .B(n68577), .X(n58574) );
  nand_x4_sg U72845 ( .A(n22793), .B(n58573), .X(n22400) );
  nand_x1_sg U72846 ( .A(n51277), .B(n57865), .X(n22793) );
  nor_x1_sg U72847 ( .A(n57334), .B(n68578), .X(n58572) );
  nand_x4_sg U72848 ( .A(n22804), .B(n58571), .X(n22401) );
  nand_x1_sg U72849 ( .A(n56739), .B(n57865), .X(n22804) );
  nor_x1_sg U72850 ( .A(n57342), .B(n58569), .X(n58570) );
  nand_x4_sg U72851 ( .A(n22815), .B(n58568), .X(n22402) );
  nand_x1_sg U72852 ( .A(n47535), .B(n57865), .X(n22815) );
  nor_x1_sg U72853 ( .A(n57342), .B(n68579), .X(n58567) );
  nand_x4_sg U72854 ( .A(n22826), .B(n58566), .X(n22403) );
  nand_x1_sg U72855 ( .A(n47651), .B(n57865), .X(n22826) );
  nor_x1_sg U72856 ( .A(n57341), .B(n68580), .X(n58565) );
  nand_x4_sg U72857 ( .A(n22837), .B(n58564), .X(n22404) );
  nand_x1_sg U72858 ( .A(n51235), .B(n57865), .X(n22837) );
  nor_x1_sg U72859 ( .A(n57341), .B(n58562), .X(n58563) );
  nand_x4_sg U72860 ( .A(n22848), .B(n58561), .X(n22405) );
  nand_x1_sg U72861 ( .A(n47671), .B(n57865), .X(n22848) );
  nor_x1_sg U72862 ( .A(n57340), .B(n68581), .X(n58560) );
  nand_x4_sg U72863 ( .A(n22859), .B(n58559), .X(n22406) );
  nand_x1_sg U72864 ( .A(n51377), .B(n57865), .X(n22859) );
  nor_x1_sg U72865 ( .A(n57340), .B(n68582), .X(n58558) );
  nand_x4_sg U72866 ( .A(n22870), .B(n58557), .X(n22407) );
  nand_x1_sg U72867 ( .A(n47665), .B(n57867), .X(n22870) );
  nor_x1_sg U72868 ( .A(n57339), .B(n58555), .X(n58556) );
  nand_x4_sg U72869 ( .A(n22881), .B(n58554), .X(n22408) );
  nand_x1_sg U72870 ( .A(n51317), .B(n57865), .X(n22881) );
  nor_x1_sg U72871 ( .A(n57339), .B(n68583), .X(n58553) );
  nand_x4_sg U72872 ( .A(n22892), .B(n58552), .X(n22409) );
  nand_x1_sg U72873 ( .A(n51379), .B(n57867), .X(n22892) );
  nor_x1_sg U72874 ( .A(n58630), .B(n68584), .X(n58551) );
  nand_x4_sg U72875 ( .A(n22903), .B(n58550), .X(n22410) );
  nand_x1_sg U72876 ( .A(n56823), .B(n57865), .X(n22903) );
  nor_x1_sg U72877 ( .A(n58630), .B(n58548), .X(n58549) );
  nand_x4_sg U72878 ( .A(n22914), .B(n58547), .X(n22411) );
  nand_x1_sg U72879 ( .A(n47667), .B(n29329), .X(n22914) );
  nor_x1_sg U72880 ( .A(n57341), .B(n58545), .X(n58546) );
  nand_x4_sg U72881 ( .A(n22925), .B(n58544), .X(n22412) );
  nand_x1_sg U72882 ( .A(n51319), .B(n57865), .X(n22925) );
  nor_x1_sg U72883 ( .A(n57342), .B(n58542), .X(n58543) );
  nand_x4_sg U72884 ( .A(n22936), .B(n58541), .X(n22413) );
  nand_x1_sg U72885 ( .A(n51423), .B(n57865), .X(n22936) );
  nor_x1_sg U72886 ( .A(n57339), .B(n68585), .X(n58540) );
  nand_x4_sg U72887 ( .A(n22947), .B(n58539), .X(n22414) );
  nand_x1_sg U72888 ( .A(n47707), .B(n57865), .X(n22947) );
  nor_x1_sg U72889 ( .A(n57340), .B(n68586), .X(n58538) );
  nand_x4_sg U72890 ( .A(n22958), .B(n58537), .X(n22415) );
  nand_x1_sg U72891 ( .A(n56859), .B(n57865), .X(n22958) );
  nor_x1_sg U72892 ( .A(n58630), .B(n58535), .X(n58536) );
  nand_x4_sg U72893 ( .A(n22969), .B(n58534), .X(n22416) );
  nand_x1_sg U72894 ( .A(n51329), .B(n57865), .X(n22969) );
  nor_x1_sg U72895 ( .A(n57338), .B(n58532), .X(n58533) );
  nand_x4_sg U72896 ( .A(n22985), .B(n58531), .X(n22422) );
  nand_x1_sg U72897 ( .A(n47549), .B(n57865), .X(n22985) );
  nor_x1_sg U72898 ( .A(n57338), .B(n58611), .X(n58530) );
  nand_x4_sg U72899 ( .A(n22998), .B(n58529), .X(n22423) );
  nand_x1_sg U72900 ( .A(n47659), .B(n57865), .X(n22998) );
  nor_x1_sg U72901 ( .A(n57337), .B(n58527), .X(n58528) );
  nand_x4_sg U72902 ( .A(n23009), .B(n58526), .X(n22424) );
  nand_x1_sg U72903 ( .A(n51299), .B(n57865), .X(n23009) );
  nor_x1_sg U72904 ( .A(n57337), .B(n68477), .X(n58525) );
  nand_x4_sg U72905 ( .A(n23020), .B(n58524), .X(n22425) );
  nand_x1_sg U72906 ( .A(n51361), .B(n57865), .X(n23020) );
  nor_x1_sg U72907 ( .A(n57336), .B(n68478), .X(n58523) );
  nand_x4_sg U72908 ( .A(n23031), .B(n58522), .X(n22426) );
  nand_x1_sg U72909 ( .A(n56809), .B(n57865), .X(n23031) );
  nor_x1_sg U72910 ( .A(n57336), .B(n58520), .X(n58521) );
  nand_x4_sg U72911 ( .A(n23042), .B(n58519), .X(n22427) );
  nand_x1_sg U72912 ( .A(n47551), .B(n57865), .X(n23042) );
  nor_x1_sg U72913 ( .A(n57335), .B(n68479), .X(n58518) );
  nand_x4_sg U72914 ( .A(n23053), .B(n58517), .X(n22428) );
  nand_x1_sg U72915 ( .A(n47661), .B(n57865), .X(n23053) );
  nor_x1_sg U72916 ( .A(n57335), .B(n68480), .X(n58516) );
  nand_x4_sg U72917 ( .A(n23064), .B(n58515), .X(n22429) );
  nand_x1_sg U72918 ( .A(n51301), .B(n57865), .X(n23064) );
  nor_x1_sg U72919 ( .A(n57337), .B(n58513), .X(n58514) );
  nand_x4_sg U72920 ( .A(n23075), .B(n58512), .X(n22430) );
  nand_x1_sg U72921 ( .A(n47669), .B(n57865), .X(n23075) );
  nor_x1_sg U72922 ( .A(n57338), .B(n68481), .X(n58511) );
  nand_x4_sg U72923 ( .A(n23086), .B(n58510), .X(n22431) );
  nand_x1_sg U72924 ( .A(n51363), .B(n57865), .X(n23086) );
  nor_x1_sg U72925 ( .A(n57335), .B(n68482), .X(n58509) );
  nand_x4_sg U72926 ( .A(n23097), .B(n58508), .X(n22432) );
  nand_x1_sg U72927 ( .A(n47663), .B(n57865), .X(n23097) );
  nor_x1_sg U72928 ( .A(n57336), .B(n58506), .X(n58507) );
  nand_x4_sg U72929 ( .A(n23108), .B(n58505), .X(n22433) );
  nand_x1_sg U72930 ( .A(n51303), .B(n57865), .X(n23108) );
  nor_x1_sg U72931 ( .A(n57334), .B(n68483), .X(n58504) );
  nand_x4_sg U72932 ( .A(n23119), .B(n58503), .X(n22434) );
  nand_x1_sg U72933 ( .A(n51257), .B(n57865), .X(n23119) );
  nor_x1_sg U72934 ( .A(n57334), .B(n68484), .X(n58502) );
  nand_x4_sg U72935 ( .A(n23130), .B(n58501), .X(n22435) );
  nand_x1_sg U72936 ( .A(n56719), .B(n57865), .X(n23130) );
  nor_x1_sg U72937 ( .A(n57333), .B(n58499), .X(n58500) );
  nand_x4_sg U72938 ( .A(n23141), .B(n58498), .X(n22436) );
  nand_x1_sg U72939 ( .A(n47629), .B(n57865), .X(n23141) );
  nor_x1_sg U72940 ( .A(n57333), .B(n58496), .X(n58497) );
  nand_x4_sg U72941 ( .A(n23152), .B(n58495), .X(n22437) );
  nand_x1_sg U72942 ( .A(n51213), .B(n57865), .X(n23152) );
  nor_x1_sg U72943 ( .A(n57332), .B(n58493), .X(n58494) );
  nand_x4_sg U72944 ( .A(n23163), .B(n58492), .X(n22438) );
  nand_x1_sg U72945 ( .A(n47683), .B(n57865), .X(n23163) );
  nor_x1_sg U72946 ( .A(n57332), .B(n68485), .X(n58491) );
  nand_x4_sg U72947 ( .A(n23174), .B(n58490), .X(n22439) );
  nand_x1_sg U72948 ( .A(n51393), .B(n57865), .X(n23174) );
  nor_x1_sg U72949 ( .A(n57331), .B(n68486), .X(n58489) );
  nand_x4_sg U72950 ( .A(n23185), .B(n58488), .X(n22440) );
  nand_x1_sg U72951 ( .A(n56835), .B(n57865), .X(n23185) );
  nor_x1_sg U72952 ( .A(n57331), .B(n67307), .X(n58487) );
  nand_x4_sg U72953 ( .A(n23196), .B(n58486), .X(n22441) );
  nand_x1_sg U72954 ( .A(n56673), .B(n57865), .X(n23196) );
  nor_x1_sg U72955 ( .A(n57330), .B(n58484), .X(n58485) );
  nor_x1_sg U72956 ( .A(n68141), .B(n26253), .X(\filter_0/n10508 ) );
  nor_x1_sg U72957 ( .A(n68140), .B(n26253), .X(\filter_0/n10504 ) );
  nor_x1_sg U72958 ( .A(n68139), .B(n26253), .X(\filter_0/n10500 ) );
  nor_x1_sg U72959 ( .A(n68138), .B(n26253), .X(\filter_0/n10496 ) );
  nor_x1_sg U72960 ( .A(n68137), .B(n26253), .X(\filter_0/n10492 ) );
  nor_x1_sg U72961 ( .A(n68136), .B(n26253), .X(\filter_0/n10488 ) );
  nor_x1_sg U72962 ( .A(n68135), .B(n26253), .X(\filter_0/n10484 ) );
  nor_x1_sg U72963 ( .A(n68134), .B(n26253), .X(\filter_0/n10480 ) );
  nor_x1_sg U72964 ( .A(n68133), .B(n26253), .X(\filter_0/n10476 ) );
  nor_x1_sg U72965 ( .A(n68132), .B(n26253), .X(\filter_0/n10472 ) );
  nor_x1_sg U72966 ( .A(n68131), .B(n26253), .X(\filter_0/n10468 ) );
  nor_x1_sg U72967 ( .A(n68130), .B(n26253), .X(\filter_0/n10464 ) );
  nor_x1_sg U72968 ( .A(n68129), .B(n26253), .X(\filter_0/n10460 ) );
  nor_x1_sg U72969 ( .A(n68121), .B(n26254), .X(\filter_0/n10428 ) );
  nor_x1_sg U72970 ( .A(n68120), .B(n26254), .X(\filter_0/n10424 ) );
  nor_x1_sg U72971 ( .A(n68119), .B(n26254), .X(\filter_0/n10420 ) );
  nor_x1_sg U72972 ( .A(n68118), .B(n26254), .X(\filter_0/n10416 ) );
  nor_x1_sg U72973 ( .A(n68117), .B(n26254), .X(\filter_0/n10412 ) );
  nor_x1_sg U72974 ( .A(n68116), .B(n26254), .X(\filter_0/n10408 ) );
  nor_x1_sg U72975 ( .A(n68115), .B(n26254), .X(\filter_0/n10404 ) );
  nor_x1_sg U72976 ( .A(n68114), .B(n26254), .X(\filter_0/n10400 ) );
  nor_x1_sg U72977 ( .A(n68113), .B(n26254), .X(\filter_0/n10396 ) );
  nor_x1_sg U72978 ( .A(n68112), .B(n26254), .X(\filter_0/n10392 ) );
  nor_x1_sg U72979 ( .A(n68111), .B(n26254), .X(\filter_0/n10388 ) );
  nor_x1_sg U72980 ( .A(n68110), .B(n26254), .X(\filter_0/n10384 ) );
  nor_x1_sg U72981 ( .A(n68109), .B(n26254), .X(\filter_0/n10380 ) );
  nor_x1_sg U72982 ( .A(n68101), .B(n26255), .X(\filter_0/n10348 ) );
  nor_x1_sg U72983 ( .A(n68100), .B(n26255), .X(\filter_0/n10344 ) );
  nor_x1_sg U72984 ( .A(n68099), .B(n26255), .X(\filter_0/n10340 ) );
  nor_x1_sg U72985 ( .A(n68098), .B(n26255), .X(\filter_0/n10336 ) );
  nor_x1_sg U72986 ( .A(n68097), .B(n26255), .X(\filter_0/n10332 ) );
  nor_x1_sg U72987 ( .A(n68096), .B(n26255), .X(\filter_0/n10328 ) );
  nor_x1_sg U72988 ( .A(n68095), .B(n26255), .X(\filter_0/n10324 ) );
  nor_x1_sg U72989 ( .A(n68094), .B(n26255), .X(\filter_0/n10320 ) );
  nor_x1_sg U72990 ( .A(n68093), .B(n26255), .X(\filter_0/n10316 ) );
  nor_x1_sg U72991 ( .A(n68092), .B(n26255), .X(\filter_0/n10312 ) );
  nor_x1_sg U72992 ( .A(n68091), .B(n26255), .X(\filter_0/n10308 ) );
  nor_x1_sg U72993 ( .A(n68090), .B(n26255), .X(\filter_0/n10304 ) );
  nor_x1_sg U72994 ( .A(n68089), .B(n26255), .X(\filter_0/n10300 ) );
  nor_x1_sg U72995 ( .A(n68081), .B(n26256), .X(\filter_0/n10268 ) );
  nor_x1_sg U72996 ( .A(n68080), .B(n26256), .X(\filter_0/n10264 ) );
  nor_x1_sg U72997 ( .A(n68079), .B(n26256), .X(\filter_0/n10260 ) );
  nor_x1_sg U72998 ( .A(n68078), .B(n26256), .X(\filter_0/n10256 ) );
  nor_x1_sg U72999 ( .A(n68077), .B(n26256), .X(\filter_0/n10252 ) );
  nor_x1_sg U73000 ( .A(n68076), .B(n26256), .X(\filter_0/n10248 ) );
  nor_x1_sg U73001 ( .A(n68075), .B(n26256), .X(\filter_0/n10244 ) );
  nor_x1_sg U73002 ( .A(n68074), .B(n26256), .X(\filter_0/n10240 ) );
  nor_x1_sg U73003 ( .A(n68073), .B(n26256), .X(\filter_0/n10236 ) );
  nor_x1_sg U73004 ( .A(n68072), .B(n26256), .X(\filter_0/n10232 ) );
  nor_x1_sg U73005 ( .A(n68071), .B(n26256), .X(\filter_0/n10228 ) );
  nor_x1_sg U73006 ( .A(n68070), .B(n26256), .X(\filter_0/n10224 ) );
  nor_x1_sg U73007 ( .A(n68069), .B(n26256), .X(\filter_0/n10220 ) );
  nor_x1_sg U73008 ( .A(n67821), .B(n26024), .X(\filter_0/n9228 ) );
  nor_x1_sg U73009 ( .A(n67820), .B(n26024), .X(\filter_0/n9224 ) );
  nor_x1_sg U73010 ( .A(n67819), .B(n26024), .X(\filter_0/n9220 ) );
  nor_x1_sg U73011 ( .A(n67818), .B(n26024), .X(\filter_0/n9216 ) );
  nor_x1_sg U73012 ( .A(n67817), .B(n26024), .X(\filter_0/n9212 ) );
  nor_x1_sg U73013 ( .A(n67816), .B(n26024), .X(\filter_0/n9208 ) );
  nor_x1_sg U73014 ( .A(n67815), .B(n26024), .X(\filter_0/n9204 ) );
  nor_x1_sg U73015 ( .A(n67814), .B(n26024), .X(\filter_0/n9200 ) );
  nor_x1_sg U73016 ( .A(n67813), .B(n26024), .X(\filter_0/n9196 ) );
  nor_x1_sg U73017 ( .A(n67812), .B(n26024), .X(\filter_0/n9192 ) );
  nor_x1_sg U73018 ( .A(n67811), .B(n26024), .X(\filter_0/n9188 ) );
  nor_x1_sg U73019 ( .A(n67810), .B(n26024), .X(\filter_0/n9184 ) );
  nor_x1_sg U73020 ( .A(n67809), .B(n26024), .X(\filter_0/n9180 ) );
  nor_x1_sg U73021 ( .A(n67801), .B(n26025), .X(\filter_0/n9148 ) );
  nor_x1_sg U73022 ( .A(n67800), .B(n26025), .X(\filter_0/n9144 ) );
  nor_x1_sg U73023 ( .A(n67799), .B(n26025), .X(\filter_0/n9140 ) );
  nor_x1_sg U73024 ( .A(n67798), .B(n26025), .X(\filter_0/n9136 ) );
  nor_x1_sg U73025 ( .A(n67797), .B(n26025), .X(\filter_0/n9132 ) );
  nor_x1_sg U73026 ( .A(n67796), .B(n26025), .X(\filter_0/n9128 ) );
  nor_x1_sg U73027 ( .A(n67795), .B(n26025), .X(\filter_0/n9124 ) );
  nor_x1_sg U73028 ( .A(n67794), .B(n26025), .X(\filter_0/n9120 ) );
  nor_x1_sg U73029 ( .A(n67793), .B(n26025), .X(\filter_0/n9116 ) );
  nor_x1_sg U73030 ( .A(n67792), .B(n26025), .X(\filter_0/n9112 ) );
  nor_x1_sg U73031 ( .A(n67791), .B(n26025), .X(\filter_0/n9108 ) );
  nor_x1_sg U73032 ( .A(n67790), .B(n26025), .X(\filter_0/n9104 ) );
  nor_x1_sg U73033 ( .A(n67789), .B(n26025), .X(\filter_0/n9100 ) );
  nor_x1_sg U73034 ( .A(n67781), .B(n26026), .X(\filter_0/n9068 ) );
  nor_x1_sg U73035 ( .A(n67780), .B(n26026), .X(\filter_0/n9064 ) );
  nor_x1_sg U73036 ( .A(n67779), .B(n26026), .X(\filter_0/n9060 ) );
  nor_x1_sg U73037 ( .A(n67778), .B(n26026), .X(\filter_0/n9056 ) );
  nor_x1_sg U73038 ( .A(n67777), .B(n26026), .X(\filter_0/n9052 ) );
  nor_x1_sg U73039 ( .A(n67776), .B(n26026), .X(\filter_0/n9048 ) );
  nor_x1_sg U73040 ( .A(n67775), .B(n26026), .X(\filter_0/n9044 ) );
  nor_x1_sg U73041 ( .A(n67774), .B(n26026), .X(\filter_0/n9040 ) );
  nor_x1_sg U73042 ( .A(n67773), .B(n26026), .X(\filter_0/n9036 ) );
  nor_x1_sg U73043 ( .A(n67772), .B(n26026), .X(\filter_0/n9032 ) );
  nor_x1_sg U73044 ( .A(n67771), .B(n26026), .X(\filter_0/n9028 ) );
  nor_x1_sg U73045 ( .A(n67770), .B(n26026), .X(\filter_0/n9024 ) );
  nor_x1_sg U73046 ( .A(n67769), .B(n26026), .X(\filter_0/n9020 ) );
  nor_x1_sg U73047 ( .A(n67761), .B(n26027), .X(\filter_0/n8988 ) );
  nor_x1_sg U73048 ( .A(n67760), .B(n26027), .X(\filter_0/n8984 ) );
  nor_x1_sg U73049 ( .A(n67759), .B(n26027), .X(\filter_0/n8980 ) );
  nor_x1_sg U73050 ( .A(n67758), .B(n26027), .X(\filter_0/n8976 ) );
  nor_x1_sg U73051 ( .A(n67757), .B(n26027), .X(\filter_0/n8972 ) );
  nor_x1_sg U73052 ( .A(n67756), .B(n26027), .X(\filter_0/n8968 ) );
  nor_x1_sg U73053 ( .A(n67755), .B(n26027), .X(\filter_0/n8964 ) );
  nor_x1_sg U73054 ( .A(n67754), .B(n26027), .X(\filter_0/n8960 ) );
  nor_x1_sg U73055 ( .A(n67753), .B(n26027), .X(\filter_0/n8956 ) );
  nor_x1_sg U73056 ( .A(n67752), .B(n26027), .X(\filter_0/n8952 ) );
  nor_x1_sg U73057 ( .A(n67751), .B(n26027), .X(\filter_0/n8948 ) );
  nor_x1_sg U73058 ( .A(n67750), .B(n26027), .X(\filter_0/n8944 ) );
  nor_x1_sg U73059 ( .A(n67749), .B(n26027), .X(\filter_0/n8940 ) );
  nor_x1_sg U73060 ( .A(n68221), .B(n26249), .X(\filter_0/n10828 ) );
  nor_x1_sg U73061 ( .A(n68220), .B(n26249), .X(\filter_0/n10824 ) );
  nor_x1_sg U73062 ( .A(n68219), .B(n26249), .X(\filter_0/n10820 ) );
  nor_x1_sg U73063 ( .A(n68218), .B(n26249), .X(\filter_0/n10816 ) );
  nor_x1_sg U73064 ( .A(n68217), .B(n26249), .X(\filter_0/n10812 ) );
  nor_x1_sg U73065 ( .A(n68216), .B(n26249), .X(\filter_0/n10808 ) );
  nor_x1_sg U73066 ( .A(n68215), .B(n26249), .X(\filter_0/n10804 ) );
  nor_x1_sg U73067 ( .A(n68214), .B(n26249), .X(\filter_0/n10800 ) );
  nor_x1_sg U73068 ( .A(n68213), .B(n26249), .X(\filter_0/n10796 ) );
  nor_x1_sg U73069 ( .A(n68212), .B(n26249), .X(\filter_0/n10792 ) );
  nor_x1_sg U73070 ( .A(n68211), .B(n26249), .X(\filter_0/n10788 ) );
  nor_x1_sg U73071 ( .A(n68210), .B(n26249), .X(\filter_0/n10784 ) );
  nor_x1_sg U73072 ( .A(n68209), .B(n26249), .X(\filter_0/n10780 ) );
  nor_x1_sg U73073 ( .A(n68201), .B(n26250), .X(\filter_0/n10748 ) );
  nor_x1_sg U73074 ( .A(n68200), .B(n26250), .X(\filter_0/n10744 ) );
  nor_x1_sg U73075 ( .A(n68199), .B(n26250), .X(\filter_0/n10740 ) );
  nor_x1_sg U73076 ( .A(n68198), .B(n26250), .X(\filter_0/n10736 ) );
  nor_x1_sg U73077 ( .A(n68197), .B(n26250), .X(\filter_0/n10732 ) );
  nor_x1_sg U73078 ( .A(n68196), .B(n26250), .X(\filter_0/n10728 ) );
  nor_x1_sg U73079 ( .A(n68195), .B(n26250), .X(\filter_0/n10724 ) );
  nor_x1_sg U73080 ( .A(n68194), .B(n26250), .X(\filter_0/n10720 ) );
  nor_x1_sg U73081 ( .A(n68193), .B(n26250), .X(\filter_0/n10716 ) );
  nor_x1_sg U73082 ( .A(n68192), .B(n26250), .X(\filter_0/n10712 ) );
  nor_x1_sg U73083 ( .A(n68191), .B(n26250), .X(\filter_0/n10708 ) );
  nor_x1_sg U73084 ( .A(n68190), .B(n26250), .X(\filter_0/n10704 ) );
  nor_x1_sg U73085 ( .A(n68189), .B(n26250), .X(\filter_0/n10700 ) );
  nor_x1_sg U73086 ( .A(n68181), .B(n26251), .X(\filter_0/n10668 ) );
  nor_x1_sg U73087 ( .A(n68180), .B(n26251), .X(\filter_0/n10664 ) );
  nor_x1_sg U73088 ( .A(n68179), .B(n26251), .X(\filter_0/n10660 ) );
  nor_x1_sg U73089 ( .A(n68178), .B(n26251), .X(\filter_0/n10656 ) );
  nor_x1_sg U73090 ( .A(n68177), .B(n26251), .X(\filter_0/n10652 ) );
  nor_x1_sg U73091 ( .A(n68176), .B(n26251), .X(\filter_0/n10648 ) );
  nor_x1_sg U73092 ( .A(n68175), .B(n26251), .X(\filter_0/n10644 ) );
  nor_x1_sg U73093 ( .A(n68174), .B(n26251), .X(\filter_0/n10640 ) );
  nor_x1_sg U73094 ( .A(n68173), .B(n26251), .X(\filter_0/n10636 ) );
  nor_x1_sg U73095 ( .A(n68172), .B(n26251), .X(\filter_0/n10632 ) );
  nor_x1_sg U73096 ( .A(n68171), .B(n26251), .X(\filter_0/n10628 ) );
  nor_x1_sg U73097 ( .A(n68170), .B(n26251), .X(\filter_0/n10624 ) );
  nor_x1_sg U73098 ( .A(n68169), .B(n26251), .X(\filter_0/n10620 ) );
  nor_x1_sg U73099 ( .A(n68161), .B(n26252), .X(\filter_0/n10588 ) );
  nor_x1_sg U73100 ( .A(n68160), .B(n26252), .X(\filter_0/n10584 ) );
  nor_x1_sg U73101 ( .A(n68159), .B(n26252), .X(\filter_0/n10580 ) );
  nor_x1_sg U73102 ( .A(n68158), .B(n26252), .X(\filter_0/n10576 ) );
  nor_x1_sg U73103 ( .A(n68157), .B(n26252), .X(\filter_0/n10572 ) );
  nor_x1_sg U73104 ( .A(n68156), .B(n26252), .X(\filter_0/n10568 ) );
  nor_x1_sg U73105 ( .A(n68155), .B(n26252), .X(\filter_0/n10564 ) );
  nor_x1_sg U73106 ( .A(n68154), .B(n26252), .X(\filter_0/n10560 ) );
  nor_x1_sg U73107 ( .A(n68153), .B(n26252), .X(\filter_0/n10556 ) );
  nor_x1_sg U73108 ( .A(n68152), .B(n26252), .X(\filter_0/n10552 ) );
  nor_x1_sg U73109 ( .A(n68151), .B(n26252), .X(\filter_0/n10548 ) );
  nor_x1_sg U73110 ( .A(n68150), .B(n26252), .X(\filter_0/n10544 ) );
  nor_x1_sg U73111 ( .A(n68149), .B(n26252), .X(\filter_0/n10540 ) );
  nor_x1_sg U73112 ( .A(n68061), .B(n26257), .X(\filter_0/n10188 ) );
  nor_x1_sg U73113 ( .A(n68060), .B(n26257), .X(\filter_0/n10184 ) );
  nor_x1_sg U73114 ( .A(n68059), .B(n26257), .X(\filter_0/n10180 ) );
  nor_x1_sg U73115 ( .A(n68058), .B(n26257), .X(\filter_0/n10176 ) );
  nor_x1_sg U73116 ( .A(n68057), .B(n26257), .X(\filter_0/n10172 ) );
  nor_x1_sg U73117 ( .A(n68056), .B(n26257), .X(\filter_0/n10168 ) );
  nor_x1_sg U73118 ( .A(n68055), .B(n26257), .X(\filter_0/n10164 ) );
  nor_x1_sg U73119 ( .A(n68054), .B(n26257), .X(\filter_0/n10160 ) );
  nor_x1_sg U73120 ( .A(n68053), .B(n26257), .X(\filter_0/n10156 ) );
  nor_x1_sg U73121 ( .A(n68052), .B(n26257), .X(\filter_0/n10152 ) );
  nor_x1_sg U73122 ( .A(n68051), .B(n26257), .X(\filter_0/n10148 ) );
  nor_x1_sg U73123 ( .A(n68050), .B(n26257), .X(\filter_0/n10144 ) );
  nor_x1_sg U73124 ( .A(n68049), .B(n26257), .X(\filter_0/n10140 ) );
  nor_x1_sg U73125 ( .A(n68041), .B(n26259), .X(\filter_0/n10108 ) );
  nor_x1_sg U73126 ( .A(n68040), .B(n26259), .X(\filter_0/n10104 ) );
  nor_x1_sg U73127 ( .A(n68039), .B(n26259), .X(\filter_0/n10100 ) );
  nor_x1_sg U73128 ( .A(n68038), .B(n26259), .X(\filter_0/n10096 ) );
  nor_x1_sg U73129 ( .A(n68037), .B(n26259), .X(\filter_0/n10092 ) );
  nor_x1_sg U73130 ( .A(n68036), .B(n26259), .X(\filter_0/n10088 ) );
  nor_x1_sg U73131 ( .A(n68035), .B(n26259), .X(\filter_0/n10084 ) );
  nor_x1_sg U73132 ( .A(n68034), .B(n26259), .X(\filter_0/n10080 ) );
  nor_x1_sg U73133 ( .A(n68033), .B(n26259), .X(\filter_0/n10076 ) );
  nor_x1_sg U73134 ( .A(n68032), .B(n26259), .X(\filter_0/n10072 ) );
  nor_x1_sg U73135 ( .A(n68031), .B(n26259), .X(\filter_0/n10068 ) );
  nor_x1_sg U73136 ( .A(n68030), .B(n26259), .X(\filter_0/n10064 ) );
  nor_x1_sg U73137 ( .A(n68029), .B(n26259), .X(\filter_0/n10060 ) );
  nor_x1_sg U73138 ( .A(n68026), .B(n26006), .X(\filter_0/n10048 ) );
  nor_x1_sg U73139 ( .A(n68025), .B(n26006), .X(\filter_0/n10044 ) );
  nor_x1_sg U73140 ( .A(n68024), .B(n26006), .X(\filter_0/n10040 ) );
  nor_x1_sg U73141 ( .A(n68023), .B(n26006), .X(\filter_0/n10036 ) );
  nor_x1_sg U73142 ( .A(n68022), .B(n26006), .X(\filter_0/n10032 ) );
  nor_x1_sg U73143 ( .A(n68021), .B(n26006), .X(\filter_0/n10028 ) );
  nor_x1_sg U73144 ( .A(n68020), .B(n26006), .X(\filter_0/n10024 ) );
  nor_x1_sg U73145 ( .A(n68019), .B(n26006), .X(\filter_0/n10020 ) );
  nor_x1_sg U73146 ( .A(n68018), .B(n26006), .X(\filter_0/n10016 ) );
  nor_x1_sg U73147 ( .A(n68017), .B(n26006), .X(\filter_0/n10012 ) );
  nor_x1_sg U73148 ( .A(n68016), .B(n26006), .X(\filter_0/n10008 ) );
  nor_x1_sg U73149 ( .A(n68009), .B(n26006), .X(\filter_0/n9980 ) );
  nor_x1_sg U73150 ( .A(n68008), .B(n26006), .X(\filter_0/n9976 ) );
  nor_x1_sg U73151 ( .A(n68007), .B(n26006), .X(\filter_0/n9972 ) );
  nor_x1_sg U73152 ( .A(n68001), .B(n26007), .X(\filter_0/n9948 ) );
  nor_x1_sg U73153 ( .A(n68000), .B(n26007), .X(\filter_0/n9944 ) );
  nor_x1_sg U73154 ( .A(n67999), .B(n26007), .X(\filter_0/n9940 ) );
  nor_x1_sg U73155 ( .A(n67998), .B(n26007), .X(\filter_0/n9936 ) );
  nor_x1_sg U73156 ( .A(n67997), .B(n26007), .X(\filter_0/n9932 ) );
  nor_x1_sg U73157 ( .A(n67996), .B(n26007), .X(\filter_0/n9928 ) );
  nor_x1_sg U73158 ( .A(n67995), .B(n26007), .X(\filter_0/n9924 ) );
  nor_x1_sg U73159 ( .A(n67994), .B(n26007), .X(\filter_0/n9920 ) );
  nor_x1_sg U73160 ( .A(n67993), .B(n26007), .X(\filter_0/n9916 ) );
  nor_x1_sg U73161 ( .A(n67992), .B(n26007), .X(\filter_0/n9912 ) );
  nor_x1_sg U73162 ( .A(n67991), .B(n26007), .X(\filter_0/n9908 ) );
  nor_x1_sg U73163 ( .A(n67990), .B(n26007), .X(\filter_0/n9904 ) );
  nor_x1_sg U73164 ( .A(n67989), .B(n26007), .X(\filter_0/n9900 ) );
  nor_x1_sg U73165 ( .A(n67901), .B(n26016), .X(\filter_0/n9548 ) );
  nor_x1_sg U73166 ( .A(n67900), .B(n26016), .X(\filter_0/n9544 ) );
  nor_x1_sg U73167 ( .A(n67899), .B(n26016), .X(\filter_0/n9540 ) );
  nor_x1_sg U73168 ( .A(n67898), .B(n26016), .X(\filter_0/n9536 ) );
  nor_x1_sg U73169 ( .A(n67897), .B(n26016), .X(\filter_0/n9532 ) );
  nor_x1_sg U73170 ( .A(n67896), .B(n26016), .X(\filter_0/n9528 ) );
  nor_x1_sg U73171 ( .A(n67895), .B(n26016), .X(\filter_0/n9524 ) );
  nor_x1_sg U73172 ( .A(n67894), .B(n26016), .X(\filter_0/n9520 ) );
  nor_x1_sg U73173 ( .A(n67893), .B(n26016), .X(\filter_0/n9516 ) );
  nor_x1_sg U73174 ( .A(n67892), .B(n26016), .X(\filter_0/n9512 ) );
  nor_x1_sg U73175 ( .A(n67891), .B(n26016), .X(\filter_0/n9508 ) );
  nor_x1_sg U73176 ( .A(n67890), .B(n26016), .X(\filter_0/n9504 ) );
  nor_x1_sg U73177 ( .A(n67889), .B(n26016), .X(\filter_0/n9500 ) );
  nor_x1_sg U73178 ( .A(n67881), .B(n26018), .X(\filter_0/n9468 ) );
  nor_x1_sg U73179 ( .A(n67880), .B(n26018), .X(\filter_0/n9464 ) );
  nor_x1_sg U73180 ( .A(n67879), .B(n26018), .X(\filter_0/n9460 ) );
  nor_x1_sg U73181 ( .A(n67878), .B(n26018), .X(\filter_0/n9456 ) );
  nor_x1_sg U73182 ( .A(n67877), .B(n26018), .X(\filter_0/n9452 ) );
  nor_x1_sg U73183 ( .A(n67876), .B(n26018), .X(\filter_0/n9448 ) );
  nor_x1_sg U73184 ( .A(n67875), .B(n26018), .X(\filter_0/n9444 ) );
  nor_x1_sg U73185 ( .A(n67874), .B(n26018), .X(\filter_0/n9440 ) );
  nor_x1_sg U73186 ( .A(n67873), .B(n26018), .X(\filter_0/n9436 ) );
  nor_x1_sg U73187 ( .A(n67872), .B(n26018), .X(\filter_0/n9432 ) );
  nor_x1_sg U73188 ( .A(n67871), .B(n26018), .X(\filter_0/n9428 ) );
  nor_x1_sg U73189 ( .A(n67870), .B(n26018), .X(\filter_0/n9424 ) );
  nor_x1_sg U73190 ( .A(n67869), .B(n26018), .X(\filter_0/n9420 ) );
  nor_x1_sg U73191 ( .A(n67861), .B(n26020), .X(\filter_0/n9388 ) );
  nor_x1_sg U73192 ( .A(n67860), .B(n26020), .X(\filter_0/n9384 ) );
  nor_x1_sg U73193 ( .A(n67859), .B(n26020), .X(\filter_0/n9380 ) );
  nor_x1_sg U73194 ( .A(n67858), .B(n26020), .X(\filter_0/n9376 ) );
  nor_x1_sg U73195 ( .A(n67857), .B(n26020), .X(\filter_0/n9372 ) );
  nor_x1_sg U73196 ( .A(n67856), .B(n26020), .X(\filter_0/n9368 ) );
  nor_x1_sg U73197 ( .A(n67855), .B(n26020), .X(\filter_0/n9364 ) );
  nor_x1_sg U73198 ( .A(n67854), .B(n26020), .X(\filter_0/n9360 ) );
  nor_x1_sg U73199 ( .A(n67853), .B(n26020), .X(\filter_0/n9356 ) );
  nor_x1_sg U73200 ( .A(n67852), .B(n26020), .X(\filter_0/n9352 ) );
  nor_x1_sg U73201 ( .A(n67851), .B(n26020), .X(\filter_0/n9348 ) );
  nor_x1_sg U73202 ( .A(n67850), .B(n26020), .X(\filter_0/n9344 ) );
  nor_x1_sg U73203 ( .A(n67849), .B(n26020), .X(\filter_0/n9340 ) );
  nor_x1_sg U73204 ( .A(n67841), .B(n26022), .X(\filter_0/n9308 ) );
  nor_x1_sg U73205 ( .A(n67840), .B(n26022), .X(\filter_0/n9304 ) );
  nor_x1_sg U73206 ( .A(n67839), .B(n26022), .X(\filter_0/n9300 ) );
  nor_x1_sg U73207 ( .A(n67838), .B(n26022), .X(\filter_0/n9296 ) );
  nor_x1_sg U73208 ( .A(n67837), .B(n26022), .X(\filter_0/n9292 ) );
  nor_x1_sg U73209 ( .A(n67836), .B(n26022), .X(\filter_0/n9288 ) );
  nor_x1_sg U73210 ( .A(n67835), .B(n26022), .X(\filter_0/n9284 ) );
  nor_x1_sg U73211 ( .A(n67834), .B(n26022), .X(\filter_0/n9280 ) );
  nor_x1_sg U73212 ( .A(n67833), .B(n26022), .X(\filter_0/n9276 ) );
  nor_x1_sg U73213 ( .A(n67832), .B(n26022), .X(\filter_0/n9272 ) );
  nor_x1_sg U73214 ( .A(n67831), .B(n26022), .X(\filter_0/n9268 ) );
  nor_x1_sg U73215 ( .A(n67830), .B(n26022), .X(\filter_0/n9264 ) );
  nor_x1_sg U73216 ( .A(n67829), .B(n26022), .X(\filter_0/n9260 ) );
  nor_x1_sg U73217 ( .A(n67741), .B(n26028), .X(\filter_0/n8908 ) );
  nor_x1_sg U73218 ( .A(n67740), .B(n26028), .X(\filter_0/n8904 ) );
  nor_x1_sg U73219 ( .A(n67739), .B(n26028), .X(\filter_0/n8900 ) );
  nor_x1_sg U73220 ( .A(n67738), .B(n26028), .X(\filter_0/n8896 ) );
  nor_x1_sg U73221 ( .A(n67737), .B(n26028), .X(\filter_0/n8892 ) );
  nor_x1_sg U73222 ( .A(n67736), .B(n26028), .X(\filter_0/n8888 ) );
  nor_x1_sg U73223 ( .A(n67735), .B(n26028), .X(\filter_0/n8884 ) );
  nor_x1_sg U73224 ( .A(n67734), .B(n26028), .X(\filter_0/n8880 ) );
  nor_x1_sg U73225 ( .A(n67733), .B(n26028), .X(\filter_0/n8876 ) );
  nor_x1_sg U73226 ( .A(n67732), .B(n26028), .X(\filter_0/n8872 ) );
  nor_x1_sg U73227 ( .A(n67731), .B(n26028), .X(\filter_0/n8868 ) );
  nor_x1_sg U73228 ( .A(n67730), .B(n26028), .X(\filter_0/n8864 ) );
  nor_x1_sg U73229 ( .A(n67729), .B(n26028), .X(\filter_0/n8860 ) );
  nor_x1_sg U73230 ( .A(n67721), .B(n26029), .X(\filter_0/n8828 ) );
  nor_x1_sg U73231 ( .A(n67720), .B(n26029), .X(\filter_0/n8824 ) );
  nor_x1_sg U73232 ( .A(n67719), .B(n26029), .X(\filter_0/n8820 ) );
  nor_x1_sg U73233 ( .A(n67718), .B(n26029), .X(\filter_0/n8816 ) );
  nor_x1_sg U73234 ( .A(n67717), .B(n26029), .X(\filter_0/n8812 ) );
  nor_x1_sg U73235 ( .A(n67716), .B(n26029), .X(\filter_0/n8808 ) );
  nor_x1_sg U73236 ( .A(n67715), .B(n26029), .X(\filter_0/n8804 ) );
  nor_x1_sg U73237 ( .A(n67714), .B(n26029), .X(\filter_0/n8800 ) );
  nor_x1_sg U73238 ( .A(n67713), .B(n26029), .X(\filter_0/n8796 ) );
  nor_x1_sg U73239 ( .A(n67712), .B(n26029), .X(\filter_0/n8792 ) );
  nor_x1_sg U73240 ( .A(n67711), .B(n26029), .X(\filter_0/n8788 ) );
  nor_x1_sg U73241 ( .A(n67710), .B(n26029), .X(\filter_0/n8784 ) );
  nor_x1_sg U73242 ( .A(n67709), .B(n26029), .X(\filter_0/n8780 ) );
  nor_x1_sg U73243 ( .A(n67701), .B(n26030), .X(\filter_0/n8748 ) );
  nor_x1_sg U73244 ( .A(n67700), .B(n26030), .X(\filter_0/n8744 ) );
  nor_x1_sg U73245 ( .A(n67699), .B(n26030), .X(\filter_0/n8740 ) );
  nor_x1_sg U73246 ( .A(n67698), .B(n26030), .X(\filter_0/n8736 ) );
  nor_x1_sg U73247 ( .A(n67697), .B(n26030), .X(\filter_0/n8732 ) );
  nor_x1_sg U73248 ( .A(n67696), .B(n26030), .X(\filter_0/n8728 ) );
  nor_x1_sg U73249 ( .A(n67695), .B(n26030), .X(\filter_0/n8724 ) );
  nor_x1_sg U73250 ( .A(n67694), .B(n26030), .X(\filter_0/n8720 ) );
  nor_x1_sg U73251 ( .A(n67693), .B(n26030), .X(\filter_0/n8716 ) );
  nor_x1_sg U73252 ( .A(n67692), .B(n26030), .X(\filter_0/n8712 ) );
  nor_x1_sg U73253 ( .A(n67691), .B(n26030), .X(\filter_0/n8708 ) );
  nor_x1_sg U73254 ( .A(n67690), .B(n26030), .X(\filter_0/n8704 ) );
  nor_x1_sg U73255 ( .A(n67689), .B(n26030), .X(\filter_0/n8700 ) );
  nor_x1_sg U73256 ( .A(n67681), .B(n26031), .X(\filter_0/n8668 ) );
  nor_x1_sg U73257 ( .A(n67680), .B(n26031), .X(\filter_0/n8664 ) );
  nor_x1_sg U73258 ( .A(n67679), .B(n26031), .X(\filter_0/n8660 ) );
  nor_x1_sg U73259 ( .A(n67678), .B(n26031), .X(\filter_0/n8656 ) );
  nor_x1_sg U73260 ( .A(n67677), .B(n26031), .X(\filter_0/n8652 ) );
  nor_x1_sg U73261 ( .A(n67676), .B(n26031), .X(\filter_0/n8648 ) );
  nor_x1_sg U73262 ( .A(n67675), .B(n26031), .X(\filter_0/n8644 ) );
  nor_x1_sg U73263 ( .A(n67674), .B(n26031), .X(\filter_0/n8640 ) );
  nor_x1_sg U73264 ( .A(n67673), .B(n26031), .X(\filter_0/n8636 ) );
  nor_x1_sg U73265 ( .A(n67672), .B(n26031), .X(\filter_0/n8632 ) );
  nor_x1_sg U73266 ( .A(n67671), .B(n26031), .X(\filter_0/n8628 ) );
  nor_x1_sg U73267 ( .A(n67670), .B(n26031), .X(\filter_0/n8624 ) );
  nor_x1_sg U73268 ( .A(n67669), .B(n26031), .X(\filter_0/n8620 ) );
  nand_x2_sg U73269 ( .A(n58471), .B(n58470), .X(n24841) );
  nand_x1_sg U73270 ( .A(n56697), .B(n57329), .X(n58471) );
  nand_x1_sg U73271 ( .A(n47773), .B(n57325), .X(n58470) );
  nand_x2_sg U73272 ( .A(n58465), .B(n58464), .X(n24931) );
  nand_x1_sg U73273 ( .A(n56739), .B(n57329), .X(n58465) );
  nand_x1_sg U73274 ( .A(n51545), .B(n57325), .X(n58464) );
  nand_x2_sg U73275 ( .A(n58459), .B(n58458), .X(n25021) );
  nand_x1_sg U73276 ( .A(n51235), .B(n57329), .X(n58459) );
  nand_x1_sg U73277 ( .A(n57071), .B(n57325), .X(n58458) );
  nand_x2_sg U73278 ( .A(n58453), .B(n58452), .X(n25111) );
  nand_x1_sg U73279 ( .A(n47665), .B(n57329), .X(n58453) );
  nand_x1_sg U73280 ( .A(n57079), .B(n57325), .X(n58452) );
  nand_x2_sg U73281 ( .A(n58447), .B(n58446), .X(n25201) );
  nand_x1_sg U73282 ( .A(n56823), .B(n57329), .X(n58447) );
  nand_x1_sg U73283 ( .A(n51553), .B(n57325), .X(n58446) );
  nand_x2_sg U73284 ( .A(n58445), .B(n58444), .X(n25231) );
  nand_x1_sg U73285 ( .A(n47667), .B(n57329), .X(n58445) );
  nand_x1_sg U73286 ( .A(n57087), .B(n57325), .X(n58444) );
  nand_x2_sg U73287 ( .A(n58443), .B(n58442), .X(n25261) );
  nand_x1_sg U73288 ( .A(n51319), .B(n57329), .X(n58443) );
  nand_x1_sg U73289 ( .A(n57089), .B(n57325), .X(n58442) );
  nand_x2_sg U73290 ( .A(n58437), .B(n58436), .X(n25351) );
  nand_x1_sg U73291 ( .A(n56859), .B(n57329), .X(n58437) );
  nand_x1_sg U73292 ( .A(n51549), .B(n57325), .X(n58436) );
  nand_x2_sg U73293 ( .A(n58435), .B(n58434), .X(n25382) );
  nand_x1_sg U73294 ( .A(n51329), .B(n57329), .X(n58435) );
  nand_x1_sg U73295 ( .A(n57081), .B(n57325), .X(n58434) );
  nand_x2_sg U73296 ( .A(n58429), .B(n58428), .X(n25443) );
  nand_x1_sg U73297 ( .A(n47659), .B(n57329), .X(n58429) );
  nand_x1_sg U73298 ( .A(n57073), .B(n57325), .X(n58428) );
  nand_x2_sg U73299 ( .A(n58423), .B(n58422), .X(n25533) );
  nand_x1_sg U73300 ( .A(n56809), .B(n57329), .X(n58423) );
  nand_x1_sg U73301 ( .A(n51547), .B(n57325), .X(n58422) );
  nand_x2_sg U73302 ( .A(n58417), .B(n58416), .X(n25623) );
  nand_x1_sg U73303 ( .A(n51301), .B(n57329), .X(n58417) );
  nand_x1_sg U73304 ( .A(n57075), .B(n57325), .X(n58416) );
  nand_x2_sg U73305 ( .A(n58411), .B(n58410), .X(n25713) );
  nand_x1_sg U73306 ( .A(n47663), .B(n57329), .X(n58411) );
  nand_x1_sg U73307 ( .A(n57077), .B(n57325), .X(n58410) );
  nand_x2_sg U73308 ( .A(n58405), .B(n58404), .X(n25803) );
  nand_x1_sg U73309 ( .A(n56719), .B(n57329), .X(n58405) );
  nand_x1_sg U73310 ( .A(n51551), .B(n57325), .X(n58404) );
  nand_x2_sg U73311 ( .A(n58403), .B(n58402), .X(n25833) );
  nand_x1_sg U73312 ( .A(n47629), .B(n57329), .X(n58403) );
  nand_x1_sg U73313 ( .A(n57083), .B(n57325), .X(n58402) );
  nand_x2_sg U73314 ( .A(n58401), .B(n58400), .X(n25863) );
  nand_x1_sg U73315 ( .A(n51213), .B(n57329), .X(n58401) );
  nand_x1_sg U73316 ( .A(n57085), .B(n57325), .X(n58400) );
  nand_x2_sg U73317 ( .A(n58395), .B(n58394), .X(n25953) );
  nand_x1_sg U73318 ( .A(n56835), .B(n57329), .X(n58395) );
  nand_x1_sg U73319 ( .A(n47759), .B(n57325), .X(n58394) );
  nand_x2_sg U73320 ( .A(n58393), .B(n58392), .X(n25984) );
  nand_x1_sg U73321 ( .A(n56673), .B(n57329), .X(n58393) );
  nand_x1_sg U73322 ( .A(n51543), .B(n57325), .X(n58392) );
  nor_x1_sg U73323 ( .A(n67981), .B(n26009), .X(\filter_0/n9868 ) );
  nor_x1_sg U73324 ( .A(n67980), .B(n26009), .X(\filter_0/n9864 ) );
  nor_x1_sg U73325 ( .A(n67979), .B(n26009), .X(\filter_0/n9860 ) );
  nor_x1_sg U73326 ( .A(n67978), .B(n26009), .X(\filter_0/n9856 ) );
  nor_x1_sg U73327 ( .A(n67977), .B(n26009), .X(\filter_0/n9852 ) );
  nor_x1_sg U73328 ( .A(n67976), .B(n26009), .X(\filter_0/n9848 ) );
  nor_x1_sg U73329 ( .A(n67975), .B(n26009), .X(\filter_0/n9844 ) );
  nor_x1_sg U73330 ( .A(n67974), .B(n26009), .X(\filter_0/n9840 ) );
  nor_x1_sg U73331 ( .A(n67973), .B(n26009), .X(\filter_0/n9836 ) );
  nor_x1_sg U73332 ( .A(n67972), .B(n26009), .X(\filter_0/n9832 ) );
  nor_x1_sg U73333 ( .A(n67971), .B(n26009), .X(\filter_0/n9828 ) );
  nor_x1_sg U73334 ( .A(n67970), .B(n26009), .X(\filter_0/n9824 ) );
  nor_x1_sg U73335 ( .A(n67969), .B(n26009), .X(\filter_0/n9820 ) );
  nor_x1_sg U73336 ( .A(n67961), .B(n26011), .X(\filter_0/n9788 ) );
  nor_x1_sg U73337 ( .A(n67960), .B(n26011), .X(\filter_0/n9784 ) );
  nor_x1_sg U73338 ( .A(n67959), .B(n26011), .X(\filter_0/n9780 ) );
  nor_x1_sg U73339 ( .A(n67958), .B(n26011), .X(\filter_0/n9776 ) );
  nor_x1_sg U73340 ( .A(n67957), .B(n26011), .X(\filter_0/n9772 ) );
  nor_x1_sg U73341 ( .A(n67956), .B(n26011), .X(\filter_0/n9768 ) );
  nor_x1_sg U73342 ( .A(n67955), .B(n26011), .X(\filter_0/n9764 ) );
  nor_x1_sg U73343 ( .A(n67954), .B(n26011), .X(\filter_0/n9760 ) );
  nor_x1_sg U73344 ( .A(n67953), .B(n26011), .X(\filter_0/n9756 ) );
  nor_x1_sg U73345 ( .A(n67952), .B(n26011), .X(\filter_0/n9752 ) );
  nor_x1_sg U73346 ( .A(n67951), .B(n26011), .X(\filter_0/n9748 ) );
  nor_x1_sg U73347 ( .A(n67950), .B(n26011), .X(\filter_0/n9744 ) );
  nor_x1_sg U73348 ( .A(n67949), .B(n26011), .X(\filter_0/n9740 ) );
  nor_x1_sg U73349 ( .A(n67941), .B(n26013), .X(\filter_0/n9708 ) );
  nor_x1_sg U73350 ( .A(n67940), .B(n26013), .X(\filter_0/n9704 ) );
  nor_x1_sg U73351 ( .A(n67939), .B(n26013), .X(\filter_0/n9700 ) );
  nor_x1_sg U73352 ( .A(n67938), .B(n26013), .X(\filter_0/n9696 ) );
  nor_x1_sg U73353 ( .A(n67937), .B(n26013), .X(\filter_0/n9692 ) );
  nor_x1_sg U73354 ( .A(n67936), .B(n26013), .X(\filter_0/n9688 ) );
  nor_x1_sg U73355 ( .A(n67935), .B(n26013), .X(\filter_0/n9684 ) );
  nor_x1_sg U73356 ( .A(n67934), .B(n26013), .X(\filter_0/n9680 ) );
  nor_x1_sg U73357 ( .A(n67933), .B(n26013), .X(\filter_0/n9676 ) );
  nor_x1_sg U73358 ( .A(n67932), .B(n26013), .X(\filter_0/n9672 ) );
  nor_x1_sg U73359 ( .A(n67931), .B(n26013), .X(\filter_0/n9668 ) );
  nor_x1_sg U73360 ( .A(n67930), .B(n26013), .X(\filter_0/n9664 ) );
  nor_x1_sg U73361 ( .A(n67929), .B(n26013), .X(\filter_0/n9660 ) );
  nor_x1_sg U73362 ( .A(n67921), .B(n26015), .X(\filter_0/n9628 ) );
  nor_x1_sg U73363 ( .A(n67920), .B(n26015), .X(\filter_0/n9624 ) );
  nor_x1_sg U73364 ( .A(n67919), .B(n26015), .X(\filter_0/n9620 ) );
  nor_x1_sg U73365 ( .A(n67918), .B(n26015), .X(\filter_0/n9616 ) );
  nor_x1_sg U73366 ( .A(n67917), .B(n26015), .X(\filter_0/n9612 ) );
  nor_x1_sg U73367 ( .A(n67916), .B(n26015), .X(\filter_0/n9608 ) );
  nor_x1_sg U73368 ( .A(n67915), .B(n26015), .X(\filter_0/n9604 ) );
  nor_x1_sg U73369 ( .A(n67914), .B(n26015), .X(\filter_0/n9600 ) );
  nor_x1_sg U73370 ( .A(n67913), .B(n26015), .X(\filter_0/n9596 ) );
  nor_x1_sg U73371 ( .A(n67912), .B(n26015), .X(\filter_0/n9592 ) );
  nor_x1_sg U73372 ( .A(n67911), .B(n26015), .X(\filter_0/n9588 ) );
  nor_x1_sg U73373 ( .A(n67910), .B(n26015), .X(\filter_0/n9584 ) );
  nor_x1_sg U73374 ( .A(n67909), .B(n26015), .X(\filter_0/n9580 ) );
  nor_x1_sg U73375 ( .A(n67661), .B(n26032), .X(\filter_0/n8588 ) );
  nor_x1_sg U73376 ( .A(n67660), .B(n26032), .X(\filter_0/n8584 ) );
  nor_x1_sg U73377 ( .A(n67659), .B(n26032), .X(\filter_0/n8580 ) );
  nor_x1_sg U73378 ( .A(n67658), .B(n26032), .X(\filter_0/n8576 ) );
  nor_x1_sg U73379 ( .A(n67657), .B(n26032), .X(\filter_0/n8572 ) );
  nor_x1_sg U73380 ( .A(n67656), .B(n26032), .X(\filter_0/n8568 ) );
  nor_x1_sg U73381 ( .A(n67655), .B(n26032), .X(\filter_0/n8564 ) );
  nor_x1_sg U73382 ( .A(n67654), .B(n26032), .X(\filter_0/n8560 ) );
  nor_x1_sg U73383 ( .A(n67653), .B(n26032), .X(\filter_0/n8556 ) );
  nor_x1_sg U73384 ( .A(n67652), .B(n26032), .X(\filter_0/n8552 ) );
  nor_x1_sg U73385 ( .A(n67651), .B(n26032), .X(\filter_0/n8548 ) );
  nor_x1_sg U73386 ( .A(n67650), .B(n26032), .X(\filter_0/n8544 ) );
  nor_x1_sg U73387 ( .A(n67649), .B(n26032), .X(\filter_0/n8540 ) );
  nor_x1_sg U73388 ( .A(n67641), .B(n26035), .X(\filter_0/n8508 ) );
  nor_x1_sg U73389 ( .A(n67640), .B(n26035), .X(\filter_0/n8504 ) );
  nor_x1_sg U73390 ( .A(n67639), .B(n26035), .X(\filter_0/n8500 ) );
  nor_x1_sg U73391 ( .A(n67638), .B(n26035), .X(\filter_0/n8496 ) );
  nor_x1_sg U73392 ( .A(n67637), .B(n26035), .X(\filter_0/n8492 ) );
  nor_x1_sg U73393 ( .A(n67636), .B(n26035), .X(\filter_0/n8488 ) );
  nor_x1_sg U73394 ( .A(n67635), .B(n26035), .X(\filter_0/n8484 ) );
  nor_x1_sg U73395 ( .A(n67634), .B(n26035), .X(\filter_0/n8480 ) );
  nor_x1_sg U73396 ( .A(n67633), .B(n26035), .X(\filter_0/n8476 ) );
  nor_x1_sg U73397 ( .A(n67632), .B(n26035), .X(\filter_0/n8472 ) );
  nor_x1_sg U73398 ( .A(n67631), .B(n26035), .X(\filter_0/n8468 ) );
  nor_x1_sg U73399 ( .A(n67630), .B(n26035), .X(\filter_0/n8464 ) );
  nor_x1_sg U73400 ( .A(n67629), .B(n26035), .X(\filter_0/n8460 ) );
  nor_x1_sg U73401 ( .A(n67621), .B(n26037), .X(\filter_0/n8428 ) );
  nor_x1_sg U73402 ( .A(n67620), .B(n26037), .X(\filter_0/n8424 ) );
  nor_x1_sg U73403 ( .A(n67619), .B(n26037), .X(\filter_0/n8420 ) );
  nor_x1_sg U73404 ( .A(n67618), .B(n26037), .X(\filter_0/n8416 ) );
  nor_x1_sg U73405 ( .A(n67617), .B(n26037), .X(\filter_0/n8412 ) );
  nor_x1_sg U73406 ( .A(n67616), .B(n26037), .X(\filter_0/n8408 ) );
  nor_x1_sg U73407 ( .A(n67615), .B(n26037), .X(\filter_0/n8404 ) );
  nor_x1_sg U73408 ( .A(n67614), .B(n26037), .X(\filter_0/n8400 ) );
  nor_x1_sg U73409 ( .A(n67613), .B(n26037), .X(\filter_0/n8396 ) );
  nor_x1_sg U73410 ( .A(n67612), .B(n26037), .X(\filter_0/n8392 ) );
  nor_x1_sg U73411 ( .A(n67611), .B(n26037), .X(\filter_0/n8388 ) );
  nor_x1_sg U73412 ( .A(n67610), .B(n26037), .X(\filter_0/n8384 ) );
  nor_x1_sg U73413 ( .A(n67609), .B(n26037), .X(\filter_0/n8380 ) );
  nor_x1_sg U73414 ( .A(n67601), .B(n26038), .X(\filter_0/n8348 ) );
  nor_x1_sg U73415 ( .A(n67600), .B(n26038), .X(\filter_0/n8344 ) );
  nor_x1_sg U73416 ( .A(n67599), .B(n26038), .X(\filter_0/n8340 ) );
  nor_x1_sg U73417 ( .A(n67598), .B(n26038), .X(\filter_0/n8336 ) );
  nor_x1_sg U73418 ( .A(n67597), .B(n26038), .X(\filter_0/n8332 ) );
  nor_x1_sg U73419 ( .A(n67596), .B(n26038), .X(\filter_0/n8328 ) );
  nor_x1_sg U73420 ( .A(n67595), .B(n26038), .X(\filter_0/n8324 ) );
  nor_x1_sg U73421 ( .A(n67594), .B(n26038), .X(\filter_0/n8320 ) );
  nor_x1_sg U73422 ( .A(n67593), .B(n26038), .X(\filter_0/n8316 ) );
  nor_x1_sg U73423 ( .A(n67592), .B(n26038), .X(\filter_0/n8312 ) );
  nor_x1_sg U73424 ( .A(n67591), .B(n26038), .X(\filter_0/n8308 ) );
  nor_x1_sg U73425 ( .A(n67590), .B(n26038), .X(\filter_0/n8304 ) );
  nor_x1_sg U73426 ( .A(n67589), .B(n26038), .X(\filter_0/n8300 ) );
  nand_x1_sg U73427 ( .A(n47743), .B(n22749), .X(n22748) );
  nand_x1_sg U73428 ( .A(n47745), .B(n57154), .X(n22763) );
  nand_x1_sg U73429 ( .A(n51489), .B(n22749), .X(n22774) );
  nand_x1_sg U73430 ( .A(n51493), .B(n57154), .X(n22785) );
  nand_x1_sg U73431 ( .A(n57015), .B(n22749), .X(n22796) );
  nand_x1_sg U73432 ( .A(n47747), .B(n57154), .X(n22807) );
  nand_x1_sg U73433 ( .A(n51491), .B(n22749), .X(n22818) );
  nand_x1_sg U73434 ( .A(n57013), .B(n57154), .X(n22829) );
  nand_x1_sg U73435 ( .A(n51515), .B(n22749), .X(n22840) );
  nand_x1_sg U73436 ( .A(n57039), .B(n57154), .X(n22851) );
  nand_x1_sg U73437 ( .A(n51503), .B(n22749), .X(n22862) );
  nand_x1_sg U73438 ( .A(n57021), .B(n57154), .X(n22873) );
  nand_x1_sg U73439 ( .A(n51517), .B(n22749), .X(n22884) );
  nand_x1_sg U73440 ( .A(n57041), .B(n57154), .X(n22895) );
  nand_x1_sg U73441 ( .A(n47757), .B(n22749), .X(n22906) );
  nand_x1_sg U73442 ( .A(n51505), .B(n57154), .X(n22917) );
  nand_x1_sg U73443 ( .A(n57027), .B(n22749), .X(n22928) );
  nand_x1_sg U73444 ( .A(n51519), .B(n57154), .X(n22939) );
  nand_x1_sg U73445 ( .A(n57043), .B(n22749), .X(n22950) );
  nand_x1_sg U73446 ( .A(n57029), .B(n57154), .X(n22961) );
  nand_x1_sg U73447 ( .A(n47749), .B(n22977), .X(n22976) );
  nand_x1_sg U73448 ( .A(n47751), .B(n57148), .X(n22990) );
  nand_x1_sg U73449 ( .A(n51495), .B(n22977), .X(n23001) );
  nand_x1_sg U73450 ( .A(n51507), .B(n57148), .X(n23012) );
  nand_x1_sg U73451 ( .A(n57031), .B(n22977), .X(n23023) );
  nand_x1_sg U73452 ( .A(n47753), .B(n57148), .X(n23034) );
  nand_x1_sg U73453 ( .A(n51497), .B(n22977), .X(n23045) );
  nand_x1_sg U73454 ( .A(n57017), .B(n57148), .X(n23056) );
  nand_x1_sg U73455 ( .A(n51509), .B(n22977), .X(n23067) );
  nand_x1_sg U73456 ( .A(n57033), .B(n57148), .X(n23078) );
  nand_x1_sg U73457 ( .A(n51499), .B(n22977), .X(n23089) );
  nand_x1_sg U73458 ( .A(n57019), .B(n57148), .X(n23100) );
  nand_x1_sg U73459 ( .A(n51511), .B(n22977), .X(n23111) );
  nand_x1_sg U73460 ( .A(n57035), .B(n57148), .X(n23122) );
  nand_x1_sg U73461 ( .A(n47755), .B(n22977), .X(n23133) );
  nand_x1_sg U73462 ( .A(n51501), .B(n57148), .X(n23144) );
  nand_x1_sg U73463 ( .A(n57023), .B(n22977), .X(n23155) );
  nand_x1_sg U73464 ( .A(n51513), .B(n57148), .X(n23166) );
  nand_x1_sg U73465 ( .A(n57037), .B(n22977), .X(n23177) );
  nand_x1_sg U73466 ( .A(n57025), .B(n57148), .X(n23188) );
  nand_x2_sg U73467 ( .A(n26148), .B(n26149), .X(n26144) );
  nand_x2_sg U73468 ( .A(n26146), .B(n26147), .X(n26145) );
  nand_x1_sg U73469 ( .A(n57107), .B(n53641), .X(n26148) );
  nand_x2_sg U73470 ( .A(n26109), .B(n26110), .X(n26105) );
  nand_x2_sg U73471 ( .A(n26107), .B(n26108), .X(n26106) );
  nand_x1_sg U73472 ( .A(n57107), .B(n53643), .X(n26109) );
  nand_x2_sg U73473 ( .A(n26240), .B(n26241), .X(n26236) );
  nand_x2_sg U73474 ( .A(n26238), .B(n26239), .X(n26237) );
  nand_x1_sg U73475 ( .A(n57107), .B(n53645), .X(n26240) );
  nand_x2_sg U73476 ( .A(n26206), .B(n26207), .X(n26202) );
  nand_x2_sg U73477 ( .A(n26204), .B(n26205), .X(n26203) );
  nand_x1_sg U73478 ( .A(n57107), .B(n53647), .X(n26206) );
  nor_x1_sg U73479 ( .A(n68146), .B(n26253), .X(\filter_0/n10528 ) );
  nor_x1_sg U73480 ( .A(n68145), .B(n26253), .X(\filter_0/n10524 ) );
  nor_x1_sg U73481 ( .A(n68144), .B(n26253), .X(\filter_0/n10520 ) );
  nor_x1_sg U73482 ( .A(n68143), .B(n26253), .X(\filter_0/n10516 ) );
  nor_x1_sg U73483 ( .A(n68142), .B(n26253), .X(\filter_0/n10512 ) );
  nor_x1_sg U73484 ( .A(n68126), .B(n26254), .X(\filter_0/n10448 ) );
  nor_x1_sg U73485 ( .A(n68125), .B(n26254), .X(\filter_0/n10444 ) );
  nor_x1_sg U73486 ( .A(n68124), .B(n26254), .X(\filter_0/n10440 ) );
  nor_x1_sg U73487 ( .A(n68123), .B(n26254), .X(\filter_0/n10436 ) );
  nor_x1_sg U73488 ( .A(n68122), .B(n26254), .X(\filter_0/n10432 ) );
  nor_x1_sg U73489 ( .A(n68106), .B(n26255), .X(\filter_0/n10368 ) );
  nor_x1_sg U73490 ( .A(n68105), .B(n26255), .X(\filter_0/n10364 ) );
  nor_x1_sg U73491 ( .A(n68104), .B(n26255), .X(\filter_0/n10360 ) );
  nor_x1_sg U73492 ( .A(n68103), .B(n26255), .X(\filter_0/n10356 ) );
  nor_x1_sg U73493 ( .A(n68102), .B(n26255), .X(\filter_0/n10352 ) );
  nor_x1_sg U73494 ( .A(n68086), .B(n26256), .X(\filter_0/n10288 ) );
  nor_x1_sg U73495 ( .A(n68085), .B(n26256), .X(\filter_0/n10284 ) );
  nor_x1_sg U73496 ( .A(n68084), .B(n26256), .X(\filter_0/n10280 ) );
  nor_x1_sg U73497 ( .A(n68083), .B(n26256), .X(\filter_0/n10276 ) );
  nor_x1_sg U73498 ( .A(n68082), .B(n26256), .X(\filter_0/n10272 ) );
  nor_x1_sg U73499 ( .A(n67826), .B(n26024), .X(\filter_0/n9248 ) );
  nor_x1_sg U73500 ( .A(n67825), .B(n26024), .X(\filter_0/n9244 ) );
  nor_x1_sg U73501 ( .A(n67824), .B(n26024), .X(\filter_0/n9240 ) );
  nor_x1_sg U73502 ( .A(n67823), .B(n26024), .X(\filter_0/n9236 ) );
  nor_x1_sg U73503 ( .A(n67822), .B(n26024), .X(\filter_0/n9232 ) );
  nor_x1_sg U73504 ( .A(n67806), .B(n26025), .X(\filter_0/n9168 ) );
  nor_x1_sg U73505 ( .A(n67805), .B(n26025), .X(\filter_0/n9164 ) );
  nor_x1_sg U73506 ( .A(n67804), .B(n26025), .X(\filter_0/n9160 ) );
  nor_x1_sg U73507 ( .A(n67803), .B(n26025), .X(\filter_0/n9156 ) );
  nor_x1_sg U73508 ( .A(n67802), .B(n26025), .X(\filter_0/n9152 ) );
  nor_x1_sg U73509 ( .A(n67786), .B(n26026), .X(\filter_0/n9088 ) );
  nor_x1_sg U73510 ( .A(n67785), .B(n26026), .X(\filter_0/n9084 ) );
  nor_x1_sg U73511 ( .A(n67784), .B(n26026), .X(\filter_0/n9080 ) );
  nor_x1_sg U73512 ( .A(n67783), .B(n26026), .X(\filter_0/n9076 ) );
  nor_x1_sg U73513 ( .A(n67782), .B(n26026), .X(\filter_0/n9072 ) );
  nor_x1_sg U73514 ( .A(n67766), .B(n26027), .X(\filter_0/n9008 ) );
  nor_x1_sg U73515 ( .A(n67765), .B(n26027), .X(\filter_0/n9004 ) );
  nor_x1_sg U73516 ( .A(n67764), .B(n26027), .X(\filter_0/n9000 ) );
  nor_x1_sg U73517 ( .A(n67763), .B(n26027), .X(\filter_0/n8996 ) );
  nor_x1_sg U73518 ( .A(n67762), .B(n26027), .X(\filter_0/n8992 ) );
  nor_x1_sg U73519 ( .A(n67093), .B(n26003), .X(\shifter_0/n10257 ) );
  nor_x1_sg U73520 ( .A(n67092), .B(n26003), .X(\shifter_0/n10245 ) );
  nor_x1_sg U73521 ( .A(n67091), .B(n26003), .X(\shifter_0/n10233 ) );
  nor_x1_sg U73522 ( .A(n67090), .B(n26003), .X(\shifter_0/n10229 ) );
  nor_x1_sg U73523 ( .A(n67089), .B(n26003), .X(\shifter_0/n10225 ) );
  nor_x1_sg U73524 ( .A(n22395), .B(n67312), .X(\shifter_0/n12737 ) );
  nor_x1_sg U73525 ( .A(n22395), .B(n67311), .X(\shifter_0/n12725 ) );
  nor_x1_sg U73526 ( .A(n22395), .B(n67310), .X(\shifter_0/n12713 ) );
  nor_x1_sg U73527 ( .A(n22395), .B(n67309), .X(\shifter_0/n12709 ) );
  nor_x1_sg U73528 ( .A(n22395), .B(n67308), .X(\shifter_0/n12705 ) );
  nor_x1_sg U73529 ( .A(n22395), .B(n67307), .X(\shifter_0/n12693 ) );
  nor_x1_sg U73530 ( .A(n68226), .B(n26249), .X(\filter_0/n8236 ) );
  nor_x1_sg U73531 ( .A(n68225), .B(n26249), .X(\filter_0/n10844 ) );
  nor_x1_sg U73532 ( .A(n68224), .B(n26249), .X(\filter_0/n10840 ) );
  nor_x1_sg U73533 ( .A(n68223), .B(n26249), .X(\filter_0/n10836 ) );
  nor_x1_sg U73534 ( .A(n68222), .B(n26249), .X(\filter_0/n10832 ) );
  nor_x1_sg U73535 ( .A(n68206), .B(n26250), .X(\filter_0/n10768 ) );
  nor_x1_sg U73536 ( .A(n68205), .B(n26250), .X(\filter_0/n10764 ) );
  nor_x1_sg U73537 ( .A(n68204), .B(n26250), .X(\filter_0/n10760 ) );
  nor_x1_sg U73538 ( .A(n68203), .B(n26250), .X(\filter_0/n10756 ) );
  nor_x1_sg U73539 ( .A(n68202), .B(n26250), .X(\filter_0/n10752 ) );
  nor_x1_sg U73540 ( .A(n68186), .B(n26251), .X(\filter_0/n10688 ) );
  nor_x1_sg U73541 ( .A(n68185), .B(n26251), .X(\filter_0/n10684 ) );
  nor_x1_sg U73542 ( .A(n68184), .B(n26251), .X(\filter_0/n10680 ) );
  nor_x1_sg U73543 ( .A(n68183), .B(n26251), .X(\filter_0/n10676 ) );
  nor_x1_sg U73544 ( .A(n68182), .B(n26251), .X(\filter_0/n10672 ) );
  nor_x1_sg U73545 ( .A(n68166), .B(n26252), .X(\filter_0/n10608 ) );
  nor_x1_sg U73546 ( .A(n68165), .B(n26252), .X(\filter_0/n10604 ) );
  nor_x1_sg U73547 ( .A(n68164), .B(n26252), .X(\filter_0/n10600 ) );
  nor_x1_sg U73548 ( .A(n68163), .B(n26252), .X(\filter_0/n10596 ) );
  nor_x1_sg U73549 ( .A(n68162), .B(n26252), .X(\filter_0/n10592 ) );
  nor_x1_sg U73550 ( .A(n68066), .B(n26257), .X(\filter_0/n10208 ) );
  nor_x1_sg U73551 ( .A(n68065), .B(n26257), .X(\filter_0/n10204 ) );
  nor_x1_sg U73552 ( .A(n68064), .B(n26257), .X(\filter_0/n10200 ) );
  nor_x1_sg U73553 ( .A(n68063), .B(n26257), .X(\filter_0/n10196 ) );
  nor_x1_sg U73554 ( .A(n68062), .B(n26257), .X(\filter_0/n10192 ) );
  nor_x1_sg U73555 ( .A(n68046), .B(n26259), .X(\filter_0/n10128 ) );
  nor_x1_sg U73556 ( .A(n68045), .B(n26259), .X(\filter_0/n10124 ) );
  nor_x1_sg U73557 ( .A(n68044), .B(n26259), .X(\filter_0/n10120 ) );
  nor_x1_sg U73558 ( .A(n68043), .B(n26259), .X(\filter_0/n10116 ) );
  nor_x1_sg U73559 ( .A(n68042), .B(n26259), .X(\filter_0/n10112 ) );
  nor_x1_sg U73560 ( .A(n68013), .B(n26006), .X(\filter_0/n9996 ) );
  nor_x1_sg U73561 ( .A(n68012), .B(n26006), .X(\filter_0/n9992 ) );
  nor_x1_sg U73562 ( .A(n68011), .B(n26006), .X(\filter_0/n9988 ) );
  nor_x1_sg U73563 ( .A(n68010), .B(n26006), .X(\filter_0/n9984 ) );
  nor_x1_sg U73564 ( .A(n68006), .B(n26007), .X(\filter_0/n9968 ) );
  nor_x1_sg U73565 ( .A(n68005), .B(n26007), .X(\filter_0/n9964 ) );
  nor_x1_sg U73566 ( .A(n68004), .B(n26007), .X(\filter_0/n9960 ) );
  nor_x1_sg U73567 ( .A(n68003), .B(n26007), .X(\filter_0/n9956 ) );
  nor_x1_sg U73568 ( .A(n68002), .B(n26007), .X(\filter_0/n9952 ) );
  nor_x1_sg U73569 ( .A(n67906), .B(n26016), .X(\filter_0/n9568 ) );
  nor_x1_sg U73570 ( .A(n67905), .B(n26016), .X(\filter_0/n9564 ) );
  nor_x1_sg U73571 ( .A(n67904), .B(n26016), .X(\filter_0/n9560 ) );
  nor_x1_sg U73572 ( .A(n67903), .B(n26016), .X(\filter_0/n9556 ) );
  nor_x1_sg U73573 ( .A(n67902), .B(n26016), .X(\filter_0/n9552 ) );
  nor_x1_sg U73574 ( .A(n67886), .B(n26018), .X(\filter_0/n9488 ) );
  nor_x1_sg U73575 ( .A(n67885), .B(n26018), .X(\filter_0/n9484 ) );
  nor_x1_sg U73576 ( .A(n67884), .B(n26018), .X(\filter_0/n9480 ) );
  nor_x1_sg U73577 ( .A(n67883), .B(n26018), .X(\filter_0/n9476 ) );
  nor_x1_sg U73578 ( .A(n67882), .B(n26018), .X(\filter_0/n9472 ) );
  nor_x1_sg U73579 ( .A(n67866), .B(n26020), .X(\filter_0/n9408 ) );
  nor_x1_sg U73580 ( .A(n67865), .B(n26020), .X(\filter_0/n9404 ) );
  nor_x1_sg U73581 ( .A(n67864), .B(n26020), .X(\filter_0/n9400 ) );
  nor_x1_sg U73582 ( .A(n67863), .B(n26020), .X(\filter_0/n9396 ) );
  nor_x1_sg U73583 ( .A(n67862), .B(n26020), .X(\filter_0/n9392 ) );
  nor_x1_sg U73584 ( .A(n67846), .B(n26022), .X(\filter_0/n9328 ) );
  nor_x1_sg U73585 ( .A(n67845), .B(n26022), .X(\filter_0/n9324 ) );
  nor_x1_sg U73586 ( .A(n67844), .B(n26022), .X(\filter_0/n9320 ) );
  nor_x1_sg U73587 ( .A(n67843), .B(n26022), .X(\filter_0/n9316 ) );
  nor_x1_sg U73588 ( .A(n67842), .B(n26022), .X(\filter_0/n9312 ) );
  nor_x1_sg U73589 ( .A(n67746), .B(n26028), .X(\filter_0/n8928 ) );
  nor_x1_sg U73590 ( .A(n67745), .B(n26028), .X(\filter_0/n8924 ) );
  nor_x1_sg U73591 ( .A(n67744), .B(n26028), .X(\filter_0/n8920 ) );
  nor_x1_sg U73592 ( .A(n67743), .B(n26028), .X(\filter_0/n8916 ) );
  nor_x1_sg U73593 ( .A(n67742), .B(n26028), .X(\filter_0/n8912 ) );
  nor_x1_sg U73594 ( .A(n67726), .B(n26029), .X(\filter_0/n8848 ) );
  nor_x1_sg U73595 ( .A(n67725), .B(n26029), .X(\filter_0/n8844 ) );
  nor_x1_sg U73596 ( .A(n67724), .B(n26029), .X(\filter_0/n8840 ) );
  nor_x1_sg U73597 ( .A(n67723), .B(n26029), .X(\filter_0/n8836 ) );
  nor_x1_sg U73598 ( .A(n67722), .B(n26029), .X(\filter_0/n8832 ) );
  nor_x1_sg U73599 ( .A(n67706), .B(n26030), .X(\filter_0/n8768 ) );
  nor_x1_sg U73600 ( .A(n67705), .B(n26030), .X(\filter_0/n8764 ) );
  nor_x1_sg U73601 ( .A(n67704), .B(n26030), .X(\filter_0/n8760 ) );
  nor_x1_sg U73602 ( .A(n67703), .B(n26030), .X(\filter_0/n8756 ) );
  nor_x1_sg U73603 ( .A(n67702), .B(n26030), .X(\filter_0/n8752 ) );
  nor_x1_sg U73604 ( .A(n67686), .B(n26031), .X(\filter_0/n8688 ) );
  nor_x1_sg U73605 ( .A(n67685), .B(n26031), .X(\filter_0/n8684 ) );
  nor_x1_sg U73606 ( .A(n67684), .B(n26031), .X(\filter_0/n8680 ) );
  nor_x1_sg U73607 ( .A(n67683), .B(n26031), .X(\filter_0/n8676 ) );
  nor_x1_sg U73608 ( .A(n67682), .B(n26031), .X(\filter_0/n8672 ) );
  nor_x1_sg U73609 ( .A(n67986), .B(n26009), .X(\filter_0/n9888 ) );
  nor_x1_sg U73610 ( .A(n67985), .B(n26009), .X(\filter_0/n9884 ) );
  nor_x1_sg U73611 ( .A(n67984), .B(n26009), .X(\filter_0/n9880 ) );
  nor_x1_sg U73612 ( .A(n67983), .B(n26009), .X(\filter_0/n9876 ) );
  nor_x1_sg U73613 ( .A(n67982), .B(n26009), .X(\filter_0/n9872 ) );
  nor_x1_sg U73614 ( .A(n67966), .B(n26011), .X(\filter_0/n9808 ) );
  nor_x1_sg U73615 ( .A(n67965), .B(n26011), .X(\filter_0/n9804 ) );
  nor_x1_sg U73616 ( .A(n67964), .B(n26011), .X(\filter_0/n9800 ) );
  nor_x1_sg U73617 ( .A(n67963), .B(n26011), .X(\filter_0/n9796 ) );
  nor_x1_sg U73618 ( .A(n67962), .B(n26011), .X(\filter_0/n9792 ) );
  nor_x1_sg U73619 ( .A(n67946), .B(n26013), .X(\filter_0/n9728 ) );
  nor_x1_sg U73620 ( .A(n67945), .B(n26013), .X(\filter_0/n9724 ) );
  nor_x1_sg U73621 ( .A(n67944), .B(n26013), .X(\filter_0/n9720 ) );
  nor_x1_sg U73622 ( .A(n67943), .B(n26013), .X(\filter_0/n9716 ) );
  nor_x1_sg U73623 ( .A(n67942), .B(n26013), .X(\filter_0/n9712 ) );
  nor_x1_sg U73624 ( .A(n67926), .B(n26015), .X(\filter_0/n9648 ) );
  nor_x1_sg U73625 ( .A(n67925), .B(n26015), .X(\filter_0/n9644 ) );
  nor_x1_sg U73626 ( .A(n67924), .B(n26015), .X(\filter_0/n9640 ) );
  nor_x1_sg U73627 ( .A(n67923), .B(n26015), .X(\filter_0/n9636 ) );
  nor_x1_sg U73628 ( .A(n67922), .B(n26015), .X(\filter_0/n9632 ) );
  nor_x1_sg U73629 ( .A(n67666), .B(n26032), .X(\filter_0/n8608 ) );
  nor_x1_sg U73630 ( .A(n67665), .B(n26032), .X(\filter_0/n8604 ) );
  nor_x1_sg U73631 ( .A(n67664), .B(n26032), .X(\filter_0/n8600 ) );
  nor_x1_sg U73632 ( .A(n67663), .B(n26032), .X(\filter_0/n8596 ) );
  nor_x1_sg U73633 ( .A(n67662), .B(n26032), .X(\filter_0/n8592 ) );
  nor_x1_sg U73634 ( .A(n67646), .B(n26035), .X(\filter_0/n8528 ) );
  nor_x1_sg U73635 ( .A(n67645), .B(n26035), .X(\filter_0/n8524 ) );
  nor_x1_sg U73636 ( .A(n67644), .B(n26035), .X(\filter_0/n8520 ) );
  nor_x1_sg U73637 ( .A(n67643), .B(n26035), .X(\filter_0/n8516 ) );
  nor_x1_sg U73638 ( .A(n67642), .B(n26035), .X(\filter_0/n8512 ) );
  nor_x1_sg U73639 ( .A(n67626), .B(n26037), .X(\filter_0/n8448 ) );
  nor_x1_sg U73640 ( .A(n67625), .B(n26037), .X(\filter_0/n8444 ) );
  nor_x1_sg U73641 ( .A(n67624), .B(n26037), .X(\filter_0/n8440 ) );
  nor_x1_sg U73642 ( .A(n67623), .B(n26037), .X(\filter_0/n8436 ) );
  nor_x1_sg U73643 ( .A(n67622), .B(n26037), .X(\filter_0/n8432 ) );
  nor_x1_sg U73644 ( .A(n67606), .B(n26038), .X(\filter_0/n8368 ) );
  nor_x1_sg U73645 ( .A(n67605), .B(n26038), .X(\filter_0/n8364 ) );
  nor_x1_sg U73646 ( .A(n67604), .B(n26038), .X(\filter_0/n8360 ) );
  nor_x1_sg U73647 ( .A(n67603), .B(n26038), .X(\filter_0/n8356 ) );
  nor_x1_sg U73648 ( .A(n67602), .B(n26038), .X(\filter_0/n8352 ) );
  nor_x1_sg U73649 ( .A(n22395), .B(n67314), .X(\shifter_0/n12761 ) );
  nor_x1_sg U73650 ( .A(n22395), .B(n67313), .X(\shifter_0/n12749 ) );
  nor_x1_sg U73651 ( .A(n58650), .B(n26003), .X(\shifter_0/n10285 ) );
  nor_x1_sg U73652 ( .A(n67095), .B(n26003), .X(\shifter_0/n10281 ) );
  nor_x1_sg U73653 ( .A(n67094), .B(n26003), .X(\shifter_0/n10269 ) );
  nor_x1_sg U73654 ( .A(n22395), .B(n67306), .X(\shifter_0/n12689 ) );
  nor_x1_sg U73655 ( .A(n67088), .B(n26003), .X(\shifter_0/n10213 ) );
  nor_x1_sg U73656 ( .A(n67087), .B(n26003), .X(\shifter_0/n10209 ) );
  nand_x2_sg U73657 ( .A(n58475), .B(n58474), .X(n24805) );
  nand_x1_sg U73658 ( .A(n47533), .B(n57329), .X(n58475) );
  nand_x1_sg U73659 ( .A(n57045), .B(n57325), .X(n58474) );
  nand_x2_sg U73660 ( .A(n58469), .B(n58468), .X(n24871) );
  nand_x1_sg U73661 ( .A(n47649), .B(n57329), .X(n58469) );
  nand_x1_sg U73662 ( .A(n56983), .B(n57325), .X(n58468) );
  nand_x2_sg U73663 ( .A(n58467), .B(n58466), .X(n24901) );
  nand_x1_sg U73664 ( .A(n51277), .B(n57329), .X(n58467) );
  nand_x1_sg U73665 ( .A(n56985), .B(n57325), .X(n58466) );
  nand_x2_sg U73666 ( .A(n58463), .B(n58462), .X(n24961) );
  nand_x1_sg U73667 ( .A(n47535), .B(n57329), .X(n58463) );
  nand_x1_sg U73668 ( .A(n56979), .B(n57325), .X(n58462) );
  nand_x2_sg U73669 ( .A(n58461), .B(n58460), .X(n24991) );
  nand_x1_sg U73670 ( .A(n47651), .B(n57329), .X(n58461) );
  nand_x1_sg U73671 ( .A(n56981), .B(n57325), .X(n58460) );
  nand_x2_sg U73672 ( .A(n58457), .B(n58456), .X(n25051) );
  nand_x1_sg U73673 ( .A(n47671), .B(n57329), .X(n58457) );
  nand_x1_sg U73674 ( .A(n57009), .B(n57325), .X(n58456) );
  nand_x2_sg U73675 ( .A(n58455), .B(n58454), .X(n25081) );
  nand_x1_sg U73676 ( .A(n51377), .B(n57329), .X(n58455) );
  nand_x1_sg U73677 ( .A(n57011), .B(n57325), .X(n58454) );
  nand_x2_sg U73678 ( .A(n58451), .B(n58450), .X(n25141) );
  nand_x1_sg U73679 ( .A(n51317), .B(n57329), .X(n58451) );
  nand_x1_sg U73680 ( .A(n57001), .B(n57325), .X(n58450) );
  nand_x2_sg U73681 ( .A(n58449), .B(n58448), .X(n25171) );
  nand_x1_sg U73682 ( .A(n51379), .B(n57329), .X(n58449) );
  nand_x1_sg U73683 ( .A(n57003), .B(n57325), .X(n58448) );
  nand_x2_sg U73684 ( .A(n58441), .B(n58440), .X(n25291) );
  nand_x1_sg U73685 ( .A(n51423), .B(n57329), .X(n58441) );
  nand_x1_sg U73686 ( .A(n56997), .B(n57325), .X(n58440) );
  nand_x2_sg U73687 ( .A(n58439), .B(n58438), .X(n25321) );
  nand_x1_sg U73688 ( .A(n47707), .B(n57329), .X(n58439) );
  nand_x1_sg U73689 ( .A(n56995), .B(n57325), .X(n58438) );
  nand_x2_sg U73690 ( .A(n58433), .B(n58432), .X(n25413) );
  nand_x1_sg U73691 ( .A(n47549), .B(n57329), .X(n58433) );
  nand_x1_sg U73692 ( .A(n57047), .B(n57325), .X(n58432) );
  nand_x2_sg U73693 ( .A(n58427), .B(n58426), .X(n25473) );
  nand_x1_sg U73694 ( .A(n51299), .B(n57329), .X(n58427) );
  nand_x1_sg U73695 ( .A(n56987), .B(n57325), .X(n58426) );
  nand_x2_sg U73696 ( .A(n58425), .B(n58424), .X(n25503) );
  nand_x1_sg U73697 ( .A(n51361), .B(n57329), .X(n58425) );
  nand_x1_sg U73698 ( .A(n56989), .B(n57325), .X(n58424) );
  nand_x2_sg U73699 ( .A(n58421), .B(n58420), .X(n25563) );
  nand_x1_sg U73700 ( .A(n47551), .B(n57329), .X(n58421) );
  nand_x1_sg U73701 ( .A(n56991), .B(n57325), .X(n58420) );
  nand_x2_sg U73702 ( .A(n58419), .B(n58418), .X(n25593) );
  nand_x1_sg U73703 ( .A(n47661), .B(n57329), .X(n58419) );
  nand_x1_sg U73704 ( .A(n56993), .B(n57325), .X(n58418) );
  nand_x2_sg U73705 ( .A(n58415), .B(n58414), .X(n25653) );
  nand_x1_sg U73706 ( .A(n47669), .B(n57329), .X(n58415) );
  nand_x1_sg U73707 ( .A(n57005), .B(n57325), .X(n58414) );
  nand_x2_sg U73708 ( .A(n58413), .B(n58412), .X(n25683) );
  nand_x1_sg U73709 ( .A(n51363), .B(n57329), .X(n58413) );
  nand_x1_sg U73710 ( .A(n57007), .B(n57325), .X(n58412) );
  nand_x2_sg U73711 ( .A(n58409), .B(n58408), .X(n25743) );
  nand_x1_sg U73712 ( .A(n51303), .B(n57329), .X(n58409) );
  nand_x1_sg U73713 ( .A(n56999), .B(n57325), .X(n58408) );
  nand_x2_sg U73714 ( .A(n58407), .B(n58406), .X(n25773) );
  nand_x1_sg U73715 ( .A(n51257), .B(n57329), .X(n58407) );
  nand_x1_sg U73716 ( .A(n56977), .B(n57325), .X(n58406) );
  nand_x2_sg U73717 ( .A(n58399), .B(n58398), .X(n25893) );
  nand_x1_sg U73718 ( .A(n47683), .B(n57329), .X(n58399) );
  nand_x1_sg U73719 ( .A(n56973), .B(n57325), .X(n58398) );
  nand_x2_sg U73720 ( .A(n58397), .B(n58396), .X(n25923) );
  nand_x1_sg U73721 ( .A(n51393), .B(n57329), .X(n58397) );
  nand_x1_sg U73722 ( .A(n56975), .B(n57325), .X(n58396) );
  nand_x2_sg U73723 ( .A(n24798), .B(n24799), .X(n24797) );
  nand_x1_sg U73724 ( .A(n47631), .B(n57322), .X(n24798) );
  nand_x1_sg U73725 ( .A(n57498), .B(n47475), .X(n24799) );
  nand_x2_sg U73726 ( .A(n24837), .B(n24838), .X(n24836) );
  nand_x1_sg U73727 ( .A(n47633), .B(n57322), .X(n24837) );
  nand_x1_sg U73728 ( .A(n57496), .B(n47389), .X(n24838) );
  nand_x2_sg U73729 ( .A(n24867), .B(n24868), .X(n24866) );
  nand_x1_sg U73730 ( .A(n51219), .B(n57322), .X(n24867) );
  nand_x1_sg U73731 ( .A(n57496), .B(n47447), .X(n24868) );
  nand_x2_sg U73732 ( .A(n24897), .B(n24898), .X(n24896) );
  nand_x1_sg U73733 ( .A(n51263), .B(n57322), .X(n24897) );
  nand_x1_sg U73734 ( .A(n57496), .B(n47477), .X(n24898) );
  nand_x2_sg U73735 ( .A(n24927), .B(n24928), .X(n24926) );
  nand_x1_sg U73736 ( .A(n56725), .B(n57322), .X(n24927) );
  nand_x1_sg U73737 ( .A(n57496), .B(n47387), .X(n24928) );
  nand_x2_sg U73738 ( .A(n24957), .B(n24958), .X(n24956) );
  nand_x1_sg U73739 ( .A(n47635), .B(n57322), .X(n24957) );
  nand_x1_sg U73740 ( .A(n57496), .B(n47304), .X(n24958) );
  nand_x2_sg U73741 ( .A(n24987), .B(n24988), .X(n24986) );
  nand_x1_sg U73742 ( .A(n51221), .B(n57322), .X(n24987) );
  nand_x1_sg U73743 ( .A(n57496), .B(n47483), .X(n24988) );
  nand_x2_sg U73744 ( .A(n25017), .B(n25018), .X(n25016) );
  nand_x1_sg U73745 ( .A(n56683), .B(n57322), .X(n25017) );
  nand_x1_sg U73746 ( .A(n57496), .B(n47455), .X(n25018) );
  nand_x2_sg U73747 ( .A(n25047), .B(n25048), .X(n25046) );
  nand_x1_sg U73748 ( .A(n51373), .B(n57322), .X(n25047) );
  nand_x1_sg U73749 ( .A(n57496), .B(n47487), .X(n25048) );
  nand_x2_sg U73750 ( .A(n25077), .B(n25078), .X(n25076) );
  nand_x1_sg U73751 ( .A(n56819), .B(n57322), .X(n25077) );
  nand_x1_sg U73752 ( .A(n57496), .B(n47467), .X(n25078) );
  nand_x2_sg U73753 ( .A(n25107), .B(n25108), .X(n25106) );
  nand_x1_sg U73754 ( .A(n51313), .B(n57322), .X(n25107) );
  nand_x1_sg U73755 ( .A(n57496), .B(n47463), .X(n25108) );
  nand_x2_sg U73756 ( .A(n25137), .B(n25138), .X(n25136) );
  nand_x1_sg U73757 ( .A(n56771), .B(n57322), .X(n25137) );
  nand_x1_sg U73758 ( .A(n57496), .B(n47453), .X(n25138) );
  nand_x2_sg U73759 ( .A(n25167), .B(n25168), .X(n25166) );
  nand_x1_sg U73760 ( .A(n51375), .B(n57322), .X(n25167) );
  nand_x1_sg U73761 ( .A(n57496), .B(n47385), .X(n25168) );
  nand_x2_sg U73762 ( .A(n25197), .B(n25198), .X(n25196) );
  nand_x1_sg U73763 ( .A(n56821), .B(n57322), .X(n25197) );
  nand_x1_sg U73764 ( .A(n57496), .B(n47325), .X(n25198) );
  nand_x2_sg U73765 ( .A(n25227), .B(n25228), .X(n25226) );
  nand_x1_sg U73766 ( .A(n51315), .B(n57322), .X(n25227) );
  nand_x1_sg U73767 ( .A(n57496), .B(n47495), .X(n25228) );
  nand_x2_sg U73768 ( .A(n25257), .B(n25258), .X(n25256) );
  nand_x1_sg U73769 ( .A(n56773), .B(n57322), .X(n25257) );
  nand_x1_sg U73770 ( .A(n57496), .B(n47302), .X(n25258) );
  nand_x2_sg U73771 ( .A(n25287), .B(n25288), .X(n25286) );
  nand_x1_sg U73772 ( .A(n56863), .B(n57322), .X(n25287) );
  nand_x1_sg U73773 ( .A(n57496), .B(n47473), .X(n25288) );
  nand_x2_sg U73774 ( .A(n25317), .B(n25318), .X(n25316) );
  nand_x1_sg U73775 ( .A(n47705), .B(n57322), .X(n25317) );
  nand_x1_sg U73776 ( .A(n57496), .B(n47323), .X(n25318) );
  nand_x2_sg U73777 ( .A(n25347), .B(n25348), .X(n25346) );
  nand_x1_sg U73778 ( .A(n51413), .B(n57322), .X(n25347) );
  nand_x1_sg U73779 ( .A(n57496), .B(n47489), .X(n25348) );
  nand_x2_sg U73780 ( .A(n25378), .B(n25379), .X(n25377) );
  nand_x1_sg U73781 ( .A(n56777), .B(n57322), .X(n25378) );
  nand_x1_sg U73782 ( .A(n57496), .B(n47465), .X(n25379) );
  nand_x2_sg U73783 ( .A(n25409), .B(n25410), .X(n25408) );
  nand_x1_sg U73784 ( .A(n47653), .B(n57322), .X(n25409) );
  nand_x1_sg U73785 ( .A(n57496), .B(n47449), .X(n25410) );
  nand_x2_sg U73786 ( .A(n25439), .B(n25440), .X(n25438) );
  nand_x1_sg U73787 ( .A(n47655), .B(n57322), .X(n25439) );
  nand_x1_sg U73788 ( .A(n57496), .B(n47383), .X(n25440) );
  nand_x2_sg U73789 ( .A(n25469), .B(n25470), .X(n25468) );
  nand_x1_sg U73790 ( .A(n51291), .B(n57322), .X(n25469) );
  nand_x1_sg U73791 ( .A(n57496), .B(n47457), .X(n25470) );
  nand_x2_sg U73792 ( .A(n25499), .B(n25500), .X(n25498) );
  nand_x1_sg U73793 ( .A(n51355), .B(n57322), .X(n25499) );
  nand_x1_sg U73794 ( .A(n57496), .B(n47479), .X(n25500) );
  nand_x2_sg U73795 ( .A(n25529), .B(n25530), .X(n25528) );
  nand_x1_sg U73796 ( .A(n56803), .B(n57322), .X(n25529) );
  nand_x1_sg U73797 ( .A(n57496), .B(n47469), .X(n25530) );
  nand_x2_sg U73798 ( .A(n25559), .B(n25560), .X(n25558) );
  nand_x1_sg U73799 ( .A(n47657), .B(n57322), .X(n25559) );
  nand_x1_sg U73800 ( .A(n57496), .B(n47451), .X(n25560) );
  nand_x2_sg U73801 ( .A(n25589), .B(n25590), .X(n25588) );
  nand_x1_sg U73802 ( .A(n51293), .B(n57322), .X(n25589) );
  nand_x1_sg U73803 ( .A(n57496), .B(n47485), .X(n25590) );
  nand_x2_sg U73804 ( .A(n25619), .B(n25620), .X(n25618) );
  nand_x1_sg U73805 ( .A(n56757), .B(n57322), .X(n25619) );
  nand_x1_sg U73806 ( .A(n57496), .B(n47459), .X(n25620) );
  nand_x2_sg U73807 ( .A(n25649), .B(n25650), .X(n25648) );
  nand_x1_sg U73808 ( .A(n51357), .B(n57322), .X(n25649) );
  nand_x1_sg U73809 ( .A(n57496), .B(n47381), .X(n25650) );
  nand_x2_sg U73810 ( .A(n25679), .B(n25680), .X(n25678) );
  nand_x1_sg U73811 ( .A(n56805), .B(n57322), .X(n25679) );
  nand_x1_sg U73812 ( .A(n57496), .B(n47321), .X(n25680) );
  nand_x2_sg U73813 ( .A(n25709), .B(n25710), .X(n25708) );
  nand_x1_sg U73814 ( .A(n51295), .B(n57322), .X(n25709) );
  nand_x1_sg U73815 ( .A(n57496), .B(n47308), .X(n25710) );
  nand_x2_sg U73816 ( .A(n25739), .B(n25740), .X(n25738) );
  nand_x1_sg U73817 ( .A(n56759), .B(n57322), .X(n25739) );
  nand_x1_sg U73818 ( .A(n57496), .B(n47291), .X(n25740) );
  nand_x2_sg U73819 ( .A(n25769), .B(n25770), .X(n25768) );
  nand_x1_sg U73820 ( .A(n51359), .B(n57322), .X(n25769) );
  nand_x1_sg U73821 ( .A(n57496), .B(n47481), .X(n25770) );
  nand_x2_sg U73822 ( .A(n25799), .B(n25800), .X(n25798) );
  nand_x1_sg U73823 ( .A(n56807), .B(n57322), .X(n25799) );
  nand_x1_sg U73824 ( .A(n57496), .B(n47471), .X(n25800) );
  nand_x2_sg U73825 ( .A(n25829), .B(n25830), .X(n25828) );
  nand_x1_sg U73826 ( .A(n51297), .B(n57322), .X(n25829) );
  nand_x1_sg U73827 ( .A(n57496), .B(n47493), .X(n25830) );
  nand_x2_sg U73828 ( .A(n25859), .B(n25860), .X(n25858) );
  nand_x1_sg U73829 ( .A(n56761), .B(n57322), .X(n25859) );
  nand_x1_sg U73830 ( .A(n57496), .B(n47461), .X(n25860) );
  nand_x2_sg U73831 ( .A(n25889), .B(n25890), .X(n25888) );
  nand_x1_sg U73832 ( .A(n56861), .B(n57322), .X(n25889) );
  nand_x1_sg U73833 ( .A(n57496), .B(n47379), .X(n25890) );
  nand_x2_sg U73834 ( .A(n25919), .B(n25920), .X(n25918) );
  nand_x1_sg U73835 ( .A(n47701), .B(n57322), .X(n25919) );
  nand_x1_sg U73836 ( .A(n57496), .B(n47377), .X(n25920) );
  nand_x2_sg U73837 ( .A(n25949), .B(n25950), .X(n25948) );
  nand_x1_sg U73838 ( .A(n51411), .B(n57322), .X(n25949) );
  nand_x1_sg U73839 ( .A(n57496), .B(n47327), .X(n25950) );
  nand_x2_sg U73840 ( .A(n25980), .B(n25981), .X(n25979) );
  nand_x1_sg U73841 ( .A(n56775), .B(n57322), .X(n25980) );
  nand_x1_sg U73842 ( .A(n57496), .B(n47306), .X(n25981) );
  nand_x1_sg U73843 ( .A(n56953), .B(n57464), .X(n23220) );
  nand_x1_sg U73844 ( .A(n56955), .B(n57464), .X(n23225) );
  nand_x1_sg U73845 ( .A(n56957), .B(n57464), .X(n23245) );
  nand_x1_sg U73846 ( .A(n56959), .B(n57464), .X(n23250) );
  nand_x1_sg U73847 ( .A(n56961), .B(n57464), .X(n23265) );
  nand_x1_sg U73848 ( .A(n56963), .B(n57464), .X(n23270) );
  nand_x1_sg U73849 ( .A(n56965), .B(n57464), .X(n23290) );
  nand_x1_sg U73850 ( .A(n56967), .B(n57464), .X(n23295) );
  nand_x1_sg U73851 ( .A(n56937), .B(n57472), .X(n23328) );
  nand_x1_sg U73852 ( .A(n56939), .B(n57472), .X(n23333) );
  nand_x1_sg U73853 ( .A(n56941), .B(n57472), .X(n23353) );
  nand_x1_sg U73854 ( .A(n56943), .B(n57472), .X(n23358) );
  nand_x1_sg U73855 ( .A(n56945), .B(n57472), .X(n23373) );
  nand_x1_sg U73856 ( .A(n56947), .B(n57472), .X(n23378) );
  nand_x1_sg U73857 ( .A(n56949), .B(n57472), .X(n23398) );
  nand_x1_sg U73858 ( .A(n56951), .B(n57472), .X(n23403) );
  nor_x1_sg U73859 ( .A(n22395), .B(n58611), .X(\shifter_0/n10205 ) );
  nand_x1_sg U73860 ( .A(n26121), .B(n51031), .X(n26156) );
  nand_x1_sg U73861 ( .A(n26122), .B(n47577), .X(n26155) );
  nand_x1_sg U73862 ( .A(n26121), .B(n51035), .X(n26120) );
  nand_x1_sg U73863 ( .A(n26122), .B(n47579), .X(n26119) );
  nand_x1_sg U73864 ( .A(n26121), .B(n51039), .X(n26248) );
  nand_x1_sg U73865 ( .A(n26122), .B(n47581), .X(n26247) );
  nand_x1_sg U73866 ( .A(n26121), .B(n51043), .X(n26214) );
  nand_x1_sg U73867 ( .A(n26122), .B(n47583), .X(n26213) );
  nand_x2_sg U73868 ( .A(n26139), .B(n26140), .X(n26138) );
  nand_x1_sg U73869 ( .A(n47497), .B(n67532), .X(n26139) );
  nand_x1_sg U73870 ( .A(n47589), .B(n67536), .X(n26140) );
  nand_x2_sg U73871 ( .A(n26100), .B(n26101), .X(n26099) );
  nand_x1_sg U73872 ( .A(n47499), .B(n67532), .X(n26100) );
  nand_x1_sg U73873 ( .A(n47591), .B(n67536), .X(n26101) );
  nand_x2_sg U73874 ( .A(n26231), .B(n26232), .X(n26230) );
  nand_x1_sg U73875 ( .A(n47501), .B(n67532), .X(n26231) );
  nand_x1_sg U73876 ( .A(n47593), .B(n67536), .X(n26232) );
  nand_x2_sg U73877 ( .A(n26197), .B(n26198), .X(n26196) );
  nand_x1_sg U73878 ( .A(n47503), .B(n67532), .X(n26197) );
  nand_x1_sg U73879 ( .A(n47595), .B(n67536), .X(n26198) );
  nor_x1_sg U73880 ( .A(n68208), .B(n26249), .X(\filter_0/n10776 ) );
  nor_x1_sg U73881 ( .A(n68207), .B(n26249), .X(\filter_0/n10772 ) );
  nor_x1_sg U73882 ( .A(n68188), .B(n26250), .X(\filter_0/n10696 ) );
  nor_x1_sg U73883 ( .A(n68187), .B(n26250), .X(\filter_0/n10692 ) );
  nor_x1_sg U73884 ( .A(n68168), .B(n26251), .X(\filter_0/n10616 ) );
  nor_x1_sg U73885 ( .A(n68167), .B(n26251), .X(\filter_0/n10612 ) );
  nor_x1_sg U73886 ( .A(n68148), .B(n26252), .X(\filter_0/n10536 ) );
  nor_x1_sg U73887 ( .A(n68147), .B(n26252), .X(\filter_0/n10532 ) );
  nor_x1_sg U73888 ( .A(n68128), .B(n26253), .X(\filter_0/n10456 ) );
  nor_x1_sg U73889 ( .A(n68127), .B(n26253), .X(\filter_0/n10452 ) );
  nor_x1_sg U73890 ( .A(n68108), .B(n26254), .X(\filter_0/n10376 ) );
  nor_x1_sg U73891 ( .A(n68107), .B(n26254), .X(\filter_0/n10372 ) );
  nor_x1_sg U73892 ( .A(n68088), .B(n26255), .X(\filter_0/n10296 ) );
  nor_x1_sg U73893 ( .A(n68087), .B(n26255), .X(\filter_0/n10292 ) );
  nor_x1_sg U73894 ( .A(n68068), .B(n26256), .X(\filter_0/n10216 ) );
  nor_x1_sg U73895 ( .A(n68067), .B(n26256), .X(\filter_0/n10212 ) );
  nor_x1_sg U73896 ( .A(n68048), .B(n26257), .X(\filter_0/n10136 ) );
  nor_x1_sg U73897 ( .A(n68047), .B(n26257), .X(\filter_0/n10132 ) );
  nor_x1_sg U73898 ( .A(n68028), .B(n26259), .X(\filter_0/n10056 ) );
  nor_x1_sg U73899 ( .A(n68027), .B(n26259), .X(\filter_0/n10052 ) );
  nor_x1_sg U73900 ( .A(n68015), .B(n26006), .X(\filter_0/n10004 ) );
  nor_x1_sg U73901 ( .A(n68014), .B(n26006), .X(\filter_0/n10000 ) );
  nor_x1_sg U73902 ( .A(n67988), .B(n26007), .X(\filter_0/n9896 ) );
  nor_x1_sg U73903 ( .A(n67987), .B(n26007), .X(\filter_0/n9892 ) );
  nor_x1_sg U73904 ( .A(n67968), .B(n26009), .X(\filter_0/n9816 ) );
  nor_x1_sg U73905 ( .A(n67967), .B(n26009), .X(\filter_0/n9812 ) );
  nor_x1_sg U73906 ( .A(n67948), .B(n26011), .X(\filter_0/n9736 ) );
  nor_x1_sg U73907 ( .A(n67947), .B(n26011), .X(\filter_0/n9732 ) );
  nor_x1_sg U73908 ( .A(n67928), .B(n26013), .X(\filter_0/n9656 ) );
  nor_x1_sg U73909 ( .A(n67927), .B(n26013), .X(\filter_0/n9652 ) );
  nor_x1_sg U73910 ( .A(n67908), .B(n26015), .X(\filter_0/n9576 ) );
  nor_x1_sg U73911 ( .A(n67907), .B(n26015), .X(\filter_0/n9572 ) );
  nor_x1_sg U73912 ( .A(n67888), .B(n26016), .X(\filter_0/n9496 ) );
  nor_x1_sg U73913 ( .A(n67887), .B(n26016), .X(\filter_0/n9492 ) );
  nor_x1_sg U73914 ( .A(n67868), .B(n26018), .X(\filter_0/n9416 ) );
  nor_x1_sg U73915 ( .A(n67867), .B(n26018), .X(\filter_0/n9412 ) );
  nor_x1_sg U73916 ( .A(n67848), .B(n26020), .X(\filter_0/n9336 ) );
  nor_x1_sg U73917 ( .A(n67847), .B(n26020), .X(\filter_0/n9332 ) );
  nor_x1_sg U73918 ( .A(n67828), .B(n26022), .X(\filter_0/n9256 ) );
  nor_x1_sg U73919 ( .A(n67827), .B(n26022), .X(\filter_0/n9252 ) );
  nor_x1_sg U73920 ( .A(n67808), .B(n26024), .X(\filter_0/n9176 ) );
  nor_x1_sg U73921 ( .A(n67807), .B(n26024), .X(\filter_0/n9172 ) );
  nor_x1_sg U73922 ( .A(n67788), .B(n26025), .X(\filter_0/n9096 ) );
  nor_x1_sg U73923 ( .A(n67787), .B(n26025), .X(\filter_0/n9092 ) );
  nor_x1_sg U73924 ( .A(n67768), .B(n26026), .X(\filter_0/n9016 ) );
  nor_x1_sg U73925 ( .A(n67767), .B(n26026), .X(\filter_0/n9012 ) );
  nor_x1_sg U73926 ( .A(n67748), .B(n26027), .X(\filter_0/n8936 ) );
  nor_x1_sg U73927 ( .A(n67747), .B(n26027), .X(\filter_0/n8932 ) );
  nor_x1_sg U73928 ( .A(n67728), .B(n26028), .X(\filter_0/n8856 ) );
  nor_x1_sg U73929 ( .A(n67727), .B(n26028), .X(\filter_0/n8852 ) );
  nor_x1_sg U73930 ( .A(n67708), .B(n26029), .X(\filter_0/n8776 ) );
  nor_x1_sg U73931 ( .A(n67707), .B(n26029), .X(\filter_0/n8772 ) );
  nor_x1_sg U73932 ( .A(n67688), .B(n26030), .X(\filter_0/n8696 ) );
  nor_x1_sg U73933 ( .A(n67687), .B(n26030), .X(\filter_0/n8692 ) );
  nor_x1_sg U73934 ( .A(n67668), .B(n26031), .X(\filter_0/n8616 ) );
  nor_x1_sg U73935 ( .A(n67667), .B(n26031), .X(\filter_0/n8612 ) );
  nor_x1_sg U73936 ( .A(n67648), .B(n26032), .X(\filter_0/n8536 ) );
  nor_x1_sg U73937 ( .A(n67647), .B(n26032), .X(\filter_0/n8532 ) );
  nor_x1_sg U73938 ( .A(n67628), .B(n26035), .X(\filter_0/n8456 ) );
  nor_x1_sg U73939 ( .A(n67627), .B(n26035), .X(\filter_0/n8452 ) );
  nor_x1_sg U73940 ( .A(n67608), .B(n26037), .X(\filter_0/n8376 ) );
  nor_x1_sg U73941 ( .A(n67607), .B(n26037), .X(\filter_0/n8372 ) );
  nor_x1_sg U73942 ( .A(n67588), .B(n26038), .X(\filter_0/n8296 ) );
  nor_x1_sg U73943 ( .A(n67587), .B(n26038), .X(\filter_0/n8292 ) );
  nor_x1_sg U73944 ( .A(n22750), .B(n22654), .X(\shifter_0/n11724 ) );
  nor_x1_sg U73945 ( .A(n22764), .B(n22656), .X(\shifter_0/n11720 ) );
  nor_x1_sg U73946 ( .A(n22775), .B(n22658), .X(\shifter_0/n11716 ) );
  nor_x1_sg U73947 ( .A(n22786), .B(n22660), .X(\shifter_0/n11712 ) );
  nor_x1_sg U73948 ( .A(n22797), .B(n22662), .X(\shifter_0/n11708 ) );
  nor_x1_sg U73949 ( .A(n22808), .B(n22664), .X(\shifter_0/n11704 ) );
  nor_x1_sg U73950 ( .A(n22819), .B(n22666), .X(\shifter_0/n11700 ) );
  nor_x1_sg U73951 ( .A(n22830), .B(n22668), .X(\shifter_0/n11696 ) );
  nor_x1_sg U73952 ( .A(n22841), .B(n22670), .X(\shifter_0/n11692 ) );
  nor_x1_sg U73953 ( .A(n22852), .B(n22672), .X(\shifter_0/n11688 ) );
  nor_x1_sg U73954 ( .A(n22863), .B(n22674), .X(\shifter_0/n11684 ) );
  nor_x1_sg U73955 ( .A(n22874), .B(n22676), .X(\shifter_0/n11680 ) );
  nor_x1_sg U73956 ( .A(n22885), .B(n22678), .X(\shifter_0/n11676 ) );
  nor_x1_sg U73957 ( .A(n22896), .B(n22680), .X(\shifter_0/n11672 ) );
  nor_x1_sg U73958 ( .A(n22907), .B(n22682), .X(\shifter_0/n11668 ) );
  nor_x1_sg U73959 ( .A(n22918), .B(n22684), .X(\shifter_0/n11664 ) );
  nor_x1_sg U73960 ( .A(n22929), .B(n22686), .X(\shifter_0/n11660 ) );
  nor_x1_sg U73961 ( .A(n22940), .B(n22688), .X(\shifter_0/n11656 ) );
  nor_x1_sg U73962 ( .A(n22951), .B(n22690), .X(\shifter_0/n11652 ) );
  nor_x1_sg U73963 ( .A(n22962), .B(n22692), .X(\shifter_0/n11648 ) );
  nor_x1_sg U73964 ( .A(n22978), .B(n22701), .X(\shifter_0/n11644 ) );
  nor_x1_sg U73965 ( .A(n22991), .B(n22703), .X(\shifter_0/n11640 ) );
  nor_x1_sg U73966 ( .A(n23002), .B(n22705), .X(\shifter_0/n11636 ) );
  nor_x1_sg U73967 ( .A(n23013), .B(n22707), .X(\shifter_0/n11632 ) );
  nor_x1_sg U73968 ( .A(n23024), .B(n22709), .X(\shifter_0/n11628 ) );
  nor_x1_sg U73969 ( .A(n23035), .B(n22711), .X(\shifter_0/n11624 ) );
  nor_x1_sg U73970 ( .A(n23046), .B(n22713), .X(\shifter_0/n11620 ) );
  nor_x1_sg U73971 ( .A(n23057), .B(n22715), .X(\shifter_0/n11616 ) );
  nor_x1_sg U73972 ( .A(n23068), .B(n22717), .X(\shifter_0/n11612 ) );
  nor_x1_sg U73973 ( .A(n23079), .B(n22719), .X(\shifter_0/n11608 ) );
  nor_x1_sg U73974 ( .A(n23090), .B(n22721), .X(\shifter_0/n11604 ) );
  nor_x1_sg U73975 ( .A(n23101), .B(n22723), .X(\shifter_0/n11600 ) );
  nor_x1_sg U73976 ( .A(n23112), .B(n22725), .X(\shifter_0/n11596 ) );
  nor_x1_sg U73977 ( .A(n23123), .B(n22727), .X(\shifter_0/n11592 ) );
  nor_x1_sg U73978 ( .A(n23134), .B(n22729), .X(\shifter_0/n11588 ) );
  nor_x1_sg U73979 ( .A(n23145), .B(n22731), .X(\shifter_0/n11584 ) );
  nor_x1_sg U73980 ( .A(n23156), .B(n22733), .X(\shifter_0/n11580 ) );
  nor_x1_sg U73981 ( .A(n23167), .B(n22735), .X(\shifter_0/n11576 ) );
  nor_x1_sg U73982 ( .A(n23178), .B(n22737), .X(\shifter_0/n11572 ) );
  nor_x1_sg U73983 ( .A(n23189), .B(n22739), .X(\shifter_0/n11568 ) );
  nand_x2_sg U73984 ( .A(n26131), .B(n26132), .X(n26130) );
  nand_x1_sg U73985 ( .A(n57106), .B(n51029), .X(n26131) );
  nand_x1_sg U73986 ( .A(n57109), .B(n53597), .X(n26132) );
  nand_x2_sg U73987 ( .A(n26089), .B(n26090), .X(n26088) );
  nand_x1_sg U73988 ( .A(n57106), .B(n51033), .X(n26089) );
  nand_x1_sg U73989 ( .A(n57109), .B(n53611), .X(n26090) );
  nand_x2_sg U73990 ( .A(n26223), .B(n26224), .X(n26222) );
  nand_x1_sg U73991 ( .A(n57106), .B(n51037), .X(n26223) );
  nand_x1_sg U73992 ( .A(n57109), .B(n53625), .X(n26224) );
  nand_x2_sg U73993 ( .A(n26189), .B(n26190), .X(n26188) );
  nand_x1_sg U73994 ( .A(n57106), .B(n51041), .X(n26189) );
  nand_x1_sg U73995 ( .A(n57109), .B(n53639), .X(n26190) );
  nand_x1_sg U73996 ( .A(n67240), .B(n57468), .X(n23207) );
  nand_x1_sg U73997 ( .A(n67238), .B(n57468), .X(n23212) );
  nand_x1_sg U73998 ( .A(n67236), .B(n57468), .X(n23217) );
  nand_x1_sg U73999 ( .A(n67230), .B(n57468), .X(n23232) );
  nand_x1_sg U74000 ( .A(n67228), .B(n57468), .X(n23237) );
  nand_x1_sg U74001 ( .A(n67226), .B(n57468), .X(n23242) );
  nand_x1_sg U74002 ( .A(n67220), .B(n57468), .X(n23257) );
  nand_x1_sg U74003 ( .A(n67218), .B(n57468), .X(n23262) );
  nand_x1_sg U74004 ( .A(n67212), .B(n57468), .X(n23277) );
  nand_x1_sg U74005 ( .A(n67210), .B(n57468), .X(n23282) );
  nand_x1_sg U74006 ( .A(n67208), .B(n57468), .X(n23287) );
  nand_x1_sg U74007 ( .A(n67202), .B(n57468), .X(n23302) );
  nand_x1_sg U74008 ( .A(n67433), .B(n57476), .X(n23315) );
  nand_x1_sg U74009 ( .A(n67431), .B(n57476), .X(n23320) );
  nand_x1_sg U74010 ( .A(n67429), .B(n57476), .X(n23325) );
  nand_x1_sg U74011 ( .A(n67423), .B(n57476), .X(n23340) );
  nand_x1_sg U74012 ( .A(n67421), .B(n57476), .X(n23345) );
  nand_x1_sg U74013 ( .A(n67419), .B(n57476), .X(n23350) );
  nand_x1_sg U74014 ( .A(n67413), .B(n57476), .X(n23365) );
  nand_x1_sg U74015 ( .A(n67411), .B(n57476), .X(n23370) );
  nand_x1_sg U74016 ( .A(n67405), .B(n57476), .X(n23385) );
  nand_x1_sg U74017 ( .A(n67403), .B(n57476), .X(n23390) );
  nand_x1_sg U74018 ( .A(n67401), .B(n57476), .X(n23395) );
  nand_x1_sg U74019 ( .A(n67395), .B(n57476), .X(n23410) );
  inv_x8_sg U74020 ( .A(n57098), .X(n57099) );
  inv_x8_sg U74021 ( .A(n57296), .X(n57100) );
  inv_x8_sg U74022 ( .A(n57101), .X(n57102) );
  nand_x8_sg U74023 ( .A(n57950), .B(n57925), .X(n57103) );
  nand_x8_sg U74024 ( .A(n57950), .B(n57925), .X(n57104) );
  inv_x8_sg U74025 ( .A(n57105), .X(n57106) );
  inv_x8_sg U74026 ( .A(n26303), .X(n57107) );
  inv_x8_sg U74027 ( .A(n57108), .X(n57109) );
  inv_x8_sg U74028 ( .A(n57110), .X(n57111) );
  inv_x8_sg U74029 ( .A(n57112), .X(n57113) );
  inv_x8_sg U74030 ( .A(n57113), .X(n57114) );
  inv_x8_sg U74031 ( .A(n25401), .X(n57115) );
  inv_x8_sg U74032 ( .A(n57115), .X(n57116) );
  inv_x8_sg U74033 ( .A(n24790), .X(n57117) );
  inv_x8_sg U74034 ( .A(n57117), .X(n57118) );
  inv_x8_sg U74035 ( .A(n57121), .X(n57119) );
  nand_x8_sg U74036 ( .A(n24777), .B(n24778), .X(n57120) );
  nand_x8_sg U74037 ( .A(n24777), .B(n24778), .X(n57121) );
  inv_x8_sg U74038 ( .A(n57124), .X(n57122) );
  nand_x8_sg U74039 ( .A(n24683), .B(n24684), .X(n57123) );
  nand_x8_sg U74040 ( .A(n24683), .B(n24684), .X(n57124) );
  inv_x8_sg U74041 ( .A(n57127), .X(n57125) );
  nand_x8_sg U74042 ( .A(n24589), .B(n24590), .X(n57126) );
  nand_x8_sg U74043 ( .A(n24589), .B(n24590), .X(n57127) );
  inv_x8_sg U74044 ( .A(n57130), .X(n57128) );
  nand_x8_sg U74045 ( .A(n24477), .B(n24478), .X(n57129) );
  nand_x8_sg U74046 ( .A(n24477), .B(n24478), .X(n57130) );
  inv_x8_sg U74047 ( .A(n24272), .X(n57131) );
  nand_x8_sg U74048 ( .A(n24368), .B(n24369), .X(n57132) );
  inv_x8_sg U74049 ( .A(n57135), .X(n57133) );
  nand_x8_sg U74050 ( .A(n24259), .B(n24260), .X(n57134) );
  nand_x8_sg U74051 ( .A(n24259), .B(n24260), .X(n57135) );
  inv_x8_sg U74052 ( .A(n57138), .X(n57136) );
  nand_x8_sg U74053 ( .A(n23931), .B(n23932), .X(n57137) );
  nand_x8_sg U74054 ( .A(n23931), .B(n23932), .X(n57138) );
  inv_x8_sg U74055 ( .A(n57141), .X(n57139) );
  nand_x8_sg U74056 ( .A(n23802), .B(n23803), .X(n57140) );
  nand_x8_sg U74057 ( .A(n23802), .B(n23803), .X(n57141) );
  inv_x8_sg U74058 ( .A(n57144), .X(n57142) );
  nand_x8_sg U74059 ( .A(n23671), .B(n23672), .X(n57143) );
  nand_x8_sg U74060 ( .A(n23671), .B(n23672), .X(n57144) );
  inv_x8_sg U74061 ( .A(n57147), .X(n57145) );
  nand_x8_sg U74062 ( .A(n23539), .B(n23540), .X(n57146) );
  nand_x8_sg U74063 ( .A(n23539), .B(n23540), .X(n57147) );
  nor_x8_sg U74064 ( .A(n22988), .B(n68588), .X(n57148) );
  nor_x8_sg U74065 ( .A(n22988), .B(n68588), .X(n22977) );
  inv_x8_sg U74066 ( .A(n57152), .X(n57149) );
  inv_x8_sg U74067 ( .A(n57150), .X(n57151) );
  nand_x8_sg U74068 ( .A(n57302), .B(n23198), .X(n57152) );
  nand_x8_sg U74069 ( .A(n57302), .B(n23198), .X(n57153) );
  nor_x8_sg U74070 ( .A(n22761), .B(n68588), .X(n57154) );
  nor_x8_sg U74071 ( .A(n22761), .B(n68588), .X(n22749) );
  inv_x8_sg U74072 ( .A(n57158), .X(n57155) );
  inv_x8_sg U74073 ( .A(n57156), .X(n57157) );
  nand_x8_sg U74074 ( .A(n57097), .B(n22971), .X(n57158) );
  nand_x8_sg U74075 ( .A(n57097), .B(n22971), .X(n57159) );
  nand_x8_sg U74076 ( .A(n22740), .B(n22741), .X(n57160) );
  nand_x8_sg U74077 ( .A(n22740), .B(n22741), .X(n57161) );
  inv_x8_sg U74078 ( .A(n57161), .X(n57162) );
  nand_x8_sg U74079 ( .A(n22693), .B(n22694), .X(n57163) );
  nand_x8_sg U74080 ( .A(n22693), .B(n22694), .X(n57164) );
  inv_x8_sg U74081 ( .A(n57164), .X(n57165) );
  inv_x8_sg U74082 ( .A(n29338), .X(n68389) );
  inv_x8_sg U74083 ( .A(n57168), .X(n57166) );
  inv_x8_sg U74084 ( .A(n57167), .X(n57168) );
  inv_x8_sg U74085 ( .A(n57169), .X(n57170) );
  inv_x8_sg U74086 ( .A(n57171), .X(n57172) );
  inv_x8_sg U74087 ( .A(n57173), .X(n57174) );
  nor_x4_sg U74088 ( .A(n57172), .B(n57854), .X(n34179) );
  inv_x8_sg U74089 ( .A(n57175), .X(n57176) );
  inv_x8_sg U74090 ( .A(n57177), .X(n57178) );
  nor_x4_sg U74091 ( .A(n57176), .B(n57854), .X(n34134) );
  nand_x8_sg U74092 ( .A(n33955), .B(n33524), .X(n57179) );
  inv_x8_sg U74093 ( .A(n57180), .X(n57181) );
  nor_x4_sg U74094 ( .A(n57179), .B(n57854), .X(n34091) );
  inv_x8_sg U74095 ( .A(n57182), .X(n57183) );
  inv_x8_sg U74096 ( .A(n57184), .X(n57185) );
  nor_x4_sg U74097 ( .A(n57183), .B(n57854), .X(n34046) );
  inv_x8_sg U74098 ( .A(n57186), .X(n57187) );
  inv_x8_sg U74099 ( .A(n57188), .X(n57189) );
  nor_x4_sg U74100 ( .A(n57187), .B(n57854), .X(n34001) );
  nand_x8_sg U74101 ( .A(n33955), .B(n33051), .X(n57190) );
  nand_x8_sg U74102 ( .A(n33955), .B(n33051), .X(n57191) );
  inv_x8_sg U74103 ( .A(n57192), .X(n57193) );
  nor_x4_sg U74104 ( .A(n33959), .B(n57855), .X(n33958) );
  nand_x8_sg U74105 ( .A(n33955), .B(n33094), .X(n57194) );
  nand_x8_sg U74106 ( .A(n33955), .B(n33094), .X(n57195) );
  inv_x8_sg U74107 ( .A(n57196), .X(n57197) );
  nor_x4_sg U74108 ( .A(n33916), .B(n57855), .X(n33915) );
  inv_x8_sg U74109 ( .A(n57198), .X(n57199) );
  inv_x8_sg U74110 ( .A(n57200), .X(n57201) );
  nor_x4_sg U74111 ( .A(n57199), .B(n57855), .X(n33871) );
  nand_x8_sg U74112 ( .A(n33265), .B(n33008), .X(n57202) );
  inv_x8_sg U74113 ( .A(n57203), .X(n57204) );
  nor_x4_sg U74114 ( .A(n57202), .B(n57855), .X(n33828) );
  nand_x8_sg U74115 ( .A(n33222), .B(n33008), .X(n57205) );
  inv_x8_sg U74116 ( .A(n57206), .X(n57207) );
  nor_x4_sg U74117 ( .A(n57205), .B(n57855), .X(n33786) );
  inv_x8_sg U74118 ( .A(n57208), .X(n57209) );
  inv_x8_sg U74119 ( .A(n57210), .X(n57211) );
  nor_x4_sg U74120 ( .A(n57209), .B(n57855), .X(n33741) );
  nand_x8_sg U74121 ( .A(n33222), .B(n33609), .X(n57212) );
  nand_x8_sg U74122 ( .A(n33222), .B(n33609), .X(n57213) );
  inv_x8_sg U74123 ( .A(n57214), .X(n57215) );
  nor_x4_sg U74124 ( .A(n33699), .B(n57855), .X(n33698) );
  nand_x8_sg U74125 ( .A(n33265), .B(n33609), .X(n57216) );
  nand_x8_sg U74126 ( .A(n33265), .B(n33609), .X(n57217) );
  inv_x8_sg U74127 ( .A(n57218), .X(n57219) );
  nor_x4_sg U74128 ( .A(n33657), .B(n57855), .X(n33656) );
  nand_x8_sg U74129 ( .A(n68230), .B(n33609), .X(n57220) );
  nand_x8_sg U74130 ( .A(n68230), .B(n33609), .X(n57221) );
  inv_x8_sg U74131 ( .A(n57222), .X(n57223) );
  nor_x4_sg U74132 ( .A(n33613), .B(n57855), .X(n33612) );
  nand_x8_sg U74133 ( .A(n68229), .B(n33609), .X(n57224) );
  inv_x8_sg U74134 ( .A(n57225), .X(n57226) );
  nor_x4_sg U74135 ( .A(n57224), .B(n57854), .X(n33569) );
  nand_x8_sg U74136 ( .A(n33309), .B(n33524), .X(n57227) );
  inv_x8_sg U74137 ( .A(n57228), .X(n57229) );
  nor_x4_sg U74138 ( .A(n57227), .B(n57854), .X(n33527) );
  nand_x8_sg U74139 ( .A(n68228), .B(n33524), .X(n57230) );
  inv_x8_sg U74140 ( .A(n57231), .X(n57232) );
  nor_x4_sg U74141 ( .A(n57230), .B(n57854), .X(n33484) );
  nand_x8_sg U74142 ( .A(n68228), .B(n33051), .X(n57233) );
  nand_x8_sg U74143 ( .A(n68228), .B(n33051), .X(n57234) );
  inv_x8_sg U74144 ( .A(n57235), .X(n57236) );
  nor_x4_sg U74145 ( .A(n33443), .B(n57854), .X(n33442) );
  nand_x8_sg U74146 ( .A(n33309), .B(n33051), .X(n57237) );
  nand_x8_sg U74147 ( .A(n33309), .B(n33051), .X(n57238) );
  inv_x8_sg U74148 ( .A(n57239), .X(n57240) );
  nor_x4_sg U74149 ( .A(n33401), .B(n57854), .X(n33400) );
  nand_x8_sg U74150 ( .A(n68231), .B(n33310), .X(n57241) );
  nand_x8_sg U74151 ( .A(n68231), .B(n33310), .X(n57242) );
  inv_x8_sg U74152 ( .A(n57243), .X(n57244) );
  nor_x4_sg U74153 ( .A(n33356), .B(n57854), .X(n33355) );
  nand_x8_sg U74154 ( .A(n68228), .B(n33310), .X(n57245) );
  nand_x8_sg U74155 ( .A(n68228), .B(n33310), .X(n57246) );
  inv_x8_sg U74156 ( .A(n57247), .X(n57248) );
  nor_x4_sg U74157 ( .A(n33314), .B(n57854), .X(n33313) );
  nand_x8_sg U74158 ( .A(n33309), .B(n33310), .X(n57249) );
  nand_x8_sg U74159 ( .A(n33309), .B(n33310), .X(n57250) );
  inv_x8_sg U74160 ( .A(n57251), .X(n57252) );
  nor_x4_sg U74161 ( .A(n33270), .B(n57854), .X(n33269) );
  nand_x8_sg U74162 ( .A(n33265), .B(n33179), .X(n57253) );
  nand_x8_sg U74163 ( .A(n33265), .B(n33179), .X(n57254) );
  inv_x8_sg U74164 ( .A(n57255), .X(n57256) );
  nor_x4_sg U74165 ( .A(n33226), .B(n57854), .X(n33225) );
  nand_x8_sg U74166 ( .A(n33222), .B(n33179), .X(n57257) );
  nand_x8_sg U74167 ( .A(n33222), .B(n33179), .X(n57258) );
  inv_x8_sg U74168 ( .A(n57259), .X(n57260) );
  nor_x4_sg U74169 ( .A(n33183), .B(n57855), .X(n33182) );
  nand_x8_sg U74170 ( .A(n68229), .B(n33179), .X(n57261) );
  nand_x8_sg U74171 ( .A(n68229), .B(n33179), .X(n57262) );
  inv_x8_sg U74172 ( .A(n57263), .X(n57264) );
  nor_x4_sg U74173 ( .A(n33140), .B(n57854), .X(n33139) );
  nand_x8_sg U74174 ( .A(n68229), .B(n32965), .X(n57265) );
  nand_x8_sg U74175 ( .A(n68229), .B(n32965), .X(n57266) );
  inv_x8_sg U74176 ( .A(n57267), .X(n57268) );
  nor_x4_sg U74177 ( .A(n33098), .B(n57854), .X(n33097) );
  nand_x8_sg U74178 ( .A(n68231), .B(n33094), .X(n57269) );
  nand_x8_sg U74179 ( .A(n68231), .B(n33094), .X(n57270) );
  inv_x8_sg U74180 ( .A(n57271), .X(n57272) );
  nor_x4_sg U74181 ( .A(n33055), .B(n57855), .X(n33054) );
  nand_x8_sg U74182 ( .A(n68231), .B(n33051), .X(n57273) );
  nand_x8_sg U74183 ( .A(n68231), .B(n33051), .X(n57274) );
  inv_x8_sg U74184 ( .A(n57275), .X(n57276) );
  nor_x4_sg U74185 ( .A(n33012), .B(n57854), .X(n33011) );
  nand_x8_sg U74186 ( .A(n68230), .B(n33008), .X(n57277) );
  nand_x8_sg U74187 ( .A(n68230), .B(n33008), .X(n57278) );
  inv_x8_sg U74188 ( .A(n57279), .X(n57280) );
  nor_x4_sg U74189 ( .A(n32969), .B(n57854), .X(n32968) );
  nand_x8_sg U74190 ( .A(n68230), .B(n32965), .X(n57281) );
  nand_x8_sg U74191 ( .A(n68230), .B(n32965), .X(n57282) );
  inv_x8_sg U74192 ( .A(n57283), .X(n57284) );
  nor_x4_sg U74193 ( .A(n32926), .B(n57855), .X(n32925) );
  inv_x8_sg U74194 ( .A(n57285), .X(n57286) );
  nor_x4_sg U74195 ( .A(n57168), .B(n47295), .X(n32881) );
  inv_x8_sg U74196 ( .A(n57287), .X(n57288) );
  nor_x4_sg U74197 ( .A(n57854), .B(n57286), .X(n32880) );
  inv_x8_sg U74198 ( .A(n57289), .X(n57290) );
  nor_x4_sg U74199 ( .A(n57168), .B(n47312), .X(n32835) );
  inv_x8_sg U74200 ( .A(n57291), .X(n57292) );
  nor_x4_sg U74201 ( .A(n57855), .B(n57290), .X(n32834) );
  inv_x8_sg U74202 ( .A(n57293), .X(n57294) );
  inv_x8_sg U74203 ( .A(n57295), .X(n57296) );
  inv_x8_sg U74204 ( .A(n57297), .X(n57298) );
  inv_x8_sg U74205 ( .A(n57299), .X(n57300) );
  inv_x8_sg U74206 ( .A(n57301), .X(n57302) );
  inv_x8_sg U74207 ( .A(n51053), .X(n57303) );
  inv_x8_sg U74208 ( .A(n57303), .X(n57304) );
  inv_x8_sg U74209 ( .A(n57305), .X(n57306) );
  inv_x8_sg U74210 ( .A(n51057), .X(n57307) );
  inv_x8_sg U74211 ( .A(n57307), .X(n57308) );
  inv_x8_sg U74212 ( .A(n57309), .X(n57310) );
  inv_x8_sg U74213 ( .A(n57312), .X(n57311) );
  inv_x8_sg U74214 ( .A(n57315), .X(n57314) );
  inv_x8_sg U74215 ( .A(n57317), .X(n57316) );
  inv_x8_sg U74216 ( .A(n57319), .X(n57318) );
  inv_x8_sg U74217 ( .A(n57321), .X(n57320) );
  inv_x8_sg U74218 ( .A(n57323), .X(n57322) );
  inv_x8_sg U74219 ( .A(n58657), .X(n57325) );
  inv_x4_sg U74220 ( .A(n57104), .X(n57326) );
  inv_x4_sg U74221 ( .A(n57103), .X(n57327) );
  inv_x8_sg U74222 ( .A(n58638), .X(n57328) );
  inv_x8_sg U74223 ( .A(n58656), .X(n57329) );
  inv_x4_sg U74224 ( .A(n57344), .X(n57330) );
  inv_x4_sg U74225 ( .A(n57344), .X(n57331) );
  inv_x4_sg U74226 ( .A(n57344), .X(n57332) );
  inv_x4_sg U74227 ( .A(n57344), .X(n57333) );
  inv_x4_sg U74228 ( .A(n57344), .X(n57334) );
  inv_x4_sg U74229 ( .A(n57344), .X(n57335) );
  inv_x4_sg U74230 ( .A(n57344), .X(n57336) );
  inv_x4_sg U74231 ( .A(n57344), .X(n57337) );
  inv_x4_sg U74232 ( .A(n57344), .X(n57338) );
  inv_x4_sg U74233 ( .A(n57344), .X(n57339) );
  inv_x4_sg U74234 ( .A(n57344), .X(n57340) );
  inv_x4_sg U74235 ( .A(n57344), .X(n57341) );
  inv_x4_sg U74236 ( .A(n57344), .X(n57342) );
  inv_x4_sg U74237 ( .A(n57344), .X(n57343) );
  inv_x8_sg U74238 ( .A(n58630), .X(n57344) );
  inv_x8_sg U74239 ( .A(n57346), .X(n57345) );
  inv_x8_sg U74240 ( .A(n58639), .X(n57348) );
  inv_x8_sg U74241 ( .A(n58639), .X(n57349) );
  inv_x8_sg U74242 ( .A(n57382), .X(n57350) );
  inv_x8_sg U74243 ( .A(n57382), .X(n57351) );
  inv_x8_sg U74244 ( .A(n57393), .X(n57352) );
  inv_x8_sg U74245 ( .A(n57386), .X(n57353) );
  inv_x8_sg U74246 ( .A(n57386), .X(n57354) );
  inv_x8_sg U74247 ( .A(n57386), .X(n57355) );
  inv_x8_sg U74248 ( .A(n57386), .X(n57356) );
  inv_x8_sg U74249 ( .A(n57385), .X(n57357) );
  inv_x8_sg U74250 ( .A(n57385), .X(n57358) );
  inv_x8_sg U74251 ( .A(n57385), .X(n57359) );
  inv_x8_sg U74252 ( .A(n57385), .X(n57360) );
  inv_x8_sg U74253 ( .A(n57384), .X(n57361) );
  inv_x8_sg U74254 ( .A(n57384), .X(n57362) );
  inv_x8_sg U74255 ( .A(n57384), .X(n57363) );
  inv_x8_sg U74256 ( .A(n57384), .X(n57364) );
  inv_x8_sg U74257 ( .A(n57383), .X(n57365) );
  inv_x8_sg U74258 ( .A(n57383), .X(n57366) );
  inv_x8_sg U74259 ( .A(n57383), .X(n57367) );
  inv_x8_sg U74260 ( .A(n57383), .X(n57368) );
  inv_x8_sg U74261 ( .A(n57386), .X(n57369) );
  inv_x8_sg U74262 ( .A(n57386), .X(n57370) );
  inv_x8_sg U74263 ( .A(n57382), .X(n57371) );
  inv_x8_sg U74264 ( .A(n57382), .X(n57372) );
  inv_x8_sg U74265 ( .A(n57392), .X(n57373) );
  inv_x8_sg U74266 ( .A(n57392), .X(n57374) );
  inv_x8_sg U74267 ( .A(n57392), .X(n57375) );
  inv_x8_sg U74268 ( .A(n57392), .X(n57376) );
  inv_x8_sg U74269 ( .A(n57382), .X(n57377) );
  inv_x8_sg U74270 ( .A(n57382), .X(n57378) );
  inv_x8_sg U74271 ( .A(n57382), .X(n57379) );
  inv_x8_sg U74272 ( .A(n57386), .X(n57380) );
  inv_x8_sg U74273 ( .A(n57382), .X(n57381) );
  inv_x8_sg U74274 ( .A(n61856), .X(n57382) );
  inv_x8_sg U74275 ( .A(n57391), .X(n57383) );
  inv_x8_sg U74276 ( .A(n57390), .X(n57384) );
  inv_x8_sg U74277 ( .A(n57389), .X(n57385) );
  inv_x8_sg U74278 ( .A(n57388), .X(n57386) );
  inv_x8_sg U74279 ( .A(n57393), .X(n57387) );
  inv_x8_sg U74280 ( .A(n57393), .X(n57388) );
  inv_x8_sg U74281 ( .A(n57392), .X(n57390) );
  inv_x8_sg U74282 ( .A(n61856), .X(n57392) );
  inv_x8_sg U74283 ( .A(n61856), .X(n57393) );
  inv_x8_sg U74284 ( .A(n57448), .X(n57394) );
  inv_x8_sg U74285 ( .A(n57436), .X(n57395) );
  inv_x8_sg U74286 ( .A(n57449), .X(n57396) );
  inv_x8_sg U74287 ( .A(n57448), .X(n57397) );
  inv_x8_sg U74288 ( .A(n57438), .X(n57398) );
  inv_x8_sg U74289 ( .A(n57438), .X(n57399) );
  inv_x8_sg U74290 ( .A(n57438), .X(n57400) );
  inv_x8_sg U74291 ( .A(n57438), .X(n57401) );
  inv_x8_sg U74292 ( .A(n57437), .X(n57402) );
  inv_x8_sg U74293 ( .A(n57437), .X(n57403) );
  inv_x8_sg U74294 ( .A(n57437), .X(n57404) );
  inv_x8_sg U74295 ( .A(n57437), .X(n57405) );
  inv_x8_sg U74296 ( .A(n57436), .X(n57406) );
  inv_x8_sg U74297 ( .A(n57436), .X(n57407) );
  inv_x8_sg U74298 ( .A(n57436), .X(n57408) );
  inv_x8_sg U74299 ( .A(n57436), .X(n57409) );
  inv_x8_sg U74300 ( .A(n57435), .X(n57410) );
  inv_x8_sg U74301 ( .A(n57435), .X(n57411) );
  inv_x8_sg U74302 ( .A(n57435), .X(n57412) );
  inv_x8_sg U74303 ( .A(n57435), .X(n57413) );
  inv_x8_sg U74304 ( .A(n57434), .X(n57414) );
  inv_x8_sg U74305 ( .A(n57434), .X(n57415) );
  inv_x8_sg U74306 ( .A(n57434), .X(n57416) );
  inv_x8_sg U74307 ( .A(n57434), .X(n57417) );
  inv_x8_sg U74308 ( .A(n57433), .X(n57418) );
  inv_x8_sg U74309 ( .A(n57433), .X(n57419) );
  inv_x8_sg U74310 ( .A(n57433), .X(n57420) );
  inv_x8_sg U74311 ( .A(n57433), .X(n57421) );
  inv_x8_sg U74312 ( .A(n57432), .X(n57422) );
  inv_x8_sg U74313 ( .A(n57432), .X(n57423) );
  inv_x8_sg U74314 ( .A(n57432), .X(n57424) );
  inv_x8_sg U74315 ( .A(n57432), .X(n57425) );
  inv_x8_sg U74316 ( .A(n57431), .X(n57426) );
  inv_x8_sg U74317 ( .A(n57431), .X(n57427) );
  inv_x8_sg U74318 ( .A(n57431), .X(n57428) );
  inv_x8_sg U74319 ( .A(n57431), .X(n57429) );
  inv_x8_sg U74320 ( .A(n57448), .X(n57430) );
  inv_x8_sg U74321 ( .A(n57446), .X(n57431) );
  inv_x8_sg U74322 ( .A(n57445), .X(n57432) );
  inv_x8_sg U74323 ( .A(n57444), .X(n57433) );
  inv_x8_sg U74324 ( .A(n57443), .X(n57434) );
  inv_x8_sg U74325 ( .A(n57442), .X(n57435) );
  inv_x8_sg U74326 ( .A(n57441), .X(n57436) );
  inv_x8_sg U74327 ( .A(n57440), .X(n57437) );
  inv_x8_sg U74328 ( .A(n57397), .X(n57438) );
  inv_x8_sg U74329 ( .A(n57447), .X(n57439) );
  inv_x8_sg U74330 ( .A(n57449), .X(n57440) );
  inv_x8_sg U74331 ( .A(n57449), .X(n57441) );
  inv_x8_sg U74332 ( .A(n57449), .X(n57442) );
  inv_x8_sg U74333 ( .A(n57449), .X(n57443) );
  inv_x8_sg U74334 ( .A(n57448), .X(n57444) );
  inv_x8_sg U74335 ( .A(n57448), .X(n57445) );
  inv_x8_sg U74336 ( .A(n57447), .X(n57446) );
  inv_x8_sg U74337 ( .A(n61858), .X(n57447) );
  inv_x8_sg U74338 ( .A(n61858), .X(n57448) );
  inv_x8_sg U74339 ( .A(n61858), .X(n57449) );
  inv_x8_sg U74340 ( .A(n68590), .X(n57450) );
  inv_x8_sg U74341 ( .A(n68591), .X(n57453) );
  inv_x8_sg U74342 ( .A(n57456), .X(n57454) );
  inv_x8_sg U74343 ( .A(n57456), .X(n57455) );
  inv_x8_sg U74344 ( .A(n57457), .X(n57456) );
  inv_x8_sg U74345 ( .A(n57460), .X(n57459) );
  inv_x8_sg U74346 ( .A(n57461), .X(n57460) );
  inv_x8_sg U74347 ( .A(n68587), .X(n57463) );
  inv_x8_sg U74348 ( .A(n57465), .X(n57464) );
  inv_x8_sg U74349 ( .A(n57469), .X(n57468) );
  inv_x8_sg U74350 ( .A(n57473), .X(n57472) );
  inv_x8_sg U74351 ( .A(n57477), .X(n57476) );
  inv_x8_sg U74352 ( .A(n57481), .X(n57480) );
  inv_x8_sg U74353 ( .A(n57485), .X(n57484) );
  inv_x8_sg U74354 ( .A(n57489), .X(n57488) );
  inv_x8_sg U74355 ( .A(n57493), .X(n57492) );
  inv_x8_sg U74356 ( .A(n57497), .X(n57496) );
  inv_x8_sg U74357 ( .A(n57500), .X(n57499) );
  inv_x8_sg U74358 ( .A(n57503), .X(n57502) );
  inv_x8_sg U74359 ( .A(n57508), .X(n57507) );
  inv_x8_sg U74360 ( .A(n57511), .X(n57510) );
  inv_x8_sg U74361 ( .A(n57514), .X(n57513) );
  inv_x8_sg U74362 ( .A(n57517), .X(n57516) );
  inv_x8_sg U74363 ( .A(n57528), .X(n57519) );
  inv_x8_sg U74364 ( .A(n57528), .X(n57520) );
  inv_x8_sg U74365 ( .A(n57528), .X(n57521) );
  inv_x8_sg U74366 ( .A(n57528), .X(n57522) );
  inv_x8_sg U74367 ( .A(n57528), .X(n57523) );
  inv_x8_sg U74368 ( .A(n57528), .X(n57524) );
  inv_x8_sg U74369 ( .A(n57528), .X(n57525) );
  inv_x8_sg U74370 ( .A(n57528), .X(n57526) );
  inv_x8_sg U74371 ( .A(n57528), .X(n57527) );
  inv_x8_sg U74372 ( .A(n57529), .X(n57528) );
  inv_x8_sg U74373 ( .A(n57549), .X(n57530) );
  inv_x8_sg U74374 ( .A(n57549), .X(n57531) );
  inv_x8_sg U74375 ( .A(n57549), .X(n57532) );
  inv_x8_sg U74376 ( .A(n57560), .X(n57533) );
  inv_x8_sg U74377 ( .A(n57560), .X(n57534) );
  inv_x8_sg U74378 ( .A(n57556), .X(n57535) );
  inv_x8_sg U74379 ( .A(n57556), .X(n57536) );
  inv_x8_sg U74380 ( .A(n57556), .X(n57537) );
  inv_x8_sg U74381 ( .A(n57556), .X(n57538) );
  inv_x8_sg U74382 ( .A(n57548), .X(n57539) );
  inv_x8_sg U74383 ( .A(n57548), .X(n57540) );
  inv_x8_sg U74384 ( .A(n57556), .X(n57541) );
  inv_x8_sg U74385 ( .A(n57548), .X(n57542) );
  inv_x8_sg U74386 ( .A(n57548), .X(n57543) );
  inv_x8_sg U74387 ( .A(n57548), .X(n57544) );
  inv_x8_sg U74388 ( .A(n57548), .X(n57545) );
  inv_x8_sg U74389 ( .A(n57549), .X(n57546) );
  inv_x8_sg U74390 ( .A(n57556), .X(n57547) );
  inv_x8_sg U74391 ( .A(n57553), .X(n57548) );
  inv_x8_sg U74392 ( .A(n57551), .X(n57549) );
  inv_x8_sg U74393 ( .A(n57560), .X(n57550) );
  inv_x8_sg U74394 ( .A(n57560), .X(n57551) );
  inv_x8_sg U74395 ( .A(n57556), .X(n57552) );
  inv_x8_sg U74396 ( .A(n57556), .X(n57553) );
  inv_x8_sg U74397 ( .A(n57555), .X(n57554) );
  inv_x8_sg U74398 ( .A(n57558), .X(n57556) );
  inv_x8_sg U74399 ( .A(n57560), .X(n57557) );
  inv_x8_sg U74400 ( .A(n57560), .X(n57558) );
  inv_x8_sg U74401 ( .A(n57561), .X(n57560) );
  inv_x8_sg U74402 ( .A(n57614), .X(n57562) );
  inv_x8_sg U74403 ( .A(n57626), .X(n57563) );
  inv_x8_sg U74404 ( .A(n57627), .X(n57564) );
  inv_x8_sg U74405 ( .A(n57626), .X(n57565) );
  inv_x8_sg U74406 ( .A(n57614), .X(n57566) );
  inv_x8_sg U74407 ( .A(n57614), .X(n57567) );
  inv_x8_sg U74408 ( .A(n57614), .X(n57568) );
  inv_x8_sg U74409 ( .A(n57614), .X(n57569) );
  inv_x8_sg U74410 ( .A(n57613), .X(n57570) );
  inv_x8_sg U74411 ( .A(n57613), .X(n57571) );
  inv_x8_sg U74412 ( .A(n57613), .X(n57572) );
  inv_x8_sg U74413 ( .A(n57613), .X(n57573) );
  inv_x8_sg U74414 ( .A(n57612), .X(n57574) );
  inv_x8_sg U74415 ( .A(n57612), .X(n57575) );
  inv_x8_sg U74416 ( .A(n57612), .X(n57576) );
  inv_x8_sg U74417 ( .A(n57611), .X(n57577) );
  inv_x8_sg U74418 ( .A(n57611), .X(n57578) );
  inv_x8_sg U74419 ( .A(n57611), .X(n57579) );
  inv_x8_sg U74420 ( .A(n57610), .X(n57580) );
  inv_x8_sg U74421 ( .A(n57610), .X(n57581) );
  inv_x8_sg U74422 ( .A(n57610), .X(n57582) );
  inv_x8_sg U74423 ( .A(n57610), .X(n57583) );
  inv_x8_sg U74424 ( .A(n57609), .X(n57584) );
  inv_x8_sg U74425 ( .A(n57609), .X(n57585) );
  inv_x8_sg U74426 ( .A(n57609), .X(n57586) );
  inv_x8_sg U74427 ( .A(n57609), .X(n57587) );
  inv_x8_sg U74428 ( .A(n57608), .X(n57588) );
  inv_x8_sg U74429 ( .A(n57608), .X(n57589) );
  inv_x8_sg U74430 ( .A(n57608), .X(n57590) );
  inv_x8_sg U74431 ( .A(n57608), .X(n57591) );
  inv_x8_sg U74432 ( .A(n57613), .X(n57592) );
  inv_x8_sg U74433 ( .A(n57610), .X(n57593) );
  inv_x8_sg U74434 ( .A(n57612), .X(n57594) );
  inv_x8_sg U74435 ( .A(n57611), .X(n57595) );
  inv_x8_sg U74436 ( .A(n57610), .X(n57596) );
  inv_x8_sg U74437 ( .A(n57608), .X(n57597) );
  inv_x8_sg U74438 ( .A(n57614), .X(n57598) );
  inv_x8_sg U74439 ( .A(n57608), .X(n57599) );
  inv_x8_sg U74440 ( .A(n57631), .X(n57600) );
  inv_x8_sg U74441 ( .A(n57607), .X(n57601) );
  inv_x8_sg U74442 ( .A(n57607), .X(n57602) );
  inv_x8_sg U74443 ( .A(n57607), .X(n57603) );
  inv_x8_sg U74444 ( .A(n57607), .X(n57604) );
  inv_x8_sg U74445 ( .A(n57607), .X(n57605) );
  inv_x8_sg U74446 ( .A(n57607), .X(n57606) );
  inv_x8_sg U74447 ( .A(n57625), .X(n57607) );
  inv_x8_sg U74448 ( .A(n57621), .X(n57608) );
  inv_x8_sg U74449 ( .A(n57620), .X(n57609) );
  inv_x8_sg U74450 ( .A(n57619), .X(n57610) );
  inv_x8_sg U74451 ( .A(n57618), .X(n57611) );
  inv_x8_sg U74452 ( .A(n57617), .X(n57612) );
  inv_x8_sg U74453 ( .A(n57616), .X(n57613) );
  inv_x8_sg U74454 ( .A(n57628), .X(n57614) );
  inv_x8_sg U74455 ( .A(n57631), .X(n57615) );
  inv_x8_sg U74456 ( .A(n57627), .X(n57616) );
  inv_x8_sg U74457 ( .A(n57627), .X(n57617) );
  inv_x8_sg U74458 ( .A(n57627), .X(n57618) );
  inv_x8_sg U74459 ( .A(n57627), .X(n57619) );
  inv_x8_sg U74460 ( .A(n57626), .X(n57620) );
  inv_x8_sg U74461 ( .A(n57626), .X(n57621) );
  inv_x8_sg U74462 ( .A(n57626), .X(n57622) );
  inv_x8_sg U74463 ( .A(n57626), .X(n57623) );
  inv_x8_sg U74464 ( .A(n57631), .X(n57624) );
  inv_x8_sg U74465 ( .A(n57631), .X(n57625) );
  inv_x8_sg U74466 ( .A(n57630), .X(n57626) );
  inv_x8_sg U74467 ( .A(n57629), .X(n57627) );
  inv_x8_sg U74468 ( .A(n57631), .X(n57628) );
  inv_x8_sg U74469 ( .A(n57631), .X(n57629) );
  inv_x8_sg U74470 ( .A(n57631), .X(n57630) );
  inv_x8_sg U74471 ( .A(n57632), .X(n57631) );
  inv_x8_sg U74472 ( .A(n57633), .X(n57632) );
  inv_x8_sg U74473 ( .A(n57719), .X(n57634) );
  inv_x8_sg U74474 ( .A(n57692), .X(n57635) );
  inv_x8_sg U74475 ( .A(n57692), .X(n57636) );
  inv_x8_sg U74476 ( .A(n57692), .X(n57637) );
  inv_x8_sg U74477 ( .A(n57692), .X(n57638) );
  inv_x8_sg U74478 ( .A(n57691), .X(n57639) );
  inv_x8_sg U74479 ( .A(n57691), .X(n57640) );
  inv_x8_sg U74480 ( .A(n57691), .X(n57641) );
  inv_x8_sg U74481 ( .A(n57690), .X(n57642) );
  inv_x8_sg U74482 ( .A(n57692), .X(n57643) );
  inv_x8_sg U74483 ( .A(n57690), .X(n57644) );
  inv_x8_sg U74484 ( .A(n57690), .X(n57645) );
  inv_x8_sg U74485 ( .A(n57690), .X(n57646) );
  inv_x8_sg U74486 ( .A(n57690), .X(n57647) );
  inv_x8_sg U74487 ( .A(n57689), .X(n57648) );
  inv_x8_sg U74488 ( .A(n57689), .X(n57649) );
  inv_x8_sg U74489 ( .A(n57689), .X(n57650) );
  inv_x8_sg U74490 ( .A(n57689), .X(n57651) );
  inv_x8_sg U74491 ( .A(n57688), .X(n57652) );
  inv_x8_sg U74492 ( .A(n57688), .X(n57653) );
  inv_x8_sg U74493 ( .A(n57688), .X(n57654) );
  inv_x8_sg U74494 ( .A(n57688), .X(n57655) );
  inv_x8_sg U74495 ( .A(n57687), .X(n57656) );
  inv_x8_sg U74496 ( .A(n57687), .X(n57657) );
  inv_x8_sg U74497 ( .A(n57687), .X(n57658) );
  inv_x8_sg U74498 ( .A(n57687), .X(n57659) );
  inv_x8_sg U74499 ( .A(n57686), .X(n57660) );
  inv_x8_sg U74500 ( .A(n57686), .X(n57661) );
  inv_x8_sg U74501 ( .A(n57686), .X(n57662) );
  inv_x8_sg U74502 ( .A(n57686), .X(n57663) );
  inv_x8_sg U74503 ( .A(n57685), .X(n57664) );
  inv_x8_sg U74504 ( .A(n57685), .X(n57665) );
  inv_x8_sg U74505 ( .A(n57685), .X(n57666) );
  inv_x8_sg U74506 ( .A(n57685), .X(n57667) );
  inv_x8_sg U74507 ( .A(n57684), .X(n57668) );
  inv_x8_sg U74508 ( .A(n57684), .X(n57669) );
  inv_x8_sg U74509 ( .A(n57684), .X(n57670) );
  inv_x8_sg U74510 ( .A(n57684), .X(n57671) );
  inv_x8_sg U74511 ( .A(n57711), .X(n57672) );
  inv_x8_sg U74512 ( .A(n57713), .X(n57673) );
  inv_x8_sg U74513 ( .A(n57683), .X(n57674) );
  inv_x8_sg U74514 ( .A(n57683), .X(n57675) );
  inv_x8_sg U74515 ( .A(n57710), .X(n57676) );
  inv_x8_sg U74516 ( .A(n57683), .X(n57677) );
  inv_x8_sg U74517 ( .A(n57713), .X(n57678) );
  inv_x8_sg U74518 ( .A(n57683), .X(n57679) );
  inv_x8_sg U74519 ( .A(n57719), .X(n57680) );
  inv_x8_sg U74520 ( .A(n57719), .X(n57681) );
  inv_x8_sg U74521 ( .A(n57721), .X(n57682) );
  inv_x8_sg U74522 ( .A(n57705), .X(n57683) );
  inv_x8_sg U74523 ( .A(n57702), .X(n57684) );
  inv_x8_sg U74524 ( .A(n57701), .X(n57685) );
  inv_x8_sg U74525 ( .A(n57700), .X(n57686) );
  inv_x8_sg U74526 ( .A(n57699), .X(n57687) );
  inv_x8_sg U74527 ( .A(n57698), .X(n57688) );
  inv_x8_sg U74528 ( .A(n57697), .X(n57689) );
  inv_x8_sg U74529 ( .A(n57696), .X(n57690) );
  inv_x8_sg U74530 ( .A(n57694), .X(n57691) );
  inv_x8_sg U74531 ( .A(n57693), .X(n57692) );
  inv_x8_sg U74532 ( .A(n57713), .X(n57693) );
  inv_x8_sg U74533 ( .A(n57713), .X(n57694) );
  inv_x8_sg U74534 ( .A(n57713), .X(n57695) );
  inv_x8_sg U74535 ( .A(n57713), .X(n57696) );
  inv_x8_sg U74536 ( .A(n57712), .X(n57697) );
  inv_x8_sg U74537 ( .A(n57712), .X(n57698) );
  inv_x8_sg U74538 ( .A(n57711), .X(n57699) );
  inv_x8_sg U74539 ( .A(n57711), .X(n57700) );
  inv_x8_sg U74540 ( .A(n57712), .X(n57701) );
  inv_x8_sg U74541 ( .A(n57711), .X(n57702) );
  inv_x8_sg U74542 ( .A(n57712), .X(n57703) );
  inv_x8_sg U74543 ( .A(n57710), .X(n57704) );
  inv_x8_sg U74544 ( .A(n57710), .X(n57705) );
  inv_x8_sg U74545 ( .A(n57710), .X(n57706) );
  inv_x8_sg U74546 ( .A(n57710), .X(n57707) );
  inv_x8_sg U74547 ( .A(n57719), .X(n57708) );
  inv_x8_sg U74548 ( .A(n57719), .X(n57709) );
  inv_x8_sg U74549 ( .A(n57718), .X(n57710) );
  inv_x8_sg U74550 ( .A(n57716), .X(n57711) );
  inv_x8_sg U74551 ( .A(n57716), .X(n57712) );
  inv_x8_sg U74552 ( .A(n57715), .X(n57713) );
  inv_x8_sg U74553 ( .A(n57719), .X(n57715) );
  inv_x8_sg U74554 ( .A(n57719), .X(n57716) );
  inv_x8_sg U74555 ( .A(n57719), .X(n57717) );
  inv_x8_sg U74556 ( .A(n57719), .X(n57718) );
  inv_x8_sg U74557 ( .A(n57720), .X(n57719) );
  inv_x8_sg U74558 ( .A(n57721), .X(n57720) );
  inv_x8_sg U74559 ( .A(n57722), .X(n57721) );
  inv_x8_sg U74560 ( .A(n57753), .X(n57724) );
  inv_x8_sg U74561 ( .A(n57753), .X(n57725) );
  inv_x8_sg U74562 ( .A(n57753), .X(n57726) );
  inv_x8_sg U74563 ( .A(n57753), .X(n57727) );
  inv_x8_sg U74564 ( .A(n57769), .X(n57728) );
  inv_x8_sg U74565 ( .A(n57752), .X(n57729) );
  inv_x8_sg U74566 ( .A(n57752), .X(n57730) );
  inv_x8_sg U74567 ( .A(n57752), .X(n57731) );
  inv_x8_sg U74568 ( .A(n57752), .X(n57732) );
  inv_x8_sg U74569 ( .A(n57753), .X(n57733) );
  inv_x8_sg U74570 ( .A(n57751), .X(n57734) );
  inv_x8_sg U74571 ( .A(n57751), .X(n57735) );
  inv_x8_sg U74572 ( .A(n57751), .X(n57736) );
  inv_x8_sg U74573 ( .A(n57753), .X(n57737) );
  inv_x8_sg U74574 ( .A(n57752), .X(n57738) );
  inv_x8_sg U74575 ( .A(n57753), .X(n57739) );
  inv_x8_sg U74576 ( .A(n57751), .X(n57740) );
  inv_x8_sg U74577 ( .A(n57751), .X(n57741) );
  inv_x8_sg U74578 ( .A(n57767), .X(n57742) );
  inv_x8_sg U74579 ( .A(n57774), .X(n57743) );
  inv_x8_sg U74580 ( .A(n57767), .X(n57744) );
  inv_x8_sg U74581 ( .A(n57751), .X(n57745) );
  inv_x8_sg U74582 ( .A(n57767), .X(n57746) );
  inv_x8_sg U74583 ( .A(n57768), .X(n57747) );
  inv_x8_sg U74584 ( .A(n57767), .X(n57748) );
  inv_x8_sg U74585 ( .A(n57768), .X(n57749) );
  inv_x8_sg U74586 ( .A(n57767), .X(n57750) );
  inv_x8_sg U74587 ( .A(n57760), .X(n57751) );
  inv_x8_sg U74588 ( .A(n57758), .X(n57752) );
  inv_x8_sg U74589 ( .A(n57754), .X(n57753) );
  inv_x8_sg U74590 ( .A(n57769), .X(n57754) );
  inv_x8_sg U74591 ( .A(n57769), .X(n57755) );
  inv_x8_sg U74592 ( .A(n57769), .X(n57756) );
  inv_x8_sg U74593 ( .A(n57769), .X(n57757) );
  inv_x8_sg U74594 ( .A(n57768), .X(n57758) );
  inv_x8_sg U74595 ( .A(n57768), .X(n57759) );
  inv_x8_sg U74596 ( .A(n57768), .X(n57760) );
  inv_x8_sg U74597 ( .A(n57768), .X(n57761) );
  inv_x8_sg U74598 ( .A(n57767), .X(n57762) );
  inv_x8_sg U74599 ( .A(n57774), .X(n57763) );
  inv_x8_sg U74600 ( .A(n57768), .X(n57764) );
  inv_x8_sg U74601 ( .A(n57767), .X(n57765) );
  inv_x8_sg U74602 ( .A(n57767), .X(n57766) );
  inv_x8_sg U74603 ( .A(n57773), .X(n57767) );
  inv_x8_sg U74604 ( .A(n57771), .X(n57768) );
  inv_x8_sg U74605 ( .A(n57770), .X(n57769) );
  inv_x8_sg U74606 ( .A(n57774), .X(n57770) );
  inv_x8_sg U74607 ( .A(n57774), .X(n57771) );
  inv_x8_sg U74608 ( .A(n57774), .X(n57772) );
  inv_x8_sg U74609 ( .A(n57774), .X(n57773) );
  inv_x8_sg U74610 ( .A(n57775), .X(n57774) );
  inv_x8_sg U74611 ( .A(n57776), .X(n57775) );
  inv_x8_sg U74612 ( .A(n57781), .X(n57779) );
  inv_x8_sg U74613 ( .A(n57781), .X(n57780) );
  inv_x8_sg U74614 ( .A(n47573), .X(n57781) );
  inv_x8_sg U74615 ( .A(n57783), .X(n57782) );
  inv_x8_sg U74616 ( .A(n57787), .X(n57786) );
  inv_x8_sg U74617 ( .A(n57792), .X(n57788) );
  inv_x8_sg U74618 ( .A(n57792), .X(n57789) );
  inv_x8_sg U74619 ( .A(n57792), .X(n57790) );
  inv_x8_sg U74620 ( .A(n57792), .X(n57791) );
  inv_x8_sg U74621 ( .A(n57793), .X(n57792) );
  inv_x8_sg U74622 ( .A(n57828), .X(n57795) );
  inv_x8_sg U74623 ( .A(n57835), .X(n57796) );
  inv_x8_sg U74624 ( .A(n57834), .X(n57797) );
  inv_x8_sg U74625 ( .A(n57834), .X(n57798) );
  inv_x8_sg U74626 ( .A(n57833), .X(n57799) );
  inv_x8_sg U74627 ( .A(n57833), .X(n57800) );
  inv_x8_sg U74628 ( .A(n57833), .X(n57801) );
  inv_x8_sg U74629 ( .A(n57833), .X(n57802) );
  inv_x8_sg U74630 ( .A(n57833), .X(n57803) );
  inv_x8_sg U74631 ( .A(n57835), .X(n57804) );
  inv_x8_sg U74632 ( .A(n57835), .X(n57805) );
  inv_x8_sg U74633 ( .A(n57832), .X(n57806) );
  inv_x8_sg U74634 ( .A(n57832), .X(n57807) );
  inv_x8_sg U74635 ( .A(n57832), .X(n57808) );
  inv_x8_sg U74636 ( .A(n57832), .X(n57809) );
  inv_x8_sg U74637 ( .A(n57831), .X(n57810) );
  inv_x8_sg U74638 ( .A(n57831), .X(n57811) );
  inv_x8_sg U74639 ( .A(n57831), .X(n57812) );
  inv_x8_sg U74640 ( .A(n57831), .X(n57813) );
  inv_x8_sg U74641 ( .A(n57830), .X(n57814) );
  inv_x8_sg U74642 ( .A(n57830), .X(n57815) );
  inv_x8_sg U74643 ( .A(n57830), .X(n57816) );
  inv_x8_sg U74644 ( .A(n57830), .X(n57817) );
  inv_x8_sg U74645 ( .A(n57831), .X(n57818) );
  inv_x8_sg U74646 ( .A(n57831), .X(n57819) );
  inv_x8_sg U74647 ( .A(n57834), .X(n57820) );
  inv_x8_sg U74648 ( .A(n57829), .X(n57821) );
  inv_x8_sg U74649 ( .A(n57828), .X(n57822) );
  inv_x8_sg U74650 ( .A(n57828), .X(n57823) );
  inv_x8_sg U74651 ( .A(n57851), .X(n57824) );
  inv_x8_sg U74652 ( .A(n57848), .X(n57825) );
  inv_x8_sg U74653 ( .A(n57848), .X(n57826) );
  inv_x8_sg U74654 ( .A(n57848), .X(n57827) );
  inv_x8_sg U74655 ( .A(n57845), .X(n57828) );
  inv_x8_sg U74656 ( .A(n57842), .X(n57830) );
  inv_x8_sg U74657 ( .A(n57841), .X(n57831) );
  inv_x8_sg U74658 ( .A(n57840), .X(n57832) );
  inv_x8_sg U74659 ( .A(n57838), .X(n57833) );
  inv_x8_sg U74660 ( .A(n57837), .X(n57834) );
  inv_x8_sg U74661 ( .A(n57836), .X(n57835) );
  inv_x8_sg U74662 ( .A(n57848), .X(n57836) );
  inv_x8_sg U74663 ( .A(n57848), .X(n57837) );
  inv_x8_sg U74664 ( .A(n57848), .X(n57838) );
  inv_x8_sg U74665 ( .A(n57848), .X(n57839) );
  inv_x8_sg U74666 ( .A(n57847), .X(n57840) );
  inv_x8_sg U74667 ( .A(n57847), .X(n57841) );
  inv_x8_sg U74668 ( .A(n57847), .X(n57842) );
  inv_x8_sg U74669 ( .A(n57847), .X(n57843) );
  inv_x8_sg U74670 ( .A(n57851), .X(n57844) );
  inv_x8_sg U74671 ( .A(n57851), .X(n57845) );
  inv_x8_sg U74672 ( .A(n57851), .X(n57846) );
  inv_x8_sg U74673 ( .A(n57850), .X(n57847) );
  inv_x8_sg U74674 ( .A(n57849), .X(n57848) );
  inv_x8_sg U74675 ( .A(n57851), .X(n57849) );
  inv_x8_sg U74676 ( .A(n57851), .X(n57850) );
  inv_x8_sg U74677 ( .A(n46203), .X(n57851) );
  inv_x8_sg U74678 ( .A(n57856), .X(n57854) );
  inv_x8_sg U74679 ( .A(n57856), .X(n57855) );
  inv_x8_sg U74680 ( .A(n32874), .X(n57856) );
  inv_x8_sg U74681 ( .A(n57102), .X(n57857) );
  inv_x8_sg U74682 ( .A(n57859), .X(n57858) );
  inv_x8_sg U74683 ( .A(n57860), .X(n57859) );
  inv_x8_sg U74684 ( .A(n57861), .X(n57860) );
  inv_x8_sg U74685 ( .A(n57863), .X(n57862) );
  inv_x8_sg U74686 ( .A(n68589), .X(n57864) );
  inv_x8_sg U74687 ( .A(n57866), .X(n57865) );
  inv_x8_sg U74688 ( .A(n57874), .X(n57870) );
  inv_x8_sg U74689 ( .A(n57874), .X(n57871) );
  inv_x8_sg U74690 ( .A(n57874), .X(n57872) );
  inv_x8_sg U74691 ( .A(n57874), .X(n57873) );
  inv_x8_sg U74692 ( .A(n57876), .X(n57874) );
  inv_x8_sg U74693 ( .A(n57881), .X(n57875) );
  inv_x8_sg U74694 ( .A(n57881), .X(n57876) );
  inv_x8_sg U74695 ( .A(n57881), .X(n57877) );
  inv_x8_sg U74696 ( .A(n57881), .X(n57878) );
  inv_x8_sg U74697 ( .A(n57881), .X(n57880) );
  inv_x8_sg U74698 ( .A(n57882), .X(n57881) );
  inv_x8_sg U74699 ( .A(n57883), .X(n57882) );
  inv_x8_sg U74700 ( .A(n57912), .X(n57886) );
  inv_x8_sg U74701 ( .A(n57912), .X(n57887) );
  inv_x8_sg U74702 ( .A(n57905), .X(n57888) );
  inv_x8_sg U74703 ( .A(n57906), .X(n57889) );
  inv_x8_sg U74704 ( .A(n57906), .X(n57890) );
  inv_x8_sg U74705 ( .A(n57906), .X(n57891) );
  inv_x8_sg U74706 ( .A(n57906), .X(n57892) );
  inv_x8_sg U74707 ( .A(n57906), .X(n57893) );
  inv_x8_sg U74708 ( .A(n57906), .X(n57894) );
  inv_x8_sg U74709 ( .A(n57912), .X(n57895) );
  inv_x8_sg U74710 ( .A(n57912), .X(n57896) );
  inv_x8_sg U74711 ( .A(n57905), .X(n57897) );
  inv_x8_sg U74712 ( .A(n57912), .X(n57898) );
  inv_x8_sg U74713 ( .A(n57912), .X(n57899) );
  inv_x8_sg U74714 ( .A(n57912), .X(n57900) );
  inv_x8_sg U74715 ( .A(n57905), .X(n57901) );
  inv_x8_sg U74716 ( .A(n57905), .X(n57902) );
  inv_x8_sg U74717 ( .A(n57905), .X(n57903) );
  inv_x8_sg U74718 ( .A(n57905), .X(n57904) );
  inv_x8_sg U74719 ( .A(n57899), .X(n57905) );
  inv_x8_sg U74720 ( .A(n57909), .X(n57906) );
  inv_x8_sg U74721 ( .A(n57912), .X(n57907) );
  inv_x8_sg U74722 ( .A(n57912), .X(n57908) );
  inv_x8_sg U74723 ( .A(n57912), .X(n57909) );
  inv_x8_sg U74724 ( .A(n57912), .X(n57910) );
  inv_x8_sg U74725 ( .A(n57912), .X(n57911) );
  inv_x8_sg U74726 ( .A(n46206), .X(n57912) );
  inv_x8_sg U74727 ( .A(n57919), .X(n57917) );
  inv_x8_sg U74728 ( .A(n57920), .X(n57918) );
  inv_x8_sg U74729 ( .A(n57920), .X(n57919) );
  inv_x8_sg U74730 ( .A(n57921), .X(n57920) );
  inv_x8_sg U74731 ( .A(n57925), .X(n57922) );
  inv_x8_sg U74732 ( .A(n57925), .X(n57923) );
  inv_x8_sg U74733 ( .A(n57925), .X(n57924) );
  inv_x8_sg U74734 ( .A(n53717), .X(n57925) );
  inv_x4_sg U74735 ( .A(n57950), .X(n57926) );
  inv_x4_sg U74736 ( .A(n57950), .X(n57927) );
  inv_x4_sg U74737 ( .A(n57946), .X(n57928) );
  inv_x4_sg U74738 ( .A(n57946), .X(n57929) );
  inv_x4_sg U74739 ( .A(n57949), .X(n57930) );
  inv_x4_sg U74740 ( .A(n57949), .X(n57931) );
  inv_x4_sg U74741 ( .A(n57949), .X(n57932) );
  inv_x4_sg U74742 ( .A(n57949), .X(n57933) );
  inv_x4_sg U74743 ( .A(n57949), .X(n57934) );
  inv_x4_sg U74744 ( .A(n57949), .X(n57935) );
  inv_x4_sg U74745 ( .A(n57949), .X(n57936) );
  inv_x4_sg U74746 ( .A(n57949), .X(n57937) );
  inv_x4_sg U74747 ( .A(n57949), .X(n57938) );
  inv_x4_sg U74748 ( .A(n57949), .X(n57939) );
  inv_x4_sg U74749 ( .A(n57949), .X(n57940) );
  inv_x4_sg U74750 ( .A(n57949), .X(n57941) );
  inv_x4_sg U74751 ( .A(n57949), .X(n57942) );
  inv_x4_sg U74752 ( .A(n57949), .X(n57943) );
  inv_x4_sg U74753 ( .A(n57949), .X(n57944) );
  inv_x4_sg U74754 ( .A(n57949), .X(n57945) );
  inv_x4_sg U74755 ( .A(n57951), .X(n57946) );
  inv_x4_sg U74756 ( .A(n57949), .X(n57948) );
  inv_x8_sg U74757 ( .A(n57951), .X(n57949) );
  inv_x8_sg U74758 ( .A(n57951), .X(n57950) );
  inv_x8_sg U74759 ( .A(n57952), .X(n57951) );
  inv_x4_sg U74760 ( .A(n46891), .X(n57952) );
  inv_x2_sg U74761 ( .A(n57953), .X(n61906) );
  nand_x8_sg U74762 ( .A(n57954), .B(n61908), .X(n30624) );
  nand_x8_sg U74763 ( .A(n58616), .B(n57296), .X(n58657) );
  nand_x8_sg U74764 ( .A(n57325), .B(n57917), .X(n58630) );
  nor_x2_sg U74765 ( .A(n58630), .B(n57956), .X(n57964) );
  nand_x8_sg U74766 ( .A(n47317), .B(n61905), .X(n61858) );
  inv_x2_sg U74767 ( .A(n32484), .X(n57968) );
  nand_x8_sg U74768 ( .A(n47615), .B(n57968), .X(n58612) );
  nand_x8_sg U74769 ( .A(n57927), .B(n57925), .X(n58639) );
  nand_x8_sg U74770 ( .A(n57923), .B(n57950), .X(n58640) );
  nor_x2_sg U74771 ( .A(n57330), .B(n68571), .X(n57984) );
  nand_x8_sg U74772 ( .A(n22467), .B(n57984), .X(n26003) );
  nand_x8_sg U74773 ( .A(n57949), .B(n57925), .X(n58638) );
  nand_x8_sg U74774 ( .A(n57326), .B(n57454), .X(n24829) );
  nand_x8_sg U74775 ( .A(n57455), .B(n57925), .X(n58125) );
  inv_x2_sg U74776 ( .A(n55311), .X(n57991) );
  inv_x2_sg U74777 ( .A(n55309), .X(n57995) );
  inv_x2_sg U74778 ( .A(n55295), .X(n58008) );
  inv_x2_sg U74779 ( .A(n55293), .X(n58012) );
  inv_x2_sg U74780 ( .A(n55291), .X(n58022) );
  inv_x2_sg U74781 ( .A(n55289), .X(n58026) );
  inv_x2_sg U74782 ( .A(n55287), .X(n58039) );
  inv_x2_sg U74783 ( .A(n55285), .X(n58043) );
  inv_x2_sg U74784 ( .A(n55315), .X(n58061) );
  inv_x2_sg U74785 ( .A(n55313), .X(n58065) );
  inv_x2_sg U74786 ( .A(n55307), .X(n58078) );
  inv_x2_sg U74787 ( .A(n55305), .X(n58082) );
  inv_x2_sg U74788 ( .A(n55303), .X(n58092) );
  inv_x2_sg U74789 ( .A(n55301), .X(n58096) );
  inv_x2_sg U74790 ( .A(n55299), .X(n58109) );
  inv_x2_sg U74791 ( .A(n55297), .X(n58113) );
  inv_x2_sg U74792 ( .A(n58127), .X(n58132) );
  inv_x2_sg U74793 ( .A(n58140), .X(n58141) );
  inv_x2_sg U74794 ( .A(n58145), .X(n58146) );
  inv_x2_sg U74795 ( .A(n58165), .X(n58166) );
  inv_x2_sg U74796 ( .A(n58170), .X(n58171) );
  inv_x2_sg U74797 ( .A(n58185), .X(n58186) );
  inv_x2_sg U74798 ( .A(n58190), .X(n58191) );
  inv_x2_sg U74799 ( .A(n58210), .X(n58211) );
  inv_x2_sg U74800 ( .A(n58215), .X(n58216) );
  inv_x2_sg U74801 ( .A(n58240), .X(n58241) );
  inv_x2_sg U74802 ( .A(n58245), .X(n58246) );
  inv_x2_sg U74803 ( .A(n58265), .X(n58266) );
  inv_x2_sg U74804 ( .A(n58270), .X(n58271) );
  inv_x2_sg U74805 ( .A(n58285), .X(n58286) );
  inv_x2_sg U74806 ( .A(n58290), .X(n58291) );
  inv_x2_sg U74807 ( .A(n58310), .X(n58311) );
  inv_x2_sg U74808 ( .A(n58315), .X(n58316) );
  nor_x2_sg U74809 ( .A(n57460), .B(n58377), .X(n58381) );
  inv_x2_sg U74810 ( .A(n58378), .X(n58379) );
  nand_x8_sg U74811 ( .A(n58381), .B(n58380), .X(n23671) );
  nor_x2_sg U74812 ( .A(n57462), .B(n58382), .X(n58386) );
  inv_x2_sg U74813 ( .A(n58383), .X(n58384) );
  nand_x8_sg U74814 ( .A(n58386), .B(n58385), .X(n23539) );
  nand_x8_sg U74815 ( .A(n57326), .B(n57296), .X(n68591) );
  nand_x8_sg U74816 ( .A(n57349), .B(n57296), .X(n68590) );
  nand_x8_sg U74817 ( .A(n58478), .B(n57296), .X(n58656) );
  inv_x2_sg U74818 ( .A(n23415), .X(n58430) );
  inv_x2_sg U74819 ( .A(n23307), .X(n58472) );
  nand_x8_sg U74820 ( .A(n57327), .B(n58479), .X(n68588) );
  nand_x8_sg U74821 ( .A(n58479), .B(n58478), .X(n68589) );
  nand_x8_sg U74822 ( .A(n57450), .B(n57917), .X(n68587) );
  nand_x8_sg U74823 ( .A(n58581), .B(n57343), .X(n58585) );
  inv_x2_sg U74824 ( .A(n58585), .X(n58482) );
  inv_x2_sg U74825 ( .A(n58583), .X(n22443) );
  inv_x2_sg U74826 ( .A(n58586), .X(n22418) );
  nor_x2_sg U74827 ( .A(n57343), .B(n22445), .X(n58587) );
  nand_x8_sg U74828 ( .A(n29338), .B(n58587), .X(n22395) );
  inv_x2_sg U74829 ( .A(n32533), .X(n58588) );
  inv_x2_sg U74830 ( .A(n32433), .X(n58599) );
  nor_x2_sg U74831 ( .A(n32415), .B(n57103), .X(n32579) );
  nor_x2_sg U74832 ( .A(n32411), .B(n58639), .X(n32580) );
  nor_x2_sg U74833 ( .A(n32405), .B(n58640), .X(n58604) );
  nor_x2_sg U74834 ( .A(n32401), .B(n57099), .X(n58603) );
  inv_x2_sg U74835 ( .A(n32499), .X(n58609) );
  nor_x2_sg U74836 ( .A(n32403), .B(n58656), .X(n58621) );
  nor_x2_sg U74837 ( .A(n32399), .B(n58657), .X(n58620) );
  inv_x2_sg U74838 ( .A(n32088), .X(n58622) );
  inv_x2_sg U74839 ( .A(n31966), .X(n58634) );
  nor_x2_sg U74840 ( .A(n31947), .B(n57104), .X(n32134) );
  nor_x2_sg U74841 ( .A(n31943), .B(n58639), .X(n32135) );
  nor_x2_sg U74842 ( .A(n31937), .B(n58640), .X(n58642) );
  nor_x2_sg U74843 ( .A(n31933), .B(n57099), .X(n58641) );
  inv_x2_sg U74844 ( .A(n32056), .X(n58648) );
  nor_x2_sg U74845 ( .A(n31935), .B(n58656), .X(n58659) );
  nor_x2_sg U74846 ( .A(n31931), .B(n58657), .X(n58658) );
  nand_x8_sg U74847 ( .A(n57430), .B(n61905), .X(n61856) );
  inv_x2_sg U74848 ( .A(ow_15[0]), .X(n58660) );
  inv_x2_sg U74849 ( .A(ow_15[1]), .X(n58665) );
  inv_x2_sg U74850 ( .A(ow_15[2]), .X(n58670) );
  inv_x2_sg U74851 ( .A(ow_15[3]), .X(n58675) );
  inv_x2_sg U74852 ( .A(ow_15[4]), .X(n58680) );
  inv_x2_sg U74853 ( .A(ow_15[5]), .X(n58685) );
  inv_x2_sg U74854 ( .A(ow_15[6]), .X(n58690) );
  inv_x2_sg U74855 ( .A(ow_15[7]), .X(n58695) );
  inv_x2_sg U74856 ( .A(ow_15[8]), .X(n58700) );
  inv_x2_sg U74857 ( .A(ow_15[9]), .X(n58705) );
  inv_x2_sg U74858 ( .A(ow_15[10]), .X(n58710) );
  inv_x2_sg U74859 ( .A(ow_15[11]), .X(n58715) );
  inv_x2_sg U74860 ( .A(ow_15[12]), .X(n58720) );
  inv_x2_sg U74861 ( .A(ow_15[13]), .X(n58725) );
  inv_x2_sg U74862 ( .A(ow_15[14]), .X(n58730) );
  inv_x2_sg U74863 ( .A(ow_15[15]), .X(n58735) );
  inv_x2_sg U74864 ( .A(ow_15[16]), .X(n58740) );
  inv_x2_sg U74865 ( .A(ow_15[17]), .X(n58745) );
  inv_x2_sg U74866 ( .A(ow_15[18]), .X(n58750) );
  inv_x2_sg U74867 ( .A(ow_15[19]), .X(n58755) );
  inv_x2_sg U74868 ( .A(ow_14[0]), .X(n58760) );
  inv_x2_sg U74869 ( .A(ow_14[1]), .X(n58765) );
  inv_x2_sg U74870 ( .A(ow_14[2]), .X(n58770) );
  inv_x2_sg U74871 ( .A(ow_14[3]), .X(n58775) );
  inv_x2_sg U74872 ( .A(ow_14[4]), .X(n58780) );
  inv_x2_sg U74873 ( .A(ow_14[5]), .X(n58785) );
  inv_x2_sg U74874 ( .A(ow_14[6]), .X(n58790) );
  inv_x2_sg U74875 ( .A(ow_14[7]), .X(n58795) );
  inv_x2_sg U74876 ( .A(ow_14[8]), .X(n58800) );
  inv_x2_sg U74877 ( .A(ow_14[9]), .X(n58805) );
  inv_x2_sg U74878 ( .A(ow_14[10]), .X(n58810) );
  inv_x2_sg U74879 ( .A(ow_14[11]), .X(n58815) );
  inv_x2_sg U74880 ( .A(ow_14[12]), .X(n58820) );
  inv_x2_sg U74881 ( .A(ow_14[13]), .X(n58825) );
  inv_x2_sg U74882 ( .A(ow_14[14]), .X(n58830) );
  inv_x2_sg U74883 ( .A(ow_14[15]), .X(n58835) );
  inv_x2_sg U74884 ( .A(ow_14[16]), .X(n58840) );
  inv_x2_sg U74885 ( .A(ow_14[17]), .X(n58845) );
  inv_x2_sg U74886 ( .A(ow_14[18]), .X(n58850) );
  inv_x2_sg U74887 ( .A(ow_14[19]), .X(n58855) );
  inv_x2_sg U74888 ( .A(ow_13[0]), .X(n58860) );
  inv_x2_sg U74889 ( .A(ow_13[1]), .X(n58865) );
  inv_x2_sg U74890 ( .A(ow_13[2]), .X(n58870) );
  inv_x2_sg U74891 ( .A(ow_13[3]), .X(n58875) );
  inv_x2_sg U74892 ( .A(ow_13[4]), .X(n58880) );
  inv_x2_sg U74893 ( .A(ow_13[5]), .X(n58885) );
  inv_x2_sg U74894 ( .A(ow_13[6]), .X(n58890) );
  inv_x2_sg U74895 ( .A(ow_13[7]), .X(n58895) );
  inv_x2_sg U74896 ( .A(ow_13[8]), .X(n58900) );
  inv_x2_sg U74897 ( .A(ow_13[9]), .X(n58905) );
  inv_x2_sg U74898 ( .A(ow_13[10]), .X(n58910) );
  inv_x2_sg U74899 ( .A(ow_13[11]), .X(n58915) );
  inv_x2_sg U74900 ( .A(ow_13[12]), .X(n58920) );
  inv_x2_sg U74901 ( .A(ow_13[13]), .X(n58925) );
  inv_x2_sg U74902 ( .A(ow_13[14]), .X(n58930) );
  inv_x2_sg U74903 ( .A(ow_13[15]), .X(n58935) );
  inv_x2_sg U74904 ( .A(ow_13[16]), .X(n58940) );
  inv_x2_sg U74905 ( .A(ow_13[17]), .X(n58945) );
  inv_x2_sg U74906 ( .A(ow_13[18]), .X(n58950) );
  inv_x2_sg U74907 ( .A(ow_13[19]), .X(n58955) );
  inv_x2_sg U74908 ( .A(ow_12[0]), .X(n58960) );
  inv_x2_sg U74909 ( .A(ow_12[1]), .X(n58965) );
  inv_x2_sg U74910 ( .A(ow_12[2]), .X(n58970) );
  inv_x2_sg U74911 ( .A(ow_12[3]), .X(n58975) );
  inv_x2_sg U74912 ( .A(ow_12[4]), .X(n58980) );
  inv_x2_sg U74913 ( .A(ow_12[5]), .X(n58985) );
  inv_x2_sg U74914 ( .A(ow_12[6]), .X(n58990) );
  inv_x2_sg U74915 ( .A(ow_12[7]), .X(n58995) );
  inv_x2_sg U74916 ( .A(ow_12[8]), .X(n59000) );
  inv_x2_sg U74917 ( .A(ow_12[9]), .X(n59005) );
  inv_x2_sg U74918 ( .A(ow_12[10]), .X(n59010) );
  inv_x2_sg U74919 ( .A(ow_12[11]), .X(n59015) );
  inv_x2_sg U74920 ( .A(ow_12[12]), .X(n59020) );
  inv_x2_sg U74921 ( .A(ow_12[13]), .X(n59025) );
  inv_x2_sg U74922 ( .A(ow_12[14]), .X(n59030) );
  inv_x2_sg U74923 ( .A(ow_12[15]), .X(n59035) );
  inv_x2_sg U74924 ( .A(ow_12[16]), .X(n59040) );
  inv_x2_sg U74925 ( .A(ow_12[17]), .X(n59045) );
  inv_x2_sg U74926 ( .A(ow_12[18]), .X(n59050) );
  inv_x2_sg U74927 ( .A(ow_12[19]), .X(n59055) );
  inv_x2_sg U74928 ( .A(ow_11[0]), .X(n59060) );
  inv_x2_sg U74929 ( .A(ow_11[1]), .X(n59065) );
  inv_x2_sg U74930 ( .A(ow_11[2]), .X(n59070) );
  inv_x2_sg U74931 ( .A(ow_11[3]), .X(n59075) );
  inv_x2_sg U74932 ( .A(ow_11[4]), .X(n59080) );
  inv_x2_sg U74933 ( .A(ow_11[5]), .X(n59085) );
  inv_x2_sg U74934 ( .A(ow_11[6]), .X(n59090) );
  inv_x2_sg U74935 ( .A(ow_11[7]), .X(n59095) );
  inv_x2_sg U74936 ( .A(ow_11[8]), .X(n59100) );
  inv_x2_sg U74937 ( .A(ow_11[9]), .X(n59105) );
  inv_x2_sg U74938 ( .A(ow_11[10]), .X(n59110) );
  inv_x2_sg U74939 ( .A(ow_11[11]), .X(n59115) );
  inv_x2_sg U74940 ( .A(ow_11[12]), .X(n59120) );
  inv_x2_sg U74941 ( .A(ow_11[13]), .X(n59125) );
  inv_x2_sg U74942 ( .A(ow_11[14]), .X(n59130) );
  inv_x2_sg U74943 ( .A(ow_11[15]), .X(n59135) );
  inv_x2_sg U74944 ( .A(ow_11[16]), .X(n59140) );
  inv_x2_sg U74945 ( .A(ow_11[17]), .X(n59145) );
  inv_x2_sg U74946 ( .A(ow_11[18]), .X(n59150) );
  inv_x2_sg U74947 ( .A(ow_11[19]), .X(n59155) );
  inv_x2_sg U74948 ( .A(ow_10[0]), .X(n59160) );
  inv_x2_sg U74949 ( .A(ow_10[1]), .X(n59165) );
  inv_x2_sg U74950 ( .A(ow_10[2]), .X(n59170) );
  inv_x2_sg U74951 ( .A(ow_10[3]), .X(n59175) );
  inv_x2_sg U74952 ( .A(ow_10[4]), .X(n59180) );
  inv_x2_sg U74953 ( .A(ow_10[5]), .X(n59185) );
  inv_x2_sg U74954 ( .A(ow_10[6]), .X(n59190) );
  inv_x2_sg U74955 ( .A(ow_10[7]), .X(n59195) );
  inv_x2_sg U74956 ( .A(ow_10[8]), .X(n59200) );
  inv_x2_sg U74957 ( .A(ow_10[9]), .X(n59205) );
  inv_x2_sg U74958 ( .A(ow_10[10]), .X(n59210) );
  inv_x2_sg U74959 ( .A(ow_10[11]), .X(n59215) );
  inv_x2_sg U74960 ( .A(ow_10[12]), .X(n59220) );
  inv_x2_sg U74961 ( .A(ow_10[13]), .X(n59225) );
  inv_x2_sg U74962 ( .A(ow_10[14]), .X(n59230) );
  inv_x2_sg U74963 ( .A(ow_10[15]), .X(n59235) );
  inv_x2_sg U74964 ( .A(ow_10[16]), .X(n59240) );
  inv_x2_sg U74965 ( .A(ow_10[17]), .X(n59245) );
  inv_x2_sg U74966 ( .A(ow_10[18]), .X(n59250) );
  inv_x2_sg U74967 ( .A(ow_10[19]), .X(n59255) );
  inv_x2_sg U74968 ( .A(ow_9[0]), .X(n59260) );
  inv_x2_sg U74969 ( .A(ow_9[1]), .X(n59265) );
  inv_x2_sg U74970 ( .A(ow_9[2]), .X(n59270) );
  inv_x2_sg U74971 ( .A(ow_9[3]), .X(n59275) );
  inv_x2_sg U74972 ( .A(ow_9[4]), .X(n59280) );
  inv_x2_sg U74973 ( .A(ow_9[5]), .X(n59285) );
  inv_x2_sg U74974 ( .A(ow_9[6]), .X(n59290) );
  inv_x2_sg U74975 ( .A(ow_9[7]), .X(n59295) );
  inv_x2_sg U74976 ( .A(ow_9[8]), .X(n59300) );
  inv_x2_sg U74977 ( .A(ow_9[9]), .X(n59305) );
  inv_x2_sg U74978 ( .A(ow_9[10]), .X(n59310) );
  inv_x2_sg U74979 ( .A(ow_9[11]), .X(n59315) );
  inv_x2_sg U74980 ( .A(ow_9[12]), .X(n59320) );
  inv_x2_sg U74981 ( .A(ow_9[13]), .X(n59325) );
  inv_x2_sg U74982 ( .A(ow_9[14]), .X(n59330) );
  inv_x2_sg U74983 ( .A(ow_9[15]), .X(n59335) );
  inv_x2_sg U74984 ( .A(ow_9[16]), .X(n59340) );
  inv_x2_sg U74985 ( .A(ow_9[17]), .X(n59345) );
  inv_x2_sg U74986 ( .A(ow_9[18]), .X(n59350) );
  inv_x2_sg U74987 ( .A(ow_9[19]), .X(n59355) );
  inv_x2_sg U74988 ( .A(ow_8[0]), .X(n59360) );
  inv_x2_sg U74989 ( .A(ow_8[1]), .X(n59365) );
  inv_x2_sg U74990 ( .A(ow_8[2]), .X(n59370) );
  inv_x2_sg U74991 ( .A(ow_8[3]), .X(n59375) );
  inv_x2_sg U74992 ( .A(ow_8[4]), .X(n59380) );
  inv_x2_sg U74993 ( .A(ow_8[5]), .X(n59385) );
  inv_x2_sg U74994 ( .A(ow_8[6]), .X(n59390) );
  inv_x2_sg U74995 ( .A(ow_8[7]), .X(n59395) );
  inv_x2_sg U74996 ( .A(ow_8[8]), .X(n59400) );
  inv_x2_sg U74997 ( .A(ow_8[9]), .X(n59405) );
  inv_x2_sg U74998 ( .A(ow_8[10]), .X(n59410) );
  inv_x2_sg U74999 ( .A(ow_8[11]), .X(n59415) );
  inv_x2_sg U75000 ( .A(ow_8[12]), .X(n59420) );
  inv_x2_sg U75001 ( .A(ow_8[13]), .X(n59425) );
  inv_x2_sg U75002 ( .A(ow_8[14]), .X(n59430) );
  inv_x2_sg U75003 ( .A(ow_8[15]), .X(n59435) );
  inv_x2_sg U75004 ( .A(ow_8[16]), .X(n59440) );
  inv_x2_sg U75005 ( .A(ow_8[17]), .X(n59445) );
  inv_x2_sg U75006 ( .A(ow_8[18]), .X(n59450) );
  inv_x2_sg U75007 ( .A(ow_8[19]), .X(n59455) );
  inv_x2_sg U75008 ( .A(ow_7[0]), .X(n59460) );
  inv_x2_sg U75009 ( .A(ow_7[1]), .X(n59465) );
  inv_x2_sg U75010 ( .A(ow_7[2]), .X(n59470) );
  inv_x2_sg U75011 ( .A(ow_7[3]), .X(n59475) );
  inv_x2_sg U75012 ( .A(ow_7[4]), .X(n59480) );
  inv_x2_sg U75013 ( .A(ow_7[5]), .X(n59485) );
  inv_x2_sg U75014 ( .A(ow_7[6]), .X(n59490) );
  inv_x2_sg U75015 ( .A(ow_7[7]), .X(n59495) );
  inv_x2_sg U75016 ( .A(ow_7[8]), .X(n59500) );
  inv_x2_sg U75017 ( .A(ow_7[9]), .X(n59505) );
  inv_x2_sg U75018 ( .A(ow_7[10]), .X(n59510) );
  inv_x2_sg U75019 ( .A(ow_7[11]), .X(n59515) );
  inv_x2_sg U75020 ( .A(ow_7[12]), .X(n59520) );
  inv_x2_sg U75021 ( .A(ow_7[13]), .X(n59525) );
  inv_x2_sg U75022 ( .A(ow_7[14]), .X(n59530) );
  inv_x2_sg U75023 ( .A(ow_7[15]), .X(n59535) );
  inv_x2_sg U75024 ( .A(ow_7[16]), .X(n59540) );
  inv_x2_sg U75025 ( .A(ow_7[17]), .X(n59545) );
  inv_x2_sg U75026 ( .A(ow_7[18]), .X(n59550) );
  inv_x2_sg U75027 ( .A(ow_7[19]), .X(n59555) );
  inv_x2_sg U75028 ( .A(ow_6[0]), .X(n59560) );
  inv_x2_sg U75029 ( .A(ow_6[1]), .X(n59565) );
  inv_x2_sg U75030 ( .A(ow_6[2]), .X(n59570) );
  inv_x2_sg U75031 ( .A(ow_6[3]), .X(n59575) );
  inv_x2_sg U75032 ( .A(ow_6[4]), .X(n59580) );
  inv_x2_sg U75033 ( .A(ow_6[5]), .X(n59585) );
  inv_x2_sg U75034 ( .A(ow_6[6]), .X(n59590) );
  inv_x2_sg U75035 ( .A(ow_6[7]), .X(n59595) );
  inv_x2_sg U75036 ( .A(ow_6[8]), .X(n59600) );
  inv_x2_sg U75037 ( .A(ow_6[9]), .X(n59605) );
  inv_x2_sg U75038 ( .A(ow_6[10]), .X(n59610) );
  inv_x2_sg U75039 ( .A(ow_6[11]), .X(n59615) );
  inv_x2_sg U75040 ( .A(ow_6[12]), .X(n59620) );
  inv_x2_sg U75041 ( .A(ow_6[13]), .X(n59625) );
  inv_x2_sg U75042 ( .A(ow_6[14]), .X(n59630) );
  inv_x2_sg U75043 ( .A(ow_6[15]), .X(n59635) );
  inv_x2_sg U75044 ( .A(ow_6[16]), .X(n59640) );
  inv_x2_sg U75045 ( .A(ow_6[17]), .X(n59645) );
  inv_x2_sg U75046 ( .A(ow_6[18]), .X(n59650) );
  inv_x2_sg U75047 ( .A(ow_6[19]), .X(n59655) );
  inv_x2_sg U75048 ( .A(ow_5[0]), .X(n59660) );
  inv_x2_sg U75049 ( .A(ow_5[1]), .X(n59665) );
  inv_x2_sg U75050 ( .A(ow_5[2]), .X(n59670) );
  inv_x2_sg U75051 ( .A(ow_5[3]), .X(n59675) );
  inv_x2_sg U75052 ( .A(ow_5[4]), .X(n59680) );
  inv_x2_sg U75053 ( .A(ow_5[5]), .X(n59685) );
  inv_x2_sg U75054 ( .A(ow_5[6]), .X(n59690) );
  inv_x2_sg U75055 ( .A(ow_5[7]), .X(n59695) );
  inv_x2_sg U75056 ( .A(ow_5[8]), .X(n59700) );
  inv_x2_sg U75057 ( .A(ow_5[9]), .X(n59705) );
  inv_x2_sg U75058 ( .A(ow_5[10]), .X(n59710) );
  inv_x2_sg U75059 ( .A(ow_5[11]), .X(n59715) );
  inv_x2_sg U75060 ( .A(ow_5[12]), .X(n59720) );
  inv_x2_sg U75061 ( .A(ow_5[13]), .X(n59725) );
  inv_x2_sg U75062 ( .A(ow_5[14]), .X(n59730) );
  inv_x2_sg U75063 ( .A(ow_5[15]), .X(n59735) );
  inv_x2_sg U75064 ( .A(ow_5[16]), .X(n59740) );
  inv_x2_sg U75065 ( .A(ow_5[17]), .X(n59745) );
  inv_x2_sg U75066 ( .A(ow_5[18]), .X(n59750) );
  inv_x2_sg U75067 ( .A(ow_5[19]), .X(n59755) );
  inv_x2_sg U75068 ( .A(ow_4[0]), .X(n59760) );
  inv_x2_sg U75069 ( .A(ow_4[1]), .X(n59765) );
  inv_x2_sg U75070 ( .A(ow_4[2]), .X(n59770) );
  inv_x2_sg U75071 ( .A(ow_4[3]), .X(n59775) );
  inv_x2_sg U75072 ( .A(ow_4[4]), .X(n59780) );
  inv_x2_sg U75073 ( .A(ow_4[5]), .X(n59785) );
  inv_x2_sg U75074 ( .A(ow_4[6]), .X(n59790) );
  inv_x2_sg U75075 ( .A(ow_4[7]), .X(n59795) );
  inv_x2_sg U75076 ( .A(ow_4[8]), .X(n59800) );
  inv_x2_sg U75077 ( .A(ow_4[9]), .X(n59805) );
  inv_x2_sg U75078 ( .A(ow_4[10]), .X(n59810) );
  inv_x2_sg U75079 ( .A(ow_4[11]), .X(n59815) );
  inv_x2_sg U75080 ( .A(ow_4[12]), .X(n59820) );
  inv_x2_sg U75081 ( .A(ow_4[13]), .X(n59825) );
  inv_x2_sg U75082 ( .A(ow_4[14]), .X(n59830) );
  inv_x2_sg U75083 ( .A(ow_4[15]), .X(n59835) );
  inv_x2_sg U75084 ( .A(ow_4[16]), .X(n59840) );
  inv_x2_sg U75085 ( .A(ow_4[17]), .X(n59845) );
  inv_x2_sg U75086 ( .A(ow_4[18]), .X(n59850) );
  inv_x2_sg U75087 ( .A(ow_4[19]), .X(n59855) );
  inv_x2_sg U75088 ( .A(ow_3[0]), .X(n59860) );
  inv_x2_sg U75089 ( .A(ow_3[1]), .X(n59865) );
  inv_x2_sg U75090 ( .A(ow_3[2]), .X(n59870) );
  inv_x2_sg U75091 ( .A(ow_3[3]), .X(n59875) );
  inv_x2_sg U75092 ( .A(ow_3[4]), .X(n59880) );
  inv_x2_sg U75093 ( .A(ow_3[5]), .X(n59885) );
  inv_x2_sg U75094 ( .A(ow_3[6]), .X(n59890) );
  inv_x2_sg U75095 ( .A(ow_3[7]), .X(n59895) );
  inv_x2_sg U75096 ( .A(ow_3[8]), .X(n59900) );
  inv_x2_sg U75097 ( .A(ow_3[9]), .X(n59905) );
  inv_x2_sg U75098 ( .A(ow_3[10]), .X(n59910) );
  inv_x2_sg U75099 ( .A(ow_3[11]), .X(n59915) );
  inv_x2_sg U75100 ( .A(ow_3[12]), .X(n59920) );
  inv_x2_sg U75101 ( .A(ow_3[13]), .X(n59925) );
  inv_x2_sg U75102 ( .A(ow_3[14]), .X(n59930) );
  inv_x2_sg U75103 ( .A(ow_3[15]), .X(n59935) );
  inv_x2_sg U75104 ( .A(ow_3[16]), .X(n59940) );
  inv_x2_sg U75105 ( .A(ow_3[17]), .X(n59945) );
  inv_x2_sg U75106 ( .A(ow_3[18]), .X(n59950) );
  inv_x2_sg U75107 ( .A(ow_3[19]), .X(n59955) );
  inv_x2_sg U75108 ( .A(ow_2[0]), .X(n59960) );
  inv_x2_sg U75109 ( .A(ow_2[1]), .X(n59965) );
  inv_x2_sg U75110 ( .A(ow_2[2]), .X(n59970) );
  inv_x2_sg U75111 ( .A(ow_2[3]), .X(n59975) );
  inv_x2_sg U75112 ( .A(ow_2[4]), .X(n59980) );
  inv_x2_sg U75113 ( .A(ow_2[5]), .X(n59985) );
  inv_x2_sg U75114 ( .A(ow_2[6]), .X(n59990) );
  inv_x2_sg U75115 ( .A(ow_2[7]), .X(n59995) );
  inv_x2_sg U75116 ( .A(ow_2[8]), .X(n60000) );
  inv_x2_sg U75117 ( .A(ow_2[9]), .X(n60005) );
  inv_x2_sg U75118 ( .A(ow_2[10]), .X(n60010) );
  inv_x2_sg U75119 ( .A(ow_2[11]), .X(n60015) );
  inv_x2_sg U75120 ( .A(ow_2[12]), .X(n60020) );
  inv_x2_sg U75121 ( .A(ow_2[13]), .X(n60025) );
  inv_x2_sg U75122 ( .A(ow_2[14]), .X(n60030) );
  inv_x2_sg U75123 ( .A(ow_2[15]), .X(n60035) );
  inv_x2_sg U75124 ( .A(ow_2[16]), .X(n60040) );
  inv_x2_sg U75125 ( .A(ow_2[17]), .X(n60045) );
  inv_x2_sg U75126 ( .A(ow_2[18]), .X(n60050) );
  inv_x2_sg U75127 ( .A(ow_2[19]), .X(n60055) );
  inv_x2_sg U75128 ( .A(ow_1[0]), .X(n60060) );
  inv_x2_sg U75129 ( .A(ow_1[1]), .X(n60065) );
  inv_x2_sg U75130 ( .A(ow_1[2]), .X(n60070) );
  inv_x2_sg U75131 ( .A(ow_1[3]), .X(n60075) );
  inv_x2_sg U75132 ( .A(ow_1[4]), .X(n60080) );
  inv_x2_sg U75133 ( .A(ow_1[5]), .X(n60085) );
  inv_x2_sg U75134 ( .A(ow_1[6]), .X(n60090) );
  inv_x2_sg U75135 ( .A(ow_1[7]), .X(n60095) );
  inv_x2_sg U75136 ( .A(ow_1[8]), .X(n60100) );
  inv_x2_sg U75137 ( .A(ow_1[9]), .X(n60105) );
  inv_x2_sg U75138 ( .A(ow_1[10]), .X(n60110) );
  inv_x2_sg U75139 ( .A(ow_1[11]), .X(n60115) );
  inv_x2_sg U75140 ( .A(ow_1[12]), .X(n60120) );
  inv_x2_sg U75141 ( .A(ow_1[13]), .X(n60125) );
  inv_x2_sg U75142 ( .A(ow_1[14]), .X(n60130) );
  inv_x2_sg U75143 ( .A(ow_1[15]), .X(n60135) );
  inv_x2_sg U75144 ( .A(ow_1[16]), .X(n60140) );
  inv_x2_sg U75145 ( .A(ow_1[17]), .X(n60145) );
  inv_x2_sg U75146 ( .A(ow_1[18]), .X(n60150) );
  inv_x2_sg U75147 ( .A(ow_1[19]), .X(n60155) );
  inv_x2_sg U75148 ( .A(ow_0[0]), .X(n60160) );
  inv_x2_sg U75149 ( .A(ow_0[1]), .X(n60165) );
  inv_x2_sg U75150 ( .A(ow_0[2]), .X(n60170) );
  inv_x2_sg U75151 ( .A(ow_0[3]), .X(n60175) );
  inv_x2_sg U75152 ( .A(ow_0[4]), .X(n60180) );
  inv_x2_sg U75153 ( .A(ow_0[5]), .X(n60185) );
  inv_x2_sg U75154 ( .A(ow_0[6]), .X(n60190) );
  inv_x2_sg U75155 ( .A(ow_0[7]), .X(n60195) );
  inv_x2_sg U75156 ( .A(ow_0[8]), .X(n60200) );
  inv_x2_sg U75157 ( .A(ow_0[9]), .X(n60205) );
  inv_x2_sg U75158 ( .A(ow_0[10]), .X(n60210) );
  inv_x2_sg U75159 ( .A(ow_0[11]), .X(n60215) );
  inv_x2_sg U75160 ( .A(ow_0[12]), .X(n60220) );
  inv_x2_sg U75161 ( .A(ow_0[13]), .X(n60225) );
  inv_x2_sg U75162 ( .A(ow_0[14]), .X(n60230) );
  inv_x2_sg U75163 ( .A(ow_0[15]), .X(n60235) );
  inv_x2_sg U75164 ( .A(ow_0[16]), .X(n60240) );
  inv_x2_sg U75165 ( .A(ow_0[17]), .X(n60245) );
  inv_x2_sg U75166 ( .A(ow_0[18]), .X(n60250) );
  inv_x2_sg U75167 ( .A(ow_0[19]), .X(n60255) );
  inv_x2_sg U75168 ( .A(oi_15[0]), .X(n60260) );
  inv_x2_sg U75169 ( .A(oi_15[1]), .X(n60265) );
  inv_x2_sg U75170 ( .A(oi_15[2]), .X(n60270) );
  inv_x2_sg U75171 ( .A(oi_15[3]), .X(n60275) );
  inv_x2_sg U75172 ( .A(oi_15[4]), .X(n60280) );
  inv_x2_sg U75173 ( .A(oi_15[5]), .X(n60285) );
  inv_x2_sg U75174 ( .A(oi_15[6]), .X(n60290) );
  inv_x2_sg U75175 ( .A(oi_15[7]), .X(n60295) );
  inv_x2_sg U75176 ( .A(oi_15[8]), .X(n60300) );
  inv_x2_sg U75177 ( .A(oi_15[9]), .X(n60305) );
  inv_x2_sg U75178 ( .A(oi_15[10]), .X(n60310) );
  inv_x2_sg U75179 ( .A(oi_15[11]), .X(n60315) );
  inv_x2_sg U75180 ( .A(oi_15[12]), .X(n60320) );
  inv_x2_sg U75181 ( .A(oi_15[13]), .X(n60325) );
  inv_x2_sg U75182 ( .A(oi_15[14]), .X(n60330) );
  inv_x2_sg U75183 ( .A(oi_15[15]), .X(n60335) );
  inv_x2_sg U75184 ( .A(oi_15[16]), .X(n60340) );
  inv_x2_sg U75185 ( .A(oi_15[17]), .X(n60345) );
  inv_x2_sg U75186 ( .A(oi_15[18]), .X(n60350) );
  inv_x2_sg U75187 ( .A(oi_15[19]), .X(n60355) );
  inv_x2_sg U75188 ( .A(oi_14[0]), .X(n60360) );
  inv_x2_sg U75189 ( .A(oi_14[1]), .X(n60365) );
  inv_x2_sg U75190 ( .A(oi_14[2]), .X(n60370) );
  inv_x2_sg U75191 ( .A(oi_14[3]), .X(n60375) );
  inv_x2_sg U75192 ( .A(oi_14[4]), .X(n60380) );
  inv_x2_sg U75193 ( .A(oi_14[5]), .X(n60385) );
  inv_x2_sg U75194 ( .A(oi_14[6]), .X(n60390) );
  inv_x2_sg U75195 ( .A(oi_14[7]), .X(n60395) );
  inv_x2_sg U75196 ( .A(oi_14[8]), .X(n60400) );
  inv_x2_sg U75197 ( .A(oi_14[9]), .X(n60405) );
  inv_x2_sg U75198 ( .A(oi_14[10]), .X(n60410) );
  inv_x2_sg U75199 ( .A(oi_14[11]), .X(n60415) );
  inv_x2_sg U75200 ( .A(oi_14[12]), .X(n60420) );
  inv_x2_sg U75201 ( .A(oi_14[13]), .X(n60425) );
  inv_x2_sg U75202 ( .A(oi_14[14]), .X(n60430) );
  inv_x2_sg U75203 ( .A(oi_14[15]), .X(n60435) );
  inv_x2_sg U75204 ( .A(oi_14[16]), .X(n60440) );
  inv_x2_sg U75205 ( .A(oi_14[17]), .X(n60445) );
  inv_x2_sg U75206 ( .A(oi_14[18]), .X(n60450) );
  inv_x2_sg U75207 ( .A(oi_14[19]), .X(n60455) );
  inv_x2_sg U75208 ( .A(oi_13[0]), .X(n60460) );
  inv_x2_sg U75209 ( .A(oi_13[1]), .X(n60465) );
  inv_x2_sg U75210 ( .A(oi_13[2]), .X(n60470) );
  inv_x2_sg U75211 ( .A(oi_13[3]), .X(n60475) );
  inv_x2_sg U75212 ( .A(oi_13[4]), .X(n60480) );
  inv_x2_sg U75213 ( .A(oi_13[5]), .X(n60485) );
  inv_x2_sg U75214 ( .A(oi_13[6]), .X(n60490) );
  inv_x2_sg U75215 ( .A(oi_13[7]), .X(n60495) );
  inv_x2_sg U75216 ( .A(oi_13[8]), .X(n60500) );
  inv_x2_sg U75217 ( .A(oi_13[9]), .X(n60505) );
  inv_x2_sg U75218 ( .A(oi_13[10]), .X(n60510) );
  inv_x2_sg U75219 ( .A(oi_13[11]), .X(n60515) );
  inv_x2_sg U75220 ( .A(oi_13[12]), .X(n60520) );
  inv_x2_sg U75221 ( .A(oi_13[13]), .X(n60525) );
  inv_x2_sg U75222 ( .A(oi_13[14]), .X(n60530) );
  inv_x2_sg U75223 ( .A(oi_13[15]), .X(n60535) );
  inv_x2_sg U75224 ( .A(oi_13[16]), .X(n60540) );
  inv_x2_sg U75225 ( .A(oi_13[17]), .X(n60545) );
  inv_x2_sg U75226 ( .A(oi_13[18]), .X(n60550) );
  inv_x2_sg U75227 ( .A(oi_13[19]), .X(n60555) );
  inv_x2_sg U75228 ( .A(oi_12[0]), .X(n60560) );
  inv_x2_sg U75229 ( .A(oi_12[1]), .X(n60565) );
  inv_x2_sg U75230 ( .A(oi_12[2]), .X(n60570) );
  inv_x2_sg U75231 ( .A(oi_12[3]), .X(n60575) );
  inv_x2_sg U75232 ( .A(oi_12[4]), .X(n60580) );
  inv_x2_sg U75233 ( .A(oi_12[5]), .X(n60585) );
  inv_x2_sg U75234 ( .A(oi_12[6]), .X(n60590) );
  inv_x2_sg U75235 ( .A(oi_12[7]), .X(n60595) );
  inv_x2_sg U75236 ( .A(oi_12[8]), .X(n60600) );
  inv_x2_sg U75237 ( .A(oi_12[9]), .X(n60605) );
  inv_x2_sg U75238 ( .A(oi_12[10]), .X(n60610) );
  inv_x2_sg U75239 ( .A(oi_12[11]), .X(n60615) );
  inv_x2_sg U75240 ( .A(oi_12[12]), .X(n60620) );
  inv_x2_sg U75241 ( .A(oi_12[13]), .X(n60625) );
  inv_x2_sg U75242 ( .A(oi_12[14]), .X(n60630) );
  inv_x2_sg U75243 ( .A(oi_12[15]), .X(n60635) );
  inv_x2_sg U75244 ( .A(oi_12[16]), .X(n60640) );
  inv_x2_sg U75245 ( .A(oi_12[17]), .X(n60645) );
  inv_x2_sg U75246 ( .A(oi_12[18]), .X(n60650) );
  inv_x2_sg U75247 ( .A(oi_12[19]), .X(n60655) );
  inv_x2_sg U75248 ( .A(oi_11[0]), .X(n60660) );
  inv_x2_sg U75249 ( .A(oi_11[1]), .X(n60665) );
  inv_x2_sg U75250 ( .A(oi_11[2]), .X(n60670) );
  inv_x2_sg U75251 ( .A(oi_11[3]), .X(n60675) );
  inv_x2_sg U75252 ( .A(oi_11[4]), .X(n60680) );
  inv_x2_sg U75253 ( .A(oi_11[5]), .X(n60685) );
  inv_x2_sg U75254 ( .A(oi_11[6]), .X(n60690) );
  inv_x2_sg U75255 ( .A(oi_11[7]), .X(n60695) );
  inv_x2_sg U75256 ( .A(oi_11[8]), .X(n60700) );
  inv_x2_sg U75257 ( .A(oi_11[9]), .X(n60705) );
  inv_x2_sg U75258 ( .A(oi_11[10]), .X(n60710) );
  inv_x2_sg U75259 ( .A(oi_11[11]), .X(n60715) );
  inv_x2_sg U75260 ( .A(oi_11[12]), .X(n60720) );
  inv_x2_sg U75261 ( .A(oi_11[13]), .X(n60725) );
  inv_x2_sg U75262 ( .A(oi_11[14]), .X(n60730) );
  inv_x2_sg U75263 ( .A(oi_11[15]), .X(n60735) );
  inv_x2_sg U75264 ( .A(oi_11[16]), .X(n60740) );
  inv_x2_sg U75265 ( .A(oi_11[17]), .X(n60745) );
  inv_x2_sg U75266 ( .A(oi_11[18]), .X(n60750) );
  inv_x2_sg U75267 ( .A(oi_11[19]), .X(n60755) );
  inv_x2_sg U75268 ( .A(oi_10[0]), .X(n60760) );
  inv_x2_sg U75269 ( .A(oi_10[1]), .X(n60765) );
  inv_x2_sg U75270 ( .A(oi_10[2]), .X(n60770) );
  inv_x2_sg U75271 ( .A(oi_10[3]), .X(n60775) );
  inv_x2_sg U75272 ( .A(oi_10[4]), .X(n60780) );
  inv_x2_sg U75273 ( .A(oi_10[5]), .X(n60785) );
  inv_x2_sg U75274 ( .A(oi_10[6]), .X(n60790) );
  inv_x2_sg U75275 ( .A(oi_10[7]), .X(n60795) );
  inv_x2_sg U75276 ( .A(oi_10[8]), .X(n60800) );
  inv_x2_sg U75277 ( .A(oi_10[9]), .X(n60805) );
  inv_x2_sg U75278 ( .A(oi_10[10]), .X(n60810) );
  inv_x2_sg U75279 ( .A(oi_10[11]), .X(n60815) );
  inv_x2_sg U75280 ( .A(oi_10[12]), .X(n60820) );
  inv_x2_sg U75281 ( .A(oi_10[13]), .X(n60825) );
  inv_x2_sg U75282 ( .A(oi_10[14]), .X(n60830) );
  inv_x2_sg U75283 ( .A(oi_10[15]), .X(n60835) );
  inv_x2_sg U75284 ( .A(oi_10[16]), .X(n60840) );
  inv_x2_sg U75285 ( .A(oi_10[17]), .X(n60845) );
  inv_x2_sg U75286 ( .A(oi_10[18]), .X(n60850) );
  inv_x2_sg U75287 ( .A(oi_10[19]), .X(n60855) );
  inv_x2_sg U75288 ( .A(oi_9[0]), .X(n60860) );
  inv_x2_sg U75289 ( .A(oi_9[1]), .X(n60865) );
  inv_x2_sg U75290 ( .A(oi_9[2]), .X(n60870) );
  inv_x2_sg U75291 ( .A(oi_9[3]), .X(n60875) );
  inv_x2_sg U75292 ( .A(oi_9[4]), .X(n60880) );
  inv_x2_sg U75293 ( .A(oi_9[5]), .X(n60885) );
  inv_x2_sg U75294 ( .A(oi_9[6]), .X(n60890) );
  inv_x2_sg U75295 ( .A(oi_9[7]), .X(n60895) );
  inv_x2_sg U75296 ( .A(oi_9[8]), .X(n60900) );
  inv_x2_sg U75297 ( .A(oi_9[9]), .X(n60905) );
  inv_x2_sg U75298 ( .A(oi_9[10]), .X(n60910) );
  inv_x2_sg U75299 ( .A(oi_9[11]), .X(n60915) );
  inv_x2_sg U75300 ( .A(oi_9[12]), .X(n60920) );
  inv_x2_sg U75301 ( .A(oi_9[13]), .X(n60925) );
  inv_x2_sg U75302 ( .A(oi_9[14]), .X(n60930) );
  inv_x2_sg U75303 ( .A(oi_9[15]), .X(n60935) );
  inv_x2_sg U75304 ( .A(oi_9[16]), .X(n60940) );
  inv_x2_sg U75305 ( .A(oi_9[17]), .X(n60945) );
  inv_x2_sg U75306 ( .A(oi_9[18]), .X(n60950) );
  inv_x2_sg U75307 ( .A(oi_9[19]), .X(n60955) );
  inv_x2_sg U75308 ( .A(oi_8[0]), .X(n60960) );
  inv_x2_sg U75309 ( .A(oi_8[1]), .X(n60965) );
  inv_x2_sg U75310 ( .A(oi_8[2]), .X(n60970) );
  inv_x2_sg U75311 ( .A(oi_8[3]), .X(n60975) );
  inv_x2_sg U75312 ( .A(oi_8[4]), .X(n60980) );
  inv_x2_sg U75313 ( .A(oi_8[5]), .X(n60985) );
  inv_x2_sg U75314 ( .A(oi_8[6]), .X(n60990) );
  inv_x2_sg U75315 ( .A(oi_8[7]), .X(n60995) );
  inv_x2_sg U75316 ( .A(oi_8[8]), .X(n61000) );
  inv_x2_sg U75317 ( .A(oi_8[9]), .X(n61005) );
  inv_x2_sg U75318 ( .A(oi_8[10]), .X(n61010) );
  inv_x2_sg U75319 ( .A(oi_8[11]), .X(n61015) );
  inv_x2_sg U75320 ( .A(oi_8[12]), .X(n61020) );
  inv_x2_sg U75321 ( .A(oi_8[13]), .X(n61025) );
  inv_x2_sg U75322 ( .A(oi_8[14]), .X(n61030) );
  inv_x2_sg U75323 ( .A(oi_8[15]), .X(n61035) );
  inv_x2_sg U75324 ( .A(oi_8[16]), .X(n61040) );
  inv_x2_sg U75325 ( .A(oi_8[17]), .X(n61045) );
  inv_x2_sg U75326 ( .A(oi_8[18]), .X(n61050) );
  inv_x2_sg U75327 ( .A(oi_8[19]), .X(n61055) );
  inv_x2_sg U75328 ( .A(oi_7[0]), .X(n61060) );
  inv_x2_sg U75329 ( .A(oi_7[1]), .X(n61065) );
  inv_x2_sg U75330 ( .A(oi_7[2]), .X(n61070) );
  inv_x2_sg U75331 ( .A(oi_7[3]), .X(n61075) );
  inv_x2_sg U75332 ( .A(oi_7[4]), .X(n61080) );
  inv_x2_sg U75333 ( .A(oi_7[5]), .X(n61085) );
  inv_x2_sg U75334 ( .A(oi_7[6]), .X(n61090) );
  inv_x2_sg U75335 ( .A(oi_7[7]), .X(n61095) );
  inv_x2_sg U75336 ( .A(oi_7[8]), .X(n61100) );
  inv_x2_sg U75337 ( .A(oi_7[9]), .X(n61105) );
  inv_x2_sg U75338 ( .A(oi_7[10]), .X(n61110) );
  inv_x2_sg U75339 ( .A(oi_7[11]), .X(n61115) );
  inv_x2_sg U75340 ( .A(oi_7[12]), .X(n61120) );
  inv_x2_sg U75341 ( .A(oi_7[13]), .X(n61125) );
  inv_x2_sg U75342 ( .A(oi_7[14]), .X(n61130) );
  inv_x2_sg U75343 ( .A(oi_7[15]), .X(n61135) );
  inv_x2_sg U75344 ( .A(oi_7[16]), .X(n61140) );
  inv_x2_sg U75345 ( .A(oi_7[17]), .X(n61145) );
  inv_x2_sg U75346 ( .A(oi_7[18]), .X(n61150) );
  inv_x2_sg U75347 ( .A(oi_7[19]), .X(n61155) );
  inv_x2_sg U75348 ( .A(oi_6[0]), .X(n61160) );
  inv_x2_sg U75349 ( .A(oi_6[1]), .X(n61165) );
  inv_x2_sg U75350 ( .A(oi_6[2]), .X(n61170) );
  inv_x2_sg U75351 ( .A(oi_6[3]), .X(n61175) );
  inv_x2_sg U75352 ( .A(oi_6[4]), .X(n61180) );
  inv_x2_sg U75353 ( .A(oi_6[5]), .X(n61185) );
  inv_x2_sg U75354 ( .A(oi_6[6]), .X(n61190) );
  inv_x2_sg U75355 ( .A(oi_6[7]), .X(n61195) );
  inv_x2_sg U75356 ( .A(oi_6[8]), .X(n61200) );
  inv_x2_sg U75357 ( .A(oi_6[9]), .X(n61205) );
  inv_x2_sg U75358 ( .A(oi_6[10]), .X(n61210) );
  inv_x2_sg U75359 ( .A(oi_6[11]), .X(n61215) );
  inv_x2_sg U75360 ( .A(oi_6[12]), .X(n61220) );
  inv_x2_sg U75361 ( .A(oi_6[13]), .X(n61225) );
  inv_x2_sg U75362 ( .A(oi_6[14]), .X(n61230) );
  inv_x2_sg U75363 ( .A(oi_6[15]), .X(n61235) );
  inv_x2_sg U75364 ( .A(oi_6[16]), .X(n61240) );
  inv_x2_sg U75365 ( .A(oi_6[17]), .X(n61245) );
  inv_x2_sg U75366 ( .A(oi_6[18]), .X(n61250) );
  inv_x2_sg U75367 ( .A(oi_6[19]), .X(n61255) );
  inv_x2_sg U75368 ( .A(oi_5[0]), .X(n61260) );
  inv_x2_sg U75369 ( .A(oi_5[1]), .X(n61265) );
  inv_x2_sg U75370 ( .A(oi_5[2]), .X(n61270) );
  inv_x2_sg U75371 ( .A(oi_5[3]), .X(n61275) );
  inv_x2_sg U75372 ( .A(oi_5[4]), .X(n61280) );
  inv_x2_sg U75373 ( .A(oi_5[5]), .X(n61285) );
  inv_x2_sg U75374 ( .A(oi_5[6]), .X(n61290) );
  inv_x2_sg U75375 ( .A(oi_5[7]), .X(n61295) );
  inv_x2_sg U75376 ( .A(oi_5[8]), .X(n61300) );
  inv_x2_sg U75377 ( .A(oi_5[9]), .X(n61305) );
  inv_x2_sg U75378 ( .A(oi_5[10]), .X(n61310) );
  inv_x2_sg U75379 ( .A(oi_5[11]), .X(n61315) );
  inv_x2_sg U75380 ( .A(oi_5[12]), .X(n61320) );
  inv_x2_sg U75381 ( .A(oi_5[13]), .X(n61325) );
  inv_x2_sg U75382 ( .A(oi_5[14]), .X(n61330) );
  inv_x2_sg U75383 ( .A(oi_5[15]), .X(n61335) );
  inv_x2_sg U75384 ( .A(oi_5[16]), .X(n61340) );
  inv_x2_sg U75385 ( .A(oi_5[17]), .X(n61345) );
  inv_x2_sg U75386 ( .A(oi_5[18]), .X(n61350) );
  inv_x2_sg U75387 ( .A(oi_5[19]), .X(n61355) );
  inv_x2_sg U75388 ( .A(oi_4[0]), .X(n61360) );
  inv_x2_sg U75389 ( .A(oi_4[1]), .X(n61365) );
  inv_x2_sg U75390 ( .A(oi_4[2]), .X(n61370) );
  inv_x2_sg U75391 ( .A(oi_4[3]), .X(n61375) );
  inv_x2_sg U75392 ( .A(oi_4[4]), .X(n61380) );
  inv_x2_sg U75393 ( .A(oi_4[5]), .X(n61385) );
  inv_x2_sg U75394 ( .A(oi_4[6]), .X(n61390) );
  inv_x2_sg U75395 ( .A(oi_4[7]), .X(n61395) );
  inv_x2_sg U75396 ( .A(oi_4[8]), .X(n61400) );
  inv_x2_sg U75397 ( .A(oi_4[9]), .X(n61405) );
  inv_x2_sg U75398 ( .A(oi_4[10]), .X(n61410) );
  inv_x2_sg U75399 ( .A(oi_4[11]), .X(n61415) );
  inv_x2_sg U75400 ( .A(oi_4[12]), .X(n61420) );
  inv_x2_sg U75401 ( .A(oi_4[13]), .X(n61425) );
  inv_x2_sg U75402 ( .A(oi_4[14]), .X(n61430) );
  inv_x2_sg U75403 ( .A(oi_4[15]), .X(n61435) );
  inv_x2_sg U75404 ( .A(oi_4[16]), .X(n61440) );
  inv_x2_sg U75405 ( .A(oi_4[17]), .X(n61445) );
  inv_x2_sg U75406 ( .A(oi_4[18]), .X(n61450) );
  inv_x2_sg U75407 ( .A(oi_4[19]), .X(n61455) );
  inv_x2_sg U75408 ( .A(oi_3[0]), .X(n61460) );
  inv_x2_sg U75409 ( .A(oi_3[1]), .X(n61465) );
  inv_x2_sg U75410 ( .A(oi_3[2]), .X(n61470) );
  inv_x2_sg U75411 ( .A(oi_3[3]), .X(n61475) );
  inv_x2_sg U75412 ( .A(oi_3[4]), .X(n61480) );
  inv_x2_sg U75413 ( .A(oi_3[5]), .X(n61485) );
  inv_x2_sg U75414 ( .A(oi_3[6]), .X(n61490) );
  inv_x2_sg U75415 ( .A(oi_3[7]), .X(n61495) );
  inv_x2_sg U75416 ( .A(oi_3[8]), .X(n61500) );
  inv_x2_sg U75417 ( .A(oi_3[9]), .X(n61505) );
  inv_x2_sg U75418 ( .A(oi_3[10]), .X(n61510) );
  inv_x2_sg U75419 ( .A(oi_3[11]), .X(n61515) );
  inv_x2_sg U75420 ( .A(oi_3[12]), .X(n61520) );
  inv_x2_sg U75421 ( .A(oi_3[13]), .X(n61525) );
  inv_x2_sg U75422 ( .A(oi_3[14]), .X(n61530) );
  inv_x2_sg U75423 ( .A(oi_3[15]), .X(n61535) );
  inv_x2_sg U75424 ( .A(oi_3[16]), .X(n61540) );
  inv_x2_sg U75425 ( .A(oi_3[17]), .X(n61545) );
  inv_x2_sg U75426 ( .A(oi_3[18]), .X(n61550) );
  inv_x2_sg U75427 ( .A(oi_3[19]), .X(n61555) );
  inv_x2_sg U75428 ( .A(oi_2[0]), .X(n61560) );
  inv_x2_sg U75429 ( .A(oi_2[1]), .X(n61565) );
  inv_x2_sg U75430 ( .A(oi_2[2]), .X(n61570) );
  inv_x2_sg U75431 ( .A(oi_2[3]), .X(n61575) );
  inv_x2_sg U75432 ( .A(oi_2[4]), .X(n61580) );
  inv_x2_sg U75433 ( .A(oi_2[5]), .X(n61585) );
  inv_x2_sg U75434 ( .A(oi_2[6]), .X(n61590) );
  inv_x2_sg U75435 ( .A(oi_2[7]), .X(n61595) );
  inv_x2_sg U75436 ( .A(oi_2[8]), .X(n61600) );
  inv_x2_sg U75437 ( .A(oi_2[9]), .X(n61605) );
  inv_x2_sg U75438 ( .A(oi_2[10]), .X(n61610) );
  inv_x2_sg U75439 ( .A(oi_2[11]), .X(n61615) );
  inv_x2_sg U75440 ( .A(oi_2[12]), .X(n61620) );
  inv_x2_sg U75441 ( .A(oi_2[13]), .X(n61625) );
  inv_x2_sg U75442 ( .A(oi_2[14]), .X(n61630) );
  inv_x2_sg U75443 ( .A(oi_2[15]), .X(n61635) );
  inv_x2_sg U75444 ( .A(oi_2[16]), .X(n61640) );
  inv_x2_sg U75445 ( .A(oi_2[17]), .X(n61645) );
  inv_x2_sg U75446 ( .A(oi_2[18]), .X(n61650) );
  inv_x2_sg U75447 ( .A(oi_2[19]), .X(n61655) );
  inv_x2_sg U75448 ( .A(oi_1[0]), .X(n61660) );
  inv_x2_sg U75449 ( .A(oi_1[1]), .X(n61665) );
  inv_x2_sg U75450 ( .A(oi_1[2]), .X(n61670) );
  inv_x2_sg U75451 ( .A(oi_1[3]), .X(n61675) );
  inv_x2_sg U75452 ( .A(oi_1[4]), .X(n61680) );
  inv_x2_sg U75453 ( .A(oi_1[5]), .X(n61685) );
  inv_x2_sg U75454 ( .A(oi_1[6]), .X(n61690) );
  inv_x2_sg U75455 ( .A(oi_1[7]), .X(n61695) );
  inv_x2_sg U75456 ( .A(oi_1[8]), .X(n61700) );
  inv_x2_sg U75457 ( .A(oi_1[9]), .X(n61705) );
  inv_x2_sg U75458 ( .A(oi_1[10]), .X(n61710) );
  inv_x2_sg U75459 ( .A(oi_1[11]), .X(n61715) );
  inv_x2_sg U75460 ( .A(oi_1[12]), .X(n61720) );
  inv_x2_sg U75461 ( .A(oi_1[13]), .X(n61725) );
  inv_x2_sg U75462 ( .A(oi_1[14]), .X(n61730) );
  inv_x2_sg U75463 ( .A(oi_1[15]), .X(n61735) );
  inv_x2_sg U75464 ( .A(oi_1[16]), .X(n61740) );
  inv_x2_sg U75465 ( .A(oi_1[17]), .X(n61745) );
  inv_x2_sg U75466 ( .A(oi_1[18]), .X(n61750) );
  inv_x2_sg U75467 ( .A(oi_1[19]), .X(n61755) );
  inv_x2_sg U75468 ( .A(oi_0[0]), .X(n61760) );
  inv_x2_sg U75469 ( .A(oi_0[1]), .X(n61765) );
  inv_x2_sg U75470 ( .A(oi_0[2]), .X(n61770) );
  inv_x2_sg U75471 ( .A(oi_0[3]), .X(n61775) );
  inv_x2_sg U75472 ( .A(oi_0[4]), .X(n61780) );
  inv_x2_sg U75473 ( .A(oi_0[5]), .X(n61785) );
  inv_x2_sg U75474 ( .A(oi_0[6]), .X(n61790) );
  inv_x2_sg U75475 ( .A(oi_0[7]), .X(n61795) );
  inv_x2_sg U75476 ( .A(oi_0[8]), .X(n61800) );
  inv_x2_sg U75477 ( .A(oi_0[9]), .X(n61805) );
  inv_x2_sg U75478 ( .A(oi_0[10]), .X(n61810) );
  inv_x2_sg U75479 ( .A(oi_0[11]), .X(n61815) );
  inv_x2_sg U75480 ( .A(oi_0[12]), .X(n61820) );
  inv_x2_sg U75481 ( .A(oi_0[13]), .X(n61825) );
  inv_x2_sg U75482 ( .A(oi_0[14]), .X(n61830) );
  inv_x2_sg U75483 ( .A(oi_0[15]), .X(n61835) );
  inv_x2_sg U75484 ( .A(oi_0[16]), .X(n61840) );
  inv_x2_sg U75485 ( .A(oi_0[17]), .X(n61845) );
  inv_x2_sg U75486 ( .A(oi_0[18]), .X(n61850) );
  inv_x2_sg U75487 ( .A(oi_0[19]), .X(n61855) );
  inv_x2_sg U80660 ( .A(n26162), .X(n67582) );
  inv_x2_sg U80661 ( .A(n26209), .X(n67543) );
  inv_x2_sg U80662 ( .A(n55069), .X(n67544) );
  inv_x2_sg U80663 ( .A(n26210), .X(n67540) );
  inv_x2_sg U80664 ( .A(n26243), .X(n67549) );
  inv_x2_sg U80665 ( .A(n55067), .X(n67550) );
  inv_x2_sg U80666 ( .A(n26244), .X(n67546) );
  inv_x2_sg U80667 ( .A(n26066), .X(n67576) );
  inv_x2_sg U80668 ( .A(n26112), .X(n67555) );
  inv_x2_sg U80669 ( .A(n55065), .X(n67556) );
  inv_x2_sg U80670 ( .A(n26115), .X(n67552) );
  inv_x2_sg U80671 ( .A(n26151), .X(n67561) );
  inv_x2_sg U80672 ( .A(n55063), .X(n67562) );
  inv_x2_sg U80673 ( .A(n26152), .X(n67558) );
  inv_x2_sg U80674 ( .A(n56595), .X(n67587) );
  inv_x2_sg U80675 ( .A(n56593), .X(n67588) );
  inv_x2_sg U80676 ( .A(n56591), .X(n67589) );
  inv_x2_sg U80677 ( .A(n56589), .X(n67590) );
  inv_x2_sg U80678 ( .A(n56587), .X(n67591) );
  inv_x2_sg U80679 ( .A(n56585), .X(n67592) );
  inv_x2_sg U80680 ( .A(n56583), .X(n67593) );
  inv_x2_sg U80681 ( .A(n56581), .X(n67594) );
  inv_x2_sg U80682 ( .A(n56579), .X(n67595) );
  inv_x2_sg U80683 ( .A(n56577), .X(n67596) );
  inv_x2_sg U80684 ( .A(n56575), .X(n67597) );
  inv_x2_sg U80685 ( .A(n56573), .X(n67598) );
  inv_x2_sg U80686 ( .A(n56571), .X(n67599) );
  inv_x2_sg U80687 ( .A(n56569), .X(n67600) );
  inv_x2_sg U80688 ( .A(n56567), .X(n67601) );
  inv_x2_sg U80689 ( .A(n56565), .X(n67602) );
  inv_x2_sg U80690 ( .A(n56563), .X(n67603) );
  inv_x2_sg U80691 ( .A(n56561), .X(n67604) );
  inv_x2_sg U80692 ( .A(n56559), .X(n67605) );
  inv_x2_sg U80693 ( .A(n56557), .X(n67606) );
  inv_x2_sg U80694 ( .A(n56555), .X(n67607) );
  inv_x2_sg U80695 ( .A(n56553), .X(n67608) );
  inv_x2_sg U80696 ( .A(n56551), .X(n67609) );
  inv_x2_sg U80697 ( .A(n56549), .X(n67610) );
  inv_x2_sg U80698 ( .A(n56547), .X(n67611) );
  inv_x2_sg U80699 ( .A(n56545), .X(n67612) );
  inv_x2_sg U80700 ( .A(n56543), .X(n67613) );
  inv_x2_sg U80701 ( .A(n56541), .X(n67614) );
  inv_x2_sg U80702 ( .A(n56539), .X(n67615) );
  inv_x2_sg U80703 ( .A(n56537), .X(n67616) );
  inv_x2_sg U80704 ( .A(n56535), .X(n67617) );
  inv_x2_sg U80705 ( .A(n56533), .X(n67618) );
  inv_x2_sg U80706 ( .A(n56531), .X(n67619) );
  inv_x2_sg U80707 ( .A(n56529), .X(n67620) );
  inv_x2_sg U80708 ( .A(n56527), .X(n67621) );
  inv_x2_sg U80709 ( .A(n56525), .X(n67622) );
  inv_x2_sg U80710 ( .A(n56523), .X(n67623) );
  inv_x2_sg U80711 ( .A(n56521), .X(n67624) );
  inv_x2_sg U80712 ( .A(n56519), .X(n67625) );
  inv_x2_sg U80713 ( .A(n56517), .X(n67626) );
  inv_x2_sg U80714 ( .A(n56515), .X(n67627) );
  inv_x2_sg U80715 ( .A(n56513), .X(n67628) );
  inv_x2_sg U80716 ( .A(n56511), .X(n67629) );
  inv_x2_sg U80717 ( .A(n56509), .X(n67630) );
  inv_x2_sg U80718 ( .A(n56507), .X(n67631) );
  inv_x2_sg U80719 ( .A(n56505), .X(n67632) );
  inv_x2_sg U80720 ( .A(n56503), .X(n67633) );
  inv_x2_sg U80721 ( .A(n56501), .X(n67634) );
  inv_x2_sg U80722 ( .A(n56499), .X(n67635) );
  inv_x2_sg U80723 ( .A(n56497), .X(n67636) );
  inv_x2_sg U80724 ( .A(n56495), .X(n67637) );
  inv_x2_sg U80725 ( .A(n56493), .X(n67638) );
  inv_x2_sg U80726 ( .A(n56491), .X(n67639) );
  inv_x2_sg U80727 ( .A(n56489), .X(n67640) );
  inv_x2_sg U80728 ( .A(n56487), .X(n67641) );
  inv_x2_sg U80729 ( .A(n56485), .X(n67642) );
  inv_x2_sg U80730 ( .A(n56483), .X(n67643) );
  inv_x2_sg U80731 ( .A(n56481), .X(n67644) );
  inv_x2_sg U80732 ( .A(n56479), .X(n67645) );
  inv_x2_sg U80733 ( .A(n56477), .X(n67646) );
  inv_x2_sg U80734 ( .A(n56475), .X(n67647) );
  inv_x2_sg U80735 ( .A(n56473), .X(n67648) );
  inv_x2_sg U80736 ( .A(n56471), .X(n67649) );
  inv_x2_sg U80737 ( .A(n56469), .X(n67650) );
  inv_x2_sg U80738 ( .A(n56467), .X(n67651) );
  inv_x2_sg U80739 ( .A(n56465), .X(n67652) );
  inv_x2_sg U80740 ( .A(n56463), .X(n67653) );
  inv_x2_sg U80741 ( .A(n56461), .X(n67654) );
  inv_x2_sg U80742 ( .A(n56459), .X(n67655) );
  inv_x2_sg U80743 ( .A(n56457), .X(n67656) );
  inv_x2_sg U80744 ( .A(n56455), .X(n67657) );
  inv_x2_sg U80745 ( .A(n56453), .X(n67658) );
  inv_x2_sg U80746 ( .A(n56451), .X(n67659) );
  inv_x2_sg U80747 ( .A(n56449), .X(n67660) );
  inv_x2_sg U80748 ( .A(n56447), .X(n67661) );
  inv_x2_sg U80749 ( .A(n56445), .X(n67662) );
  inv_x2_sg U80750 ( .A(n56443), .X(n67663) );
  inv_x2_sg U80751 ( .A(n56441), .X(n67664) );
  inv_x2_sg U80752 ( .A(n56439), .X(n67665) );
  inv_x2_sg U80753 ( .A(n56437), .X(n67666) );
  inv_x2_sg U80754 ( .A(n56435), .X(n67667) );
  inv_x2_sg U80755 ( .A(n56433), .X(n67668) );
  inv_x2_sg U80756 ( .A(n56431), .X(n67669) );
  inv_x2_sg U80757 ( .A(n56429), .X(n67670) );
  inv_x2_sg U80758 ( .A(n56427), .X(n67671) );
  inv_x2_sg U80759 ( .A(n56425), .X(n67672) );
  inv_x2_sg U80760 ( .A(n56423), .X(n67673) );
  inv_x2_sg U80761 ( .A(n56421), .X(n67674) );
  inv_x2_sg U80762 ( .A(n56419), .X(n67675) );
  inv_x2_sg U80763 ( .A(n56417), .X(n67676) );
  inv_x2_sg U80764 ( .A(n56415), .X(n67677) );
  inv_x2_sg U80765 ( .A(n56413), .X(n67678) );
  inv_x2_sg U80766 ( .A(n56411), .X(n67679) );
  inv_x2_sg U80767 ( .A(n56409), .X(n67680) );
  inv_x2_sg U80768 ( .A(n56407), .X(n67681) );
  inv_x2_sg U80769 ( .A(n56405), .X(n67682) );
  inv_x2_sg U80770 ( .A(n56403), .X(n67683) );
  inv_x2_sg U80771 ( .A(n56401), .X(n67684) );
  inv_x2_sg U80772 ( .A(n56399), .X(n67685) );
  inv_x2_sg U80773 ( .A(n56397), .X(n67686) );
  inv_x2_sg U80774 ( .A(n56395), .X(n67687) );
  inv_x2_sg U80775 ( .A(n56393), .X(n67688) );
  inv_x2_sg U80776 ( .A(n56391), .X(n67689) );
  inv_x2_sg U80777 ( .A(n56389), .X(n67690) );
  inv_x2_sg U80778 ( .A(n56387), .X(n67691) );
  inv_x2_sg U80779 ( .A(n56385), .X(n67692) );
  inv_x2_sg U80780 ( .A(n56383), .X(n67693) );
  inv_x2_sg U80781 ( .A(n56381), .X(n67694) );
  inv_x2_sg U80782 ( .A(n56379), .X(n67695) );
  inv_x2_sg U80783 ( .A(n56377), .X(n67696) );
  inv_x2_sg U80784 ( .A(n56375), .X(n67697) );
  inv_x2_sg U80785 ( .A(n56373), .X(n67698) );
  inv_x2_sg U80786 ( .A(n56371), .X(n67699) );
  inv_x2_sg U80787 ( .A(n56369), .X(n67700) );
  inv_x2_sg U80788 ( .A(n56367), .X(n67701) );
  inv_x2_sg U80789 ( .A(n56365), .X(n67702) );
  inv_x2_sg U80790 ( .A(n56363), .X(n67703) );
  inv_x2_sg U80791 ( .A(n56361), .X(n67704) );
  inv_x2_sg U80792 ( .A(n56359), .X(n67705) );
  inv_x2_sg U80793 ( .A(n56357), .X(n67706) );
  inv_x2_sg U80794 ( .A(n56355), .X(n67707) );
  inv_x2_sg U80795 ( .A(n56353), .X(n67708) );
  inv_x2_sg U80796 ( .A(n56351), .X(n67709) );
  inv_x2_sg U80797 ( .A(n56349), .X(n67710) );
  inv_x2_sg U80798 ( .A(n56347), .X(n67711) );
  inv_x2_sg U80799 ( .A(n56345), .X(n67712) );
  inv_x2_sg U80800 ( .A(n56343), .X(n67713) );
  inv_x2_sg U80801 ( .A(n56341), .X(n67714) );
  inv_x2_sg U80802 ( .A(n56339), .X(n67715) );
  inv_x2_sg U80803 ( .A(n56337), .X(n67716) );
  inv_x2_sg U80804 ( .A(n56335), .X(n67717) );
  inv_x2_sg U80805 ( .A(n56333), .X(n67718) );
  inv_x2_sg U80806 ( .A(n56331), .X(n67719) );
  inv_x2_sg U80807 ( .A(n56329), .X(n67720) );
  inv_x2_sg U80808 ( .A(n56327), .X(n67721) );
  inv_x2_sg U80809 ( .A(n56325), .X(n67722) );
  inv_x2_sg U80810 ( .A(n56323), .X(n67723) );
  inv_x2_sg U80811 ( .A(n56321), .X(n67724) );
  inv_x2_sg U80812 ( .A(n56319), .X(n67725) );
  inv_x2_sg U80813 ( .A(n56317), .X(n67726) );
  inv_x2_sg U80814 ( .A(n56315), .X(n67727) );
  inv_x2_sg U80815 ( .A(n56313), .X(n67728) );
  inv_x2_sg U80816 ( .A(n56311), .X(n67729) );
  inv_x2_sg U80817 ( .A(n56309), .X(n67730) );
  inv_x2_sg U80818 ( .A(n56307), .X(n67731) );
  inv_x2_sg U80819 ( .A(n56305), .X(n67732) );
  inv_x2_sg U80820 ( .A(n56303), .X(n67733) );
  inv_x2_sg U80821 ( .A(n56301), .X(n67734) );
  inv_x2_sg U80822 ( .A(n56299), .X(n67735) );
  inv_x2_sg U80823 ( .A(n56297), .X(n67736) );
  inv_x2_sg U80824 ( .A(n56295), .X(n67737) );
  inv_x2_sg U80825 ( .A(n56293), .X(n67738) );
  inv_x2_sg U80826 ( .A(n56291), .X(n67739) );
  inv_x2_sg U80827 ( .A(n56289), .X(n67740) );
  inv_x2_sg U80828 ( .A(n56287), .X(n67741) );
  inv_x2_sg U80829 ( .A(n56285), .X(n67742) );
  inv_x2_sg U80830 ( .A(n56283), .X(n67743) );
  inv_x2_sg U80831 ( .A(n56281), .X(n67744) );
  inv_x2_sg U80832 ( .A(n56279), .X(n67745) );
  inv_x2_sg U80833 ( .A(n56277), .X(n67746) );
  inv_x2_sg U80834 ( .A(n56275), .X(n67747) );
  inv_x2_sg U80835 ( .A(n56273), .X(n67748) );
  inv_x2_sg U80836 ( .A(n56271), .X(n67749) );
  inv_x2_sg U80837 ( .A(n56269), .X(n67750) );
  inv_x2_sg U80838 ( .A(n56267), .X(n67751) );
  inv_x2_sg U80839 ( .A(n56265), .X(n67752) );
  inv_x2_sg U80840 ( .A(n56263), .X(n67753) );
  inv_x2_sg U80841 ( .A(n56261), .X(n67754) );
  inv_x2_sg U80842 ( .A(n56259), .X(n67755) );
  inv_x2_sg U80843 ( .A(n56257), .X(n67756) );
  inv_x2_sg U80844 ( .A(n56255), .X(n67757) );
  inv_x2_sg U80845 ( .A(n56253), .X(n67758) );
  inv_x2_sg U80846 ( .A(n56251), .X(n67759) );
  inv_x2_sg U80847 ( .A(n56249), .X(n67760) );
  inv_x2_sg U80848 ( .A(n56247), .X(n67761) );
  inv_x2_sg U80849 ( .A(n56245), .X(n67762) );
  inv_x2_sg U80850 ( .A(n56243), .X(n67763) );
  inv_x2_sg U80851 ( .A(n56241), .X(n67764) );
  inv_x2_sg U80852 ( .A(n56239), .X(n67765) );
  inv_x2_sg U80853 ( .A(n56237), .X(n67766) );
  inv_x2_sg U80854 ( .A(n56235), .X(n67767) );
  inv_x2_sg U80855 ( .A(n56233), .X(n67768) );
  inv_x2_sg U80856 ( .A(n56231), .X(n67769) );
  inv_x2_sg U80857 ( .A(n56229), .X(n67770) );
  inv_x2_sg U80858 ( .A(n56227), .X(n67771) );
  inv_x2_sg U80859 ( .A(n56225), .X(n67772) );
  inv_x2_sg U80860 ( .A(n56223), .X(n67773) );
  inv_x2_sg U80861 ( .A(n56221), .X(n67774) );
  inv_x2_sg U80862 ( .A(n56219), .X(n67775) );
  inv_x2_sg U80863 ( .A(n56217), .X(n67776) );
  inv_x2_sg U80864 ( .A(n56215), .X(n67777) );
  inv_x2_sg U80865 ( .A(n56213), .X(n67778) );
  inv_x2_sg U80866 ( .A(n56211), .X(n67779) );
  inv_x2_sg U80867 ( .A(n56209), .X(n67780) );
  inv_x2_sg U80868 ( .A(n56207), .X(n67781) );
  inv_x2_sg U80869 ( .A(n56205), .X(n67782) );
  inv_x2_sg U80870 ( .A(n56203), .X(n67783) );
  inv_x2_sg U80871 ( .A(n56201), .X(n67784) );
  inv_x2_sg U80872 ( .A(n56199), .X(n67785) );
  inv_x2_sg U80873 ( .A(n56197), .X(n67786) );
  inv_x2_sg U80874 ( .A(n56195), .X(n67787) );
  inv_x2_sg U80875 ( .A(n56193), .X(n67788) );
  inv_x2_sg U80876 ( .A(n56191), .X(n67789) );
  inv_x2_sg U80877 ( .A(n56189), .X(n67790) );
  inv_x2_sg U80878 ( .A(n56187), .X(n67791) );
  inv_x2_sg U80879 ( .A(n56185), .X(n67792) );
  inv_x2_sg U80880 ( .A(n56183), .X(n67793) );
  inv_x2_sg U80881 ( .A(n56181), .X(n67794) );
  inv_x2_sg U80882 ( .A(n56179), .X(n67795) );
  inv_x2_sg U80883 ( .A(n56177), .X(n67796) );
  inv_x2_sg U80884 ( .A(n56175), .X(n67797) );
  inv_x2_sg U80885 ( .A(n56173), .X(n67798) );
  inv_x2_sg U80886 ( .A(n56171), .X(n67799) );
  inv_x2_sg U80887 ( .A(n56169), .X(n67800) );
  inv_x2_sg U80888 ( .A(n56167), .X(n67801) );
  inv_x2_sg U80889 ( .A(n56165), .X(n67802) );
  inv_x2_sg U80890 ( .A(n56163), .X(n67803) );
  inv_x2_sg U80891 ( .A(n56161), .X(n67804) );
  inv_x2_sg U80892 ( .A(n56159), .X(n67805) );
  inv_x2_sg U80893 ( .A(n56157), .X(n67806) );
  inv_x2_sg U80894 ( .A(n56155), .X(n67807) );
  inv_x2_sg U80895 ( .A(n56153), .X(n67808) );
  inv_x2_sg U80896 ( .A(n56151), .X(n67809) );
  inv_x2_sg U80897 ( .A(n56149), .X(n67810) );
  inv_x2_sg U80898 ( .A(n56147), .X(n67811) );
  inv_x2_sg U80899 ( .A(n56145), .X(n67812) );
  inv_x2_sg U80900 ( .A(n56143), .X(n67813) );
  inv_x2_sg U80901 ( .A(n56141), .X(n67814) );
  inv_x2_sg U80902 ( .A(n56139), .X(n67815) );
  inv_x2_sg U80903 ( .A(n56137), .X(n67816) );
  inv_x2_sg U80904 ( .A(n56135), .X(n67817) );
  inv_x2_sg U80905 ( .A(n56133), .X(n67818) );
  inv_x2_sg U80906 ( .A(n56131), .X(n67819) );
  inv_x2_sg U80907 ( .A(n56129), .X(n67820) );
  inv_x2_sg U80908 ( .A(n56127), .X(n67821) );
  inv_x2_sg U80909 ( .A(n56125), .X(n67822) );
  inv_x2_sg U80910 ( .A(n56123), .X(n67823) );
  inv_x2_sg U80911 ( .A(n56121), .X(n67824) );
  inv_x2_sg U80912 ( .A(n56119), .X(n67825) );
  inv_x2_sg U80913 ( .A(n56117), .X(n67826) );
  inv_x2_sg U80914 ( .A(n56115), .X(n67827) );
  inv_x2_sg U80915 ( .A(n56113), .X(n67828) );
  inv_x2_sg U80916 ( .A(n56111), .X(n67829) );
  inv_x2_sg U80917 ( .A(n56109), .X(n67830) );
  inv_x2_sg U80918 ( .A(n56107), .X(n67831) );
  inv_x2_sg U80919 ( .A(n56105), .X(n67832) );
  inv_x2_sg U80920 ( .A(n56103), .X(n67833) );
  inv_x2_sg U80921 ( .A(n56101), .X(n67834) );
  inv_x2_sg U80922 ( .A(n56099), .X(n67835) );
  inv_x2_sg U80923 ( .A(n56097), .X(n67836) );
  inv_x2_sg U80924 ( .A(n56095), .X(n67837) );
  inv_x2_sg U80925 ( .A(n56093), .X(n67838) );
  inv_x2_sg U80926 ( .A(n56091), .X(n67839) );
  inv_x2_sg U80927 ( .A(n56089), .X(n67840) );
  inv_x2_sg U80928 ( .A(n56087), .X(n67841) );
  inv_x2_sg U80929 ( .A(n56085), .X(n67842) );
  inv_x2_sg U80930 ( .A(n56083), .X(n67843) );
  inv_x2_sg U80931 ( .A(n56081), .X(n67844) );
  inv_x2_sg U80932 ( .A(n56079), .X(n67845) );
  inv_x2_sg U80933 ( .A(n56077), .X(n67846) );
  inv_x2_sg U80934 ( .A(n56075), .X(n67847) );
  inv_x2_sg U80935 ( .A(n56073), .X(n67848) );
  inv_x2_sg U80936 ( .A(n56071), .X(n67849) );
  inv_x2_sg U80937 ( .A(n56069), .X(n67850) );
  inv_x2_sg U80938 ( .A(n56067), .X(n67851) );
  inv_x2_sg U80939 ( .A(n56065), .X(n67852) );
  inv_x2_sg U80940 ( .A(n56063), .X(n67853) );
  inv_x2_sg U80941 ( .A(n56061), .X(n67854) );
  inv_x2_sg U80942 ( .A(n56059), .X(n67855) );
  inv_x2_sg U80943 ( .A(n56057), .X(n67856) );
  inv_x2_sg U80944 ( .A(n56055), .X(n67857) );
  inv_x2_sg U80945 ( .A(n56053), .X(n67858) );
  inv_x2_sg U80946 ( .A(n56051), .X(n67859) );
  inv_x2_sg U80947 ( .A(n56049), .X(n67860) );
  inv_x2_sg U80948 ( .A(n56047), .X(n67861) );
  inv_x2_sg U80949 ( .A(n56045), .X(n67862) );
  inv_x2_sg U80950 ( .A(n56043), .X(n67863) );
  inv_x2_sg U80951 ( .A(n56041), .X(n67864) );
  inv_x2_sg U80952 ( .A(n56039), .X(n67865) );
  inv_x2_sg U80953 ( .A(n56037), .X(n67866) );
  inv_x2_sg U80954 ( .A(n56035), .X(n67867) );
  inv_x2_sg U80955 ( .A(n56033), .X(n67868) );
  inv_x2_sg U80956 ( .A(n56031), .X(n67869) );
  inv_x2_sg U80957 ( .A(n56029), .X(n67870) );
  inv_x2_sg U80958 ( .A(n56027), .X(n67871) );
  inv_x2_sg U80959 ( .A(n56025), .X(n67872) );
  inv_x2_sg U80960 ( .A(n56023), .X(n67873) );
  inv_x2_sg U80961 ( .A(n56021), .X(n67874) );
  inv_x2_sg U80962 ( .A(n56019), .X(n67875) );
  inv_x2_sg U80963 ( .A(n56017), .X(n67876) );
  inv_x2_sg U80964 ( .A(n56015), .X(n67877) );
  inv_x2_sg U80965 ( .A(n56013), .X(n67878) );
  inv_x2_sg U80966 ( .A(n56011), .X(n67879) );
  inv_x2_sg U80967 ( .A(n56009), .X(n67880) );
  inv_x2_sg U80968 ( .A(n56007), .X(n67881) );
  inv_x2_sg U80969 ( .A(n56005), .X(n67882) );
  inv_x2_sg U80970 ( .A(n56003), .X(n67883) );
  inv_x2_sg U80971 ( .A(n56001), .X(n67884) );
  inv_x2_sg U80972 ( .A(n55999), .X(n67885) );
  inv_x2_sg U80973 ( .A(n55997), .X(n67886) );
  inv_x2_sg U80974 ( .A(n55995), .X(n67887) );
  inv_x2_sg U80975 ( .A(n55993), .X(n67888) );
  inv_x2_sg U80976 ( .A(n55991), .X(n67889) );
  inv_x2_sg U80977 ( .A(n55989), .X(n67890) );
  inv_x2_sg U80978 ( .A(n55987), .X(n67891) );
  inv_x2_sg U80979 ( .A(n55985), .X(n67892) );
  inv_x2_sg U80980 ( .A(n55983), .X(n67893) );
  inv_x2_sg U80981 ( .A(n55981), .X(n67894) );
  inv_x2_sg U80982 ( .A(n55979), .X(n67895) );
  inv_x2_sg U80983 ( .A(n55977), .X(n67896) );
  inv_x2_sg U80984 ( .A(n55975), .X(n67897) );
  inv_x2_sg U80985 ( .A(n55973), .X(n67898) );
  inv_x2_sg U80986 ( .A(n55971), .X(n67899) );
  inv_x2_sg U80987 ( .A(n55969), .X(n67900) );
  inv_x2_sg U80988 ( .A(n55967), .X(n67901) );
  inv_x2_sg U80989 ( .A(n55965), .X(n67902) );
  inv_x2_sg U80990 ( .A(n55963), .X(n67903) );
  inv_x2_sg U80991 ( .A(n55961), .X(n67904) );
  inv_x2_sg U80992 ( .A(n55959), .X(n67905) );
  inv_x2_sg U80993 ( .A(n55957), .X(n67906) );
  inv_x2_sg U80994 ( .A(n55955), .X(n67907) );
  inv_x2_sg U80995 ( .A(n55953), .X(n67908) );
  inv_x2_sg U80996 ( .A(n55951), .X(n67909) );
  inv_x2_sg U80997 ( .A(n55949), .X(n67910) );
  inv_x2_sg U80998 ( .A(n55947), .X(n67911) );
  inv_x2_sg U80999 ( .A(n55945), .X(n67912) );
  inv_x2_sg U81000 ( .A(n55943), .X(n67913) );
  inv_x2_sg U81001 ( .A(n55941), .X(n67914) );
  inv_x2_sg U81002 ( .A(n55939), .X(n67915) );
  inv_x2_sg U81003 ( .A(n55937), .X(n67916) );
  inv_x2_sg U81004 ( .A(n55935), .X(n67917) );
  inv_x2_sg U81005 ( .A(n55933), .X(n67918) );
  inv_x2_sg U81006 ( .A(n55931), .X(n67919) );
  inv_x2_sg U81007 ( .A(n55929), .X(n67920) );
  inv_x2_sg U81008 ( .A(n55927), .X(n67921) );
  inv_x2_sg U81009 ( .A(n55925), .X(n67922) );
  inv_x2_sg U81010 ( .A(n55923), .X(n67923) );
  inv_x2_sg U81011 ( .A(n55921), .X(n67924) );
  inv_x2_sg U81012 ( .A(n55919), .X(n67925) );
  inv_x2_sg U81013 ( .A(n55917), .X(n67926) );
  inv_x2_sg U81014 ( .A(n55915), .X(n67927) );
  inv_x2_sg U81015 ( .A(n55913), .X(n67928) );
  inv_x2_sg U81016 ( .A(n55911), .X(n67929) );
  inv_x2_sg U81017 ( .A(n55909), .X(n67930) );
  inv_x2_sg U81018 ( .A(n55907), .X(n67931) );
  inv_x2_sg U81019 ( .A(n55905), .X(n67932) );
  inv_x2_sg U81020 ( .A(n55903), .X(n67933) );
  inv_x2_sg U81021 ( .A(n55901), .X(n67934) );
  inv_x2_sg U81022 ( .A(n55899), .X(n67935) );
  inv_x2_sg U81023 ( .A(n55897), .X(n67936) );
  inv_x2_sg U81024 ( .A(n55895), .X(n67937) );
  inv_x2_sg U81025 ( .A(n55893), .X(n67938) );
  inv_x2_sg U81026 ( .A(n55891), .X(n67939) );
  inv_x2_sg U81027 ( .A(n55889), .X(n67940) );
  inv_x2_sg U81028 ( .A(n55887), .X(n67941) );
  inv_x2_sg U81029 ( .A(n55885), .X(n67942) );
  inv_x2_sg U81030 ( .A(n55883), .X(n67943) );
  inv_x2_sg U81031 ( .A(n55881), .X(n67944) );
  inv_x2_sg U81032 ( .A(n55879), .X(n67945) );
  inv_x2_sg U81033 ( .A(n55877), .X(n67946) );
  inv_x2_sg U81034 ( .A(n55875), .X(n67947) );
  inv_x2_sg U81035 ( .A(n55873), .X(n67948) );
  inv_x2_sg U81036 ( .A(n55871), .X(n67949) );
  inv_x2_sg U81037 ( .A(n55869), .X(n67950) );
  inv_x2_sg U81038 ( .A(n55867), .X(n67951) );
  inv_x2_sg U81039 ( .A(n55865), .X(n67952) );
  inv_x2_sg U81040 ( .A(n55863), .X(n67953) );
  inv_x2_sg U81041 ( .A(n55861), .X(n67954) );
  inv_x2_sg U81042 ( .A(n55859), .X(n67955) );
  inv_x2_sg U81043 ( .A(n55857), .X(n67956) );
  inv_x2_sg U81044 ( .A(n55855), .X(n67957) );
  inv_x2_sg U81045 ( .A(n55853), .X(n67958) );
  inv_x2_sg U81046 ( .A(n55851), .X(n67959) );
  inv_x2_sg U81047 ( .A(n55849), .X(n67960) );
  inv_x2_sg U81048 ( .A(n55847), .X(n67961) );
  inv_x2_sg U81049 ( .A(n55845), .X(n67962) );
  inv_x2_sg U81050 ( .A(n55843), .X(n67963) );
  inv_x2_sg U81051 ( .A(n55841), .X(n67964) );
  inv_x2_sg U81052 ( .A(n55839), .X(n67965) );
  inv_x2_sg U81053 ( .A(n55837), .X(n67966) );
  inv_x2_sg U81054 ( .A(n55835), .X(n67967) );
  inv_x2_sg U81055 ( .A(n55833), .X(n67968) );
  inv_x2_sg U81056 ( .A(n55831), .X(n67969) );
  inv_x2_sg U81057 ( .A(n55829), .X(n67970) );
  inv_x2_sg U81058 ( .A(n55827), .X(n67971) );
  inv_x2_sg U81059 ( .A(n55825), .X(n67972) );
  inv_x2_sg U81060 ( .A(n55823), .X(n67973) );
  inv_x2_sg U81061 ( .A(n55821), .X(n67974) );
  inv_x2_sg U81062 ( .A(n55819), .X(n67975) );
  inv_x2_sg U81063 ( .A(n55817), .X(n67976) );
  inv_x2_sg U81064 ( .A(n55815), .X(n67977) );
  inv_x2_sg U81065 ( .A(n55813), .X(n67978) );
  inv_x2_sg U81066 ( .A(n55811), .X(n67979) );
  inv_x2_sg U81067 ( .A(n55809), .X(n67980) );
  inv_x2_sg U81068 ( .A(n55807), .X(n67981) );
  inv_x2_sg U81069 ( .A(n55805), .X(n67982) );
  inv_x2_sg U81070 ( .A(n55803), .X(n67983) );
  inv_x2_sg U81071 ( .A(n55801), .X(n67984) );
  inv_x2_sg U81072 ( .A(n55799), .X(n67985) );
  inv_x2_sg U81073 ( .A(n55797), .X(n67986) );
  inv_x2_sg U81074 ( .A(n55795), .X(n67987) );
  inv_x2_sg U81075 ( .A(n55793), .X(n67988) );
  inv_x2_sg U81076 ( .A(n55791), .X(n67989) );
  inv_x2_sg U81077 ( .A(n55789), .X(n67990) );
  inv_x2_sg U81078 ( .A(n55787), .X(n67991) );
  inv_x2_sg U81079 ( .A(n55785), .X(n67992) );
  inv_x2_sg U81080 ( .A(n55783), .X(n67993) );
  inv_x2_sg U81081 ( .A(n55781), .X(n67994) );
  inv_x2_sg U81082 ( .A(n55779), .X(n67995) );
  inv_x2_sg U81083 ( .A(n55777), .X(n67996) );
  inv_x2_sg U81084 ( .A(n55775), .X(n67997) );
  inv_x2_sg U81085 ( .A(n55773), .X(n67998) );
  inv_x2_sg U81086 ( .A(n55771), .X(n67999) );
  inv_x2_sg U81087 ( .A(n55769), .X(n68000) );
  inv_x2_sg U81088 ( .A(n55767), .X(n68001) );
  inv_x2_sg U81089 ( .A(n55765), .X(n68002) );
  inv_x2_sg U81090 ( .A(n55763), .X(n68003) );
  inv_x2_sg U81091 ( .A(n55761), .X(n68004) );
  inv_x2_sg U81092 ( .A(n55759), .X(n68005) );
  inv_x2_sg U81093 ( .A(n55757), .X(n68006) );
  inv_x2_sg U81094 ( .A(n55755), .X(n68007) );
  inv_x2_sg U81095 ( .A(n55753), .X(n68008) );
  inv_x2_sg U81096 ( .A(n55751), .X(n68009) );
  inv_x2_sg U81097 ( .A(n55749), .X(n68010) );
  inv_x2_sg U81098 ( .A(n55747), .X(n68011) );
  inv_x2_sg U81099 ( .A(n55745), .X(n68012) );
  inv_x2_sg U81100 ( .A(n55743), .X(n68013) );
  inv_x2_sg U81101 ( .A(n55741), .X(n68014) );
  inv_x2_sg U81102 ( .A(n55739), .X(n68015) );
  inv_x2_sg U81103 ( .A(n55737), .X(n68016) );
  inv_x2_sg U81104 ( .A(n55735), .X(n68017) );
  inv_x2_sg U81105 ( .A(n55733), .X(n68018) );
  inv_x2_sg U81106 ( .A(n55731), .X(n68019) );
  inv_x2_sg U81107 ( .A(n55729), .X(n68020) );
  inv_x2_sg U81108 ( .A(n55727), .X(n68021) );
  inv_x2_sg U81109 ( .A(n55725), .X(n68022) );
  inv_x2_sg U81110 ( .A(n55723), .X(n68023) );
  inv_x2_sg U81111 ( .A(n55721), .X(n68024) );
  inv_x2_sg U81112 ( .A(n55719), .X(n68025) );
  inv_x2_sg U81113 ( .A(n55717), .X(n68026) );
  inv_x2_sg U81114 ( .A(n55715), .X(n68027) );
  inv_x2_sg U81115 ( .A(n55713), .X(n68028) );
  inv_x2_sg U81116 ( .A(n55711), .X(n68029) );
  inv_x2_sg U81117 ( .A(n55709), .X(n68030) );
  inv_x2_sg U81118 ( .A(n55707), .X(n68031) );
  inv_x2_sg U81119 ( .A(n55705), .X(n68032) );
  inv_x2_sg U81120 ( .A(n55703), .X(n68033) );
  inv_x2_sg U81121 ( .A(n55701), .X(n68034) );
  inv_x2_sg U81122 ( .A(n55699), .X(n68035) );
  inv_x2_sg U81123 ( .A(n55697), .X(n68036) );
  inv_x2_sg U81124 ( .A(n55695), .X(n68037) );
  inv_x2_sg U81125 ( .A(n55693), .X(n68038) );
  inv_x2_sg U81126 ( .A(n55691), .X(n68039) );
  inv_x2_sg U81127 ( .A(n55689), .X(n68040) );
  inv_x2_sg U81128 ( .A(n55687), .X(n68041) );
  inv_x2_sg U81129 ( .A(n55685), .X(n68042) );
  inv_x2_sg U81130 ( .A(n55683), .X(n68043) );
  inv_x2_sg U81131 ( .A(n55681), .X(n68044) );
  inv_x2_sg U81132 ( .A(n55679), .X(n68045) );
  inv_x2_sg U81133 ( .A(n55677), .X(n68046) );
  inv_x2_sg U81134 ( .A(n55675), .X(n68047) );
  inv_x2_sg U81135 ( .A(n55673), .X(n68048) );
  inv_x2_sg U81136 ( .A(n55671), .X(n68049) );
  inv_x2_sg U81137 ( .A(n55669), .X(n68050) );
  inv_x2_sg U81138 ( .A(n55667), .X(n68051) );
  inv_x2_sg U81139 ( .A(n55665), .X(n68052) );
  inv_x2_sg U81140 ( .A(n55663), .X(n68053) );
  inv_x2_sg U81141 ( .A(n55661), .X(n68054) );
  inv_x2_sg U81142 ( .A(n55659), .X(n68055) );
  inv_x2_sg U81143 ( .A(n55657), .X(n68056) );
  inv_x2_sg U81144 ( .A(n55655), .X(n68057) );
  inv_x2_sg U81145 ( .A(n55653), .X(n68058) );
  inv_x2_sg U81146 ( .A(n55651), .X(n68059) );
  inv_x2_sg U81147 ( .A(n55649), .X(n68060) );
  inv_x2_sg U81148 ( .A(n55647), .X(n68061) );
  inv_x2_sg U81149 ( .A(n55645), .X(n68062) );
  inv_x2_sg U81150 ( .A(n55643), .X(n68063) );
  inv_x2_sg U81151 ( .A(n55641), .X(n68064) );
  inv_x2_sg U81152 ( .A(n55639), .X(n68065) );
  inv_x2_sg U81153 ( .A(n55637), .X(n68066) );
  inv_x2_sg U81154 ( .A(n55635), .X(n68067) );
  inv_x2_sg U81155 ( .A(n55633), .X(n68068) );
  inv_x2_sg U81156 ( .A(n55631), .X(n68069) );
  inv_x2_sg U81157 ( .A(n55629), .X(n68070) );
  inv_x2_sg U81158 ( .A(n55627), .X(n68071) );
  inv_x2_sg U81159 ( .A(n55625), .X(n68072) );
  inv_x2_sg U81160 ( .A(n55623), .X(n68073) );
  inv_x2_sg U81161 ( .A(n55621), .X(n68074) );
  inv_x2_sg U81162 ( .A(n55619), .X(n68075) );
  inv_x2_sg U81163 ( .A(n55617), .X(n68076) );
  inv_x2_sg U81164 ( .A(n55615), .X(n68077) );
  inv_x2_sg U81165 ( .A(n55613), .X(n68078) );
  inv_x2_sg U81166 ( .A(n55611), .X(n68079) );
  inv_x2_sg U81167 ( .A(n55609), .X(n68080) );
  inv_x2_sg U81168 ( .A(n55607), .X(n68081) );
  inv_x2_sg U81169 ( .A(n55605), .X(n68082) );
  inv_x2_sg U81170 ( .A(n55603), .X(n68083) );
  inv_x2_sg U81171 ( .A(n55601), .X(n68084) );
  inv_x2_sg U81172 ( .A(n55599), .X(n68085) );
  inv_x2_sg U81173 ( .A(n55597), .X(n68086) );
  inv_x2_sg U81174 ( .A(n55595), .X(n68087) );
  inv_x2_sg U81175 ( .A(n55593), .X(n68088) );
  inv_x2_sg U81176 ( .A(n55591), .X(n68089) );
  inv_x2_sg U81177 ( .A(n55589), .X(n68090) );
  inv_x2_sg U81178 ( .A(n55587), .X(n68091) );
  inv_x2_sg U81179 ( .A(n55585), .X(n68092) );
  inv_x2_sg U81180 ( .A(n55583), .X(n68093) );
  inv_x2_sg U81181 ( .A(n55581), .X(n68094) );
  inv_x2_sg U81182 ( .A(n55579), .X(n68095) );
  inv_x2_sg U81183 ( .A(n55577), .X(n68096) );
  inv_x2_sg U81184 ( .A(n55575), .X(n68097) );
  inv_x2_sg U81185 ( .A(n55573), .X(n68098) );
  inv_x2_sg U81186 ( .A(n55571), .X(n68099) );
  inv_x2_sg U81187 ( .A(n55569), .X(n68100) );
  inv_x2_sg U81188 ( .A(n55567), .X(n68101) );
  inv_x2_sg U81189 ( .A(n55565), .X(n68102) );
  inv_x2_sg U81190 ( .A(n55563), .X(n68103) );
  inv_x2_sg U81191 ( .A(n55561), .X(n68104) );
  inv_x2_sg U81192 ( .A(n55559), .X(n68105) );
  inv_x2_sg U81193 ( .A(n55557), .X(n68106) );
  inv_x2_sg U81194 ( .A(n55555), .X(n68107) );
  inv_x2_sg U81195 ( .A(n55553), .X(n68108) );
  inv_x2_sg U81196 ( .A(n55551), .X(n68109) );
  inv_x2_sg U81197 ( .A(n55549), .X(n68110) );
  inv_x2_sg U81198 ( .A(n55547), .X(n68111) );
  inv_x2_sg U81199 ( .A(n55545), .X(n68112) );
  inv_x2_sg U81200 ( .A(n55543), .X(n68113) );
  inv_x2_sg U81201 ( .A(n55541), .X(n68114) );
  inv_x2_sg U81202 ( .A(n55539), .X(n68115) );
  inv_x2_sg U81203 ( .A(n55537), .X(n68116) );
  inv_x2_sg U81204 ( .A(n55535), .X(n68117) );
  inv_x2_sg U81205 ( .A(n55533), .X(n68118) );
  inv_x2_sg U81206 ( .A(n55531), .X(n68119) );
  inv_x2_sg U81207 ( .A(n55529), .X(n68120) );
  inv_x2_sg U81208 ( .A(n55527), .X(n68121) );
  inv_x2_sg U81209 ( .A(n55525), .X(n68122) );
  inv_x2_sg U81210 ( .A(n55523), .X(n68123) );
  inv_x2_sg U81211 ( .A(n55521), .X(n68124) );
  inv_x2_sg U81212 ( .A(n55519), .X(n68125) );
  inv_x2_sg U81213 ( .A(n55517), .X(n68126) );
  inv_x2_sg U81214 ( .A(n55515), .X(n68127) );
  inv_x2_sg U81215 ( .A(n55513), .X(n68128) );
  inv_x2_sg U81216 ( .A(n55511), .X(n68129) );
  inv_x2_sg U81217 ( .A(n55509), .X(n68130) );
  inv_x2_sg U81218 ( .A(n55507), .X(n68131) );
  inv_x2_sg U81219 ( .A(n55505), .X(n68132) );
  inv_x2_sg U81220 ( .A(n55503), .X(n68133) );
  inv_x2_sg U81221 ( .A(n55501), .X(n68134) );
  inv_x2_sg U81222 ( .A(n55499), .X(n68135) );
  inv_x2_sg U81223 ( .A(n55497), .X(n68136) );
  inv_x2_sg U81224 ( .A(n55495), .X(n68137) );
  inv_x2_sg U81225 ( .A(n55493), .X(n68138) );
  inv_x2_sg U81226 ( .A(n55491), .X(n68139) );
  inv_x2_sg U81227 ( .A(n55489), .X(n68140) );
  inv_x2_sg U81228 ( .A(n55487), .X(n68141) );
  inv_x2_sg U81229 ( .A(n55485), .X(n68142) );
  inv_x2_sg U81230 ( .A(n55483), .X(n68143) );
  inv_x2_sg U81231 ( .A(n55481), .X(n68144) );
  inv_x2_sg U81232 ( .A(n55479), .X(n68145) );
  inv_x2_sg U81233 ( .A(n55477), .X(n68146) );
  inv_x2_sg U81234 ( .A(n55475), .X(n68147) );
  inv_x2_sg U81235 ( .A(n55473), .X(n68148) );
  inv_x2_sg U81236 ( .A(n55471), .X(n68149) );
  inv_x2_sg U81237 ( .A(n55469), .X(n68150) );
  inv_x2_sg U81238 ( .A(n55467), .X(n68151) );
  inv_x2_sg U81239 ( .A(n55465), .X(n68152) );
  inv_x2_sg U81240 ( .A(n55463), .X(n68153) );
  inv_x2_sg U81241 ( .A(n55461), .X(n68154) );
  inv_x2_sg U81242 ( .A(n55459), .X(n68155) );
  inv_x2_sg U81243 ( .A(n55457), .X(n68156) );
  inv_x2_sg U81244 ( .A(n55455), .X(n68157) );
  inv_x2_sg U81245 ( .A(n55453), .X(n68158) );
  inv_x2_sg U81246 ( .A(n55451), .X(n68159) );
  inv_x2_sg U81247 ( .A(n55449), .X(n68160) );
  inv_x2_sg U81248 ( .A(n55447), .X(n68161) );
  inv_x2_sg U81249 ( .A(n55445), .X(n68162) );
  inv_x2_sg U81250 ( .A(n55443), .X(n68163) );
  inv_x2_sg U81251 ( .A(n55441), .X(n68164) );
  inv_x2_sg U81252 ( .A(n55439), .X(n68165) );
  inv_x2_sg U81253 ( .A(n55437), .X(n68166) );
  inv_x2_sg U81254 ( .A(n55435), .X(n68167) );
  inv_x2_sg U81255 ( .A(n55433), .X(n68168) );
  inv_x2_sg U81256 ( .A(n55431), .X(n68169) );
  inv_x2_sg U81257 ( .A(n55429), .X(n68170) );
  inv_x2_sg U81258 ( .A(n55427), .X(n68171) );
  inv_x2_sg U81259 ( .A(n55425), .X(n68172) );
  inv_x2_sg U81260 ( .A(n55423), .X(n68173) );
  inv_x2_sg U81261 ( .A(n55421), .X(n68174) );
  inv_x2_sg U81262 ( .A(n55419), .X(n68175) );
  inv_x2_sg U81263 ( .A(n55417), .X(n68176) );
  inv_x2_sg U81264 ( .A(n55415), .X(n68177) );
  inv_x2_sg U81265 ( .A(n55413), .X(n68178) );
  inv_x2_sg U81266 ( .A(n55411), .X(n68179) );
  inv_x2_sg U81267 ( .A(n55409), .X(n68180) );
  inv_x2_sg U81268 ( .A(n55407), .X(n68181) );
  inv_x2_sg U81269 ( .A(n55405), .X(n68182) );
  inv_x2_sg U81270 ( .A(n55403), .X(n68183) );
  inv_x2_sg U81271 ( .A(n55401), .X(n68184) );
  inv_x2_sg U81272 ( .A(n55399), .X(n68185) );
  inv_x2_sg U81273 ( .A(n55397), .X(n68186) );
  inv_x2_sg U81274 ( .A(n55395), .X(n68187) );
  inv_x2_sg U81275 ( .A(n55393), .X(n68188) );
  inv_x2_sg U81276 ( .A(n55391), .X(n68189) );
  inv_x2_sg U81277 ( .A(n55389), .X(n68190) );
  inv_x2_sg U81278 ( .A(n55387), .X(n68191) );
  inv_x2_sg U81279 ( .A(n55385), .X(n68192) );
  inv_x2_sg U81280 ( .A(n55383), .X(n68193) );
  inv_x2_sg U81281 ( .A(n55381), .X(n68194) );
  inv_x2_sg U81282 ( .A(n55379), .X(n68195) );
  inv_x2_sg U81283 ( .A(n55377), .X(n68196) );
  inv_x2_sg U81284 ( .A(n55375), .X(n68197) );
  inv_x2_sg U81285 ( .A(n55373), .X(n68198) );
  inv_x2_sg U81286 ( .A(n55371), .X(n68199) );
  inv_x2_sg U81287 ( .A(n55369), .X(n68200) );
  inv_x2_sg U81288 ( .A(n55367), .X(n68201) );
  inv_x2_sg U81289 ( .A(n55365), .X(n68202) );
  inv_x2_sg U81290 ( .A(n55363), .X(n68203) );
  inv_x2_sg U81291 ( .A(n55361), .X(n68204) );
  inv_x2_sg U81292 ( .A(n55359), .X(n68205) );
  inv_x2_sg U81293 ( .A(n55357), .X(n68206) );
  inv_x2_sg U81294 ( .A(n55355), .X(n68207) );
  inv_x2_sg U81295 ( .A(n55353), .X(n68208) );
  inv_x2_sg U81296 ( .A(n55351), .X(n68209) );
  inv_x2_sg U81297 ( .A(n55349), .X(n68210) );
  inv_x2_sg U81298 ( .A(n55347), .X(n68211) );
  inv_x2_sg U81299 ( .A(n55345), .X(n68212) );
  inv_x2_sg U81300 ( .A(n55343), .X(n68213) );
  inv_x2_sg U81301 ( .A(n55341), .X(n68214) );
  inv_x2_sg U81302 ( .A(n55339), .X(n68215) );
  inv_x2_sg U81303 ( .A(n55337), .X(n68216) );
  inv_x2_sg U81304 ( .A(n55335), .X(n68217) );
  inv_x2_sg U81305 ( .A(n55333), .X(n68218) );
  inv_x2_sg U81306 ( .A(n55331), .X(n68219) );
  inv_x2_sg U81307 ( .A(n55329), .X(n68220) );
  inv_x2_sg U81308 ( .A(n55327), .X(n68221) );
  inv_x2_sg U81309 ( .A(n55325), .X(n68222) );
  inv_x2_sg U81310 ( .A(n55323), .X(n68223) );
  inv_x2_sg U81311 ( .A(n55321), .X(n68224) );
  inv_x2_sg U81312 ( .A(n55319), .X(n68225) );
  inv_x2_sg U81313 ( .A(n55317), .X(n68226) );
  inv_x2_sg U81314 ( .A(n26269), .X(n67564) );
  inv_x2_sg U81315 ( .A(n26296), .X(n67566) );
  inv_x2_sg U81316 ( .A(n51059), .X(n67567) );
  inv_x2_sg U81317 ( .A(n26305), .X(n67569) );
  inv_x2_sg U81318 ( .A(n51063), .X(n67571) );
  inv_x2_sg U81319 ( .A(n51061), .X(n67572) );
  inv_x2_sg U81320 ( .A(n57081), .X(n67087) );
  inv_x2_sg U81321 ( .A(n51549), .X(n67088) );
  inv_x2_sg U81322 ( .A(n57089), .X(n67089) );
  inv_x2_sg U81323 ( .A(n57087), .X(n67090) );
  inv_x2_sg U81324 ( .A(n51553), .X(n67091) );
  inv_x2_sg U81325 ( .A(n57079), .X(n67092) );
  inv_x2_sg U81326 ( .A(n57071), .X(n67093) );
  inv_x2_sg U81327 ( .A(n51545), .X(n67094) );
  inv_x2_sg U81328 ( .A(n47773), .X(n67095) );
  inv_x2_sg U81329 ( .A(n26002), .X(n67475) );
  inv_x2_sg U81330 ( .A(n25911), .X(n67476) );
  inv_x2_sg U81331 ( .A(n25881), .X(n67477) );
  inv_x2_sg U81332 ( .A(n25851), .X(n67478) );
  inv_x2_sg U81333 ( .A(n25761), .X(n67479) );
  inv_x2_sg U81334 ( .A(n25731), .X(n67480) );
  inv_x2_sg U81335 ( .A(n25641), .X(n67481) );
  inv_x2_sg U81336 ( .A(n25611), .X(n67482) );
  inv_x2_sg U81337 ( .A(n25581), .X(n67483) );
  inv_x2_sg U81338 ( .A(n25491), .X(n67484) );
  inv_x2_sg U81339 ( .A(n25461), .X(n67485) );
  inv_x2_sg U81340 ( .A(n25431), .X(n67486) );
  inv_x2_sg U81341 ( .A(n25400), .X(n67282) );
  inv_x2_sg U81342 ( .A(n25309), .X(n67283) );
  inv_x2_sg U81343 ( .A(n25279), .X(n67284) );
  inv_x2_sg U81344 ( .A(n25249), .X(n67285) );
  inv_x2_sg U81345 ( .A(n25159), .X(n67286) );
  inv_x2_sg U81346 ( .A(n25129), .X(n67287) );
  inv_x2_sg U81347 ( .A(n25039), .X(n67288) );
  inv_x2_sg U81348 ( .A(n25009), .X(n67289) );
  inv_x2_sg U81349 ( .A(n24979), .X(n67290) );
  inv_x2_sg U81350 ( .A(n24889), .X(n67291) );
  inv_x2_sg U81351 ( .A(n24859), .X(n67292) );
  inv_x2_sg U81352 ( .A(n24828), .X(n67293) );
  inv_x2_sg U81353 ( .A(n51543), .X(n67306) );
  inv_x2_sg U81354 ( .A(n57085), .X(n67308) );
  inv_x2_sg U81355 ( .A(n57083), .X(n67309) );
  inv_x2_sg U81356 ( .A(n51551), .X(n67310) );
  inv_x2_sg U81357 ( .A(n57077), .X(n67311) );
  inv_x2_sg U81358 ( .A(n57075), .X(n67312) );
  inv_x2_sg U81359 ( .A(n51547), .X(n67313) );
  inv_x2_sg U81360 ( .A(n57073), .X(n67314) );
  inv_x2_sg U81361 ( .A(n32041), .X(n68267) );
  inv_x2_sg U81362 ( .A(n35839), .X(n68269) );
  inv_x2_sg U81363 ( .A(n51065), .X(n68270) );
  inv_x2_sg U81364 ( .A(n32428), .X(n68407) );
  inv_x2_sg U81365 ( .A(n32450), .X(n68416) );
  inv_x2_sg U81366 ( .A(n32453), .X(n68417) );
  inv_x2_sg U81367 ( .A(n32458), .X(n68418) );
  inv_x2_sg U81368 ( .A(n32461), .X(n68419) );
  inv_x2_sg U81369 ( .A(n32433), .X(n68420) );
  inv_x2_sg U81370 ( .A(n32626), .X(n68421) );
  inv_x2_sg U81371 ( .A(n32629), .X(n68422) );
  inv_x2_sg U81372 ( .A(n32634), .X(n68423) );
  inv_x2_sg U81373 ( .A(n32637), .X(n68424) );
  inv_x2_sg U81374 ( .A(n32513), .X(n68425) );
  inv_x2_sg U81375 ( .A(n32587), .X(n68434) );
  inv_x2_sg U81376 ( .A(n32590), .X(n68435) );
  inv_x2_sg U81377 ( .A(n32595), .X(n68436) );
  inv_x2_sg U81378 ( .A(n32598), .X(n68437) );
  inv_x2_sg U81379 ( .A(n32567), .X(n68438) );
  inv_x2_sg U81380 ( .A(n32570), .X(n68439) );
  inv_x2_sg U81381 ( .A(n32575), .X(n68440) );
  inv_x2_sg U81382 ( .A(n32578), .X(n68441) );
  inv_x2_sg U81383 ( .A(n32721), .X(n68443) );
  inv_x2_sg U81384 ( .A(n32728), .X(n68444) );
  inv_x2_sg U81385 ( .A(n32731), .X(n68445) );
  inv_x2_sg U81386 ( .A(n32736), .X(n68446) );
  inv_x2_sg U81387 ( .A(n32739), .X(n68447) );
  inv_x2_sg U81388 ( .A(n32749), .X(n68449) );
  inv_x2_sg U81389 ( .A(n32752), .X(n68450) );
  inv_x2_sg U81390 ( .A(n32757), .X(n68451) );
  inv_x2_sg U81391 ( .A(n32760), .X(n68452) );
  inv_x2_sg U81392 ( .A(n32779), .X(n68453) );
  inv_x2_sg U81393 ( .A(n32786), .X(n68454) );
  inv_x2_sg U81394 ( .A(n32789), .X(n68455) );
  inv_x2_sg U81395 ( .A(n32794), .X(n68456) );
  inv_x2_sg U81396 ( .A(n32797), .X(n68457) );
  inv_x2_sg U81397 ( .A(n32709), .X(n68459) );
  inv_x2_sg U81398 ( .A(n32712), .X(n68460) );
  inv_x2_sg U81399 ( .A(n32717), .X(n68461) );
  inv_x2_sg U81400 ( .A(n32720), .X(n68462) );
  inv_x2_sg U81401 ( .A(n32520), .X(n68463) );
  inv_x2_sg U81402 ( .A(n32767), .X(n68464) );
  inv_x2_sg U81403 ( .A(n32770), .X(n68465) );
  inv_x2_sg U81404 ( .A(n32775), .X(n68466) );
  inv_x2_sg U81405 ( .A(n32778), .X(n68467) );
  inv_x2_sg U81406 ( .A(n32673), .X(n68468) );
  inv_x2_sg U81407 ( .A(n32676), .X(n68469) );
  inv_x2_sg U81408 ( .A(n32681), .X(n68470) );
  inv_x2_sg U81409 ( .A(n32684), .X(n68471) );
  inv_x2_sg U81410 ( .A(n32691), .X(n68473) );
  inv_x2_sg U81411 ( .A(n32694), .X(n68474) );
  inv_x2_sg U81412 ( .A(n32699), .X(n68475) );
  inv_x2_sg U81413 ( .A(n32702), .X(n68476) );
  inv_x2_sg U81414 ( .A(n31961), .X(n68496) );
  inv_x2_sg U81415 ( .A(n32008), .X(n68505) );
  inv_x2_sg U81416 ( .A(n32011), .X(n68506) );
  inv_x2_sg U81417 ( .A(n32016), .X(n68507) );
  inv_x2_sg U81418 ( .A(n32019), .X(n68508) );
  inv_x2_sg U81419 ( .A(n31966), .X(n68509) );
  inv_x2_sg U81420 ( .A(n32181), .X(n68510) );
  inv_x2_sg U81421 ( .A(n32184), .X(n68511) );
  inv_x2_sg U81422 ( .A(n32189), .X(n68512) );
  inv_x2_sg U81423 ( .A(n32192), .X(n68513) );
  inv_x2_sg U81424 ( .A(n32067), .X(n68514) );
  inv_x2_sg U81425 ( .A(n32142), .X(n68525) );
  inv_x2_sg U81426 ( .A(n32145), .X(n68526) );
  inv_x2_sg U81427 ( .A(n32150), .X(n68527) );
  inv_x2_sg U81428 ( .A(n32153), .X(n68528) );
  inv_x2_sg U81429 ( .A(n32122), .X(n68530) );
  inv_x2_sg U81430 ( .A(n32125), .X(n68531) );
  inv_x2_sg U81431 ( .A(n32130), .X(n68532) );
  inv_x2_sg U81432 ( .A(n32133), .X(n68533) );
  inv_x2_sg U81433 ( .A(n32276), .X(n68536) );
  inv_x2_sg U81434 ( .A(n32283), .X(n68537) );
  inv_x2_sg U81435 ( .A(n32286), .X(n68538) );
  inv_x2_sg U81436 ( .A(n32291), .X(n68539) );
  inv_x2_sg U81437 ( .A(n32294), .X(n68540) );
  inv_x2_sg U81438 ( .A(n32304), .X(n68542) );
  inv_x2_sg U81439 ( .A(n32307), .X(n68543) );
  inv_x2_sg U81440 ( .A(n32312), .X(n68544) );
  inv_x2_sg U81441 ( .A(n32315), .X(n68545) );
  inv_x2_sg U81442 ( .A(n32334), .X(n68546) );
  inv_x2_sg U81443 ( .A(n32341), .X(n68547) );
  inv_x2_sg U81444 ( .A(n32344), .X(n68548) );
  inv_x2_sg U81445 ( .A(n32349), .X(n68549) );
  inv_x2_sg U81446 ( .A(n32352), .X(n68550) );
  inv_x2_sg U81447 ( .A(n32264), .X(n68552) );
  inv_x2_sg U81448 ( .A(n32267), .X(n68553) );
  inv_x2_sg U81449 ( .A(n32272), .X(n68554) );
  inv_x2_sg U81450 ( .A(n32275), .X(n68555) );
  inv_x2_sg U81451 ( .A(n32075), .X(n68556) );
  inv_x2_sg U81452 ( .A(n32322), .X(n68557) );
  inv_x2_sg U81453 ( .A(n32325), .X(n68558) );
  inv_x2_sg U81454 ( .A(n32330), .X(n68559) );
  inv_x2_sg U81455 ( .A(n32333), .X(n68560) );
  inv_x2_sg U81456 ( .A(n32228), .X(n68561) );
  inv_x2_sg U81457 ( .A(n32231), .X(n68562) );
  inv_x2_sg U81458 ( .A(n32236), .X(n68563) );
  inv_x2_sg U81459 ( .A(n32239), .X(n68564) );
  inv_x2_sg U81460 ( .A(n32246), .X(n68566) );
  inv_x2_sg U81461 ( .A(n32249), .X(n68567) );
  inv_x2_sg U81462 ( .A(n32254), .X(n68568) );
  inv_x2_sg U81463 ( .A(n32257), .X(n68569) );
endmodule

