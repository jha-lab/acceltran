
module fifo ( clk, reset, data_in, rd_en, wr_en, empty, full, data_out );
  input [19:0] data_in;
  output [19:0] data_out;
  input clk, reset, rd_en, wr_en;
  output empty, full;
  wire   \buff_mem[19][19] , \buff_mem[19][18] , \buff_mem[19][17] ,
         \buff_mem[19][16] , \buff_mem[19][15] , \buff_mem[19][14] ,
         \buff_mem[19][13] , \buff_mem[19][12] , \buff_mem[19][11] ,
         \buff_mem[19][10] , \buff_mem[19][9] , \buff_mem[19][8] ,
         \buff_mem[19][7] , \buff_mem[19][6] , \buff_mem[19][5] ,
         \buff_mem[19][4] , \buff_mem[19][3] , \buff_mem[19][2] ,
         \buff_mem[19][1] , \buff_mem[19][0] , \buff_mem[18][19] ,
         \buff_mem[18][18] , \buff_mem[18][17] , \buff_mem[18][16] ,
         \buff_mem[18][15] , \buff_mem[18][14] , \buff_mem[18][13] ,
         \buff_mem[18][12] , \buff_mem[18][11] , \buff_mem[18][10] ,
         \buff_mem[18][9] , \buff_mem[18][8] , \buff_mem[18][7] ,
         \buff_mem[18][6] , \buff_mem[18][5] , \buff_mem[18][4] ,
         \buff_mem[18][3] , \buff_mem[18][2] , \buff_mem[18][1] ,
         \buff_mem[18][0] , \buff_mem[17][19] , \buff_mem[17][18] ,
         \buff_mem[17][17] , \buff_mem[17][16] , \buff_mem[17][15] ,
         \buff_mem[17][14] , \buff_mem[17][13] , \buff_mem[17][12] ,
         \buff_mem[17][11] , \buff_mem[17][10] , \buff_mem[17][9] ,
         \buff_mem[17][8] , \buff_mem[17][7] , \buff_mem[17][6] ,
         \buff_mem[17][5] , \buff_mem[17][4] , \buff_mem[17][3] ,
         \buff_mem[17][2] , \buff_mem[17][1] , \buff_mem[17][0] ,
         \buff_mem[16][19] , \buff_mem[16][18] , \buff_mem[16][17] ,
         \buff_mem[16][16] , \buff_mem[16][15] , \buff_mem[16][14] ,
         \buff_mem[16][13] , \buff_mem[16][12] , \buff_mem[16][11] ,
         \buff_mem[16][10] , \buff_mem[16][9] , \buff_mem[16][8] ,
         \buff_mem[16][7] , \buff_mem[16][6] , \buff_mem[16][5] ,
         \buff_mem[16][4] , \buff_mem[16][3] , \buff_mem[16][2] ,
         \buff_mem[16][1] , \buff_mem[16][0] , \buff_mem[15][19] ,
         \buff_mem[15][18] , \buff_mem[15][17] , \buff_mem[15][16] ,
         \buff_mem[15][15] , \buff_mem[15][14] , \buff_mem[15][13] ,
         \buff_mem[15][12] , \buff_mem[15][11] , \buff_mem[15][10] ,
         \buff_mem[15][9] , \buff_mem[15][8] , \buff_mem[15][7] ,
         \buff_mem[15][6] , \buff_mem[15][5] , \buff_mem[15][4] ,
         \buff_mem[15][3] , \buff_mem[15][2] , \buff_mem[15][1] ,
         \buff_mem[15][0] , \buff_mem[14][19] , \buff_mem[14][18] ,
         \buff_mem[14][17] , \buff_mem[14][16] , \buff_mem[14][15] ,
         \buff_mem[14][14] , \buff_mem[14][13] , \buff_mem[14][12] ,
         \buff_mem[14][11] , \buff_mem[14][10] , \buff_mem[14][9] ,
         \buff_mem[14][8] , \buff_mem[14][7] , \buff_mem[14][6] ,
         \buff_mem[14][5] , \buff_mem[14][4] , \buff_mem[14][3] ,
         \buff_mem[14][2] , \buff_mem[14][1] , \buff_mem[14][0] ,
         \buff_mem[13][19] , \buff_mem[13][18] , \buff_mem[13][17] ,
         \buff_mem[13][16] , \buff_mem[13][15] , \buff_mem[13][14] ,
         \buff_mem[13][13] , \buff_mem[13][12] , \buff_mem[13][11] ,
         \buff_mem[13][10] , \buff_mem[13][9] , \buff_mem[13][8] ,
         \buff_mem[13][7] , \buff_mem[13][6] , \buff_mem[13][5] ,
         \buff_mem[13][4] , \buff_mem[13][3] , \buff_mem[13][2] ,
         \buff_mem[13][1] , \buff_mem[13][0] , \buff_mem[12][19] ,
         \buff_mem[12][18] , \buff_mem[12][17] , \buff_mem[12][16] ,
         \buff_mem[12][15] , \buff_mem[12][14] , \buff_mem[12][13] ,
         \buff_mem[12][12] , \buff_mem[12][11] , \buff_mem[12][10] ,
         \buff_mem[12][9] , \buff_mem[12][8] , \buff_mem[12][7] ,
         \buff_mem[12][6] , \buff_mem[12][5] , \buff_mem[12][4] ,
         \buff_mem[12][3] , \buff_mem[12][2] , \buff_mem[12][1] ,
         \buff_mem[12][0] , \buff_mem[11][19] , \buff_mem[11][18] ,
         \buff_mem[11][17] , \buff_mem[11][16] , \buff_mem[11][15] ,
         \buff_mem[11][14] , \buff_mem[11][13] , \buff_mem[11][12] ,
         \buff_mem[11][11] , \buff_mem[11][10] , \buff_mem[11][9] ,
         \buff_mem[11][8] , \buff_mem[11][7] , \buff_mem[11][6] ,
         \buff_mem[11][5] , \buff_mem[11][4] , \buff_mem[11][3] ,
         \buff_mem[11][2] , \buff_mem[11][1] , \buff_mem[11][0] ,
         \buff_mem[10][19] , \buff_mem[10][18] , \buff_mem[10][17] ,
         \buff_mem[10][16] , \buff_mem[10][15] , \buff_mem[10][14] ,
         \buff_mem[10][13] , \buff_mem[10][12] , \buff_mem[10][11] ,
         \buff_mem[10][10] , \buff_mem[10][9] , \buff_mem[10][8] ,
         \buff_mem[10][7] , \buff_mem[10][6] , \buff_mem[10][5] ,
         \buff_mem[10][4] , \buff_mem[10][3] , \buff_mem[10][2] ,
         \buff_mem[10][1] , \buff_mem[10][0] , \buff_mem[9][19] ,
         \buff_mem[9][18] , \buff_mem[9][17] , \buff_mem[9][16] ,
         \buff_mem[9][15] , \buff_mem[9][14] , \buff_mem[9][13] ,
         \buff_mem[9][12] , \buff_mem[9][11] , \buff_mem[9][10] ,
         \buff_mem[9][9] , \buff_mem[9][8] , \buff_mem[9][7] ,
         \buff_mem[9][6] , \buff_mem[9][5] , \buff_mem[9][4] ,
         \buff_mem[9][3] , \buff_mem[9][2] , \buff_mem[9][1] ,
         \buff_mem[9][0] , \buff_mem[8][19] , \buff_mem[8][18] ,
         \buff_mem[8][17] , \buff_mem[8][16] , \buff_mem[8][15] ,
         \buff_mem[8][14] , \buff_mem[8][13] , \buff_mem[8][12] ,
         \buff_mem[8][11] , \buff_mem[8][10] , \buff_mem[8][9] ,
         \buff_mem[8][8] , \buff_mem[8][7] , \buff_mem[8][6] ,
         \buff_mem[8][5] , \buff_mem[8][4] , \buff_mem[8][3] ,
         \buff_mem[8][2] , \buff_mem[8][1] , \buff_mem[8][0] ,
         \buff_mem[7][19] , \buff_mem[7][18] , \buff_mem[7][17] ,
         \buff_mem[7][16] , \buff_mem[7][15] , \buff_mem[7][14] ,
         \buff_mem[7][13] , \buff_mem[7][12] , \buff_mem[7][11] ,
         \buff_mem[7][10] , \buff_mem[7][9] , \buff_mem[7][8] ,
         \buff_mem[7][7] , \buff_mem[7][6] , \buff_mem[7][5] ,
         \buff_mem[7][4] , \buff_mem[7][3] , \buff_mem[7][2] ,
         \buff_mem[7][1] , \buff_mem[7][0] , \buff_mem[6][19] ,
         \buff_mem[6][18] , \buff_mem[6][17] , \buff_mem[6][16] ,
         \buff_mem[6][15] , \buff_mem[6][14] , \buff_mem[6][13] ,
         \buff_mem[6][12] , \buff_mem[6][11] , \buff_mem[6][10] ,
         \buff_mem[6][9] , \buff_mem[6][8] , \buff_mem[6][7] ,
         \buff_mem[6][6] , \buff_mem[6][5] , \buff_mem[6][4] ,
         \buff_mem[6][3] , \buff_mem[6][2] , \buff_mem[6][1] ,
         \buff_mem[6][0] , \buff_mem[5][19] , \buff_mem[5][18] ,
         \buff_mem[5][17] , \buff_mem[5][16] , \buff_mem[5][15] ,
         \buff_mem[5][14] , \buff_mem[5][13] , \buff_mem[5][12] ,
         \buff_mem[5][11] , \buff_mem[5][10] , \buff_mem[5][9] ,
         \buff_mem[5][8] , \buff_mem[5][7] , \buff_mem[5][6] ,
         \buff_mem[5][5] , \buff_mem[5][4] , \buff_mem[5][3] ,
         \buff_mem[5][2] , \buff_mem[5][1] , \buff_mem[5][0] ,
         \buff_mem[4][19] , \buff_mem[4][18] , \buff_mem[4][17] ,
         \buff_mem[4][16] , \buff_mem[4][15] , \buff_mem[4][14] ,
         \buff_mem[4][13] , \buff_mem[4][12] , \buff_mem[4][11] ,
         \buff_mem[4][10] , \buff_mem[4][9] , \buff_mem[4][8] ,
         \buff_mem[4][7] , \buff_mem[4][6] , \buff_mem[4][5] ,
         \buff_mem[4][4] , \buff_mem[4][3] , \buff_mem[4][2] ,
         \buff_mem[4][1] , \buff_mem[4][0] , \buff_mem[3][19] ,
         \buff_mem[3][18] , \buff_mem[3][17] , \buff_mem[3][16] ,
         \buff_mem[3][15] , \buff_mem[3][14] , \buff_mem[3][13] ,
         \buff_mem[3][12] , \buff_mem[3][11] , \buff_mem[3][10] ,
         \buff_mem[3][9] , \buff_mem[3][8] , \buff_mem[3][7] ,
         \buff_mem[3][6] , \buff_mem[3][5] , \buff_mem[3][4] ,
         \buff_mem[3][3] , \buff_mem[3][2] , \buff_mem[3][1] ,
         \buff_mem[3][0] , \buff_mem[2][19] , \buff_mem[2][18] ,
         \buff_mem[2][17] , \buff_mem[2][16] , \buff_mem[2][15] ,
         \buff_mem[2][14] , \buff_mem[2][13] , \buff_mem[2][12] ,
         \buff_mem[2][11] , \buff_mem[2][10] , \buff_mem[2][9] ,
         \buff_mem[2][8] , \buff_mem[2][7] , \buff_mem[2][6] ,
         \buff_mem[2][5] , \buff_mem[2][4] , \buff_mem[2][3] ,
         \buff_mem[2][2] , \buff_mem[2][1] , \buff_mem[2][0] ,
         \buff_mem[1][19] , \buff_mem[1][18] , \buff_mem[1][17] ,
         \buff_mem[1][16] , \buff_mem[1][15] , \buff_mem[1][14] ,
         \buff_mem[1][13] , \buff_mem[1][12] , \buff_mem[1][11] ,
         \buff_mem[1][10] , \buff_mem[1][9] , \buff_mem[1][8] ,
         \buff_mem[1][7] , \buff_mem[1][6] , \buff_mem[1][5] ,
         \buff_mem[1][4] , \buff_mem[1][3] , \buff_mem[1][2] ,
         \buff_mem[1][1] , \buff_mem[1][0] , \buff_mem[0][19] ,
         \buff_mem[0][18] , \buff_mem[0][17] , \buff_mem[0][16] ,
         \buff_mem[0][15] , \buff_mem[0][14] , \buff_mem[0][13] ,
         \buff_mem[0][12] , \buff_mem[0][11] , \buff_mem[0][10] ,
         \buff_mem[0][9] , \buff_mem[0][8] , \buff_mem[0][7] ,
         \buff_mem[0][6] , \buff_mem[0][5] , \buff_mem[0][4] ,
         \buff_mem[0][3] , \buff_mem[0][2] , \buff_mem[0][1] ,
         \buff_mem[0][0] , N142, N143, N144, N145, N146, N147, N148, N149,
         N150, N151, N152, N153, N154, N155, N156, N157, N158, N159, N160,
         N161, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n3235, n3236, n3258, n3260, n3261, n3262, n3263,
         n3266, n3269, n3272, n3273, n3275, n3276, n3277, n3278, n3282, n3286,
         n3287, n3288, n3290, n3311, n3333, n3334, n3335, n3336, n3337, n3338,
         n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348,
         n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3358, n3359,
         n3360, n3361, n3362, n3366, n3371, n3373, n3374, n3375, n3376, n3377,
         n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387,
         n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397,
         n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407,
         n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417,
         n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427,
         n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437,
         n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447,
         n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457,
         n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467,
         n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477,
         n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487,
         n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497,
         n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507,
         n3508, n3509, n3510, n3511, n3512, n3514, n3515, n3517, n3518, n3519,
         n3520, n3521, n3522, n3524, n3525, n3526, n3527, n3528, n3530, n3531,
         n3533, n3534, n3536, n3537, n3539, n3540, n3541, n3542, n3543, n3545,
         n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3554, n3555, n3557,
         n3558, n3560, n3561, n3563, n3564, n3566, n3567, n3569, n3570, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3580, n3581, n3582, n3583,
         n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593,
         n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603,
         n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613,
         n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623,
         n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633,
         n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643,
         n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653,
         n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3664,
         n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674,
         n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684,
         n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694,
         n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704,
         n3705, n3706, n3707, n3709, n3710, n3711, n3712, n3713, n3714, n3715,
         n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725,
         n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735,
         n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745,
         n3746, n3747, n3748, n3749, n3751, n3752, n3753, n3754, n3755, n3756,
         n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766,
         n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776,
         n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786,
         n3787, n3788, n3789, n3790, n3791, n3793, n3794, n3795, n3796, n3797,
         n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807,
         n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817,
         n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827,
         n3828, n3829, n3830, n3831, n3832, n3833, n3835, n3836, n3837, n3838,
         n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848,
         n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858,
         n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868,
         n3869, n3870, n3871, n3872, n3873, n3875, n3876, n3877, n3879, n3880,
         n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890,
         n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900,
         n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910,
         n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920,
         n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930,
         n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940,
         n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950,
         n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960,
         n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970,
         n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980,
         n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990,
         n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000,
         n4001, n4002, n4003, n4005, n4006, n4007, n4008, n4009, n4010, n4011,
         n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021,
         n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031,
         n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041,
         n4042, n4043, n4044, n4045, n4046, n4047, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4091, n4092, n4093,
         n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103,
         n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113,
         n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123,
         n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4133, n4134,
         n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144,
         n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154,
         n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164,
         n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4175,
         n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185,
         n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195,
         n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205,
         n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4215, n4216,
         n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226,
         n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236,
         n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246,
         n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256,
         n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266,
         n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276,
         n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286,
         n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296,
         n4297, n4298, n4299, n4300, n4301, n4303, n4304, n4305, n4306, n4307,
         n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317,
         n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327,
         n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337,
         n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347,
         n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357,
         n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367,
         n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377,
         n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387,
         n4388, n4389, n4390, n4392, n4393, n4394, n4395, n4396, n4397, n4398,
         n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408,
         n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4418, n4419,
         n4420, n4422, n4423, n4426, n4427, n4428, n4429, n4432, n4433, n4434,
         n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4445,
         n4446, n4448, n4449, n4450, n4453, n4454, n4455, n4456, n4458, n4459,
         n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469,
         n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479,
         n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489,
         n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499,
         n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509,
         n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519,
         n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529,
         n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539,
         n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549,
         n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559,
         n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569,
         n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579,
         n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589,
         n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599,
         n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609,
         n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619,
         n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629,
         n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639,
         n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649,
         n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659,
         n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669,
         n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679,
         n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689,
         n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699,
         n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709,
         n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719,
         n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729,
         n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739,
         n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749,
         n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759,
         n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769,
         n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779,
         n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789,
         n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799,
         n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809,
         n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819,
         n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829,
         n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839,
         n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849,
         n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859,
         n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869,
         n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879,
         n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889,
         n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899,
         n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909,
         n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919,
         n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929,
         n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939,
         n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949,
         n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959,
         n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969,
         n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979,
         n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989,
         n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999,
         n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009,
         n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019,
         n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029,
         n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039,
         n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049,
         n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059,
         n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069,
         n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079,
         n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089,
         n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099,
         n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109,
         n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119,
         n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129,
         n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139,
         n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149,
         n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159,
         n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169,
         n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179,
         n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189,
         n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199,
         n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209,
         n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219,
         n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229,
         n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239,
         n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249,
         n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259,
         n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269,
         n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279,
         n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289,
         n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299,
         n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309,
         n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319,
         n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329,
         n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339,
         n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349,
         n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359,
         n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369,
         n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379,
         n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389,
         n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399,
         n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409,
         n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419,
         n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429,
         n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439,
         n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449,
         n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459,
         n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469,
         n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479,
         n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489,
         n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499,
         n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509,
         n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519,
         n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529,
         n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539,
         n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549,
         n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559,
         n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569,
         n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579,
         n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589,
         n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599,
         n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609,
         n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619,
         n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629,
         n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639,
         n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649,
         n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659,
         n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669,
         n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679,
         n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689,
         n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699,
         n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709,
         n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719,
         n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729,
         n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739,
         n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749,
         n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759,
         n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769,
         n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779,
         n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789,
         n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799,
         n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809,
         n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819,
         n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829,
         n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839,
         n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849,
         n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859,
         n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869,
         n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879,
         n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889,
         n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899,
         n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909,
         n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919,
         n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929,
         n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939,
         n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949,
         n5950, n5951, n5952, n5953, n5954, n5955, n5956;
  wire   [4:0] rd_ptr;
  wire   [4:0] wr_ptr;

  dff_sg \rd_ptr_reg[0]  ( .D(n2375), .CP(clk), .Q(rd_ptr[0]) );
  dff_sg full_reg ( .D(n2374), .CP(clk), .Q(full) );
  dff_sg \wr_ptr_reg[0]  ( .D(n2373), .CP(clk), .Q(wr_ptr[0]) );
  dff_sg \wr_ptr_reg[1]  ( .D(n2372), .CP(clk), .Q(wr_ptr[1]) );
  dff_sg \wr_ptr_reg[2]  ( .D(n2371), .CP(clk), .Q(wr_ptr[2]) );
  dff_sg \wr_ptr_reg[3]  ( .D(n2370), .CP(clk), .Q(wr_ptr[3]) );
  dff_sg \wr_ptr_reg[4]  ( .D(n2369), .CP(clk), .Q(wr_ptr[4]) );
  dff_sg empty_reg ( .D(n2368), .CP(clk), .Q(empty) );
  dff_sg \rd_ptr_reg[1]  ( .D(n1967), .CP(clk), .Q(rd_ptr[1]) );
  dff_sg \rd_ptr_reg[2]  ( .D(n1966), .CP(clk), .Q(rd_ptr[2]) );
  dff_sg \rd_ptr_reg[3]  ( .D(n1965), .CP(clk), .Q(rd_ptr[3]) );
  dff_sg \rd_ptr_reg[4]  ( .D(n1964), .CP(clk), .Q(rd_ptr[4]) );
  dff_sg \buff_mem_reg[3][13]  ( .D(n2294), .CP(clk), .Q(\buff_mem[3][13] ) );
  dff_sg \buff_mem_reg[2][13]  ( .D(n2314), .CP(clk), .Q(\buff_mem[2][13] ) );
  dff_sg \buff_mem_reg[1][13]  ( .D(n2334), .CP(clk), .Q(\buff_mem[1][13] ) );
  dff_sg \buff_mem_reg[0][13]  ( .D(n2354), .CP(clk), .Q(\buff_mem[0][13] ) );
  dff_sg \buff_mem_reg[19][13]  ( .D(n1974), .CP(clk), .Q(\buff_mem[19][13] )
         );
  dff_sg \buff_mem_reg[18][13]  ( .D(n1994), .CP(clk), .Q(\buff_mem[18][13] )
         );
  dff_sg \buff_mem_reg[17][13]  ( .D(n2014), .CP(clk), .Q(\buff_mem[17][13] )
         );
  dff_sg \buff_mem_reg[16][13]  ( .D(n2034), .CP(clk), .Q(\buff_mem[16][13] )
         );
  dff_sg \buff_mem_reg[11][13]  ( .D(n2134), .CP(clk), .Q(\buff_mem[11][13] )
         );
  dff_sg \buff_mem_reg[10][13]  ( .D(n2154), .CP(clk), .Q(\buff_mem[10][13] )
         );
  dff_sg \buff_mem_reg[9][13]  ( .D(n2174), .CP(clk), .Q(\buff_mem[9][13] ) );
  dff_sg \buff_mem_reg[8][13]  ( .D(n2194), .CP(clk), .Q(\buff_mem[8][13] ) );
  dff_sg \buff_mem_reg[3][12]  ( .D(n2295), .CP(clk), .Q(\buff_mem[3][12] ) );
  dff_sg \buff_mem_reg[2][12]  ( .D(n2315), .CP(clk), .Q(\buff_mem[2][12] ) );
  dff_sg \buff_mem_reg[1][12]  ( .D(n2335), .CP(clk), .Q(\buff_mem[1][12] ) );
  dff_sg \buff_mem_reg[0][12]  ( .D(n2355), .CP(clk), .Q(\buff_mem[0][12] ) );
  dff_sg \buff_mem_reg[19][12]  ( .D(n1975), .CP(clk), .Q(\buff_mem[19][12] )
         );
  dff_sg \buff_mem_reg[18][12]  ( .D(n1995), .CP(clk), .Q(\buff_mem[18][12] )
         );
  dff_sg \buff_mem_reg[17][12]  ( .D(n2015), .CP(clk), .Q(\buff_mem[17][12] )
         );
  dff_sg \buff_mem_reg[16][12]  ( .D(n2035), .CP(clk), .Q(\buff_mem[16][12] )
         );
  dff_sg \buff_mem_reg[11][12]  ( .D(n2135), .CP(clk), .Q(\buff_mem[11][12] )
         );
  dff_sg \buff_mem_reg[10][12]  ( .D(n2155), .CP(clk), .Q(\buff_mem[10][12] )
         );
  dff_sg \buff_mem_reg[9][12]  ( .D(n2175), .CP(clk), .Q(\buff_mem[9][12] ) );
  dff_sg \buff_mem_reg[8][12]  ( .D(n2195), .CP(clk), .Q(\buff_mem[8][12] ) );
  dff_sg \buff_mem_reg[3][11]  ( .D(n2296), .CP(clk), .Q(\buff_mem[3][11] ) );
  dff_sg \buff_mem_reg[2][11]  ( .D(n2316), .CP(clk), .Q(\buff_mem[2][11] ) );
  dff_sg \buff_mem_reg[1][11]  ( .D(n2336), .CP(clk), .Q(\buff_mem[1][11] ) );
  dff_sg \buff_mem_reg[0][11]  ( .D(n2356), .CP(clk), .Q(\buff_mem[0][11] ) );
  dff_sg \buff_mem_reg[19][11]  ( .D(n1976), .CP(clk), .Q(\buff_mem[19][11] )
         );
  dff_sg \buff_mem_reg[18][11]  ( .D(n1996), .CP(clk), .Q(\buff_mem[18][11] )
         );
  dff_sg \buff_mem_reg[17][11]  ( .D(n2016), .CP(clk), .Q(\buff_mem[17][11] )
         );
  dff_sg \buff_mem_reg[16][11]  ( .D(n2036), .CP(clk), .Q(\buff_mem[16][11] )
         );
  dff_sg \buff_mem_reg[11][11]  ( .D(n2136), .CP(clk), .Q(\buff_mem[11][11] )
         );
  dff_sg \buff_mem_reg[10][11]  ( .D(n2156), .CP(clk), .Q(\buff_mem[10][11] )
         );
  dff_sg \buff_mem_reg[9][11]  ( .D(n2176), .CP(clk), .Q(\buff_mem[9][11] ) );
  dff_sg \buff_mem_reg[8][11]  ( .D(n2196), .CP(clk), .Q(\buff_mem[8][11] ) );
  dff_sg \buff_mem_reg[3][10]  ( .D(n2297), .CP(clk), .Q(\buff_mem[3][10] ) );
  dff_sg \buff_mem_reg[2][10]  ( .D(n2317), .CP(clk), .Q(\buff_mem[2][10] ) );
  dff_sg \buff_mem_reg[1][10]  ( .D(n2337), .CP(clk), .Q(\buff_mem[1][10] ) );
  dff_sg \buff_mem_reg[0][10]  ( .D(n2357), .CP(clk), .Q(\buff_mem[0][10] ) );
  dff_sg \buff_mem_reg[19][10]  ( .D(n1977), .CP(clk), .Q(\buff_mem[19][10] )
         );
  dff_sg \buff_mem_reg[18][10]  ( .D(n1997), .CP(clk), .Q(\buff_mem[18][10] )
         );
  dff_sg \buff_mem_reg[17][10]  ( .D(n2017), .CP(clk), .Q(\buff_mem[17][10] )
         );
  dff_sg \buff_mem_reg[16][10]  ( .D(n2037), .CP(clk), .Q(\buff_mem[16][10] )
         );
  dff_sg \buff_mem_reg[11][10]  ( .D(n2137), .CP(clk), .Q(\buff_mem[11][10] )
         );
  dff_sg \buff_mem_reg[10][10]  ( .D(n2157), .CP(clk), .Q(\buff_mem[10][10] )
         );
  dff_sg \buff_mem_reg[9][10]  ( .D(n2177), .CP(clk), .Q(\buff_mem[9][10] ) );
  dff_sg \buff_mem_reg[8][10]  ( .D(n2197), .CP(clk), .Q(\buff_mem[8][10] ) );
  dff_sg \buff_mem_reg[3][9]  ( .D(n2298), .CP(clk), .Q(\buff_mem[3][9] ) );
  dff_sg \buff_mem_reg[2][9]  ( .D(n2318), .CP(clk), .Q(\buff_mem[2][9] ) );
  dff_sg \buff_mem_reg[1][9]  ( .D(n2338), .CP(clk), .Q(\buff_mem[1][9] ) );
  dff_sg \buff_mem_reg[0][9]  ( .D(n2358), .CP(clk), .Q(\buff_mem[0][9] ) );
  dff_sg \buff_mem_reg[19][9]  ( .D(n1978), .CP(clk), .Q(\buff_mem[19][9] ) );
  dff_sg \buff_mem_reg[18][9]  ( .D(n1998), .CP(clk), .Q(\buff_mem[18][9] ) );
  dff_sg \buff_mem_reg[17][9]  ( .D(n2018), .CP(clk), .Q(\buff_mem[17][9] ) );
  dff_sg \buff_mem_reg[16][9]  ( .D(n2038), .CP(clk), .Q(\buff_mem[16][9] ) );
  dff_sg \buff_mem_reg[11][9]  ( .D(n2138), .CP(clk), .Q(\buff_mem[11][9] ) );
  dff_sg \buff_mem_reg[10][9]  ( .D(n2158), .CP(clk), .Q(\buff_mem[10][9] ) );
  dff_sg \buff_mem_reg[9][9]  ( .D(n2178), .CP(clk), .Q(\buff_mem[9][9] ) );
  dff_sg \buff_mem_reg[8][9]  ( .D(n2198), .CP(clk), .Q(\buff_mem[8][9] ) );
  dff_sg \buff_mem_reg[3][8]  ( .D(n2299), .CP(clk), .Q(\buff_mem[3][8] ) );
  dff_sg \buff_mem_reg[2][8]  ( .D(n2319), .CP(clk), .Q(\buff_mem[2][8] ) );
  dff_sg \buff_mem_reg[1][8]  ( .D(n2339), .CP(clk), .Q(\buff_mem[1][8] ) );
  dff_sg \buff_mem_reg[0][8]  ( .D(n2359), .CP(clk), .Q(\buff_mem[0][8] ) );
  dff_sg \buff_mem_reg[19][8]  ( .D(n1979), .CP(clk), .Q(\buff_mem[19][8] ) );
  dff_sg \buff_mem_reg[18][8]  ( .D(n1999), .CP(clk), .Q(\buff_mem[18][8] ) );
  dff_sg \buff_mem_reg[17][8]  ( .D(n2019), .CP(clk), .Q(\buff_mem[17][8] ) );
  dff_sg \buff_mem_reg[16][8]  ( .D(n2039), .CP(clk), .Q(\buff_mem[16][8] ) );
  dff_sg \buff_mem_reg[11][8]  ( .D(n2139), .CP(clk), .Q(\buff_mem[11][8] ) );
  dff_sg \buff_mem_reg[10][8]  ( .D(n2159), .CP(clk), .Q(\buff_mem[10][8] ) );
  dff_sg \buff_mem_reg[9][8]  ( .D(n2179), .CP(clk), .Q(\buff_mem[9][8] ) );
  dff_sg \buff_mem_reg[8][8]  ( .D(n2199), .CP(clk), .Q(\buff_mem[8][8] ) );
  dff_sg \buff_mem_reg[3][7]  ( .D(n2300), .CP(clk), .Q(\buff_mem[3][7] ) );
  dff_sg \buff_mem_reg[2][7]  ( .D(n2320), .CP(clk), .Q(\buff_mem[2][7] ) );
  dff_sg \buff_mem_reg[1][7]  ( .D(n2340), .CP(clk), .Q(\buff_mem[1][7] ) );
  dff_sg \buff_mem_reg[0][7]  ( .D(n2360), .CP(clk), .Q(\buff_mem[0][7] ) );
  dff_sg \buff_mem_reg[19][7]  ( .D(n1980), .CP(clk), .Q(\buff_mem[19][7] ) );
  dff_sg \buff_mem_reg[18][7]  ( .D(n2000), .CP(clk), .Q(\buff_mem[18][7] ) );
  dff_sg \buff_mem_reg[17][7]  ( .D(n2020), .CP(clk), .Q(\buff_mem[17][7] ) );
  dff_sg \buff_mem_reg[16][7]  ( .D(n2040), .CP(clk), .Q(\buff_mem[16][7] ) );
  dff_sg \buff_mem_reg[11][7]  ( .D(n2140), .CP(clk), .Q(\buff_mem[11][7] ) );
  dff_sg \buff_mem_reg[10][7]  ( .D(n2160), .CP(clk), .Q(\buff_mem[10][7] ) );
  dff_sg \buff_mem_reg[9][7]  ( .D(n2180), .CP(clk), .Q(\buff_mem[9][7] ) );
  dff_sg \buff_mem_reg[8][7]  ( .D(n2200), .CP(clk), .Q(\buff_mem[8][7] ) );
  dff_sg \buff_mem_reg[3][6]  ( .D(n2301), .CP(clk), .Q(\buff_mem[3][6] ) );
  dff_sg \buff_mem_reg[2][6]  ( .D(n2321), .CP(clk), .Q(\buff_mem[2][6] ) );
  dff_sg \buff_mem_reg[1][6]  ( .D(n2341), .CP(clk), .Q(\buff_mem[1][6] ) );
  dff_sg \buff_mem_reg[0][6]  ( .D(n2361), .CP(clk), .Q(\buff_mem[0][6] ) );
  dff_sg \buff_mem_reg[19][6]  ( .D(n1981), .CP(clk), .Q(\buff_mem[19][6] ) );
  dff_sg \buff_mem_reg[18][6]  ( .D(n2001), .CP(clk), .Q(\buff_mem[18][6] ) );
  dff_sg \buff_mem_reg[17][6]  ( .D(n2021), .CP(clk), .Q(\buff_mem[17][6] ) );
  dff_sg \buff_mem_reg[16][6]  ( .D(n2041), .CP(clk), .Q(\buff_mem[16][6] ) );
  dff_sg \buff_mem_reg[11][6]  ( .D(n2141), .CP(clk), .Q(\buff_mem[11][6] ) );
  dff_sg \buff_mem_reg[10][6]  ( .D(n2161), .CP(clk), .Q(\buff_mem[10][6] ) );
  dff_sg \buff_mem_reg[9][6]  ( .D(n2181), .CP(clk), .Q(\buff_mem[9][6] ) );
  dff_sg \buff_mem_reg[8][6]  ( .D(n2201), .CP(clk), .Q(\buff_mem[8][6] ) );
  dff_sg \buff_mem_reg[3][5]  ( .D(n2302), .CP(clk), .Q(\buff_mem[3][5] ) );
  dff_sg \buff_mem_reg[2][5]  ( .D(n2322), .CP(clk), .Q(\buff_mem[2][5] ) );
  dff_sg \buff_mem_reg[1][5]  ( .D(n2342), .CP(clk), .Q(\buff_mem[1][5] ) );
  dff_sg \buff_mem_reg[0][5]  ( .D(n2362), .CP(clk), .Q(\buff_mem[0][5] ) );
  dff_sg \buff_mem_reg[19][5]  ( .D(n1982), .CP(clk), .Q(\buff_mem[19][5] ) );
  dff_sg \buff_mem_reg[18][5]  ( .D(n2002), .CP(clk), .Q(\buff_mem[18][5] ) );
  dff_sg \buff_mem_reg[17][5]  ( .D(n2022), .CP(clk), .Q(\buff_mem[17][5] ) );
  dff_sg \buff_mem_reg[16][5]  ( .D(n2042), .CP(clk), .Q(\buff_mem[16][5] ) );
  dff_sg \buff_mem_reg[11][5]  ( .D(n2142), .CP(clk), .Q(\buff_mem[11][5] ) );
  dff_sg \buff_mem_reg[10][5]  ( .D(n2162), .CP(clk), .Q(\buff_mem[10][5] ) );
  dff_sg \buff_mem_reg[9][5]  ( .D(n2182), .CP(clk), .Q(\buff_mem[9][5] ) );
  dff_sg \buff_mem_reg[8][5]  ( .D(n2202), .CP(clk), .Q(\buff_mem[8][5] ) );
  dff_sg \buff_mem_reg[3][4]  ( .D(n2303), .CP(clk), .Q(\buff_mem[3][4] ) );
  dff_sg \buff_mem_reg[2][4]  ( .D(n2323), .CP(clk), .Q(\buff_mem[2][4] ) );
  dff_sg \buff_mem_reg[1][4]  ( .D(n2343), .CP(clk), .Q(\buff_mem[1][4] ) );
  dff_sg \buff_mem_reg[0][4]  ( .D(n2363), .CP(clk), .Q(\buff_mem[0][4] ) );
  dff_sg \buff_mem_reg[19][4]  ( .D(n1983), .CP(clk), .Q(\buff_mem[19][4] ) );
  dff_sg \buff_mem_reg[18][4]  ( .D(n2003), .CP(clk), .Q(\buff_mem[18][4] ) );
  dff_sg \buff_mem_reg[17][4]  ( .D(n2023), .CP(clk), .Q(\buff_mem[17][4] ) );
  dff_sg \buff_mem_reg[16][4]  ( .D(n2043), .CP(clk), .Q(\buff_mem[16][4] ) );
  dff_sg \buff_mem_reg[11][4]  ( .D(n2143), .CP(clk), .Q(\buff_mem[11][4] ) );
  dff_sg \buff_mem_reg[10][4]  ( .D(n2163), .CP(clk), .Q(\buff_mem[10][4] ) );
  dff_sg \buff_mem_reg[9][4]  ( .D(n2183), .CP(clk), .Q(\buff_mem[9][4] ) );
  dff_sg \buff_mem_reg[8][4]  ( .D(n2203), .CP(clk), .Q(\buff_mem[8][4] ) );
  dff_sg \buff_mem_reg[3][3]  ( .D(n2304), .CP(clk), .Q(\buff_mem[3][3] ) );
  dff_sg \buff_mem_reg[2][3]  ( .D(n2324), .CP(clk), .Q(\buff_mem[2][3] ) );
  dff_sg \buff_mem_reg[1][3]  ( .D(n2344), .CP(clk), .Q(\buff_mem[1][3] ) );
  dff_sg \buff_mem_reg[0][3]  ( .D(n2364), .CP(clk), .Q(\buff_mem[0][3] ) );
  dff_sg \buff_mem_reg[19][3]  ( .D(n1984), .CP(clk), .Q(\buff_mem[19][3] ) );
  dff_sg \buff_mem_reg[18][3]  ( .D(n2004), .CP(clk), .Q(\buff_mem[18][3] ) );
  dff_sg \buff_mem_reg[17][3]  ( .D(n2024), .CP(clk), .Q(\buff_mem[17][3] ) );
  dff_sg \buff_mem_reg[16][3]  ( .D(n2044), .CP(clk), .Q(\buff_mem[16][3] ) );
  dff_sg \buff_mem_reg[11][3]  ( .D(n2144), .CP(clk), .Q(\buff_mem[11][3] ) );
  dff_sg \buff_mem_reg[10][3]  ( .D(n2164), .CP(clk), .Q(\buff_mem[10][3] ) );
  dff_sg \buff_mem_reg[9][3]  ( .D(n2184), .CP(clk), .Q(\buff_mem[9][3] ) );
  dff_sg \buff_mem_reg[8][3]  ( .D(n2204), .CP(clk), .Q(\buff_mem[8][3] ) );
  dff_sg \buff_mem_reg[3][2]  ( .D(n2305), .CP(clk), .Q(\buff_mem[3][2] ) );
  dff_sg \buff_mem_reg[2][2]  ( .D(n2325), .CP(clk), .Q(\buff_mem[2][2] ) );
  dff_sg \buff_mem_reg[1][2]  ( .D(n2345), .CP(clk), .Q(\buff_mem[1][2] ) );
  dff_sg \buff_mem_reg[0][2]  ( .D(n2365), .CP(clk), .Q(\buff_mem[0][2] ) );
  dff_sg \buff_mem_reg[19][2]  ( .D(n1985), .CP(clk), .Q(\buff_mem[19][2] ) );
  dff_sg \buff_mem_reg[18][2]  ( .D(n2005), .CP(clk), .Q(\buff_mem[18][2] ) );
  dff_sg \buff_mem_reg[17][2]  ( .D(n2025), .CP(clk), .Q(\buff_mem[17][2] ) );
  dff_sg \buff_mem_reg[16][2]  ( .D(n2045), .CP(clk), .Q(\buff_mem[16][2] ) );
  dff_sg \buff_mem_reg[11][2]  ( .D(n2145), .CP(clk), .Q(\buff_mem[11][2] ) );
  dff_sg \buff_mem_reg[10][2]  ( .D(n2165), .CP(clk), .Q(\buff_mem[10][2] ) );
  dff_sg \buff_mem_reg[9][2]  ( .D(n2185), .CP(clk), .Q(\buff_mem[9][2] ) );
  dff_sg \buff_mem_reg[8][2]  ( .D(n2205), .CP(clk), .Q(\buff_mem[8][2] ) );
  dff_sg \buff_mem_reg[3][1]  ( .D(n2306), .CP(clk), .Q(\buff_mem[3][1] ) );
  dff_sg \buff_mem_reg[2][1]  ( .D(n2326), .CP(clk), .Q(\buff_mem[2][1] ) );
  dff_sg \buff_mem_reg[1][1]  ( .D(n2346), .CP(clk), .Q(\buff_mem[1][1] ) );
  dff_sg \buff_mem_reg[0][1]  ( .D(n2366), .CP(clk), .Q(\buff_mem[0][1] ) );
  dff_sg \buff_mem_reg[19][1]  ( .D(n1986), .CP(clk), .Q(\buff_mem[19][1] ) );
  dff_sg \buff_mem_reg[18][1]  ( .D(n2006), .CP(clk), .Q(\buff_mem[18][1] ) );
  dff_sg \buff_mem_reg[17][1]  ( .D(n2026), .CP(clk), .Q(\buff_mem[17][1] ) );
  dff_sg \buff_mem_reg[16][1]  ( .D(n2046), .CP(clk), .Q(\buff_mem[16][1] ) );
  dff_sg \buff_mem_reg[11][1]  ( .D(n2146), .CP(clk), .Q(\buff_mem[11][1] ) );
  dff_sg \buff_mem_reg[10][1]  ( .D(n2166), .CP(clk), .Q(\buff_mem[10][1] ) );
  dff_sg \buff_mem_reg[9][1]  ( .D(n2186), .CP(clk), .Q(\buff_mem[9][1] ) );
  dff_sg \buff_mem_reg[8][1]  ( .D(n2206), .CP(clk), .Q(\buff_mem[8][1] ) );
  dff_sg \buff_mem_reg[3][0]  ( .D(n2307), .CP(clk), .Q(\buff_mem[3][0] ) );
  dff_sg \buff_mem_reg[2][0]  ( .D(n2327), .CP(clk), .Q(\buff_mem[2][0] ) );
  dff_sg \buff_mem_reg[1][0]  ( .D(n2347), .CP(clk), .Q(\buff_mem[1][0] ) );
  dff_sg \buff_mem_reg[0][0]  ( .D(n2367), .CP(clk), .Q(\buff_mem[0][0] ) );
  dff_sg \buff_mem_reg[19][0]  ( .D(n1987), .CP(clk), .Q(\buff_mem[19][0] ) );
  dff_sg \buff_mem_reg[18][0]  ( .D(n2007), .CP(clk), .Q(\buff_mem[18][0] ) );
  dff_sg \buff_mem_reg[17][0]  ( .D(n2027), .CP(clk), .Q(\buff_mem[17][0] ) );
  dff_sg \buff_mem_reg[16][0]  ( .D(n2047), .CP(clk), .Q(\buff_mem[16][0] ) );
  dff_sg \buff_mem_reg[11][0]  ( .D(n2147), .CP(clk), .Q(\buff_mem[11][0] ) );
  dff_sg \buff_mem_reg[10][0]  ( .D(n2167), .CP(clk), .Q(\buff_mem[10][0] ) );
  dff_sg \buff_mem_reg[9][0]  ( .D(n2187), .CP(clk), .Q(\buff_mem[9][0] ) );
  dff_sg \buff_mem_reg[8][0]  ( .D(n2207), .CP(clk), .Q(\buff_mem[8][0] ) );
  dff_sg \buff_mem_reg[3][19]  ( .D(n2288), .CP(clk), .Q(\buff_mem[3][19] ) );
  dff_sg \buff_mem_reg[2][19]  ( .D(n2308), .CP(clk), .Q(\buff_mem[2][19] ) );
  dff_sg \buff_mem_reg[1][19]  ( .D(n2328), .CP(clk), .Q(\buff_mem[1][19] ) );
  dff_sg \buff_mem_reg[0][19]  ( .D(n2348), .CP(clk), .Q(\buff_mem[0][19] ) );
  dff_sg \buff_mem_reg[19][19]  ( .D(n1968), .CP(clk), .Q(\buff_mem[19][19] )
         );
  dff_sg \buff_mem_reg[18][19]  ( .D(n1988), .CP(clk), .Q(\buff_mem[18][19] )
         );
  dff_sg \buff_mem_reg[17][19]  ( .D(n2008), .CP(clk), .Q(\buff_mem[17][19] )
         );
  dff_sg \buff_mem_reg[16][19]  ( .D(n2028), .CP(clk), .Q(\buff_mem[16][19] )
         );
  dff_sg \buff_mem_reg[11][19]  ( .D(n2128), .CP(clk), .Q(\buff_mem[11][19] )
         );
  dff_sg \buff_mem_reg[10][19]  ( .D(n2148), .CP(clk), .Q(\buff_mem[10][19] )
         );
  dff_sg \buff_mem_reg[9][19]  ( .D(n2168), .CP(clk), .Q(\buff_mem[9][19] ) );
  dff_sg \buff_mem_reg[8][19]  ( .D(n2188), .CP(clk), .Q(\buff_mem[8][19] ) );
  dff_sg \buff_mem_reg[3][18]  ( .D(n2289), .CP(clk), .Q(\buff_mem[3][18] ) );
  dff_sg \buff_mem_reg[2][18]  ( .D(n2309), .CP(clk), .Q(\buff_mem[2][18] ) );
  dff_sg \buff_mem_reg[1][18]  ( .D(n2329), .CP(clk), .Q(\buff_mem[1][18] ) );
  dff_sg \buff_mem_reg[0][18]  ( .D(n2349), .CP(clk), .Q(\buff_mem[0][18] ) );
  dff_sg \buff_mem_reg[19][18]  ( .D(n1969), .CP(clk), .Q(\buff_mem[19][18] )
         );
  dff_sg \buff_mem_reg[18][18]  ( .D(n1989), .CP(clk), .Q(\buff_mem[18][18] )
         );
  dff_sg \buff_mem_reg[17][18]  ( .D(n2009), .CP(clk), .Q(\buff_mem[17][18] )
         );
  dff_sg \buff_mem_reg[16][18]  ( .D(n2029), .CP(clk), .Q(\buff_mem[16][18] )
         );
  dff_sg \buff_mem_reg[11][18]  ( .D(n2129), .CP(clk), .Q(\buff_mem[11][18] )
         );
  dff_sg \buff_mem_reg[10][18]  ( .D(n2149), .CP(clk), .Q(\buff_mem[10][18] )
         );
  dff_sg \buff_mem_reg[9][18]  ( .D(n2169), .CP(clk), .Q(\buff_mem[9][18] ) );
  dff_sg \buff_mem_reg[8][18]  ( .D(n2189), .CP(clk), .Q(\buff_mem[8][18] ) );
  dff_sg \buff_mem_reg[3][17]  ( .D(n2290), .CP(clk), .Q(\buff_mem[3][17] ) );
  dff_sg \buff_mem_reg[2][17]  ( .D(n2310), .CP(clk), .Q(\buff_mem[2][17] ) );
  dff_sg \buff_mem_reg[1][17]  ( .D(n2330), .CP(clk), .Q(\buff_mem[1][17] ) );
  dff_sg \buff_mem_reg[0][17]  ( .D(n2350), .CP(clk), .Q(\buff_mem[0][17] ) );
  dff_sg \buff_mem_reg[19][17]  ( .D(n1970), .CP(clk), .Q(\buff_mem[19][17] )
         );
  dff_sg \buff_mem_reg[18][17]  ( .D(n1990), .CP(clk), .Q(\buff_mem[18][17] )
         );
  dff_sg \buff_mem_reg[17][17]  ( .D(n2010), .CP(clk), .Q(\buff_mem[17][17] )
         );
  dff_sg \buff_mem_reg[16][17]  ( .D(n2030), .CP(clk), .Q(\buff_mem[16][17] )
         );
  dff_sg \buff_mem_reg[11][17]  ( .D(n2130), .CP(clk), .Q(\buff_mem[11][17] )
         );
  dff_sg \buff_mem_reg[10][17]  ( .D(n2150), .CP(clk), .Q(\buff_mem[10][17] )
         );
  dff_sg \buff_mem_reg[9][17]  ( .D(n2170), .CP(clk), .Q(\buff_mem[9][17] ) );
  dff_sg \buff_mem_reg[8][17]  ( .D(n2190), .CP(clk), .Q(\buff_mem[8][17] ) );
  dff_sg \buff_mem_reg[3][16]  ( .D(n2291), .CP(clk), .Q(\buff_mem[3][16] ) );
  dff_sg \buff_mem_reg[2][16]  ( .D(n2311), .CP(clk), .Q(\buff_mem[2][16] ) );
  dff_sg \buff_mem_reg[1][16]  ( .D(n2331), .CP(clk), .Q(\buff_mem[1][16] ) );
  dff_sg \buff_mem_reg[0][16]  ( .D(n2351), .CP(clk), .Q(\buff_mem[0][16] ) );
  dff_sg \buff_mem_reg[19][16]  ( .D(n1971), .CP(clk), .Q(\buff_mem[19][16] )
         );
  dff_sg \buff_mem_reg[18][16]  ( .D(n1991), .CP(clk), .Q(\buff_mem[18][16] )
         );
  dff_sg \buff_mem_reg[17][16]  ( .D(n2011), .CP(clk), .Q(\buff_mem[17][16] )
         );
  dff_sg \buff_mem_reg[16][16]  ( .D(n2031), .CP(clk), .Q(\buff_mem[16][16] )
         );
  dff_sg \buff_mem_reg[11][16]  ( .D(n2131), .CP(clk), .Q(\buff_mem[11][16] )
         );
  dff_sg \buff_mem_reg[10][16]  ( .D(n2151), .CP(clk), .Q(\buff_mem[10][16] )
         );
  dff_sg \buff_mem_reg[9][16]  ( .D(n2171), .CP(clk), .Q(\buff_mem[9][16] ) );
  dff_sg \buff_mem_reg[8][16]  ( .D(n2191), .CP(clk), .Q(\buff_mem[8][16] ) );
  dff_sg \buff_mem_reg[3][15]  ( .D(n2292), .CP(clk), .Q(\buff_mem[3][15] ) );
  dff_sg \buff_mem_reg[2][15]  ( .D(n2312), .CP(clk), .Q(\buff_mem[2][15] ) );
  dff_sg \buff_mem_reg[1][15]  ( .D(n2332), .CP(clk), .Q(\buff_mem[1][15] ) );
  dff_sg \buff_mem_reg[0][15]  ( .D(n2352), .CP(clk), .Q(\buff_mem[0][15] ) );
  dff_sg \buff_mem_reg[19][15]  ( .D(n1972), .CP(clk), .Q(\buff_mem[19][15] )
         );
  dff_sg \buff_mem_reg[18][15]  ( .D(n1992), .CP(clk), .Q(\buff_mem[18][15] )
         );
  dff_sg \buff_mem_reg[17][15]  ( .D(n2012), .CP(clk), .Q(\buff_mem[17][15] )
         );
  dff_sg \buff_mem_reg[16][15]  ( .D(n2032), .CP(clk), .Q(\buff_mem[16][15] )
         );
  dff_sg \buff_mem_reg[11][15]  ( .D(n2132), .CP(clk), .Q(\buff_mem[11][15] )
         );
  dff_sg \buff_mem_reg[10][15]  ( .D(n2152), .CP(clk), .Q(\buff_mem[10][15] )
         );
  dff_sg \buff_mem_reg[9][15]  ( .D(n2172), .CP(clk), .Q(\buff_mem[9][15] ) );
  dff_sg \buff_mem_reg[8][15]  ( .D(n2192), .CP(clk), .Q(\buff_mem[8][15] ) );
  dff_sg \buff_mem_reg[15][19]  ( .D(n2048), .CP(clk), .Q(\buff_mem[15][19] )
         );
  dff_sg \buff_mem_reg[15][18]  ( .D(n2049), .CP(clk), .Q(\buff_mem[15][18] )
         );
  dff_sg \buff_mem_reg[15][17]  ( .D(n2050), .CP(clk), .Q(\buff_mem[15][17] )
         );
  dff_sg \buff_mem_reg[15][16]  ( .D(n2051), .CP(clk), .Q(\buff_mem[15][16] )
         );
  dff_sg \buff_mem_reg[15][15]  ( .D(n2052), .CP(clk), .Q(\buff_mem[15][15] )
         );
  dff_sg \buff_mem_reg[15][13]  ( .D(n2054), .CP(clk), .Q(\buff_mem[15][13] )
         );
  dff_sg \buff_mem_reg[15][12]  ( .D(n2055), .CP(clk), .Q(\buff_mem[15][12] )
         );
  dff_sg \buff_mem_reg[15][11]  ( .D(n2056), .CP(clk), .Q(\buff_mem[15][11] )
         );
  dff_sg \buff_mem_reg[15][10]  ( .D(n2057), .CP(clk), .Q(\buff_mem[15][10] )
         );
  dff_sg \buff_mem_reg[15][9]  ( .D(n2058), .CP(clk), .Q(\buff_mem[15][9] ) );
  dff_sg \buff_mem_reg[15][8]  ( .D(n2059), .CP(clk), .Q(\buff_mem[15][8] ) );
  dff_sg \buff_mem_reg[15][7]  ( .D(n2060), .CP(clk), .Q(\buff_mem[15][7] ) );
  dff_sg \buff_mem_reg[15][6]  ( .D(n2061), .CP(clk), .Q(\buff_mem[15][6] ) );
  dff_sg \buff_mem_reg[15][5]  ( .D(n2062), .CP(clk), .Q(\buff_mem[15][5] ) );
  dff_sg \buff_mem_reg[15][4]  ( .D(n2063), .CP(clk), .Q(\buff_mem[15][4] ) );
  dff_sg \buff_mem_reg[15][3]  ( .D(n2064), .CP(clk), .Q(\buff_mem[15][3] ) );
  dff_sg \buff_mem_reg[15][2]  ( .D(n2065), .CP(clk), .Q(\buff_mem[15][2] ) );
  dff_sg \buff_mem_reg[15][1]  ( .D(n2066), .CP(clk), .Q(\buff_mem[15][1] ) );
  dff_sg \buff_mem_reg[15][0]  ( .D(n2067), .CP(clk), .Q(\buff_mem[15][0] ) );
  dff_sg \buff_mem_reg[14][19]  ( .D(n2068), .CP(clk), .Q(\buff_mem[14][19] )
         );
  dff_sg \buff_mem_reg[14][18]  ( .D(n2069), .CP(clk), .Q(\buff_mem[14][18] )
         );
  dff_sg \buff_mem_reg[14][17]  ( .D(n2070), .CP(clk), .Q(\buff_mem[14][17] )
         );
  dff_sg \buff_mem_reg[14][16]  ( .D(n2071), .CP(clk), .Q(\buff_mem[14][16] )
         );
  dff_sg \buff_mem_reg[14][15]  ( .D(n2072), .CP(clk), .Q(\buff_mem[14][15] )
         );
  dff_sg \buff_mem_reg[14][13]  ( .D(n2074), .CP(clk), .Q(\buff_mem[14][13] )
         );
  dff_sg \buff_mem_reg[14][12]  ( .D(n2075), .CP(clk), .Q(\buff_mem[14][12] )
         );
  dff_sg \buff_mem_reg[14][11]  ( .D(n2076), .CP(clk), .Q(\buff_mem[14][11] )
         );
  dff_sg \buff_mem_reg[14][10]  ( .D(n2077), .CP(clk), .Q(\buff_mem[14][10] )
         );
  dff_sg \buff_mem_reg[14][9]  ( .D(n2078), .CP(clk), .Q(\buff_mem[14][9] ) );
  dff_sg \buff_mem_reg[14][8]  ( .D(n2079), .CP(clk), .Q(\buff_mem[14][8] ) );
  dff_sg \buff_mem_reg[14][7]  ( .D(n2080), .CP(clk), .Q(\buff_mem[14][7] ) );
  dff_sg \buff_mem_reg[14][6]  ( .D(n2081), .CP(clk), .Q(\buff_mem[14][6] ) );
  dff_sg \buff_mem_reg[14][5]  ( .D(n2082), .CP(clk), .Q(\buff_mem[14][5] ) );
  dff_sg \buff_mem_reg[14][4]  ( .D(n2083), .CP(clk), .Q(\buff_mem[14][4] ) );
  dff_sg \buff_mem_reg[14][3]  ( .D(n2084), .CP(clk), .Q(\buff_mem[14][3] ) );
  dff_sg \buff_mem_reg[14][2]  ( .D(n2085), .CP(clk), .Q(\buff_mem[14][2] ) );
  dff_sg \buff_mem_reg[14][1]  ( .D(n2086), .CP(clk), .Q(\buff_mem[14][1] ) );
  dff_sg \buff_mem_reg[14][0]  ( .D(n2087), .CP(clk), .Q(\buff_mem[14][0] ) );
  dff_sg \buff_mem_reg[13][19]  ( .D(n2088), .CP(clk), .Q(\buff_mem[13][19] )
         );
  dff_sg \buff_mem_reg[13][18]  ( .D(n2089), .CP(clk), .Q(\buff_mem[13][18] )
         );
  dff_sg \buff_mem_reg[13][17]  ( .D(n2090), .CP(clk), .Q(\buff_mem[13][17] )
         );
  dff_sg \buff_mem_reg[13][16]  ( .D(n2091), .CP(clk), .Q(\buff_mem[13][16] )
         );
  dff_sg \buff_mem_reg[13][15]  ( .D(n2092), .CP(clk), .Q(\buff_mem[13][15] )
         );
  dff_sg \buff_mem_reg[13][13]  ( .D(n2094), .CP(clk), .Q(\buff_mem[13][13] )
         );
  dff_sg \buff_mem_reg[13][12]  ( .D(n2095), .CP(clk), .Q(\buff_mem[13][12] )
         );
  dff_sg \buff_mem_reg[13][11]  ( .D(n2096), .CP(clk), .Q(\buff_mem[13][11] )
         );
  dff_sg \buff_mem_reg[13][10]  ( .D(n2097), .CP(clk), .Q(\buff_mem[13][10] )
         );
  dff_sg \buff_mem_reg[13][9]  ( .D(n2098), .CP(clk), .Q(\buff_mem[13][9] ) );
  dff_sg \buff_mem_reg[13][8]  ( .D(n2099), .CP(clk), .Q(\buff_mem[13][8] ) );
  dff_sg \buff_mem_reg[13][7]  ( .D(n2100), .CP(clk), .Q(\buff_mem[13][7] ) );
  dff_sg \buff_mem_reg[13][6]  ( .D(n2101), .CP(clk), .Q(\buff_mem[13][6] ) );
  dff_sg \buff_mem_reg[13][5]  ( .D(n2102), .CP(clk), .Q(\buff_mem[13][5] ) );
  dff_sg \buff_mem_reg[13][4]  ( .D(n2103), .CP(clk), .Q(\buff_mem[13][4] ) );
  dff_sg \buff_mem_reg[13][3]  ( .D(n2104), .CP(clk), .Q(\buff_mem[13][3] ) );
  dff_sg \buff_mem_reg[13][2]  ( .D(n2105), .CP(clk), .Q(\buff_mem[13][2] ) );
  dff_sg \buff_mem_reg[13][1]  ( .D(n2106), .CP(clk), .Q(\buff_mem[13][1] ) );
  dff_sg \buff_mem_reg[13][0]  ( .D(n2107), .CP(clk), .Q(\buff_mem[13][0] ) );
  dff_sg \buff_mem_reg[12][19]  ( .D(n2108), .CP(clk), .Q(\buff_mem[12][19] )
         );
  dff_sg \buff_mem_reg[12][18]  ( .D(n2109), .CP(clk), .Q(\buff_mem[12][18] )
         );
  dff_sg \buff_mem_reg[12][17]  ( .D(n2110), .CP(clk), .Q(\buff_mem[12][17] )
         );
  dff_sg \buff_mem_reg[12][16]  ( .D(n2111), .CP(clk), .Q(\buff_mem[12][16] )
         );
  dff_sg \buff_mem_reg[12][15]  ( .D(n2112), .CP(clk), .Q(\buff_mem[12][15] )
         );
  dff_sg \buff_mem_reg[12][13]  ( .D(n2114), .CP(clk), .Q(\buff_mem[12][13] )
         );
  dff_sg \buff_mem_reg[12][12]  ( .D(n2115), .CP(clk), .Q(\buff_mem[12][12] )
         );
  dff_sg \buff_mem_reg[12][11]  ( .D(n2116), .CP(clk), .Q(\buff_mem[12][11] )
         );
  dff_sg \buff_mem_reg[12][10]  ( .D(n2117), .CP(clk), .Q(\buff_mem[12][10] )
         );
  dff_sg \buff_mem_reg[12][9]  ( .D(n2118), .CP(clk), .Q(\buff_mem[12][9] ) );
  dff_sg \buff_mem_reg[12][8]  ( .D(n2119), .CP(clk), .Q(\buff_mem[12][8] ) );
  dff_sg \buff_mem_reg[12][7]  ( .D(n2120), .CP(clk), .Q(\buff_mem[12][7] ) );
  dff_sg \buff_mem_reg[12][6]  ( .D(n2121), .CP(clk), .Q(\buff_mem[12][6] ) );
  dff_sg \buff_mem_reg[12][5]  ( .D(n2122), .CP(clk), .Q(\buff_mem[12][5] ) );
  dff_sg \buff_mem_reg[12][4]  ( .D(n2123), .CP(clk), .Q(\buff_mem[12][4] ) );
  dff_sg \buff_mem_reg[12][3]  ( .D(n2124), .CP(clk), .Q(\buff_mem[12][3] ) );
  dff_sg \buff_mem_reg[12][2]  ( .D(n2125), .CP(clk), .Q(\buff_mem[12][2] ) );
  dff_sg \buff_mem_reg[12][1]  ( .D(n2126), .CP(clk), .Q(\buff_mem[12][1] ) );
  dff_sg \buff_mem_reg[12][0]  ( .D(n2127), .CP(clk), .Q(\buff_mem[12][0] ) );
  dff_sg \buff_mem_reg[7][19]  ( .D(n2208), .CP(clk), .Q(\buff_mem[7][19] ) );
  dff_sg \buff_mem_reg[7][18]  ( .D(n2209), .CP(clk), .Q(\buff_mem[7][18] ) );
  dff_sg \buff_mem_reg[7][17]  ( .D(n2210), .CP(clk), .Q(\buff_mem[7][17] ) );
  dff_sg \buff_mem_reg[7][16]  ( .D(n2211), .CP(clk), .Q(\buff_mem[7][16] ) );
  dff_sg \buff_mem_reg[7][15]  ( .D(n2212), .CP(clk), .Q(\buff_mem[7][15] ) );
  dff_sg \buff_mem_reg[7][13]  ( .D(n2214), .CP(clk), .Q(\buff_mem[7][13] ) );
  dff_sg \buff_mem_reg[7][12]  ( .D(n2215), .CP(clk), .Q(\buff_mem[7][12] ) );
  dff_sg \buff_mem_reg[7][11]  ( .D(n2216), .CP(clk), .Q(\buff_mem[7][11] ) );
  dff_sg \buff_mem_reg[7][10]  ( .D(n2217), .CP(clk), .Q(\buff_mem[7][10] ) );
  dff_sg \buff_mem_reg[7][9]  ( .D(n2218), .CP(clk), .Q(\buff_mem[7][9] ) );
  dff_sg \buff_mem_reg[7][8]  ( .D(n2219), .CP(clk), .Q(\buff_mem[7][8] ) );
  dff_sg \buff_mem_reg[7][7]  ( .D(n2220), .CP(clk), .Q(\buff_mem[7][7] ) );
  dff_sg \buff_mem_reg[7][6]  ( .D(n2221), .CP(clk), .Q(\buff_mem[7][6] ) );
  dff_sg \buff_mem_reg[7][5]  ( .D(n2222), .CP(clk), .Q(\buff_mem[7][5] ) );
  dff_sg \buff_mem_reg[7][4]  ( .D(n2223), .CP(clk), .Q(\buff_mem[7][4] ) );
  dff_sg \buff_mem_reg[7][3]  ( .D(n2224), .CP(clk), .Q(\buff_mem[7][3] ) );
  dff_sg \buff_mem_reg[7][2]  ( .D(n2225), .CP(clk), .Q(\buff_mem[7][2] ) );
  dff_sg \buff_mem_reg[7][1]  ( .D(n2226), .CP(clk), .Q(\buff_mem[7][1] ) );
  dff_sg \buff_mem_reg[7][0]  ( .D(n2227), .CP(clk), .Q(\buff_mem[7][0] ) );
  dff_sg \buff_mem_reg[6][19]  ( .D(n2228), .CP(clk), .Q(\buff_mem[6][19] ) );
  dff_sg \buff_mem_reg[6][18]  ( .D(n2229), .CP(clk), .Q(\buff_mem[6][18] ) );
  dff_sg \buff_mem_reg[6][17]  ( .D(n2230), .CP(clk), .Q(\buff_mem[6][17] ) );
  dff_sg \buff_mem_reg[6][16]  ( .D(n2231), .CP(clk), .Q(\buff_mem[6][16] ) );
  dff_sg \buff_mem_reg[6][15]  ( .D(n2232), .CP(clk), .Q(\buff_mem[6][15] ) );
  dff_sg \buff_mem_reg[6][13]  ( .D(n2234), .CP(clk), .Q(\buff_mem[6][13] ) );
  dff_sg \buff_mem_reg[6][12]  ( .D(n2235), .CP(clk), .Q(\buff_mem[6][12] ) );
  dff_sg \buff_mem_reg[6][11]  ( .D(n2236), .CP(clk), .Q(\buff_mem[6][11] ) );
  dff_sg \buff_mem_reg[6][10]  ( .D(n2237), .CP(clk), .Q(\buff_mem[6][10] ) );
  dff_sg \buff_mem_reg[6][9]  ( .D(n2238), .CP(clk), .Q(\buff_mem[6][9] ) );
  dff_sg \buff_mem_reg[6][8]  ( .D(n2239), .CP(clk), .Q(\buff_mem[6][8] ) );
  dff_sg \buff_mem_reg[6][7]  ( .D(n2240), .CP(clk), .Q(\buff_mem[6][7] ) );
  dff_sg \buff_mem_reg[6][6]  ( .D(n2241), .CP(clk), .Q(\buff_mem[6][6] ) );
  dff_sg \buff_mem_reg[6][5]  ( .D(n2242), .CP(clk), .Q(\buff_mem[6][5] ) );
  dff_sg \buff_mem_reg[6][4]  ( .D(n2243), .CP(clk), .Q(\buff_mem[6][4] ) );
  dff_sg \buff_mem_reg[6][3]  ( .D(n2244), .CP(clk), .Q(\buff_mem[6][3] ) );
  dff_sg \buff_mem_reg[6][2]  ( .D(n2245), .CP(clk), .Q(\buff_mem[6][2] ) );
  dff_sg \buff_mem_reg[6][1]  ( .D(n2246), .CP(clk), .Q(\buff_mem[6][1] ) );
  dff_sg \buff_mem_reg[6][0]  ( .D(n2247), .CP(clk), .Q(\buff_mem[6][0] ) );
  dff_sg \buff_mem_reg[5][19]  ( .D(n2248), .CP(clk), .Q(\buff_mem[5][19] ) );
  dff_sg \buff_mem_reg[5][18]  ( .D(n2249), .CP(clk), .Q(\buff_mem[5][18] ) );
  dff_sg \buff_mem_reg[5][17]  ( .D(n2250), .CP(clk), .Q(\buff_mem[5][17] ) );
  dff_sg \buff_mem_reg[5][16]  ( .D(n2251), .CP(clk), .Q(\buff_mem[5][16] ) );
  dff_sg \buff_mem_reg[5][15]  ( .D(n2252), .CP(clk), .Q(\buff_mem[5][15] ) );
  dff_sg \buff_mem_reg[5][13]  ( .D(n2254), .CP(clk), .Q(\buff_mem[5][13] ) );
  dff_sg \buff_mem_reg[5][12]  ( .D(n2255), .CP(clk), .Q(\buff_mem[5][12] ) );
  dff_sg \buff_mem_reg[5][11]  ( .D(n2256), .CP(clk), .Q(\buff_mem[5][11] ) );
  dff_sg \buff_mem_reg[5][10]  ( .D(n2257), .CP(clk), .Q(\buff_mem[5][10] ) );
  dff_sg \buff_mem_reg[5][9]  ( .D(n2258), .CP(clk), .Q(\buff_mem[5][9] ) );
  dff_sg \buff_mem_reg[5][8]  ( .D(n2259), .CP(clk), .Q(\buff_mem[5][8] ) );
  dff_sg \buff_mem_reg[5][7]  ( .D(n2260), .CP(clk), .Q(\buff_mem[5][7] ) );
  dff_sg \buff_mem_reg[5][6]  ( .D(n2261), .CP(clk), .Q(\buff_mem[5][6] ) );
  dff_sg \buff_mem_reg[5][5]  ( .D(n2262), .CP(clk), .Q(\buff_mem[5][5] ) );
  dff_sg \buff_mem_reg[5][4]  ( .D(n2263), .CP(clk), .Q(\buff_mem[5][4] ) );
  dff_sg \buff_mem_reg[5][3]  ( .D(n2264), .CP(clk), .Q(\buff_mem[5][3] ) );
  dff_sg \buff_mem_reg[5][2]  ( .D(n2265), .CP(clk), .Q(\buff_mem[5][2] ) );
  dff_sg \buff_mem_reg[5][1]  ( .D(n2266), .CP(clk), .Q(\buff_mem[5][1] ) );
  dff_sg \buff_mem_reg[5][0]  ( .D(n2267), .CP(clk), .Q(\buff_mem[5][0] ) );
  dff_sg \buff_mem_reg[4][13]  ( .D(n2274), .CP(clk), .Q(\buff_mem[4][13] ) );
  dff_sg \buff_mem_reg[4][12]  ( .D(n2275), .CP(clk), .Q(\buff_mem[4][12] ) );
  dff_sg \buff_mem_reg[4][11]  ( .D(n2276), .CP(clk), .Q(\buff_mem[4][11] ) );
  dff_sg \buff_mem_reg[4][10]  ( .D(n2277), .CP(clk), .Q(\buff_mem[4][10] ) );
  dff_sg \buff_mem_reg[4][9]  ( .D(n2278), .CP(clk), .Q(\buff_mem[4][9] ) );
  dff_sg \buff_mem_reg[4][8]  ( .D(n2279), .CP(clk), .Q(\buff_mem[4][8] ) );
  dff_sg \buff_mem_reg[4][7]  ( .D(n2280), .CP(clk), .Q(\buff_mem[4][7] ) );
  dff_sg \buff_mem_reg[4][6]  ( .D(n2281), .CP(clk), .Q(\buff_mem[4][6] ) );
  dff_sg \buff_mem_reg[4][5]  ( .D(n2282), .CP(clk), .Q(\buff_mem[4][5] ) );
  dff_sg \buff_mem_reg[4][4]  ( .D(n2283), .CP(clk), .Q(\buff_mem[4][4] ) );
  dff_sg \buff_mem_reg[4][3]  ( .D(n2284), .CP(clk), .Q(\buff_mem[4][3] ) );
  dff_sg \buff_mem_reg[4][2]  ( .D(n2285), .CP(clk), .Q(\buff_mem[4][2] ) );
  dff_sg \buff_mem_reg[4][1]  ( .D(n2286), .CP(clk), .Q(\buff_mem[4][1] ) );
  dff_sg \buff_mem_reg[4][0]  ( .D(n2287), .CP(clk), .Q(\buff_mem[4][0] ) );
  dff_sg \buff_mem_reg[4][19]  ( .D(n2268), .CP(clk), .Q(\buff_mem[4][19] ) );
  dff_sg \buff_mem_reg[4][18]  ( .D(n2269), .CP(clk), .Q(\buff_mem[4][18] ) );
  dff_sg \buff_mem_reg[4][17]  ( .D(n2270), .CP(clk), .Q(\buff_mem[4][17] ) );
  dff_sg \buff_mem_reg[4][16]  ( .D(n2271), .CP(clk), .Q(\buff_mem[4][16] ) );
  dff_sg \buff_mem_reg[4][15]  ( .D(n2272), .CP(clk), .Q(\buff_mem[4][15] ) );
  dff_sg \buff_mem_reg[3][14]  ( .D(n2293), .CP(clk), .Q(\buff_mem[3][14] ) );
  dff_sg \buff_mem_reg[2][14]  ( .D(n2313), .CP(clk), .Q(\buff_mem[2][14] ) );
  dff_sg \buff_mem_reg[1][14]  ( .D(n2333), .CP(clk), .Q(\buff_mem[1][14] ) );
  dff_sg \buff_mem_reg[0][14]  ( .D(n2353), .CP(clk), .Q(\buff_mem[0][14] ) );
  dff_sg \buff_mem_reg[19][14]  ( .D(n1973), .CP(clk), .Q(\buff_mem[19][14] )
         );
  dff_sg \buff_mem_reg[18][14]  ( .D(n1993), .CP(clk), .Q(\buff_mem[18][14] )
         );
  dff_sg \buff_mem_reg[17][14]  ( .D(n2013), .CP(clk), .Q(\buff_mem[17][14] )
         );
  dff_sg \buff_mem_reg[16][14]  ( .D(n2033), .CP(clk), .Q(\buff_mem[16][14] )
         );
  dff_sg \buff_mem_reg[15][14]  ( .D(n2053), .CP(clk), .Q(\buff_mem[15][14] )
         );
  dff_sg \buff_mem_reg[14][14]  ( .D(n2073), .CP(clk), .Q(\buff_mem[14][14] )
         );
  dff_sg \buff_mem_reg[13][14]  ( .D(n2093), .CP(clk), .Q(\buff_mem[13][14] )
         );
  dff_sg \buff_mem_reg[12][14]  ( .D(n2113), .CP(clk), .Q(\buff_mem[12][14] )
         );
  dff_sg \buff_mem_reg[11][14]  ( .D(n2133), .CP(clk), .Q(\buff_mem[11][14] )
         );
  dff_sg \buff_mem_reg[10][14]  ( .D(n2153), .CP(clk), .Q(\buff_mem[10][14] )
         );
  dff_sg \buff_mem_reg[9][14]  ( .D(n2173), .CP(clk), .Q(\buff_mem[9][14] ) );
  dff_sg \buff_mem_reg[8][14]  ( .D(n2193), .CP(clk), .Q(\buff_mem[8][14] ) );
  dff_sg \buff_mem_reg[7][14]  ( .D(n2213), .CP(clk), .Q(\buff_mem[7][14] ) );
  dff_sg \buff_mem_reg[6][14]  ( .D(n2233), .CP(clk), .Q(\buff_mem[6][14] ) );
  dff_sg \buff_mem_reg[5][14]  ( .D(n2253), .CP(clk), .Q(\buff_mem[5][14] ) );
  dff_sg \buff_mem_reg[4][14]  ( .D(n2273), .CP(clk), .Q(\buff_mem[4][14] ) );
  dff_sg \data_out_reg[19]  ( .D(N161), .CP(clk), .Q(data_out[19]) );
  dff_sg \data_out_reg[18]  ( .D(N160), .CP(clk), .Q(data_out[18]) );
  dff_sg \data_out_reg[17]  ( .D(N159), .CP(clk), .Q(data_out[17]) );
  dff_sg \data_out_reg[16]  ( .D(N158), .CP(clk), .Q(data_out[16]) );
  dff_sg \data_out_reg[15]  ( .D(N157), .CP(clk), .Q(data_out[15]) );
  dff_sg \data_out_reg[14]  ( .D(N156), .CP(clk), .Q(data_out[14]) );
  dff_sg \data_out_reg[13]  ( .D(N155), .CP(clk), .Q(data_out[13]) );
  dff_sg \data_out_reg[12]  ( .D(N154), .CP(clk), .Q(data_out[12]) );
  dff_sg \data_out_reg[11]  ( .D(N153), .CP(clk), .Q(data_out[11]) );
  dff_sg \data_out_reg[10]  ( .D(N152), .CP(clk), .Q(data_out[10]) );
  dff_sg \data_out_reg[9]  ( .D(N151), .CP(clk), .Q(data_out[9]) );
  dff_sg \data_out_reg[8]  ( .D(N150), .CP(clk), .Q(data_out[8]) );
  dff_sg \data_out_reg[7]  ( .D(N149), .CP(clk), .Q(data_out[7]) );
  dff_sg \data_out_reg[6]  ( .D(N148), .CP(clk), .Q(data_out[6]) );
  dff_sg \data_out_reg[5]  ( .D(N147), .CP(clk), .Q(data_out[5]) );
  dff_sg \data_out_reg[4]  ( .D(N146), .CP(clk), .Q(data_out[4]) );
  dff_sg \data_out_reg[3]  ( .D(N145), .CP(clk), .Q(data_out[3]) );
  dff_sg \data_out_reg[2]  ( .D(N144), .CP(clk), .Q(data_out[2]) );
  dff_sg \data_out_reg[1]  ( .D(N143), .CP(clk), .Q(data_out[1]) );
  dff_sg \data_out_reg[0]  ( .D(N142), .CP(clk), .Q(data_out[0]) );
  nor_x1_sg U4799 ( .A(n5169), .B(n5170), .X(n5167) );
  nor_x1_sg U4800 ( .A(n5129), .B(n5130), .X(n5128) );
  nor_x1_sg U4801 ( .A(n5090), .B(n5091), .X(n5089) );
  nor_x1_sg U4802 ( .A(n5051), .B(n5052), .X(n5050) );
  nor_x1_sg U4803 ( .A(n5012), .B(n5013), .X(n5011) );
  nor_x1_sg U4804 ( .A(n4973), .B(n4974), .X(n4972) );
  nor_x1_sg U4805 ( .A(n4934), .B(n4935), .X(n4933) );
  nor_x1_sg U4806 ( .A(n4895), .B(n4896), .X(n4894) );
  nor_x1_sg U4807 ( .A(n4856), .B(n4857), .X(n4855) );
  nor_x1_sg U4808 ( .A(n4817), .B(n4818), .X(n4816) );
  nor_x1_sg U4809 ( .A(n4778), .B(n4779), .X(n4777) );
  nor_x1_sg U4810 ( .A(n4739), .B(n4740), .X(n4738) );
  nor_x1_sg U4811 ( .A(n4700), .B(n4701), .X(n4699) );
  nor_x1_sg U4812 ( .A(n4661), .B(n4662), .X(n4660) );
  nor_x1_sg U4813 ( .A(n4622), .B(n4623), .X(n4621) );
  nor_x1_sg U4814 ( .A(n4583), .B(n4584), .X(n4582) );
  nor_x1_sg U4815 ( .A(n4544), .B(n4545), .X(n4543) );
  nor_x1_sg U4816 ( .A(n4505), .B(n4506), .X(n4504) );
  nor_x1_sg U4817 ( .A(n4466), .B(n4467), .X(n4465) );
  nor_x1_sg U4818 ( .A(n4409), .B(n4410), .X(n4408) );
  inv_x8_sg U4819 ( .A(data_in[14]), .X(n5892) );
  inv_x1_sg U4820 ( .A(n5727), .X(n5728) );
  inv_x1_sg U4821 ( .A(n5951), .X(n5660) );
  inv_x1_sg U4822 ( .A(n5655), .X(n5657) );
  inv_x8_sg U4823 ( .A(data_in[16]), .X(n3269) );
  inv_x8_sg U4824 ( .A(data_in[19]), .X(n3266) );
  inv_x8_sg U4825 ( .A(data_in[0]), .X(n5919) );
  inv_x8_sg U4826 ( .A(data_in[1]), .X(n5908) );
  inv_x8_sg U4827 ( .A(data_in[2]), .X(n5894) );
  inv_x8_sg U4828 ( .A(data_in[3]), .X(n3282) );
  inv_x8_sg U4829 ( .A(data_in[4]), .X(n5890) );
  inv_x8_sg U4830 ( .A(data_in[5]), .X(n5910) );
  inv_x8_sg U4831 ( .A(data_in[8]), .X(n3277) );
  inv_x1_sg U4832 ( .A(n5216), .X(n5354) );
  inv_x8_sg U4833 ( .A(data_in[9]), .X(n3276) );
  inv_x1_sg U4834 ( .A(n5355), .X(n5350) );
  inv_x8_sg U4835 ( .A(data_in[10]), .X(n3275) );
  inv_x8_sg U4836 ( .A(data_in[11]), .X(n5909) );
  inv_x8_sg U4837 ( .A(data_in[12]), .X(n3273) );
  inv_x1_sg U4838 ( .A(n3920), .X(n5347) );
  inv_x1_sg U4839 ( .A(n5780), .X(n5781) );
  inv_x8_sg U4840 ( .A(data_in[13]), .X(n3272) );
  inv_x1_sg U4841 ( .A(n5668), .X(n5669) );
  nand_x1_sg U4842 ( .A(n5844), .B(n5190), .X(n5186) );
  nand_x1_sg U4843 ( .A(n5864), .B(n5201), .X(n5197) );
  nand_x1_sg U4844 ( .A(n5865), .B(n5155), .X(n5151) );
  nand_x1_sg U4845 ( .A(n5845), .B(n5145), .X(n5141) );
  nand_x1_sg U4846 ( .A(n5866), .B(n5116), .X(n5112) );
  nand_x1_sg U4847 ( .A(n5846), .B(n5106), .X(n5102) );
  nand_x1_sg U4848 ( .A(n5847), .B(n5067), .X(n5063) );
  nand_x1_sg U4849 ( .A(n5867), .B(n5077), .X(n5073) );
  nand_x1_sg U4850 ( .A(n5868), .B(n5038), .X(n5034) );
  nand_x1_sg U4851 ( .A(n5848), .B(n5028), .X(n5024) );
  nand_x1_sg U4852 ( .A(n5869), .B(n4999), .X(n4995) );
  nand_x1_sg U4853 ( .A(n5849), .B(n4989), .X(n4985) );
  nand_x1_sg U4854 ( .A(n5870), .B(n4960), .X(n4956) );
  nand_x1_sg U4855 ( .A(n5850), .B(n4950), .X(n4946) );
  nand_x1_sg U4856 ( .A(n5871), .B(n4921), .X(n4917) );
  nand_x1_sg U4857 ( .A(n5851), .B(n4911), .X(n4907) );
  nand_x1_sg U4858 ( .A(n5872), .B(n4882), .X(n4878) );
  nand_x1_sg U4859 ( .A(n5852), .B(n4872), .X(n4868) );
  nand_x1_sg U4860 ( .A(n5853), .B(n4833), .X(n4829) );
  nand_x1_sg U4861 ( .A(n5873), .B(n4843), .X(n4839) );
  nand_x1_sg U4862 ( .A(n5874), .B(n4804), .X(n4800) );
  nand_x1_sg U4863 ( .A(n5854), .B(n4794), .X(n4790) );
  nand_x1_sg U4864 ( .A(n5875), .B(n4765), .X(n4761) );
  nand_x1_sg U4865 ( .A(n5855), .B(n4755), .X(n4751) );
  nand_x1_sg U4866 ( .A(n5876), .B(n4726), .X(n4722) );
  nand_x1_sg U4867 ( .A(n5856), .B(n4716), .X(n4712) );
  nand_x1_sg U4868 ( .A(n5857), .B(n4677), .X(n4673) );
  nand_x1_sg U4869 ( .A(n5877), .B(n4687), .X(n4683) );
  nand_x1_sg U4870 ( .A(n5858), .B(n4638), .X(n4634) );
  nand_x1_sg U4871 ( .A(n5878), .B(n4648), .X(n4644) );
  nand_x1_sg U4872 ( .A(n5879), .B(n4609), .X(n4605) );
  nand_x1_sg U4873 ( .A(n5859), .B(n4599), .X(n4595) );
  nand_x1_sg U4874 ( .A(n5860), .B(n4560), .X(n4556) );
  nand_x1_sg U4875 ( .A(n5880), .B(n4570), .X(n4566) );
  nand_x1_sg U4876 ( .A(n5881), .B(n4531), .X(n4527) );
  nand_x1_sg U4877 ( .A(n5861), .B(n4521), .X(n4517) );
  nand_x1_sg U4878 ( .A(n5862), .B(n4482), .X(n4478) );
  nand_x1_sg U4879 ( .A(n5882), .B(n4492), .X(n4488) );
  nand_x1_sg U4880 ( .A(n5883), .B(n4446), .X(n4440) );
  nand_x1_sg U4881 ( .A(n5863), .B(n4432), .X(n4426) );
  nand_x1_sg U4882 ( .A(n4404), .B(n4405), .X(n3512) );
  inv_x1_sg U4883 ( .A(n3497), .X(n3290) );
  nand_x1_sg U4884 ( .A(n4394), .B(n4395), .X(n3509) );
  inv_x1_sg U4885 ( .A(n3462), .X(n3358) );
  nand_x1_sg U4886 ( .A(n3477), .B(n3478), .X(n3456) );
  nand_x2_sg U4887 ( .A(n5195), .B(n5196), .X(n5169) );
  nand_x2_sg U4888 ( .A(n5171), .B(n5172), .X(n5170) );
  nand_x2_sg U4889 ( .A(n5131), .B(n5132), .X(n5130) );
  nand_x2_sg U4890 ( .A(n5149), .B(n5150), .X(n5129) );
  nand_x2_sg U4891 ( .A(n5092), .B(n5093), .X(n5091) );
  nand_x2_sg U4892 ( .A(n5110), .B(n5111), .X(n5090) );
  nand_x2_sg U4893 ( .A(n5071), .B(n5072), .X(n5051) );
  nand_x2_sg U4894 ( .A(n5053), .B(n5054), .X(n5052) );
  nand_x2_sg U4895 ( .A(n5014), .B(n5015), .X(n5013) );
  nand_x2_sg U4896 ( .A(n5032), .B(n5033), .X(n5012) );
  nand_x2_sg U4897 ( .A(n4975), .B(n4976), .X(n4974) );
  nand_x2_sg U4898 ( .A(n4993), .B(n4994), .X(n4973) );
  nand_x2_sg U4899 ( .A(n4936), .B(n4937), .X(n4935) );
  nand_x2_sg U4900 ( .A(n4954), .B(n4955), .X(n4934) );
  nand_x2_sg U4901 ( .A(n4897), .B(n4898), .X(n4896) );
  nand_x2_sg U4902 ( .A(n4915), .B(n4916), .X(n4895) );
  nand_x2_sg U4903 ( .A(n4858), .B(n4859), .X(n4857) );
  nand_x2_sg U4904 ( .A(n4876), .B(n4877), .X(n4856) );
  nand_x2_sg U4905 ( .A(n4837), .B(n4838), .X(n4817) );
  nand_x2_sg U4906 ( .A(n4819), .B(n4820), .X(n4818) );
  nand_x2_sg U4907 ( .A(n4780), .B(n4781), .X(n4779) );
  nand_x2_sg U4908 ( .A(n4798), .B(n4799), .X(n4778) );
  nand_x2_sg U4909 ( .A(n4741), .B(n4742), .X(n4740) );
  nand_x2_sg U4910 ( .A(n4759), .B(n4760), .X(n4739) );
  nand_x2_sg U4911 ( .A(n4702), .B(n4703), .X(n4701) );
  nand_x2_sg U4912 ( .A(n4720), .B(n4721), .X(n4700) );
  nand_x2_sg U4913 ( .A(n4681), .B(n4682), .X(n4661) );
  nand_x2_sg U4914 ( .A(n4663), .B(n4664), .X(n4662) );
  nand_x2_sg U4915 ( .A(n4642), .B(n4643), .X(n4622) );
  nand_x2_sg U4916 ( .A(n4624), .B(n4625), .X(n4623) );
  nand_x2_sg U4917 ( .A(n4585), .B(n4586), .X(n4584) );
  nand_x2_sg U4918 ( .A(n4603), .B(n4604), .X(n4583) );
  nand_x2_sg U4919 ( .A(n4564), .B(n4565), .X(n4544) );
  nand_x2_sg U4920 ( .A(n4546), .B(n4547), .X(n4545) );
  nand_x2_sg U4921 ( .A(n4507), .B(n4508), .X(n4506) );
  nand_x2_sg U4922 ( .A(n4525), .B(n4526), .X(n4505) );
  nand_x2_sg U4923 ( .A(n4486), .B(n4487), .X(n4466) );
  nand_x2_sg U4924 ( .A(n4468), .B(n4469), .X(n4467) );
  nand_x2_sg U4925 ( .A(n4411), .B(n4412), .X(n4410) );
  nand_x2_sg U4926 ( .A(n4438), .B(n4439), .X(n4409) );
  inv_x16_sg U4927 ( .A(reset), .X(n5214) );
  inv_x16_sg U4928 ( .A(reset), .X(n5215) );
  inv_x16_sg U4929 ( .A(reset), .X(n5825) );
  nand_x16_sg U4930 ( .A(n5825), .B(n3618), .X(n5803) );
  nand_x16_sg U4931 ( .A(n5215), .B(n4129), .X(n5951) );
  nand_x4_sg U4932 ( .A(n5899), .B(n4001), .X(n5780) );
  nand_x4_sg U4933 ( .A(n5927), .B(n3831), .X(n5727) );
  nand_x4_sg U4934 ( .A(n5901), .B(n3702), .X(n5668) );
  nand_x4_sg U4935 ( .A(n5896), .B(n3959), .X(n5216) );
  nand_x1_sg U4936 ( .A(n3260), .B(n5323), .X(n3959) );
  inv_x1_sg U4937 ( .A(n5177), .X(n5217) );
  inv_x1_sg U4938 ( .A(n5217), .X(n5218) );
  inv_x1_sg U4939 ( .A(n3576), .X(n5219) );
  inv_x1_sg U4940 ( .A(n5219), .X(n5220) );
  inv_x1_sg U4941 ( .A(wr_ptr[4]), .X(n5221) );
  inv_x1_sg U4942 ( .A(n5221), .X(n5222) );
  inv_x1_sg U4943 ( .A(rd_ptr[0]), .X(n5223) );
  inv_x1_sg U4944 ( .A(n5223), .X(n5224) );
  inv_x1_sg U4945 ( .A(n5947), .X(n5225) );
  inv_x1_sg U4946 ( .A(n5357), .X(n5226) );
  inv_x1_sg U4947 ( .A(n5945), .X(n5227) );
  inv_x1_sg U4948 ( .A(n5362), .X(n5228) );
  inv_x1_sg U4949 ( .A(n5944), .X(n5229) );
  inv_x1_sg U4950 ( .A(n5367), .X(n5230) );
  inv_x1_sg U4951 ( .A(n3541), .X(n5231) );
  inv_x1_sg U4952 ( .A(n5372), .X(n5232) );
  inv_x1_sg U4953 ( .A(n3574), .X(n5233) );
  inv_x1_sg U4954 ( .A(n5233), .X(n5234) );
  inv_x1_sg U4955 ( .A(n5937), .X(n5235) );
  inv_x1_sg U4956 ( .A(n5235), .X(n5236) );
  inv_x1_sg U4957 ( .A(n4445), .X(n5237) );
  inv_x1_sg U4958 ( .A(n5237), .X(n5238) );
  inv_x1_sg U4959 ( .A(n5903), .X(n5239) );
  inv_x1_sg U4960 ( .A(n5392), .X(n5240) );
  inv_x1_sg U4961 ( .A(n5902), .X(n5241) );
  inv_x1_sg U4962 ( .A(n5397), .X(n5242) );
  inv_x1_sg U4963 ( .A(n5904), .X(n5243) );
  inv_x1_sg U4964 ( .A(n5402), .X(n5244) );
  inv_x1_sg U4965 ( .A(n5905), .X(n5245) );
  inv_x1_sg U4966 ( .A(n5407), .X(n5246) );
  inv_x1_sg U4967 ( .A(n5922), .X(n5247) );
  inv_x1_sg U4968 ( .A(n5419), .X(n5248) );
  inv_x1_sg U4969 ( .A(n5923), .X(n5249) );
  inv_x1_sg U4970 ( .A(n5424), .X(n5250) );
  inv_x1_sg U4971 ( .A(n5924), .X(n5251) );
  inv_x1_sg U4972 ( .A(n5429), .X(n5252) );
  inv_x1_sg U4973 ( .A(n5925), .X(n5253) );
  inv_x1_sg U4974 ( .A(n5434), .X(n5254) );
  inv_x1_sg U4975 ( .A(n5926), .X(n5255) );
  inv_x1_sg U4976 ( .A(n5439), .X(n5256) );
  inv_x1_sg U4977 ( .A(n4418), .X(n5257) );
  inv_x1_sg U4978 ( .A(n5257), .X(n5258) );
  inv_x1_sg U4979 ( .A(n5940), .X(n5259) );
  inv_x1_sg U4980 ( .A(n5259), .X(n5260) );
  inv_x1_sg U4981 ( .A(n5939), .X(n5261) );
  inv_x1_sg U4982 ( .A(n5261), .X(n5262) );
  inv_x1_sg U4983 ( .A(n5936), .X(n5263) );
  inv_x1_sg U4984 ( .A(n5263), .X(n5264) );
  inv_x1_sg U4985 ( .A(n4437), .X(n5265) );
  inv_x1_sg U4986 ( .A(n5265), .X(n5266) );
  inv_x1_sg U4987 ( .A(n5933), .X(n5267) );
  inv_x1_sg U4988 ( .A(n5267), .X(n5268) );
  inv_x1_sg U4989 ( .A(n5932), .X(n5269) );
  inv_x1_sg U4990 ( .A(n5269), .X(n5270) );
  inv_x1_sg U4991 ( .A(n5935), .X(n5271) );
  inv_x1_sg U4992 ( .A(n5271), .X(n5272) );
  inv_x1_sg U4993 ( .A(n4460), .X(n5273) );
  inv_x1_sg U4994 ( .A(n5273), .X(n5274) );
  inv_x1_sg U4995 ( .A(n4433), .X(n5275) );
  inv_x1_sg U4996 ( .A(n5275), .X(n5276) );
  inv_x1_sg U4997 ( .A(n5934), .X(n5277) );
  inv_x1_sg U4998 ( .A(n5277), .X(n5278) );
  inv_x1_sg U4999 ( .A(n5931), .X(n5279) );
  inv_x1_sg U5000 ( .A(n5279), .X(n5280) );
  inv_x1_sg U5001 ( .A(n5948), .X(n5281) );
  inv_x1_sg U5002 ( .A(n5519), .X(n5282) );
  inv_x1_sg U5003 ( .A(n3520), .X(n5283) );
  inv_x1_sg U5004 ( .A(n5524), .X(n5284) );
  inv_x1_sg U5005 ( .A(n3526), .X(n5285) );
  inv_x1_sg U5006 ( .A(n5529), .X(n5286) );
  inv_x1_sg U5007 ( .A(n3550), .X(n5287) );
  inv_x1_sg U5008 ( .A(n5534), .X(n5288) );
  inv_x1_sg U5009 ( .A(n3920), .X(n5289) );
  inv_x1_sg U5010 ( .A(n5760), .X(n5290) );
  inv_x1_sg U5011 ( .A(n5727), .X(n5291) );
  inv_x1_sg U5012 ( .A(n5668), .X(n5292) );
  inv_x1_sg U5013 ( .A(n5740), .X(n5293) );
  inv_x1_sg U5014 ( .A(n5570), .X(n5294) );
  inv_x1_sg U5015 ( .A(n4260), .X(n5295) );
  inv_x1_sg U5016 ( .A(n5750), .X(n5296) );
  inv_x1_sg U5017 ( .A(n5949), .X(n5297) );
  inv_x1_sg U5018 ( .A(n5654), .X(n5298) );
  inv_x1_sg U5019 ( .A(n5770), .X(n5299) );
  inv_x1_sg U5020 ( .A(n5886), .X(n5300) );
  inv_x1_sg U5021 ( .A(n5681), .X(n5301) );
  inv_x1_sg U5022 ( .A(n5953), .X(n5302) );
  inv_x1_sg U5023 ( .A(n3621), .X(n5303) );
  inv_x1_sg U5024 ( .A(n5804), .X(n5304) );
  inv_x1_sg U5025 ( .A(n5885), .X(n5305) );
  inv_x1_sg U5026 ( .A(n5712), .X(n5306) );
  inv_x1_sg U5027 ( .A(n5793), .X(n5307) );
  inv_x1_sg U5028 ( .A(n5780), .X(n5308) );
  inv_x1_sg U5029 ( .A(n3547), .X(n5309) );
  inv_x1_sg U5030 ( .A(n5643), .X(n5310) );
  inv_x1_sg U5031 ( .A(n5946), .X(n5311) );
  inv_x1_sg U5032 ( .A(n5648), .X(n5312) );
  nand_x4_sg U5033 ( .A(n5214), .B(n4383), .X(n4344) );
  nand_x2_sg U5034 ( .A(n5900), .B(n4299), .X(n4260) );
  nand_x2_sg U5035 ( .A(n5929), .B(n4213), .X(n5949) );
  nand_x2_sg U5036 ( .A(n5900), .B(n3789), .X(n5886) );
  nand_x2_sg U5037 ( .A(n5901), .B(n3660), .X(n3621) );
  inv_x1_sg U5038 ( .A(n4396), .X(n5313) );
  inv_x1_sg U5039 ( .A(rd_ptr[1]), .X(n5314) );
  inv_x1_sg U5040 ( .A(n3371), .X(n5315) );
  inv_x1_sg U5041 ( .A(n5315), .X(n5316) );
  inv_x1_sg U5042 ( .A(n3465), .X(n5317) );
  inv_x1_sg U5043 ( .A(n5317), .X(n5318) );
  nor_x1_sg U5044 ( .A(reset), .B(empty), .X(n5319) );
  inv_x1_sg U5045 ( .A(n3468), .X(n5320) );
  inv_x1_sg U5046 ( .A(n5320), .X(n5321) );
  inv_x1_sg U5047 ( .A(n3469), .X(n5322) );
  inv_x1_sg U5048 ( .A(n5322), .X(n5323) );
  inv_x1_sg U5049 ( .A(wr_ptr[2]), .X(n5324) );
  inv_x1_sg U5050 ( .A(n5324), .X(n5325) );
  inv_x1_sg U5051 ( .A(n5833), .X(n5326) );
  inv_x1_sg U5052 ( .A(n5663), .X(n5327) );
  inv_x1_sg U5053 ( .A(n5676), .X(n5328) );
  inv_x1_sg U5054 ( .A(n5698), .X(n5329) );
  inv_x1_sg U5055 ( .A(n5722), .X(n5330) );
  inv_x1_sg U5056 ( .A(n5735), .X(n5331) );
  inv_x1_sg U5057 ( .A(n5788), .X(n5332) );
  inv_x1_sg U5058 ( .A(n4406), .X(n5333) );
  inv_x1_sg U5059 ( .A(n5812), .X(n5334) );
  inv_x1_sg U5060 ( .A(n5888), .X(n5335) );
  inv_x1_sg U5061 ( .A(n5335), .X(n5336) );
  inv_x1_sg U5062 ( .A(rd_ptr[4]), .X(n5337) );
  inv_x1_sg U5063 ( .A(n5337), .X(n5338) );
  inv_x1_sg U5064 ( .A(rd_ptr[2]), .X(n5339) );
  inv_x1_sg U5065 ( .A(n5339), .X(n5340) );
  inv_x1_sg U5066 ( .A(wr_ptr[3]), .X(n5341) );
  inv_x1_sg U5067 ( .A(n5341), .X(n5342) );
  inv_x1_sg U5068 ( .A(n5834), .X(n5343) );
  inv_x1_sg U5069 ( .A(rd_ptr[4]), .X(n5344) );
  inv_x1_sg U5070 ( .A(n3474), .X(n5345) );
  inv_x1_sg U5071 ( .A(n5820), .X(n5346) );
  inv_x1_sg U5072 ( .A(n5347), .X(n5348) );
  inv_x1_sg U5073 ( .A(n5347), .X(n5349) );
  inv_x1_sg U5074 ( .A(n5350), .X(n5351) );
  inv_x1_sg U5075 ( .A(n5350), .X(n5352) );
  inv_x1_sg U5076 ( .A(n5350), .X(n5353) );
  inv_x1_sg U5077 ( .A(n5354), .X(n5355) );
  inv_x1_sg U5078 ( .A(n5354), .X(n5356) );
  inv_x1_sg U5079 ( .A(n5947), .X(n5357) );
  inv_x1_sg U5080 ( .A(n5357), .X(n5358) );
  inv_x1_sg U5081 ( .A(n5357), .X(n5359) );
  inv_x1_sg U5082 ( .A(n5357), .X(n5360) );
  inv_x1_sg U5083 ( .A(n5225), .X(n5361) );
  inv_x1_sg U5084 ( .A(n5945), .X(n5362) );
  inv_x1_sg U5085 ( .A(n5362), .X(n5363) );
  inv_x1_sg U5086 ( .A(n5362), .X(n5364) );
  inv_x1_sg U5087 ( .A(n5362), .X(n5365) );
  inv_x1_sg U5088 ( .A(n5227), .X(n5366) );
  inv_x1_sg U5089 ( .A(n5944), .X(n5367) );
  inv_x1_sg U5090 ( .A(n5367), .X(n5368) );
  inv_x1_sg U5091 ( .A(n5367), .X(n5369) );
  inv_x1_sg U5092 ( .A(n5367), .X(n5370) );
  inv_x1_sg U5093 ( .A(n5229), .X(n5371) );
  inv_x1_sg U5094 ( .A(n3541), .X(n5372) );
  inv_x1_sg U5095 ( .A(n5372), .X(n5373) );
  inv_x1_sg U5096 ( .A(n5372), .X(n5374) );
  inv_x1_sg U5097 ( .A(n5372), .X(n5375) );
  inv_x1_sg U5098 ( .A(n5231), .X(n5376) );
  inv_x1_sg U5099 ( .A(n3574), .X(n5377) );
  inv_x1_sg U5100 ( .A(n5377), .X(n5378) );
  inv_x1_sg U5101 ( .A(n5377), .X(n5379) );
  inv_x1_sg U5102 ( .A(n5377), .X(n5380) );
  inv_x1_sg U5103 ( .A(n5377), .X(n5381) );
  inv_x1_sg U5104 ( .A(n5937), .X(n5382) );
  inv_x1_sg U5105 ( .A(n5382), .X(n5383) );
  inv_x1_sg U5106 ( .A(n5382), .X(n5384) );
  inv_x1_sg U5107 ( .A(n5382), .X(n5385) );
  inv_x1_sg U5108 ( .A(n5382), .X(n5386) );
  inv_x1_sg U5109 ( .A(n4445), .X(n5387) );
  inv_x1_sg U5110 ( .A(n5387), .X(n5388) );
  inv_x1_sg U5111 ( .A(n5387), .X(n5389) );
  inv_x1_sg U5112 ( .A(n5387), .X(n5390) );
  inv_x1_sg U5113 ( .A(n5387), .X(n5391) );
  inv_x1_sg U5114 ( .A(n5903), .X(n5392) );
  inv_x1_sg U5115 ( .A(n5392), .X(n5393) );
  inv_x1_sg U5116 ( .A(n5392), .X(n5394) );
  inv_x1_sg U5117 ( .A(n5392), .X(n5395) );
  inv_x1_sg U5118 ( .A(n5239), .X(n5396) );
  inv_x1_sg U5119 ( .A(n5902), .X(n5397) );
  inv_x1_sg U5120 ( .A(n5397), .X(n5398) );
  inv_x1_sg U5121 ( .A(n5397), .X(n5399) );
  inv_x1_sg U5122 ( .A(n5397), .X(n5400) );
  inv_x1_sg U5123 ( .A(n5241), .X(n5401) );
  inv_x1_sg U5124 ( .A(n5904), .X(n5402) );
  inv_x1_sg U5125 ( .A(n5402), .X(n5403) );
  inv_x1_sg U5126 ( .A(n5402), .X(n5404) );
  inv_x1_sg U5127 ( .A(n5402), .X(n5405) );
  inv_x1_sg U5128 ( .A(n5243), .X(n5406) );
  inv_x1_sg U5129 ( .A(n5905), .X(n5407) );
  inv_x1_sg U5130 ( .A(n5407), .X(n5408) );
  inv_x1_sg U5131 ( .A(n5407), .X(n5409) );
  inv_x1_sg U5132 ( .A(n5407), .X(n5410) );
  inv_x1_sg U5133 ( .A(n5245), .X(n5411) );
  inv_x1_sg U5134 ( .A(n5413), .X(n5412) );
  inv_x1_sg U5135 ( .A(n5914), .X(n5413) );
  inv_x1_sg U5136 ( .A(n5914), .X(n5414) );
  inv_x1_sg U5137 ( .A(n5413), .X(n5415) );
  inv_x1_sg U5138 ( .A(n5413), .X(n5416) );
  inv_x1_sg U5139 ( .A(n5414), .X(n5417) );
  inv_x1_sg U5140 ( .A(n5413), .X(n5418) );
  inv_x1_sg U5141 ( .A(n5922), .X(n5419) );
  inv_x1_sg U5142 ( .A(n5419), .X(n5420) );
  inv_x1_sg U5143 ( .A(n5419), .X(n5421) );
  inv_x1_sg U5144 ( .A(n5419), .X(n5422) );
  inv_x1_sg U5145 ( .A(n5247), .X(n5423) );
  inv_x1_sg U5146 ( .A(n5923), .X(n5424) );
  inv_x1_sg U5147 ( .A(n5424), .X(n5425) );
  inv_x1_sg U5148 ( .A(n5424), .X(n5426) );
  inv_x1_sg U5149 ( .A(n5424), .X(n5427) );
  inv_x1_sg U5150 ( .A(n5249), .X(n5428) );
  inv_x1_sg U5151 ( .A(n5924), .X(n5429) );
  inv_x1_sg U5152 ( .A(n5429), .X(n5430) );
  inv_x1_sg U5153 ( .A(n5429), .X(n5431) );
  inv_x1_sg U5154 ( .A(n5429), .X(n5432) );
  inv_x1_sg U5155 ( .A(n5251), .X(n5433) );
  inv_x1_sg U5156 ( .A(n5925), .X(n5434) );
  inv_x1_sg U5157 ( .A(n5434), .X(n5435) );
  inv_x1_sg U5158 ( .A(n5434), .X(n5436) );
  inv_x1_sg U5159 ( .A(n5434), .X(n5437) );
  inv_x1_sg U5160 ( .A(n5253), .X(n5438) );
  inv_x1_sg U5161 ( .A(n5926), .X(n5439) );
  inv_x1_sg U5162 ( .A(n5439), .X(n5440) );
  inv_x1_sg U5163 ( .A(n5439), .X(n5441) );
  inv_x1_sg U5164 ( .A(n5439), .X(n5442) );
  inv_x1_sg U5165 ( .A(n5255), .X(n5443) );
  inv_x1_sg U5166 ( .A(n4418), .X(n5444) );
  inv_x1_sg U5167 ( .A(n5444), .X(n5445) );
  inv_x1_sg U5168 ( .A(n5444), .X(n5446) );
  inv_x1_sg U5169 ( .A(n5444), .X(n5447) );
  inv_x1_sg U5170 ( .A(n5444), .X(n5448) );
  inv_x1_sg U5171 ( .A(n5940), .X(n5449) );
  inv_x1_sg U5172 ( .A(n5449), .X(n5450) );
  inv_x1_sg U5173 ( .A(n5449), .X(n5451) );
  inv_x1_sg U5174 ( .A(n5449), .X(n5452) );
  inv_x1_sg U5175 ( .A(n5449), .X(n5453) );
  inv_x1_sg U5176 ( .A(n5456), .X(n5454) );
  inv_x1_sg U5177 ( .A(n5938), .X(n5455) );
  inv_x1_sg U5178 ( .A(n5938), .X(n5456) );
  inv_x1_sg U5179 ( .A(n5455), .X(n5457) );
  inv_x1_sg U5180 ( .A(n5456), .X(n5458) );
  inv_x1_sg U5181 ( .A(n5456), .X(n5459) );
  inv_x1_sg U5182 ( .A(n5456), .X(n5460) );
  inv_x1_sg U5183 ( .A(n5939), .X(n5461) );
  inv_x1_sg U5184 ( .A(n5461), .X(n5462) );
  inv_x1_sg U5185 ( .A(n5461), .X(n5463) );
  inv_x1_sg U5186 ( .A(n5461), .X(n5464) );
  inv_x1_sg U5187 ( .A(n5461), .X(n5465) );
  inv_x1_sg U5188 ( .A(n5936), .X(n5466) );
  inv_x1_sg U5189 ( .A(n5466), .X(n5467) );
  inv_x1_sg U5190 ( .A(n5466), .X(n5468) );
  inv_x1_sg U5191 ( .A(n5466), .X(n5469) );
  inv_x1_sg U5192 ( .A(n5466), .X(n5470) );
  inv_x1_sg U5193 ( .A(n4437), .X(n5471) );
  inv_x1_sg U5194 ( .A(n5471), .X(n5472) );
  inv_x1_sg U5195 ( .A(n5471), .X(n5473) );
  inv_x1_sg U5196 ( .A(n5471), .X(n5474) );
  inv_x1_sg U5197 ( .A(n5471), .X(n5475) );
  inv_x1_sg U5198 ( .A(n4464), .X(n5476) );
  inv_x1_sg U5199 ( .A(n5476), .X(n5477) );
  inv_x1_sg U5200 ( .A(n5476), .X(n5478) );
  inv_x1_sg U5201 ( .A(n5476), .X(n5479) );
  inv_x1_sg U5202 ( .A(n4464), .X(n5480) );
  inv_x1_sg U5203 ( .A(n5480), .X(n5481) );
  inv_x1_sg U5204 ( .A(n5480), .X(n5482) );
  inv_x1_sg U5205 ( .A(n5480), .X(n5483) );
  inv_x1_sg U5206 ( .A(n5933), .X(n5484) );
  inv_x1_sg U5207 ( .A(n5484), .X(n5485) );
  inv_x1_sg U5208 ( .A(n5484), .X(n5486) );
  inv_x1_sg U5209 ( .A(n5484), .X(n5487) );
  inv_x1_sg U5210 ( .A(n5484), .X(n5488) );
  inv_x1_sg U5211 ( .A(n5932), .X(n5489) );
  inv_x1_sg U5212 ( .A(n5489), .X(n5490) );
  inv_x1_sg U5213 ( .A(n5489), .X(n5491) );
  inv_x1_sg U5214 ( .A(n5489), .X(n5492) );
  inv_x1_sg U5215 ( .A(n5489), .X(n5493) );
  inv_x1_sg U5216 ( .A(n5935), .X(n5494) );
  inv_x1_sg U5217 ( .A(n5494), .X(n5495) );
  inv_x1_sg U5218 ( .A(n5494), .X(n5496) );
  inv_x1_sg U5219 ( .A(n5494), .X(n5497) );
  inv_x1_sg U5220 ( .A(n5494), .X(n5498) );
  inv_x1_sg U5221 ( .A(n4460), .X(n5499) );
  inv_x1_sg U5222 ( .A(n5499), .X(n5500) );
  inv_x1_sg U5223 ( .A(n5499), .X(n5501) );
  inv_x1_sg U5224 ( .A(n5499), .X(n5502) );
  inv_x1_sg U5225 ( .A(n5499), .X(n5503) );
  inv_x1_sg U5226 ( .A(n4433), .X(n5504) );
  inv_x1_sg U5227 ( .A(n5504), .X(n5505) );
  inv_x1_sg U5228 ( .A(n5504), .X(n5506) );
  inv_x1_sg U5229 ( .A(n5504), .X(n5507) );
  inv_x1_sg U5230 ( .A(n5504), .X(n5508) );
  inv_x1_sg U5231 ( .A(n5934), .X(n5509) );
  inv_x1_sg U5232 ( .A(n5509), .X(n5510) );
  inv_x1_sg U5233 ( .A(n5509), .X(n5511) );
  inv_x1_sg U5234 ( .A(n5509), .X(n5512) );
  inv_x1_sg U5235 ( .A(n5509), .X(n5513) );
  inv_x1_sg U5236 ( .A(n5931), .X(n5514) );
  inv_x1_sg U5237 ( .A(n5514), .X(n5515) );
  inv_x1_sg U5238 ( .A(n5514), .X(n5516) );
  inv_x1_sg U5239 ( .A(n5514), .X(n5517) );
  inv_x1_sg U5240 ( .A(n5514), .X(n5518) );
  inv_x1_sg U5241 ( .A(n5948), .X(n5519) );
  inv_x1_sg U5242 ( .A(n5519), .X(n5520) );
  inv_x1_sg U5243 ( .A(n5519), .X(n5521) );
  inv_x1_sg U5244 ( .A(n5519), .X(n5522) );
  inv_x1_sg U5245 ( .A(n5281), .X(n5523) );
  inv_x1_sg U5246 ( .A(n3520), .X(n5524) );
  inv_x1_sg U5247 ( .A(n5524), .X(n5525) );
  inv_x1_sg U5248 ( .A(n5524), .X(n5526) );
  inv_x1_sg U5249 ( .A(n5524), .X(n5527) );
  inv_x1_sg U5250 ( .A(n5283), .X(n5528) );
  inv_x1_sg U5251 ( .A(n3526), .X(n5529) );
  inv_x1_sg U5252 ( .A(n5529), .X(n5530) );
  inv_x1_sg U5253 ( .A(n5529), .X(n5531) );
  inv_x1_sg U5254 ( .A(n5529), .X(n5532) );
  inv_x1_sg U5255 ( .A(n5285), .X(n5533) );
  inv_x1_sg U5256 ( .A(n3550), .X(n5534) );
  inv_x1_sg U5257 ( .A(n5534), .X(n5535) );
  inv_x1_sg U5258 ( .A(n5534), .X(n5536) );
  inv_x1_sg U5259 ( .A(n5534), .X(n5537) );
  inv_x1_sg U5260 ( .A(n5287), .X(n5538) );
  inv_x1_sg U5261 ( .A(n5541), .X(n5539) );
  inv_x1_sg U5262 ( .A(n4462), .X(n5540) );
  inv_x1_sg U5263 ( .A(n4462), .X(n5541) );
  inv_x1_sg U5264 ( .A(n5540), .X(n5542) );
  inv_x1_sg U5265 ( .A(n5541), .X(n5543) );
  inv_x1_sg U5266 ( .A(n5541), .X(n5544) );
  inv_x1_sg U5267 ( .A(n5541), .X(n5545) );
  inv_x1_sg U5268 ( .A(n5216), .X(n5546) );
  inv_x1_sg U5269 ( .A(n3920), .X(n5547) );
  inv_x1_sg U5270 ( .A(n5216), .X(n5548) );
  inv_x1_sg U5271 ( .A(n5216), .X(n5549) );
  inv_x1_sg U5272 ( .A(n5764), .X(n5550) );
  inv_x1_sg U5273 ( .A(n5550), .X(n5551) );
  inv_x1_sg U5274 ( .A(n5550), .X(n5552) );
  inv_x1_sg U5275 ( .A(n5550), .X(n5553) );
  inv_x1_sg U5276 ( .A(n5550), .X(n5554) );
  inv_x1_sg U5277 ( .A(n5731), .X(n5555) );
  inv_x1_sg U5278 ( .A(n5555), .X(n5556) );
  inv_x1_sg U5279 ( .A(n5555), .X(n5557) );
  inv_x1_sg U5280 ( .A(n5555), .X(n5558) );
  inv_x1_sg U5281 ( .A(n5555), .X(n5559) );
  inv_x1_sg U5282 ( .A(n5672), .X(n5560) );
  inv_x1_sg U5283 ( .A(n5560), .X(n5561) );
  inv_x1_sg U5284 ( .A(n5560), .X(n5562) );
  inv_x1_sg U5285 ( .A(n5560), .X(n5563) );
  inv_x1_sg U5286 ( .A(n5560), .X(n5564) );
  inv_x1_sg U5287 ( .A(n5744), .X(n5565) );
  inv_x1_sg U5288 ( .A(n5565), .X(n5566) );
  inv_x1_sg U5289 ( .A(n5565), .X(n5567) );
  inv_x1_sg U5290 ( .A(n5565), .X(n5568) );
  inv_x1_sg U5291 ( .A(n5565), .X(n5569) );
  inv_x1_sg U5292 ( .A(n5827), .X(n5570) );
  inv_x1_sg U5293 ( .A(n5570), .X(n5571) );
  inv_x1_sg U5294 ( .A(n5570), .X(n5572) );
  inv_x1_sg U5295 ( .A(n5570), .X(n5573) );
  inv_x1_sg U5296 ( .A(n4344), .X(n5574) );
  inv_x1_sg U5297 ( .A(n5828), .X(n5575) );
  inv_x1_sg U5298 ( .A(n5575), .X(n5576) );
  inv_x1_sg U5299 ( .A(n5575), .X(n5577) );
  inv_x1_sg U5300 ( .A(n5575), .X(n5578) );
  inv_x1_sg U5301 ( .A(n5575), .X(n5579) );
  inv_x1_sg U5302 ( .A(n5754), .X(n5580) );
  inv_x1_sg U5303 ( .A(n5580), .X(n5581) );
  inv_x1_sg U5304 ( .A(n5580), .X(n5582) );
  inv_x1_sg U5305 ( .A(n5580), .X(n5583) );
  inv_x1_sg U5306 ( .A(n5580), .X(n5584) );
  inv_x1_sg U5307 ( .A(n5829), .X(n5585) );
  inv_x1_sg U5308 ( .A(n5585), .X(n5586) );
  inv_x1_sg U5309 ( .A(n5585), .X(n5587) );
  inv_x1_sg U5310 ( .A(n5585), .X(n5588) );
  inv_x1_sg U5311 ( .A(n5585), .X(n5589) );
  inv_x1_sg U5312 ( .A(n5661), .X(n5590) );
  inv_x1_sg U5313 ( .A(n5662), .X(n5591) );
  inv_x1_sg U5314 ( .A(n5656), .X(n5592) );
  inv_x1_sg U5315 ( .A(n5951), .X(n5593) );
  inv_x1_sg U5316 ( .A(n5774), .X(n5594) );
  inv_x1_sg U5317 ( .A(n5594), .X(n5595) );
  inv_x1_sg U5318 ( .A(n5594), .X(n5596) );
  inv_x1_sg U5319 ( .A(n5594), .X(n5597) );
  inv_x1_sg U5320 ( .A(n5594), .X(n5598) );
  inv_x1_sg U5321 ( .A(n5830), .X(n5599) );
  inv_x1_sg U5322 ( .A(n5599), .X(n5600) );
  inv_x1_sg U5323 ( .A(n5599), .X(n5601) );
  inv_x1_sg U5324 ( .A(n5599), .X(n5602) );
  inv_x1_sg U5325 ( .A(n5599), .X(n5603) );
  inv_x1_sg U5326 ( .A(n5685), .X(n5604) );
  inv_x1_sg U5327 ( .A(n5604), .X(n5605) );
  inv_x1_sg U5328 ( .A(n5604), .X(n5606) );
  inv_x1_sg U5329 ( .A(n5604), .X(n5607) );
  inv_x1_sg U5330 ( .A(n5604), .X(n5608) );
  inv_x1_sg U5331 ( .A(n5953), .X(n5609) );
  inv_x1_sg U5332 ( .A(n5703), .X(n5610) );
  inv_x1_sg U5333 ( .A(n5953), .X(n5611) );
  inv_x1_sg U5334 ( .A(n5703), .X(n5612) );
  inv_x1_sg U5335 ( .A(n5837), .X(n5613) );
  inv_x1_sg U5336 ( .A(n5613), .X(n5614) );
  inv_x1_sg U5337 ( .A(n5613), .X(n5615) );
  inv_x1_sg U5338 ( .A(n5613), .X(n5616) );
  inv_x1_sg U5339 ( .A(n5613), .X(n5617) );
  inv_x1_sg U5340 ( .A(n5811), .X(n5618) );
  inv_x1_sg U5341 ( .A(n5618), .X(n5619) );
  inv_x1_sg U5342 ( .A(n5618), .X(n5620) );
  inv_x1_sg U5343 ( .A(n5618), .X(n5621) );
  inv_x1_sg U5344 ( .A(n5618), .X(n5622) );
  inv_x1_sg U5345 ( .A(n5838), .X(n5623) );
  inv_x1_sg U5346 ( .A(n5623), .X(n5624) );
  inv_x1_sg U5347 ( .A(n5623), .X(n5625) );
  inv_x1_sg U5348 ( .A(n5623), .X(n5626) );
  inv_x1_sg U5349 ( .A(n5623), .X(n5627) );
  inv_x1_sg U5350 ( .A(n5716), .X(n5628) );
  inv_x1_sg U5351 ( .A(n5628), .X(n5629) );
  inv_x1_sg U5352 ( .A(n5628), .X(n5630) );
  inv_x1_sg U5353 ( .A(n5628), .X(n5631) );
  inv_x1_sg U5354 ( .A(n5628), .X(n5632) );
  inv_x1_sg U5355 ( .A(n5797), .X(n5633) );
  inv_x1_sg U5356 ( .A(n5633), .X(n5634) );
  inv_x1_sg U5357 ( .A(n5633), .X(n5635) );
  inv_x1_sg U5358 ( .A(n5633), .X(n5636) );
  inv_x1_sg U5359 ( .A(n5633), .X(n5637) );
  inv_x1_sg U5360 ( .A(n5784), .X(n5638) );
  inv_x1_sg U5361 ( .A(n5638), .X(n5639) );
  inv_x1_sg U5362 ( .A(n5638), .X(n5640) );
  inv_x1_sg U5363 ( .A(n5638), .X(n5641) );
  inv_x1_sg U5364 ( .A(n5638), .X(n5642) );
  inv_x1_sg U5365 ( .A(n3547), .X(n5643) );
  inv_x1_sg U5366 ( .A(n5643), .X(n5644) );
  inv_x1_sg U5367 ( .A(n5643), .X(n5645) );
  inv_x1_sg U5368 ( .A(n5643), .X(n5646) );
  inv_x1_sg U5369 ( .A(n5309), .X(n5647) );
  inv_x1_sg U5370 ( .A(n5946), .X(n5648) );
  inv_x1_sg U5371 ( .A(n5648), .X(n5649) );
  inv_x1_sg U5372 ( .A(n5648), .X(n5650) );
  inv_x1_sg U5373 ( .A(n5648), .X(n5651) );
  inv_x1_sg U5374 ( .A(n5311), .X(n5652) );
  inv_x4_sg U5375 ( .A(n5951), .X(n5653) );
  inv_x1_sg U5376 ( .A(n5653), .X(n5654) );
  inv_x1_sg U5377 ( .A(n5653), .X(n5655) );
  inv_x1_sg U5378 ( .A(n5653), .X(n5656) );
  inv_x1_sg U5379 ( .A(n5657), .X(n5658) );
  inv_x1_sg U5380 ( .A(n5657), .X(n5659) );
  inv_x1_sg U5381 ( .A(n5660), .X(n5661) );
  inv_x1_sg U5382 ( .A(n5660), .X(n5662) );
  inv_x1_sg U5383 ( .A(n4344), .X(n5663) );
  inv_x1_sg U5384 ( .A(n5827), .X(n5664) );
  inv_x1_sg U5385 ( .A(n5663), .X(n5665) );
  inv_x1_sg U5386 ( .A(n5663), .X(n5666) );
  inv_x1_sg U5387 ( .A(n5663), .X(n5667) );
  inv_x1_sg U5388 ( .A(n5669), .X(n5670) );
  inv_x1_sg U5389 ( .A(n5669), .X(n5671) );
  inv_x4_sg U5390 ( .A(n5893), .X(n5672) );
  inv_x1_sg U5391 ( .A(n5672), .X(n5673) );
  inv_x1_sg U5392 ( .A(n5672), .X(n5674) );
  inv_x1_sg U5393 ( .A(n5672), .X(n5675) );
  inv_x1_sg U5394 ( .A(n5885), .X(n5676) );
  inv_x1_sg U5395 ( .A(n5838), .X(n5677) );
  inv_x1_sg U5396 ( .A(n5676), .X(n5678) );
  inv_x1_sg U5397 ( .A(n5676), .X(n5679) );
  inv_x1_sg U5398 ( .A(n5676), .X(n5680) );
  nand_x4_sg U5399 ( .A(n5901), .B(n3873), .X(n5681) );
  inv_x1_sg U5400 ( .A(n5685), .X(n5682) );
  inv_x1_sg U5401 ( .A(n5686), .X(n5683) );
  inv_x1_sg U5402 ( .A(n5686), .X(n5684) );
  inv_x4_sg U5403 ( .A(n5954), .X(n5685) );
  inv_x1_sg U5404 ( .A(n5682), .X(n5686) );
  inv_x1_sg U5405 ( .A(n5685), .X(n5687) );
  inv_x1_sg U5406 ( .A(n5685), .X(n5688) );
  inv_x1_sg U5407 ( .A(n5686), .X(n5689) );
  inv_x1_sg U5408 ( .A(n5686), .X(n5690) );
  nand_x8_sg U5409 ( .A(n5839), .B(n3873), .X(n5954) );
  inv_x1_sg U5410 ( .A(n4399), .X(n5691) );
  inv_x1_sg U5411 ( .A(n4399), .X(n5692) );
  inv_x1_sg U5412 ( .A(n5691), .X(n5693) );
  inv_x1_sg U5413 ( .A(n5691), .X(n5694) );
  inv_x1_sg U5414 ( .A(n5692), .X(n5695) );
  inv_x1_sg U5415 ( .A(n5692), .X(n5696) );
  inv_x1_sg U5416 ( .A(n5692), .X(n5697) );
  inv_x1_sg U5417 ( .A(n4260), .X(n5698) );
  inv_x1_sg U5418 ( .A(n5828), .X(n5699) );
  inv_x1_sg U5419 ( .A(n5698), .X(n5700) );
  inv_x1_sg U5420 ( .A(n5698), .X(n5701) );
  inv_x1_sg U5421 ( .A(n5698), .X(n5702) );
  nand_x1_sg U5422 ( .A(n5839), .B(n3917), .X(n5703) );
  inv_x1_sg U5423 ( .A(n5703), .X(n5704) );
  inv_x1_sg U5424 ( .A(n5704), .X(n5705) );
  inv_x1_sg U5425 ( .A(n5704), .X(n5706) );
  inv_x1_sg U5426 ( .A(n5704), .X(n5707) );
  inv_x1_sg U5427 ( .A(n5953), .X(n5708) );
  inv_x1_sg U5428 ( .A(n5708), .X(n5709) );
  inv_x1_sg U5429 ( .A(n5708), .X(n5710) );
  inv_x1_sg U5430 ( .A(n5708), .X(n5711) );
  nand_x1_sg U5431 ( .A(n5928), .B(n3917), .X(n5953) );
  nand_x4_sg U5432 ( .A(n5928), .B(n4171), .X(n5712) );
  inv_x1_sg U5433 ( .A(n5716), .X(n5713) );
  inv_x1_sg U5434 ( .A(n5717), .X(n5714) );
  inv_x1_sg U5435 ( .A(n5717), .X(n5715) );
  inv_x4_sg U5436 ( .A(n5950), .X(n5716) );
  inv_x1_sg U5437 ( .A(n5713), .X(n5717) );
  inv_x1_sg U5438 ( .A(n5716), .X(n5718) );
  inv_x1_sg U5439 ( .A(n5716), .X(n5719) );
  inv_x1_sg U5440 ( .A(n5717), .X(n5720) );
  inv_x1_sg U5441 ( .A(n5717), .X(n5721) );
  nand_x8_sg U5442 ( .A(n5927), .B(n4171), .X(n5950) );
  inv_x1_sg U5443 ( .A(n5949), .X(n5722) );
  inv_x1_sg U5444 ( .A(n5829), .X(n5723) );
  inv_x1_sg U5445 ( .A(n5722), .X(n5724) );
  inv_x1_sg U5446 ( .A(n5722), .X(n5725) );
  inv_x1_sg U5447 ( .A(n5722), .X(n5726) );
  inv_x1_sg U5448 ( .A(n5728), .X(n5729) );
  inv_x1_sg U5449 ( .A(n5728), .X(n5730) );
  inv_x4_sg U5450 ( .A(n5955), .X(n5731) );
  inv_x1_sg U5451 ( .A(n5731), .X(n5732) );
  inv_x1_sg U5452 ( .A(n5731), .X(n5733) );
  inv_x1_sg U5453 ( .A(n5731), .X(n5734) );
  inv_x1_sg U5454 ( .A(n5886), .X(n5735) );
  inv_x1_sg U5455 ( .A(n5830), .X(n5736) );
  inv_x1_sg U5456 ( .A(n5735), .X(n5737) );
  inv_x1_sg U5457 ( .A(n5735), .X(n5738) );
  inv_x1_sg U5458 ( .A(n5735), .X(n5739) );
  nand_x4_sg U5459 ( .A(n5930), .B(n3575), .X(n5740) );
  inv_x1_sg U5460 ( .A(n5744), .X(n5741) );
  inv_x1_sg U5461 ( .A(n5745), .X(n5742) );
  inv_x1_sg U5462 ( .A(n5745), .X(n5743) );
  inv_x4_sg U5463 ( .A(n3517), .X(n5744) );
  inv_x1_sg U5464 ( .A(n5741), .X(n5745) );
  inv_x1_sg U5465 ( .A(n5744), .X(n5746) );
  inv_x1_sg U5466 ( .A(n5744), .X(n5747) );
  inv_x1_sg U5467 ( .A(n5745), .X(n5748) );
  inv_x1_sg U5468 ( .A(n5745), .X(n5749) );
  nand_x8_sg U5469 ( .A(n5896), .B(n3575), .X(n3517) );
  nand_x4_sg U5470 ( .A(n5895), .B(n4043), .X(n5750) );
  inv_x1_sg U5471 ( .A(n5754), .X(n5751) );
  inv_x1_sg U5472 ( .A(n5755), .X(n5752) );
  inv_x1_sg U5473 ( .A(n5755), .X(n5753) );
  inv_x4_sg U5474 ( .A(n5952), .X(n5754) );
  inv_x1_sg U5475 ( .A(n5751), .X(n5755) );
  inv_x1_sg U5476 ( .A(n5754), .X(n5756) );
  inv_x1_sg U5477 ( .A(n5754), .X(n5757) );
  inv_x1_sg U5478 ( .A(n5755), .X(n5758) );
  inv_x1_sg U5479 ( .A(n5755), .X(n5759) );
  nand_x8_sg U5480 ( .A(n5897), .B(n4043), .X(n5952) );
  nand_x4_sg U5481 ( .A(n5898), .B(n4257), .X(n5760) );
  inv_x1_sg U5482 ( .A(n5764), .X(n5761) );
  inv_x1_sg U5483 ( .A(n5765), .X(n5762) );
  inv_x1_sg U5484 ( .A(n5765), .X(n5763) );
  inv_x4_sg U5485 ( .A(n4218), .X(n5764) );
  inv_x1_sg U5486 ( .A(n5761), .X(n5765) );
  inv_x1_sg U5487 ( .A(n5764), .X(n5766) );
  inv_x1_sg U5488 ( .A(n5764), .X(n5767) );
  inv_x1_sg U5489 ( .A(n5765), .X(n5768) );
  inv_x1_sg U5490 ( .A(n5765), .X(n5769) );
  nand_x8_sg U5491 ( .A(n5899), .B(n4257), .X(n4218) );
  nand_x4_sg U5492 ( .A(n5839), .B(n4087), .X(n5770) );
  inv_x1_sg U5493 ( .A(n5774), .X(n5771) );
  inv_x1_sg U5494 ( .A(n5775), .X(n5772) );
  inv_x1_sg U5495 ( .A(n5775), .X(n5773) );
  inv_x4_sg U5496 ( .A(n5889), .X(n5774) );
  inv_x1_sg U5497 ( .A(n5771), .X(n5775) );
  inv_x1_sg U5498 ( .A(n5774), .X(n5776) );
  inv_x1_sg U5499 ( .A(n5774), .X(n5777) );
  inv_x1_sg U5500 ( .A(n5775), .X(n5778) );
  inv_x1_sg U5501 ( .A(n5775), .X(n5779) );
  nand_x8_sg U5502 ( .A(n5928), .B(n4087), .X(n5889) );
  inv_x1_sg U5503 ( .A(n5781), .X(n5782) );
  inv_x1_sg U5504 ( .A(n5781), .X(n5783) );
  inv_x4_sg U5505 ( .A(n3962), .X(n5784) );
  inv_x1_sg U5506 ( .A(n5784), .X(n5785) );
  inv_x1_sg U5507 ( .A(n5784), .X(n5786) );
  inv_x1_sg U5508 ( .A(n5784), .X(n5787) );
  inv_x1_sg U5509 ( .A(n3621), .X(n5788) );
  inv_x1_sg U5510 ( .A(n5837), .X(n5789) );
  inv_x1_sg U5511 ( .A(n5788), .X(n5790) );
  inv_x1_sg U5512 ( .A(n5788), .X(n5791) );
  inv_x1_sg U5513 ( .A(n5788), .X(n5792) );
  nand_x4_sg U5514 ( .A(n5929), .B(n3747), .X(n5793) );
  inv_x1_sg U5515 ( .A(n5797), .X(n5794) );
  inv_x1_sg U5516 ( .A(n5798), .X(n5795) );
  inv_x1_sg U5517 ( .A(n5798), .X(n5796) );
  inv_x4_sg U5518 ( .A(n5956), .X(n5797) );
  inv_x1_sg U5519 ( .A(n5794), .X(n5798) );
  inv_x1_sg U5520 ( .A(n5797), .X(n5799) );
  inv_x1_sg U5521 ( .A(n5797), .X(n5800) );
  inv_x1_sg U5522 ( .A(n5798), .X(n5801) );
  inv_x1_sg U5523 ( .A(n5798), .X(n5802) );
  nand_x8_sg U5524 ( .A(n5930), .B(n3747), .X(n5956) );
  inv_x1_sg U5525 ( .A(n5807), .X(n5804) );
  inv_x1_sg U5526 ( .A(n5811), .X(n5805) );
  inv_x1_sg U5527 ( .A(n5811), .X(n5806) );
  inv_x4_sg U5528 ( .A(n5803), .X(n5807) );
  inv_x1_sg U5529 ( .A(n5807), .X(n5808) );
  inv_x1_sg U5530 ( .A(n5807), .X(n5809) );
  inv_x1_sg U5531 ( .A(n5807), .X(n5810) );
  inv_x2_sg U5532 ( .A(n5803), .X(n5811) );
  inv_x1_sg U5533 ( .A(n5333), .X(n5812) );
  inv_x1_sg U5534 ( .A(n5812), .X(n5813) );
  inv_x1_sg U5535 ( .A(n5812), .X(n5814) );
  inv_x1_sg U5536 ( .A(n4406), .X(n5815) );
  inv_x1_sg U5537 ( .A(n5812), .X(n5816) );
  inv_x1_sg U5538 ( .A(n5943), .X(n5817) );
  inv_x1_sg U5539 ( .A(n5943), .X(n5818) );
  inv_x1_sg U5540 ( .A(n5817), .X(n5819) );
  inv_x1_sg U5541 ( .A(n5817), .X(n5820) );
  inv_x1_sg U5542 ( .A(n5817), .X(n5821) );
  inv_x1_sg U5543 ( .A(n5818), .X(n5822) );
  inv_x1_sg U5544 ( .A(n5818), .X(n5823) );
  inv_x1_sg U5545 ( .A(n5818), .X(n5824) );
  nand_x8_sg U5546 ( .A(n5900), .B(n4001), .X(n3962) );
  nand_x8_sg U5547 ( .A(n5895), .B(n3831), .X(n5955) );
  nand_x8_sg U5548 ( .A(n5898), .B(n3959), .X(n3920) );
  inv_x16_sg U5549 ( .A(reset), .X(n5839) );
  nor_x1_sg U5550 ( .A(n3276), .B(n5820), .X(n5946) );
  nor_x1_sg U5551 ( .A(n3275), .B(n5823), .X(n3547) );
  nor_x1_sg U5552 ( .A(n5890), .B(n5821), .X(n5947) );
  nor_x1_sg U5553 ( .A(n3273), .B(n5820), .X(n5945) );
  nor_x1_sg U5554 ( .A(n3269), .B(n5822), .X(n5944) );
  nor_x1_sg U5555 ( .A(n3277), .B(n5819), .X(n3541) );
  nor_x1_sg U5556 ( .A(n3266), .B(n5822), .X(n3574) );
  nor_x1_sg U5557 ( .A(n3335), .B(n5181), .X(n5937) );
  nor_x1_sg U5558 ( .A(n5191), .B(n3335), .X(n4445) );
  nor_x1_sg U5559 ( .A(n5836), .B(reset), .X(n3465) );
  nor_x1_sg U5560 ( .A(n5181), .B(n5831), .X(n4399) );
  inv_x1_sg U5561 ( .A(wr_ptr[4]), .X(n5826) );
  inv_x1_sg U5562 ( .A(n4344), .X(n5827) );
  inv_x1_sg U5563 ( .A(n4260), .X(n5828) );
  inv_x1_sg U5564 ( .A(n5949), .X(n5829) );
  inv_x1_sg U5565 ( .A(n5886), .X(n5830) );
  inv_x1_sg U5566 ( .A(n4396), .X(n5831) );
  inv_x1_sg U5567 ( .A(rd_ptr[1]), .X(n5832) );
  inv_x1_sg U5568 ( .A(wr_ptr[0]), .X(n5833) );
  inv_x1_sg U5569 ( .A(wr_ptr[1]), .X(n5834) );
  inv_x1_sg U5570 ( .A(n3474), .X(n5835) );
  inv_x1_sg U5571 ( .A(n5943), .X(n5836) );
  inv_x1_sg U5572 ( .A(n3621), .X(n5837) );
  inv_x1_sg U5573 ( .A(n5885), .X(n5838) );
  nand_x1_sg U5574 ( .A(n3875), .B(n3705), .X(n5840) );
  nand_x1_sg U5575 ( .A(n4215), .B(n3705), .X(n5841) );
  inv_x1_sg U5576 ( .A(n5843), .X(n5842) );
  nand_x4_sg U5577 ( .A(n5897), .B(n4341), .X(n5885) );
  nand_x16_sg U5578 ( .A(n5319), .B(rd_en), .X(n5843) );
  nor_x1_sg U5579 ( .A(reset), .B(empty), .X(n5168) );
  nand_x4_sg U5580 ( .A(n4386), .B(n4387), .X(n5943) );
  inv_x1_sg U5581 ( .A(n5192), .X(n5844) );
  inv_x1_sg U5582 ( .A(n5146), .X(n5845) );
  inv_x1_sg U5583 ( .A(n5107), .X(n5846) );
  inv_x1_sg U5584 ( .A(n5068), .X(n5847) );
  inv_x1_sg U5585 ( .A(n5029), .X(n5848) );
  inv_x1_sg U5586 ( .A(n4990), .X(n5849) );
  inv_x1_sg U5587 ( .A(n4951), .X(n5850) );
  inv_x1_sg U5588 ( .A(n4912), .X(n5851) );
  inv_x1_sg U5589 ( .A(n4873), .X(n5852) );
  inv_x1_sg U5590 ( .A(n4834), .X(n5853) );
  inv_x1_sg U5591 ( .A(n4795), .X(n5854) );
  inv_x1_sg U5592 ( .A(n4756), .X(n5855) );
  inv_x1_sg U5593 ( .A(n4717), .X(n5856) );
  inv_x1_sg U5594 ( .A(n4678), .X(n5857) );
  inv_x1_sg U5595 ( .A(n4639), .X(n5858) );
  inv_x1_sg U5596 ( .A(n4600), .X(n5859) );
  inv_x1_sg U5597 ( .A(n4561), .X(n5860) );
  inv_x1_sg U5598 ( .A(n4522), .X(n5861) );
  inv_x1_sg U5599 ( .A(n4483), .X(n5862) );
  inv_x1_sg U5600 ( .A(n4434), .X(n5863) );
  inv_x1_sg U5601 ( .A(n5203), .X(n5864) );
  inv_x1_sg U5602 ( .A(n5156), .X(n5865) );
  inv_x1_sg U5603 ( .A(n5117), .X(n5866) );
  inv_x1_sg U5604 ( .A(n5078), .X(n5867) );
  inv_x1_sg U5605 ( .A(n5039), .X(n5868) );
  inv_x1_sg U5606 ( .A(n5000), .X(n5869) );
  inv_x1_sg U5607 ( .A(n4961), .X(n5870) );
  inv_x1_sg U5608 ( .A(n4922), .X(n5871) );
  inv_x1_sg U5609 ( .A(n4883), .X(n5872) );
  inv_x1_sg U5610 ( .A(n4844), .X(n5873) );
  inv_x1_sg U5611 ( .A(n4805), .X(n5874) );
  inv_x1_sg U5612 ( .A(n4766), .X(n5875) );
  inv_x1_sg U5613 ( .A(n4727), .X(n5876) );
  inv_x1_sg U5614 ( .A(n4688), .X(n5877) );
  inv_x1_sg U5615 ( .A(n4649), .X(n5878) );
  inv_x1_sg U5616 ( .A(n4610), .X(n5879) );
  inv_x1_sg U5617 ( .A(n4571), .X(n5880) );
  inv_x1_sg U5618 ( .A(n4532), .X(n5881) );
  inv_x1_sg U5619 ( .A(n4493), .X(n5882) );
  inv_x1_sg U5620 ( .A(n4448), .X(n5883) );
  inv_x8_sg U5621 ( .A(data_in[7]), .X(n3278) );
  inv_x8_sg U5622 ( .A(data_in[18]), .X(n5884) );
  inv_x8_sg U5623 ( .A(reset), .X(n5929) );
  inv_x16_sg U5624 ( .A(reset), .X(n5928) );
  nand_x8_sg U5625 ( .A(n5214), .B(n3702), .X(n5893) );
  inv_x1_sg U5626 ( .A(n5841), .X(n5887) );
  nand_x1_sg U5627 ( .A(rd_ptr[0]), .B(n5832), .X(n5888) );
  inv_x8_sg U5628 ( .A(data_in[6]), .X(n5891) );
  nor_x1_sg U5629 ( .A(n5894), .B(n5820), .X(n5903) );
  inv_x16_sg U5630 ( .A(reset), .X(n5895) );
  inv_x16_sg U5631 ( .A(reset), .X(n5896) );
  inv_x16_sg U5632 ( .A(reset), .X(n5897) );
  inv_x16_sg U5633 ( .A(reset), .X(n5898) );
  inv_x16_sg U5634 ( .A(reset), .X(n5899) );
  inv_x16_sg U5635 ( .A(reset), .X(n5900) );
  inv_x16_sg U5636 ( .A(reset), .X(n5901) );
  inv_x16_sg U5637 ( .A(reset), .X(n5927) );
  inv_x16_sg U5638 ( .A(reset), .X(n5930) );
  nor_x1_sg U5639 ( .A(n5891), .B(n5824), .X(n5902) );
  nor_x1_sg U5640 ( .A(n5884), .B(n5822), .X(n5904) );
  nor_x1_sg U5641 ( .A(n5892), .B(n5819), .X(n5905) );
  inv_x1_sg U5642 ( .A(n5921), .X(n5906) );
  inv_x1_sg U5643 ( .A(rd_ptr[2]), .X(n5907) );
  inv_x8_sg U5644 ( .A(data_in[17]), .X(n5911) );
  inv_x8_sg U5645 ( .A(data_in[15]), .X(n5912) );
  nand_x16_sg U5646 ( .A(n5319), .B(rd_en), .X(n5942) );
  nor_x1_sg U5647 ( .A(n5842), .B(reset), .X(n5913) );
  nand_x1_sg U5648 ( .A(n5178), .B(n5184), .X(n5914) );
  nand_x1_sg U5649 ( .A(rd_ptr[2]), .B(n3371), .X(n5181) );
  nand_x1_sg U5650 ( .A(rd_ptr[3]), .B(n5907), .X(n5191) );
  inv_x1_sg U5651 ( .A(wr_ptr[2]), .X(n5915) );
  inv_x1_sg U5652 ( .A(n4407), .X(n5916) );
  inv_x1_sg U5653 ( .A(n5920), .X(n5917) );
  nand_x16_sg U5654 ( .A(n5168), .B(rd_en), .X(n4407) );
  inv_x1_sg U5655 ( .A(n5178), .X(n5918) );
  nand_x1_sg U5656 ( .A(n5832), .B(n3333), .X(n5177) );
  inv_x8_sg U5657 ( .A(wr_en), .X(n3287) );
  inv_x8_sg U5658 ( .A(rd_en), .X(n3286) );
  nand_x16_sg U5659 ( .A(n5319), .B(rd_en), .X(n5920) );
  nand_x16_sg U5660 ( .A(n5168), .B(rd_en), .X(n5921) );
  nand_x16_sg U5661 ( .A(n5319), .B(rd_en), .X(n5941) );
  nor_x1_sg U5662 ( .A(n3272), .B(n5821), .X(n5922) );
  nor_x1_sg U5663 ( .A(n3278), .B(n5823), .X(n5923) );
  nor_x1_sg U5664 ( .A(n5910), .B(n5821), .X(n5924) );
  nor_x1_sg U5665 ( .A(n5911), .B(n5823), .X(n5925) );
  nor_x1_sg U5666 ( .A(n5912), .B(n5824), .X(n5926) );
  inv_x1_sg U5667 ( .A(n5840), .X(n3261) );
  inv_x1_sg U5668 ( .A(n4044), .X(n3260) );
  inv_x1_sg U5669 ( .A(n4384), .X(n3258) );
  inv_x1_sg U5670 ( .A(n3703), .X(n3262) );
  inv_x1_sg U5671 ( .A(n3500), .X(n3334) );
  inv_x1_sg U5672 ( .A(n3508), .X(n3311) );
  inv_x1_sg U5673 ( .A(n3455), .X(n3360) );
  nand_x1_sg U5674 ( .A(n3502), .B(n3503), .X(n3448) );
  nor_x1_sg U5675 ( .A(n4388), .B(n3287), .X(n4386) );
  inv_x1_sg U5676 ( .A(n5213), .X(n3336) );
  nand_x1_sg U5677 ( .A(n5204), .B(n5205), .X(n5203) );
  nand_x1_sg U5678 ( .A(n5193), .B(n5194), .X(n5192) );
  inv_x1_sg U5679 ( .A(n5166), .X(n3337) );
  nand_x1_sg U5680 ( .A(n5157), .B(n5158), .X(n5156) );
  nand_x1_sg U5681 ( .A(n5147), .B(n5148), .X(n5146) );
  inv_x1_sg U5682 ( .A(n5127), .X(n3338) );
  nand_x1_sg U5683 ( .A(n5118), .B(n5119), .X(n5117) );
  nand_x1_sg U5684 ( .A(n5108), .B(n5109), .X(n5107) );
  inv_x1_sg U5685 ( .A(n5088), .X(n3339) );
  nand_x1_sg U5686 ( .A(n5079), .B(n5080), .X(n5078) );
  nand_x1_sg U5687 ( .A(n5069), .B(n5070), .X(n5068) );
  inv_x1_sg U5688 ( .A(n5049), .X(n3340) );
  nand_x1_sg U5689 ( .A(n5040), .B(n5041), .X(n5039) );
  nand_x1_sg U5690 ( .A(n5030), .B(n5031), .X(n5029) );
  inv_x1_sg U5691 ( .A(n5010), .X(n3341) );
  nand_x1_sg U5692 ( .A(n5001), .B(n5002), .X(n5000) );
  nand_x1_sg U5693 ( .A(n4991), .B(n4992), .X(n4990) );
  inv_x1_sg U5694 ( .A(n4971), .X(n3342) );
  nand_x1_sg U5695 ( .A(n4962), .B(n4963), .X(n4961) );
  nand_x1_sg U5696 ( .A(n4952), .B(n4953), .X(n4951) );
  inv_x1_sg U5697 ( .A(n4932), .X(n3343) );
  nand_x1_sg U5698 ( .A(n4923), .B(n4924), .X(n4922) );
  nand_x1_sg U5699 ( .A(n4913), .B(n4914), .X(n4912) );
  inv_x1_sg U5700 ( .A(n4893), .X(n3344) );
  nand_x1_sg U5701 ( .A(n4884), .B(n4885), .X(n4883) );
  nand_x1_sg U5702 ( .A(n4874), .B(n4875), .X(n4873) );
  inv_x1_sg U5703 ( .A(n4854), .X(n3345) );
  nand_x1_sg U5704 ( .A(n4845), .B(n4846), .X(n4844) );
  nand_x1_sg U5705 ( .A(n4835), .B(n4836), .X(n4834) );
  inv_x1_sg U5706 ( .A(n4815), .X(n3346) );
  nand_x1_sg U5707 ( .A(n4806), .B(n4807), .X(n4805) );
  nand_x1_sg U5708 ( .A(n4796), .B(n4797), .X(n4795) );
  inv_x1_sg U5709 ( .A(n4776), .X(n3347) );
  nand_x1_sg U5710 ( .A(n4767), .B(n4768), .X(n4766) );
  nand_x1_sg U5711 ( .A(n4757), .B(n4758), .X(n4756) );
  inv_x1_sg U5712 ( .A(n4737), .X(n3348) );
  nand_x1_sg U5713 ( .A(n4728), .B(n4729), .X(n4727) );
  nand_x1_sg U5714 ( .A(n4718), .B(n4719), .X(n4717) );
  inv_x1_sg U5715 ( .A(n4698), .X(n3349) );
  nand_x1_sg U5716 ( .A(n4689), .B(n4690), .X(n4688) );
  nand_x1_sg U5717 ( .A(n4679), .B(n4680), .X(n4678) );
  inv_x1_sg U5718 ( .A(n4659), .X(n3350) );
  nand_x1_sg U5719 ( .A(n4650), .B(n4651), .X(n4649) );
  nand_x1_sg U5720 ( .A(n4640), .B(n4641), .X(n4639) );
  inv_x1_sg U5721 ( .A(n4620), .X(n3351) );
  nand_x1_sg U5722 ( .A(n4611), .B(n4612), .X(n4610) );
  nand_x1_sg U5723 ( .A(n4601), .B(n4602), .X(n4600) );
  inv_x1_sg U5724 ( .A(n4581), .X(n3352) );
  nand_x1_sg U5725 ( .A(n4572), .B(n4573), .X(n4571) );
  nand_x1_sg U5726 ( .A(n4562), .B(n4563), .X(n4561) );
  inv_x1_sg U5727 ( .A(n4542), .X(n3353) );
  nand_x1_sg U5728 ( .A(n4533), .B(n4534), .X(n4532) );
  nand_x1_sg U5729 ( .A(n4523), .B(n4524), .X(n4522) );
  inv_x1_sg U5730 ( .A(n4503), .X(n3354) );
  nand_x1_sg U5731 ( .A(n4494), .B(n4495), .X(n4493) );
  nand_x1_sg U5732 ( .A(n4484), .B(n4485), .X(n4483) );
  inv_x1_sg U5733 ( .A(n4463), .X(n3355) );
  nand_x1_sg U5734 ( .A(n4449), .B(n4450), .X(n4448) );
  nand_x1_sg U5735 ( .A(n4435), .B(n4436), .X(n4434) );
  nor_x1_sg U5736 ( .A(n4399), .B(n4400), .X(n3497) );
  nand_x1_sg U5737 ( .A(n3448), .B(n3501), .X(n3491) );
  nand_x1_sg U5738 ( .A(n3493), .B(n3494), .X(n3492) );
  nand_x1_sg U5739 ( .A(n3495), .B(n3496), .X(n3494) );
  nor_x1_sg U5740 ( .A(n3504), .B(n3505), .X(n3489) );
  nor_x1_sg U5741 ( .A(n3482), .B(n3483), .X(n3462) );
  nor_x1_sg U5742 ( .A(n3472), .B(n3473), .X(n3459) );
  nand_x1_sg U5743 ( .A(n3460), .B(n3461), .X(n3450) );
  nand_x1_sg U5744 ( .A(n3452), .B(n3453), .X(n3451) );
  nor_x1_sg U5745 ( .A(n5206), .B(n5207), .X(n5195) );
  nand_x1_sg U5746 ( .A(n5210), .B(n5211), .X(n5206) );
  nor_x1_sg U5747 ( .A(n5197), .B(n5198), .X(n5196) );
  nand_x1_sg U5748 ( .A(n5199), .B(n5200), .X(n5198) );
  nor_x1_sg U5749 ( .A(n5173), .B(n5174), .X(n5172) );
  nand_x1_sg U5750 ( .A(n5179), .B(n5180), .X(n5173) );
  nor_x1_sg U5751 ( .A(n5186), .B(n5187), .X(n5171) );
  nand_x1_sg U5752 ( .A(n5188), .B(n5189), .X(n5187) );
  nor_x1_sg U5753 ( .A(n5159), .B(n5160), .X(n5149) );
  nand_x1_sg U5754 ( .A(n5163), .B(n5164), .X(n5159) );
  nor_x1_sg U5755 ( .A(n5151), .B(n5152), .X(n5150) );
  nand_x1_sg U5756 ( .A(n5153), .B(n5154), .X(n5152) );
  nor_x1_sg U5757 ( .A(n5133), .B(n5134), .X(n5132) );
  nand_x1_sg U5758 ( .A(n5137), .B(n5138), .X(n5133) );
  nor_x1_sg U5759 ( .A(n5141), .B(n5142), .X(n5131) );
  nand_x1_sg U5760 ( .A(n5143), .B(n5144), .X(n5142) );
  nor_x1_sg U5761 ( .A(n5120), .B(n5121), .X(n5110) );
  nand_x1_sg U5762 ( .A(n5124), .B(n5125), .X(n5120) );
  nor_x1_sg U5763 ( .A(n5112), .B(n5113), .X(n5111) );
  nand_x1_sg U5764 ( .A(n5114), .B(n5115), .X(n5113) );
  nor_x1_sg U5765 ( .A(n5094), .B(n5095), .X(n5093) );
  nand_x1_sg U5766 ( .A(n5098), .B(n5099), .X(n5094) );
  nor_x1_sg U5767 ( .A(n5102), .B(n5103), .X(n5092) );
  nand_x1_sg U5768 ( .A(n5104), .B(n5105), .X(n5103) );
  nor_x1_sg U5769 ( .A(n5081), .B(n5082), .X(n5071) );
  nand_x1_sg U5770 ( .A(n5085), .B(n5086), .X(n5081) );
  nor_x1_sg U5771 ( .A(n5073), .B(n5074), .X(n5072) );
  nand_x1_sg U5772 ( .A(n5075), .B(n5076), .X(n5074) );
  nor_x1_sg U5773 ( .A(n5055), .B(n5056), .X(n5054) );
  nand_x1_sg U5774 ( .A(n5059), .B(n5060), .X(n5055) );
  nor_x1_sg U5775 ( .A(n5063), .B(n5064), .X(n5053) );
  nand_x1_sg U5776 ( .A(n5065), .B(n5066), .X(n5064) );
  nor_x1_sg U5777 ( .A(n5042), .B(n5043), .X(n5032) );
  nand_x1_sg U5778 ( .A(n5046), .B(n5047), .X(n5042) );
  nor_x1_sg U5779 ( .A(n5034), .B(n5035), .X(n5033) );
  nand_x1_sg U5780 ( .A(n5036), .B(n5037), .X(n5035) );
  nor_x1_sg U5781 ( .A(n5016), .B(n5017), .X(n5015) );
  nand_x1_sg U5782 ( .A(n5020), .B(n5021), .X(n5016) );
  nor_x1_sg U5783 ( .A(n5024), .B(n5025), .X(n5014) );
  nand_x1_sg U5784 ( .A(n5026), .B(n5027), .X(n5025) );
  nor_x1_sg U5785 ( .A(n5003), .B(n5004), .X(n4993) );
  nand_x1_sg U5786 ( .A(n5007), .B(n5008), .X(n5003) );
  nor_x1_sg U5787 ( .A(n4995), .B(n4996), .X(n4994) );
  nand_x1_sg U5788 ( .A(n4997), .B(n4998), .X(n4996) );
  nor_x1_sg U5789 ( .A(n4977), .B(n4978), .X(n4976) );
  nand_x1_sg U5790 ( .A(n4981), .B(n4982), .X(n4977) );
  nor_x1_sg U5791 ( .A(n4985), .B(n4986), .X(n4975) );
  nand_x1_sg U5792 ( .A(n4987), .B(n4988), .X(n4986) );
  nor_x1_sg U5793 ( .A(n4964), .B(n4965), .X(n4954) );
  nand_x1_sg U5794 ( .A(n4968), .B(n4969), .X(n4964) );
  nor_x1_sg U5795 ( .A(n4956), .B(n4957), .X(n4955) );
  nand_x1_sg U5796 ( .A(n4958), .B(n4959), .X(n4957) );
  nor_x1_sg U5797 ( .A(n4938), .B(n4939), .X(n4937) );
  nand_x1_sg U5798 ( .A(n4942), .B(n4943), .X(n4938) );
  nor_x1_sg U5799 ( .A(n4946), .B(n4947), .X(n4936) );
  nand_x1_sg U5800 ( .A(n4948), .B(n4949), .X(n4947) );
  nor_x1_sg U5801 ( .A(n4925), .B(n4926), .X(n4915) );
  nand_x1_sg U5802 ( .A(n4929), .B(n4930), .X(n4925) );
  nor_x1_sg U5803 ( .A(n4917), .B(n4918), .X(n4916) );
  nand_x1_sg U5804 ( .A(n4919), .B(n4920), .X(n4918) );
  nor_x1_sg U5805 ( .A(n4899), .B(n4900), .X(n4898) );
  nand_x1_sg U5806 ( .A(n4903), .B(n4904), .X(n4899) );
  nor_x1_sg U5807 ( .A(n4907), .B(n4908), .X(n4897) );
  nand_x1_sg U5808 ( .A(n4909), .B(n4910), .X(n4908) );
  nor_x1_sg U5809 ( .A(n4886), .B(n4887), .X(n4876) );
  nand_x1_sg U5810 ( .A(n4890), .B(n4891), .X(n4886) );
  nor_x1_sg U5811 ( .A(n4878), .B(n4879), .X(n4877) );
  nand_x1_sg U5812 ( .A(n4880), .B(n4881), .X(n4879) );
  nor_x1_sg U5813 ( .A(n4860), .B(n4861), .X(n4859) );
  nand_x1_sg U5814 ( .A(n4864), .B(n4865), .X(n4860) );
  nor_x1_sg U5815 ( .A(n4868), .B(n4869), .X(n4858) );
  nand_x1_sg U5816 ( .A(n4870), .B(n4871), .X(n4869) );
  nor_x1_sg U5817 ( .A(n4847), .B(n4848), .X(n4837) );
  nand_x1_sg U5818 ( .A(n4851), .B(n4852), .X(n4847) );
  nor_x1_sg U5819 ( .A(n4839), .B(n4840), .X(n4838) );
  nand_x1_sg U5820 ( .A(n4841), .B(n4842), .X(n4840) );
  nor_x1_sg U5821 ( .A(n4821), .B(n4822), .X(n4820) );
  nand_x1_sg U5822 ( .A(n4825), .B(n4826), .X(n4821) );
  nor_x1_sg U5823 ( .A(n4829), .B(n4830), .X(n4819) );
  nand_x1_sg U5824 ( .A(n4831), .B(n4832), .X(n4830) );
  nor_x1_sg U5825 ( .A(n4808), .B(n4809), .X(n4798) );
  nand_x1_sg U5826 ( .A(n4812), .B(n4813), .X(n4808) );
  nor_x1_sg U5827 ( .A(n4800), .B(n4801), .X(n4799) );
  nand_x1_sg U5828 ( .A(n4802), .B(n4803), .X(n4801) );
  nor_x1_sg U5829 ( .A(n4782), .B(n4783), .X(n4781) );
  nand_x1_sg U5830 ( .A(n4786), .B(n4787), .X(n4782) );
  nor_x1_sg U5831 ( .A(n4790), .B(n4791), .X(n4780) );
  nand_x1_sg U5832 ( .A(n4792), .B(n4793), .X(n4791) );
  nor_x1_sg U5833 ( .A(n4769), .B(n4770), .X(n4759) );
  nand_x1_sg U5834 ( .A(n4773), .B(n4774), .X(n4769) );
  nor_x1_sg U5835 ( .A(n4761), .B(n4762), .X(n4760) );
  nand_x1_sg U5836 ( .A(n4763), .B(n4764), .X(n4762) );
  nor_x1_sg U5837 ( .A(n4743), .B(n4744), .X(n4742) );
  nand_x1_sg U5838 ( .A(n4747), .B(n4748), .X(n4743) );
  nor_x1_sg U5839 ( .A(n4751), .B(n4752), .X(n4741) );
  nand_x1_sg U5840 ( .A(n4753), .B(n4754), .X(n4752) );
  nor_x1_sg U5841 ( .A(n4730), .B(n4731), .X(n4720) );
  nand_x1_sg U5842 ( .A(n4734), .B(n4735), .X(n4730) );
  nor_x1_sg U5843 ( .A(n4722), .B(n4723), .X(n4721) );
  nand_x1_sg U5844 ( .A(n4724), .B(n4725), .X(n4723) );
  nor_x1_sg U5845 ( .A(n4704), .B(n4705), .X(n4703) );
  nand_x1_sg U5846 ( .A(n4708), .B(n4709), .X(n4704) );
  nor_x1_sg U5847 ( .A(n4712), .B(n4713), .X(n4702) );
  nand_x1_sg U5848 ( .A(n4714), .B(n4715), .X(n4713) );
  nor_x1_sg U5849 ( .A(n4691), .B(n4692), .X(n4681) );
  nand_x1_sg U5850 ( .A(n4695), .B(n4696), .X(n4691) );
  nor_x1_sg U5851 ( .A(n4683), .B(n4684), .X(n4682) );
  nand_x1_sg U5852 ( .A(n4685), .B(n4686), .X(n4684) );
  nor_x1_sg U5853 ( .A(n4665), .B(n4666), .X(n4664) );
  nand_x1_sg U5854 ( .A(n4669), .B(n4670), .X(n4665) );
  nor_x1_sg U5855 ( .A(n4673), .B(n4674), .X(n4663) );
  nand_x1_sg U5856 ( .A(n4675), .B(n4676), .X(n4674) );
  nor_x1_sg U5857 ( .A(n4652), .B(n4653), .X(n4642) );
  nand_x1_sg U5858 ( .A(n4656), .B(n4657), .X(n4652) );
  nor_x1_sg U5859 ( .A(n4644), .B(n4645), .X(n4643) );
  nand_x1_sg U5860 ( .A(n4646), .B(n4647), .X(n4645) );
  nor_x1_sg U5861 ( .A(n4626), .B(n4627), .X(n4625) );
  nand_x1_sg U5862 ( .A(n4630), .B(n4631), .X(n4626) );
  nor_x1_sg U5863 ( .A(n4634), .B(n4635), .X(n4624) );
  nand_x1_sg U5864 ( .A(n4636), .B(n4637), .X(n4635) );
  nor_x1_sg U5865 ( .A(n4613), .B(n4614), .X(n4603) );
  nand_x1_sg U5866 ( .A(n4617), .B(n4618), .X(n4613) );
  nor_x1_sg U5867 ( .A(n4605), .B(n4606), .X(n4604) );
  nand_x1_sg U5868 ( .A(n4607), .B(n4608), .X(n4606) );
  nor_x1_sg U5869 ( .A(n4587), .B(n4588), .X(n4586) );
  nand_x1_sg U5870 ( .A(n4591), .B(n4592), .X(n4587) );
  nor_x1_sg U5871 ( .A(n4595), .B(n4596), .X(n4585) );
  nand_x1_sg U5872 ( .A(n4597), .B(n4598), .X(n4596) );
  nor_x1_sg U5873 ( .A(n4574), .B(n4575), .X(n4564) );
  nand_x1_sg U5874 ( .A(n4578), .B(n4579), .X(n4574) );
  nor_x1_sg U5875 ( .A(n4566), .B(n4567), .X(n4565) );
  nand_x1_sg U5876 ( .A(n4568), .B(n4569), .X(n4567) );
  nor_x1_sg U5877 ( .A(n4548), .B(n4549), .X(n4547) );
  nand_x1_sg U5878 ( .A(n4552), .B(n4553), .X(n4548) );
  nor_x1_sg U5879 ( .A(n4556), .B(n4557), .X(n4546) );
  nand_x1_sg U5880 ( .A(n4558), .B(n4559), .X(n4557) );
  nor_x1_sg U5881 ( .A(n4535), .B(n4536), .X(n4525) );
  nand_x1_sg U5882 ( .A(n4539), .B(n4540), .X(n4535) );
  nor_x1_sg U5883 ( .A(n4527), .B(n4528), .X(n4526) );
  nand_x1_sg U5884 ( .A(n4529), .B(n4530), .X(n4528) );
  nor_x1_sg U5885 ( .A(n4509), .B(n4510), .X(n4508) );
  nand_x1_sg U5886 ( .A(n4513), .B(n4514), .X(n4509) );
  nor_x1_sg U5887 ( .A(n4517), .B(n4518), .X(n4507) );
  nand_x1_sg U5888 ( .A(n4519), .B(n4520), .X(n4518) );
  nor_x1_sg U5889 ( .A(n4496), .B(n4497), .X(n4486) );
  nand_x1_sg U5890 ( .A(n4500), .B(n4501), .X(n4496) );
  nor_x1_sg U5891 ( .A(n4488), .B(n4489), .X(n4487) );
  nand_x1_sg U5892 ( .A(n4490), .B(n4491), .X(n4489) );
  nor_x1_sg U5893 ( .A(n4470), .B(n4471), .X(n4469) );
  nand_x1_sg U5894 ( .A(n4474), .B(n4475), .X(n4470) );
  nor_x1_sg U5895 ( .A(n4478), .B(n4479), .X(n4468) );
  nand_x1_sg U5896 ( .A(n4480), .B(n4481), .X(n4479) );
  nor_x1_sg U5897 ( .A(n4453), .B(n4454), .X(n4438) );
  nand_x1_sg U5898 ( .A(n4458), .B(n4459), .X(n4453) );
  nor_x1_sg U5899 ( .A(n4440), .B(n4441), .X(n4439) );
  nand_x1_sg U5900 ( .A(n4442), .B(n4443), .X(n4441) );
  nor_x1_sg U5901 ( .A(n4413), .B(n4414), .X(n4412) );
  nand_x1_sg U5902 ( .A(n4419), .B(n4420), .X(n4413) );
  nor_x1_sg U5903 ( .A(n4426), .B(n4427), .X(n4411) );
  nand_x1_sg U5904 ( .A(n4428), .B(n4429), .X(n4427) );
  inv_x1_sg U5905 ( .A(n3487), .X(n3236) );
  nand_x2_sg U5906 ( .A(n3489), .B(n3490), .X(n3488) );
  nor_x1_sg U5907 ( .A(n3491), .B(n3492), .X(n3490) );
  nor_x1_sg U5908 ( .A(n3450), .B(n3451), .X(n3440) );
  inv_x1_sg U5909 ( .A(n3511), .X(n3288) );
  nand_x2_sg U5910 ( .A(n3440), .B(n3441), .X(n3439) );
  nand_x1_sg U5911 ( .A(n3235), .B(n3485), .X(n2368) );
  inv_x1_sg U5912 ( .A(n3486), .X(n3235) );
  nand_x1_sg U5913 ( .A(n4402), .B(n4403), .X(n1964) );
  nand_x1_sg U5914 ( .A(n3334), .B(n3498), .X(n3493) );
  nand_x1_sg U5915 ( .A(n3436), .B(n3437), .X(n2374) );
  inv_x1_sg U5916 ( .A(n3438), .X(n3263) );
  nand_x1_sg U5917 ( .A(n3861), .B(n3862), .X(n2213) );
  nand_x1_sg U5918 ( .A(n4031), .B(n4032), .X(n2133) );
  nand_x1_sg U5919 ( .A(n3690), .B(n3691), .X(n2293) );
  nand_x1_sg U5920 ( .A(n5246), .B(n5674), .X(n3690) );
  nand_x1_sg U5921 ( .A(n3832), .B(n3833), .X(n2227) );
  nand_x1_sg U5922 ( .A(n3835), .B(n3836), .X(n2226) );
  nand_x1_sg U5923 ( .A(n3837), .B(n3838), .X(n2225) );
  nand_x1_sg U5924 ( .A(n3839), .B(n3840), .X(n2224) );
  nand_x1_sg U5925 ( .A(n3841), .B(n3842), .X(n2223) );
  nand_x1_sg U5926 ( .A(n3843), .B(n3844), .X(n2222) );
  nand_x1_sg U5927 ( .A(n3845), .B(n3846), .X(n2221) );
  nand_x1_sg U5928 ( .A(n3847), .B(n3848), .X(n2220) );
  nand_x1_sg U5929 ( .A(n3849), .B(n3850), .X(n2219) );
  nand_x1_sg U5930 ( .A(n3851), .B(n3852), .X(n2218) );
  nand_x1_sg U5931 ( .A(n3853), .B(n3854), .X(n2217) );
  nand_x1_sg U5932 ( .A(n3855), .B(n3856), .X(n2216) );
  nand_x1_sg U5933 ( .A(n3857), .B(n3858), .X(n2215) );
  nand_x1_sg U5934 ( .A(n3859), .B(n3860), .X(n2214) );
  nand_x1_sg U5935 ( .A(n3863), .B(n3864), .X(n2212) );
  nand_x1_sg U5936 ( .A(n3865), .B(n3866), .X(n2211) );
  nand_x1_sg U5937 ( .A(n3867), .B(n3868), .X(n2210) );
  nand_x1_sg U5938 ( .A(n3869), .B(n3870), .X(n2209) );
  nand_x1_sg U5939 ( .A(n3871), .B(n3872), .X(n2208) );
  nand_x1_sg U5940 ( .A(n4175), .B(n4176), .X(n2066) );
  nand_x1_sg U5941 ( .A(n4179), .B(n4180), .X(n2064) );
  nand_x1_sg U5942 ( .A(n4183), .B(n4184), .X(n2062) );
  nand_x1_sg U5943 ( .A(n4187), .B(n4188), .X(n2060) );
  nand_x1_sg U5944 ( .A(n4191), .B(n4192), .X(n2058) );
  nand_x1_sg U5945 ( .A(n4195), .B(n4196), .X(n2056) );
  nand_x1_sg U5946 ( .A(n4199), .B(n4200), .X(n2054) );
  nand_x1_sg U5947 ( .A(n4203), .B(n4204), .X(n2052) );
  nand_x1_sg U5948 ( .A(n4207), .B(n4208), .X(n2050) );
  nand_x1_sg U5949 ( .A(n4033), .B(n4034), .X(n2132) );
  nand_x1_sg U5950 ( .A(n3692), .B(n3693), .X(n2292) );
  nand_x1_sg U5951 ( .A(n4035), .B(n4036), .X(n2131) );
  nand_x1_sg U5952 ( .A(n3694), .B(n3695), .X(n2291) );
  nand_x1_sg U5953 ( .A(n4037), .B(n4038), .X(n2130) );
  nand_x1_sg U5954 ( .A(n3696), .B(n3697), .X(n2290) );
  nand_x1_sg U5955 ( .A(n4039), .B(n4040), .X(n2129) );
  nand_x1_sg U5956 ( .A(n3698), .B(n3699), .X(n2289) );
  nand_x1_sg U5957 ( .A(n4041), .B(n4042), .X(n2128) );
  nand_x1_sg U5958 ( .A(n3700), .B(n3701), .X(n2288) );
  nand_x1_sg U5959 ( .A(n4002), .B(n4003), .X(n2147) );
  nand_x1_sg U5960 ( .A(n3661), .B(n3662), .X(n2307) );
  nand_x1_sg U5961 ( .A(n4005), .B(n4006), .X(n2146) );
  nand_x1_sg U5962 ( .A(n3664), .B(n3665), .X(n2306) );
  nand_x1_sg U5963 ( .A(n4007), .B(n4008), .X(n2145) );
  nand_x1_sg U5964 ( .A(n3666), .B(n3667), .X(n2305) );
  nand_x1_sg U5965 ( .A(n4009), .B(n4010), .X(n2144) );
  nand_x1_sg U5966 ( .A(n3668), .B(n3669), .X(n2304) );
  nand_x1_sg U5967 ( .A(n4011), .B(n4012), .X(n2143) );
  nand_x1_sg U5968 ( .A(n3670), .B(n3671), .X(n2303) );
  nand_x1_sg U5969 ( .A(n4013), .B(n4014), .X(n2142) );
  nand_x1_sg U5970 ( .A(n3672), .B(n3673), .X(n2302) );
  nand_x1_sg U5971 ( .A(n4015), .B(n4016), .X(n2141) );
  nand_x1_sg U5972 ( .A(n3674), .B(n3675), .X(n2301) );
  nand_x1_sg U5973 ( .A(n4017), .B(n4018), .X(n2140) );
  nand_x1_sg U5974 ( .A(n3676), .B(n3677), .X(n2300) );
  nand_x1_sg U5975 ( .A(n4019), .B(n4020), .X(n2139) );
  nand_x1_sg U5976 ( .A(n3678), .B(n3679), .X(n2299) );
  nand_x1_sg U5977 ( .A(n4021), .B(n4022), .X(n2138) );
  nand_x1_sg U5978 ( .A(n3680), .B(n3681), .X(n2298) );
  nand_x1_sg U5979 ( .A(n4023), .B(n4024), .X(n2137) );
  nand_x1_sg U5980 ( .A(n3682), .B(n3683), .X(n2297) );
  nand_x1_sg U5981 ( .A(n4025), .B(n4026), .X(n2136) );
  nand_x1_sg U5982 ( .A(n3684), .B(n3685), .X(n2296) );
  nand_x1_sg U5983 ( .A(n4027), .B(n4028), .X(n2135) );
  nand_x1_sg U5984 ( .A(n3686), .B(n3687), .X(n2295) );
  nand_x1_sg U5985 ( .A(n4029), .B(n4030), .X(n2134) );
  nand_x1_sg U5986 ( .A(n3688), .B(n3689), .X(n2294) );
  nand_x1_sg U5987 ( .A(n3739), .B(n3740), .X(n2271) );
  nand_x1_sg U5988 ( .A(n3743), .B(n3744), .X(n2269) );
  nand_x1_sg U5989 ( .A(n3745), .B(n3746), .X(n2268) );
  nand_x1_sg U5990 ( .A(n3706), .B(n3707), .X(n2287) );
  nand_x1_sg U5991 ( .A(n3711), .B(n3712), .X(n2285) );
  nand_x1_sg U5992 ( .A(n3715), .B(n3716), .X(n2283) );
  nand_x1_sg U5993 ( .A(n3719), .B(n3720), .X(n2281) );
  nand_x1_sg U5994 ( .A(n3723), .B(n3724), .X(n2279) );
  nand_x1_sg U5995 ( .A(n3727), .B(n3728), .X(n2277) );
  nand_x1_sg U5996 ( .A(n3731), .B(n3732), .X(n2275) );
  nand_x1_sg U5997 ( .A(n4088), .B(n4089), .X(n2107) );
  nand_x1_sg U5998 ( .A(n4093), .B(n4094), .X(n2105) );
  nand_x1_sg U5999 ( .A(n4097), .B(n4098), .X(n2103) );
  nand_x1_sg U6000 ( .A(n4101), .B(n4102), .X(n2101) );
  nand_x1_sg U6001 ( .A(n4105), .B(n4106), .X(n2099) );
  nand_x1_sg U6002 ( .A(n4109), .B(n4110), .X(n2097) );
  nand_x1_sg U6003 ( .A(n4113), .B(n4114), .X(n2095) );
  nand_x1_sg U6004 ( .A(n4121), .B(n4122), .X(n2091) );
  nand_x1_sg U6005 ( .A(n4125), .B(n4126), .X(n2089) );
  nand_x1_sg U6006 ( .A(n4127), .B(n4128), .X(n2088) );
  nand_x1_sg U6007 ( .A(n3993), .B(n3994), .X(n2151) );
  nand_x1_sg U6008 ( .A(n3997), .B(n3998), .X(n2149) );
  nand_x1_sg U6009 ( .A(n3999), .B(n4000), .X(n2148) );
  nand_x1_sg U6010 ( .A(n3960), .B(n3961), .X(n2167) );
  nand_x1_sg U6011 ( .A(n3965), .B(n3966), .X(n2165) );
  nand_x1_sg U6012 ( .A(n3969), .B(n3970), .X(n2163) );
  nand_x1_sg U6013 ( .A(n3973), .B(n3974), .X(n2161) );
  nand_x1_sg U6014 ( .A(n3977), .B(n3978), .X(n2159) );
  nand_x1_sg U6015 ( .A(n3981), .B(n3982), .X(n2157) );
  nand_x1_sg U6016 ( .A(n3985), .B(n3986), .X(n2155) );
  nand_x1_sg U6017 ( .A(n3748), .B(n3749), .X(n2267) );
  nand_x1_sg U6018 ( .A(n3753), .B(n3754), .X(n2265) );
  nand_x1_sg U6019 ( .A(n3757), .B(n3758), .X(n2263) );
  nand_x1_sg U6020 ( .A(n3761), .B(n3762), .X(n2261) );
  nand_x1_sg U6021 ( .A(n3765), .B(n3766), .X(n2259) );
  nand_x1_sg U6022 ( .A(n3769), .B(n3770), .X(n2257) );
  nand_x1_sg U6023 ( .A(n3773), .B(n3774), .X(n2255) );
  nand_x1_sg U6024 ( .A(n3781), .B(n3782), .X(n2251) );
  nand_x1_sg U6025 ( .A(n3785), .B(n3786), .X(n2249) );
  nand_x1_sg U6026 ( .A(n3787), .B(n3788), .X(n2248) );
  nand_x1_sg U6027 ( .A(n4046), .B(n4047), .X(n2127) );
  nand_x1_sg U6028 ( .A(n4051), .B(n4052), .X(n2125) );
  nand_x1_sg U6029 ( .A(n4055), .B(n4056), .X(n2123) );
  nand_x1_sg U6030 ( .A(n4059), .B(n4060), .X(n2121) );
  nand_x1_sg U6031 ( .A(n4063), .B(n4064), .X(n2119) );
  nand_x1_sg U6032 ( .A(n4067), .B(n4068), .X(n2117) );
  nand_x1_sg U6033 ( .A(n4071), .B(n4072), .X(n2115) );
  nand_x1_sg U6034 ( .A(n4079), .B(n4080), .X(n2111) );
  nand_x1_sg U6035 ( .A(n4083), .B(n4084), .X(n2109) );
  nand_x1_sg U6036 ( .A(n4085), .B(n4086), .X(n2108) );
  nand_x1_sg U6037 ( .A(n3737), .B(n3738), .X(n2272) );
  nand_x1_sg U6038 ( .A(n3741), .B(n3742), .X(n2270) );
  nand_x1_sg U6039 ( .A(n3709), .B(n3710), .X(n2286) );
  nand_x1_sg U6040 ( .A(n3713), .B(n3714), .X(n2284) );
  nand_x1_sg U6041 ( .A(n3717), .B(n3718), .X(n2282) );
  nand_x1_sg U6042 ( .A(n3721), .B(n3722), .X(n2280) );
  nand_x1_sg U6043 ( .A(n3725), .B(n3726), .X(n2278) );
  nand_x1_sg U6044 ( .A(n3729), .B(n3730), .X(n2276) );
  nand_x1_sg U6045 ( .A(n3733), .B(n3734), .X(n2274) );
  nand_x1_sg U6046 ( .A(n3751), .B(n3752), .X(n2266) );
  nand_x1_sg U6047 ( .A(n3755), .B(n3756), .X(n2264) );
  nand_x1_sg U6048 ( .A(n3759), .B(n3760), .X(n2262) );
  nand_x1_sg U6049 ( .A(n3763), .B(n3764), .X(n2260) );
  nand_x1_sg U6050 ( .A(n3767), .B(n3768), .X(n2258) );
  nand_x1_sg U6051 ( .A(n3771), .B(n3772), .X(n2256) );
  nand_x1_sg U6052 ( .A(n3775), .B(n3776), .X(n2254) );
  nand_x1_sg U6053 ( .A(n3779), .B(n3780), .X(n2252) );
  nand_x1_sg U6054 ( .A(n3783), .B(n3784), .X(n2250) );
  nand_x1_sg U6055 ( .A(n3793), .B(n3794), .X(n2246) );
  nand_x1_sg U6056 ( .A(n3797), .B(n3798), .X(n2244) );
  nand_x1_sg U6057 ( .A(n3801), .B(n3802), .X(n2242) );
  nand_x1_sg U6058 ( .A(n3805), .B(n3806), .X(n2240) );
  nand_x1_sg U6059 ( .A(n3809), .B(n3810), .X(n2238) );
  nand_x1_sg U6060 ( .A(n3813), .B(n3814), .X(n2236) );
  nand_x1_sg U6061 ( .A(n3817), .B(n3818), .X(n2234) );
  nand_x1_sg U6062 ( .A(n3821), .B(n3822), .X(n2232) );
  nand_x1_sg U6063 ( .A(n3825), .B(n3826), .X(n2230) );
  nand_x1_sg U6064 ( .A(n4049), .B(n4050), .X(n2126) );
  nand_x1_sg U6065 ( .A(n4053), .B(n4054), .X(n2124) );
  nand_x1_sg U6066 ( .A(n4057), .B(n4058), .X(n2122) );
  nand_x1_sg U6067 ( .A(n4061), .B(n4062), .X(n2120) );
  nand_x1_sg U6068 ( .A(n4065), .B(n4066), .X(n2118) );
  nand_x1_sg U6069 ( .A(n4069), .B(n4070), .X(n2116) );
  nand_x1_sg U6070 ( .A(n4073), .B(n4074), .X(n2114) );
  nand_x1_sg U6071 ( .A(n4077), .B(n4078), .X(n2112) );
  nand_x1_sg U6072 ( .A(n4081), .B(n4082), .X(n2110) );
  nand_x1_sg U6073 ( .A(n4091), .B(n4092), .X(n2106) );
  nand_x1_sg U6074 ( .A(n4095), .B(n4096), .X(n2104) );
  nand_x1_sg U6075 ( .A(n4099), .B(n4100), .X(n2102) );
  nand_x1_sg U6076 ( .A(n4103), .B(n4104), .X(n2100) );
  nand_x1_sg U6077 ( .A(n4107), .B(n4108), .X(n2098) );
  nand_x1_sg U6078 ( .A(n4111), .B(n4112), .X(n2096) );
  nand_x1_sg U6079 ( .A(n4115), .B(n4116), .X(n2094) );
  nand_x1_sg U6080 ( .A(n4119), .B(n4120), .X(n2092) );
  nand_x1_sg U6081 ( .A(n4123), .B(n4124), .X(n2090) );
  nand_x1_sg U6082 ( .A(n4133), .B(n4134), .X(n2086) );
  nand_x1_sg U6083 ( .A(n4137), .B(n4138), .X(n2084) );
  nand_x1_sg U6084 ( .A(n4141), .B(n4142), .X(n2082) );
  nand_x1_sg U6085 ( .A(n4145), .B(n4146), .X(n2080) );
  nand_x1_sg U6086 ( .A(n4149), .B(n4150), .X(n2078) );
  nand_x1_sg U6087 ( .A(n4153), .B(n4154), .X(n2076) );
  nand_x1_sg U6088 ( .A(n4157), .B(n4158), .X(n2074) );
  nand_x1_sg U6089 ( .A(n4161), .B(n4162), .X(n2072) );
  nand_x1_sg U6090 ( .A(n4165), .B(n4166), .X(n2070) );
  nand_x1_sg U6091 ( .A(n3907), .B(n3908), .X(n2192) );
  nand_x1_sg U6092 ( .A(n3949), .B(n3950), .X(n2172) );
  nand_x1_sg U6093 ( .A(n3991), .B(n3992), .X(n2152) );
  nand_x1_sg U6094 ( .A(n3911), .B(n3912), .X(n2190) );
  nand_x1_sg U6095 ( .A(n3953), .B(n3954), .X(n2170) );
  nand_x1_sg U6096 ( .A(n3995), .B(n3996), .X(n2150) );
  nand_x1_sg U6097 ( .A(n3879), .B(n3880), .X(n2206) );
  nand_x1_sg U6098 ( .A(n3921), .B(n3922), .X(n2186) );
  nand_x1_sg U6099 ( .A(n3963), .B(n3964), .X(n2166) );
  nand_x1_sg U6100 ( .A(n3883), .B(n3884), .X(n2204) );
  nand_x1_sg U6101 ( .A(n3925), .B(n3926), .X(n2184) );
  nand_x1_sg U6102 ( .A(n3967), .B(n3968), .X(n2164) );
  nand_x1_sg U6103 ( .A(n3887), .B(n3888), .X(n2202) );
  nand_x1_sg U6104 ( .A(n3929), .B(n3930), .X(n2182) );
  nand_x1_sg U6105 ( .A(n3971), .B(n3972), .X(n2162) );
  nand_x1_sg U6106 ( .A(n3891), .B(n3892), .X(n2200) );
  nand_x1_sg U6107 ( .A(n3933), .B(n3934), .X(n2180) );
  nand_x1_sg U6108 ( .A(n3975), .B(n3976), .X(n2160) );
  nand_x1_sg U6109 ( .A(n3895), .B(n3896), .X(n2198) );
  nand_x1_sg U6110 ( .A(n3937), .B(n3938), .X(n2178) );
  nand_x1_sg U6111 ( .A(n3979), .B(n3980), .X(n2158) );
  nand_x1_sg U6112 ( .A(n3899), .B(n3900), .X(n2196) );
  nand_x1_sg U6113 ( .A(n3941), .B(n3942), .X(n2176) );
  nand_x1_sg U6114 ( .A(n3983), .B(n3984), .X(n2156) );
  nand_x1_sg U6115 ( .A(n3903), .B(n3904), .X(n2194) );
  nand_x1_sg U6116 ( .A(n3945), .B(n3946), .X(n2174) );
  nand_x1_sg U6117 ( .A(n3987), .B(n3988), .X(n2154) );
  nand_x1_sg U6118 ( .A(n3819), .B(n3820), .X(n2233) );
  nand_x1_sg U6119 ( .A(n3905), .B(n3906), .X(n2193) );
  nand_x1_sg U6120 ( .A(n3947), .B(n3948), .X(n2173) );
  nand_x1_sg U6121 ( .A(n4159), .B(n4160), .X(n2073) );
  nand_x1_sg U6122 ( .A(n4201), .B(n4202), .X(n2053) );
  nand_x1_sg U6123 ( .A(n3790), .B(n3791), .X(n2247) );
  nand_x1_sg U6124 ( .A(n3795), .B(n3796), .X(n2245) );
  nand_x1_sg U6125 ( .A(n3799), .B(n3800), .X(n2243) );
  nand_x1_sg U6126 ( .A(n3803), .B(n3804), .X(n2241) );
  nand_x1_sg U6127 ( .A(n3807), .B(n3808), .X(n2239) );
  nand_x1_sg U6128 ( .A(n3811), .B(n3812), .X(n2237) );
  nand_x1_sg U6129 ( .A(n3815), .B(n3816), .X(n2235) );
  nand_x1_sg U6130 ( .A(n3823), .B(n3824), .X(n2231) );
  nand_x1_sg U6131 ( .A(n3827), .B(n3828), .X(n2229) );
  nand_x1_sg U6132 ( .A(n3829), .B(n3830), .X(n2228) );
  nand_x1_sg U6133 ( .A(n4130), .B(n4131), .X(n2087) );
  nand_x1_sg U6134 ( .A(n4135), .B(n4136), .X(n2085) );
  nand_x1_sg U6135 ( .A(n4139), .B(n4140), .X(n2083) );
  nand_x1_sg U6136 ( .A(n4143), .B(n4144), .X(n2081) );
  nand_x1_sg U6137 ( .A(n4147), .B(n4148), .X(n2079) );
  nand_x1_sg U6138 ( .A(n4151), .B(n4152), .X(n2077) );
  nand_x1_sg U6139 ( .A(n4155), .B(n4156), .X(n2075) );
  nand_x1_sg U6140 ( .A(n4163), .B(n4164), .X(n2071) );
  nand_x1_sg U6141 ( .A(n4167), .B(n4168), .X(n2069) );
  nand_x1_sg U6142 ( .A(n4169), .B(n4170), .X(n2068) );
  nand_x1_sg U6143 ( .A(n4172), .B(n4173), .X(n2067) );
  nand_x1_sg U6144 ( .A(n4177), .B(n4178), .X(n2065) );
  nand_x1_sg U6145 ( .A(n4181), .B(n4182), .X(n2063) );
  nand_x1_sg U6146 ( .A(n4185), .B(n4186), .X(n2061) );
  nand_x1_sg U6147 ( .A(n4189), .B(n4190), .X(n2059) );
  nand_x1_sg U6148 ( .A(n4193), .B(n4194), .X(n2057) );
  nand_x1_sg U6149 ( .A(n4197), .B(n4198), .X(n2055) );
  nand_x1_sg U6150 ( .A(n4205), .B(n4206), .X(n2051) );
  nand_x1_sg U6151 ( .A(n4209), .B(n4210), .X(n2049) );
  nand_x1_sg U6152 ( .A(n4211), .B(n4212), .X(n2048) );
  nand_x1_sg U6153 ( .A(n3909), .B(n3910), .X(n2191) );
  nand_x1_sg U6154 ( .A(n3951), .B(n3952), .X(n2171) );
  nand_x1_sg U6155 ( .A(n3913), .B(n3914), .X(n2189) );
  nand_x1_sg U6156 ( .A(n3955), .B(n3956), .X(n2169) );
  nand_x1_sg U6157 ( .A(n3915), .B(n3916), .X(n2188) );
  nand_x1_sg U6158 ( .A(n3957), .B(n3958), .X(n2168) );
  nand_x1_sg U6159 ( .A(n3876), .B(n3877), .X(n2207) );
  nand_x1_sg U6160 ( .A(n3918), .B(n3919), .X(n2187) );
  nand_x1_sg U6161 ( .A(n3881), .B(n3882), .X(n2205) );
  nand_x1_sg U6162 ( .A(n3923), .B(n3924), .X(n2185) );
  nand_x1_sg U6163 ( .A(n3885), .B(n3886), .X(n2203) );
  nand_x1_sg U6164 ( .A(n3927), .B(n3928), .X(n2183) );
  nand_x1_sg U6165 ( .A(n3889), .B(n3890), .X(n2201) );
  nand_x1_sg U6166 ( .A(n3931), .B(n3932), .X(n2181) );
  nand_x1_sg U6167 ( .A(n3893), .B(n3894), .X(n2199) );
  nand_x1_sg U6168 ( .A(n3935), .B(n3936), .X(n2179) );
  nand_x1_sg U6169 ( .A(n3897), .B(n3898), .X(n2197) );
  nand_x1_sg U6170 ( .A(n3939), .B(n3940), .X(n2177) );
  nand_x1_sg U6171 ( .A(n3901), .B(n3902), .X(n2195) );
  nand_x1_sg U6172 ( .A(n3943), .B(n3944), .X(n2175) );
  nand_x1_sg U6173 ( .A(n3777), .B(n3778), .X(n2253) );
  nand_x1_sg U6174 ( .A(n5246), .B(n5331), .X(n3777) );
  nand_x1_sg U6175 ( .A(n4075), .B(n4076), .X(n2113) );
  nand_x1_sg U6176 ( .A(n5409), .B(n5777), .X(n4075) );
  nand_x1_sg U6177 ( .A(n3735), .B(n3736), .X(n2273) );
  nand_x1_sg U6178 ( .A(n5410), .B(n5801), .X(n3735) );
  nand_x1_sg U6179 ( .A(n3989), .B(n3990), .X(n2153) );
  nand_x1_sg U6180 ( .A(n5408), .B(n5785), .X(n3989) );
  nand_x1_sg U6181 ( .A(n4117), .B(n4118), .X(n2093) );
  nand_x1_sg U6182 ( .A(n5408), .B(n5654), .X(n4117) );
  nand_x1_sg U6183 ( .A(n3560), .B(n3561), .X(n2352) );
  nand_x1_sg U6184 ( .A(n3608), .B(n3609), .X(n2332) );
  nand_x1_sg U6185 ( .A(n3650), .B(n3651), .X(n2312) );
  nand_x1_sg U6186 ( .A(n3566), .B(n3567), .X(n2350) );
  nand_x1_sg U6187 ( .A(n3612), .B(n3613), .X(n2330) );
  nand_x1_sg U6188 ( .A(n3654), .B(n3655), .X(n2310) );
  nand_x1_sg U6189 ( .A(n3518), .B(n3519), .X(n2366) );
  nand_x1_sg U6190 ( .A(n3580), .B(n3581), .X(n2346) );
  nand_x1_sg U6191 ( .A(n3622), .B(n3623), .X(n2326) );
  nand_x1_sg U6192 ( .A(n3524), .B(n3525), .X(n2364) );
  nand_x1_sg U6193 ( .A(n3584), .B(n3585), .X(n2344) );
  nand_x1_sg U6194 ( .A(n3626), .B(n3627), .X(n2324) );
  nand_x1_sg U6195 ( .A(n3530), .B(n3531), .X(n2362) );
  nand_x1_sg U6196 ( .A(n3588), .B(n3589), .X(n2342) );
  nand_x1_sg U6197 ( .A(n3630), .B(n3631), .X(n2322) );
  nand_x1_sg U6198 ( .A(n3536), .B(n3537), .X(n2360) );
  nand_x1_sg U6199 ( .A(n3592), .B(n3593), .X(n2340) );
  nand_x1_sg U6200 ( .A(n3634), .B(n3635), .X(n2320) );
  nand_x1_sg U6201 ( .A(n3542), .B(n3543), .X(n2358) );
  nand_x1_sg U6202 ( .A(n3596), .B(n3597), .X(n2338) );
  nand_x1_sg U6203 ( .A(n3638), .B(n3639), .X(n2318) );
  nand_x1_sg U6204 ( .A(n3548), .B(n3549), .X(n2356) );
  nand_x1_sg U6205 ( .A(n3600), .B(n3601), .X(n2336) );
  nand_x1_sg U6206 ( .A(n3642), .B(n3643), .X(n2316) );
  nand_x1_sg U6207 ( .A(n3554), .B(n3555), .X(n2354) );
  nand_x1_sg U6208 ( .A(n3604), .B(n3605), .X(n2334) );
  nand_x1_sg U6209 ( .A(n3646), .B(n3647), .X(n2314) );
  nand_x1_sg U6210 ( .A(n3557), .B(n3558), .X(n2353) );
  nand_x1_sg U6211 ( .A(n3606), .B(n3607), .X(n2333) );
  nand_x1_sg U6212 ( .A(n3648), .B(n3649), .X(n2313) );
  nand_x1_sg U6213 ( .A(n3563), .B(n3564), .X(n2351) );
  nand_x1_sg U6214 ( .A(n3610), .B(n3611), .X(n2331) );
  nand_x1_sg U6215 ( .A(n3652), .B(n3653), .X(n2311) );
  nand_x1_sg U6216 ( .A(n3569), .B(n3570), .X(n2349) );
  nand_x1_sg U6217 ( .A(n3614), .B(n3615), .X(n2329) );
  nand_x1_sg U6218 ( .A(n3656), .B(n3657), .X(n2309) );
  nand_x1_sg U6219 ( .A(n3572), .B(n3573), .X(n2348) );
  nand_x1_sg U6220 ( .A(n3616), .B(n3617), .X(n2328) );
  nand_x1_sg U6221 ( .A(n3658), .B(n3659), .X(n2308) );
  nand_x1_sg U6222 ( .A(n3514), .B(n3515), .X(n2367) );
  nand_x1_sg U6223 ( .A(n3577), .B(n3578), .X(n2347) );
  nand_x1_sg U6224 ( .A(n3619), .B(n3620), .X(n2327) );
  nand_x1_sg U6225 ( .A(n3521), .B(n3522), .X(n2365) );
  nand_x1_sg U6226 ( .A(n3582), .B(n3583), .X(n2345) );
  nand_x1_sg U6227 ( .A(n3624), .B(n3625), .X(n2325) );
  nand_x1_sg U6228 ( .A(n3527), .B(n3528), .X(n2363) );
  nand_x1_sg U6229 ( .A(n3586), .B(n3587), .X(n2343) );
  nand_x1_sg U6230 ( .A(n3628), .B(n3629), .X(n2323) );
  nand_x1_sg U6231 ( .A(n3533), .B(n3534), .X(n2361) );
  nand_x1_sg U6232 ( .A(n3590), .B(n3591), .X(n2341) );
  nand_x1_sg U6233 ( .A(n3632), .B(n3633), .X(n2321) );
  nand_x1_sg U6234 ( .A(n3539), .B(n3540), .X(n2359) );
  nand_x1_sg U6235 ( .A(n3594), .B(n3595), .X(n2339) );
  nand_x1_sg U6236 ( .A(n3636), .B(n3637), .X(n2319) );
  nand_x1_sg U6237 ( .A(n3545), .B(n3546), .X(n2357) );
  nand_x1_sg U6238 ( .A(n3598), .B(n3599), .X(n2337) );
  nand_x1_sg U6239 ( .A(n3640), .B(n3641), .X(n2317) );
  nand_x1_sg U6240 ( .A(n3551), .B(n3552), .X(n2355) );
  nand_x1_sg U6241 ( .A(n3602), .B(n3603), .X(n2335) );
  nand_x1_sg U6242 ( .A(n3644), .B(n3645), .X(n2315) );
  nand_x1_sg U6243 ( .A(n4371), .B(n4372), .X(n1973) );
  nand_x1_sg U6244 ( .A(n4373), .B(n4374), .X(n1972) );
  nand_x1_sg U6245 ( .A(n4375), .B(n4376), .X(n1971) );
  nand_x1_sg U6246 ( .A(n4377), .B(n4378), .X(n1970) );
  nand_x1_sg U6247 ( .A(n4379), .B(n4380), .X(n1969) );
  nand_x1_sg U6248 ( .A(n4342), .B(n4343), .X(n1987) );
  nand_x1_sg U6249 ( .A(n4345), .B(n4346), .X(n1986) );
  nand_x1_sg U6250 ( .A(n4347), .B(n4348), .X(n1985) );
  nand_x1_sg U6251 ( .A(n4349), .B(n4350), .X(n1984) );
  nand_x1_sg U6252 ( .A(n4351), .B(n4352), .X(n1983) );
  nand_x1_sg U6253 ( .A(n4353), .B(n4354), .X(n1982) );
  nand_x1_sg U6254 ( .A(n4355), .B(n4356), .X(n1981) );
  nand_x1_sg U6255 ( .A(n4357), .B(n4358), .X(n1980) );
  nand_x1_sg U6256 ( .A(n4359), .B(n4360), .X(n1979) );
  nand_x1_sg U6257 ( .A(n4361), .B(n4362), .X(n1978) );
  nand_x1_sg U6258 ( .A(n4363), .B(n4364), .X(n1977) );
  nand_x1_sg U6259 ( .A(n4365), .B(n4366), .X(n1976) );
  nand_x1_sg U6260 ( .A(n4367), .B(n4368), .X(n1975) );
  nand_x1_sg U6261 ( .A(n4369), .B(n4370), .X(n1974) );
  nand_x1_sg U6262 ( .A(n4381), .B(n4382), .X(n1968) );
  nand_x1_sg U6263 ( .A(n4247), .B(n4248), .X(n2032) );
  nand_x1_sg U6264 ( .A(n4289), .B(n4290), .X(n2012) );
  nand_x1_sg U6265 ( .A(n4331), .B(n4332), .X(n1992) );
  nand_x1_sg U6266 ( .A(n4251), .B(n4252), .X(n2030) );
  nand_x1_sg U6267 ( .A(n4293), .B(n4294), .X(n2010) );
  nand_x1_sg U6268 ( .A(n4335), .B(n4336), .X(n1990) );
  nand_x1_sg U6269 ( .A(n4219), .B(n4220), .X(n2046) );
  nand_x1_sg U6270 ( .A(n4261), .B(n4262), .X(n2026) );
  nand_x1_sg U6271 ( .A(n4303), .B(n4304), .X(n2006) );
  nand_x1_sg U6272 ( .A(n4223), .B(n4224), .X(n2044) );
  nand_x1_sg U6273 ( .A(n4265), .B(n4266), .X(n2024) );
  nand_x1_sg U6274 ( .A(n4307), .B(n4308), .X(n2004) );
  nand_x1_sg U6275 ( .A(n4227), .B(n4228), .X(n2042) );
  nand_x1_sg U6276 ( .A(n4269), .B(n4270), .X(n2022) );
  nand_x1_sg U6277 ( .A(n4311), .B(n4312), .X(n2002) );
  nand_x1_sg U6278 ( .A(n4231), .B(n4232), .X(n2040) );
  nand_x1_sg U6279 ( .A(n4273), .B(n4274), .X(n2020) );
  nand_x1_sg U6280 ( .A(n4315), .B(n4316), .X(n2000) );
  nand_x1_sg U6281 ( .A(n4235), .B(n4236), .X(n2038) );
  nand_x1_sg U6282 ( .A(n4277), .B(n4278), .X(n2018) );
  nand_x1_sg U6283 ( .A(n4319), .B(n4320), .X(n1998) );
  nand_x1_sg U6284 ( .A(n4239), .B(n4240), .X(n2036) );
  nand_x1_sg U6285 ( .A(n4281), .B(n4282), .X(n2016) );
  nand_x1_sg U6286 ( .A(n4323), .B(n4324), .X(n1996) );
  nand_x1_sg U6287 ( .A(n4243), .B(n4244), .X(n2034) );
  nand_x1_sg U6288 ( .A(n4285), .B(n4286), .X(n2014) );
  nand_x1_sg U6289 ( .A(n4327), .B(n4328), .X(n1994) );
  nand_x1_sg U6290 ( .A(n4245), .B(n4246), .X(n2033) );
  nand_x1_sg U6291 ( .A(n4287), .B(n4288), .X(n2013) );
  nand_x1_sg U6292 ( .A(n4329), .B(n4330), .X(n1993) );
  nand_x1_sg U6293 ( .A(n4249), .B(n4250), .X(n2031) );
  nand_x1_sg U6294 ( .A(n4291), .B(n4292), .X(n2011) );
  nand_x1_sg U6295 ( .A(n4333), .B(n4334), .X(n1991) );
  nand_x1_sg U6296 ( .A(n4253), .B(n4254), .X(n2029) );
  nand_x1_sg U6297 ( .A(n4295), .B(n4296), .X(n2009) );
  nand_x1_sg U6298 ( .A(n4337), .B(n4338), .X(n1989) );
  nand_x1_sg U6299 ( .A(n4255), .B(n4256), .X(n2028) );
  nand_x1_sg U6300 ( .A(n4297), .B(n4298), .X(n2008) );
  nand_x1_sg U6301 ( .A(n4339), .B(n4340), .X(n1988) );
  nand_x1_sg U6302 ( .A(n4216), .B(n4217), .X(n2047) );
  nand_x1_sg U6303 ( .A(n4258), .B(n4259), .X(n2027) );
  nand_x1_sg U6304 ( .A(n4300), .B(n4301), .X(n2007) );
  nand_x1_sg U6305 ( .A(n4221), .B(n4222), .X(n2045) );
  nand_x1_sg U6306 ( .A(n4263), .B(n4264), .X(n2025) );
  nand_x1_sg U6307 ( .A(n4305), .B(n4306), .X(n2005) );
  nand_x1_sg U6308 ( .A(n4225), .B(n4226), .X(n2043) );
  nand_x1_sg U6309 ( .A(n4267), .B(n4268), .X(n2023) );
  nand_x1_sg U6310 ( .A(n4309), .B(n4310), .X(n2003) );
  nand_x1_sg U6311 ( .A(n4229), .B(n4230), .X(n2041) );
  nand_x1_sg U6312 ( .A(n4271), .B(n4272), .X(n2021) );
  nand_x1_sg U6313 ( .A(n4313), .B(n4314), .X(n2001) );
  nand_x1_sg U6314 ( .A(n4233), .B(n4234), .X(n2039) );
  nand_x1_sg U6315 ( .A(n4275), .B(n4276), .X(n2019) );
  nand_x1_sg U6316 ( .A(n4317), .B(n4318), .X(n1999) );
  nand_x1_sg U6317 ( .A(n4237), .B(n4238), .X(n2037) );
  nand_x1_sg U6318 ( .A(n4279), .B(n4280), .X(n2017) );
  nand_x1_sg U6319 ( .A(n4321), .B(n4322), .X(n1997) );
  nand_x1_sg U6320 ( .A(n4241), .B(n4242), .X(n2035) );
  nand_x1_sg U6321 ( .A(n4283), .B(n4284), .X(n2015) );
  nand_x1_sg U6322 ( .A(n4325), .B(n4326), .X(n1995) );
  nand_x1_sg U6323 ( .A(n4397), .B(n4398), .X(n1965) );
  nand_x1_sg U6324 ( .A(n3480), .B(n3481), .X(n2369) );
  nand_x1_sg U6325 ( .A(n4392), .B(n4393), .X(n1966) );
  nand_x1_sg U6326 ( .A(n4389), .B(n4390), .X(n1967) );
  nand_x1_sg U6327 ( .A(n3445), .B(n3446), .X(n3444) );
  nand_x1_sg U6328 ( .A(n3475), .B(n3476), .X(n2370) );
  nand_x1_sg U6329 ( .A(n3470), .B(n3471), .X(n2371) );
  nand_x1_sg U6330 ( .A(n3433), .B(n3434), .X(n2375) );
  nand_x1_sg U6331 ( .A(n3466), .B(n3467), .X(n2372) );
  nand_x1_sg U6332 ( .A(n3463), .B(n3464), .X(n2373) );
  nand_x1_sg U6333 ( .A(n5208), .B(n5209), .X(n5207) );
  nand_x1_sg U6334 ( .A(n5161), .B(n5162), .X(n5160) );
  nand_x1_sg U6335 ( .A(n5083), .B(n5084), .X(n5082) );
  nand_x1_sg U6336 ( .A(n5044), .B(n5045), .X(n5043) );
  nand_x1_sg U6337 ( .A(n4966), .B(n4967), .X(n4965) );
  nand_x1_sg U6338 ( .A(n4927), .B(n4928), .X(n4926) );
  nand_x1_sg U6339 ( .A(n4849), .B(n4850), .X(n4848) );
  nand_x1_sg U6340 ( .A(n4810), .B(n4811), .X(n4809) );
  nand_x1_sg U6341 ( .A(n4732), .B(n4733), .X(n4731) );
  nand_x1_sg U6342 ( .A(n4693), .B(n4694), .X(n4692) );
  nand_x1_sg U6343 ( .A(n4615), .B(n4616), .X(n4614) );
  nand_x1_sg U6344 ( .A(n4576), .B(n4577), .X(n4575) );
  nand_x1_sg U6345 ( .A(n4498), .B(n4499), .X(n4497) );
  nand_x1_sg U6346 ( .A(n4455), .B(n4456), .X(n4454) );
  nand_x1_sg U6347 ( .A(n5122), .B(n5123), .X(n5121) );
  nand_x1_sg U6348 ( .A(n5005), .B(n5006), .X(n5004) );
  nand_x1_sg U6349 ( .A(n4888), .B(n4889), .X(n4887) );
  nand_x1_sg U6350 ( .A(n4771), .B(n4772), .X(n4770) );
  nand_x1_sg U6351 ( .A(n4654), .B(n4655), .X(n4653) );
  nand_x1_sg U6352 ( .A(n4537), .B(n4538), .X(n4536) );
  nand_x1_sg U6353 ( .A(n5096), .B(n5097), .X(n5095) );
  nand_x1_sg U6354 ( .A(n4979), .B(n4980), .X(n4978) );
  nand_x1_sg U6355 ( .A(n4862), .B(n4863), .X(n4861) );
  nand_x1_sg U6356 ( .A(n4745), .B(n4746), .X(n4744) );
  nand_x1_sg U6357 ( .A(n4628), .B(n4629), .X(n4627) );
  nand_x1_sg U6358 ( .A(n4511), .B(n4512), .X(n4510) );
  nand_x1_sg U6359 ( .A(n3506), .B(n5916), .X(n3505) );
  nand_x1_sg U6360 ( .A(n3510), .B(n3288), .X(n3504) );
  nor_x1_sg U6361 ( .A(n3507), .B(n3311), .X(n3506) );
  nor_x1_sg U6362 ( .A(n5918), .B(n5218), .X(n4418) );
  nand_x1_sg U6363 ( .A(n3262), .B(n5345), .X(n3702) );
  nand_x1_sg U6364 ( .A(n5887), .B(n5835), .X(n4213) );
  inv_x1_sg U6365 ( .A(n3447), .X(n3356) );
  nand_x1_sg U6366 ( .A(n3258), .B(n5835), .X(n4383) );
  nor_x1_sg U6367 ( .A(n5314), .B(n3333), .X(n4396) );
  nor_x1_sg U6368 ( .A(n5831), .B(n5907), .X(n4401) );
  nor_x1_sg U6369 ( .A(n3512), .B(n5826), .X(n3511) );
  nand_x1_sg U6370 ( .A(n3465), .B(n3488), .X(n3487) );
  nand_x1_sg U6371 ( .A(n3512), .B(n5826), .X(n3510) );
  nor_x1_sg U6372 ( .A(n3371), .B(n4401), .X(n4400) );
  nand_x1_sg U6373 ( .A(n3497), .B(n3366), .X(n3495) );
  nor_x1_sg U6374 ( .A(n5918), .B(n5336), .X(n5940) );
  nor_x1_sg U6375 ( .A(n5167), .B(n5941), .X(N142) );
  nor_x1_sg U6376 ( .A(n5128), .B(n5942), .X(N143) );
  nor_x1_sg U6377 ( .A(n5050), .B(n5941), .X(N145) );
  nor_x1_sg U6378 ( .A(n5011), .B(n5941), .X(N146) );
  nor_x1_sg U6379 ( .A(n4933), .B(n4407), .X(N148) );
  nor_x1_sg U6380 ( .A(n4894), .B(n5843), .X(N149) );
  nor_x1_sg U6381 ( .A(n4816), .B(n4407), .X(N151) );
  nor_x1_sg U6382 ( .A(n4777), .B(n5920), .X(N152) );
  nor_x1_sg U6383 ( .A(n4699), .B(n4407), .X(N154) );
  nor_x1_sg U6384 ( .A(n4660), .B(n5920), .X(N155) );
  nor_x1_sg U6385 ( .A(n4582), .B(n5921), .X(N157) );
  nor_x1_sg U6386 ( .A(n4543), .B(n5942), .X(N158) );
  nor_x1_sg U6387 ( .A(n4465), .B(n5843), .X(N160) );
  nor_x1_sg U6388 ( .A(n4408), .B(n5942), .X(N161) );
  nor_x1_sg U6389 ( .A(n5089), .B(n5843), .X(N144) );
  nor_x1_sg U6390 ( .A(n4972), .B(n5941), .X(N147) );
  nor_x1_sg U6391 ( .A(n4855), .B(n5921), .X(N150) );
  nor_x1_sg U6392 ( .A(n4738), .B(n5921), .X(N153) );
  nor_x1_sg U6393 ( .A(n4621), .B(n5942), .X(N156) );
  nor_x1_sg U6394 ( .A(n4504), .B(n5920), .X(N159) );
  nand_x1_sg U6395 ( .A(n5178), .B(n4396), .X(n5938) );
  nand_x1_sg U6396 ( .A(n5915), .B(n3509), .X(n3508) );
  nor_x1_sg U6397 ( .A(n5218), .B(n5181), .X(n5939) );
  nor_x1_sg U6398 ( .A(n5336), .B(n5181), .X(n5936) );
  nor_x1_sg U6399 ( .A(n5915), .B(n3509), .X(n3507) );
  nor_x1_sg U6400 ( .A(n5191), .B(n5177), .X(n4437) );
  inv_x1_sg U6401 ( .A(n5184), .X(n3335) );
  nand_x1_sg U6402 ( .A(n3335), .B(n5888), .X(n3499) );
  nand_x1_sg U6403 ( .A(n3435), .B(n3439), .X(n3438) );
  nor_x1_sg U6404 ( .A(n3442), .B(n3443), .X(n3441) );
  inv_x1_sg U6405 ( .A(n3484), .X(n3359) );
  inv_x1_sg U6406 ( .A(n3479), .X(n3361) );
  nor_x1_sg U6407 ( .A(n5888), .B(n5337), .X(n4464) );
  nor_x1_sg U6408 ( .A(n5336), .B(n5202), .X(n5933) );
  nor_x1_sg U6409 ( .A(n5202), .B(n5177), .X(n5932) );
  nor_x1_sg U6410 ( .A(n5191), .B(n5313), .X(n5935) );
  nor_x1_sg U6411 ( .A(n5313), .B(n5344), .X(n4460) );
  nor_x1_sg U6412 ( .A(n5191), .B(n5336), .X(n4433) );
  nor_x1_sg U6413 ( .A(n3335), .B(n5202), .X(n5934) );
  nor_x1_sg U6414 ( .A(n5316), .B(n3456), .X(n3454) );
  nand_x1_sg U6415 ( .A(n5316), .B(n3456), .X(n3455) );
  nor_x1_sg U6416 ( .A(n5177), .B(n5344), .X(n5931) );
  nor_x1_sg U6417 ( .A(n5907), .B(n3362), .X(n3457) );
  inv_x1_sg U6418 ( .A(n3459), .X(n3362) );
  nand_x1_sg U6419 ( .A(n3261), .B(n3469), .X(n3789) );
  nand_x1_sg U6420 ( .A(n5887), .B(n5323), .X(n4129) );
  nand_x1_sg U6421 ( .A(n3261), .B(n5321), .X(n3831) );
  nand_x1_sg U6422 ( .A(n5887), .B(n3468), .X(n4171) );
  nand_x1_sg U6423 ( .A(n3260), .B(n5321), .X(n4001) );
  nand_x1_sg U6424 ( .A(n3261), .B(n3576), .X(n3747) );
  nand_x1_sg U6425 ( .A(n5887), .B(n3576), .X(n4087) );
  nand_x1_sg U6426 ( .A(n3260), .B(n5220), .X(n3917) );
  nand_x1_sg U6427 ( .A(n3704), .B(n3705), .X(n3703) );
  nor_x1_sg U6428 ( .A(n5324), .B(n3366), .X(n4215) );
  nand_x1_sg U6429 ( .A(n3468), .B(n3262), .X(n3660) );
  nand_x1_sg U6430 ( .A(n3261), .B(n5345), .X(n3873) );
  nand_x1_sg U6431 ( .A(n3260), .B(n5345), .X(n4043) );
  nand_x1_sg U6432 ( .A(n3469), .B(n3262), .X(n3618) );
  nand_x1_sg U6433 ( .A(n5220), .B(n3262), .X(n3575) );
  nor_x1_sg U6434 ( .A(n5321), .B(n5323), .X(n3447) );
  nand_x1_sg U6435 ( .A(n3258), .B(n3468), .X(n4341) );
  nand_x1_sg U6436 ( .A(n3258), .B(n3469), .X(n4299) );
  nand_x1_sg U6437 ( .A(n4385), .B(n3704), .X(n4384) );
  nor_x1_sg U6438 ( .A(n5826), .B(n5819), .X(n4385) );
  nand_x1_sg U6439 ( .A(n3258), .B(n3576), .X(n4257) );
  nor_x1_sg U6440 ( .A(n5919), .B(n5822), .X(n5948) );
  nor_x1_sg U6441 ( .A(n5908), .B(n5824), .X(n3520) );
  nor_x1_sg U6442 ( .A(n3282), .B(n5819), .X(n3526) );
  nor_x1_sg U6443 ( .A(n5909), .B(n5821), .X(n3550) );
  nand_x1_sg U6444 ( .A(n4401), .B(rd_ptr[3]), .X(n4406) );
  inv_x1_sg U6445 ( .A(rd_ptr[0]), .X(n3333) );
  nand_x1_sg U6446 ( .A(empty), .B(n3236), .X(n3485) );
  nor_x1_sg U6447 ( .A(n3236), .B(n3435), .X(n3486) );
  nand_x1_sg U6448 ( .A(n5338), .B(n4406), .X(n4405) );
  nand_x1_sg U6449 ( .A(n5813), .B(n5344), .X(n4404) );
  nand_x1_sg U6450 ( .A(n5342), .B(n3290), .X(n3496) );
  nand_x1_sg U6451 ( .A(n5343), .B(n3499), .X(n3498) );
  nand_x1_sg U6452 ( .A(n5814), .B(n5338), .X(n3501) );
  nor_x1_sg U6453 ( .A(n5185), .B(n5340), .X(n5178) );
  nand_x1_sg U6454 ( .A(n5337), .B(n3371), .X(n5185) );
  nand_x1_sg U6455 ( .A(n5175), .B(n5176), .X(n5174) );
  nand_x1_sg U6456 ( .A(n5465), .B(\buff_mem[4][0] ), .X(n5180) );
  nand_x1_sg U6457 ( .A(n5135), .B(n5136), .X(n5134) );
  nand_x1_sg U6458 ( .A(n5463), .B(\buff_mem[4][1] ), .X(n5138) );
  nand_x1_sg U6459 ( .A(n5057), .B(n5058), .X(n5056) );
  nand_x1_sg U6460 ( .A(n5464), .B(\buff_mem[4][3] ), .X(n5060) );
  nand_x1_sg U6461 ( .A(n5018), .B(n5019), .X(n5017) );
  nand_x1_sg U6462 ( .A(n5465), .B(\buff_mem[4][4] ), .X(n5021) );
  nand_x1_sg U6463 ( .A(n4940), .B(n4941), .X(n4939) );
  nand_x1_sg U6464 ( .A(n5463), .B(\buff_mem[4][6] ), .X(n4943) );
  nand_x1_sg U6465 ( .A(n4901), .B(n4902), .X(n4900) );
  nand_x1_sg U6466 ( .A(n5462), .B(\buff_mem[4][7] ), .X(n4904) );
  nand_x1_sg U6467 ( .A(n4823), .B(n4824), .X(n4822) );
  nand_x1_sg U6468 ( .A(n5462), .B(\buff_mem[4][9] ), .X(n4826) );
  nand_x1_sg U6469 ( .A(n4784), .B(n4785), .X(n4783) );
  nand_x1_sg U6470 ( .A(n5262), .B(\buff_mem[4][10] ), .X(n4787) );
  nand_x1_sg U6471 ( .A(n4706), .B(n4707), .X(n4705) );
  nand_x1_sg U6472 ( .A(n5464), .B(\buff_mem[4][12] ), .X(n4709) );
  nand_x1_sg U6473 ( .A(n4667), .B(n4668), .X(n4666) );
  nand_x1_sg U6474 ( .A(n5465), .B(\buff_mem[4][13] ), .X(n4670) );
  nand_x1_sg U6475 ( .A(n4589), .B(n4590), .X(n4588) );
  nand_x1_sg U6476 ( .A(n5262), .B(\buff_mem[4][15] ), .X(n4592) );
  nand_x1_sg U6477 ( .A(n4550), .B(n4551), .X(n4549) );
  nand_x1_sg U6478 ( .A(n5462), .B(\buff_mem[4][16] ), .X(n4553) );
  nand_x1_sg U6479 ( .A(n4472), .B(n4473), .X(n4471) );
  nand_x1_sg U6480 ( .A(n5462), .B(\buff_mem[4][18] ), .X(n4475) );
  nand_x1_sg U6481 ( .A(n4415), .B(n4416), .X(n4414) );
  nand_x1_sg U6482 ( .A(n5464), .B(\buff_mem[4][19] ), .X(n4420) );
  nand_x1_sg U6483 ( .A(n5453), .B(\buff_mem[1][0] ), .X(n5176) );
  nand_x1_sg U6484 ( .A(n5453), .B(\buff_mem[1][1] ), .X(n5136) );
  nand_x1_sg U6485 ( .A(n5260), .B(\buff_mem[1][3] ), .X(n5058) );
  nand_x1_sg U6486 ( .A(n5453), .B(\buff_mem[1][4] ), .X(n5019) );
  nand_x1_sg U6487 ( .A(n5452), .B(\buff_mem[1][6] ), .X(n4941) );
  nand_x1_sg U6488 ( .A(n5450), .B(\buff_mem[1][7] ), .X(n4902) );
  nand_x1_sg U6489 ( .A(n5451), .B(\buff_mem[1][9] ), .X(n4824) );
  nand_x1_sg U6490 ( .A(n5260), .B(\buff_mem[1][10] ), .X(n4785) );
  nand_x1_sg U6491 ( .A(n5452), .B(\buff_mem[1][12] ), .X(n4707) );
  nand_x1_sg U6492 ( .A(n5451), .B(\buff_mem[1][13] ), .X(n4668) );
  nand_x1_sg U6493 ( .A(n5450), .B(\buff_mem[1][15] ), .X(n4590) );
  nand_x1_sg U6494 ( .A(n5452), .B(\buff_mem[1][16] ), .X(n4551) );
  nand_x1_sg U6495 ( .A(n5451), .B(\buff_mem[1][18] ), .X(n4473) );
  nand_x1_sg U6496 ( .A(n5260), .B(\buff_mem[1][19] ), .X(n4416) );
  nand_x1_sg U6497 ( .A(n5448), .B(\buff_mem[0][0] ), .X(n5175) );
  nand_x1_sg U6498 ( .A(n5446), .B(\buff_mem[0][1] ), .X(n5135) );
  nand_x1_sg U6499 ( .A(n5258), .B(\buff_mem[0][3] ), .X(n5057) );
  nand_x1_sg U6500 ( .A(n5448), .B(\buff_mem[0][4] ), .X(n5018) );
  nand_x1_sg U6501 ( .A(n5447), .B(\buff_mem[0][6] ), .X(n4940) );
  nand_x1_sg U6502 ( .A(n5445), .B(\buff_mem[0][7] ), .X(n4901) );
  nand_x1_sg U6503 ( .A(n5446), .B(\buff_mem[0][9] ), .X(n4823) );
  nand_x1_sg U6504 ( .A(n5446), .B(\buff_mem[0][10] ), .X(n4784) );
  nand_x1_sg U6505 ( .A(n5448), .B(\buff_mem[0][12] ), .X(n4706) );
  nand_x1_sg U6506 ( .A(n5446), .B(\buff_mem[0][13] ), .X(n4667) );
  nand_x1_sg U6507 ( .A(n5258), .B(\buff_mem[0][15] ), .X(n4589) );
  nand_x1_sg U6508 ( .A(n5447), .B(\buff_mem[0][16] ), .X(n4550) );
  nand_x1_sg U6509 ( .A(n5448), .B(\buff_mem[0][18] ), .X(n4472) );
  nand_x1_sg U6510 ( .A(n5445), .B(\buff_mem[0][19] ), .X(n4415) );
  nand_x1_sg U6511 ( .A(n5258), .B(\buff_mem[0][2] ), .X(n5096) );
  nand_x1_sg U6512 ( .A(n5447), .B(\buff_mem[0][5] ), .X(n4979) );
  nand_x1_sg U6513 ( .A(n5445), .B(\buff_mem[0][8] ), .X(n4862) );
  nand_x1_sg U6514 ( .A(n5258), .B(\buff_mem[0][11] ), .X(n4745) );
  nand_x1_sg U6515 ( .A(n5445), .B(\buff_mem[0][14] ), .X(n4628) );
  nand_x1_sg U6516 ( .A(n5447), .B(\buff_mem[0][17] ), .X(n4511) );
  nand_x1_sg U6517 ( .A(n5464), .B(\buff_mem[4][2] ), .X(n5099) );
  nand_x1_sg U6518 ( .A(n5463), .B(\buff_mem[4][5] ), .X(n4982) );
  nand_x1_sg U6519 ( .A(n5262), .B(\buff_mem[4][8] ), .X(n4865) );
  nand_x1_sg U6520 ( .A(n5262), .B(\buff_mem[4][11] ), .X(n4748) );
  nand_x1_sg U6521 ( .A(n5465), .B(\buff_mem[4][14] ), .X(n4631) );
  nand_x1_sg U6522 ( .A(n5463), .B(\buff_mem[4][17] ), .X(n4514) );
  nand_x1_sg U6523 ( .A(n5450), .B(\buff_mem[1][2] ), .X(n5097) );
  nand_x1_sg U6524 ( .A(n5450), .B(\buff_mem[1][5] ), .X(n4980) );
  nand_x1_sg U6525 ( .A(n5451), .B(\buff_mem[1][8] ), .X(n4863) );
  nand_x1_sg U6526 ( .A(n5260), .B(\buff_mem[1][11] ), .X(n4746) );
  nand_x1_sg U6527 ( .A(n5452), .B(\buff_mem[1][14] ), .X(n4629) );
  nand_x1_sg U6528 ( .A(n5453), .B(\buff_mem[1][17] ), .X(n4512) );
  nand_x1_sg U6529 ( .A(\buff_mem[15][0] ), .B(n5333), .X(n5209) );
  nand_x1_sg U6530 ( .A(\buff_mem[15][1] ), .B(n5816), .X(n5162) );
  nand_x1_sg U6531 ( .A(\buff_mem[15][2] ), .B(n5814), .X(n5123) );
  nand_x1_sg U6532 ( .A(\buff_mem[15][3] ), .B(n5333), .X(n5084) );
  nand_x1_sg U6533 ( .A(\buff_mem[15][4] ), .B(n5814), .X(n5045) );
  nand_x1_sg U6534 ( .A(\buff_mem[15][5] ), .B(n5813), .X(n5006) );
  nand_x1_sg U6535 ( .A(\buff_mem[15][6] ), .B(n5816), .X(n4967) );
  nand_x1_sg U6536 ( .A(\buff_mem[15][7] ), .B(n5813), .X(n4928) );
  nand_x1_sg U6537 ( .A(\buff_mem[15][8] ), .B(n5334), .X(n4889) );
  nand_x1_sg U6538 ( .A(\buff_mem[15][9] ), .B(n5333), .X(n4850) );
  nand_x1_sg U6539 ( .A(\buff_mem[15][10] ), .B(n5334), .X(n4811) );
  nand_x1_sg U6540 ( .A(\buff_mem[15][11] ), .B(n5815), .X(n4772) );
  nand_x1_sg U6541 ( .A(\buff_mem[15][12] ), .B(n5813), .X(n4733) );
  nand_x1_sg U6542 ( .A(\buff_mem[15][13] ), .B(n5815), .X(n4694) );
  nand_x1_sg U6543 ( .A(\buff_mem[15][14] ), .B(n5815), .X(n4655) );
  nand_x1_sg U6544 ( .A(\buff_mem[15][15] ), .B(n5814), .X(n4616) );
  nand_x1_sg U6545 ( .A(\buff_mem[15][16] ), .B(n5815), .X(n4577) );
  nand_x1_sg U6546 ( .A(\buff_mem[15][17] ), .B(n5816), .X(n4538) );
  nand_x1_sg U6547 ( .A(\buff_mem[15][18] ), .B(n5334), .X(n4499) );
  nand_x1_sg U6548 ( .A(\buff_mem[15][19] ), .B(n5816), .X(n4456) );
  nand_x1_sg U6549 ( .A(n5500), .B(\buff_mem[19][0] ), .X(n5211) );
  nand_x1_sg U6550 ( .A(n5503), .B(\buff_mem[19][1] ), .X(n5164) );
  nand_x1_sg U6551 ( .A(n5501), .B(\buff_mem[19][3] ), .X(n5086) );
  nand_x1_sg U6552 ( .A(n5503), .B(\buff_mem[19][4] ), .X(n5047) );
  nand_x1_sg U6553 ( .A(n5502), .B(\buff_mem[19][6] ), .X(n4969) );
  nand_x1_sg U6554 ( .A(n5274), .B(\buff_mem[19][7] ), .X(n4930) );
  nand_x1_sg U6555 ( .A(n5503), .B(\buff_mem[19][9] ), .X(n4852) );
  nand_x1_sg U6556 ( .A(n5500), .B(\buff_mem[19][10] ), .X(n4813) );
  nand_x1_sg U6557 ( .A(n5500), .B(\buff_mem[19][12] ), .X(n4735) );
  nand_x1_sg U6558 ( .A(n5502), .B(\buff_mem[19][13] ), .X(n4696) );
  nand_x1_sg U6559 ( .A(n5274), .B(\buff_mem[19][15] ), .X(n4618) );
  nand_x1_sg U6560 ( .A(n5502), .B(\buff_mem[19][16] ), .X(n4579) );
  nand_x1_sg U6561 ( .A(n5503), .B(\buff_mem[19][18] ), .X(n4501) );
  nand_x1_sg U6562 ( .A(n5501), .B(\buff_mem[19][19] ), .X(n4459) );
  nand_x1_sg U6563 ( .A(n5501), .B(\buff_mem[19][2] ), .X(n5125) );
  nand_x1_sg U6564 ( .A(n5502), .B(\buff_mem[19][5] ), .X(n5008) );
  nand_x1_sg U6565 ( .A(n5274), .B(\buff_mem[19][8] ), .X(n4891) );
  nand_x1_sg U6566 ( .A(n5501), .B(\buff_mem[19][11] ), .X(n4774) );
  nand_x1_sg U6567 ( .A(n5274), .B(\buff_mem[19][14] ), .X(n4657) );
  nand_x1_sg U6568 ( .A(n5500), .B(\buff_mem[19][17] ), .X(n4540) );
  nor_x1_sg U6569 ( .A(n5182), .B(n5183), .X(n5179) );
  nor_x1_sg U6570 ( .A(n3412), .B(n5454), .X(n5183) );
  nor_x1_sg U6571 ( .A(n3413), .B(n5417), .X(n5182) );
  inv_x1_sg U6572 ( .A(\buff_mem[3][0] ), .X(n3412) );
  nor_x1_sg U6573 ( .A(n5139), .B(n5140), .X(n5137) );
  nor_x1_sg U6574 ( .A(n3409), .B(n5458), .X(n5140) );
  nor_x1_sg U6575 ( .A(n3410), .B(n5416), .X(n5139) );
  inv_x1_sg U6576 ( .A(\buff_mem[3][1] ), .X(n3409) );
  nor_x1_sg U6577 ( .A(n5061), .B(n5062), .X(n5059) );
  nor_x1_sg U6578 ( .A(n3403), .B(n5459), .X(n5062) );
  nor_x1_sg U6579 ( .A(n3404), .B(n5417), .X(n5061) );
  inv_x1_sg U6580 ( .A(\buff_mem[3][3] ), .X(n3403) );
  nor_x1_sg U6581 ( .A(n5022), .B(n5023), .X(n5020) );
  nor_x1_sg U6582 ( .A(n3400), .B(n5454), .X(n5023) );
  nor_x1_sg U6583 ( .A(n3401), .B(n5418), .X(n5022) );
  inv_x1_sg U6584 ( .A(\buff_mem[3][4] ), .X(n3400) );
  nor_x1_sg U6585 ( .A(n4944), .B(n4945), .X(n4942) );
  nor_x1_sg U6586 ( .A(n3394), .B(n5459), .X(n4945) );
  nor_x1_sg U6587 ( .A(n3395), .B(n5415), .X(n4944) );
  inv_x1_sg U6588 ( .A(\buff_mem[3][6] ), .X(n3394) );
  nor_x1_sg U6589 ( .A(n4905), .B(n4906), .X(n4903) );
  nor_x1_sg U6590 ( .A(n3391), .B(n5457), .X(n4906) );
  nor_x1_sg U6591 ( .A(n3392), .B(n5417), .X(n4905) );
  inv_x1_sg U6592 ( .A(\buff_mem[3][7] ), .X(n3391) );
  nor_x1_sg U6593 ( .A(n4827), .B(n4828), .X(n4825) );
  nor_x1_sg U6594 ( .A(n3385), .B(n5457), .X(n4828) );
  nor_x1_sg U6595 ( .A(n3386), .B(n5415), .X(n4827) );
  inv_x1_sg U6596 ( .A(\buff_mem[3][9] ), .X(n3385) );
  nor_x1_sg U6597 ( .A(n4788), .B(n4789), .X(n4786) );
  nor_x1_sg U6598 ( .A(n3382), .B(n5460), .X(n4789) );
  nor_x1_sg U6599 ( .A(n3383), .B(n5418), .X(n4788) );
  inv_x1_sg U6600 ( .A(\buff_mem[3][10] ), .X(n3382) );
  nor_x1_sg U6601 ( .A(n4710), .B(n4711), .X(n4708) );
  nor_x1_sg U6602 ( .A(n3376), .B(n5457), .X(n4711) );
  nor_x1_sg U6603 ( .A(n3377), .B(n5415), .X(n4710) );
  inv_x1_sg U6604 ( .A(\buff_mem[3][12] ), .X(n3376) );
  nor_x1_sg U6605 ( .A(n4671), .B(n4672), .X(n4669) );
  nor_x1_sg U6606 ( .A(n3373), .B(n5458), .X(n4672) );
  nor_x1_sg U6607 ( .A(n3374), .B(n5412), .X(n4671) );
  inv_x1_sg U6608 ( .A(\buff_mem[3][13] ), .X(n3373) );
  nor_x1_sg U6609 ( .A(n4593), .B(n4594), .X(n4591) );
  nor_x1_sg U6610 ( .A(n3427), .B(n5459), .X(n4594) );
  nor_x1_sg U6611 ( .A(n3428), .B(n5412), .X(n4593) );
  inv_x1_sg U6612 ( .A(\buff_mem[3][15] ), .X(n3427) );
  nor_x1_sg U6613 ( .A(n4554), .B(n4555), .X(n4552) );
  nor_x1_sg U6614 ( .A(n3424), .B(n5458), .X(n4555) );
  nor_x1_sg U6615 ( .A(n3425), .B(n5415), .X(n4554) );
  inv_x1_sg U6616 ( .A(\buff_mem[3][16] ), .X(n3424) );
  nor_x1_sg U6617 ( .A(n4476), .B(n4477), .X(n4474) );
  nor_x1_sg U6618 ( .A(n3418), .B(n5454), .X(n4477) );
  nor_x1_sg U6619 ( .A(n3419), .B(n5416), .X(n4476) );
  inv_x1_sg U6620 ( .A(\buff_mem[3][18] ), .X(n3418) );
  nor_x1_sg U6621 ( .A(n4422), .B(n4423), .X(n4419) );
  nor_x1_sg U6622 ( .A(n3415), .B(n5460), .X(n4423) );
  nor_x1_sg U6623 ( .A(n3416), .B(n5412), .X(n4422) );
  inv_x1_sg U6624 ( .A(\buff_mem[3][19] ), .X(n3415) );
  nand_x1_sg U6625 ( .A(n5383), .B(\buff_mem[6][2] ), .X(n5105) );
  nand_x1_sg U6626 ( .A(n5236), .B(\buff_mem[6][5] ), .X(n4988) );
  nand_x1_sg U6627 ( .A(n5384), .B(\buff_mem[6][8] ), .X(n4871) );
  nand_x1_sg U6628 ( .A(n5236), .B(\buff_mem[6][11] ), .X(n4754) );
  nand_x1_sg U6629 ( .A(n5386), .B(\buff_mem[6][14] ), .X(n4637) );
  nand_x1_sg U6630 ( .A(n5385), .B(\buff_mem[6][17] ), .X(n4520) );
  nand_x1_sg U6631 ( .A(\buff_mem[8][0] ), .B(n5473), .X(n5194) );
  nand_x1_sg U6632 ( .A(\buff_mem[7][0] ), .B(n5693), .X(n5193) );
  nand_x1_sg U6633 ( .A(\buff_mem[8][1] ), .B(n5472), .X(n5148) );
  nand_x1_sg U6634 ( .A(\buff_mem[7][1] ), .B(n5695), .X(n5147) );
  nand_x1_sg U6635 ( .A(\buff_mem[8][2] ), .B(n5472), .X(n5109) );
  nand_x1_sg U6636 ( .A(\buff_mem[7][2] ), .B(n5696), .X(n5108) );
  nand_x1_sg U6637 ( .A(\buff_mem[8][3] ), .B(n5473), .X(n5070) );
  nand_x1_sg U6638 ( .A(\buff_mem[7][3] ), .B(n5693), .X(n5069) );
  nand_x1_sg U6639 ( .A(\buff_mem[8][4] ), .B(n5474), .X(n5031) );
  nand_x1_sg U6640 ( .A(\buff_mem[7][4] ), .B(n5696), .X(n5030) );
  nand_x1_sg U6641 ( .A(\buff_mem[8][5] ), .B(n5266), .X(n4992) );
  nand_x1_sg U6642 ( .A(\buff_mem[7][5] ), .B(n5697), .X(n4991) );
  nand_x1_sg U6643 ( .A(\buff_mem[8][6] ), .B(n5472), .X(n4953) );
  nand_x1_sg U6644 ( .A(\buff_mem[7][6] ), .B(n5694), .X(n4952) );
  nand_x1_sg U6645 ( .A(\buff_mem[8][7] ), .B(n5474), .X(n4914) );
  nand_x1_sg U6646 ( .A(\buff_mem[7][7] ), .B(n5697), .X(n4913) );
  nand_x1_sg U6647 ( .A(\buff_mem[8][8] ), .B(n5475), .X(n4875) );
  nand_x1_sg U6648 ( .A(\buff_mem[7][8] ), .B(n5697), .X(n4874) );
  nand_x1_sg U6649 ( .A(\buff_mem[8][9] ), .B(n5266), .X(n4836) );
  nand_x1_sg U6650 ( .A(\buff_mem[7][9] ), .B(n5694), .X(n4835) );
  nand_x1_sg U6651 ( .A(\buff_mem[8][10] ), .B(n5475), .X(n4797) );
  nand_x1_sg U6652 ( .A(\buff_mem[7][10] ), .B(n5697), .X(n4796) );
  nand_x1_sg U6653 ( .A(\buff_mem[8][11] ), .B(n5474), .X(n4758) );
  nand_x1_sg U6654 ( .A(\buff_mem[7][11] ), .B(n5695), .X(n4757) );
  nand_x1_sg U6655 ( .A(\buff_mem[8][12] ), .B(n5473), .X(n4719) );
  nand_x1_sg U6656 ( .A(\buff_mem[7][12] ), .B(n5695), .X(n4718) );
  nand_x1_sg U6657 ( .A(\buff_mem[8][13] ), .B(n5473), .X(n4680) );
  nand_x1_sg U6658 ( .A(\buff_mem[7][13] ), .B(n5695), .X(n4679) );
  nand_x1_sg U6659 ( .A(\buff_mem[8][14] ), .B(n5475), .X(n4641) );
  nand_x1_sg U6660 ( .A(\buff_mem[7][14] ), .B(n5694), .X(n4640) );
  nand_x1_sg U6661 ( .A(\buff_mem[8][15] ), .B(n5266), .X(n4602) );
  nand_x1_sg U6662 ( .A(\buff_mem[7][15] ), .B(n5693), .X(n4601) );
  nand_x1_sg U6663 ( .A(\buff_mem[8][16] ), .B(n5474), .X(n4563) );
  nand_x1_sg U6664 ( .A(\buff_mem[7][16] ), .B(n5696), .X(n4562) );
  nand_x1_sg U6665 ( .A(\buff_mem[8][17] ), .B(n5472), .X(n4524) );
  nand_x1_sg U6666 ( .A(\buff_mem[7][17] ), .B(n5693), .X(n4523) );
  nand_x1_sg U6667 ( .A(\buff_mem[8][18] ), .B(n5266), .X(n4485) );
  nand_x1_sg U6668 ( .A(\buff_mem[7][18] ), .B(n5694), .X(n4484) );
  nand_x1_sg U6669 ( .A(\buff_mem[8][19] ), .B(n5475), .X(n4436) );
  nand_x1_sg U6670 ( .A(\buff_mem[7][19] ), .B(n5696), .X(n4435) );
  nand_x1_sg U6671 ( .A(n5385), .B(\buff_mem[6][0] ), .X(n5189) );
  nand_x1_sg U6672 ( .A(n5383), .B(\buff_mem[6][1] ), .X(n5144) );
  nand_x1_sg U6673 ( .A(n5384), .B(\buff_mem[6][3] ), .X(n5066) );
  nand_x1_sg U6674 ( .A(n5386), .B(\buff_mem[6][4] ), .X(n5027) );
  nand_x1_sg U6675 ( .A(n5384), .B(\buff_mem[6][6] ), .X(n4949) );
  nand_x1_sg U6676 ( .A(n5236), .B(\buff_mem[6][7] ), .X(n4910) );
  nand_x1_sg U6677 ( .A(n5386), .B(\buff_mem[6][9] ), .X(n4832) );
  nand_x1_sg U6678 ( .A(n5383), .B(\buff_mem[6][10] ), .X(n4793) );
  nand_x1_sg U6679 ( .A(n5236), .B(\buff_mem[6][12] ), .X(n4715) );
  nand_x1_sg U6680 ( .A(n5385), .B(\buff_mem[6][13] ), .X(n4676) );
  nand_x1_sg U6681 ( .A(n5384), .B(\buff_mem[6][15] ), .X(n4598) );
  nand_x1_sg U6682 ( .A(n5386), .B(\buff_mem[6][16] ), .X(n4559) );
  nand_x1_sg U6683 ( .A(n5385), .B(\buff_mem[6][18] ), .X(n4481) );
  nand_x1_sg U6684 ( .A(n5383), .B(\buff_mem[6][19] ), .X(n4429) );
  nor_x1_sg U6685 ( .A(n5100), .B(n5101), .X(n5098) );
  nor_x1_sg U6686 ( .A(n3406), .B(n5460), .X(n5101) );
  nor_x1_sg U6687 ( .A(n3407), .B(n5416), .X(n5100) );
  inv_x1_sg U6688 ( .A(\buff_mem[3][2] ), .X(n3406) );
  nor_x1_sg U6689 ( .A(n4983), .B(n4984), .X(n4981) );
  nor_x1_sg U6690 ( .A(n3397), .B(n5459), .X(n4984) );
  nor_x1_sg U6691 ( .A(n3398), .B(n5418), .X(n4983) );
  inv_x1_sg U6692 ( .A(\buff_mem[3][5] ), .X(n3397) );
  nor_x1_sg U6693 ( .A(n4866), .B(n4867), .X(n4864) );
  nor_x1_sg U6694 ( .A(n3388), .B(n5460), .X(n4867) );
  nor_x1_sg U6695 ( .A(n3389), .B(n5412), .X(n4866) );
  inv_x1_sg U6696 ( .A(\buff_mem[3][8] ), .X(n3388) );
  nor_x1_sg U6697 ( .A(n4749), .B(n4750), .X(n4747) );
  nor_x1_sg U6698 ( .A(n3379), .B(n5454), .X(n4750) );
  nor_x1_sg U6699 ( .A(n3380), .B(n5418), .X(n4749) );
  inv_x1_sg U6700 ( .A(\buff_mem[3][11] ), .X(n3379) );
  nor_x1_sg U6701 ( .A(n4632), .B(n4633), .X(n4630) );
  nor_x1_sg U6702 ( .A(n3430), .B(n5458), .X(n4633) );
  nor_x1_sg U6703 ( .A(n3431), .B(n5417), .X(n4632) );
  inv_x1_sg U6704 ( .A(\buff_mem[3][14] ), .X(n3430) );
  nor_x1_sg U6705 ( .A(n4515), .B(n4516), .X(n4513) );
  nor_x1_sg U6706 ( .A(n3421), .B(n5457), .X(n4516) );
  nor_x1_sg U6707 ( .A(n3422), .B(n5416), .X(n4515) );
  inv_x1_sg U6708 ( .A(\buff_mem[3][17] ), .X(n3421) );
  nand_x1_sg U6709 ( .A(n4396), .B(n5907), .X(n4394) );
  nand_x1_sg U6710 ( .A(n5340), .B(n5831), .X(n4395) );
  nand_x1_sg U6711 ( .A(n5338), .B(n5913), .X(n4402) );
  nand_x1_sg U6712 ( .A(n5906), .B(n3512), .X(n4403) );
  nand_x1_sg U6713 ( .A(n5468), .B(\buff_mem[5][0] ), .X(n5188) );
  nand_x1_sg U6714 ( .A(n5469), .B(\buff_mem[5][1] ), .X(n5143) );
  nand_x1_sg U6715 ( .A(n5467), .B(\buff_mem[5][3] ), .X(n5065) );
  nand_x1_sg U6716 ( .A(n5470), .B(\buff_mem[5][4] ), .X(n5026) );
  nand_x1_sg U6717 ( .A(n5264), .B(\buff_mem[5][6] ), .X(n4948) );
  nand_x1_sg U6718 ( .A(n5469), .B(\buff_mem[5][7] ), .X(n4909) );
  nand_x1_sg U6719 ( .A(n5470), .B(\buff_mem[5][9] ), .X(n4831) );
  nand_x1_sg U6720 ( .A(n5467), .B(\buff_mem[5][10] ), .X(n4792) );
  nand_x1_sg U6721 ( .A(n5467), .B(\buff_mem[5][12] ), .X(n4714) );
  nand_x1_sg U6722 ( .A(n5468), .B(\buff_mem[5][13] ), .X(n4675) );
  nand_x1_sg U6723 ( .A(n5264), .B(\buff_mem[5][15] ), .X(n4597) );
  nand_x1_sg U6724 ( .A(n5470), .B(\buff_mem[5][16] ), .X(n4558) );
  nand_x1_sg U6725 ( .A(n5468), .B(\buff_mem[5][18] ), .X(n4480) );
  nand_x1_sg U6726 ( .A(n5264), .B(\buff_mem[5][19] ), .X(n4428) );
  inv_x1_sg U6727 ( .A(rd_ptr[3]), .X(n3371) );
  nand_x1_sg U6728 ( .A(n5264), .B(\buff_mem[5][2] ), .X(n5104) );
  nand_x1_sg U6729 ( .A(n5469), .B(\buff_mem[5][5] ), .X(n4987) );
  nand_x1_sg U6730 ( .A(n5469), .B(\buff_mem[5][8] ), .X(n4870) );
  nand_x1_sg U6731 ( .A(n5467), .B(\buff_mem[5][11] ), .X(n4753) );
  nand_x1_sg U6732 ( .A(n5468), .B(\buff_mem[5][14] ), .X(n4636) );
  nand_x1_sg U6733 ( .A(n5470), .B(\buff_mem[5][17] ), .X(n4519) );
  nor_x1_sg U6734 ( .A(n5832), .B(rd_ptr[0]), .X(n5184) );
  nor_x1_sg U6735 ( .A(n3499), .B(n5343), .X(n3500) );
  nand_x1_sg U6736 ( .A(wr_ptr[1]), .B(wr_ptr[0]), .X(n3474) );
  nand_x1_sg U6737 ( .A(n5342), .B(n3361), .X(n3484) );
  nand_x1_sg U6738 ( .A(wr_ptr[2]), .B(n5835), .X(n3479) );
  nor_x1_sg U6739 ( .A(n3484), .B(wr_ptr[4]), .X(n3482) );
  nor_x1_sg U6740 ( .A(n5826), .B(n3359), .X(n3483) );
  nand_x1_sg U6741 ( .A(n3462), .B(n5338), .X(n3461) );
  nand_x1_sg U6742 ( .A(n3358), .B(n5344), .X(n3460) );
  nand_x1_sg U6743 ( .A(n5346), .B(n3438), .X(n3436) );
  nand_x1_sg U6744 ( .A(full), .B(n3263), .X(n3437) );
  nand_x1_sg U6745 ( .A(\buff_mem[17][0] ), .B(n5477), .X(n5213) );
  nand_x1_sg U6746 ( .A(\buff_mem[17][1] ), .B(n5478), .X(n5166) );
  nand_x1_sg U6747 ( .A(\buff_mem[17][3] ), .B(n5477), .X(n5088) );
  nand_x1_sg U6748 ( .A(\buff_mem[17][4] ), .B(n5478), .X(n5049) );
  nand_x1_sg U6749 ( .A(\buff_mem[17][6] ), .B(n5482), .X(n4971) );
  nand_x1_sg U6750 ( .A(\buff_mem[17][7] ), .B(n5483), .X(n4932) );
  nand_x1_sg U6751 ( .A(\buff_mem[17][9] ), .B(n5482), .X(n4854) );
  nand_x1_sg U6752 ( .A(\buff_mem[17][10] ), .B(n5481), .X(n4815) );
  nand_x1_sg U6753 ( .A(\buff_mem[17][12] ), .B(n5479), .X(n4737) );
  nand_x1_sg U6754 ( .A(\buff_mem[17][13] ), .B(n5481), .X(n4698) );
  nand_x1_sg U6755 ( .A(\buff_mem[17][15] ), .B(n5483), .X(n4620) );
  nand_x1_sg U6756 ( .A(\buff_mem[17][16] ), .B(n5479), .X(n4581) );
  nand_x1_sg U6757 ( .A(\buff_mem[17][18] ), .B(n5479), .X(n4503) );
  nand_x1_sg U6758 ( .A(\buff_mem[17][19] ), .B(n5481), .X(n4463) );
  nor_x1_sg U6759 ( .A(n3336), .B(n5212), .X(n5210) );
  nor_x1_sg U6760 ( .A(n3414), .B(n5539), .X(n5212) );
  inv_x1_sg U6761 ( .A(\buff_mem[18][0] ), .X(n3414) );
  nor_x1_sg U6762 ( .A(n3337), .B(n5165), .X(n5163) );
  nor_x1_sg U6763 ( .A(n3411), .B(n5545), .X(n5165) );
  inv_x1_sg U6764 ( .A(\buff_mem[18][1] ), .X(n3411) );
  nor_x1_sg U6765 ( .A(n3339), .B(n5087), .X(n5085) );
  nor_x1_sg U6766 ( .A(n3405), .B(n5543), .X(n5087) );
  inv_x1_sg U6767 ( .A(\buff_mem[18][3] ), .X(n3405) );
  nor_x1_sg U6768 ( .A(n3340), .B(n5048), .X(n5046) );
  nor_x1_sg U6769 ( .A(n3402), .B(n5544), .X(n5048) );
  inv_x1_sg U6770 ( .A(\buff_mem[18][4] ), .X(n3402) );
  nor_x1_sg U6771 ( .A(n3342), .B(n4970), .X(n4968) );
  nor_x1_sg U6772 ( .A(n3396), .B(n5542), .X(n4970) );
  inv_x1_sg U6773 ( .A(\buff_mem[18][6] ), .X(n3396) );
  nor_x1_sg U6774 ( .A(n3343), .B(n4931), .X(n4929) );
  nor_x1_sg U6775 ( .A(n3393), .B(n5543), .X(n4931) );
  inv_x1_sg U6776 ( .A(\buff_mem[18][7] ), .X(n3393) );
  nor_x1_sg U6777 ( .A(n3345), .B(n4853), .X(n4851) );
  nor_x1_sg U6778 ( .A(n3387), .B(n5543), .X(n4853) );
  inv_x1_sg U6779 ( .A(\buff_mem[18][9] ), .X(n3387) );
  nor_x1_sg U6780 ( .A(n3346), .B(n4814), .X(n4812) );
  nor_x1_sg U6781 ( .A(n3384), .B(n5545), .X(n4814) );
  inv_x1_sg U6782 ( .A(\buff_mem[18][10] ), .X(n3384) );
  nor_x1_sg U6783 ( .A(n3348), .B(n4736), .X(n4734) );
  nor_x1_sg U6784 ( .A(n3378), .B(n5545), .X(n4736) );
  inv_x1_sg U6785 ( .A(\buff_mem[18][12] ), .X(n3378) );
  nor_x1_sg U6786 ( .A(n3349), .B(n4697), .X(n4695) );
  nor_x1_sg U6787 ( .A(n3375), .B(n5539), .X(n4697) );
  inv_x1_sg U6788 ( .A(\buff_mem[18][13] ), .X(n3375) );
  nor_x1_sg U6789 ( .A(n3351), .B(n4619), .X(n4617) );
  nor_x1_sg U6790 ( .A(n3429), .B(n5542), .X(n4619) );
  inv_x1_sg U6791 ( .A(\buff_mem[18][15] ), .X(n3429) );
  nor_x1_sg U6792 ( .A(n3352), .B(n4580), .X(n4578) );
  nor_x1_sg U6793 ( .A(n3426), .B(n5543), .X(n4580) );
  inv_x1_sg U6794 ( .A(\buff_mem[18][16] ), .X(n3426) );
  nor_x1_sg U6795 ( .A(n3354), .B(n4502), .X(n4500) );
  nor_x1_sg U6796 ( .A(n3420), .B(n5539), .X(n4502) );
  inv_x1_sg U6797 ( .A(\buff_mem[18][18] ), .X(n3420) );
  nor_x1_sg U6798 ( .A(n3355), .B(n4461), .X(n4458) );
  nor_x1_sg U6799 ( .A(n3417), .B(n5545), .X(n4461) );
  inv_x1_sg U6800 ( .A(\buff_mem[18][19] ), .X(n3417) );
  nand_x1_sg U6801 ( .A(n5315), .B(n5913), .X(n4397) );
  nand_x1_sg U6802 ( .A(n5906), .B(n3290), .X(n4398) );
  nand_x1_sg U6803 ( .A(\buff_mem[17][2] ), .B(n5478), .X(n5127) );
  nand_x1_sg U6804 ( .A(\buff_mem[17][5] ), .B(n5477), .X(n5010) );
  nand_x1_sg U6805 ( .A(\buff_mem[17][8] ), .B(n5482), .X(n4893) );
  nand_x1_sg U6806 ( .A(\buff_mem[17][11] ), .B(n5477), .X(n4776) );
  nand_x1_sg U6807 ( .A(\buff_mem[17][14] ), .B(n5478), .X(n4659) );
  nand_x1_sg U6808 ( .A(\buff_mem[17][17] ), .B(n5483), .X(n4542) );
  nor_x1_sg U6809 ( .A(n3338), .B(n5126), .X(n5124) );
  nor_x1_sg U6810 ( .A(n3408), .B(n5542), .X(n5126) );
  inv_x1_sg U6811 ( .A(\buff_mem[18][2] ), .X(n3408) );
  nor_x1_sg U6812 ( .A(n3341), .B(n5009), .X(n5007) );
  nor_x1_sg U6813 ( .A(n3399), .B(n5544), .X(n5009) );
  inv_x1_sg U6814 ( .A(\buff_mem[18][5] ), .X(n3399) );
  nor_x1_sg U6815 ( .A(n3344), .B(n4892), .X(n4890) );
  nor_x1_sg U6816 ( .A(n3390), .B(n5542), .X(n4892) );
  inv_x1_sg U6817 ( .A(\buff_mem[18][8] ), .X(n3390) );
  nor_x1_sg U6818 ( .A(n3347), .B(n4775), .X(n4773) );
  nor_x1_sg U6819 ( .A(n3381), .B(n5544), .X(n4775) );
  inv_x1_sg U6820 ( .A(\buff_mem[18][11] ), .X(n3381) );
  nor_x1_sg U6821 ( .A(n3350), .B(n4658), .X(n4656) );
  nor_x1_sg U6822 ( .A(n3432), .B(n5539), .X(n4658) );
  inv_x1_sg U6823 ( .A(\buff_mem[18][14] ), .X(n3432) );
  nor_x1_sg U6824 ( .A(n3353), .B(n4541), .X(n4539) );
  nor_x1_sg U6825 ( .A(n3423), .B(n5544), .X(n4541) );
  inv_x1_sg U6826 ( .A(\buff_mem[18][17] ), .X(n3423) );
  nand_x1_sg U6827 ( .A(n5498), .B(\buff_mem[11][0] ), .X(n5200) );
  nand_x1_sg U6828 ( .A(n5495), .B(\buff_mem[11][1] ), .X(n5154) );
  nand_x1_sg U6829 ( .A(n5498), .B(\buff_mem[11][3] ), .X(n5076) );
  nand_x1_sg U6830 ( .A(n5498), .B(\buff_mem[11][4] ), .X(n5037) );
  nand_x1_sg U6831 ( .A(n5496), .B(\buff_mem[11][6] ), .X(n4959) );
  nand_x1_sg U6832 ( .A(n5272), .B(\buff_mem[11][7] ), .X(n4920) );
  nand_x1_sg U6833 ( .A(n5495), .B(\buff_mem[11][9] ), .X(n4842) );
  nand_x1_sg U6834 ( .A(n5272), .B(\buff_mem[11][10] ), .X(n4803) );
  nand_x1_sg U6835 ( .A(n5496), .B(\buff_mem[11][12] ), .X(n4725) );
  nand_x1_sg U6836 ( .A(n5497), .B(\buff_mem[11][13] ), .X(n4686) );
  nand_x1_sg U6837 ( .A(n5496), .B(\buff_mem[11][15] ), .X(n4608) );
  nand_x1_sg U6838 ( .A(n5272), .B(\buff_mem[11][16] ), .X(n4569) );
  nand_x1_sg U6839 ( .A(n5497), .B(\buff_mem[11][18] ), .X(n4491) );
  nand_x1_sg U6840 ( .A(n5272), .B(\buff_mem[11][19] ), .X(n4443) );
  nand_x1_sg U6841 ( .A(\buff_mem[12][0] ), .B(n5270), .X(n5204) );
  nand_x1_sg U6842 ( .A(\buff_mem[13][0] ), .B(n5486), .X(n5205) );
  nand_x1_sg U6843 ( .A(\buff_mem[12][1] ), .B(n5490), .X(n5157) );
  nand_x1_sg U6844 ( .A(\buff_mem[13][1] ), .B(n5268), .X(n5158) );
  nand_x1_sg U6845 ( .A(\buff_mem[12][3] ), .B(n5491), .X(n5079) );
  nand_x1_sg U6846 ( .A(\buff_mem[13][3] ), .B(n5485), .X(n5080) );
  nand_x1_sg U6847 ( .A(\buff_mem[12][4] ), .B(n5492), .X(n5040) );
  nand_x1_sg U6848 ( .A(\buff_mem[13][4] ), .B(n5486), .X(n5041) );
  nand_x1_sg U6849 ( .A(\buff_mem[12][6] ), .B(n5270), .X(n4962) );
  nand_x1_sg U6850 ( .A(\buff_mem[13][6] ), .B(n5268), .X(n4963) );
  nand_x1_sg U6851 ( .A(\buff_mem[12][7] ), .B(n5492), .X(n4923) );
  nand_x1_sg U6852 ( .A(\buff_mem[13][7] ), .B(n5485), .X(n4924) );
  nand_x1_sg U6853 ( .A(\buff_mem[12][9] ), .B(n5270), .X(n4845) );
  nand_x1_sg U6854 ( .A(\buff_mem[13][9] ), .B(n5268), .X(n4846) );
  nand_x1_sg U6855 ( .A(\buff_mem[12][10] ), .B(n5490), .X(n4806) );
  nand_x1_sg U6856 ( .A(\buff_mem[13][10] ), .B(n5268), .X(n4807) );
  nand_x1_sg U6857 ( .A(\buff_mem[12][12] ), .B(n5491), .X(n4728) );
  nand_x1_sg U6858 ( .A(\buff_mem[13][12] ), .B(n5487), .X(n4729) );
  nand_x1_sg U6859 ( .A(\buff_mem[12][13] ), .B(n5270), .X(n4689) );
  nand_x1_sg U6860 ( .A(\buff_mem[13][13] ), .B(n5488), .X(n4690) );
  nand_x1_sg U6861 ( .A(\buff_mem[12][15] ), .B(n5490), .X(n4611) );
  nand_x1_sg U6862 ( .A(\buff_mem[13][15] ), .B(n5486), .X(n4612) );
  nand_x1_sg U6863 ( .A(\buff_mem[12][16] ), .B(n5491), .X(n4572) );
  nand_x1_sg U6864 ( .A(\buff_mem[13][16] ), .B(n5488), .X(n4573) );
  nand_x1_sg U6865 ( .A(\buff_mem[12][18] ), .B(n5490), .X(n4494) );
  nand_x1_sg U6866 ( .A(\buff_mem[13][18] ), .B(n5486), .X(n4495) );
  nand_x1_sg U6867 ( .A(\buff_mem[12][19] ), .B(n5493), .X(n4449) );
  nand_x1_sg U6868 ( .A(\buff_mem[13][19] ), .B(n5487), .X(n4450) );
  nand_x1_sg U6869 ( .A(n5507), .B(\buff_mem[9][0] ), .X(n5190) );
  nand_x1_sg U6870 ( .A(n5506), .B(\buff_mem[9][1] ), .X(n5145) );
  nand_x1_sg U6871 ( .A(n5505), .B(\buff_mem[9][3] ), .X(n5067) );
  nand_x1_sg U6872 ( .A(n5508), .B(\buff_mem[9][4] ), .X(n5028) );
  nand_x1_sg U6873 ( .A(n5276), .B(\buff_mem[9][6] ), .X(n4950) );
  nand_x1_sg U6874 ( .A(n5276), .B(\buff_mem[9][7] ), .X(n4911) );
  nand_x1_sg U6875 ( .A(n5507), .B(\buff_mem[9][9] ), .X(n4833) );
  nand_x1_sg U6876 ( .A(n5506), .B(\buff_mem[9][10] ), .X(n4794) );
  nand_x1_sg U6877 ( .A(n5505), .B(\buff_mem[9][12] ), .X(n4716) );
  nand_x1_sg U6878 ( .A(n5507), .B(\buff_mem[9][13] ), .X(n4677) );
  nand_x1_sg U6879 ( .A(n5506), .B(\buff_mem[9][15] ), .X(n4599) );
  nand_x1_sg U6880 ( .A(n5508), .B(\buff_mem[9][16] ), .X(n4560) );
  nand_x1_sg U6881 ( .A(n5508), .B(\buff_mem[9][18] ), .X(n4482) );
  nand_x1_sg U6882 ( .A(n5505), .B(\buff_mem[9][19] ), .X(n4432) );
  nand_x1_sg U6883 ( .A(rd_ptr[2]), .B(rd_ptr[3]), .X(n5202) );
  nand_x1_sg U6884 ( .A(n5391), .B(\buff_mem[10][0] ), .X(n5199) );
  nand_x1_sg U6885 ( .A(n5390), .B(\buff_mem[10][1] ), .X(n5153) );
  nand_x1_sg U6886 ( .A(n5238), .B(\buff_mem[10][3] ), .X(n5075) );
  nand_x1_sg U6887 ( .A(n5391), .B(\buff_mem[10][4] ), .X(n5036) );
  nand_x1_sg U6888 ( .A(n5391), .B(\buff_mem[10][6] ), .X(n4958) );
  nand_x1_sg U6889 ( .A(n5388), .B(\buff_mem[10][7] ), .X(n4919) );
  nand_x1_sg U6890 ( .A(n5389), .B(\buff_mem[10][9] ), .X(n4841) );
  nand_x1_sg U6891 ( .A(n5388), .B(\buff_mem[10][10] ), .X(n4802) );
  nand_x1_sg U6892 ( .A(n5390), .B(\buff_mem[10][12] ), .X(n4724) );
  nand_x1_sg U6893 ( .A(n5389), .B(\buff_mem[10][13] ), .X(n4685) );
  nand_x1_sg U6894 ( .A(n5238), .B(\buff_mem[10][15] ), .X(n4607) );
  nand_x1_sg U6895 ( .A(n5388), .B(\buff_mem[10][16] ), .X(n4568) );
  nand_x1_sg U6896 ( .A(n5238), .B(\buff_mem[10][18] ), .X(n4490) );
  nand_x1_sg U6897 ( .A(n5389), .B(\buff_mem[10][19] ), .X(n4442) );
  nand_x1_sg U6898 ( .A(n5497), .B(\buff_mem[11][2] ), .X(n5115) );
  nand_x1_sg U6899 ( .A(n5498), .B(\buff_mem[11][5] ), .X(n4998) );
  nand_x1_sg U6900 ( .A(n5495), .B(\buff_mem[11][8] ), .X(n4881) );
  nand_x1_sg U6901 ( .A(n5495), .B(\buff_mem[11][11] ), .X(n4764) );
  nand_x1_sg U6902 ( .A(n5496), .B(\buff_mem[11][14] ), .X(n4647) );
  nand_x1_sg U6903 ( .A(n5497), .B(\buff_mem[11][17] ), .X(n4530) );
  nand_x1_sg U6904 ( .A(\buff_mem[12][2] ), .B(n5491), .X(n5118) );
  nand_x1_sg U6905 ( .A(\buff_mem[13][2] ), .B(n5487), .X(n5119) );
  nand_x1_sg U6906 ( .A(\buff_mem[12][5] ), .B(n5493), .X(n5001) );
  nand_x1_sg U6907 ( .A(\buff_mem[13][5] ), .B(n5487), .X(n5002) );
  nand_x1_sg U6908 ( .A(\buff_mem[12][8] ), .B(n5492), .X(n4884) );
  nand_x1_sg U6909 ( .A(\buff_mem[13][8] ), .B(n5485), .X(n4885) );
  nand_x1_sg U6910 ( .A(\buff_mem[12][11] ), .B(n5493), .X(n4767) );
  nand_x1_sg U6911 ( .A(\buff_mem[13][11] ), .B(n5488), .X(n4768) );
  nand_x1_sg U6912 ( .A(\buff_mem[12][14] ), .B(n5492), .X(n4650) );
  nand_x1_sg U6913 ( .A(\buff_mem[13][14] ), .B(n5488), .X(n4651) );
  nand_x1_sg U6914 ( .A(\buff_mem[12][17] ), .B(n5493), .X(n4533) );
  nand_x1_sg U6915 ( .A(\buff_mem[13][17] ), .B(n5485), .X(n4534) );
  nand_x1_sg U6916 ( .A(n5276), .B(\buff_mem[9][2] ), .X(n5106) );
  nand_x1_sg U6917 ( .A(n5505), .B(\buff_mem[9][5] ), .X(n4989) );
  nand_x1_sg U6918 ( .A(n5506), .B(\buff_mem[9][8] ), .X(n4872) );
  nand_x1_sg U6919 ( .A(n5276), .B(\buff_mem[9][11] ), .X(n4755) );
  nand_x1_sg U6920 ( .A(n5508), .B(\buff_mem[9][14] ), .X(n4638) );
  nand_x1_sg U6921 ( .A(n5507), .B(\buff_mem[9][17] ), .X(n4521) );
  nand_x1_sg U6922 ( .A(n5390), .B(\buff_mem[10][2] ), .X(n5114) );
  nand_x1_sg U6923 ( .A(n5391), .B(\buff_mem[10][5] ), .X(n4997) );
  nand_x1_sg U6924 ( .A(n5390), .B(\buff_mem[10][8] ), .X(n4880) );
  nand_x1_sg U6925 ( .A(n5389), .B(\buff_mem[10][11] ), .X(n4763) );
  nand_x1_sg U6926 ( .A(n5238), .B(\buff_mem[10][14] ), .X(n4646) );
  nand_x1_sg U6927 ( .A(n5388), .B(\buff_mem[10][17] ), .X(n4529) );
  nand_x1_sg U6928 ( .A(n5513), .B(\buff_mem[14][0] ), .X(n5201) );
  nand_x1_sg U6929 ( .A(n5510), .B(\buff_mem[14][1] ), .X(n5155) );
  nand_x1_sg U6930 ( .A(n5510), .B(\buff_mem[14][3] ), .X(n5077) );
  nand_x1_sg U6931 ( .A(n5513), .B(\buff_mem[14][4] ), .X(n5038) );
  nand_x1_sg U6932 ( .A(n5511), .B(\buff_mem[14][6] ), .X(n4960) );
  nand_x1_sg U6933 ( .A(n5511), .B(\buff_mem[14][7] ), .X(n4921) );
  nand_x1_sg U6934 ( .A(n5510), .B(\buff_mem[14][9] ), .X(n4843) );
  nand_x1_sg U6935 ( .A(n5278), .B(\buff_mem[14][10] ), .X(n4804) );
  nand_x1_sg U6936 ( .A(n5513), .B(\buff_mem[14][12] ), .X(n4726) );
  nand_x1_sg U6937 ( .A(n5511), .B(\buff_mem[14][13] ), .X(n4687) );
  nand_x1_sg U6938 ( .A(n5512), .B(\buff_mem[14][15] ), .X(n4609) );
  nand_x1_sg U6939 ( .A(n5278), .B(\buff_mem[14][16] ), .X(n4570) );
  nand_x1_sg U6940 ( .A(n5512), .B(\buff_mem[14][18] ), .X(n4492) );
  nand_x1_sg U6941 ( .A(n5278), .B(\buff_mem[14][19] ), .X(n4446) );
  nand_x1_sg U6942 ( .A(n5513), .B(\buff_mem[14][2] ), .X(n5116) );
  nand_x1_sg U6943 ( .A(n5510), .B(\buff_mem[14][5] ), .X(n4999) );
  nand_x1_sg U6944 ( .A(n5512), .B(\buff_mem[14][8] ), .X(n4882) );
  nand_x1_sg U6945 ( .A(n5512), .B(\buff_mem[14][11] ), .X(n4765) );
  nand_x1_sg U6946 ( .A(n5278), .B(\buff_mem[14][14] ), .X(n4648) );
  nand_x1_sg U6947 ( .A(n5511), .B(\buff_mem[14][17] ), .X(n4531) );
  nand_x1_sg U6948 ( .A(n5342), .B(n3479), .X(n3478) );
  nand_x1_sg U6949 ( .A(n3361), .B(n3366), .X(n3477) );
  nor_x1_sg U6950 ( .A(n3457), .B(n3458), .X(n3452) );
  nor_x1_sg U6951 ( .A(n3454), .B(n3360), .X(n3453) );
  nor_x1_sg U6952 ( .A(n5340), .B(n3459), .X(n3458) );
  nor_x1_sg U6953 ( .A(n3474), .B(n5325), .X(n3472) );
  nor_x1_sg U6954 ( .A(n5915), .B(n5835), .X(n3473) );
  nand_x1_sg U6955 ( .A(n5517), .B(\buff_mem[16][0] ), .X(n5208) );
  nand_x1_sg U6956 ( .A(n5518), .B(\buff_mem[16][1] ), .X(n5161) );
  nand_x1_sg U6957 ( .A(n5517), .B(\buff_mem[16][3] ), .X(n5083) );
  nand_x1_sg U6958 ( .A(n5280), .B(\buff_mem[16][4] ), .X(n5044) );
  nand_x1_sg U6959 ( .A(n5517), .B(\buff_mem[16][6] ), .X(n4966) );
  nand_x1_sg U6960 ( .A(n5518), .B(\buff_mem[16][7] ), .X(n4927) );
  nand_x1_sg U6961 ( .A(n5518), .B(\buff_mem[16][9] ), .X(n4849) );
  nand_x1_sg U6962 ( .A(n5515), .B(\buff_mem[16][10] ), .X(n4810) );
  nand_x1_sg U6963 ( .A(n5280), .B(\buff_mem[16][12] ), .X(n4732) );
  nand_x1_sg U6964 ( .A(n5517), .B(\buff_mem[16][13] ), .X(n4693) );
  nand_x1_sg U6965 ( .A(n5515), .B(\buff_mem[16][15] ), .X(n4615) );
  nand_x1_sg U6966 ( .A(n5516), .B(\buff_mem[16][16] ), .X(n4576) );
  nand_x1_sg U6967 ( .A(n5516), .B(\buff_mem[16][18] ), .X(n4498) );
  nand_x1_sg U6968 ( .A(n5516), .B(\buff_mem[16][19] ), .X(n4455) );
  nand_x1_sg U6969 ( .A(n5280), .B(\buff_mem[16][2] ), .X(n5122) );
  nand_x1_sg U6970 ( .A(n5518), .B(\buff_mem[16][5] ), .X(n5005) );
  nand_x1_sg U6971 ( .A(n5280), .B(\buff_mem[16][8] ), .X(n4888) );
  nand_x1_sg U6972 ( .A(n5516), .B(\buff_mem[16][11] ), .X(n4771) );
  nand_x1_sg U6973 ( .A(n5515), .B(\buff_mem[16][14] ), .X(n4654) );
  nand_x1_sg U6974 ( .A(n5515), .B(\buff_mem[16][17] ), .X(n4537) );
  nor_x1_sg U6975 ( .A(n5823), .B(wr_ptr[4]), .X(n3705) );
  nor_x1_sg U6976 ( .A(empty), .B(n3286), .X(n4388) );
  nand_x1_sg U6977 ( .A(n3448), .B(n3449), .X(n3442) );
  nand_x1_sg U6978 ( .A(n5222), .B(n3359), .X(n3449) );
  nor_x1_sg U6979 ( .A(wr_ptr[3]), .B(n5915), .X(n3875) );
  nand_x1_sg U6980 ( .A(n4045), .B(n3705), .X(n4044) );
  nor_x1_sg U6981 ( .A(n5325), .B(n3366), .X(n4045) );
  nand_x1_sg U6982 ( .A(\buff_mem[4][14] ), .B(n5634), .X(n3736) );
  nand_x1_sg U6983 ( .A(\buff_mem[10][14] ), .B(n5641), .X(n3990) );
  nand_x1_sg U6984 ( .A(\buff_mem[12][14] ), .B(n5597), .X(n4076) );
  nand_x1_sg U6985 ( .A(\buff_mem[13][14] ), .B(n5590), .X(n4118) );
  nand_x1_sg U6986 ( .A(n5256), .B(n5800), .X(n3737) );
  nand_x1_sg U6987 ( .A(\buff_mem[4][15] ), .B(n5637), .X(n3738) );
  nand_x1_sg U6988 ( .A(n5368), .B(n5802), .X(n3739) );
  nand_x1_sg U6989 ( .A(\buff_mem[4][16] ), .B(n5307), .X(n3740) );
  nand_x1_sg U6990 ( .A(n5436), .B(n5799), .X(n3741) );
  nand_x1_sg U6991 ( .A(\buff_mem[4][17] ), .B(n5637), .X(n3742) );
  nand_x1_sg U6992 ( .A(n5244), .B(n5799), .X(n3743) );
  nand_x1_sg U6993 ( .A(\buff_mem[4][18] ), .B(n5634), .X(n3744) );
  nand_x1_sg U6994 ( .A(n5379), .B(n5799), .X(n3745) );
  nand_x1_sg U6995 ( .A(\buff_mem[4][19] ), .B(n5307), .X(n3746) );
  nand_x1_sg U6996 ( .A(n5521), .B(n5793), .X(n3706) );
  nand_x1_sg U6997 ( .A(\buff_mem[4][0] ), .B(n5635), .X(n3707) );
  nand_x1_sg U6998 ( .A(n5526), .B(n5796), .X(n3709) );
  nand_x1_sg U6999 ( .A(\buff_mem[4][1] ), .B(n5636), .X(n3710) );
  nand_x1_sg U7000 ( .A(n5393), .B(n5800), .X(n3711) );
  nand_x1_sg U7001 ( .A(\buff_mem[4][2] ), .B(n5634), .X(n3712) );
  nand_x1_sg U7002 ( .A(n5531), .B(n5799), .X(n3713) );
  nand_x1_sg U7003 ( .A(\buff_mem[4][3] ), .B(n5636), .X(n3714) );
  nand_x1_sg U7004 ( .A(n5358), .B(n5793), .X(n3715) );
  nand_x1_sg U7005 ( .A(\buff_mem[4][4] ), .B(n5636), .X(n3716) );
  nand_x1_sg U7006 ( .A(n5430), .B(n5795), .X(n3717) );
  nand_x1_sg U7007 ( .A(\buff_mem[4][5] ), .B(n5635), .X(n3718) );
  nand_x1_sg U7008 ( .A(n5400), .B(n5801), .X(n3719) );
  nand_x1_sg U7009 ( .A(\buff_mem[4][6] ), .B(n5637), .X(n3720) );
  nand_x1_sg U7010 ( .A(n5425), .B(n5800), .X(n3721) );
  nand_x1_sg U7011 ( .A(\buff_mem[4][7] ), .B(n5634), .X(n3722) );
  nand_x1_sg U7012 ( .A(n5373), .B(n5794), .X(n3723) );
  nand_x1_sg U7013 ( .A(\buff_mem[4][8] ), .B(n5307), .X(n3724) );
  nand_x1_sg U7014 ( .A(n5650), .B(n5800), .X(n3725) );
  nand_x1_sg U7015 ( .A(\buff_mem[4][9] ), .B(n5637), .X(n3726) );
  nand_x1_sg U7016 ( .A(n5644), .B(n5802), .X(n3727) );
  nand_x1_sg U7017 ( .A(\buff_mem[4][10] ), .B(n5635), .X(n3728) );
  nand_x1_sg U7018 ( .A(n5288), .B(n5793), .X(n3729) );
  nand_x1_sg U7019 ( .A(\buff_mem[4][11] ), .B(n5635), .X(n3730) );
  nand_x1_sg U7020 ( .A(n5365), .B(n5796), .X(n3731) );
  nand_x1_sg U7021 ( .A(\buff_mem[4][12] ), .B(n5636), .X(n3732) );
  nand_x1_sg U7022 ( .A(n5421), .B(n5794), .X(n3733) );
  nand_x1_sg U7023 ( .A(\buff_mem[4][13] ), .B(n5307), .X(n3734) );
  nand_x1_sg U7024 ( .A(n5522), .B(n5770), .X(n4046) );
  nand_x1_sg U7025 ( .A(\buff_mem[12][0] ), .B(n5299), .X(n4047) );
  nand_x1_sg U7026 ( .A(n5528), .B(n5778), .X(n4049) );
  nand_x1_sg U7027 ( .A(\buff_mem[12][1] ), .B(n5597), .X(n4050) );
  nand_x1_sg U7028 ( .A(n5393), .B(n5776), .X(n4051) );
  nand_x1_sg U7029 ( .A(\buff_mem[12][2] ), .B(n5596), .X(n4052) );
  nand_x1_sg U7030 ( .A(n5533), .B(n5776), .X(n4053) );
  nand_x1_sg U7031 ( .A(\buff_mem[12][3] ), .B(n5595), .X(n4054) );
  nand_x1_sg U7032 ( .A(n5361), .B(n5772), .X(n4055) );
  nand_x1_sg U7033 ( .A(\buff_mem[12][4] ), .B(n5597), .X(n4056) );
  nand_x1_sg U7034 ( .A(n5430), .B(n5776), .X(n4057) );
  nand_x1_sg U7035 ( .A(\buff_mem[12][5] ), .B(n5598), .X(n4058) );
  nand_x1_sg U7036 ( .A(n5398), .B(n5770), .X(n4059) );
  nand_x1_sg U7037 ( .A(\buff_mem[12][6] ), .B(n5595), .X(n4060) );
  nand_x1_sg U7038 ( .A(n5425), .B(n5779), .X(n4061) );
  nand_x1_sg U7039 ( .A(\buff_mem[12][7] ), .B(n5598), .X(n4062) );
  nand_x1_sg U7040 ( .A(n5373), .B(n5771), .X(n4063) );
  nand_x1_sg U7041 ( .A(\buff_mem[12][8] ), .B(n5595), .X(n4064) );
  nand_x1_sg U7042 ( .A(n5651), .B(n5776), .X(n4065) );
  nand_x1_sg U7043 ( .A(\buff_mem[12][9] ), .B(n5598), .X(n4066) );
  nand_x1_sg U7044 ( .A(n5645), .B(n5778), .X(n4067) );
  nand_x1_sg U7045 ( .A(\buff_mem[12][10] ), .B(n5596), .X(n4068) );
  nand_x1_sg U7046 ( .A(n5536), .B(n5770), .X(n4069) );
  nand_x1_sg U7047 ( .A(\buff_mem[12][11] ), .B(n5598), .X(n4070) );
  nand_x1_sg U7048 ( .A(n5363), .B(n5773), .X(n4071) );
  nand_x1_sg U7049 ( .A(\buff_mem[12][12] ), .B(n5299), .X(n4072) );
  nand_x1_sg U7050 ( .A(n5423), .B(n5773), .X(n4073) );
  nand_x1_sg U7051 ( .A(\buff_mem[12][13] ), .B(n5595), .X(n4074) );
  nand_x1_sg U7052 ( .A(n5256), .B(n5777), .X(n4077) );
  nand_x1_sg U7053 ( .A(\buff_mem[12][15] ), .B(n5299), .X(n4078) );
  nand_x1_sg U7054 ( .A(n5370), .B(n5779), .X(n4079) );
  nand_x1_sg U7055 ( .A(\buff_mem[12][16] ), .B(n5597), .X(n4080) );
  nand_x1_sg U7056 ( .A(n5254), .B(n5771), .X(n4081) );
  nand_x1_sg U7057 ( .A(\buff_mem[12][17] ), .B(n5596), .X(n4082) );
  nand_x1_sg U7058 ( .A(n5405), .B(n5777), .X(n4083) );
  nand_x1_sg U7059 ( .A(\buff_mem[12][18] ), .B(n5596), .X(n4084) );
  nand_x1_sg U7060 ( .A(n5380), .B(n5777), .X(n4085) );
  nand_x1_sg U7061 ( .A(\buff_mem[12][19] ), .B(n5299), .X(n4086) );
  nand_x1_sg U7062 ( .A(n5522), .B(n5661), .X(n4088) );
  nand_x1_sg U7063 ( .A(\buff_mem[13][0] ), .B(n5593), .X(n4089) );
  nand_x1_sg U7064 ( .A(n5527), .B(n5658), .X(n4091) );
  nand_x1_sg U7065 ( .A(\buff_mem[13][1] ), .B(n5590), .X(n4092) );
  nand_x1_sg U7066 ( .A(n5240), .B(n5658), .X(n4093) );
  nand_x1_sg U7067 ( .A(\buff_mem[13][2] ), .B(n5593), .X(n4094) );
  nand_x1_sg U7068 ( .A(n5530), .B(n5655), .X(n4095) );
  nand_x1_sg U7069 ( .A(\buff_mem[13][3] ), .B(n5591), .X(n4096) );
  nand_x1_sg U7070 ( .A(n5226), .B(n5654), .X(n4097) );
  nand_x1_sg U7071 ( .A(\buff_mem[13][4] ), .B(n5298), .X(n4098) );
  nand_x1_sg U7072 ( .A(n5252), .B(n5662), .X(n4099) );
  nand_x1_sg U7073 ( .A(\buff_mem[13][5] ), .B(n5591), .X(n4100) );
  nand_x1_sg U7074 ( .A(n5401), .B(n5661), .X(n4101) );
  nand_x1_sg U7075 ( .A(\buff_mem[13][6] ), .B(n5590), .X(n4102) );
  nand_x1_sg U7076 ( .A(n5250), .B(n5656), .X(n4103) );
  nand_x1_sg U7077 ( .A(\buff_mem[13][7] ), .B(n5591), .X(n4104) );
  nand_x1_sg U7078 ( .A(n5376), .B(n5659), .X(n4105) );
  nand_x1_sg U7079 ( .A(\buff_mem[13][8] ), .B(n5590), .X(n4106) );
  nand_x1_sg U7080 ( .A(n5649), .B(n5662), .X(n4107) );
  nand_x1_sg U7081 ( .A(\buff_mem[13][9] ), .B(n5593), .X(n4108) );
  nand_x1_sg U7082 ( .A(n5310), .B(n5662), .X(n4109) );
  nand_x1_sg U7083 ( .A(\buff_mem[13][10] ), .B(n5593), .X(n4110) );
  nand_x1_sg U7084 ( .A(n5288), .B(n5654), .X(n4111) );
  nand_x1_sg U7085 ( .A(\buff_mem[13][11] ), .B(n5592), .X(n4112) );
  nand_x1_sg U7086 ( .A(n5364), .B(n5655), .X(n4113) );
  nand_x1_sg U7087 ( .A(\buff_mem[13][12] ), .B(n5298), .X(n4114) );
  nand_x1_sg U7088 ( .A(n5420), .B(n5659), .X(n4115) );
  nand_x1_sg U7089 ( .A(\buff_mem[13][13] ), .B(n5591), .X(n4116) );
  nand_x1_sg U7090 ( .A(n5442), .B(n5656), .X(n4119) );
  nand_x1_sg U7091 ( .A(\buff_mem[13][15] ), .B(n5592), .X(n4120) );
  nand_x1_sg U7092 ( .A(n5371), .B(n5661), .X(n4121) );
  nand_x1_sg U7093 ( .A(\buff_mem[13][16] ), .B(n5298), .X(n4122) );
  nand_x1_sg U7094 ( .A(n5438), .B(n5656), .X(n4123) );
  nand_x1_sg U7095 ( .A(\buff_mem[13][17] ), .B(n5592), .X(n4124) );
  nand_x1_sg U7096 ( .A(n5406), .B(n5655), .X(n4125) );
  nand_x1_sg U7097 ( .A(\buff_mem[13][18] ), .B(n5592), .X(n4126) );
  nand_x1_sg U7098 ( .A(n5234), .B(n5659), .X(n4127) );
  nand_x1_sg U7099 ( .A(\buff_mem[13][19] ), .B(n5298), .X(n4128) );
  nand_x1_sg U7100 ( .A(n5440), .B(n5782), .X(n3991) );
  nand_x1_sg U7101 ( .A(\buff_mem[10][15] ), .B(n5640), .X(n3992) );
  nand_x1_sg U7102 ( .A(n5371), .B(n5787), .X(n3993) );
  nand_x1_sg U7103 ( .A(\buff_mem[10][16] ), .B(n5641), .X(n3994) );
  nand_x1_sg U7104 ( .A(n5254), .B(n5785), .X(n3995) );
  nand_x1_sg U7105 ( .A(\buff_mem[10][17] ), .B(n5640), .X(n3996) );
  nand_x1_sg U7106 ( .A(n5404), .B(n5782), .X(n3997) );
  nand_x1_sg U7107 ( .A(\buff_mem[10][18] ), .B(n5308), .X(n3998) );
  nand_x1_sg U7108 ( .A(n5378), .B(n5783), .X(n3999) );
  nand_x1_sg U7109 ( .A(\buff_mem[10][19] ), .B(n5641), .X(n4000) );
  nand_x1_sg U7110 ( .A(n5521), .B(n5787), .X(n3960) );
  nand_x1_sg U7111 ( .A(\buff_mem[10][0] ), .B(n5639), .X(n3961) );
  nand_x1_sg U7112 ( .A(n5525), .B(n5783), .X(n3963) );
  nand_x1_sg U7113 ( .A(\buff_mem[10][1] ), .B(n5641), .X(n3964) );
  nand_x1_sg U7114 ( .A(n5393), .B(n5787), .X(n3965) );
  nand_x1_sg U7115 ( .A(\buff_mem[10][2] ), .B(n5639), .X(n3966) );
  nand_x1_sg U7116 ( .A(n5532), .B(n5780), .X(n3967) );
  nand_x1_sg U7117 ( .A(\buff_mem[10][3] ), .B(n5640), .X(n3968) );
  nand_x1_sg U7118 ( .A(n5361), .B(n5785), .X(n3969) );
  nand_x1_sg U7119 ( .A(\buff_mem[10][4] ), .B(n5308), .X(n3970) );
  nand_x1_sg U7120 ( .A(n5430), .B(n5786), .X(n3971) );
  nand_x1_sg U7121 ( .A(\buff_mem[10][5] ), .B(n5640), .X(n3972) );
  nand_x1_sg U7122 ( .A(n5242), .B(n5785), .X(n3973) );
  nand_x1_sg U7123 ( .A(\buff_mem[10][6] ), .B(n5308), .X(n3974) );
  nand_x1_sg U7124 ( .A(n5427), .B(n5787), .X(n3975) );
  nand_x1_sg U7125 ( .A(\buff_mem[10][7] ), .B(n5639), .X(n3976) );
  nand_x1_sg U7126 ( .A(n5375), .B(n5782), .X(n3977) );
  nand_x1_sg U7127 ( .A(\buff_mem[10][8] ), .B(n5642), .X(n3978) );
  nand_x1_sg U7128 ( .A(n5312), .B(n5783), .X(n3979) );
  nand_x1_sg U7129 ( .A(\buff_mem[10][9] ), .B(n5642), .X(n3980) );
  nand_x1_sg U7130 ( .A(n5647), .B(n5786), .X(n3981) );
  nand_x1_sg U7131 ( .A(\buff_mem[10][10] ), .B(n5642), .X(n3982) );
  nand_x1_sg U7132 ( .A(n5535), .B(n5786), .X(n3983) );
  nand_x1_sg U7133 ( .A(\buff_mem[10][11] ), .B(n5639), .X(n3984) );
  nand_x1_sg U7134 ( .A(n5228), .B(n5786), .X(n3985) );
  nand_x1_sg U7135 ( .A(\buff_mem[10][12] ), .B(n5642), .X(n3986) );
  nand_x1_sg U7136 ( .A(n5248), .B(n5782), .X(n3987) );
  nand_x1_sg U7137 ( .A(\buff_mem[10][13] ), .B(n5308), .X(n3988) );
  nand_x1_sg U7138 ( .A(\buff_mem[3][14] ), .B(n5562), .X(n3691) );
  nand_x1_sg U7139 ( .A(n5441), .B(n5673), .X(n3692) );
  nand_x1_sg U7140 ( .A(\buff_mem[3][15] ), .B(n5562), .X(n3693) );
  nand_x1_sg U7141 ( .A(n5368), .B(n5674), .X(n3694) );
  nand_x1_sg U7142 ( .A(\buff_mem[3][16] ), .B(n5292), .X(n3695) );
  nand_x1_sg U7143 ( .A(n5435), .B(n5675), .X(n3696) );
  nand_x1_sg U7144 ( .A(\buff_mem[3][17] ), .B(n5563), .X(n3697) );
  nand_x1_sg U7145 ( .A(n5404), .B(n5671), .X(n3698) );
  nand_x1_sg U7146 ( .A(\buff_mem[3][18] ), .B(n5561), .X(n3699) );
  nand_x1_sg U7147 ( .A(n5381), .B(n5675), .X(n3700) );
  nand_x1_sg U7148 ( .A(\buff_mem[3][19] ), .B(n5292), .X(n3701) );
  nand_x1_sg U7149 ( .A(n5522), .B(n5675), .X(n3661) );
  nand_x1_sg U7150 ( .A(\buff_mem[3][0] ), .B(n5564), .X(n3662) );
  nand_x1_sg U7151 ( .A(n5527), .B(n5668), .X(n3664) );
  nand_x1_sg U7152 ( .A(\buff_mem[3][1] ), .B(n5563), .X(n3665) );
  nand_x1_sg U7153 ( .A(n5396), .B(n5670), .X(n3666) );
  nand_x1_sg U7154 ( .A(\buff_mem[3][2] ), .B(n5564), .X(n3667) );
  nand_x1_sg U7155 ( .A(n5286), .B(n5670), .X(n3668) );
  nand_x1_sg U7156 ( .A(\buff_mem[3][3] ), .B(n5562), .X(n3669) );
  nand_x1_sg U7157 ( .A(n5358), .B(n5674), .X(n3670) );
  nand_x1_sg U7158 ( .A(\buff_mem[3][4] ), .B(n5292), .X(n3671) );
  nand_x1_sg U7159 ( .A(n5432), .B(n5670), .X(n3672) );
  nand_x1_sg U7160 ( .A(\buff_mem[3][5] ), .B(n5562), .X(n3673) );
  nand_x1_sg U7161 ( .A(n5242), .B(n5674), .X(n3674) );
  nand_x1_sg U7162 ( .A(\buff_mem[3][6] ), .B(n5561), .X(n3675) );
  nand_x1_sg U7163 ( .A(n5426), .B(n5673), .X(n3676) );
  nand_x1_sg U7164 ( .A(\buff_mem[3][7] ), .B(n5563), .X(n3677) );
  nand_x1_sg U7165 ( .A(n5375), .B(n5675), .X(n3678) );
  nand_x1_sg U7166 ( .A(\buff_mem[3][8] ), .B(n5561), .X(n3679) );
  nand_x1_sg U7167 ( .A(n5651), .B(n5673), .X(n3680) );
  nand_x1_sg U7168 ( .A(\buff_mem[3][9] ), .B(n5564), .X(n3681) );
  nand_x1_sg U7169 ( .A(n5644), .B(n5673), .X(n3682) );
  nand_x1_sg U7170 ( .A(\buff_mem[3][10] ), .B(n5564), .X(n3683) );
  nand_x1_sg U7171 ( .A(n5537), .B(n5670), .X(n3684) );
  nand_x1_sg U7172 ( .A(\buff_mem[3][11] ), .B(n5561), .X(n3685) );
  nand_x1_sg U7173 ( .A(n5364), .B(n5671), .X(n3686) );
  nand_x1_sg U7174 ( .A(\buff_mem[3][12] ), .B(n5292), .X(n3687) );
  nand_x1_sg U7175 ( .A(n5422), .B(n5671), .X(n3688) );
  nand_x1_sg U7176 ( .A(\buff_mem[3][13] ), .B(n5563), .X(n3689) );
  nand_x1_sg U7177 ( .A(\buff_mem[5][14] ), .B(n5600), .X(n3778) );
  nand_x1_sg U7178 ( .A(n5410), .B(n5733), .X(n3819) );
  nand_x1_sg U7179 ( .A(\buff_mem[6][14] ), .B(n5557), .X(n3820) );
  nand_x1_sg U7180 ( .A(n5409), .B(n5709), .X(n3905) );
  nand_x1_sg U7181 ( .A(\buff_mem[8][14] ), .B(n5610), .X(n3906) );
  nand_x1_sg U7182 ( .A(n5408), .B(n5356), .X(n3947) );
  nand_x1_sg U7183 ( .A(\buff_mem[9][14] ), .B(n5548), .X(n3948) );
  nand_x1_sg U7184 ( .A(n5409), .B(n5715), .X(n4159) );
  nand_x1_sg U7185 ( .A(\buff_mem[14][14] ), .B(n5631), .X(n4160) );
  nand_x1_sg U7186 ( .A(n5523), .B(n5738), .X(n3748) );
  nand_x1_sg U7187 ( .A(\buff_mem[5][0] ), .B(n5601), .X(n3749) );
  nand_x1_sg U7188 ( .A(n5528), .B(n5737), .X(n3751) );
  nand_x1_sg U7189 ( .A(\buff_mem[5][1] ), .B(n5603), .X(n3752) );
  nand_x1_sg U7190 ( .A(n5240), .B(n5737), .X(n3753) );
  nand_x1_sg U7191 ( .A(\buff_mem[5][2] ), .B(n5601), .X(n3754) );
  nand_x1_sg U7192 ( .A(n5533), .B(n5737), .X(n3755) );
  nand_x1_sg U7193 ( .A(\buff_mem[5][3] ), .B(n5602), .X(n3756) );
  nand_x1_sg U7194 ( .A(n5358), .B(n5739), .X(n3757) );
  nand_x1_sg U7195 ( .A(\buff_mem[5][4] ), .B(n5602), .X(n3758) );
  nand_x1_sg U7196 ( .A(n5252), .B(n5331), .X(n3759) );
  nand_x1_sg U7197 ( .A(\buff_mem[5][5] ), .B(n5603), .X(n3760) );
  nand_x1_sg U7198 ( .A(n5401), .B(n5331), .X(n3761) );
  nand_x1_sg U7199 ( .A(\buff_mem[5][6] ), .B(n5600), .X(n3762) );
  nand_x1_sg U7200 ( .A(n5428), .B(n5739), .X(n3763) );
  nand_x1_sg U7201 ( .A(\buff_mem[5][7] ), .B(n5601), .X(n3764) );
  nand_x1_sg U7202 ( .A(n5373), .B(n5736), .X(n3765) );
  nand_x1_sg U7203 ( .A(\buff_mem[5][8] ), .B(n5300), .X(n3766) );
  nand_x1_sg U7204 ( .A(n5312), .B(n5739), .X(n3767) );
  nand_x1_sg U7205 ( .A(\buff_mem[5][9] ), .B(n5300), .X(n3768) );
  nand_x1_sg U7206 ( .A(n5647), .B(n5331), .X(n3769) );
  nand_x1_sg U7207 ( .A(\buff_mem[5][10] ), .B(n5300), .X(n3770) );
  nand_x1_sg U7208 ( .A(n5535), .B(n5738), .X(n3771) );
  nand_x1_sg U7209 ( .A(\buff_mem[5][11] ), .B(n5602), .X(n3772) );
  nand_x1_sg U7210 ( .A(n5366), .B(n5736), .X(n3773) );
  nand_x1_sg U7211 ( .A(\buff_mem[5][12] ), .B(n5300), .X(n3774) );
  nand_x1_sg U7212 ( .A(n5423), .B(n5738), .X(n3775) );
  nand_x1_sg U7213 ( .A(\buff_mem[5][13] ), .B(n5600), .X(n3776) );
  nand_x1_sg U7214 ( .A(n5443), .B(n5739), .X(n3779) );
  nand_x1_sg U7215 ( .A(\buff_mem[5][15] ), .B(n5603), .X(n3780) );
  nand_x1_sg U7216 ( .A(n5371), .B(n5736), .X(n3781) );
  nand_x1_sg U7217 ( .A(\buff_mem[5][16] ), .B(n5600), .X(n3782) );
  nand_x1_sg U7218 ( .A(n5436), .B(n5738), .X(n3783) );
  nand_x1_sg U7219 ( .A(\buff_mem[5][17] ), .B(n5601), .X(n3784) );
  nand_x1_sg U7220 ( .A(n5404), .B(n5737), .X(n3785) );
  nand_x1_sg U7221 ( .A(\buff_mem[5][18] ), .B(n5603), .X(n3786) );
  nand_x1_sg U7222 ( .A(n5378), .B(n5736), .X(n3787) );
  nand_x1_sg U7223 ( .A(\buff_mem[5][19] ), .B(n5602), .X(n3788) );
  nand_x1_sg U7224 ( .A(n5282), .B(n5734), .X(n3790) );
  nand_x1_sg U7225 ( .A(\buff_mem[6][0] ), .B(n5557), .X(n3791) );
  nand_x1_sg U7226 ( .A(n5284), .B(n5734), .X(n3793) );
  nand_x1_sg U7227 ( .A(\buff_mem[6][1] ), .B(n5557), .X(n3794) );
  nand_x1_sg U7228 ( .A(n5240), .B(n5730), .X(n3795) );
  nand_x1_sg U7229 ( .A(\buff_mem[6][2] ), .B(n5558), .X(n3796) );
  nand_x1_sg U7230 ( .A(n5286), .B(n5732), .X(n3797) );
  nand_x1_sg U7231 ( .A(\buff_mem[6][3] ), .B(n5559), .X(n3798) );
  nand_x1_sg U7232 ( .A(n5361), .B(n5734), .X(n3799) );
  nand_x1_sg U7233 ( .A(\buff_mem[6][4] ), .B(n5291), .X(n3800) );
  nand_x1_sg U7234 ( .A(n5252), .B(n5729), .X(n3801) );
  nand_x1_sg U7235 ( .A(\buff_mem[6][5] ), .B(n5558), .X(n3802) );
  nand_x1_sg U7236 ( .A(n5398), .B(n5733), .X(n3803) );
  nand_x1_sg U7237 ( .A(\buff_mem[6][6] ), .B(n5559), .X(n3804) );
  nand_x1_sg U7238 ( .A(n5428), .B(n5729), .X(n3805) );
  nand_x1_sg U7239 ( .A(\buff_mem[6][7] ), .B(n5291), .X(n3806) );
  nand_x1_sg U7240 ( .A(n5376), .B(n5732), .X(n3807) );
  nand_x1_sg U7241 ( .A(\buff_mem[6][8] ), .B(n5291), .X(n3808) );
  nand_x1_sg U7242 ( .A(n5649), .B(n5733), .X(n3809) );
  nand_x1_sg U7243 ( .A(\buff_mem[6][9] ), .B(n5559), .X(n3810) );
  nand_x1_sg U7244 ( .A(n5647), .B(n5732), .X(n3811) );
  nand_x1_sg U7245 ( .A(\buff_mem[6][10] ), .B(n5559), .X(n3812) );
  nand_x1_sg U7246 ( .A(n5535), .B(n5729), .X(n3813) );
  nand_x1_sg U7247 ( .A(\buff_mem[6][11] ), .B(n5556), .X(n3814) );
  nand_x1_sg U7248 ( .A(n5365), .B(n5730), .X(n3815) );
  nand_x1_sg U7249 ( .A(\buff_mem[6][12] ), .B(n5556), .X(n3816) );
  nand_x1_sg U7250 ( .A(n5248), .B(n5733), .X(n3817) );
  nand_x1_sg U7251 ( .A(\buff_mem[6][13] ), .B(n5558), .X(n3818) );
  nand_x1_sg U7252 ( .A(n5256), .B(n5727), .X(n3821) );
  nand_x1_sg U7253 ( .A(\buff_mem[6][15] ), .B(n5558), .X(n3822) );
  nand_x1_sg U7254 ( .A(n5369), .B(n5734), .X(n3823) );
  nand_x1_sg U7255 ( .A(\buff_mem[6][16] ), .B(n5556), .X(n3824) );
  nand_x1_sg U7256 ( .A(n5436), .B(n5732), .X(n3825) );
  nand_x1_sg U7257 ( .A(\buff_mem[6][17] ), .B(n5557), .X(n3826) );
  nand_x1_sg U7258 ( .A(n5403), .B(n5730), .X(n3827) );
  nand_x1_sg U7259 ( .A(\buff_mem[6][18] ), .B(n5556), .X(n3828) );
  nand_x1_sg U7260 ( .A(n5381), .B(n5729), .X(n3829) );
  nand_x1_sg U7261 ( .A(\buff_mem[6][19] ), .B(n5291), .X(n3830) );
  nand_x1_sg U7262 ( .A(n5521), .B(n5712), .X(n4130) );
  nand_x1_sg U7263 ( .A(\buff_mem[14][0] ), .B(n5630), .X(n4131) );
  nand_x1_sg U7264 ( .A(n5525), .B(n5713), .X(n4133) );
  nand_x1_sg U7265 ( .A(\buff_mem[14][1] ), .B(n5629), .X(n4134) );
  nand_x1_sg U7266 ( .A(n5394), .B(n5718), .X(n4135) );
  nand_x1_sg U7267 ( .A(\buff_mem[14][2] ), .B(n5632), .X(n4136) );
  nand_x1_sg U7268 ( .A(n5531), .B(n5720), .X(n4137) );
  nand_x1_sg U7269 ( .A(\buff_mem[14][3] ), .B(n5629), .X(n4138) );
  nand_x1_sg U7270 ( .A(n5226), .B(n5718), .X(n4139) );
  nand_x1_sg U7271 ( .A(\buff_mem[14][4] ), .B(n5631), .X(n4140) );
  nand_x1_sg U7272 ( .A(n5431), .B(n5715), .X(n4141) );
  nand_x1_sg U7273 ( .A(\buff_mem[14][5] ), .B(n5630), .X(n4142) );
  nand_x1_sg U7274 ( .A(n5400), .B(n5720), .X(n4143) );
  nand_x1_sg U7275 ( .A(\buff_mem[14][6] ), .B(n5306), .X(n4144) );
  nand_x1_sg U7276 ( .A(n5427), .B(n5719), .X(n4145) );
  nand_x1_sg U7277 ( .A(\buff_mem[14][7] ), .B(n5631), .X(n4146) );
  nand_x1_sg U7278 ( .A(n5374), .B(n5719), .X(n4147) );
  nand_x1_sg U7279 ( .A(\buff_mem[14][8] ), .B(n5306), .X(n4148) );
  nand_x1_sg U7280 ( .A(n5650), .B(n5712), .X(n4149) );
  nand_x1_sg U7281 ( .A(\buff_mem[14][9] ), .B(n5630), .X(n4150) );
  nand_x1_sg U7282 ( .A(n5644), .B(n5713), .X(n4151) );
  nand_x1_sg U7283 ( .A(\buff_mem[14][10] ), .B(n5632), .X(n4152) );
  nand_x1_sg U7284 ( .A(n5288), .B(n5719), .X(n4153) );
  nand_x1_sg U7285 ( .A(\buff_mem[14][11] ), .B(n5632), .X(n4154) );
  nand_x1_sg U7286 ( .A(n5363), .B(n5721), .X(n4155) );
  nand_x1_sg U7287 ( .A(\buff_mem[14][12] ), .B(n5306), .X(n4156) );
  nand_x1_sg U7288 ( .A(n5421), .B(n5712), .X(n4157) );
  nand_x1_sg U7289 ( .A(\buff_mem[14][13] ), .B(n5630), .X(n4158) );
  nand_x1_sg U7290 ( .A(n5441), .B(n5718), .X(n4161) );
  nand_x1_sg U7291 ( .A(\buff_mem[14][15] ), .B(n5629), .X(n4162) );
  nand_x1_sg U7292 ( .A(n5230), .B(n5718), .X(n4163) );
  nand_x1_sg U7293 ( .A(\buff_mem[14][16] ), .B(n5631), .X(n4164) );
  nand_x1_sg U7294 ( .A(n5437), .B(n5714), .X(n4165) );
  nand_x1_sg U7295 ( .A(\buff_mem[14][17] ), .B(n5629), .X(n4166) );
  nand_x1_sg U7296 ( .A(n5405), .B(n5721), .X(n4167) );
  nand_x1_sg U7297 ( .A(\buff_mem[14][18] ), .B(n5632), .X(n4168) );
  nand_x1_sg U7298 ( .A(n5234), .B(n5719), .X(n4169) );
  nand_x1_sg U7299 ( .A(\buff_mem[14][19] ), .B(n5306), .X(n4170) );
  nand_x1_sg U7300 ( .A(n5441), .B(n5710), .X(n3907) );
  nand_x1_sg U7301 ( .A(\buff_mem[8][15] ), .B(n5302), .X(n3908) );
  nand_x1_sg U7302 ( .A(n5440), .B(n5356), .X(n3949) );
  nand_x1_sg U7303 ( .A(\buff_mem[9][15] ), .B(n5548), .X(n3950) );
  nand_x1_sg U7304 ( .A(n5368), .B(n5705), .X(n3909) );
  nand_x1_sg U7305 ( .A(\buff_mem[8][16] ), .B(n5612), .X(n3910) );
  nand_x1_sg U7306 ( .A(n5369), .B(n5352), .X(n3951) );
  nand_x1_sg U7307 ( .A(\buff_mem[9][16] ), .B(n5548), .X(n3952) );
  nand_x1_sg U7308 ( .A(n5436), .B(n5710), .X(n3911) );
  nand_x1_sg U7309 ( .A(\buff_mem[8][17] ), .B(n5609), .X(n3912) );
  nand_x1_sg U7310 ( .A(n5435), .B(n5348), .X(n3953) );
  nand_x1_sg U7311 ( .A(\buff_mem[9][17] ), .B(n5547), .X(n3954) );
  nand_x1_sg U7312 ( .A(n5403), .B(n5711), .X(n3913) );
  nand_x1_sg U7313 ( .A(\buff_mem[8][18] ), .B(n5610), .X(n3914) );
  nand_x1_sg U7314 ( .A(n5406), .B(n5355), .X(n3955) );
  nand_x1_sg U7315 ( .A(\buff_mem[9][18] ), .B(n5549), .X(n3956) );
  nand_x1_sg U7316 ( .A(n5380), .B(n5707), .X(n3915) );
  nand_x1_sg U7317 ( .A(\buff_mem[8][19] ), .B(n5611), .X(n3916) );
  nand_x1_sg U7318 ( .A(n5234), .B(n5349), .X(n3957) );
  nand_x1_sg U7319 ( .A(\buff_mem[9][19] ), .B(n5547), .X(n3958) );
  nand_x1_sg U7320 ( .A(n5520), .B(n5707), .X(n3876) );
  nand_x1_sg U7321 ( .A(\buff_mem[8][0] ), .B(n5609), .X(n3877) );
  nand_x1_sg U7322 ( .A(n5523), .B(n5352), .X(n3918) );
  nand_x1_sg U7323 ( .A(\buff_mem[9][0] ), .B(n5548), .X(n3919) );
  nand_x1_sg U7324 ( .A(n5526), .B(n5707), .X(n3879) );
  nand_x1_sg U7325 ( .A(\buff_mem[8][1] ), .B(n5610), .X(n3880) );
  nand_x1_sg U7326 ( .A(n5527), .B(n5353), .X(n3921) );
  nand_x1_sg U7327 ( .A(\buff_mem[9][1] ), .B(n5547), .X(n3922) );
  nand_x1_sg U7328 ( .A(n5394), .B(n5705), .X(n3881) );
  nand_x1_sg U7329 ( .A(\buff_mem[8][2] ), .B(n5611), .X(n3882) );
  nand_x1_sg U7330 ( .A(n5395), .B(n5349), .X(n3923) );
  nand_x1_sg U7331 ( .A(\buff_mem[9][2] ), .B(n5549), .X(n3924) );
  nand_x1_sg U7332 ( .A(n5532), .B(n5706), .X(n3883) );
  nand_x1_sg U7333 ( .A(\buff_mem[8][3] ), .B(n5609), .X(n3884) );
  nand_x1_sg U7334 ( .A(n5531), .B(n5348), .X(n3925) );
  nand_x1_sg U7335 ( .A(\buff_mem[9][3] ), .B(n5546), .X(n3926) );
  nand_x1_sg U7336 ( .A(n5360), .B(n5706), .X(n3885) );
  nand_x1_sg U7337 ( .A(\buff_mem[8][4] ), .B(n5302), .X(n3886) );
  nand_x1_sg U7338 ( .A(n5360), .B(n5356), .X(n3927) );
  nand_x1_sg U7339 ( .A(\buff_mem[9][4] ), .B(n5549), .X(n3928) );
  nand_x1_sg U7340 ( .A(n5431), .B(n5711), .X(n3887) );
  nand_x1_sg U7341 ( .A(\buff_mem[8][5] ), .B(n5610), .X(n3888) );
  nand_x1_sg U7342 ( .A(n5432), .B(n5353), .X(n3929) );
  nand_x1_sg U7343 ( .A(\buff_mem[9][5] ), .B(n5546), .X(n3930) );
  nand_x1_sg U7344 ( .A(n5398), .B(n5711), .X(n3889) );
  nand_x1_sg U7345 ( .A(\buff_mem[8][6] ), .B(n5302), .X(n3890) );
  nand_x1_sg U7346 ( .A(n5399), .B(n5348), .X(n3931) );
  nand_x1_sg U7347 ( .A(\buff_mem[9][6] ), .B(n5289), .X(n3932) );
  nand_x1_sg U7348 ( .A(n5425), .B(n5706), .X(n3891) );
  nand_x1_sg U7349 ( .A(\buff_mem[8][7] ), .B(n5302), .X(n3892) );
  nand_x1_sg U7350 ( .A(n5426), .B(n5349), .X(n3933) );
  nand_x1_sg U7351 ( .A(\buff_mem[9][7] ), .B(n5546), .X(n3934) );
  nand_x1_sg U7352 ( .A(n5373), .B(n5705), .X(n3893) );
  nand_x1_sg U7353 ( .A(\buff_mem[8][8] ), .B(n5612), .X(n3894) );
  nand_x1_sg U7354 ( .A(n5232), .B(n5351), .X(n3935) );
  nand_x1_sg U7355 ( .A(\buff_mem[9][8] ), .B(n5549), .X(n3936) );
  nand_x1_sg U7356 ( .A(n5649), .B(n5709), .X(n3895) );
  nand_x1_sg U7357 ( .A(\buff_mem[8][9] ), .B(n5612), .X(n3896) );
  nand_x1_sg U7358 ( .A(n5651), .B(n5356), .X(n3937) );
  nand_x1_sg U7359 ( .A(\buff_mem[9][9] ), .B(n5289), .X(n3938) );
  nand_x1_sg U7360 ( .A(n5646), .B(n5710), .X(n3897) );
  nand_x1_sg U7361 ( .A(\buff_mem[8][10] ), .B(n5612), .X(n3898) );
  nand_x1_sg U7362 ( .A(n5646), .B(n5351), .X(n3939) );
  nand_x1_sg U7363 ( .A(\buff_mem[9][10] ), .B(n5289), .X(n3940) );
  nand_x1_sg U7364 ( .A(n5536), .B(n5705), .X(n3899) );
  nand_x1_sg U7365 ( .A(\buff_mem[8][11] ), .B(n5611), .X(n3900) );
  nand_x1_sg U7366 ( .A(n5537), .B(n5348), .X(n3941) );
  nand_x1_sg U7367 ( .A(\buff_mem[9][11] ), .B(n5547), .X(n3942) );
  nand_x1_sg U7368 ( .A(n5366), .B(n5709), .X(n3901) );
  nand_x1_sg U7369 ( .A(\buff_mem[8][12] ), .B(n5611), .X(n3902) );
  nand_x1_sg U7370 ( .A(n5364), .B(n3920), .X(n3943) );
  nand_x1_sg U7371 ( .A(\buff_mem[9][12] ), .B(n5546), .X(n3944) );
  nand_x1_sg U7372 ( .A(n5421), .B(n5706), .X(n3903) );
  nand_x1_sg U7373 ( .A(\buff_mem[8][13] ), .B(n5609), .X(n3904) );
  nand_x1_sg U7374 ( .A(n5422), .B(n5349), .X(n3945) );
  nand_x1_sg U7375 ( .A(\buff_mem[9][13] ), .B(n5289), .X(n3946) );
  nand_x1_sg U7376 ( .A(n5411), .B(n5724), .X(n4201) );
  nand_x1_sg U7377 ( .A(\buff_mem[15][14] ), .B(n5588), .X(n4202) );
  nand_x1_sg U7378 ( .A(n5282), .B(n5723), .X(n4172) );
  nand_x1_sg U7379 ( .A(\buff_mem[15][0] ), .B(n5587), .X(n4173) );
  nand_x1_sg U7380 ( .A(n5284), .B(n5725), .X(n4175) );
  nand_x1_sg U7381 ( .A(\buff_mem[15][1] ), .B(n5588), .X(n4176) );
  nand_x1_sg U7382 ( .A(n5394), .B(n5725), .X(n4177) );
  nand_x1_sg U7383 ( .A(\buff_mem[15][2] ), .B(n5586), .X(n4178) );
  nand_x1_sg U7384 ( .A(n5533), .B(n5725), .X(n4179) );
  nand_x1_sg U7385 ( .A(\buff_mem[15][3] ), .B(n5588), .X(n4180) );
  nand_x1_sg U7386 ( .A(n5359), .B(n5726), .X(n4181) );
  nand_x1_sg U7387 ( .A(\buff_mem[15][4] ), .B(n5586), .X(n4182) );
  nand_x1_sg U7388 ( .A(n5433), .B(n5724), .X(n4183) );
  nand_x1_sg U7389 ( .A(\buff_mem[15][5] ), .B(n5588), .X(n4184) );
  nand_x1_sg U7390 ( .A(n5400), .B(n5723), .X(n4185) );
  nand_x1_sg U7391 ( .A(\buff_mem[15][6] ), .B(n5586), .X(n4186) );
  nand_x1_sg U7392 ( .A(n5427), .B(n5725), .X(n4187) );
  nand_x1_sg U7393 ( .A(\buff_mem[15][7] ), .B(n5587), .X(n4188) );
  nand_x1_sg U7394 ( .A(n5376), .B(n5330), .X(n4189) );
  nand_x1_sg U7395 ( .A(\buff_mem[15][8] ), .B(n5589), .X(n4190) );
  nand_x1_sg U7396 ( .A(n5652), .B(n5726), .X(n4191) );
  nand_x1_sg U7397 ( .A(\buff_mem[15][9] ), .B(n5297), .X(n4192) );
  nand_x1_sg U7398 ( .A(n5644), .B(n5330), .X(n4193) );
  nand_x1_sg U7399 ( .A(\buff_mem[15][10] ), .B(n5297), .X(n4194) );
  nand_x1_sg U7400 ( .A(n5288), .B(n5724), .X(n4195) );
  nand_x1_sg U7401 ( .A(\buff_mem[15][11] ), .B(n5589), .X(n4196) );
  nand_x1_sg U7402 ( .A(n5228), .B(n5330), .X(n4197) );
  nand_x1_sg U7403 ( .A(\buff_mem[15][12] ), .B(n5297), .X(n4198) );
  nand_x1_sg U7404 ( .A(n5421), .B(n5726), .X(n4199) );
  nand_x1_sg U7405 ( .A(\buff_mem[15][13] ), .B(n5587), .X(n4200) );
  nand_x1_sg U7406 ( .A(n5256), .B(n5726), .X(n4203) );
  nand_x1_sg U7407 ( .A(\buff_mem[15][15] ), .B(n5587), .X(n4204) );
  nand_x1_sg U7408 ( .A(n5230), .B(n5723), .X(n4205) );
  nand_x1_sg U7409 ( .A(\buff_mem[15][16] ), .B(n5297), .X(n4206) );
  nand_x1_sg U7410 ( .A(n5438), .B(n5330), .X(n4207) );
  nand_x1_sg U7411 ( .A(\buff_mem[15][17] ), .B(n5589), .X(n4208) );
  nand_x1_sg U7412 ( .A(n5406), .B(n5724), .X(n4209) );
  nand_x1_sg U7413 ( .A(\buff_mem[15][18] ), .B(n5589), .X(n4210) );
  nand_x1_sg U7414 ( .A(n5381), .B(n5723), .X(n4211) );
  nand_x1_sg U7415 ( .A(\buff_mem[15][19] ), .B(n5586), .X(n4212) );
  nand_x1_sg U7416 ( .A(n5408), .B(n5332), .X(n3648) );
  nand_x1_sg U7417 ( .A(\buff_mem[2][14] ), .B(n5615), .X(n3649) );
  nand_x1_sg U7418 ( .A(n5440), .B(n5792), .X(n3650) );
  nand_x1_sg U7419 ( .A(\buff_mem[2][15] ), .B(n5616), .X(n3651) );
  nand_x1_sg U7420 ( .A(n5369), .B(n5789), .X(n3652) );
  nand_x1_sg U7421 ( .A(\buff_mem[2][16] ), .B(n5303), .X(n3653) );
  nand_x1_sg U7422 ( .A(n5438), .B(n5791), .X(n3654) );
  nand_x1_sg U7423 ( .A(\buff_mem[2][17] ), .B(n5617), .X(n3655) );
  nand_x1_sg U7424 ( .A(n5244), .B(n5332), .X(n3656) );
  nand_x1_sg U7425 ( .A(\buff_mem[2][18] ), .B(n5614), .X(n3657) );
  nand_x1_sg U7426 ( .A(n5379), .B(n5789), .X(n3658) );
  nand_x1_sg U7427 ( .A(\buff_mem[2][19] ), .B(n5614), .X(n3659) );
  nand_x1_sg U7428 ( .A(n5522), .B(n5791), .X(n3619) );
  nand_x1_sg U7429 ( .A(\buff_mem[2][0] ), .B(n5615), .X(n3620) );
  nand_x1_sg U7430 ( .A(n5525), .B(n5791), .X(n3622) );
  nand_x1_sg U7431 ( .A(\buff_mem[2][1] ), .B(n5617), .X(n3623) );
  nand_x1_sg U7432 ( .A(n5396), .B(n5332), .X(n3624) );
  nand_x1_sg U7433 ( .A(\buff_mem[2][2] ), .B(n5616), .X(n3625) );
  nand_x1_sg U7434 ( .A(n5530), .B(n5790), .X(n3626) );
  nand_x1_sg U7435 ( .A(\buff_mem[2][3] ), .B(n5615), .X(n3627) );
  nand_x1_sg U7436 ( .A(n5359), .B(n5332), .X(n3628) );
  nand_x1_sg U7437 ( .A(\buff_mem[2][4] ), .B(n5614), .X(n3629) );
  nand_x1_sg U7438 ( .A(n5431), .B(n5792), .X(n3630) );
  nand_x1_sg U7439 ( .A(\buff_mem[2][5] ), .B(n5615), .X(n3631) );
  nand_x1_sg U7440 ( .A(n5401), .B(n5791), .X(n3632) );
  nand_x1_sg U7441 ( .A(\buff_mem[2][6] ), .B(n5614), .X(n3633) );
  nand_x1_sg U7442 ( .A(n5425), .B(n5790), .X(n3634) );
  nand_x1_sg U7443 ( .A(\buff_mem[2][7] ), .B(n5616), .X(n3635) );
  nand_x1_sg U7444 ( .A(n5374), .B(n5789), .X(n3636) );
  nand_x1_sg U7445 ( .A(\buff_mem[2][8] ), .B(n5303), .X(n3637) );
  nand_x1_sg U7446 ( .A(n5649), .B(n5792), .X(n3638) );
  nand_x1_sg U7447 ( .A(\buff_mem[2][9] ), .B(n5303), .X(n3639) );
  nand_x1_sg U7448 ( .A(n5310), .B(n5792), .X(n3640) );
  nand_x1_sg U7449 ( .A(\buff_mem[2][10] ), .B(n5303), .X(n3641) );
  nand_x1_sg U7450 ( .A(n5538), .B(n5790), .X(n3642) );
  nand_x1_sg U7451 ( .A(\buff_mem[2][11] ), .B(n5616), .X(n3643) );
  nand_x1_sg U7452 ( .A(n5366), .B(n5789), .X(n3644) );
  nand_x1_sg U7453 ( .A(\buff_mem[2][12] ), .B(n5617), .X(n3645) );
  nand_x1_sg U7454 ( .A(n5423), .B(n5790), .X(n3646) );
  nand_x1_sg U7455 ( .A(\buff_mem[2][13] ), .B(n5617), .X(n3647) );
  nand_x1_sg U7456 ( .A(n5410), .B(n5681), .X(n3861) );
  nand_x1_sg U7457 ( .A(\buff_mem[7][14] ), .B(n5301), .X(n3862) );
  nand_x1_sg U7458 ( .A(n5246), .B(n5757), .X(n4031) );
  nand_x1_sg U7459 ( .A(\buff_mem[11][14] ), .B(n5581), .X(n4032) );
  nand_x1_sg U7460 ( .A(n5523), .B(n5687), .X(n3832) );
  nand_x1_sg U7461 ( .A(\buff_mem[7][0] ), .B(n5607), .X(n3833) );
  nand_x1_sg U7462 ( .A(n5525), .B(n5688), .X(n3835) );
  nand_x1_sg U7463 ( .A(\buff_mem[7][1] ), .B(n5301), .X(n3836) );
  nand_x1_sg U7464 ( .A(n5395), .B(n5684), .X(n3837) );
  nand_x1_sg U7465 ( .A(\buff_mem[7][2] ), .B(n5301), .X(n3838) );
  nand_x1_sg U7466 ( .A(n5530), .B(n5681), .X(n3839) );
  nand_x1_sg U7467 ( .A(\buff_mem[7][3] ), .B(n5606), .X(n3840) );
  nand_x1_sg U7468 ( .A(n5359), .B(n5683), .X(n3841) );
  nand_x1_sg U7469 ( .A(\buff_mem[7][4] ), .B(n5607), .X(n3842) );
  nand_x1_sg U7470 ( .A(n5432), .B(n5690), .X(n3843) );
  nand_x1_sg U7471 ( .A(\buff_mem[7][5] ), .B(n5607), .X(n3844) );
  nand_x1_sg U7472 ( .A(n5399), .B(n5690), .X(n3845) );
  nand_x1_sg U7473 ( .A(\buff_mem[7][6] ), .B(n5608), .X(n3846) );
  nand_x1_sg U7474 ( .A(n5427), .B(n5687), .X(n3847) );
  nand_x1_sg U7475 ( .A(\buff_mem[7][7] ), .B(n5605), .X(n3848) );
  nand_x1_sg U7476 ( .A(n5232), .B(n5688), .X(n3849) );
  nand_x1_sg U7477 ( .A(\buff_mem[7][8] ), .B(n5605), .X(n3850) );
  nand_x1_sg U7478 ( .A(n5652), .B(n5682), .X(n3851) );
  nand_x1_sg U7479 ( .A(\buff_mem[7][9] ), .B(n5606), .X(n3852) );
  nand_x1_sg U7480 ( .A(n5645), .B(n5687), .X(n3853) );
  nand_x1_sg U7481 ( .A(\buff_mem[7][10] ), .B(n5608), .X(n3854) );
  nand_x1_sg U7482 ( .A(n5535), .B(n5681), .X(n3855) );
  nand_x1_sg U7483 ( .A(\buff_mem[7][11] ), .B(n5605), .X(n3856) );
  nand_x1_sg U7484 ( .A(n5228), .B(n5687), .X(n3857) );
  nand_x1_sg U7485 ( .A(\buff_mem[7][12] ), .B(n5606), .X(n3858) );
  nand_x1_sg U7486 ( .A(n5420), .B(n5689), .X(n3859) );
  nand_x1_sg U7487 ( .A(\buff_mem[7][13] ), .B(n5608), .X(n3860) );
  nand_x1_sg U7488 ( .A(n5442), .B(n5684), .X(n3863) );
  nand_x1_sg U7489 ( .A(\buff_mem[7][15] ), .B(n5301), .X(n3864) );
  nand_x1_sg U7490 ( .A(n5230), .B(n5689), .X(n3865) );
  nand_x1_sg U7491 ( .A(\buff_mem[7][16] ), .B(n5606), .X(n3866) );
  nand_x1_sg U7492 ( .A(n5437), .B(n5688), .X(n3867) );
  nand_x1_sg U7493 ( .A(\buff_mem[7][17] ), .B(n5607), .X(n3868) );
  nand_x1_sg U7494 ( .A(n5404), .B(n5682), .X(n3869) );
  nand_x1_sg U7495 ( .A(\buff_mem[7][18] ), .B(n5605), .X(n3870) );
  nand_x1_sg U7496 ( .A(n5379), .B(n5688), .X(n3871) );
  nand_x1_sg U7497 ( .A(\buff_mem[7][19] ), .B(n5608), .X(n3872) );
  nand_x1_sg U7498 ( .A(n5443), .B(n5759), .X(n4033) );
  nand_x1_sg U7499 ( .A(\buff_mem[11][15] ), .B(n5296), .X(n4034) );
  nand_x1_sg U7500 ( .A(n5370), .B(n5757), .X(n4035) );
  nand_x1_sg U7501 ( .A(\buff_mem[11][16] ), .B(n5583), .X(n4036) );
  nand_x1_sg U7502 ( .A(n5435), .B(n5751), .X(n4037) );
  nand_x1_sg U7503 ( .A(\buff_mem[11][17] ), .B(n5584), .X(n4038) );
  nand_x1_sg U7504 ( .A(n5403), .B(n5753), .X(n4039) );
  nand_x1_sg U7505 ( .A(\buff_mem[11][18] ), .B(n5582), .X(n4040) );
  nand_x1_sg U7506 ( .A(n5380), .B(n5757), .X(n4041) );
  nand_x1_sg U7507 ( .A(\buff_mem[11][19] ), .B(n5296), .X(n4042) );
  nand_x1_sg U7508 ( .A(n5520), .B(n5757), .X(n4002) );
  nand_x1_sg U7509 ( .A(\buff_mem[11][0] ), .B(n5296), .X(n4003) );
  nand_x1_sg U7510 ( .A(n5526), .B(n5750), .X(n4005) );
  nand_x1_sg U7511 ( .A(\buff_mem[11][1] ), .B(n5582), .X(n4006) );
  nand_x1_sg U7512 ( .A(n5394), .B(n5756), .X(n4007) );
  nand_x1_sg U7513 ( .A(\buff_mem[11][2] ), .B(n5583), .X(n4008) );
  nand_x1_sg U7514 ( .A(n5532), .B(n5750), .X(n4009) );
  nand_x1_sg U7515 ( .A(\buff_mem[11][3] ), .B(n5581), .X(n4010) );
  nand_x1_sg U7516 ( .A(n5360), .B(n5758), .X(n4011) );
  nand_x1_sg U7517 ( .A(\buff_mem[11][4] ), .B(n5583), .X(n4012) );
  nand_x1_sg U7518 ( .A(n5252), .B(n5756), .X(n4013) );
  nand_x1_sg U7519 ( .A(\buff_mem[11][5] ), .B(n5582), .X(n4014) );
  nand_x1_sg U7520 ( .A(n5242), .B(n5751), .X(n4015) );
  nand_x1_sg U7521 ( .A(\buff_mem[11][6] ), .B(n5583), .X(n4016) );
  nand_x1_sg U7522 ( .A(n5250), .B(n5756), .X(n4017) );
  nand_x1_sg U7523 ( .A(\buff_mem[11][7] ), .B(n5584), .X(n4018) );
  nand_x1_sg U7524 ( .A(n5232), .B(n5758), .X(n4019) );
  nand_x1_sg U7525 ( .A(\buff_mem[11][8] ), .B(n5581), .X(n4020) );
  nand_x1_sg U7526 ( .A(n5650), .B(n5750), .X(n4021) );
  nand_x1_sg U7527 ( .A(\buff_mem[11][9] ), .B(n5582), .X(n4022) );
  nand_x1_sg U7528 ( .A(n5646), .B(n5756), .X(n4023) );
  nand_x1_sg U7529 ( .A(\buff_mem[11][10] ), .B(n5584), .X(n4024) );
  nand_x1_sg U7530 ( .A(n5536), .B(n5759), .X(n4025) );
  nand_x1_sg U7531 ( .A(\buff_mem[11][11] ), .B(n5584), .X(n4026) );
  nand_x1_sg U7532 ( .A(n5363), .B(n5752), .X(n4027) );
  nand_x1_sg U7533 ( .A(\buff_mem[11][12] ), .B(n5296), .X(n4028) );
  nand_x1_sg U7534 ( .A(n5420), .B(n5753), .X(n4029) );
  nand_x1_sg U7535 ( .A(\buff_mem[11][13] ), .B(n5581), .X(n4030) );
  nand_x1_sg U7536 ( .A(n5409), .B(n5743), .X(n3557) );
  nand_x1_sg U7537 ( .A(\buff_mem[0][14] ), .B(n5293), .X(n3558) );
  nand_x1_sg U7538 ( .A(n5411), .B(n5806), .X(n3606) );
  nand_x1_sg U7539 ( .A(\buff_mem[1][14] ), .B(n5619), .X(n3607) );
  nand_x1_sg U7540 ( .A(n5441), .B(n5747), .X(n3560) );
  nand_x1_sg U7541 ( .A(\buff_mem[0][15] ), .B(n5566), .X(n3561) );
  nand_x1_sg U7542 ( .A(n5442), .B(n5805), .X(n3608) );
  nand_x1_sg U7543 ( .A(\buff_mem[1][15] ), .B(n5619), .X(n3609) );
  nand_x1_sg U7544 ( .A(n5230), .B(n5746), .X(n3563) );
  nand_x1_sg U7545 ( .A(\buff_mem[0][16] ), .B(n5293), .X(n3564) );
  nand_x1_sg U7546 ( .A(n5368), .B(n5810), .X(n3610) );
  nand_x1_sg U7547 ( .A(\buff_mem[1][16] ), .B(n5621), .X(n3611) );
  nand_x1_sg U7548 ( .A(n5435), .B(n5749), .X(n3566) );
  nand_x1_sg U7549 ( .A(\buff_mem[0][17] ), .B(n5566), .X(n3567) );
  nand_x1_sg U7550 ( .A(n5437), .B(n5809), .X(n3612) );
  nand_x1_sg U7551 ( .A(\buff_mem[1][17] ), .B(n5620), .X(n3613) );
  nand_x1_sg U7552 ( .A(n5244), .B(n5747), .X(n3569) );
  nand_x1_sg U7553 ( .A(\buff_mem[0][18] ), .B(n5569), .X(n3570) );
  nand_x1_sg U7554 ( .A(n5405), .B(n5805), .X(n3614) );
  nand_x1_sg U7555 ( .A(\buff_mem[1][18] ), .B(n5620), .X(n3615) );
  nand_x1_sg U7556 ( .A(n5381), .B(n5746), .X(n3572) );
  nand_x1_sg U7557 ( .A(\buff_mem[0][19] ), .B(n5293), .X(n3573) );
  nand_x1_sg U7558 ( .A(n5378), .B(n5804), .X(n3616) );
  nand_x1_sg U7559 ( .A(\buff_mem[1][19] ), .B(n5622), .X(n3617) );
  nand_x1_sg U7560 ( .A(n5520), .B(n5746), .X(n3514) );
  nand_x1_sg U7561 ( .A(\buff_mem[0][0] ), .B(n5567), .X(n3515) );
  nand_x1_sg U7562 ( .A(n5521), .B(n5808), .X(n3577) );
  nand_x1_sg U7563 ( .A(\buff_mem[1][0] ), .B(n5304), .X(n3578) );
  nand_x1_sg U7564 ( .A(n5526), .B(n5748), .X(n3518) );
  nand_x1_sg U7565 ( .A(\buff_mem[0][1] ), .B(n5567), .X(n3519) );
  nand_x1_sg U7566 ( .A(n5528), .B(n5810), .X(n3580) );
  nand_x1_sg U7567 ( .A(\buff_mem[1][1] ), .B(n5621), .X(n3581) );
  nand_x1_sg U7568 ( .A(n5240), .B(n5740), .X(n3521) );
  nand_x1_sg U7569 ( .A(\buff_mem[0][2] ), .B(n5568), .X(n3522) );
  nand_x1_sg U7570 ( .A(n5395), .B(n5810), .X(n3582) );
  nand_x1_sg U7571 ( .A(\buff_mem[1][2] ), .B(n5619), .X(n3583) );
  nand_x1_sg U7572 ( .A(n5532), .B(n5749), .X(n3524) );
  nand_x1_sg U7573 ( .A(\buff_mem[0][3] ), .B(n5569), .X(n3525) );
  nand_x1_sg U7574 ( .A(n5286), .B(n5808), .X(n3584) );
  nand_x1_sg U7575 ( .A(\buff_mem[1][3] ), .B(n5304), .X(n3585) );
  nand_x1_sg U7576 ( .A(n5226), .B(n5741), .X(n3527) );
  nand_x1_sg U7577 ( .A(\buff_mem[0][4] ), .B(n5568), .X(n3528) );
  nand_x1_sg U7578 ( .A(n5226), .B(n5808), .X(n3586) );
  nand_x1_sg U7579 ( .A(\buff_mem[1][4] ), .B(n5304), .X(n3587) );
  nand_x1_sg U7580 ( .A(n5433), .B(n5740), .X(n3530) );
  nand_x1_sg U7581 ( .A(\buff_mem[0][5] ), .B(n5567), .X(n3531) );
  nand_x1_sg U7582 ( .A(n5433), .B(n5809), .X(n3588) );
  nand_x1_sg U7583 ( .A(\buff_mem[1][5] ), .B(n5620), .X(n3589) );
  nand_x1_sg U7584 ( .A(n5398), .B(n5742), .X(n3533) );
  nand_x1_sg U7585 ( .A(\buff_mem[0][6] ), .B(n5569), .X(n3534) );
  nand_x1_sg U7586 ( .A(n5399), .B(n5805), .X(n3590) );
  nand_x1_sg U7587 ( .A(\buff_mem[1][6] ), .B(n5620), .X(n3591) );
  nand_x1_sg U7588 ( .A(n5426), .B(n5741), .X(n3536) );
  nand_x1_sg U7589 ( .A(\buff_mem[0][7] ), .B(n5293), .X(n3537) );
  nand_x1_sg U7590 ( .A(n5426), .B(n5809), .X(n3592) );
  nand_x1_sg U7591 ( .A(\buff_mem[1][7] ), .B(n5621), .X(n3593) );
  nand_x1_sg U7592 ( .A(n5374), .B(n5747), .X(n3539) );
  nand_x1_sg U7593 ( .A(\buff_mem[0][8] ), .B(n5568), .X(n3540) );
  nand_x1_sg U7594 ( .A(n5374), .B(n5810), .X(n3594) );
  nand_x1_sg U7595 ( .A(\buff_mem[1][8] ), .B(n5622), .X(n3595) );
  nand_x1_sg U7596 ( .A(n5312), .B(n5746), .X(n3542) );
  nand_x1_sg U7597 ( .A(\buff_mem[0][9] ), .B(n5569), .X(n3543) );
  nand_x1_sg U7598 ( .A(n5650), .B(n5809), .X(n3596) );
  nand_x1_sg U7599 ( .A(\buff_mem[1][9] ), .B(n5622), .X(n3597) );
  nand_x1_sg U7600 ( .A(n5310), .B(n5748), .X(n3545) );
  nand_x1_sg U7601 ( .A(\buff_mem[0][10] ), .B(n5567), .X(n3546) );
  nand_x1_sg U7602 ( .A(n5645), .B(n5806), .X(n3598) );
  nand_x1_sg U7603 ( .A(\buff_mem[1][10] ), .B(n5622), .X(n3599) );
  nand_x1_sg U7604 ( .A(n5537), .B(n5743), .X(n3548) );
  nand_x1_sg U7605 ( .A(\buff_mem[0][11] ), .B(n5568), .X(n3549) );
  nand_x1_sg U7606 ( .A(n5537), .B(n5808), .X(n3600) );
  nand_x1_sg U7607 ( .A(\buff_mem[1][11] ), .B(n5304), .X(n3601) );
  nand_x1_sg U7608 ( .A(n5363), .B(n5740), .X(n3551) );
  nand_x1_sg U7609 ( .A(\buff_mem[0][12] ), .B(n5566), .X(n3552) );
  nand_x1_sg U7610 ( .A(n5365), .B(n5804), .X(n3602) );
  nand_x1_sg U7611 ( .A(\buff_mem[1][12] ), .B(n5621), .X(n3603) );
  nand_x1_sg U7612 ( .A(n5248), .B(n5747), .X(n3554) );
  nand_x1_sg U7613 ( .A(\buff_mem[0][13] ), .B(n5566), .X(n3555) );
  nand_x1_sg U7614 ( .A(n5422), .B(n5806), .X(n3604) );
  nand_x1_sg U7615 ( .A(\buff_mem[1][13] ), .B(n5619), .X(n3605) );
  nor_x1_sg U7616 ( .A(n5834), .B(wr_ptr[0]), .X(n3468) );
  nand_x1_sg U7617 ( .A(n5836), .B(n3444), .X(n3443) );
  nand_x1_sg U7618 ( .A(n3447), .B(n5832), .X(n3445) );
  nand_x1_sg U7619 ( .A(rd_ptr[1]), .B(n3356), .X(n3446) );
  nor_x1_sg U7620 ( .A(n5833), .B(wr_ptr[1]), .X(n3469) );
  nand_x1_sg U7621 ( .A(n5318), .B(n5222), .X(n3480) );
  nand_x1_sg U7622 ( .A(n5836), .B(n3358), .X(n3481) );
  nand_x1_sg U7623 ( .A(n5410), .B(n5328), .X(n4329) );
  nand_x1_sg U7624 ( .A(\buff_mem[18][14] ), .B(n5624), .X(n4330) );
  nand_x1_sg U7625 ( .A(n5443), .B(n5678), .X(n4331) );
  nand_x1_sg U7626 ( .A(\buff_mem[18][15] ), .B(n5624), .X(n4332) );
  nand_x1_sg U7627 ( .A(n5370), .B(n5328), .X(n4333) );
  nand_x1_sg U7628 ( .A(\buff_mem[18][16] ), .B(n5624), .X(n4334) );
  nand_x1_sg U7629 ( .A(n5437), .B(n5678), .X(n4335) );
  nand_x1_sg U7630 ( .A(\buff_mem[18][17] ), .B(n5627), .X(n4336) );
  nand_x1_sg U7631 ( .A(n5403), .B(n5680), .X(n4337) );
  nand_x1_sg U7632 ( .A(\buff_mem[18][18] ), .B(n5626), .X(n4338) );
  nand_x1_sg U7633 ( .A(n5380), .B(n5677), .X(n4339) );
  nand_x1_sg U7634 ( .A(\buff_mem[18][19] ), .B(n5305), .X(n4340) );
  nand_x1_sg U7635 ( .A(n5520), .B(n5677), .X(n4300) );
  nand_x1_sg U7636 ( .A(\buff_mem[18][0] ), .B(n5625), .X(n4301) );
  nand_x1_sg U7637 ( .A(n5527), .B(n5678), .X(n4303) );
  nand_x1_sg U7638 ( .A(\buff_mem[18][1] ), .B(n5627), .X(n4304) );
  nand_x1_sg U7639 ( .A(n5396), .B(n5679), .X(n4305) );
  nand_x1_sg U7640 ( .A(\buff_mem[18][2] ), .B(n5626), .X(n4306) );
  nand_x1_sg U7641 ( .A(n5530), .B(n5679), .X(n4307) );
  nand_x1_sg U7642 ( .A(\buff_mem[18][3] ), .B(n5626), .X(n4308) );
  nand_x1_sg U7643 ( .A(n5359), .B(n5680), .X(n4309) );
  nand_x1_sg U7644 ( .A(\buff_mem[18][4] ), .B(n5624), .X(n4310) );
  nand_x1_sg U7645 ( .A(n5432), .B(n5679), .X(n4311) );
  nand_x1_sg U7646 ( .A(\buff_mem[18][5] ), .B(n5625), .X(n4312) );
  nand_x1_sg U7647 ( .A(n5399), .B(n5677), .X(n4313) );
  nand_x1_sg U7648 ( .A(\buff_mem[18][6] ), .B(n5626), .X(n4314) );
  nand_x1_sg U7649 ( .A(n5250), .B(n5328), .X(n4315) );
  nand_x1_sg U7650 ( .A(\buff_mem[18][7] ), .B(n5627), .X(n4316) );
  nand_x1_sg U7651 ( .A(n5375), .B(n5677), .X(n4317) );
  nand_x1_sg U7652 ( .A(\buff_mem[18][8] ), .B(n5305), .X(n4318) );
  nand_x1_sg U7653 ( .A(n5312), .B(n5680), .X(n4319) );
  nand_x1_sg U7654 ( .A(\buff_mem[18][9] ), .B(n5305), .X(n4320) );
  nand_x1_sg U7655 ( .A(n5645), .B(n5328), .X(n4321) );
  nand_x1_sg U7656 ( .A(\buff_mem[18][10] ), .B(n5305), .X(n4322) );
  nand_x1_sg U7657 ( .A(n5538), .B(n5678), .X(n4323) );
  nand_x1_sg U7658 ( .A(\buff_mem[18][11] ), .B(n5625), .X(n4324) );
  nand_x1_sg U7659 ( .A(n5228), .B(n5680), .X(n4325) );
  nand_x1_sg U7660 ( .A(\buff_mem[18][12] ), .B(n5627), .X(n4326) );
  nand_x1_sg U7661 ( .A(n5422), .B(n5679), .X(n4327) );
  nand_x1_sg U7662 ( .A(\buff_mem[18][13] ), .B(n5625), .X(n4328) );
  inv_x1_sg U7663 ( .A(wr_ptr[3]), .X(n3366) );
  nand_x1_sg U7664 ( .A(n5411), .B(n5699), .X(n4287) );
  nand_x1_sg U7665 ( .A(\buff_mem[17][14] ), .B(n5579), .X(n4288) );
  nand_x1_sg U7666 ( .A(n5442), .B(n5701), .X(n4289) );
  nand_x1_sg U7667 ( .A(\buff_mem[17][15] ), .B(n5578), .X(n4290) );
  nand_x1_sg U7668 ( .A(n5370), .B(n5329), .X(n4291) );
  nand_x1_sg U7669 ( .A(\buff_mem[17][16] ), .B(n5577), .X(n4292) );
  nand_x1_sg U7670 ( .A(n5254), .B(n5701), .X(n4293) );
  nand_x1_sg U7671 ( .A(\buff_mem[17][17] ), .B(n5579), .X(n4294) );
  nand_x1_sg U7672 ( .A(n5405), .B(n5702), .X(n4295) );
  nand_x1_sg U7673 ( .A(\buff_mem[17][18] ), .B(n5577), .X(n4296) );
  nand_x1_sg U7674 ( .A(n5379), .B(n5700), .X(n4297) );
  nand_x1_sg U7675 ( .A(\buff_mem[17][19] ), .B(n5577), .X(n4298) );
  nand_x1_sg U7676 ( .A(n5282), .B(n5700), .X(n4258) );
  nand_x1_sg U7677 ( .A(\buff_mem[17][0] ), .B(n5578), .X(n4259) );
  nand_x1_sg U7678 ( .A(n5284), .B(n5699), .X(n4261) );
  nand_x1_sg U7679 ( .A(\buff_mem[17][1] ), .B(n5577), .X(n4262) );
  nand_x1_sg U7680 ( .A(n5395), .B(n5700), .X(n4263) );
  nand_x1_sg U7681 ( .A(\buff_mem[17][2] ), .B(n5295), .X(n4264) );
  nand_x1_sg U7682 ( .A(n5531), .B(n5329), .X(n4265) );
  nand_x1_sg U7683 ( .A(\buff_mem[17][3] ), .B(n5578), .X(n4266) );
  nand_x1_sg U7684 ( .A(n5360), .B(n5702), .X(n4267) );
  nand_x1_sg U7685 ( .A(\buff_mem[17][4] ), .B(n5576), .X(n4268) );
  nand_x1_sg U7686 ( .A(n5431), .B(n5699), .X(n4269) );
  nand_x1_sg U7687 ( .A(\buff_mem[17][5] ), .B(n5576), .X(n4270) );
  nand_x1_sg U7688 ( .A(n5400), .B(n5701), .X(n4271) );
  nand_x1_sg U7689 ( .A(\buff_mem[17][6] ), .B(n5579), .X(n4272) );
  nand_x1_sg U7690 ( .A(n5250), .B(n5329), .X(n4273) );
  nand_x1_sg U7691 ( .A(\buff_mem[17][7] ), .B(n5578), .X(n4274) );
  nand_x1_sg U7692 ( .A(n5375), .B(n5700), .X(n4275) );
  nand_x1_sg U7693 ( .A(\buff_mem[17][8] ), .B(n5576), .X(n4276) );
  nand_x1_sg U7694 ( .A(n5652), .B(n5702), .X(n4277) );
  nand_x1_sg U7695 ( .A(\buff_mem[17][9] ), .B(n5295), .X(n4278) );
  nand_x1_sg U7696 ( .A(n5310), .B(n5329), .X(n4279) );
  nand_x1_sg U7697 ( .A(\buff_mem[17][10] ), .B(n5295), .X(n4280) );
  nand_x1_sg U7698 ( .A(n5538), .B(n5699), .X(n4281) );
  nand_x1_sg U7699 ( .A(\buff_mem[17][11] ), .B(n5579), .X(n4282) );
  nand_x1_sg U7700 ( .A(n5365), .B(n5702), .X(n4283) );
  nand_x1_sg U7701 ( .A(\buff_mem[17][12] ), .B(n5576), .X(n4284) );
  nand_x1_sg U7702 ( .A(n5420), .B(n5701), .X(n4285) );
  nand_x1_sg U7703 ( .A(\buff_mem[17][13] ), .B(n5295), .X(n4286) );
  nand_x1_sg U7704 ( .A(n5523), .B(n5666), .X(n4343) );
  nand_x1_sg U7705 ( .A(\buff_mem[19][0] ), .B(n5574), .X(n4342) );
  nand_x1_sg U7706 ( .A(n5411), .B(n5327), .X(n4372) );
  nand_x1_sg U7707 ( .A(\buff_mem[19][14] ), .B(n5574), .X(n4371) );
  nand_x1_sg U7708 ( .A(n5443), .B(n5667), .X(n4374) );
  nand_x1_sg U7709 ( .A(\buff_mem[19][15] ), .B(n5571), .X(n4373) );
  nand_x1_sg U7710 ( .A(n5371), .B(n5664), .X(n4376) );
  nand_x1_sg U7711 ( .A(\buff_mem[19][16] ), .B(n5572), .X(n4375) );
  nand_x1_sg U7712 ( .A(n5438), .B(n5666), .X(n4378) );
  nand_x1_sg U7713 ( .A(\buff_mem[19][17] ), .B(n5571), .X(n4377) );
  nand_x1_sg U7714 ( .A(n5406), .B(n5664), .X(n4380) );
  nand_x1_sg U7715 ( .A(\buff_mem[19][18] ), .B(n5573), .X(n4379) );
  nand_x1_sg U7716 ( .A(n5528), .B(n5665), .X(n4346) );
  nand_x1_sg U7717 ( .A(\buff_mem[19][1] ), .B(n5572), .X(n4345) );
  nand_x1_sg U7718 ( .A(n5396), .B(n5664), .X(n4348) );
  nand_x1_sg U7719 ( .A(\buff_mem[19][2] ), .B(n5571), .X(n4347) );
  nand_x1_sg U7720 ( .A(n5533), .B(n5667), .X(n4350) );
  nand_x1_sg U7721 ( .A(\buff_mem[19][3] ), .B(n5574), .X(n4349) );
  nand_x1_sg U7722 ( .A(n5361), .B(n5327), .X(n4352) );
  nand_x1_sg U7723 ( .A(\buff_mem[19][4] ), .B(n5572), .X(n4351) );
  nand_x1_sg U7724 ( .A(n5433), .B(n5327), .X(n4354) );
  nand_x1_sg U7725 ( .A(\buff_mem[19][5] ), .B(n5294), .X(n4353) );
  nand_x1_sg U7726 ( .A(n5401), .B(n5666), .X(n4356) );
  nand_x1_sg U7727 ( .A(\buff_mem[19][6] ), .B(n5573), .X(n4355) );
  nand_x1_sg U7728 ( .A(n5428), .B(n5665), .X(n4358) );
  nand_x1_sg U7729 ( .A(\buff_mem[19][7] ), .B(n5573), .X(n4357) );
  nand_x1_sg U7730 ( .A(n5376), .B(n5665), .X(n4360) );
  nand_x1_sg U7731 ( .A(\buff_mem[19][8] ), .B(n5572), .X(n4359) );
  nand_x1_sg U7732 ( .A(n5652), .B(n5665), .X(n4362) );
  nand_x1_sg U7733 ( .A(\buff_mem[19][9] ), .B(n5571), .X(n4361) );
  nand_x1_sg U7734 ( .A(n5647), .B(n5666), .X(n4364) );
  nand_x1_sg U7735 ( .A(\buff_mem[19][10] ), .B(n5574), .X(n4363) );
  nand_x1_sg U7736 ( .A(n5538), .B(n5327), .X(n4366) );
  nand_x1_sg U7737 ( .A(\buff_mem[19][11] ), .B(n5294), .X(n4365) );
  nand_x1_sg U7738 ( .A(n5366), .B(n5667), .X(n4368) );
  nand_x1_sg U7739 ( .A(\buff_mem[19][12] ), .B(n5294), .X(n4367) );
  nand_x1_sg U7740 ( .A(n5423), .B(n5667), .X(n4370) );
  nand_x1_sg U7741 ( .A(\buff_mem[19][13] ), .B(n5573), .X(n4369) );
  nand_x1_sg U7742 ( .A(n5340), .B(n3435), .X(n4392) );
  nand_x1_sg U7743 ( .A(n5906), .B(n3509), .X(n4393) );
  nand_x1_sg U7744 ( .A(n5246), .B(n5766), .X(n4245) );
  nand_x1_sg U7745 ( .A(\buff_mem[16][14] ), .B(n5552), .X(n4246) );
  nand_x1_sg U7746 ( .A(n5440), .B(n5763), .X(n4247) );
  nand_x1_sg U7747 ( .A(\buff_mem[16][15] ), .B(n5553), .X(n4248) );
  nand_x1_sg U7748 ( .A(n5369), .B(n5768), .X(n4249) );
  nand_x1_sg U7749 ( .A(\buff_mem[16][16] ), .B(n5551), .X(n4250) );
  nand_x1_sg U7750 ( .A(n5254), .B(n5767), .X(n4251) );
  nand_x1_sg U7751 ( .A(\buff_mem[16][17] ), .B(n5554), .X(n4252) );
  nand_x1_sg U7752 ( .A(n5244), .B(n5763), .X(n4253) );
  nand_x1_sg U7753 ( .A(\buff_mem[16][18] ), .B(n5552), .X(n4254) );
  nand_x1_sg U7754 ( .A(n5378), .B(n5767), .X(n4255) );
  nand_x1_sg U7755 ( .A(\buff_mem[16][19] ), .B(n5553), .X(n4256) );
  nand_x1_sg U7756 ( .A(n5282), .B(n5767), .X(n4216) );
  nand_x1_sg U7757 ( .A(\buff_mem[16][0] ), .B(n5554), .X(n4217) );
  nand_x1_sg U7758 ( .A(n5284), .B(n5766), .X(n4219) );
  nand_x1_sg U7759 ( .A(\buff_mem[16][1] ), .B(n5554), .X(n4220) );
  nand_x1_sg U7760 ( .A(n5393), .B(n5760), .X(n4221) );
  nand_x1_sg U7761 ( .A(\buff_mem[16][2] ), .B(n5553), .X(n4222) );
  nand_x1_sg U7762 ( .A(n5286), .B(n5760), .X(n4223) );
  nand_x1_sg U7763 ( .A(\buff_mem[16][3] ), .B(n5551), .X(n4224) );
  nand_x1_sg U7764 ( .A(n5358), .B(n5768), .X(n4225) );
  nand_x1_sg U7765 ( .A(\buff_mem[16][4] ), .B(n5553), .X(n4226) );
  nand_x1_sg U7766 ( .A(n5430), .B(n5761), .X(n4227) );
  nand_x1_sg U7767 ( .A(\buff_mem[16][5] ), .B(n5551), .X(n4228) );
  nand_x1_sg U7768 ( .A(n5242), .B(n5760), .X(n4229) );
  nand_x1_sg U7769 ( .A(\buff_mem[16][6] ), .B(n5552), .X(n4230) );
  nand_x1_sg U7770 ( .A(n5428), .B(n5769), .X(n4231) );
  nand_x1_sg U7771 ( .A(\buff_mem[16][7] ), .B(n5290), .X(n4232) );
  nand_x1_sg U7772 ( .A(n5232), .B(n5767), .X(n4233) );
  nand_x1_sg U7773 ( .A(\buff_mem[16][8] ), .B(n5290), .X(n4234) );
  nand_x1_sg U7774 ( .A(n5651), .B(n5761), .X(n4235) );
  nand_x1_sg U7775 ( .A(\buff_mem[16][9] ), .B(n5552), .X(n4236) );
  nand_x1_sg U7776 ( .A(n5646), .B(n5766), .X(n4237) );
  nand_x1_sg U7777 ( .A(\buff_mem[16][10] ), .B(n5554), .X(n4238) );
  nand_x1_sg U7778 ( .A(n5536), .B(n5769), .X(n4239) );
  nand_x1_sg U7779 ( .A(\buff_mem[16][11] ), .B(n5551), .X(n4240) );
  nand_x1_sg U7780 ( .A(n5364), .B(n5762), .X(n4241) );
  nand_x1_sg U7781 ( .A(\buff_mem[16][12] ), .B(n5290), .X(n4242) );
  nand_x1_sg U7782 ( .A(n5248), .B(n5766), .X(n4243) );
  nand_x1_sg U7783 ( .A(\buff_mem[16][13] ), .B(n5290), .X(n4244) );
  nand_x1_sg U7784 ( .A(n5234), .B(n5664), .X(n4381) );
  nand_x1_sg U7785 ( .A(\buff_mem[19][19] ), .B(n5294), .X(n4382) );
  nor_x1_sg U7786 ( .A(wr_ptr[0]), .B(wr_ptr[1]), .X(n3576) );
  nand_x1_sg U7787 ( .A(n5184), .B(rd_ptr[4]), .X(n4462) );
  nand_x1_sg U7788 ( .A(rd_ptr[1]), .B(n5913), .X(n4389) );
  nand_x1_sg U7789 ( .A(n5917), .B(n3499), .X(n4390) );
  nor_x1_sg U7790 ( .A(wr_ptr[3]), .B(wr_ptr[2]), .X(n3704) );
  nor_x1_sg U7791 ( .A(reset), .B(full), .X(n4387) );
  nand_x1_sg U7792 ( .A(n3465), .B(n5342), .X(n3475) );
  nand_x1_sg U7793 ( .A(n5346), .B(n3456), .X(n3476) );
  nand_x1_sg U7794 ( .A(n5318), .B(n5325), .X(n3470) );
  nand_x1_sg U7795 ( .A(n5836), .B(n3362), .X(n3471) );
  nand_x1_sg U7796 ( .A(n5318), .B(n5343), .X(n3466) );
  nand_x1_sg U7797 ( .A(n5346), .B(n3356), .X(n3467) );
  nor_x1_sg U7798 ( .A(n5916), .B(reset), .X(n3435) );
  nand_x1_sg U7799 ( .A(n5326), .B(n3333), .X(n3503) );
  nand_x1_sg U7800 ( .A(n5224), .B(n5833), .X(n3502) );
  nand_x1_sg U7801 ( .A(n5906), .B(n3333), .X(n3433) );
  nand_x1_sg U7802 ( .A(n5224), .B(n5913), .X(n3434) );
  nand_x1_sg U7803 ( .A(n5346), .B(n5833), .X(n3463) );
  nand_x1_sg U7804 ( .A(n3465), .B(n5326), .X(n3464) );
  inv_x1_sg U7805 ( .A(\buff_mem[2][0] ), .X(n3413) );
  inv_x1_sg U7806 ( .A(\buff_mem[2][1] ), .X(n3410) );
  inv_x1_sg U7807 ( .A(\buff_mem[2][2] ), .X(n3407) );
  inv_x1_sg U7808 ( .A(\buff_mem[2][3] ), .X(n3404) );
  inv_x1_sg U7809 ( .A(\buff_mem[2][4] ), .X(n3401) );
  inv_x1_sg U7810 ( .A(\buff_mem[2][5] ), .X(n3398) );
  inv_x1_sg U7811 ( .A(\buff_mem[2][6] ), .X(n3395) );
  inv_x1_sg U7812 ( .A(\buff_mem[2][7] ), .X(n3392) );
  inv_x1_sg U7813 ( .A(\buff_mem[2][8] ), .X(n3389) );
  inv_x1_sg U7814 ( .A(\buff_mem[2][9] ), .X(n3386) );
  inv_x1_sg U7815 ( .A(\buff_mem[2][10] ), .X(n3383) );
  inv_x1_sg U7816 ( .A(\buff_mem[2][11] ), .X(n3380) );
  inv_x1_sg U7817 ( .A(\buff_mem[2][12] ), .X(n3377) );
  inv_x1_sg U7818 ( .A(\buff_mem[2][13] ), .X(n3374) );
  inv_x1_sg U7819 ( .A(\buff_mem[2][14] ), .X(n3431) );
  inv_x1_sg U7820 ( .A(\buff_mem[2][15] ), .X(n3428) );
  inv_x1_sg U7821 ( .A(\buff_mem[2][16] ), .X(n3425) );
  inv_x1_sg U7822 ( .A(\buff_mem[2][17] ), .X(n3422) );
  inv_x1_sg U7823 ( .A(\buff_mem[2][18] ), .X(n3419) );
  inv_x1_sg U7824 ( .A(\buff_mem[2][19] ), .X(n3416) );
endmodule

