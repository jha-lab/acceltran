
module loss ( clk, reset, model, .yHat({\yHat[15][19] , \yHat[15][18] , 
        \yHat[15][17] , \yHat[15][16] , \yHat[15][15] , \yHat[15][14] , 
        \yHat[15][13] , \yHat[15][12] , \yHat[15][11] , \yHat[15][10] , 
        \yHat[15][9] , \yHat[15][8] , \yHat[15][7] , \yHat[15][6] , 
        \yHat[15][5] , \yHat[15][4] , \yHat[15][3] , \yHat[15][2] , 
        \yHat[15][1] , \yHat[15][0] , \yHat[14][19] , \yHat[14][18] , 
        \yHat[14][17] , \yHat[14][16] , \yHat[14][15] , \yHat[14][14] , 
        \yHat[14][13] , \yHat[14][12] , \yHat[14][11] , \yHat[14][10] , 
        \yHat[14][9] , \yHat[14][8] , \yHat[14][7] , \yHat[14][6] , 
        \yHat[14][5] , \yHat[14][4] , \yHat[14][3] , \yHat[14][2] , 
        \yHat[14][1] , \yHat[14][0] , \yHat[13][19] , \yHat[13][18] , 
        \yHat[13][17] , \yHat[13][16] , \yHat[13][15] , \yHat[13][14] , 
        \yHat[13][13] , \yHat[13][12] , \yHat[13][11] , \yHat[13][10] , 
        \yHat[13][9] , \yHat[13][8] , \yHat[13][7] , \yHat[13][6] , 
        \yHat[13][5] , \yHat[13][4] , \yHat[13][3] , \yHat[13][2] , 
        \yHat[13][1] , \yHat[13][0] , \yHat[12][19] , \yHat[12][18] , 
        \yHat[12][17] , \yHat[12][16] , \yHat[12][15] , \yHat[12][14] , 
        \yHat[12][13] , \yHat[12][12] , \yHat[12][11] , \yHat[12][10] , 
        \yHat[12][9] , \yHat[12][8] , \yHat[12][7] , \yHat[12][6] , 
        \yHat[12][5] , \yHat[12][4] , \yHat[12][3] , \yHat[12][2] , 
        \yHat[12][1] , \yHat[12][0] , \yHat[11][19] , \yHat[11][18] , 
        \yHat[11][17] , \yHat[11][16] , \yHat[11][15] , \yHat[11][14] , 
        \yHat[11][13] , \yHat[11][12] , \yHat[11][11] , \yHat[11][10] , 
        \yHat[11][9] , \yHat[11][8] , \yHat[11][7] , \yHat[11][6] , 
        \yHat[11][5] , \yHat[11][4] , \yHat[11][3] , \yHat[11][2] , 
        \yHat[11][1] , \yHat[11][0] , \yHat[10][19] , \yHat[10][18] , 
        \yHat[10][17] , \yHat[10][16] , \yHat[10][15] , \yHat[10][14] , 
        \yHat[10][13] , \yHat[10][12] , \yHat[10][11] , \yHat[10][10] , 
        \yHat[10][9] , \yHat[10][8] , \yHat[10][7] , \yHat[10][6] , 
        \yHat[10][5] , \yHat[10][4] , \yHat[10][3] , \yHat[10][2] , 
        \yHat[10][1] , \yHat[10][0] , \yHat[9][19] , \yHat[9][18] , 
        \yHat[9][17] , \yHat[9][16] , \yHat[9][15] , \yHat[9][14] , 
        \yHat[9][13] , \yHat[9][12] , \yHat[9][11] , \yHat[9][10] , 
        \yHat[9][9] , \yHat[9][8] , \yHat[9][7] , \yHat[9][6] , \yHat[9][5] , 
        \yHat[9][4] , \yHat[9][3] , \yHat[9][2] , \yHat[9][1] , \yHat[9][0] , 
        \yHat[8][19] , \yHat[8][18] , \yHat[8][17] , \yHat[8][16] , 
        \yHat[8][15] , \yHat[8][14] , \yHat[8][13] , \yHat[8][12] , 
        \yHat[8][11] , \yHat[8][10] , \yHat[8][9] , \yHat[8][8] , \yHat[8][7] , 
        \yHat[8][6] , \yHat[8][5] , \yHat[8][4] , \yHat[8][3] , \yHat[8][2] , 
        \yHat[8][1] , \yHat[8][0] , \yHat[7][19] , \yHat[7][18] , 
        \yHat[7][17] , \yHat[7][16] , \yHat[7][15] , \yHat[7][14] , 
        \yHat[7][13] , \yHat[7][12] , \yHat[7][11] , \yHat[7][10] , 
        \yHat[7][9] , \yHat[7][8] , \yHat[7][7] , \yHat[7][6] , \yHat[7][5] , 
        \yHat[7][4] , \yHat[7][3] , \yHat[7][2] , \yHat[7][1] , \yHat[7][0] , 
        \yHat[6][19] , \yHat[6][18] , \yHat[6][17] , \yHat[6][16] , 
        \yHat[6][15] , \yHat[6][14] , \yHat[6][13] , \yHat[6][12] , 
        \yHat[6][11] , \yHat[6][10] , \yHat[6][9] , \yHat[6][8] , \yHat[6][7] , 
        \yHat[6][6] , \yHat[6][5] , \yHat[6][4] , \yHat[6][3] , \yHat[6][2] , 
        \yHat[6][1] , \yHat[6][0] , \yHat[5][19] , \yHat[5][18] , 
        \yHat[5][17] , \yHat[5][16] , \yHat[5][15] , \yHat[5][14] , 
        \yHat[5][13] , \yHat[5][12] , \yHat[5][11] , \yHat[5][10] , 
        \yHat[5][9] , \yHat[5][8] , \yHat[5][7] , \yHat[5][6] , \yHat[5][5] , 
        \yHat[5][4] , \yHat[5][3] , \yHat[5][2] , \yHat[5][1] , \yHat[5][0] , 
        \yHat[4][19] , \yHat[4][18] , \yHat[4][17] , \yHat[4][16] , 
        \yHat[4][15] , \yHat[4][14] , \yHat[4][13] , \yHat[4][12] , 
        \yHat[4][11] , \yHat[4][10] , \yHat[4][9] , \yHat[4][8] , \yHat[4][7] , 
        \yHat[4][6] , \yHat[4][5] , \yHat[4][4] , \yHat[4][3] , \yHat[4][2] , 
        \yHat[4][1] , \yHat[4][0] , \yHat[3][19] , \yHat[3][18] , 
        \yHat[3][17] , \yHat[3][16] , \yHat[3][15] , \yHat[3][14] , 
        \yHat[3][13] , \yHat[3][12] , \yHat[3][11] , \yHat[3][10] , 
        \yHat[3][9] , \yHat[3][8] , \yHat[3][7] , \yHat[3][6] , \yHat[3][5] , 
        \yHat[3][4] , \yHat[3][3] , \yHat[3][2] , \yHat[3][1] , \yHat[3][0] , 
        \yHat[2][19] , \yHat[2][18] , \yHat[2][17] , \yHat[2][16] , 
        \yHat[2][15] , \yHat[2][14] , \yHat[2][13] , \yHat[2][12] , 
        \yHat[2][11] , \yHat[2][10] , \yHat[2][9] , \yHat[2][8] , \yHat[2][7] , 
        \yHat[2][6] , \yHat[2][5] , \yHat[2][4] , \yHat[2][3] , \yHat[2][2] , 
        \yHat[2][1] , \yHat[2][0] , \yHat[1][19] , \yHat[1][18] , 
        \yHat[1][17] , \yHat[1][16] , \yHat[1][15] , \yHat[1][14] , 
        \yHat[1][13] , \yHat[1][12] , \yHat[1][11] , \yHat[1][10] , 
        \yHat[1][9] , \yHat[1][8] , \yHat[1][7] , \yHat[1][6] , \yHat[1][5] , 
        \yHat[1][4] , \yHat[1][3] , \yHat[1][2] , \yHat[1][1] , \yHat[1][0] , 
        \yHat[0][19] , \yHat[0][18] , \yHat[0][17] , \yHat[0][16] , 
        \yHat[0][15] , \yHat[0][14] , \yHat[0][13] , \yHat[0][12] , 
        \yHat[0][11] , \yHat[0][10] , \yHat[0][9] , \yHat[0][8] , \yHat[0][7] , 
        \yHat[0][6] , \yHat[0][5] , \yHat[0][4] , \yHat[0][3] , \yHat[0][2] , 
        \yHat[0][1] , \yHat[0][0] }), .y({\y[15][19] , \y[15][18] , 
        \y[15][17] , \y[15][16] , \y[15][15] , \y[15][14] , \y[15][13] , 
        \y[15][12] , \y[15][11] , \y[15][10] , \y[15][9] , \y[15][8] , 
        \y[15][7] , \y[15][6] , \y[15][5] , \y[15][4] , \y[15][3] , \y[15][2] , 
        \y[15][1] , \y[15][0] , \y[14][19] , \y[14][18] , \y[14][17] , 
        \y[14][16] , \y[14][15] , \y[14][14] , \y[14][13] , \y[14][12] , 
        \y[14][11] , \y[14][10] , \y[14][9] , \y[14][8] , \y[14][7] , 
        \y[14][6] , \y[14][5] , \y[14][4] , \y[14][3] , \y[14][2] , \y[14][1] , 
        \y[14][0] , \y[13][19] , \y[13][18] , \y[13][17] , \y[13][16] , 
        \y[13][15] , \y[13][14] , \y[13][13] , \y[13][12] , \y[13][11] , 
        \y[13][10] , \y[13][9] , \y[13][8] , \y[13][7] , \y[13][6] , 
        \y[13][5] , \y[13][4] , \y[13][3] , \y[13][2] , \y[13][1] , \y[13][0] , 
        \y[12][19] , \y[12][18] , \y[12][17] , \y[12][16] , \y[12][15] , 
        \y[12][14] , \y[12][13] , \y[12][12] , \y[12][11] , \y[12][10] , 
        \y[12][9] , \y[12][8] , \y[12][7] , \y[12][6] , \y[12][5] , \y[12][4] , 
        \y[12][3] , \y[12][2] , \y[12][1] , \y[12][0] , \y[11][19] , 
        \y[11][18] , \y[11][17] , \y[11][16] , \y[11][15] , \y[11][14] , 
        \y[11][13] , \y[11][12] , \y[11][11] , \y[11][10] , \y[11][9] , 
        \y[11][8] , \y[11][7] , \y[11][6] , \y[11][5] , \y[11][4] , \y[11][3] , 
        \y[11][2] , \y[11][1] , \y[11][0] , \y[10][19] , \y[10][18] , 
        \y[10][17] , \y[10][16] , \y[10][15] , \y[10][14] , \y[10][13] , 
        \y[10][12] , \y[10][11] , \y[10][10] , \y[10][9] , \y[10][8] , 
        \y[10][7] , \y[10][6] , \y[10][5] , \y[10][4] , \y[10][3] , \y[10][2] , 
        \y[10][1] , \y[10][0] , \y[9][19] , \y[9][18] , \y[9][17] , \y[9][16] , 
        \y[9][15] , \y[9][14] , \y[9][13] , \y[9][12] , \y[9][11] , \y[9][10] , 
        \y[9][9] , \y[9][8] , \y[9][7] , \y[9][6] , \y[9][5] , \y[9][4] , 
        \y[9][3] , \y[9][2] , \y[9][1] , \y[9][0] , \y[8][19] , \y[8][18] , 
        \y[8][17] , \y[8][16] , \y[8][15] , \y[8][14] , \y[8][13] , \y[8][12] , 
        \y[8][11] , \y[8][10] , \y[8][9] , \y[8][8] , \y[8][7] , \y[8][6] , 
        \y[8][5] , \y[8][4] , \y[8][3] , \y[8][2] , \y[8][1] , \y[8][0] , 
        \y[7][19] , \y[7][18] , \y[7][17] , \y[7][16] , \y[7][15] , \y[7][14] , 
        \y[7][13] , \y[7][12] , \y[7][11] , \y[7][10] , \y[7][9] , \y[7][8] , 
        \y[7][7] , \y[7][6] , \y[7][5] , \y[7][4] , \y[7][3] , \y[7][2] , 
        \y[7][1] , \y[7][0] , \y[6][19] , \y[6][18] , \y[6][17] , \y[6][16] , 
        \y[6][15] , \y[6][14] , \y[6][13] , \y[6][12] , \y[6][11] , \y[6][10] , 
        \y[6][9] , \y[6][8] , \y[6][7] , \y[6][6] , \y[6][5] , \y[6][4] , 
        \y[6][3] , \y[6][2] , \y[6][1] , \y[6][0] , \y[5][19] , \y[5][18] , 
        \y[5][17] , \y[5][16] , \y[5][15] , \y[5][14] , \y[5][13] , \y[5][12] , 
        \y[5][11] , \y[5][10] , \y[5][9] , \y[5][8] , \y[5][7] , \y[5][6] , 
        \y[5][5] , \y[5][4] , \y[5][3] , \y[5][2] , \y[5][1] , \y[5][0] , 
        \y[4][19] , \y[4][18] , \y[4][17] , \y[4][16] , \y[4][15] , \y[4][14] , 
        \y[4][13] , \y[4][12] , \y[4][11] , \y[4][10] , \y[4][9] , \y[4][8] , 
        \y[4][7] , \y[4][6] , \y[4][5] , \y[4][4] , \y[4][3] , \y[4][2] , 
        \y[4][1] , \y[4][0] , \y[3][19] , \y[3][18] , \y[3][17] , \y[3][16] , 
        \y[3][15] , \y[3][14] , \y[3][13] , \y[3][12] , \y[3][11] , \y[3][10] , 
        \y[3][9] , \y[3][8] , \y[3][7] , \y[3][6] , \y[3][5] , \y[3][4] , 
        \y[3][3] , \y[3][2] , \y[3][1] , \y[3][0] , \y[2][19] , \y[2][18] , 
        \y[2][17] , \y[2][16] , \y[2][15] , \y[2][14] , \y[2][13] , \y[2][12] , 
        \y[2][11] , \y[2][10] , \y[2][9] , \y[2][8] , \y[2][7] , \y[2][6] , 
        \y[2][5] , \y[2][4] , \y[2][3] , \y[2][2] , \y[2][1] , \y[2][0] , 
        \y[1][19] , \y[1][18] , \y[1][17] , \y[1][16] , \y[1][15] , \y[1][14] , 
        \y[1][13] , \y[1][12] , \y[1][11] , \y[1][10] , \y[1][9] , \y[1][8] , 
        \y[1][7] , \y[1][6] , \y[1][5] , \y[1][4] , \y[1][3] , \y[1][2] , 
        \y[1][1] , \y[1][0] , \y[0][19] , \y[0][18] , \y[0][17] , \y[0][16] , 
        \y[0][15] , \y[0][14] , \y[0][13] , \y[0][12] , \y[0][11] , \y[0][10] , 
        \y[0][9] , \y[0][8] , \y[0][7] , \y[0][6] , \y[0][5] , \y[0][4] , 
        \y[0][3] , \y[0][2] , \y[0][1] , \y[0][0] }), num, input_ready, 
        output_taken, state, out );
  input [3:0] num;
  output [1:0] state;
  output [19:0] out;
  input clk, reset, model, \yHat[15][19] , \yHat[15][18] , \yHat[15][17] ,
         \yHat[15][16] , \yHat[15][15] , \yHat[15][14] , \yHat[15][13] ,
         \yHat[15][12] , \yHat[15][11] , \yHat[15][10] , \yHat[15][9] ,
         \yHat[15][8] , \yHat[15][7] , \yHat[15][6] , \yHat[15][5] ,
         \yHat[15][4] , \yHat[15][3] , \yHat[15][2] , \yHat[15][1] ,
         \yHat[15][0] , \yHat[14][19] , \yHat[14][18] , \yHat[14][17] ,
         \yHat[14][16] , \yHat[14][15] , \yHat[14][14] , \yHat[14][13] ,
         \yHat[14][12] , \yHat[14][11] , \yHat[14][10] , \yHat[14][9] ,
         \yHat[14][8] , \yHat[14][7] , \yHat[14][6] , \yHat[14][5] ,
         \yHat[14][4] , \yHat[14][3] , \yHat[14][2] , \yHat[14][1] ,
         \yHat[14][0] , \yHat[13][19] , \yHat[13][18] , \yHat[13][17] ,
         \yHat[13][16] , \yHat[13][15] , \yHat[13][14] , \yHat[13][13] ,
         \yHat[13][12] , \yHat[13][11] , \yHat[13][10] , \yHat[13][9] ,
         \yHat[13][8] , \yHat[13][7] , \yHat[13][6] , \yHat[13][5] ,
         \yHat[13][4] , \yHat[13][3] , \yHat[13][2] , \yHat[13][1] ,
         \yHat[13][0] , \yHat[12][19] , \yHat[12][18] , \yHat[12][17] ,
         \yHat[12][16] , \yHat[12][15] , \yHat[12][14] , \yHat[12][13] ,
         \yHat[12][12] , \yHat[12][11] , \yHat[12][10] , \yHat[12][9] ,
         \yHat[12][8] , \yHat[12][7] , \yHat[12][6] , \yHat[12][5] ,
         \yHat[12][4] , \yHat[12][3] , \yHat[12][2] , \yHat[12][1] ,
         \yHat[12][0] , \yHat[11][19] , \yHat[11][18] , \yHat[11][17] ,
         \yHat[11][16] , \yHat[11][15] , \yHat[11][14] , \yHat[11][13] ,
         \yHat[11][12] , \yHat[11][11] , \yHat[11][10] , \yHat[11][9] ,
         \yHat[11][8] , \yHat[11][7] , \yHat[11][6] , \yHat[11][5] ,
         \yHat[11][4] , \yHat[11][3] , \yHat[11][2] , \yHat[11][1] ,
         \yHat[11][0] , \yHat[10][19] , \yHat[10][18] , \yHat[10][17] ,
         \yHat[10][16] , \yHat[10][15] , \yHat[10][14] , \yHat[10][13] ,
         \yHat[10][12] , \yHat[10][11] , \yHat[10][10] , \yHat[10][9] ,
         \yHat[10][8] , \yHat[10][7] , \yHat[10][6] , \yHat[10][5] ,
         \yHat[10][4] , \yHat[10][3] , \yHat[10][2] , \yHat[10][1] ,
         \yHat[10][0] , \yHat[9][19] , \yHat[9][18] , \yHat[9][17] ,
         \yHat[9][16] , \yHat[9][15] , \yHat[9][14] , \yHat[9][13] ,
         \yHat[9][12] , \yHat[9][11] , \yHat[9][10] , \yHat[9][9] ,
         \yHat[9][8] , \yHat[9][7] , \yHat[9][6] , \yHat[9][5] , \yHat[9][4] ,
         \yHat[9][3] , \yHat[9][2] , \yHat[9][1] , \yHat[9][0] , \yHat[8][19] ,
         \yHat[8][18] , \yHat[8][17] , \yHat[8][16] , \yHat[8][15] ,
         \yHat[8][14] , \yHat[8][13] , \yHat[8][12] , \yHat[8][11] ,
         \yHat[8][10] , \yHat[8][9] , \yHat[8][8] , \yHat[8][7] , \yHat[8][6] ,
         \yHat[8][5] , \yHat[8][4] , \yHat[8][3] , \yHat[8][2] , \yHat[8][1] ,
         \yHat[8][0] , \yHat[7][19] , \yHat[7][18] , \yHat[7][17] ,
         \yHat[7][16] , \yHat[7][15] , \yHat[7][14] , \yHat[7][13] ,
         \yHat[7][12] , \yHat[7][11] , \yHat[7][10] , \yHat[7][9] ,
         \yHat[7][8] , \yHat[7][7] , \yHat[7][6] , \yHat[7][5] , \yHat[7][4] ,
         \yHat[7][3] , \yHat[7][2] , \yHat[7][1] , \yHat[7][0] , \yHat[6][19] ,
         \yHat[6][18] , \yHat[6][17] , \yHat[6][16] , \yHat[6][15] ,
         \yHat[6][14] , \yHat[6][13] , \yHat[6][12] , \yHat[6][11] ,
         \yHat[6][10] , \yHat[6][9] , \yHat[6][8] , \yHat[6][7] , \yHat[6][6] ,
         \yHat[6][5] , \yHat[6][4] , \yHat[6][3] , \yHat[6][2] , \yHat[6][1] ,
         \yHat[6][0] , \yHat[5][19] , \yHat[5][18] , \yHat[5][17] ,
         \yHat[5][16] , \yHat[5][15] , \yHat[5][14] , \yHat[5][13] ,
         \yHat[5][12] , \yHat[5][11] , \yHat[5][10] , \yHat[5][9] ,
         \yHat[5][8] , \yHat[5][7] , \yHat[5][6] , \yHat[5][5] , \yHat[5][4] ,
         \yHat[5][3] , \yHat[5][2] , \yHat[5][1] , \yHat[5][0] , \yHat[4][19] ,
         \yHat[4][18] , \yHat[4][17] , \yHat[4][16] , \yHat[4][15] ,
         \yHat[4][14] , \yHat[4][13] , \yHat[4][12] , \yHat[4][11] ,
         \yHat[4][10] , \yHat[4][9] , \yHat[4][8] , \yHat[4][7] , \yHat[4][6] ,
         \yHat[4][5] , \yHat[4][4] , \yHat[4][3] , \yHat[4][2] , \yHat[4][1] ,
         \yHat[4][0] , \yHat[3][19] , \yHat[3][18] , \yHat[3][17] ,
         \yHat[3][16] , \yHat[3][15] , \yHat[3][14] , \yHat[3][13] ,
         \yHat[3][12] , \yHat[3][11] , \yHat[3][10] , \yHat[3][9] ,
         \yHat[3][8] , \yHat[3][7] , \yHat[3][6] , \yHat[3][5] , \yHat[3][4] ,
         \yHat[3][3] , \yHat[3][2] , \yHat[3][1] , \yHat[3][0] , \yHat[2][19] ,
         \yHat[2][18] , \yHat[2][17] , \yHat[2][16] , \yHat[2][15] ,
         \yHat[2][14] , \yHat[2][13] , \yHat[2][12] , \yHat[2][11] ,
         \yHat[2][10] , \yHat[2][9] , \yHat[2][8] , \yHat[2][7] , \yHat[2][6] ,
         \yHat[2][5] , \yHat[2][4] , \yHat[2][3] , \yHat[2][2] , \yHat[2][1] ,
         \yHat[2][0] , \yHat[1][19] , \yHat[1][18] , \yHat[1][17] ,
         \yHat[1][16] , \yHat[1][15] , \yHat[1][14] , \yHat[1][13] ,
         \yHat[1][12] , \yHat[1][11] , \yHat[1][10] , \yHat[1][9] ,
         \yHat[1][8] , \yHat[1][7] , \yHat[1][6] , \yHat[1][5] , \yHat[1][4] ,
         \yHat[1][3] , \yHat[1][2] , \yHat[1][1] , \yHat[1][0] , \yHat[0][19] ,
         \yHat[0][18] , \yHat[0][17] , \yHat[0][16] , \yHat[0][15] ,
         \yHat[0][14] , \yHat[0][13] , \yHat[0][12] , \yHat[0][11] ,
         \yHat[0][10] , \yHat[0][9] , \yHat[0][8] , \yHat[0][7] , \yHat[0][6] ,
         \yHat[0][5] , \yHat[0][4] , \yHat[0][3] , \yHat[0][2] , \yHat[0][1] ,
         \yHat[0][0] , \y[15][19] , \y[15][18] , \y[15][17] , \y[15][16] ,
         \y[15][15] , \y[15][14] , \y[15][13] , \y[15][12] , \y[15][11] ,
         \y[15][10] , \y[15][9] , \y[15][8] , \y[15][7] , \y[15][6] ,
         \y[15][5] , \y[15][4] , \y[15][3] , \y[15][2] , \y[15][1] ,
         \y[15][0] , \y[14][19] , \y[14][18] , \y[14][17] , \y[14][16] ,
         \y[14][15] , \y[14][14] , \y[14][13] , \y[14][12] , \y[14][11] ,
         \y[14][10] , \y[14][9] , \y[14][8] , \y[14][7] , \y[14][6] ,
         \y[14][5] , \y[14][4] , \y[14][3] , \y[14][2] , \y[14][1] ,
         \y[14][0] , \y[13][19] , \y[13][18] , \y[13][17] , \y[13][16] ,
         \y[13][15] , \y[13][14] , \y[13][13] , \y[13][12] , \y[13][11] ,
         \y[13][10] , \y[13][9] , \y[13][8] , \y[13][7] , \y[13][6] ,
         \y[13][5] , \y[13][4] , \y[13][3] , \y[13][2] , \y[13][1] ,
         \y[13][0] , \y[12][19] , \y[12][18] , \y[12][17] , \y[12][16] ,
         \y[12][15] , \y[12][14] , \y[12][13] , \y[12][12] , \y[12][11] ,
         \y[12][10] , \y[12][9] , \y[12][8] , \y[12][7] , \y[12][6] ,
         \y[12][5] , \y[12][4] , \y[12][3] , \y[12][2] , \y[12][1] ,
         \y[12][0] , \y[11][19] , \y[11][18] , \y[11][17] , \y[11][16] ,
         \y[11][15] , \y[11][14] , \y[11][13] , \y[11][12] , \y[11][11] ,
         \y[11][10] , \y[11][9] , \y[11][8] , \y[11][7] , \y[11][6] ,
         \y[11][5] , \y[11][4] , \y[11][3] , \y[11][2] , \y[11][1] ,
         \y[11][0] , \y[10][19] , \y[10][18] , \y[10][17] , \y[10][16] ,
         \y[10][15] , \y[10][14] , \y[10][13] , \y[10][12] , \y[10][11] ,
         \y[10][10] , \y[10][9] , \y[10][8] , \y[10][7] , \y[10][6] ,
         \y[10][5] , \y[10][4] , \y[10][3] , \y[10][2] , \y[10][1] ,
         \y[10][0] , \y[9][19] , \y[9][18] , \y[9][17] , \y[9][16] ,
         \y[9][15] , \y[9][14] , \y[9][13] , \y[9][12] , \y[9][11] ,
         \y[9][10] , \y[9][9] , \y[9][8] , \y[9][7] , \y[9][6] , \y[9][5] ,
         \y[9][4] , \y[9][3] , \y[9][2] , \y[9][1] , \y[9][0] , \y[8][19] ,
         \y[8][18] , \y[8][17] , \y[8][16] , \y[8][15] , \y[8][14] ,
         \y[8][13] , \y[8][12] , \y[8][11] , \y[8][10] , \y[8][9] , \y[8][8] ,
         \y[8][7] , \y[8][6] , \y[8][5] , \y[8][4] , \y[8][3] , \y[8][2] ,
         \y[8][1] , \y[8][0] , \y[7][19] , \y[7][18] , \y[7][17] , \y[7][16] ,
         \y[7][15] , \y[7][14] , \y[7][13] , \y[7][12] , \y[7][11] ,
         \y[7][10] , \y[7][9] , \y[7][8] , \y[7][7] , \y[7][6] , \y[7][5] ,
         \y[7][4] , \y[7][3] , \y[7][2] , \y[7][1] , \y[7][0] , \y[6][19] ,
         \y[6][18] , \y[6][17] , \y[6][16] , \y[6][15] , \y[6][14] ,
         \y[6][13] , \y[6][12] , \y[6][11] , \y[6][10] , \y[6][9] , \y[6][8] ,
         \y[6][7] , \y[6][6] , \y[6][5] , \y[6][4] , \y[6][3] , \y[6][2] ,
         \y[6][1] , \y[6][0] , \y[5][19] , \y[5][18] , \y[5][17] , \y[5][16] ,
         \y[5][15] , \y[5][14] , \y[5][13] , \y[5][12] , \y[5][11] ,
         \y[5][10] , \y[5][9] , \y[5][8] , \y[5][7] , \y[5][6] , \y[5][5] ,
         \y[5][4] , \y[5][3] , \y[5][2] , \y[5][1] , \y[5][0] , \y[4][19] ,
         \y[4][18] , \y[4][17] , \y[4][16] , \y[4][15] , \y[4][14] ,
         \y[4][13] , \y[4][12] , \y[4][11] , \y[4][10] , \y[4][9] , \y[4][8] ,
         \y[4][7] , \y[4][6] , \y[4][5] , \y[4][4] , \y[4][3] , \y[4][2] ,
         \y[4][1] , \y[4][0] , \y[3][19] , \y[3][18] , \y[3][17] , \y[3][16] ,
         \y[3][15] , \y[3][14] , \y[3][13] , \y[3][12] , \y[3][11] ,
         \y[3][10] , \y[3][9] , \y[3][8] , \y[3][7] , \y[3][6] , \y[3][5] ,
         \y[3][4] , \y[3][3] , \y[3][2] , \y[3][1] , \y[3][0] , \y[2][19] ,
         \y[2][18] , \y[2][17] , \y[2][16] , \y[2][15] , \y[2][14] ,
         \y[2][13] , \y[2][12] , \y[2][11] , \y[2][10] , \y[2][9] , \y[2][8] ,
         \y[2][7] , \y[2][6] , \y[2][5] , \y[2][4] , \y[2][3] , \y[2][2] ,
         \y[2][1] , \y[2][0] , \y[1][19] , \y[1][18] , \y[1][17] , \y[1][16] ,
         \y[1][15] , \y[1][14] , \y[1][13] , \y[1][12] , \y[1][11] ,
         \y[1][10] , \y[1][9] , \y[1][8] , \y[1][7] , \y[1][6] , \y[1][5] ,
         \y[1][4] , \y[1][3] , \y[1][2] , \y[1][1] , \y[1][0] , \y[0][19] ,
         \y[0][18] , \y[0][17] , \y[0][16] , \y[0][15] , \y[0][14] ,
         \y[0][13] , \y[0][12] , \y[0][11] , \y[0][10] , \y[0][9] , \y[0][8] ,
         \y[0][7] , \y[0][6] , \y[0][5] , \y[0][4] , \y[0][3] , \y[0][2] ,
         \y[0][1] , \y[0][0] , input_ready, output_taken;
  wire   done, \reg_yHat[14][19] , \reg_yHat[14][18] , \reg_yHat[14][17] ,
         \reg_yHat[14][16] , \reg_yHat[14][15] , \reg_yHat[14][14] ,
         \reg_yHat[14][13] , \reg_yHat[14][12] , \reg_yHat[14][11] ,
         \reg_yHat[14][10] , \reg_yHat[14][9] , \reg_yHat[14][8] ,
         \reg_yHat[14][7] , \reg_yHat[14][6] , \reg_yHat[14][5] ,
         \reg_yHat[14][4] , \reg_yHat[14][3] , \reg_yHat[14][2] ,
         \reg_yHat[14][1] , \reg_yHat[14][0] , \reg_yHat[13][19] ,
         \reg_yHat[13][18] , \reg_yHat[13][17] , \reg_yHat[13][16] ,
         \reg_yHat[13][15] , \reg_yHat[13][14] , \reg_yHat[13][13] ,
         \reg_yHat[13][12] , \reg_yHat[13][11] , \reg_yHat[13][10] ,
         \reg_yHat[13][9] , \reg_yHat[13][8] , \reg_yHat[13][7] ,
         \reg_yHat[13][6] , \reg_yHat[13][5] , \reg_yHat[13][4] ,
         \reg_yHat[13][3] , \reg_yHat[13][2] , \reg_yHat[13][1] ,
         \reg_yHat[13][0] , \reg_yHat[12][19] , \reg_yHat[12][18] ,
         \reg_yHat[12][17] , \reg_yHat[12][16] , \reg_yHat[12][15] ,
         \reg_yHat[12][14] , \reg_yHat[12][13] , \reg_yHat[12][12] ,
         \reg_yHat[12][11] , \reg_yHat[12][10] , \reg_yHat[12][9] ,
         \reg_yHat[12][8] , \reg_yHat[12][7] , \reg_yHat[12][6] ,
         \reg_yHat[12][5] , \reg_yHat[12][4] , \reg_yHat[12][3] ,
         \reg_yHat[12][2] , \reg_yHat[12][1] , \reg_yHat[12][0] ,
         \reg_yHat[11][19] , \reg_yHat[11][18] , \reg_yHat[11][17] ,
         \reg_yHat[11][16] , \reg_yHat[11][15] , \reg_yHat[11][14] ,
         \reg_yHat[11][13] , \reg_yHat[11][12] , \reg_yHat[11][11] ,
         \reg_yHat[11][10] , \reg_yHat[11][9] , \reg_yHat[11][8] ,
         \reg_yHat[11][7] , \reg_yHat[11][6] , \reg_yHat[11][5] ,
         \reg_yHat[11][4] , \reg_yHat[11][3] , \reg_yHat[11][2] ,
         \reg_yHat[11][1] , \reg_yHat[11][0] , \reg_yHat[10][19] ,
         \reg_yHat[10][18] , \reg_yHat[10][17] , \reg_yHat[10][16] ,
         \reg_yHat[10][15] , \reg_yHat[10][14] , \reg_yHat[10][13] ,
         \reg_yHat[10][12] , \reg_yHat[10][11] , \reg_yHat[10][10] ,
         \reg_yHat[10][9] , \reg_yHat[10][8] , \reg_yHat[10][7] ,
         \reg_yHat[10][6] , \reg_yHat[10][5] , \reg_yHat[10][4] ,
         \reg_yHat[10][3] , \reg_yHat[10][2] , \reg_yHat[10][1] ,
         \reg_yHat[10][0] , \reg_yHat[9][19] , \reg_yHat[9][18] ,
         \reg_yHat[9][17] , \reg_yHat[9][16] , \reg_yHat[9][15] ,
         \reg_yHat[9][14] , \reg_yHat[9][13] , \reg_yHat[9][12] ,
         \reg_yHat[9][11] , \reg_yHat[9][10] , \reg_yHat[9][9] ,
         \reg_yHat[9][8] , \reg_yHat[9][7] , \reg_yHat[9][6] ,
         \reg_yHat[9][5] , \reg_yHat[9][4] , \reg_yHat[9][3] ,
         \reg_yHat[9][2] , \reg_yHat[9][1] , \reg_yHat[9][0] ,
         \reg_yHat[8][19] , \reg_yHat[8][18] , \reg_yHat[8][17] ,
         \reg_yHat[8][16] , \reg_yHat[8][15] , \reg_yHat[8][14] ,
         \reg_yHat[8][13] , \reg_yHat[8][12] , \reg_yHat[8][11] ,
         \reg_yHat[8][10] , \reg_yHat[8][9] , \reg_yHat[8][8] ,
         \reg_yHat[8][7] , \reg_yHat[8][6] , \reg_yHat[8][5] ,
         \reg_yHat[8][4] , \reg_yHat[8][3] , \reg_yHat[8][2] ,
         \reg_yHat[8][1] , \reg_yHat[8][0] , \reg_yHat[7][19] ,
         \reg_yHat[7][18] , \reg_yHat[7][17] , \reg_yHat[7][16] ,
         \reg_yHat[7][15] , \reg_yHat[7][14] , \reg_yHat[7][13] ,
         \reg_yHat[7][12] , \reg_yHat[7][11] , \reg_yHat[7][10] ,
         \reg_yHat[7][9] , \reg_yHat[7][8] , \reg_yHat[7][7] ,
         \reg_yHat[7][6] , \reg_yHat[7][5] , \reg_yHat[7][4] ,
         \reg_yHat[7][3] , \reg_yHat[7][2] , \reg_yHat[7][1] ,
         \reg_yHat[7][0] , \reg_yHat[6][19] , \reg_yHat[6][18] ,
         \reg_yHat[6][17] , \reg_yHat[6][16] , \reg_yHat[6][15] ,
         \reg_yHat[6][14] , \reg_yHat[6][13] , \reg_yHat[6][12] ,
         \reg_yHat[6][11] , \reg_yHat[6][10] , \reg_yHat[6][9] ,
         \reg_yHat[6][8] , \reg_yHat[6][7] , \reg_yHat[6][6] ,
         \reg_yHat[6][5] , \reg_yHat[6][4] , \reg_yHat[6][3] ,
         \reg_yHat[6][2] , \reg_yHat[6][1] , \reg_yHat[6][0] ,
         \reg_yHat[5][19] , \reg_yHat[5][18] , \reg_yHat[5][17] ,
         \reg_yHat[5][16] , \reg_yHat[5][15] , \reg_yHat[5][14] ,
         \reg_yHat[5][13] , \reg_yHat[5][12] , \reg_yHat[5][11] ,
         \reg_yHat[5][10] , \reg_yHat[5][9] , \reg_yHat[5][8] ,
         \reg_yHat[5][7] , \reg_yHat[5][6] , \reg_yHat[5][5] ,
         \reg_yHat[5][4] , \reg_yHat[5][3] , \reg_yHat[5][2] ,
         \reg_yHat[5][1] , \reg_yHat[5][0] , \reg_yHat[4][19] ,
         \reg_yHat[4][18] , \reg_yHat[4][17] , \reg_yHat[4][16] ,
         \reg_yHat[4][15] , \reg_yHat[4][14] , \reg_yHat[4][13] ,
         \reg_yHat[4][12] , \reg_yHat[4][11] , \reg_yHat[4][10] ,
         \reg_yHat[4][9] , \reg_yHat[4][8] , \reg_yHat[4][7] ,
         \reg_yHat[4][6] , \reg_yHat[4][5] , \reg_yHat[4][4] ,
         \reg_yHat[4][3] , \reg_yHat[4][2] , \reg_yHat[4][1] ,
         \reg_yHat[4][0] , \reg_yHat[3][19] , \reg_yHat[3][18] ,
         \reg_yHat[3][17] , \reg_yHat[3][16] , \reg_yHat[3][15] ,
         \reg_yHat[3][14] , \reg_yHat[3][13] , \reg_yHat[3][12] ,
         \reg_yHat[3][11] , \reg_yHat[3][10] , \reg_yHat[3][9] ,
         \reg_yHat[3][8] , \reg_yHat[3][7] , \reg_yHat[3][6] ,
         \reg_yHat[3][5] , \reg_yHat[3][4] , \reg_yHat[3][3] ,
         \reg_yHat[3][2] , \reg_yHat[3][1] , \reg_yHat[3][0] ,
         \reg_yHat[2][19] , \reg_yHat[2][18] , \reg_yHat[2][17] ,
         \reg_yHat[2][16] , \reg_yHat[2][15] , \reg_yHat[2][14] ,
         \reg_yHat[2][13] , \reg_yHat[2][12] , \reg_yHat[2][11] ,
         \reg_yHat[2][10] , \reg_yHat[2][9] , \reg_yHat[2][8] ,
         \reg_yHat[2][7] , \reg_yHat[2][6] , \reg_yHat[2][5] ,
         \reg_yHat[2][4] , \reg_yHat[2][3] , \reg_yHat[2][2] ,
         \reg_yHat[2][1] , \reg_yHat[2][0] , \reg_yHat[1][19] ,
         \reg_yHat[1][18] , \reg_yHat[1][17] , \reg_yHat[1][16] ,
         \reg_yHat[1][15] , \reg_yHat[1][14] , \reg_yHat[1][13] ,
         \reg_yHat[1][12] , \reg_yHat[1][11] , \reg_yHat[1][10] ,
         \reg_yHat[1][9] , \reg_yHat[1][8] , \reg_yHat[1][7] ,
         \reg_yHat[1][6] , \reg_yHat[1][5] , \reg_yHat[1][4] ,
         \reg_yHat[1][3] , \reg_yHat[1][2] , \reg_yHat[1][1] ,
         \reg_yHat[1][0] , \reg_yHat[0][19] , \reg_yHat[0][18] ,
         \reg_yHat[0][17] , \reg_yHat[0][16] , \reg_yHat[0][15] ,
         \reg_yHat[0][14] , \reg_yHat[0][13] , \reg_yHat[0][12] ,
         \reg_yHat[0][11] , \reg_yHat[0][10] , \reg_yHat[0][9] ,
         \reg_yHat[0][8] , \reg_yHat[0][7] , \reg_yHat[0][6] ,
         \reg_yHat[0][5] , \reg_yHat[0][4] , \reg_yHat[0][3] ,
         \reg_yHat[0][2] , \reg_yHat[0][1] , \reg_yHat[0][0] , \reg_y[14][19] ,
         \reg_y[14][18] , \reg_y[14][17] , \reg_y[14][16] , \reg_y[14][15] ,
         \reg_y[14][14] , \reg_y[14][13] , \reg_y[14][12] , \reg_y[14][11] ,
         \reg_y[14][10] , \reg_y[14][9] , \reg_y[14][8] , \reg_y[14][7] ,
         \reg_y[14][6] , \reg_y[14][5] , \reg_y[14][4] , \reg_y[14][3] ,
         \reg_y[14][2] , \reg_y[14][1] , \reg_y[14][0] , \reg_y[13][19] ,
         \reg_y[13][18] , \reg_y[13][17] , \reg_y[13][16] , \reg_y[13][15] ,
         \reg_y[13][14] , \reg_y[13][13] , \reg_y[13][12] , \reg_y[13][11] ,
         \reg_y[13][10] , \reg_y[13][9] , \reg_y[13][8] , \reg_y[13][7] ,
         \reg_y[13][6] , \reg_y[13][5] , \reg_y[13][4] , \reg_y[13][3] ,
         \reg_y[13][2] , \reg_y[13][1] , \reg_y[13][0] , \reg_y[12][19] ,
         \reg_y[12][18] , \reg_y[12][17] , \reg_y[12][16] , \reg_y[12][15] ,
         \reg_y[12][14] , \reg_y[12][13] , \reg_y[12][12] , \reg_y[12][11] ,
         \reg_y[12][10] , \reg_y[12][9] , \reg_y[12][8] , \reg_y[12][7] ,
         \reg_y[12][6] , \reg_y[12][5] , \reg_y[12][4] , \reg_y[12][3] ,
         \reg_y[12][2] , \reg_y[12][1] , \reg_y[12][0] , \reg_y[11][19] ,
         \reg_y[11][18] , \reg_y[11][17] , \reg_y[11][16] , \reg_y[11][15] ,
         \reg_y[11][14] , \reg_y[11][13] , \reg_y[11][12] , \reg_y[11][11] ,
         \reg_y[11][10] , \reg_y[11][9] , \reg_y[11][8] , \reg_y[11][7] ,
         \reg_y[11][6] , \reg_y[11][5] , \reg_y[11][4] , \reg_y[11][3] ,
         \reg_y[11][2] , \reg_y[11][1] , \reg_y[11][0] , \reg_y[10][19] ,
         \reg_y[10][18] , \reg_y[10][17] , \reg_y[10][16] , \reg_y[10][15] ,
         \reg_y[10][14] , \reg_y[10][13] , \reg_y[10][12] , \reg_y[10][11] ,
         \reg_y[10][10] , \reg_y[10][9] , \reg_y[10][8] , \reg_y[10][7] ,
         \reg_y[10][6] , \reg_y[10][5] , \reg_y[10][4] , \reg_y[10][3] ,
         \reg_y[10][2] , \reg_y[10][1] , \reg_y[10][0] , \reg_y[9][19] ,
         \reg_y[9][18] , \reg_y[9][17] , \reg_y[9][16] , \reg_y[9][15] ,
         \reg_y[9][14] , \reg_y[9][13] , \reg_y[9][12] , \reg_y[9][11] ,
         \reg_y[9][10] , \reg_y[9][9] , \reg_y[9][8] , \reg_y[9][7] ,
         \reg_y[9][6] , \reg_y[9][5] , \reg_y[9][4] , \reg_y[9][3] ,
         \reg_y[9][2] , \reg_y[9][1] , \reg_y[9][0] , \reg_y[8][19] ,
         \reg_y[8][18] , \reg_y[8][17] , \reg_y[8][16] , \reg_y[8][15] ,
         \reg_y[8][14] , \reg_y[8][13] , \reg_y[8][12] , \reg_y[8][11] ,
         \reg_y[8][10] , \reg_y[8][9] , \reg_y[8][8] , \reg_y[8][7] ,
         \reg_y[8][6] , \reg_y[8][5] , \reg_y[8][4] , \reg_y[8][3] ,
         \reg_y[8][2] , \reg_y[8][1] , \reg_y[8][0] , \reg_y[7][19] ,
         \reg_y[7][18] , \reg_y[7][17] , \reg_y[7][16] , \reg_y[7][15] ,
         \reg_y[7][14] , \reg_y[7][13] , \reg_y[7][12] , \reg_y[7][11] ,
         \reg_y[7][10] , \reg_y[7][9] , \reg_y[7][8] , \reg_y[7][7] ,
         \reg_y[7][6] , \reg_y[7][5] , \reg_y[7][4] , \reg_y[7][3] ,
         \reg_y[7][2] , \reg_y[7][1] , \reg_y[7][0] , \reg_y[6][19] ,
         \reg_y[6][18] , \reg_y[6][17] , \reg_y[6][16] , \reg_y[6][15] ,
         \reg_y[6][14] , \reg_y[6][13] , \reg_y[6][12] , \reg_y[6][11] ,
         \reg_y[6][10] , \reg_y[6][9] , \reg_y[6][8] , \reg_y[6][7] ,
         \reg_y[6][6] , \reg_y[6][5] , \reg_y[6][4] , \reg_y[6][3] ,
         \reg_y[6][2] , \reg_y[6][1] , \reg_y[6][0] , \reg_y[5][19] ,
         \reg_y[5][18] , \reg_y[5][17] , \reg_y[5][16] , \reg_y[5][15] ,
         \reg_y[5][14] , \reg_y[5][13] , \reg_y[5][12] , \reg_y[5][11] ,
         \reg_y[5][10] , \reg_y[5][9] , \reg_y[5][8] , \reg_y[5][7] ,
         \reg_y[5][6] , \reg_y[5][5] , \reg_y[5][4] , \reg_y[5][3] ,
         \reg_y[5][2] , \reg_y[5][1] , \reg_y[5][0] , \reg_y[4][19] ,
         \reg_y[4][18] , \reg_y[4][17] , \reg_y[4][16] , \reg_y[4][15] ,
         \reg_y[4][14] , \reg_y[4][13] , \reg_y[4][12] , \reg_y[4][11] ,
         \reg_y[4][10] , \reg_y[4][9] , \reg_y[4][8] , \reg_y[4][7] ,
         \reg_y[4][6] , \reg_y[4][5] , \reg_y[4][4] , \reg_y[4][3] ,
         \reg_y[4][2] , \reg_y[4][1] , \reg_y[4][0] , \reg_y[3][19] ,
         \reg_y[3][18] , \reg_y[3][17] , \reg_y[3][16] , \reg_y[3][15] ,
         \reg_y[3][14] , \reg_y[3][13] , \reg_y[3][12] , \reg_y[3][11] ,
         \reg_y[3][10] , \reg_y[3][9] , \reg_y[3][8] , \reg_y[3][7] ,
         \reg_y[3][6] , \reg_y[3][5] , \reg_y[3][4] , \reg_y[3][3] ,
         \reg_y[3][2] , \reg_y[3][1] , \reg_y[3][0] , \reg_y[2][19] ,
         \reg_y[2][18] , \reg_y[2][17] , \reg_y[2][16] , \reg_y[2][15] ,
         \reg_y[2][14] , \reg_y[2][13] , \reg_y[2][12] , \reg_y[2][11] ,
         \reg_y[2][10] , \reg_y[2][9] , \reg_y[2][8] , \reg_y[2][7] ,
         \reg_y[2][6] , \reg_y[2][5] , \reg_y[2][4] , \reg_y[2][3] ,
         \reg_y[2][2] , \reg_y[2][1] , \reg_y[2][0] , \reg_y[1][19] ,
         \reg_y[1][18] , \reg_y[1][17] , \reg_y[1][16] , \reg_y[1][15] ,
         \reg_y[1][14] , \reg_y[1][13] , \reg_y[1][12] , \reg_y[1][11] ,
         \reg_y[1][10] , \reg_y[1][9] , \reg_y[1][8] , \reg_y[1][7] ,
         \reg_y[1][6] , \reg_y[1][5] , \reg_y[1][4] , \reg_y[1][3] ,
         \reg_y[1][2] , \reg_y[1][1] , \reg_y[1][0] , \reg_y[0][19] ,
         \reg_y[0][18] , \reg_y[0][17] , \reg_y[0][16] , \reg_y[0][15] ,
         \reg_y[0][14] , \reg_y[0][13] , \reg_y[0][12] , \reg_y[0][11] ,
         \reg_y[0][10] , \reg_y[0][9] , \reg_y[0][8] , \reg_y[0][7] ,
         \reg_y[0][6] , \reg_y[0][5] , \reg_y[0][4] , \reg_y[0][3] ,
         \reg_y[0][2] , \reg_y[0][1] , \reg_y[0][0] , reg_model, n1353, n1354,
         n1355, n1356, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
         n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
         n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
         n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
         n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
         n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
         n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
         n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
         n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
         n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
         n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
         n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
         n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
         n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
         n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
         n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
         n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
         n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
         n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
         n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
         n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
         n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
         n1995, n1996, n1997, n1998, n1999, n36862, n36863, n36864, n36865,
         n36866, n36867, n36868, n36869, n36870, n36871, n36872, n36873,
         n36874, n36875, n36876, n36877, n36878, n36879, n36880, n36881,
         n36882, n36883, n36884, n36885, n36886, n36887, n36888, n36889,
         n36890, n36891, n36892, n36893, n36894, n36895, n36896, n36897,
         n36898, n36899, n36900, n36901, n36902, n36903, n36904, n36905,
         n36906, n36908, n36909, n36910, n36912, n36913, n36914, n36915,
         n36916, n36917, n36918, n36919, n36920, n36921, n36922, n36923,
         n36924, n36925, n36926, n36927, n36928, n36929, n36930, n36931,
         n36932, n36933, n36934, n36935, n36936, n36937, n36938, n36939,
         n36940, n36941, n36942, n36943, n36944, n36945, n36946, n36947,
         n36948, n36949, n36950, n36951, n36952, n36953, n36954, n36955,
         n36956, n36957, n36958, n36959, n36960, n36961, n36962, n36963,
         n36964, n36965, n36966, n36967, n36968, n36969, n36970, n36971,
         n36972, n36973, n36974, n36975, n36976, n36977, n36978, n36979,
         n36980, n36981, n36982, n36983, n36984, n36985, n36986, n36987,
         n36988, n36989, n36990, n36991, n36992, n36993, n36994, n36995,
         n36996, n36997, n36998, n36999, n37000, n37001, n37002, n37003,
         n37004, n37005, n37006, n37007, n37008, n37009, n37010, n37011,
         n37012, n37013, n37014, n37015, n37016, n37017, n37018, n37019,
         n37020, n37021, n37022, n37023, n37024, n37025, n37026, n37027,
         n37028, n37029, n37030, n37031, n37032, n37033, n37034, n37035,
         n37036, n37037, n37038, n37039, n37040, n37041, n37042, n37043,
         n37044, n37045, n37046, n37047, n37048, n37049, n37050, n37051,
         n37052, n37053, n37054, n37055, n37056, n37057, n37058, n37059,
         n37060, n37061, n37062, n37063, n37064, n37065, n37066, n37067,
         n37068, n37069, n37070, n37071, n37072, n37073, n37074, n37075,
         n37076, n37077, n37078, n37079, n37080, n37081, n37082, n37083,
         n37084, n37085, n37086, n37087, n37088, n37089, n37090, n37091,
         n37092, n37093, n37094, n37095, n37096, n37097, n37098, n37099,
         n37100, n37101, n37102, n37103, n37104, n37105, n37106, n37107,
         n37108, n37109, n37110, n37111, n37112, n37113, n37114, n37115,
         n37116, n37117, n37118, n37119, n37120, n37121, n37122, n37123,
         n37124, n37125, n37126, n37127, n37128, n37129, n37130, n37131,
         n37132, n37133, n37134, n37135, n37136, n37137, n37138, n37139,
         n37140, n37141, n37142, n37143, n37144, n37145, n37146, n37147,
         n37148, n37149, n37150, n37151, n37152, n37153, n37154, n37155,
         n37156, n37157, n37158, n37159, n37160, n37161, n37162, n37163,
         n37164, n37165, n37166, n37167, n37168, n37169, n37170, n37171,
         n37172, n37173, n37174, n37175, n37176, n37177, n37178, n37179,
         n37180, n37181, n37182, n37183, n37184, n37185, n37186, n37187,
         n37188, n37189, n37190, n37191, n37192, n37193, n37194, n37195,
         n37196, n37197, n37198, n37199, n37200, n37201, n37202, n37203,
         n37204, n37205, n37206, n37207, n37208, n37209, n37210, n37211,
         n37212, n37213, n37214, n37215, n37216, n37217, n37218, n37219,
         n37220, n37221, n37222, n37223, n37224, n37225, n37226, n37227,
         n37228, n37229, n37230, n37231, n37232, n37233, n37234, n37235,
         n37236, n37237, n37238, n37239, n37240, n37241, n37242, n37243,
         n37244, n37245, n37246, n37247, n37248, n37249, n37250, n37251,
         n37252, n37253, n37254, n37255, n37256, n37257, n37258, n37259,
         n37260, n37261, n37262, n37263, n37264, n37265, n37266, n37267,
         n37268, n37269, n37270, n37271, n37272, n37273, n37274, n37275,
         n37276, n37277, n37278, n37279, n37280, n37281, n37282, n37283,
         n37284, n37285, n37286, n37287, n37288, n37289, n37290, n37291,
         n37292, n37293, n37294, n37295, n37296, n37297, n37298, n37299,
         n37300, n37301, n37302, n37303, n37304, n37305, n37306, n37307,
         n37308, n37309, n37310, n37311, n37312, n37313, n37314, n37315,
         n37316, n37317, n37318, n37319, n37320, n37321, n37322, n37323,
         n37324, n37325, n37326, n37327, n37328, n37329, n37330, n37331,
         n37332, n37333, n37334, n37335, n37336, n37337, n37338, n37339,
         n37340, n37341, n37342, n37343, n37344, n37345, n37346, n37347,
         n37348, n37349, n37350, n37351, n37352, n37353, n37354, n37355,
         n37356, n37357, n37358, n37359, n37360, n37361, n37362, n37363,
         n37364, n37365, n37366, n37367, n37368, n37369, n37370, n37371,
         n37372, n37373, n37374, n37375, n37376, n37377, n37378, n37379,
         n37380, n37381, n37382, n37383, n37384, n37385, n37386, n37387,
         n37388, n37389, n37390, n37391, n37392, n37393, n37394, n37395,
         n37396, n37397, n37398, n37399, n37400, n37401, n37402, n37403,
         n37404, n37405, n37406, n37407, n37408, n37409, n37410, n37411,
         n37412, n37413, n37414, n37415, n37416, n37417, n37418, n37419,
         n37420, n37421, n37422, n37423, n37424, n37425, n37426, n37427,
         n37428, n37429, n37430, n37431, n37432, n37433, n37434, n37435,
         n37436, n37437, n37438, n37439, n37440, n37441, n37442, n37443,
         n37444, n37445, n37446, n37447, n37448, n37449, n37450, n37451,
         n37452, n37453, n37454, n37455, n37456, n37457, n37458, n37459,
         n37460, n37461, n37462, n37463, n37464, n37465, n37466, n37467,
         n37468, n37469, n37470, n37471, n37472, n37473, n37474, n37475,
         n37476, n37477, n37478, n37479, n37480, n37481, n37482, n37483,
         n37484, n37485, n37486, n37487, n37488, n37489, n37490, n37491,
         n37492, n37493, n37494, n37495, n37496, n37497, n37498, n37499,
         n37500, n37501, n37502, n37503, n37504, n37505, n37506, n37507,
         n37508, n37509, n37510, n37511, n37512, n37513, n37514, n37515,
         n37516, n37517, n37518, n37519, n37520, n37521, n37522, n37523,
         n37524, n37525, n37526, n37527, n37528, n37529, n37530, n37531,
         n37532, n37533, n37534, n37535, n37536, n37537, n37538, n37539,
         n37540, n37541, n37542, n37543, n37544, n37545, n37546, n37547,
         n37548, n37549, n37550, n37551, n37552, n37553, n37554, n37555,
         n37556, n37557, n37558, n37559, n37560, n37561, n37562, n37563,
         n37564, n37565, n37566, n37567, n37568, n37569, n37570, n37571,
         n37572, n37573, n37574, n37575, n37576, n37577, n37578, n37579,
         n37580, n37581, n37582, n37583, n37584, n37585, n37586, n37587,
         n37588, n37589, n37590, n37591, n37592, n37593, n37594, n37595,
         n37596, n37597, n37598, n37599, n37600, n37601, n37602, n37603,
         n37604, n37605, n37606, n37607, n37608, n37609, n37610, n37611,
         n37612, n37613, n37614, n37615, n37616, n37617, n37618, n37619,
         n37620, n37621, n37622, n37623, n37624, n37625, n37626, n37627,
         n37628, n37629, n37630, n37631, n37632, n37633, n37634, n37635,
         n37636, n37637, n37638, n37639, n37640, n37641, n37642, n37643,
         n37644, n37645, n37646, n37647, n37648, n37649, n37650, n37651,
         n37652, n37653, n37654, n37655, n37656, n37657, n37658, n37659,
         n37660, n37661, n37662, n37663, n37664, n37665, n37666, n37667,
         n37668, n37669, n37670, n37671, n37672, n37673, n37674, n37675,
         n37676, n37677, n37678, n37679, n37680, n37681, n37682, n37683,
         n37684, n37685, n37686, n37687, n37688, n37689, n37690, n37691,
         n37692, n37693, n37694, n37695, n37696, n37697, n37698, n37699,
         n37700, n37701, n37702, n37703, n37704, n37705, n37706, n37707,
         n37708, n37709, n37710, n37711, n37712, n37713, n37714, n37715,
         n37716, n37717, n37718, n37719, n37720, n37721, n37722, n37723,
         n37724, n37725, n37726, n37727, n37728, n37729, n37730, n37731,
         n37732, n37733, n37734, n37735, n37736, n37737, n37738, n37739,
         n37740, n37741, n37742, n37743, n37744, n37745, n37746, n37747,
         n37748, n37749, n37750, n37751, n37752, n37753, n37754, n37755,
         n37756, n37757, n37758, n37759, n37760, n37761, n37762, n37763,
         n37764, n37765, n37766, n37767, n37768, n37769, n37770, n37771,
         n37772, n37773, n37774, n37775, n37776, n37777, n37778, n37779,
         n37780, n37781, n37782, n37783, n37784, n37785, n37786, n37787,
         n37788, n37789, n37790, n37791, n37792, n37793, n37794, n37795,
         n37796, n37797, n37798, n37799, n37800, n37801, n37802, n37803,
         n37804, n37805, n37806, n37807, n37808, n37809, n37810, n37811,
         n37812, n37813, n37814, n37815, n37816, n37817, n37818, n37819,
         n37820, n37821, n37822, n37823, n37824, n37825, n37826, n37827,
         n37828, n37829, n37830, n37831, n37832, n37833, n37834, n37835,
         n37836, n37837, n37838, n37839, n37840, n37841, n37842, n37843,
         n37844, n37845, n37846, n37847, n37848, n37849, n37850, n37851,
         n37852, n37853, n37854, n37855, n37856, n37857, n37858, n37859,
         n37860, n37861, n37862, n37863, n37864, n37865, n37866, n37867,
         n37868, n37869, n37870, n37871, n37872, n37873, n37874, n37875,
         n37876, n37877, n37878, n37879, n37880, n37881, n37882, n37883,
         n37884, n37885, n37886, n37887, n37888, n37889, n37890, n37891,
         n37892, n37893, n37894, n37895, n37896, n37897, n37898, n37899,
         n37900, n37901, n37902, n37903, n37904, n37905, n37906, n37907,
         n37908, n37909, n37910, n37911, n37912, n37913, n37914, n37915,
         n37916, n37917, n37918, n37919, n37920, n37921, n37922, n37923,
         n37924, n37925, n37926, n37927, n37928, n37929, n37930, n37931,
         n37932, n37933, n37934, n37935, n37936, n37937, n37938, n37939,
         n37940, n37941, n37942, n37943, n37944, n37945, n37946, n37947,
         n37948, n37949, n37950, n37951, n37952, n37953, n37954, n37955,
         n37956, n37957, n37958, n37959, n37960, n37961, n37962, n37963,
         n37964, n37965, n37966, n37967, n37968, n37969, n37970, n37971,
         n37972, n37973, n37974, n37975, n37976, n37977, n37978, n37979,
         n37980, n37981, n37982, n37983, n37984, n37985, n37986, n37987,
         n37988, n37989, n37990, n37991, n37992, n37993, n37994, n37995,
         n37996, n37997, n37998, n37999, n38000, n38001, n38002, n38003,
         n38004, n38005, n38006, n38007, n38008, n38009, n38010, n38011,
         n38012, n38013, n38014, n38015, n38016, n38017, n38018, n38019,
         n38020, n38021, n38022, n38023, n38024, n38025, n38026, n38027,
         n38028, n38029, n38030, n38031, n38032, n38033, n38034, n38035,
         n38036, n38037, n38038, n38039, n38040, n38041, n38042, n38043,
         n38044, n38045, n38046, n38047, n38048, n38049, n38050, n38051,
         n38052, n38053, n38054, n38055, n38056, n38057, n38058, n38059,
         n38060, n38061, n38062, n38063, n38064, n38065, n38066, n38067,
         n38068, n38069, n38070, n38071, n38072, n38073, n38074, n38075,
         n38076, n38077, n38078, n38079, n38080, n38081, n38082, n38083,
         n38084, n38085, n38086, n38087, n38088, n38089, n38090, n38091,
         n38092, n38093, n38094, n38095, n38096, n38097, n38098, n38099,
         n38100, n38101, n38102, n38103, n38104, n38105, n38106, n38107,
         n38108, n38109, n38110, n38111, n38112, n38113, n38114, n38115,
         n38116, n38117, n38118, n38119, n38120, n9999, n9998, n9997, n9996,
         n9995, n9994, n9993, n9992, n9991, n9990, n9989, n9988, n9987, n9986,
         n9985, n9984, n9983, n9982, n9981, n9980, n9979, n9978, n9977, n9976,
         n9975, n9974, n9973, n9972, n9971, n9970, n9969, n9968, n9967, n9966,
         n9965, n9964, n9963, n9962, n9961, n9960, n9959, n9958, n9957, n9956,
         n9955, n9954, n9953, n9952, n9951, n9950, n9949, n9948, n9947, n9946,
         n9945, n9944, n9943, n9942, n9941, n9940, n9939, n9938, n9937, n9936,
         n9935, n9934, n9933, n9932, n9931, n9930, n9929, n9928, n9927, n9926,
         n9925, n9924, n9923, n9922, n9921, n9920, n9919, n9918, n9917, n9916,
         n9915, n9914, n9913, n9912, n9911, n9910, n9909, n9908, n9907, n9906,
         n9905, n9904, n9903, n9902, n9900, n9899, n9898, n9897, n9896, n9895,
         n9894, n9893, n9892, n9891, n9890, n9889, n9888, n9887, n9886, n9885,
         n9884, n9883, n9882, n9881, n9880, n9879, n9878, n9877, n9876, n9875,
         n9874, n9873, n9872, n9871, n9870, n9869, n9868, n9867, n9866, n9865,
         n9864, n9863, n9862, n9861, n9860, n9859, n9858, n9857, n9856, n9855,
         n9854, n9853, n9852, n9851, n9850, n9849, n9848, n9847, n9846, n9845,
         n9844, n9843, n9842, n9841, n9840, n9839, n9838, n9837, n9836, n9835,
         n9834, n9833, n9832, n9831, n9830, n9829, n9828, n9827, n9826, n9825,
         n9824, n9823, n9822, n9821, n9820, n9819, n9818, n9817, n9816, n9815,
         n9814, n9813, n9812, n9811, n9810, n9809, n9808, n9807, n9806, n9805,
         n9804, n9802, n9801, n9800, n9799, n9798, n9797, n9796, n9795, n9794,
         n9793, n9792, n9791, n9790, n9789, n9788, n9787, n9786, n9785, n9784,
         n9783, n9782, n9781, n9780, n9779, n9778, n9777, n9776, n9775, n9774,
         n9773, n9772, n9771, n9770, n9769, n9768, n9767, n9766, n9765, n9764,
         n9763, n9762, n9761, n9760, n9759, n9758, n9757, n9756, n9755, n9754,
         n9753, n9752, n9751, n9750, n9749, n9748, n9747, n9746, n9745, n9744,
         n9743, n9742, n9741, n9740, n9739, n9738, n9737, n9736, n9735, n9734,
         n9733, n9732, n9731, n9730, n9729, n9728, n9727, n9726, n9725, n9724,
         n9723, n9722, n9721, n9720, n9719, n9718, n9717, n9716, n9715, n9714,
         n9713, n9712, n9711, n9710, n9709, n9708, n9707, n9706, n9705, n9704,
         n9703, n9702, n9701, n9700, n9699, n9698, n9697, n9696, n9695, n9694,
         n9693, n9692, n9691, n9690, n9689, n9688, n9687, n9686, n9685, n9684,
         n9683, n9682, n9681, n9680, n9679, n9678, n9677, n9676, n9675, n9674,
         n9673, n9672, n9671, n9670, n9669, n9668, n9667, n9666, n9665, n9664,
         n9663, n9662, n9661, n9660, n9659, n9658, n9657, n9656, n9655, n9654,
         n9653, n9652, n9651, n9650, n9649, n9648, n9647, n9646, n9645, n9644,
         n9643, n9642, n9641, n9640, n9639, n9638, n9637, n9636, n9635, n9634,
         n9633, n9632, n9631, n9630, n9629, n9628, n9627, n9626, n9625, n9624,
         n9623, n9622, n9621, n9620, n9619, n9618, n9617, n9616, n9615, n9614,
         n9613, n9612, n9611, n9609, n9608, n9607, n9606, n9605, n9604, n9603,
         n9602, n9601, n9600, n9599, n9598, n9597, n9596, n9595, n9594, n9593,
         n9592, n9591, n9590, n9589, n9588, n9587, n9586, n9585, n9584, n9583,
         n9582, n9581, n9580, n9579, n9578, n9577, n9576, n9575, n9574, n9573,
         n9572, n9571, n9570, n9569, n9568, n9567, n9566, n9565, n9564, n9563,
         n9562, n9561, n9560, n9559, n9558, n9557, n9556, n9555, n9554, n9553,
         n9552, n9551, n9550, n9549, n9548, n9547, n9546, n9545, n9544, n9543,
         n9542, n9541, n9540, n9539, n9538, n9537, n9536, n9535, n9534, n9533,
         n9532, n9531, n9530, n9529, n9528, n9527, n9526, n9525, n9524, n9523,
         n9522, n9521, n9520, n9519, n9518, n9517, n9516, n9515, n9514, n9513,
         n9512, n9511, n9510, n9509, n9508, n9507, n9506, n9505, n9504, n9503,
         n9502, n9501, n9500, n9499, n9498, n9497, n9496, n9495, n9494, n9493,
         n9491, n9490, n9489, n9488, n9487, n9486, n9485, n9484, n9483, n9482,
         n9481, n9480, n9479, n9478, n9477, n9476, n9475, n9474, n9473, n9472,
         n9471, n9470, n9469, n9468, n9467, n9466, n9465, n9464, n9463, n9462,
         n9461, n9460, n9459, n9458, n9457, n9456, n9455, n9454, n9452, n9451,
         n9450, n9449, n9448, n9447, n9445, n9444, n9443, n9442, n9441, n9440,
         n9439, n9438, n9437, n9436, n9435, n9434, n9433, n9432, n9431, n9430,
         n9429, n9428, n9427, n9425, n9424, n9423, n9422, n9421, n9420, n9419,
         n9418, n9417, n9416, n9415, n9414, n9413, n9412, n9411, n9410, n9409,
         n9408, n9407, n9406, n9405, n9404, n9403, n9402, n9400, n9399, n9398,
         n9397, n9396, n9395, n9394, n9393, n9392, n9391, n9390, n9389, n9388,
         n9387, n9386, n9385, n9384, n9383, n9382, n9381, n9380, n9379, n9378,
         n9377, n9376, n9375, n9374, n9373, n9372, n9371, n9370, n9369, n9368,
         n9367, n9366, n9365, n9364, n9363, n9362, n9361, n9360, n9359, n9358,
         n9357, n9356, n9355, n9354, n9353, n9352, n9351, n9350, n9349, n9348,
         n9347, n9346, n9345, n9344, n9343, n9342, n9341, n9340, n9339, n9338,
         n9337, n9336, n9335, n9334, n9333, n9332, n9331, n9330, n9329, n9328,
         n9327, n9326, n9325, n9324, n9323, n9322, n9321, n9320, n9319, n9318,
         n9317, n9316, n9315, n9314, n9313, n9312, n9311, n9310, n9309, n9308,
         n9307, n9306, n9305, n9304, n9303, n9302, n9301, n9300, n9299, n9298,
         n9297, n9296, n9295, n9294, n9293, n9292, n9291, n9290, n9289, n9288,
         n9287, n9286, n9285, n9284, n9283, n9282, n9280, n9279, n9278, n9277,
         n9276, n9275, n9274, n9273, n9272, n9271, n9270, n9269, n9268, n9267,
         n9266, n9265, n9264, n9263, n9262, n9261, n9260, n9259, n9258, n9257,
         n9256, n9255, n9254, n9253, n9252, n9251, n9250, n9249, n9248, n9247,
         n9246, n9245, n9244, n9243, n9242, n9241, n9240, n9239, n9238, n9237,
         n9236, n9235, n9234, n9233, n9232, n9231, n9230, n9229, n9228, n9227,
         n9226, n9225, n9224, n9223, n9222, n9221, n9220, n9219, n9218, n9217,
         n9216, n9215, n9214, n9213, n9212, n9211, n9210, n9209, n9208, n9207,
         n9206, n9205, n9204, n9203, n9202, n9201, n9200, n9199, n9198, n9197,
         n9196, n9195, n9194, n9193, n9192, n9191, n9190, n9189, n9188, n9187,
         n9186, n9185, n9184, n9183, n9182, n9181, n9180, n9179, n9178, n9177,
         n9176, n9175, n9174, n9173, n9172, n9171, n9170, n9169, n9168, n9167,
         n9166, n9165, n9164, n9163, n9162, n9161, n9160, n9159, n9158, n9157,
         n9156, n9155, n9154, n9153, n9152, n9151, n9150, n9149, n9148, n9147,
         n9146, n9145, n9144, n9143, n9142, n9141, n9140, n9139, n9138, n9137,
         n9136, n9135, n9134, n9133, n9132, n9131, n9130, n9129, n9128, n9127,
         n9126, n9125, n9124, n9123, n9122, n9121, n9120, n9119, n9118, n9117,
         n9116, n9115, n9114, n9113, n9112, n9111, n9110, n9109, n9108, n9107,
         n9106, n9105, n9104, n9103, n9102, n9101, n9100, n9099, n9098, n9097,
         n9096, n9095, n9094, n9093, n9092, n9091, n9090, n9089, n9088, n9087,
         n9086, n9085, n9084, n9083, n9082, n9081, n9080, n9079, n9078, n9077,
         n9076, n9075, n9074, n9073, n9072, n9071, n9070, n9069, n9068, n9067,
         n9066, n9065, n9064, n9063, n9062, n9061, n9060, n9059, n9058, n9057,
         n9056, n9055, n9054, n9053, n9052, n9051, n9050, n9049, n9048, n9047,
         n9046, n9045, n9044, n9043, n9042, n9041, n9040, n9039, n9038, n9037,
         n9036, n9035, n9034, n9033, n9032, n9031, n9030, n9029, n9028, n9027,
         n9026, n9025, n9024, n9023, n9022, n9021, n9020, n9019, n9018, n9017,
         n9016, n9015, n9014, n9013, n9012, n9011, n9010, n9009, n9008, n9007,
         n9006, n9005, n9004, n9003, n9002, n9001, n9000, n8999, n8998, n8997,
         n8996, n8995, n8994, n8993, n8992, n8991, n8990, n8989, n8988, n8987,
         n8986, n8985, n8984, n8982, n8981, n8980, n8979, n8978, n8977, n8976,
         n8975, n8974, n8973, n8972, n8971, n8970, n8969, n8968, n8967, n8966,
         n8965, n8964, n8963, n8962, n8961, n8960, n8959, n8958, n8957, n8956,
         n8955, n8954, n8953, n8952, n8951, n8950, n8949, n8948, n8947, n8946,
         n8945, n8944, n8943, n8942, n8941, n8940, n8939, n8938, n8937, n8936,
         n8935, n8934, n8933, n8932, n8931, n8930, n8929, n8928, n8927, n8926,
         n8925, n8924, n8923, n8922, n8921, n8920, n8919, n8918, n8917, n8916,
         n8915, n8914, n8913, n8912, n8911, n8910, n8909, n8908, n8907, n8906,
         n8905, n8904, n8903, n8902, n8901, n8900, n8899, n8898, n8897, n8896,
         n8895, n8894, n8893, n8892, n8891, n8890, n8889, n8888, n8887, n8886,
         n8885, n8884, n8883, n8882, n8881, n8880, n8879, n8878, n8877, n8876,
         n8875, n8874, n8873, n8872, n8871, n8870, n8869, n8868, n8867, n8866,
         n8865, n8864, n8863, n8862, n8861, n8860, n8859, n8858, n8857, n8856,
         n8855, n8854, n8853, n8852, n8851, n8850, n8849, n8848, n8847, n8846,
         n8845, n8844, n8843, n8842, n8841, n8840, n8839, n8838, n8837, n8836,
         n8835, n8834, n8833, n8832, n8831, n8830, n8829, n8828, n8827, n8826,
         n8825, n8824, n8823, n8822, n8821, n8820, n8819, n8818, n8817, n8816,
         n8815, n8814, n8813, n8812, n8811, n8810, n8809, n8808, n8807, n8806,
         n8805, n8804, n8803, n8802, n8801, n8800, n8799, n8798, n8797, n8796,
         n8795, n8794, n8793, n8792, n8791, n8789, n8788, n8787, n8786, n8785,
         n8784, n8783, n8782, n8781, n8780, n8779, n8778, n8777, n8776, n8775,
         n8774, n8773, n8772, n8771, n8770, n8769, n8768, n8767, n8766, n8765,
         n8764, n8763, n8762, n8761, n8760, n8759, n8758, n8757, n8756, n8755,
         n8754, n8753, n8752, n8751, n8750, n8749, n8748, n8747, n8746, n8745,
         n8744, n8743, n8742, n8741, n8740, n8739, n8738, n8737, n8736, n8735,
         n8734, n8733, n8732, n8731, n8730, n8729, n8728, n8727, n8726, n8725,
         n8724, n8723, n8722, n8721, n8720, n8718, n8717, n8716, n8715, n8714,
         n8713, n8712, n8711, n8710, n8709, n8708, n8707, n8706, n8705, n8704,
         n8703, n8702, n8701, n8700, n8699, n8698, n8697, n8696, n8695, n8694,
         n8693, n8692, n8691, n8690, n8689, n8688, n8687, n8686, n8685, n8684,
         n8683, n8682, n8681, n8680, n8679, n8678, n8677, n8676, n8675, n8674,
         n8673, n8671, n8670, n8669, n8668, n8667, n8666, n8665, n8664, n8663,
         n8662, n8661, n8660, n8659, n8658, n8657, n8656, n8655, n8654, n8653,
         n8652, n8651, n8650, n8649, n8648, n8647, n8646, n8645, n8644, n8643,
         n8642, n8641, n8640, n8639, n8638, n8637, n8636, n8635, n8634, n8632,
         n8631, n8630, n8629, n8628, n8627, n8625, n8624, n8623, n8622, n8621,
         n8620, n8619, n8618, n8617, n8616, n8615, n8614, n8613, n8612, n8611,
         n8610, n8609, n8608, n8607, n8605, n8604, n8603, n8602, n8601, n8600,
         n8599, n8598, n8597, n8596, n8595, n8594, n8593, n8592, n8591, n8590,
         n8589, n8588, n8587, n8586, n8585, n8584, n8583, n8582, n8580, n8579,
         n8578, n8577, n8576, n8575, n8574, n8573, n8572, n8571, n8570, n8569,
         n8568, n8567, n8566, n8565, n8564, n8563, n8562, n8561, n8560, n8559,
         n8558, n8557, n8556, n8555, n8554, n8553, n8552, n8551, n8550, n8549,
         n8548, n8547, n8546, n8545, n8544, n8543, n8542, n8541, n8540, n8539,
         n8538, n8537, n8536, n8535, n8534, n8533, n8532, n8531, n8530, n8529,
         n8528, n8527, n8526, n8525, n8524, n8523, n8522, n8521, n8520, n8519,
         n8518, n8517, n8516, n8515, n8514, n8513, n8512, n8511, n8510, n8509,
         n8508, n8507, n8506, n8505, n8504, n8503, n8502, n8501, n8500, n8499,
         n8498, n8497, n8496, n8495, n8494, n8493, n8492, n8491, n8490, n8489,
         n8488, n8487, n8486, n8485, n8484, n8483, n8482, n8481, n8480, n8479,
         n8478, n8477, n8476, n8475, n8474, n8473, n8472, n8471, n8470, n8469,
         n8468, n8467, n8466, n8465, n8464, n8463, n8462, n8460, n8459, n8458,
         n8457, n8456, n8455, n8454, n8453, n8452, n8451, n8450, n8449, n8448,
         n8447, n8446, n8445, n8444, n8443, n8442, n8441, n8440, n8439, n8438,
         n8437, n8436, n8435, n8434, n8433, n8432, n8431, n8430, n8429, n8428,
         n8427, n8426, n8425, n8424, n8423, n8422, n8421, n8420, n8419, n8418,
         n8417, n8416, n8415, n8414, n8413, n8412, n8411, n8410, n8409, n8408,
         n8407, n8406, n8405, n8404, n8403, n8402, n8401, n8400, n8399, n8398,
         n8397, n8396, n8395, n8394, n8393, n8392, n8391, n8390, n8389, n8388,
         n8387, n8386, n8385, n8384, n8383, n8382, n8381, n8380, n8379, n8378,
         n8377, n8376, n8375, n8374, n8373, n8372, n8371, n8370, n8369, n8368,
         n8367, n8366, n8365, n8364, n8363, n8362, n8361, n8360, n8359, n8358,
         n8357, n8356, n8355, n8354, n8353, n8352, n8351, n8350, n8349, n8348,
         n8347, n8346, n8345, n8344, n8343, n8342, n8341, n8340, n8339, n8338,
         n8337, n8336, n8335, n8334, n8333, n8332, n8331, n8330, n8329, n8328,
         n8327, n8326, n8325, n8324, n8323, n8322, n8321, n8320, n8319, n8318,
         n8317, n8316, n8315, n8314, n8313, n8312, n8311, n8310, n8309, n8308,
         n8307, n8306, n8305, n8304, n8303, n8302, n8301, n8300, n8299, n8298,
         n8297, n8296, n8295, n8294, n8293, n8292, n8291, n8290, n8289, n8288,
         n8287, n8286, n8285, n8284, n8283, n8282, n8281, n8280, n8279, n8278,
         n8277, n8276, n8275, n8274, n8273, n8272, n8271, n8270, n8269, n8268,
         n8267, n8266, n8265, n8264, n8262, n8261, n8260, n8259, n8258, n8257,
         n8256, n8255, n8254, n8253, n8252, n8251, n8250, n8249, n8248, n8247,
         n8246, n8245, n8244, n8243, n8242, n8241, n8240, n8239, n8238, n8237,
         n8236, n8235, n8234, n8233, n8232, n8231, n8230, n8229, n8228, n8227,
         n8226, n8225, n8224, n8223, n8222, n8221, n8220, n8219, n8218, n8217,
         n8216, n8215, n8214, n8213, n8212, n8211, n8210, n8209, n8208, n8207,
         n8206, n8205, n8204, n8203, n8202, n8201, n8200, n8199, n8198, n8197,
         n8196, n8195, n8194, n8193, n8192, n8191, n8190, n8189, n8188, n8187,
         n8186, n8185, n8184, n8183, n8182, n8181, n8180, n8179, n8178, n8177,
         n8176, n8175, n8174, n8173, n8172, n8171, n8170, n8169, n8168, n8167,
         n8166, n8164, n8163, n8162, n8161, n8160, n8159, n8158, n8157, n8156,
         n8155, n8154, n8153, n8152, n8151, n8150, n8149, n8148, n8147, n8146,
         n8145, n8144, n8143, n8142, n8141, n8140, n8139, n8138, n8137, n8136,
         n8135, n8134, n8133, n8132, n8131, n8130, n8129, n8128, n8127, n8126,
         n8125, n8124, n8123, n8122, n8121, n8120, n8119, n8117, n8116, n8115,
         n8114, n8113, n8112, n8111, n8110, n8109, n8108, n8107, n8106, n8105,
         n8104, n8103, n8102, n8101, n8100, n8099, n8098, n8097, n8096, n8095,
         n8094, n8093, n8092, n8091, n8090, n8089, n8088, n8087, n8086, n8085,
         n8084, n8083, n8082, n8081, n8080, n8079, n8078, n8077, n8076, n8075,
         n8074, n8073, n8072, n8071, n8070, n8069, n8068, n8067, n8066, n8065,
         n8064, n8063, n8062, n8061, n8060, n8059, n8058, n8057, n8056, n8055,
         n8054, n8053, n8052, n8051, n8050, n8049, n8048, n8047, n8046, n8045,
         n8044, n8043, n8042, n8041, n8040, n8039, n8038, n8037, n8036, n8035,
         n8034, n8033, n8032, n8031, n8030, n8029, n8028, n8027, n8026, n8025,
         n8024, n8023, n8022, n8021, n8020, n8019, n8018, n8017, n8016, n8015,
         n8014, n8013, n8012, n8011, n8010, n8009, n8008, n8007, n8006, n8005,
         n8004, n8003, n8002, n8001, n8000, n7999, n7998, n7997, n7996, n7995,
         n7994, n7993, n7992, n7991, n7990, n7989, n7988, n7987, n7986, n7985,
         n7984, n7983, n7982, n7981, n7980, n7979, n7978, n7977, n7976, n7975,
         n7974, n7973, n7971, n7970, n7969, n7968, n7967, n7966, n7965, n7964,
         n7963, n7962, n7961, n7960, n7959, n7958, n7957, n7956, n7955, n7954,
         n7953, n7952, n7951, n7950, n7949, n7948, n7947, n7946, n7945, n7944,
         n7943, n7942, n7941, n7940, n7939, n7938, n7937, n7936, n7935, n7934,
         n7933, n7932, n7931, n7930, n7929, n7928, n7927, n7926, n7925, n7924,
         n7923, n7922, n7921, n7920, n7919, n7918, n7917, n7916, n7915, n7914,
         n7913, n7912, n7911, n7910, n7909, n7908, n7907, n7906, n7905, n7904,
         n7903, n7902, n7900, n7899, n7898, n7897, n7896, n7895, n7894, n7893,
         n7892, n7891, n7890, n7889, n7888, n7887, n7886, n7885, n7884, n7883,
         n7882, n7881, n7880, n7879, n7878, n7877, n7876, n7875, n7874, n7873,
         n7872, n7871, n7870, n7869, n7868, n7867, n7866, n7865, n7864, n7863,
         n7862, n7861, n7860, n7859, n7858, n7857, n7856, n7855, n7853, n7852,
         n7851, n7850, n7849, n7848, n7847, n7846, n7845, n7844, n7843, n7842,
         n7841, n7840, n7839, n7838, n7837, n7836, n7835, n7834, n7833, n7832,
         n7831, n7830, n7829, n7828, n7827, n7826, n7825, n7824, n7823, n7822,
         n7821, n7820, n7819, n7818, n7817, n7816, n7814, n7813, n7812, n7811,
         n7810, n7809, n7807, n7806, n7805, n7804, n7803, n7802, n7801, n7800,
         n7799, n7798, n7797, n7796, n7795, n7794, n7793, n7792, n7791, n7790,
         n7789, n7787, n7786, n7785, n7784, n7783, n7782, n7781, n7780, n7779,
         n7778, n7777, n7776, n7775, n7774, n7773, n7772, n7771, n7770, n7769,
         n7768, n7767, n7766, n7765, n7764, n7762, n7761, n7760, n7759, n7758,
         n7757, n7756, n7755, n7754, n7753, n7752, n7751, n7750, n7749, n7748,
         n7747, n7746, n7745, n7744, n7743, n7742, n7741, n7740, n7739, n7738,
         n7737, n7736, n7735, n7734, n7733, n7732, n7731, n7730, n7729, n7728,
         n7727, n7726, n7725, n7724, n7723, n7722, n7721, n7720, n7719, n7718,
         n7717, n7716, n7715, n7714, n7713, n7712, n7711, n7710, n7709, n7708,
         n7707, n7706, n7705, n7704, n7703, n7702, n7701, n7700, n7699, n7698,
         n7697, n7696, n7695, n7694, n7693, n7692, n7691, n7690, n7689, n7688,
         n7687, n7686, n7685, n7684, n7683, n7682, n7681, n7680, n7679, n7678,
         n7677, n7676, n7675, n7674, n7673, n7672, n7671, n7670, n7669, n7668,
         n7667, n7666, n7665, n7664, n7663, n7662, n7661, n7660, n7659, n7658,
         n7657, n7656, n7655, n7654, n7653, n7652, n7651, n7650, n7649, n7648,
         n7647, n7646, n7645, n7644, n7642, n7641, n7640, n7639, n7638, n7637,
         n7636, n7635, n7634, n7633, n7632, n7631, n7630, n7629, n7628, n7627,
         n7626, n7625, n7624, n7623, n7622, n7621, n7620, n7619, n7618, n7617,
         n7616, n7615, n7614, n7613, n7612, n7611, n7610, n7609, n7608, n7607,
         n7606, n7605, n7604, n7603, n7602, n7601, n7600, n7599, n7598, n7597,
         n7596, n7595, n7594, n7593, n7592, n7591, n7590, n7589, n7588, n7587,
         n7586, n7585, n7584, n7583, n7582, n7581, n7580, n7579, n7578, n7577,
         n7576, n7575, n7574, n7573, n7572, n7571, n7570, n7569, n7568, n7567,
         n7566, n7565, n7564, n7563, n7562, n7561, n7560, n7559, n7558, n7557,
         n7556, n7555, n7554, n7553, n7552, n7551, n7550, n7549, n7548, n7547,
         n7546, n7545, n7544, n7543, n7542, n7541, n7540, n7539, n7538, n7537,
         n7536, n7535, n7534, n7533, n7532, n7531, n7530, n7529, n7528, n7527,
         n7526, n7525, n7524, n7523, n7522, n7521, n7520, n7519, n7518, n7517,
         n7516, n7515, n7514, n7513, n7512, n7511, n7510, n7509, n7508, n7507,
         n7506, n7505, n7504, n7503, n7502, n7501, n7500, n7499, n7498, n7497,
         n7496, n7495, n7494, n7493, n7492, n7491, n7490, n7489, n7488, n7487,
         n7486, n7485, n7484, n7483, n7482, n7481, n7480, n7479, n7478, n7477,
         n7476, n7475, n7474, n7473, n7472, n7471, n7470, n7469, n7468, n7467,
         n7466, n7465, n7464, n7463, n7462, n7461, n7460, n7459, n7458, n7457,
         n7456, n7455, n7454, n7453, n7452, n7451, n7450, n7449, n7448, n7447,
         n7446, n7445, n7444, n7443, n7442, n7441, n7440, n7439, n7438, n7437,
         n7436, n7435, n7434, n7433, n7432, n7431, n7430, n7429, n7428, n7427,
         n7426, n7425, n7424, n7423, n7422, n7421, n7420, n7419, n7418, n7417,
         n7416, n7415, n7414, n7413, n7412, n7411, n7410, n7409, n7408, n7407,
         n7406, n7405, n7404, n7403, n7402, n7401, n7400, n7399, n7398, n7397,
         n7396, n7395, n7394, n7393, n7392, n7391, n7390, n7389, n7388, n7387,
         n7386, n7385, n7384, n7383, n7382, n7381, n7380, n7379, n7378, n7377,
         n7376, n7375, n7374, n7373, n7372, n7371, n7370, n7369, n7368, n7367,
         n7366, n7365, n7364, n7363, n7362, n7361, n7360, n7359, n7358, n7357,
         n7356, n7355, n7354, n7353, n7352, n7351, n7350, n7349, n7348, n7346,
         n7345, n7344, n7343, n7342, n7341, n7340, n7339, n7338, n7337, n7336,
         n7335, n7334, n7333, n7332, n7331, n7330, n7329, n7328, n7327, n7326,
         n7325, n7324, n7323, n7322, n7321, n7320, n7319, n7318, n7317, n7316,
         n7315, n7314, n7313, n7312, n7311, n7310, n7309, n7308, n7307, n7306,
         n7305, n7304, n7303, n7302, n7301, n7300, n7299, n7298, n7297, n7296,
         n7295, n7294, n7293, n7292, n7291, n7290, n7289, n7288, n7287, n7286,
         n7285, n7283, n7282, n7281, n7280, n7279, n7278, n7277, n7276, n7275,
         n7274, n7273, n7272, n7271, n7270, n7269, n7268, n7267, n7266, n7265,
         n7264, n7263, n7262, n7260, n7259, n7258, n7257, n7256, n7255, n7254,
         n7253, n7252, n7251, n7250, n7249, n7248, n7247, n7246, n7245, n7244,
         n7243, n7242, n7241, n7240, n7239, n7238, n7237, n7236, n7235, n7234,
         n7233, n7232, n7231, n7230, n7229, n7228, n7227, n7226, n7225, n7224,
         n7223, n7222, n7221, n7220, n7219, n7218, n7217, n7215, n7214, n7213,
         n7212, n7211, n7210, n7209, n7208, n7207, n7206, n7205, n7204, n7203,
         n7202, n7201, n7200, n7199, n7198, n7197, n7196, n7195, n7194, n7193,
         n7192, n7191, n7190, n7189, n7188, n7187, n7186, n7185, n7184, n7183,
         n7182, n7181, n7180, n7179, n7178, n7177, n7176, n7175, n7174, n7173,
         n7172, n7171, n7170, n7169, n7168, n7167, n7166, n7165, n7164, n7163,
         n7162, n7161, n7160, n7159, n7158, n7157, n7156, n7155, n7154, n7153,
         n7152, n7151, n7150, n7149, n7148, n7147, n7146, n7145, n7144, n7143,
         n7142, n7141, n7140, n7139, n7138, n7137, n7136, n7135, n7134, n7133,
         n7132, n7131, n7130, n7129, n7128, n7127, n7126, n7125, n7124, n7123,
         n7122, n7121, n7120, n7119, n7118, n7117, n7116, n7115, n7114, n7113,
         n7112, n7111, n7110, n7109, n7108, n7107, n7106, n7105, n7104, n7103,
         n7102, n7101, n7100, n7099, n7098, n7097, n7096, n7095, n7094, n7093,
         n7092, n7091, n7090, n7089, n7088, n7087, n7086, n7085, n7084, n7082,
         n7081, n7080, n7079, n7078, n7077, n7076, n7075, n7074, n7073, n7072,
         n7071, n7070, n7069, n7068, n7067, n7066, n7065, n7064, n7063, n7062,
         n7061, n7060, n7059, n7058, n7057, n7056, n7055, n7054, n7053, n7052,
         n7051, n7050, n7049, n7048, n7047, n7046, n7045, n7044, n7043, n7042,
         n7041, n7040, n7039, n7038, n7037, n7035, n7034, n7033, n7032, n7031,
         n7030, n7029, n7028, n7027, n7026, n7025, n7024, n7023, n7022, n7021,
         n7020, n7019, n7018, n7017, n7016, n7015, n7014, n7013, n7012, n7011,
         n7010, n7009, n7008, n7007, n7006, n7005, n7004, n7003, n7002, n7001,
         n7000, n6999, n6997, n6996, n6995, n6994, n6993, n6992, n6991, n6990,
         n6989, n6988, n6987, n6986, n6985, n6984, n6983, n6982, n6981, n6980,
         n6979, n6978, n6977, n6976, n6975, n6974, n6973, n6972, n6971, n6970,
         n6969, n6968, n6967, n6966, n6965, n6964, n6963, n6962, n6961, n6960,
         n6959, n6958, n6957, n6956, n6955, n6954, n6953, n6952, n6951, n6950,
         n6949, n6948, n6947, n6945, n6944, n6943, n6942, n6941, n6940, n6939,
         n6938, n6937, n6936, n6935, n6934, n6933, n6932, n6931, n6930, n6929,
         n6928, n6927, n6926, n6925, n6924, n6923, n6922, n6921, n6920, n6919,
         n6918, n6917, n6916, n6915, n6914, n6913, n6912, n6911, n6910, n6909,
         n6908, n6907, n6906, n6905, n6904, n6903, n6902, n6901, n6900, n6899,
         n6898, n6897, n6896, n6895, n6894, n6893, n6892, n6891, n6890, n6889,
         n6888, n6887, n6886, n6885, n6884, n6883, n6882, n6881, n6880, n6879,
         n6878, n6877, n6876, n6875, n6874, n6873, n6872, n6871, n6870, n6869,
         n6868, n6867, n6866, n6865, n6864, n6863, n6862, n6861, n6860, n6859,
         n6858, n6857, n6856, n6855, n6854, n6853, n6852, n6851, n6850, n6849,
         n6848, n6847, n6846, n6845, n6844, n6843, n6842, n6841, n6840, n6839,
         n6838, n6837, n6836, n6835, n6834, n6833, n6832, n6831, n6830, n6829,
         n6828, n6827, n6826, n6825, n6824, n6823, n6822, n6821, n6820, n6819,
         n6818, n6817, n6816, n6815, n6814, n6813, n6812, n6811, n6810, n6809,
         n6808, n6807, n6806, n6805, n6804, n6803, n6802, n6801, n6800, n6799,
         n6798, n6797, n6796, n6795, n6794, n6793, n6792, n6791, n6790, n6789,
         n6788, n6787, n6786, n6785, n6784, n6783, n6782, n6781, n6780, n6779,
         n6778, n6777, n6776, n6775, n6774, n6773, n6772, n6771, n6770, n6769,
         n6768, n6767, n6766, n6765, n6764, n6763, n6762, n6761, n6760, n6759,
         n6758, n6757, n6756, n6755, n6754, n6753, n6752, n6751, n6750, n6749,
         n6748, n6747, n6746, n6745, n6744, n6743, n6742, n6741, n6740, n6739,
         n6738, n6737, n6736, n6735, n6734, n6733, n6732, n6731, n6730, n6729,
         n6728, n6727, n6726, n6725, n6724, n6723, n6722, n6721, n6720, n6719,
         n6718, n6717, n6716, n6715, n6714, n6713, n6712, n6711, n6710, n6709,
         n6708, n6707, n6706, n6705, n6704, n6703, n6702, n6701, n6700, n6699,
         n6698, n6697, n6696, n6695, n6694, n6693, n6692, n6691, n6690, n6689,
         n6687, n6686, n6685, n6684, n6683, n6680, n6679, n6678, n6677, n6676,
         n6675, n6674, n6673, n6672, n6671, n6670, n6669, n6668, n6667, n6666,
         n6665, n6664, n6663, n6662, n6661, n6660, n6659, n6658, n6657, n6655,
         n6654, n6653, n6652, n6651, n6650, n6649, n6648, n6647, n6646, n6645,
         n6644, n6643, n6642, n6641, n6639, n6638, n6637, n6636, n6635, n6633,
         n6632, n6631, n6630, n6629, n6628, n6627, n6626, n6625, n6624, n6623,
         n6622, n6621, n6620, n6619, n6617, n6616, n6615, n6614, n6613, n6612,
         n6611, n6609, n6608, n6607, n6606, n6605, n6604, n6603, n6602, n6601,
         n6600, n6599, n6598, n6597, n6596, n6594, n6593, n6592, n6591, n6590,
         n6588, n6587, n6586, n6585, n6584, n6583, n6582, n6581, n6580, n6579,
         n6578, n6577, n6576, n6575, n6573, n6572, n6571, n6570, n6569, n6568,
         n6567, n6565, n6564, n6563, n6562, n6561, n6560, n6559, n6558, n6557,
         n6556, n6555, n6554, n6553, n6552, n6550, n6549, n6548, n6547, n6546,
         n6544, n6543, n6542, n6541, n6540, n6539, n6538, n6537, n6536, n6535,
         n6534, n6533, n6532, n6531, n6530, n6528, n6527, n6526, n6525, n6524,
         n6523, n6522, n6520, n6519, n6518, n6517, n6516, n6515, n6514, n6513,
         n6512, n6511, n6510, n6509, n6508, n6507, n6505, n6504, n6503, n6502,
         n6501, n6499, n6498, n6497, n6496, n6495, n6494, n6493, n6492, n6491,
         n6490, n6489, n6488, n6487, n6486, n6484, n6483, n6482, n6481, n6480,
         n6479, n6478, n6476, n6475, n6474, n6473, n6472, n6471, n6470, n6469,
         n6468, n6467, n6466, n6465, n6464, n6463, n6461, n6460, n6459, n6458,
         n6457, n6455, n6454, n6453, n6452, n6451, n6450, n6449, n6448, n6447,
         n6446, n6445, n6444, n6443, n6442, n6441, n6439, n6438, n6437, n6436,
         n6435, n6434, n6433, n6431, n6430, n6429, n6428, n6427, n6426, n6425,
         n6424, n6423, n6422, n6421, n6420, n6419, n6418, n6416, n6415, n6414,
         n6413, n6412, n6410, n6409, n6408, n6407, n6406, n6405, n6404, n6403,
         n6402, n6401, n6400, n6399, n6398, n6397, n6395, n6394, n6393, n6392,
         n6391, n6390, n6389, n6387, n6386, n6385, n6384, n6383, n6382, n6381,
         n6380, n6379, n6378, n6377, n6376, n6375, n6374, n6372, n6371, n6370,
         n6369, n6368, n6366, n6365, n6364, n6363, n6362, n6361, n6360, n6359,
         n6358, n6357, n6356, n6355, n6354, n6353, n6352, n6350, n6349, n6348,
         n6347, n6346, n6345, n6344, n6342, n6341, n6340, n6339, n6338, n6337,
         n6336, n6335, n6334, n6333, n6332, n6331, n6330, n6329, n6327, n6326,
         n6325, n6324, n6323, n6321, n6320, n6319, n6318, n6317, n6316, n6315,
         n6314, n6313, n6312, n6311, n6310, n6309, n6308, n6306, n6305, n6304,
         n6303, n6302, n6301, n6300, n6298, n6297, n6296, n6295, n6294, n6293,
         n6292, n6291, n6290, n6289, n6288, n6287, n6286, n6285, n6283, n6282,
         n6281, n6280, n6279, n6277, n6276, n6275, n6274, n6273, n6272, n6271,
         n6270, n6269, n6268, n6267, n6266, n6265, n6264, n6263, n6261, n6260,
         n6259, n6258, n6257, n6256, n6255, n6253, n6252, n6251, n6250, n6249,
         n6248, n6247, n6246, n6245, n6244, n6243, n6242, n6241, n6240, n6238,
         n6237, n6236, n6235, n6234, n6232, n6231, n6230, n6229, n6228, n6227,
         n6226, n6225, n6224, n6223, n6222, n6221, n6220, n6219, n6218, n6217,
         n6216, n6215, n6214, n6213, n6212, n6211, n6210, n6209, n6208, n6207,
         n6206, n6205, n6204, n6203, n6202, n6201, n6200, n6199, n6198, n6197,
         n6196, n6195, n6194, n6193, n6192, n6191, n6190, n6189, n6188, n6186,
         n6185, n6184, n6183, n6182, n6181, n6180, n6178, n6177, n6176, n6175,
         n6174, n6173, n6172, n6171, n6170, n6169, n6168, n6167, n6166, n6165,
         n6164, n6163, n6162, n6161, n6160, n6159, n6158, n6157, n6156, n6155,
         n6154, n6153, n6152, n6151, n6150, n6149, n6148, n6147, n6146, n6145,
         n6144, n6143, n6142, n6140, n6139, n6138, n6137, n6136, n6135, n6134,
         n6133, n6132, n6131, n6130, n6129, n6128, n6127, n6126, n6125, n6124,
         n6123, n6122, n6121, n6120, n6119, n6118, n6117, n6116, n6115, n6114,
         n6113, n6112, n6111, n6110, n6109, n6108, n6107, n6106, n6105, n6104,
         n6103, n6102, n6101, n6100, n6099, n6098, n6097, n6096, n6095, n6094,
         n6093, n6092, n6091, n6090, n6089, n6087, n6086, n6085, n6084, n6083,
         n6082, n6081, n6080, n6079, n6078, n6077, n6076, n6075, n6074, n6073,
         n6071, n6070, n6069, n6068, n6067, n6066, n6065, n6064, n6063, n6062,
         n6061, n6060, n6059, n6058, n6057, n6055, n6054, n6053, n6051, n6050,
         n6049, n6048, n6047, n6045, n6044, n6043, n6042, n6041, n6040, n6039,
         n6038, n6037, n6036, n6035, n6034, n6033, n6032, n6031, n6030, n6029,
         n6028, n6027, n6026, n6025, n6024, n6023, n6022, n6021, n6020, n6018,
         n6017, n6016, n6015, n6014, n6013, n6012, n6011, n6010, n6009, n6008,
         n6006, n6005, n6003, n6002, n6001, n6000, n5999, n5998, n5997, n5996,
         n5995, n5994, n5993, n5992, n5991, n5990, n5987, n5985, n5984, n5983,
         n5982, n5981, n5980, n5979, n5978, n5977, n5976, n5974, n5973, n5972,
         n5971, n5970, n5969, n5968, n5967, n5966, n5965, n5964, n5963, n5962,
         n5961, n5960, n5959, n5958, n5957, n5956, n5955, n5954, n5953, n5952,
         n5951, n5950, n5949, n5948, n5947, n5946, n5945, n5944, n5943, n5942,
         n5941, n5940, n5939, n5938, n5937, n5936, n5935, n5934, n5933, n5932,
         n5931, n5930, n5929, n5928, n5927, n5926, n5925, n5924, n5923, n5922,
         n5921, n5920, n5919, n5918, n5917, n5916, n5915, n5914, n5913, n5912,
         n5911, n5910, n5909, n5908, n5907, n5906, n5905, n5904, n5903, n5902,
         n5901, n5900, n5899, n5898, n5897, n5896, n5895, n5894, n5893, n5892,
         n5891, n5890, n5889, n5888, n5887, n5886, n5885, n5884, n5883, n5882,
         n5881, n5880, n5879, n5878, n5877, n5876, n5875, n5874, n5873, n5872,
         n5871, n5870, n5869, n5868, n5867, n5866, n5865, n5864, n5863, n5862,
         n5861, n5860, n5859, n5858, n5856, n5855, n5854, n5853, n5852, n5851,
         n5850, n5849, n5848, n5847, n5846, n5845, n5844, n5843, n5842, n5841,
         n5840, n5839, n5838, n5837, n5836, n5835, n5834, n5833, n5832, n5831,
         n5830, n5829, n5828, n5827, n5826, n5825, n5824, n5823, n5822, n5821,
         n5820, n5819, n5818, n5817, n5816, n5815, n5814, n5813, n5812, n5811,
         n5810, n5809, n5808, n5807, n5806, n5805, n5804, n5803, n5802, n5801,
         n5800, n5799, n5798, n5797, n5796, n5795, n5794, n5793, n5792, n5791,
         n5790, n5789, n5788, n5787, n5786, n5785, n5784, n5783, n5782, n5781,
         n5780, n5779, n5778, n5777, n5776, n5775, n5774, n5773, n5772, n5771,
         n5769, n5768, n5767, n5766, n5765, n5764, n5763, n5762, n5761, n5760,
         n5759, n5758, n5757, n5756, n5755, n5754, n5753, n5752, n5751, n5750,
         n5749, n5748, n5747, n5745, n5744, n5743, n5742, n5741, n5740, n5739,
         n5738, n5737, n5736, n5735, n5734, n5732, n5731, n5730, n5729, n5728,
         n5727, n5726, n5725, n5724, n5723, n5722, n5721, n5720, n5719, n5718,
         n5717, n5716, n5715, n5714, n5713, n5712, n5711, n5710, n5709, n5708,
         n5707, n5706, n5705, n5704, n5703, n5702, n5700, n5699, n5698, n5697,
         n5696, n5695, n5694, n5693, n5692, n5691, n5690, n5689, n5687, n5685,
         n5684, n5683, n5682, n5681, n5680, n5679, n5678, n5677, n5676, n5675,
         n5674, n5673, n5672, n5671, n5670, n5669, n5668, n5667, n5666, n5665,
         n5664, n5663, n5662, n5661, n5660, n5659, n5658, n5657, n5656, n5655,
         n5654, n5653, n5652, n5651, n5650, n5649, n5648, n5647, n5646, n5645,
         n5644, n5643, n5642, n5628, n5627, n5626, n5625, n5624, n5623, n5622,
         n5621, n5620, n5619, n5618, n5617, n5616, n5615, n5614, n5613, n5612,
         n5611, n5610, n5609, n5608, n5607, n5606, n5605, n5604, n5603, n5602,
         n5601, n5600, n5599, n5598, n5597, n5596, n5595, n5594, n5593, n5592,
         n5591, n5590, n5589, n5588, n5587, n5586, n5585, n5584, n5583, n5582,
         n5581, n5580, n5579, n5578, n5577, n5576, n5575, n5574, n5573, n5572,
         n5571, n5570, n5569, n5568, n5567, n5566, n5556, n5555, n5554, n5553,
         n5552, n5551, n5550, n5549, n5548, n5547, n5546, n5545, n5544, n5543,
         n5542, n5541, n5540, n5539, n5538, n5537, n5536, n5534, n5533, n5532,
         n5531, n5530, n5529, n5528, n5527, n5526, n5525, n5524, n5523, n5522,
         n5521, n5520, n5519, n5518, n5517, n5516, n5514, n5513, n5512, n5511,
         n5510, n5509, n5508, n5507, n5506, n5505, n5504, n5503, n5502, n5501,
         n5500, n5499, n5498, n5497, n5496, n5494, n5493, n5492, n5491, n5490,
         n5480, n5479, n5478, n5477, n5476, n5475, n5474, n5473, n5472, n5471,
         n5470, n5469, n5468, n5467, n5466, n5465, n5464, n5463, n5462, n5461,
         n5460, n5459, n5458, n5457, n5456, n5455, n5454, n5453, n5452, n5451,
         n5450, n5449, n5448, n5447, n5446, n5445, n5444, n5443, n5442, n5441,
         n5440, n5439, n5438, n5437, n5436, n5435, n5434, n5433, n5432, n5431,
         n5430, n5429, n5428, n5427, n5426, n5425, n5424, n5423, n5422, n5421,
         n5420, n5419, n5418, n5417, n5415, n5414, n5413, n5412, n5411, n5410,
         n5409, n5408, n5406, n5404, n5402, n5400, n5399, n5398, n5397, n5396,
         n5395, n5394, n5393, n5392, n5391, n5390, n5389, n5388, n5387, n5386,
         n5385, n5384, n5383, n5382, n5381, n5380, n5379, n5378, n5377, n5376,
         n5375, n5374, n5373, n5372, n5371, n5370, n5369, n5368, n5367, n5366,
         n5365, n5364, n5363, n5362, n5361, n5360, n5359, n5358, n5357, n5356,
         n5355, n5354, n5353, n5352, n5351, n5350, n5349, n5348, n5347, n5346,
         n5345, n5344, n5343, n5342, n5341, n5340, n5339, n5338, n5337, n5336,
         n5335, n5334, n5333, n5332, n5331, n5330, n5329, n5328, n5327, n5326,
         n5325, n5324, n5323, n5322, n5321, n5320, n5319, n5318, n5317, n5316,
         n5315, n5314, n5313, n5312, n5311, n5310, n5309, n5308, n5307, n5306,
         n5305, n5304, n5303, n5302, n5301, n5300, n5299, n5298, n5297, n5296,
         n5295, n5294, n5293, n5292, n5291, n5290, n5289, n5288, n5287, n5286,
         n5285, n5284, n5283, n5282, n5281, n5280, n5279, n5278, n5277, n5276,
         n5275, n5274, n5273, n5272, n5271, n5270, n5269, n5268, n5267, n5266,
         n5265, n5264, n5263, n5262, n5261, n5260, n5259, n5258, n5257, n5256,
         n5255, n5254, n5253, n5252, n5251, n5250, n5249, n5248, n5247, n5246,
         n5245, n5244, n5243, n5242, n5241, n5240, n5239, n5238, n5237, n5236,
         n5235, n5234, n5233, n5232, n5231, n5230, n5229, n5228, n5227, n5226,
         n5225, n5224, n5223, n5222, n5221, n5220, n5219, n5218, n5217, n5216,
         n5215, n5214, n5213, n5212, n5211, n5210, n5209, n5208, n5207, n5206,
         n5205, n5204, n5203, n5202, n5201, n5200, n5199, n5198, n5197, n5196,
         n5195, n5194, n5193, n5192, n5191, n5190, n5189, n5188, n5187, n5186,
         n5185, n5184, n5183, n5182, n5181, n5180, n5179, n5178, n5177, n5176,
         n5175, n5174, n5173, n5172, n5171, n5170, n5169, n5168, n5167, n5166,
         n5165, n5164, n5163, n5162, n5161, n5160, n5159, n5158, n5157, n5156,
         n5155, n5154, n5153, n5152, n5151, n5149, n5148, n5147, n5146, n5145,
         n5144, n5143, n5142, n5141, n5140, n5139, n5138, n5137, n5136, n5135,
         n5134, n5133, n5132, n5131, n5130, n5129, n5128, n5127, n5126, n5125,
         n5124, n5123, n5122, n5121, n5120, n5119, n5118, n5117, n5116, n5115,
         n5114, n5113, n5112, n5111, n5110, n5109, n5108, n5107, n5106, n5105,
         n5104, n5103, n5102, n29275, n29274, n29273, n29272, n29271, n29270,
         n29269, n29268, n29267, n29266, n29265, n29264, n29263, n29262,
         n29261, n29260, n29259, n29258, n29257, n29256, n29255, n29254,
         n29253, n29252, n29251, n29250, n29249, n29248, n29247, n29246,
         n29245, n29244, n29243, n29242, n29241, n29240, n29239, n29238,
         n29237, n29236, n29235, n29234, n29233, n29232, n29231, n29230,
         n29229, n29228, n29227, n29226, n29225, n29224, n29223, n29222,
         n29221, n29220, n29219, n29218, n29217, n29216, n29215, n29214,
         n29213, n29212, n29211, n29210, n29209, n29208, n29207, n29206,
         n29205, n29204, n29203, n29202, n29201, n29200, n29199, n29198,
         n29197, n29196, n29195, n29194, n29193, n29192, n29191, n29190,
         n29189, n29188, n29187, n29186, n29185, n29184, n29183, n29182,
         n29181, n29180, n29179, n29178, n29177, n29176, n29175, n29174,
         n29173, n29172, n29171, n29170, n29169, n29168, n29167, n29166,
         n29165, n29164, n29163, n29162, n29161, n29160, n29159, n29158,
         n29157, n29156, n29155, n29154, n29153, n29152, n29151, n29150,
         n29149, n29148, n29147, n29146, n29145, n29144, n29143, n29142,
         n29141, n29140, n29139, n29138, n29137, n29136, n29135, n29134,
         n29133, n29132, n29131, n29130, n29129, n29128, n29127, n29126,
         n29125, n29124, n29123, n29122, n29121, n29120, n29119, n29118,
         n29117, n29116, n29115, n29114, n29113, n29112, n29111, n29110,
         n29109, n29108, n29107, n29106, n29105, n29104, n29103, n29102,
         n29101, n29100, n29099, n29098, n29097, n29096, n29095, n29094,
         n29093, n29092, n29091, n29090, n29089, n29088, n29087, n29086,
         n29085, n29084, n29083, n29082, n29081, n29080, n29079, n29078,
         n29077, n29076, n29075, n29074, n29073, n29072, n29071, n29070,
         n29069, n29068, n29067, n29066, n29065, n29064, n29063, n29062,
         n29061, n29060, n29059, n29058, n29057, n29056, n29055, n29054,
         n29053, n29052, n29051, n29050, n29049, n29048, n29047, n29046,
         n29045, n29044, n29043, n29042, n29041, n29040, n29039, n29038,
         n29037, n29036, n29035, n29034, n29033, n29032, n29031, n29030,
         n29029, n29028, n29027, n29026, n29025, n29024, n29023, n29022,
         n29021, n29020, n29019, n29018, n29017, n29016, n29015, n29014,
         n29013, n29012, n29011, n29010, n29009, n29008, n29007, n29006,
         n29005, n29004, n29003, n29002, n29001, n29000, n28999, n28998,
         n28997, n28996, n28995, n28994, n28993, n28992, n28991, n28990,
         n28989, n28988, n28987, n28986, n28985, n28984, n28983, n28982,
         n28981, n28980, n28979, n28978, n28977, n28976, n28975, n28974,
         n28973, n28972, n28971, n28970, n28969, n28968, n28967, n28966,
         n28965, n28964, n28963, n28962, n28961, n28960, n28959, n28958,
         n28957, n28956, n28955, n28954, n28953, n28952, n28951, n28950,
         n28949, n28948, n28947, n28946, n28945, n28944, n28943, n28942,
         n28941, n28940, n28939, n28938, n28937, n28936, n28935, n28934,
         n28933, n28932, n28931, n28930, n28929, n28928, n28927, n28926,
         n28925, n28924, n28923, n28922, n28921, n28920, n28919, n28918,
         n28917, n28916, n28915, n28914, n28913, n28912, n28911, n28910,
         n28909, n28908, n28907, n28906, n28905, n28904, n28903, n28902,
         n28901, n28900, n28899, n28898, n28897, n28896, n28895, n28894,
         n28893, n28892, n28891, n28890, n28889, n28888, n28887, n28886,
         n28885, n28884, n28883, n28882, n28881, n28880, n28879, n28878,
         n28877, n28876, n28875, n28874, n28873, n28872, n28871, n28870,
         n28869, n28868, n28867, n28866, n28865, n28864, n28863, n28862,
         n28861, n28860, n28859, n28858, n28857, n28856, n28855, n28854,
         n28853, n28852, n28851, n28850, n28849, n28848, n28847, n28846,
         n28845, n28844, n28843, n28842, n28841, n28840, n28839, n28838,
         n28837, n28836, n28835, n28834, n28833, n28832, n28831, n28830,
         n28829, n28828, n28827, n28826, n28825, n28824, n28823, n28822,
         n28821, n28820, n28819, n28818, n28817, n28816, n28815, n28814,
         n28813, n28812, n28811, n28810, n28809, n28808, n28807, n28806,
         n28805, n28804, n28803, n28802, n28801, n28800, n28799, n28798,
         n28797, n28796, n28795, n28794, n28793, n28792, n28791, n28790,
         n28789, n28788, n28787, n28786, n28785, n28784, n28783, n28782,
         n28781, n28780, n28779, n28778, n28777, n28776, n28775, n28774,
         n28773, n28772, n28771, n28770, n28769, n28768, n28767, n28766,
         n28765, n28764, n28763, n28762, n28761, n28760, n28759, n28758,
         n28757, n28756, n28755, n28754, n28753, n28752, n28751, n28750,
         n28749, n28748, n28747, n28746, n28745, n28744, n28743, n28742,
         n28741, n28740, n28739, n28738, n28737, n28736, n28735, n28734,
         n28733, n28732, n28731, n28730, n28729, n28728, n28727, n28726,
         n28725, n28724, n28723, n28722, n28721, n28720, n28719, n28718,
         n28717, n28716, n28715, n28714, n28713, n28712, n28711, n28710,
         n28709, n28708, n28707, n28706, n28705, n28704, n28703, n28702,
         n28701, n28700, n28699, n28698, n28697, n28696, n28695, n28694,
         n28693, n28692, n28691, n28690, n28689, n28688, n28687, n28686,
         n28685, n28684, n28683, n28682, n28681, n28680, n28679, n28678,
         n28677, n28676, n28675, n28674, n28673, n28672, n28671, n28670,
         n28669, n28668, n28667, n28666, n28665, n28664, n28663, n28662,
         n28661, n28660, n28659, n28658, n28657, n28656, n28655, n28654,
         n28653, n28652, n28651, n28650, n28649, n28648, n28647, n28646,
         n28645, n28644, n28643, n28642, n28641, n28640, n28639, n28638,
         n28637, n28636, n28635, n28634, n28633, n28632, n28631, n28630,
         n28629, n28628, n28627, n28626, n28625, n28624, n28623, n28622,
         n28621, n28620, n28619, n28618, n28617, n28616, n28615, n28614,
         n28613, n28612, n28611, n28610, n28609, n28608, n28607, n28606,
         n28605, n28604, n28603, n28602, n28601, n28600, n28599, n28598,
         n28597, n28596, n28595, n28594, n28593, n28592, n28591, n28590,
         n28589, n28588, n28587, n28586, n28585, n28584, n28583, n28582,
         n28581, n28580, n28579, n28578, n28577, n28576, n28575, n28574,
         n28573, n28572, n28571, n28570, n28569, n28568, n28567, n28566,
         n28565, n28564, n28563, n28562, n28561, n28560, n28559, n28558,
         n28557, n28556, n28555, n28554, n28553, n28552, n28551, n28550,
         n28549, n28548, n28547, n28546, n28545, n28544, n28543, n28542,
         n28541, n28540, n28539, n28538, n28537, n28536, n28535, n28534,
         n28533, n28532, n28531, n28530, n28529, n28528, n28527, n28526,
         n28525, n28524, n28523, n28522, n28521, n28520, n28519, n28518,
         n28517, n28516, n28515, n28514, n28513, n28512, n28511, n28510,
         n28509, n28508, n28507, n28506, n28505, n28504, n28503, n28502,
         n28501, n28500, n28499, n28498, n28497, n28496, n28495, n28494,
         n28493, n28492, n28491, n28490, n28489, n28488, n28487, n28486,
         n28485, n28484, n28483, n28482, n28481, n28480, n28479, n28478,
         n28477, n28476, n28475, n28474, n28473, n28472, n28471, n28470,
         n28469, n28468, n28467, n28466, n28465, n28464, n28463, n28462,
         n28461, n28460, n28459, n28458, n28457, n28456, n28455, n28454,
         n28453, n28452, n28451, n28450, n28449, n28448, n28447, n28446,
         n28445, n28444, n28443, n28442, n28441, n28440, n28439, n28438,
         n28437, n28436, n28435, n28434, n28433, n28432, n28431, n28430,
         n28429, n28428, n28427, n28426, n28425, n28424, n28423, n28422,
         n28421, n28420, n28419, n28418, n28417, n28416, n28415, n28414,
         n28413, n28412, n28411, n28410, n28409, n28408, n28407, n28406,
         n28405, n28404, n28403, n28402, n28401, n28400, n28399, n28398,
         n28397, n28396, n28395, n28394, n28393, n28392, n28391, n28390,
         n28389, n28388, n28387, n28386, n28385, n28384, n28383, n28382,
         n28381, n28380, n28379, n28378, n28377, n28376, n28375, n28374,
         n28373, n28372, n28371, n28370, n28369, n28368, n28367, n28366,
         n28365, n28364, n28363, n28362, n28361, n28360, n28359, n28358,
         n28357, n28356, n28355, n28354, n28353, n28352, n28351, n28350,
         n28349, n28348, n28347, n28346, n28345, n28344, n28343, n28342,
         n28341, n28340, n28339, n28338, n28337, n28336, n28335, n28334,
         n28333, n28332, n28331, n28330, n28329, n28328, n28327, n28326,
         n28325, n28324, n28323, n28322, n28321, n28320, n28319, n28318,
         n28317, n28316, n28315, n28314, n28313, n28312, n28311, n28310,
         n28309, n28308, n28307, n28306, n28305, n28304, n28303, n28302,
         n28301, n28300, n28299, n28298, n28297, n28296, n28295, n28294,
         n28293, n28292, n28291, n28290, n28289, n28288, n28287, n28286,
         n28285, n28284, n28283, n28282, n28281, n28280, n28279, n28278,
         n28277, n28276, n28275, n28274, n28273, n28272, n28271, n28270,
         n28269, n28268, n28267, n28266, n28265, n28264, n28263, n28262,
         n28261, n28260, n28259, n28258, n28257, n28256, n28255, n28254,
         n28253, n28252, n28251, n28250, n28249, n28248, n28247, n28246,
         n28245, n28244, n28243, n28242, n28241, n28240, n28239, n28238,
         n28237, n28236, n28235, n28234, n28233, n28232, n28231, n28230,
         n28229, n28228, n28227, n28226, n28225, n28224, n28223, n28222,
         n28221, n28220, n28219, n28218, n28217, n28216, n28215, n28214,
         n28213, n28212, n28211, n28210, n28209, n28208, n28207, n28206,
         n28205, n28204, n28203, n28202, n28201, n28200, n28199, n28198,
         n28197, n28196, n28195, n28194, n28193, n28192, n28191, n28190,
         n28189, n28188, n28187, n28186, n28185, n28184, n28183, n28182,
         n28181, n28180, n28179, n28178, n28177, n28176, n28175, n28174,
         n28173, n28172, n28171, n28170, n28169, n28168, n28167, n28166,
         n28165, n28164, n28163, n28162, n28161, n28160, n28159, n28158,
         n28157, n28156, n28155, n28154, n28153, n28152, n28151, n28150,
         n28149, n28148, n28147, n28146, n28145, n28144, n28143, n28142,
         n28141, n28140, n28139, n28138, n28137, n28136, n28135, n28134,
         n28133, n28132, n28131, n28130, n28129, n28128, n28127, n28126,
         n28125, n28124, n28123, n28122, n28121, n28120, n28119, n28118,
         n28117, n28116, n28115, n28114, n28113, n28112, n28111, n28110,
         n28109, n28108, n28107, n28106, n28105, n28104, n28103, n28102,
         n28101, n28100, n28099, n28098, n28097, n28096, n28095, n28094,
         n28093, n28092, n28091, n28090, n28089, n28088, n28087, n28086,
         n28085, n28084, n28083, n28082, n28081, n28080, n28079, n28078,
         n28077, n28076, n28075, n28074, n28073, n28072, n28071, n28070,
         n28069, n28068, n28067, n28066, n28065, n28064, n28063, n28062,
         n28061, n28060, n28059, n28058, n28057, n28056, n28055, n28054,
         n28053, n28052, n28051, n28050, n28049, n28048, n28047, n28046,
         n28045, n28044, n28043, n28042, n28041, n28040, n28039, n28038,
         n28037, n28036, n28035, n28034, n28033, n28032, n28031, n28030,
         n28029, n28028, n28027, n28026, n28025, n28024, n28023, n28022,
         n28021, n28020, n28019, n28018, n28017, n28016, n28015, n28014,
         n28013, n28012, n28011, n28010, n28009, n28008, n28007, n28006,
         n28005, n28004, n28003, n28002, n28001, n28000, n27999, n27998,
         n27997, n27996, n27995, n27994, n27993, n27992, n27991, n27990,
         n27989, n27988, n27987, n27986, n27985, n27984, n27983, n27982,
         n27981, n27980, n27979, n27978, n27977, n27976, n27975, n27974,
         n27973, n27972, n27971, n27970, n27969, n27968, n27967, n27966,
         n27965, n27964, n27963, n27962, n27961, n27960, n27959, n27958,
         n27957, n27956, n27955, n27954, n27953, n27952, n27951, n27950,
         n27949, n27948, n27947, n27946, n27945, n27944, n27943, n27942,
         n27941, n27940, n27939, n27938, n27937, n27936, n27935, n27934,
         n27933, n27932, n27931, n27930, n27929, n27928, n27927, n27926,
         n27925, n27924, n27923, n27922, n27921, n27920, n27919, n27918,
         n27917, n27916, n27915, n27914, n27913, n27912, n27911, n27910,
         n27909, n27908, n27907, n27906, n27905, n27904, n27903, n27902,
         n27901, n27900, n27899, n27898, n27897, n27896, n27895, n27894,
         n27893, n27892, n27891, n27890, n27889, n27888, n27887, n27886,
         n27885, n27884, n27883, n27882, n27881, n27880, n27879, n27878,
         n27877, n27876, n27875, n27874, n27873, n27872, n27871, n27870,
         n27869, n27868, n27867, n27866, n27865, n27864, n27863, n27862,
         n27861, n27860, n27859, n27858, n27857, n27856, n27855, n27854,
         n27853, n27852, n27851, n27850, n27849, n27848, n27847, n27846,
         n27845, n27844, n27843, n27842, n27841, n27840, n27839, n27838,
         n27837, n27836, n27835, n27834, n27833, n27832, n27831, n27830,
         n27829, n27828, n27827, n27826, n27825, n27824, n27823, n27822,
         n27821, n27820, n27819, n27818, n27817, n27816, n27815, n27814,
         n27813, n27812, n27811, n27810, n27809, n27808, n27807, n27806,
         n27805, n27804, n27803, n27802, n27801, n27800, n27799, n27798,
         n27797, n27796, n27795, n27794, n27793, n27792, n27791, n27790,
         n27789, n27788, n27787, n27786, n27785, n27784, n27783, n27782,
         n27781, n27780, n27779, n27778, n27777, n27776, n27775, n27774,
         n27773, n27772, n27771, n27770, n27769, n27768, n27767, n27766,
         n27765, n27764, n27763, n27762, n27761, n27760, n27759, n27758,
         n27757, n27756, n27755, n27754, n27753, n27752, n27751, n27750,
         n27749, n27748, n27747, n27746, n27745, n27744, n27743, n27742,
         n27741, n27740, n27739, n27738, n27737, n27736, n27735, n27734,
         n27733, n27732, n27731, n27730, n27729, n27728, n27727, n27726,
         n27725, n27724, n27723, n27722, n27721, n27720, n27719, n27718,
         n27717, n27716, n27715, n27714, n27713, n27712, n27711, n27710,
         n27709, n27708, n27707, n27706, n27705, n27704, n27703, n27702,
         n27701, n27700, n27699, n27698, n27697, n27696, n27695, n27694,
         n27693, n27692, n27691, n27690, n27689, n27688, n27687, n27686,
         n27685, n27684, n27683, n27682, n27681, n27680, n27679, n27678,
         n27677, n27676, n27675, n27674, n27673, n27672, n27671, n27670,
         n27669, n27668, n27667, n27666, n27665, n27664, n27663, n27662,
         n27661, n27660, n27659, n27658, n27657, n27656, n27655, n27654,
         n27653, n27652, n27651, n27650, n27649, n27648, n27647, n27646,
         n27645, n27644, n27643, n27642, n27641, n27640, n27639, n27638,
         n27637, n27636, n27635, n27634, n27633, n27632, n27631, n27630,
         n27629, n27628, n27627, n27626, n27625, n27624, n27623, n27622,
         n27621, n27620, n27619, n27618, n27617, n27616, n27615, n27614,
         n27613, n27612, n27611, n27610, n27609, n27608, n27607, n27606,
         n27605, n27604, n27603, n27602, n27601, n27600, n27599, n27598,
         n27597, n27596, n27595, n27594, n27593, n27592, n27591, n27590,
         n27589, n27588, n27587, n27586, n27585, n27584, n27583, n27582,
         n27581, n27580, n27579, n27578, n27577, n27576, n27575, n27574,
         n27573, n27572, n27571, n27570, n27569, n27568, n27567, n27566,
         n27565, n27564, n27563, n27562, n27561, n27560, n27559, n27558,
         n27557, n27556, n27555, n27554, n27553, n27552, n27551, n27550,
         n27549, n27548, n27547, n27546, n27545, n27544, n27543, n27542,
         n27541, n27540, n27539, n27538, n27537, n27536, n27535, n27534,
         n27533, n27532, n27531, n27530, n27529, n27528, n27527, n27526,
         n27525, n27524, n27523, n27522, n27521, n27520, n27519, n27518,
         n27517, n27516, n27515, n27514, n27513, n27512, n27511, n27510,
         n27509, n27508, n27507, n27506, n27505, n27504, n27503, n27502,
         n27501, n27500, n27499, n27498, n27497, n27496, n27495, n27494,
         n27493, n27492, n27491, n27490, n27489, n27488, n27487, n27486,
         n27485, n27484, n27483, n27482, n27481, n27480, n27479, n27478,
         n27477, n27476, n27475, n27474, n27473, n27472, n27471, n27470,
         n27469, n27468, n27467, n27466, n27465, n27464, n27463, n27462,
         n27461, n27460, n27459, n27458, n27457, n27456, n27455, n27454,
         n27453, n27452, n27451, n27450, n27449, n27448, n27447, n27446,
         n27445, n27444, n27443, n27442, n27441, n27440, n27439, n27438,
         n27437, n27436, n27435, n27434, n27433, n27432, n27431, n27430,
         n27429, n27428, n27427, n27426, n27425, n27424, n27423, n27422,
         n27421, n27420, n27419, n27418, n27417, n27416, n27415, n27414,
         n27413, n27412, n27411, n27410, n27409, n27408, n27407, n27406,
         n27405, n27404, n27403, n27402, n27401, n27400, n27399, n27398,
         n27397, n27396, n27395, n27394, n27393, n27392, n27391, n27390,
         n27389, n27388, n27387, n27386, n27385, n27384, n27383, n27382,
         n27381, n27380, n27379, n27378, n27377, n27376, n27375, n27374,
         n27373, n27372, n27371, n27370, n27369, n27368, n27367, n27366,
         n27365, n27364, n27363, n27362, n27361, n27360, n27359, n27358,
         n27357, n27356, n27355, n27354, n27353, n27352, n27351, n27350,
         n27349, n27348, n27347, n27346, n27345, n27344, n27343, n27342,
         n27341, n27340, n27339, n27338, n27337, n27336, n27335, n27334,
         n27333, n27332, n27331, n27330, n27329, n27328, n27327, n27326,
         n27325, n27324, n27323, n27322, n27321, n27320, n27319, n27318,
         n27317, n27316, n27315, n27314, n27313, n27312, n27311, n27310,
         n27309, n27308, n27307, n27306, n27305, n27304, n27303, n27302,
         n27301, n27300, n27299, n27298, n27297, n27296, n27295, n27294,
         n27293, n27292, n27291, n27290, n27289, n27288, n27287, n27286,
         n27285, n27284, n27283, n27282, n27281, n27280, n27279, n27278,
         n27277, n27276, n27275, n27274, n27273, n27272, n27271, n27270,
         n27269, n27268, n27267, n27266, n27265, n27264, n27263, n27262,
         n27261, n27260, n27259, n27258, n27257, n27256, n27255, n27254,
         n27253, n27252, n27251, n27250, n27249, n27248, n27247, n27246,
         n27245, n27244, n27243, n27242, n27241, n27240, n27239, n27238,
         n27237, n27236, n27235, n27234, n27233, n27232, n27231, n27230,
         n27229, n27228, n27227, n27226, n27225, n27224, n27223, n27222,
         n27221, n27220, n27219, n27218, n27217, n27216, n27215, n27214,
         n27213, n27212, n27211, n27210, n27209, n27208, n27207, n27206,
         n27205, n27204, n27203, n27202, n27201, n27200, n27199, n27198,
         n27197, n27196, n27195, n27194, n27193, n27192, n27191, n27190,
         n27189, n27188, n27187, n27186, n27185, n27184, n27183, n27182,
         n27181, n27180, n27179, n27178, n27177, n27176, n27175, n27174,
         n27173, n27172, n27171, n27170, n27169, n27168, n27167, n27166,
         n27165, n27164, n27163, n27162, n27161, n27160, n27159, n27158,
         n27157, n27156, n27155, n27154, n27153, n27152, n27151, n27150,
         n27149, n27148, n27147, n27146, n27145, n27144, n27143, n27142,
         n27141, n27140, n27139, n27138, n27137, n27136, n27135, n27134,
         n27133, n27132, n27131, n27130, n27129, n27128, n27127, n27126,
         n27125, n27124, n27123, n27122, n27121, n27120, n27119, n27118,
         n27117, n27116, n27115, n27114, n27113, n27112, n27111, n27110,
         n27109, n27108, n27107, n27106, n27105, n27104, n27103, n27102,
         n27101, n27100, n27099, n27098, n27097, n27096, n27095, n27094,
         n27093, n27092, n27091, n27090, n27089, n27088, n27087, n27086,
         n27085, n27084, n27083, n27082, n27081, n27080, n27079, n27078,
         n27077, n27076, n27075, n27074, n27073, n27072, n27071, n27070,
         n27069, n27068, n27067, n27066, n27065, n27064, n27063, n27062,
         n27061, n27060, n27059, n27058, n27057, n27056, n27055, n27054,
         n27053, n27052, n27051, n27050, n27049, n27048, n27047, n27046,
         n27045, n27044, n27043, n27042, n27041, n27040, n27039, n27038,
         n27037, n27036, n27035, n27034, n27033, n27032, n27031, n27030,
         n27029, n27028, n27027, n27026, n27025, n27024, n27023, n27022,
         n27021, n27020, n27019, n27018, n27017, n27016, n27015, n27014,
         n27013, n27012, n27011, n27010, n27009, n27008, n27007, n27006,
         n27005, n27004, n27003, n27002, n27001, n27000, n26999, n26998,
         n26997, n26996, n26995, n26994, n26993, n26992, n26991, n26990,
         n26989, n26988, n26987, n26986, n26985, n26984, n26983, n26982,
         n26981, n26980, n26979, n26978, n26977, n26976, n26975, n26974,
         n26973, n26972, n26971, n26970, n26969, n26968, n26967, n26966,
         n26965, n26964, n26963, n26962, n26961, n26960, n26959, n26958,
         n26957, n26956, n26955, n26954, n26953, n26952, n26951, n26950,
         n26949, n26948, n26947, n26946, n26945, n26944, n26943, n26942,
         n26941, n26940, n26939, n26938, n26937, n26936, n26935, n26934,
         n26933, n26932, n26931, n26930, n26929, n26928, n26927, n26926,
         n26925, n26924, n26923, n26922, n26921, n26920, n26919, n26918,
         n26917, n26916, n26915, n26914, n26913, n26912, n26911, n26910,
         n26909, n26908, n26907, n26906, n26905, n26904, n26903, n26902,
         n26901, n26900, n26899, n26898, n26897, n26896, n26895, n26894,
         n26893, n26892, n26891, n26890, n26889, n26888, n26887, n26886,
         n26885, n26884, n26883, n26882, n26881, n26880, n26879, n26878,
         n26877, n26876, n26875, n26874, n26873, n26872, n26871, n26870,
         n26869, n26868, n26867, n26866, n26865, n26864, n26863, n26862,
         n26861, n26860, n26859, n26858, n26857, n26856, n26855, n26854,
         n26853, n26852, n26851, n26850, n26849, n26848, n26847, n26846,
         n26845, n26844, n26843, n26842, n26841, n26840, n26839, n26838,
         n26837, n26836, n26835, n26834, n26833, n26832, n26831, n26830,
         n26829, n26828, n26827, n26826, n26825, n26824, n26823, n26822,
         n26821, n26820, n26819, n26818, n26817, n26816, n26815, n26814,
         n26813, n26812, n26811, n26810, n26809, n26808, n26807, n26806,
         n26805, n26804, n26803, n26802, n26801, n26800, n26799, n26798,
         n26797, n26796, n26795, n26794, n26793, n26792, n26791, n26790,
         n26789, n26788, n26787, n26786, n26785, n26784, n26783, n26782,
         n26781, n26780, n26779, n26778, n26777, n26776, n26775, n26774,
         n26773, n26772, n26771, n26770, n26769, n26768, n26767, n26766,
         n26765, n26764, n26763, n26762, n26761, n26760, n26759, n26758,
         n26757, n26756, n26755, n26754, n26753, n26752, n26751, n26750,
         n26749, n26748, n26747, n26746, n26745, n26744, n26743, n26742,
         n26741, n26740, n26739, n26738, n26737, n26736, n26735, n26734,
         n26733, n26732, n26731, n26730, n26729, n26728, n26727, n26726,
         n26725, n26724, n26723, n26722, n26721, n26720, n26719, n26718,
         n26717, n26716, n26715, n26714, n26713, n26712, n26711, n26710,
         n26709, n26708, n26707, n26706, n26705, n26704, n26703, n26702,
         n26701, n26700, n26699, n26698, n26697, n26696, n26695, n26694,
         n26693, n26692, n26691, n26690, n26689, n26688, n26687, n26686,
         n26685, n26684, n26683, n26682, n26681, n26680, n26679, n26678,
         n26677, n26676, n26675, n26674, n26673, n26672, n26671, n26670,
         n26669, n26668, n26667, n26666, n26665, n26664, n26663, n26662,
         n26661, n26660, n26659, n26658, n26657, n26656, n26655, n26654,
         n26653, n26652, n26651, n26650, n26649, n26648, n26646, n26645,
         n26644, n26643, n26642, n26641, n26640, n26639, n26638, n26637,
         n26636, n26635, n26634, n26633, n26632, n26631, n26630, n26629,
         n26628, n26627, n26626, n26625, n26624, n26623, n26622, n26621,
         n26620, n26619, n26618, n26617, n26616, n26615, n26614, n26613,
         n26612, n26611, n26610, n26609, n26608, n26607, n26606, n26605,
         n26604, n26603, n26602, n26601, n26600, n26599, n26598, n26597,
         n26596, n26595, n26594, n26593, n26592, n26591, n26590, n26589,
         n26588, n26587, n26586, n26585, n26584, n26583, n26582, n26581,
         n26580, n26579, n26578, n26577, n26576, n26575, n26574, n26573,
         n26572, n26571, n26570, n26569, n26568, n26567, n26566, n26565,
         n26564, n26563, n26562, n26561, n26560, n26559, n26558, n26557,
         n26556, n26555, n26554, n26553, n26552, n26551, n26550, n26549,
         n26548, n26547, n26546, n26545, n26544, n26543, n26542, n26541,
         n26540, n26539, n26538, n26537, n26536, n26535, n26534, n26533,
         n26532, n26531, n26530, n26529, n26528, n26527, n26526, n26525,
         n26524, n26523, n26522, n26521, n26520, n26519, n26518, n26517,
         n26516, n26515, n26514, n26513, n26512, n26511, n26510, n26509,
         n26508, n26507, n26506, n26505, n26504, n26503, n26502, n26501,
         n26500, n26499, n26498, n26497, n26496, n26495, n26494, n26493,
         n26492, n26491, n26490, n26489, n26488, n26487, n26486, n26485,
         n26484, n26483, n26482, n26481, n26480, n26479, n26478, n26476,
         n26475, n26474, n26473, n26472, n26471, n26470, n26469, n26468,
         n26467, n26466, n26465, n26464, n26463, n26462, n26461, n26460,
         n26459, n26458, n26457, n26456, n26455, n26454, n26453, n26452,
         n26451, n26450, n26449, n26448, n26447, n26446, n26445, n26444,
         n26443, n26442, n26441, n26440, n26439, n26438, n26437, n26436,
         n26435, n26434, n26433, n26432, n26431, n26430, n26429, n26428,
         n26427, n26426, n26425, n26424, n26423, n26422, n26421, n26420,
         n26419, n26418, n26417, n26416, n26415, n26414, n26413, n26412,
         n26411, n26410, n26409, n26408, n26407, n26406, n26405, n26404,
         n26403, n26402, n26401, n26400, n26399, n26398, n26397, n26396,
         n26395, n26394, n26393, n26392, n26391, n26390, n26389, n26388,
         n26387, n26386, n26385, n26384, n26383, n26382, n26381, n26380,
         n26379, n26378, n26377, n26376, n26375, n26374, n26373, n26372,
         n26371, n26370, n26368, n26367, n26366, n26365, n26364, n26363,
         n26362, n26361, n26360, n26359, n26358, n26357, n26356, n26355,
         n26354, n26353, n26352, n26351, n26350, n26349, n26348, n26347,
         n26346, n26345, n26344, n26343, n26342, n26341, n26340, n26339,
         n26338, n26337, n26336, n26335, n26334, n26333, n26332, n26331,
         n26330, n26329, n26328, n26327, n26326, n26325, n26324, n26323,
         n26322, n26321, n26320, n26319, n26318, n26317, n26316, n26315,
         n26314, n26313, n26312, n26311, n26310, n26309, n26308, n26307,
         n26306, n26305, n26304, n26303, n26302, n26301, n26300, n26299,
         n26298, n26297, n26296, n26295, n26294, n26293, n26292, n26291,
         n26290, n26289, n26288, n26287, n26286, n26285, n26284, n26283,
         n26282, n26281, n26280, n26279, n26278, n26277, n26276, n26275,
         n26274, n26273, n26272, n26271, n26270, n26269, n26268, n26267,
         n26266, n26265, n26264, n26263, n26262, n26261, n26260, n26259,
         n26258, n26257, n26256, n26255, n26254, n26253, n26252, n26251,
         n26250, n26249, n26248, n26247, n26246, n26245, n26244, n26243,
         n26242, n26241, n26240, n26239, n26238, n26237, n26236, n26235,
         n26234, n26233, n26232, n26231, n26230, n26229, n26228, n26227,
         n26226, n26225, n26224, n26223, n26222, n26221, n26220, n26219,
         n26218, n26217, n26216, n26215, n26214, n26213, n26212, n26211,
         n26210, n26209, n26208, n26207, n26206, n26205, n26204, n26203,
         n26202, n26201, n26200, n26199, n26198, n26197, n26196, n26195,
         n26194, n26193, n26192, n26191, n26190, n26189, n26188, n26187,
         n26186, n26185, n26184, n26183, n26182, n26181, n26180, n26179,
         n26178, n26177, n26176, n26175, n26174, n26173, n26172, n26171,
         n26170, n26169, n26168, n26167, n26166, n26165, n26164, n26163,
         n26162, n26161, n26160, n26159, n26158, n26157, n26156, n26155,
         n26154, n26153, n26152, n26151, n26150, n26149, n26148, n26147,
         n26146, n26145, n26144, n26143, n26142, n26141, n26140, n26139,
         n26138, n26137, n26136, n26135, n26134, n26133, n26132, n26131,
         n26130, n26129, n26128, n26127, n26126, n26125, n26124, n26123,
         n26122, n26121, n26120, n26119, n26118, n26117, n26116, n26115,
         n26114, n26113, n26112, n26111, n26110, n26109, n26108, n26107,
         n26106, n26105, n26104, n26103, n26102, n26101, n26100, n26099,
         n26098, n26097, n26096, n26095, n26094, n26093, n26092, n26091,
         n26090, n26089, n26088, n26087, n26086, n26085, n26084, n26083,
         n26082, n26081, n26080, n26079, n26078, n26077, n26076, n26075,
         n26074, n26073, n26072, n26071, n26070, n26069, n26068, n26067,
         n26066, n26065, n26064, n26063, n26062, n26061, n26060, n26059,
         n26058, n26057, n26056, n26055, n26054, n26053, n26052, n26051,
         n26050, n26049, n26048, n26047, n26046, n26045, n26044, n26043,
         n26042, n26041, n26040, n26039, n26038, n26037, n26036, n26035,
         n26034, n26033, n26032, n26031, n26030, n26029, n26028, n26027,
         n26026, n26025, n26024, n26022, n26021, n26020, n26019, n26018,
         n26017, n26016, n26015, n26014, n26013, n26012, n26011, n26010,
         n26009, n26008, n26007, n26006, n26005, n26004, n26003, n26002,
         n26001, n26000, n25999, n25998, n25997, n25996, n25995, n25994,
         n25993, n25992, n25991, n25990, n25989, n25988, n25987, n25986,
         n25985, n25984, n25983, n25982, n25981, n25980, n25979, n25978,
         n25977, n25976, n25975, n25974, n25973, n25972, n25971, n25970,
         n25969, n25968, n25967, n25966, n25965, n25964, n25963, n25962,
         n25961, n25960, n25959, n25958, n25957, n25956, n25955, n25954,
         n25953, n25952, n25951, n25950, n25949, n25948, n25947, n25946,
         n25945, n25944, n25943, n25942, n25941, n25940, n25939, n25938,
         n25937, n25936, n25935, n25934, n25933, n25932, n25931, n25930,
         n25929, n25928, n25927, n25926, n25925, n25924, n25923, n25921,
         n25920, n25919, n25918, n25917, n25916, n25915, n25914, n25913,
         n25912, n25911, n25910, n25909, n25908, n25907, n25906, n25905,
         n25904, n25903, n25902, n25901, n25900, n25899, n25898, n25897,
         n25896, n25895, n25894, n25893, n25892, n25891, n25890, n25889,
         n25888, n25887, n25886, n25885, n25884, n25883, n25882, n25881,
         n25880, n25879, n25878, n25877, n25876, n25875, n25874, n25873,
         n25872, n25871, n25870, n25869, n25868, n25867, n25866, n25865,
         n25864, n25863, n25862, n25861, n25860, n25859, n25858, n25857,
         n25856, n25855, n25854, n25853, n25852, n25851, n25850, n25849,
         n25848, n25847, n25846, n25845, n25844, n25843, n25842, n25841,
         n25840, n25839, n25838, n25837, n25836, n25835, n25834, n25833,
         n25832, n25831, n25830, n25829, n25828, n25827, n25826, n25825,
         n25824, n25823, n25822, n25821, n25820, n25819, n25818, n25817,
         n25816, n25815, n25814, n25813, n25812, n25811, n25810, n25808,
         n25807, n25806, n25805, n25804, n25803, n25802, n25801, n25800,
         n25799, n25798, n25797, n25796, n25795, n25794, n25793, n25792,
         n25791, n25790, n25789, n25788, n25787, n25786, n25785, n25784,
         n25783, n25782, n25781, n25780, n25779, n25778, n25777, n25776,
         n25775, n25774, n25773, n25772, n25771, n25770, n25769, n25768,
         n25767, n25766, n25765, n25764, n25763, n25762, n25761, n25760,
         n25759, n25758, n25757, n25756, n25755, n25754, n25753, n25752,
         n25751, n25750, n25749, n25748, n25747, n25746, n25745, n25744,
         n25743, n25742, n25741, n25740, n25739, n25738, n25737, n25736,
         n25735, n25734, n25733, n25732, n25731, n25730, n25729, n25728,
         n25727, n25726, n25725, n25724, n25723, n25722, n25721, n25720,
         n25719, n25718, n25717, n25716, n25715, n25714, n25713, n25712,
         n25711, n25710, n25709, n25708, n25707, n25706, n25705, n25704,
         n25703, n25702, n25701, n25700, n25699, n25698, n25697, n25696,
         n25695, n25694, n25693, n25692, n25691, n25690, n25689, n25688,
         n25687, n25686, n25685, n25684, n25683, n25682, n25681, n25680,
         n25679, n25678, n25677, n25676, n25675, n25674, n25673, n25672,
         n25671, n25670, n25669, n25668, n25667, n25666, n25665, n25664,
         n25663, n25662, n25661, n25660, n25659, n25658, n25657, n25656,
         n25655, n25654, n25653, n25652, n25651, n25650, n25649, n25648,
         n25647, n25646, n25645, n25644, n25643, n25642, n25641, n25640,
         n25639, n25638, n25637, n25636, n25635, n25634, n25633, n25632,
         n25631, n25630, n25629, n25628, n25627, n25626, n25625, n25624,
         n25623, n25622, n25621, n25620, n25619, n25618, n25617, n25616,
         n25615, n25614, n25613, n25612, n25611, n25610, n25609, n25608,
         n25607, n25606, n25605, n25604, n25603, n25602, n25601, n25600,
         n25599, n25598, n25597, n25596, n25595, n25594, n25593, n25592,
         n25591, n25590, n25589, n25588, n25587, n25586, n25585, n25584,
         n25583, n25582, n25581, n25580, n25579, n25578, n25577, n25576,
         n25575, n25574, n25573, n25572, n25571, n25570, n25569, n25568,
         n25567, n25566, n25565, n25564, n25563, n25562, n25561, n25560,
         n25559, n25558, n25557, n25556, n25555, n25554, n25553, n25552,
         n25551, n25550, n25549, n25548, n25547, n25546, n25545, n25544,
         n25543, n25542, n25541, n25540, n25539, n25538, n25537, n25536,
         n25535, n25534, n25533, n25531, n25530, n25529, n25528, n25527,
         n25526, n25525, n25524, n25523, n25522, n25521, n25520, n25519,
         n25518, n25517, n25516, n25515, n25514, n25513, n25512, n25511,
         n25510, n25509, n25508, n25507, n25506, n25505, n25504, n25503,
         n25502, n25501, n25500, n25499, n25498, n25497, n25496, n25495,
         n25494, n25493, n25492, n25491, n25490, n25489, n25488, n25487,
         n25486, n25485, n25484, n25483, n25482, n25481, n25480, n25479,
         n25478, n25477, n25476, n25475, n25474, n25473, n25472, n25471,
         n25470, n25469, n25468, n25467, n25466, n25465, n25464, n25463,
         n25462, n25461, n25460, n25459, n25458, n25457, n25456, n25455,
         n25454, n25453, n25452, n25451, n25450, n25449, n25448, n25447,
         n25446, n25445, n25444, n25443, n25442, n25441, n25440, n25439,
         n25438, n25437, n25436, n25435, n25434, n25433, n25432, n25431,
         n25430, n25429, n25428, n25427, n25426, n25425, n25424, n25423,
         n25422, n25421, n25420, n25419, n25418, n25417, n25416, n25415,
         n25414, n25413, n25412, n25411, n25410, n25409, n25408, n25407,
         n25406, n25405, n25404, n25403, n25402, n25401, n25400, n25399,
         n25398, n25397, n25396, n25395, n25394, n25393, n25392, n25391,
         n25390, n25389, n25388, n25387, n25386, n25385, n25384, n25383,
         n25382, n25381, n25380, n25379, n25378, n25377, n25376, n25375,
         n25374, n25373, n25372, n25371, n25370, n25369, n25368, n25367,
         n25366, n25365, n25364, n25363, n25362, n25360, n25359, n25358,
         n25357, n25356, n25355, n25354, n25353, n25352, n25351, n25350,
         n25349, n25348, n25347, n25346, n25345, n25344, n25343, n25342,
         n25341, n25340, n25339, n25338, n25337, n25336, n25335, n25334,
         n25333, n25332, n25331, n25330, n25329, n25328, n25327, n25326,
         n25325, n25324, n25323, n25322, n25321, n25320, n25319, n25318,
         n25317, n25316, n25315, n25314, n25313, n25312, n25311, n25310,
         n25309, n25308, n25307, n25306, n25305, n25304, n25303, n25302,
         n25301, n25300, n25299, n25298, n25297, n25296, n25295, n25294,
         n25293, n25292, n25291, n25290, n25289, n25288, n25287, n25286,
         n25285, n25284, n25283, n25282, n25281, n25280, n25279, n25278,
         n25277, n25276, n25275, n25274, n25273, n25272, n25271, n25270,
         n25269, n25268, n25267, n25266, n25265, n25264, n25263, n25262,
         n25261, n25260, n25259, n25258, n25257, n25256, n25255, n25254,
         n25252, n25251, n25250, n25249, n25248, n25247, n25246, n25245,
         n25244, n25243, n25242, n25241, n25240, n25239, n25238, n25237,
         n25236, n25235, n25234, n25233, n25232, n25231, n25230, n25229,
         n25228, n25227, n25226, n25225, n25224, n25223, n25222, n25221,
         n25220, n25219, n25218, n25217, n25216, n25215, n25214, n25213,
         n25212, n25211, n25210, n25209, n25208, n25207, n25206, n25205,
         n25204, n25203, n25202, n25201, n25200, n25199, n25198, n25197,
         n25196, n25195, n25194, n25193, n25192, n25191, n25190, n25189,
         n25188, n25187, n25186, n25185, n25184, n25183, n25182, n25181,
         n25180, n25179, n25178, n25177, n25176, n25175, n25174, n25173,
         n25172, n25171, n25170, n25169, n25168, n25167, n25166, n25165,
         n25164, n25163, n25162, n25161, n25160, n25159, n25158, n25157,
         n25156, n25155, n25154, n25153, n25152, n25151, n25150, n25149,
         n25148, n25147, n25146, n25145, n25144, n25143, n25142, n25141,
         n25140, n25139, n25138, n25137, n25136, n25135, n25134, n25133,
         n25132, n25131, n25130, n25129, n25128, n25127, n25126, n25125,
         n25124, n25123, n25122, n25121, n25120, n25119, n25118, n25117,
         n25116, n25115, n25114, n25113, n25112, n25111, n25110, n25109,
         n25108, n25107, n25106, n25105, n25104, n25103, n25102, n25101,
         n25100, n25099, n25098, n25097, n25096, n25095, n25094, n25093,
         n25092, n25091, n25090, n25089, n25088, n25087, n25086, n25085,
         n25084, n25083, n25082, n25081, n25080, n25079, n25078, n25077,
         n25076, n25075, n25074, n25073, n25072, n25071, n25070, n25069,
         n25068, n25067, n25066, n25065, n25064, n25063, n25062, n25061,
         n25060, n25059, n25058, n25057, n25056, n25055, n25054, n25053,
         n25052, n25051, n25050, n25049, n25048, n25047, n25046, n25045,
         n25044, n25043, n25042, n25041, n25040, n25039, n25038, n25037,
         n25036, n25035, n25034, n25033, n25032, n25031, n25030, n25029,
         n25028, n25027, n25026, n25025, n25024, n25023, n25022, n25021,
         n25020, n25019, n25018, n25017, n25016, n25015, n25014, n25013,
         n25012, n25011, n25010, n25009, n25008, n25007, n25006, n25005,
         n25004, n25003, n25002, n25001, n25000, n24999, n24998, n24997,
         n24996, n24995, n24994, n24993, n24992, n24991, n24990, n24989,
         n24988, n24987, n24986, n24985, n24984, n24983, n24982, n24981,
         n24980, n24979, n24978, n24977, n24976, n24975, n24973, n24972,
         n24971, n24970, n24969, n24968, n24967, n24966, n24965, n24964,
         n24963, n24962, n24961, n24960, n24959, n24958, n24957, n24956,
         n24955, n24954, n24953, n24952, n24951, n24950, n24949, n24948,
         n24947, n24946, n24945, n24944, n24943, n24942, n24941, n24940,
         n24939, n24938, n24937, n24936, n24935, n24934, n24933, n24932,
         n24931, n24930, n24929, n24928, n24927, n24926, n24925, n24924,
         n24923, n24922, n24921, n24920, n24919, n24918, n24917, n24916,
         n24915, n24914, n24913, n24912, n24911, n24910, n24909, n24908,
         n24907, n24906, n24905, n24904, n24903, n24902, n24901, n24900,
         n24899, n24898, n24897, n24896, n24895, n24894, n24893, n24892,
         n24891, n24890, n24889, n24888, n24887, n24886, n24885, n24884,
         n24883, n24882, n24881, n24880, n24879, n24878, n24877, n24876,
         n24875, n24874, n24873, n24872, n24871, n24870, n24869, n24868,
         n24867, n24866, n24865, n24864, n24863, n24862, n24861, n24860,
         n24859, n24858, n24857, n24856, n24855, n24854, n24853, n24852,
         n24851, n24850, n24849, n24848, n24847, n24846, n24845, n24844,
         n24843, n24842, n24841, n24840, n24839, n24838, n24837, n24836,
         n24835, n24834, n24833, n24832, n24831, n24830, n24829, n24828,
         n24827, n24826, n24825, n24824, n24823, n24822, n24821, n24820,
         n24819, n24818, n24817, n24816, n24815, n24814, n24813, n24812,
         n24811, n24810, n24809, n24808, n24807, n24806, n24805, n24804,
         n24803, n24802, n24801, n24800, n24799, n24798, n24797, n24796,
         n24795, n24794, n24793, n24792, n24791, n24790, n24789, n24788,
         n24787, n24786, n24785, n24784, n24783, n24782, n24781, n24780,
         n24779, n24778, n24777, n24776, n24775, n24774, n24773, n24772,
         n24771, n24770, n24769, n24768, n24767, n24766, n24765, n24764,
         n24763, n24762, n24761, n24760, n24759, n24758, n24757, n24756,
         n24755, n24754, n24753, n24752, n24751, n24750, n24749, n24748,
         n24747, n24746, n24745, n24744, n24743, n24742, n24741, n24740,
         n24739, n24738, n24737, n24736, n24735, n24734, n24733, n24732,
         n24731, n24730, n24729, n24728, n24727, n24726, n24725, n24724,
         n24723, n24722, n24721, n24720, n24719, n24718, n24717, n24716,
         n24715, n24714, n24713, n24712, n24711, n24710, n24709, n24708,
         n24707, n24706, n24705, n24704, n24703, n24702, n24701, n24700,
         n24699, n24698, n24697, n24696, n24694, n24693, n24692, n24691,
         n24690, n24689, n24688, n24687, n24686, n24685, n24684, n24683,
         n24682, n24681, n24680, n24679, n24678, n24677, n24676, n24675,
         n24674, n24673, n24672, n24671, n24670, n24669, n24668, n24667,
         n24666, n24665, n24664, n24663, n24662, n24661, n24660, n24659,
         n24658, n24657, n24656, n24655, n24654, n24653, n24652, n24651,
         n24650, n24649, n24648, n24647, n24646, n24645, n24644, n24643,
         n24642, n24641, n24640, n24639, n24638, n24637, n24636, n24635,
         n24634, n24633, n24632, n24631, n24630, n24629, n24628, n24627,
         n24626, n24625, n24624, n24623, n24622, n24621, n24620, n24619,
         n24618, n24617, n24616, n24615, n24614, n24613, n24612, n24611,
         n24610, n24609, n24608, n24607, n24606, n24605, n24604, n24603,
         n24602, n24601, n24600, n24599, n24598, n24597, n24596, n24595,
         n24594, n24593, n24592, n24591, n24590, n24589, n24588, n24587,
         n24586, n24585, n24584, n24583, n24582, n24581, n24580, n24579,
         n24578, n24577, n24576, n24575, n24574, n24573, n24572, n24571,
         n24570, n24569, n24568, n24567, n24566, n24565, n24564, n24563,
         n24562, n24561, n24560, n24559, n24558, n24557, n24556, n24555,
         n24554, n24553, n24552, n24551, n24550, n24549, n24548, n24547,
         n24546, n24545, n24544, n24543, n24542, n24541, n24540, n24539,
         n24538, n24537, n24536, n24535, n24534, n24533, n24532, n24531,
         n24530, n24529, n24528, n24527, n24526, n24525, n24524, n24523,
         n24522, n24521, n24520, n24519, n24518, n24517, n24516, n24515,
         n24514, n24513, n24512, n24511, n24510, n24509, n24508, n24507,
         n24506, n24505, n24504, n24503, n24502, n24501, n24500, n24499,
         n24498, n24497, n24496, n24495, n24494, n24493, n24492, n24491,
         n24490, n24489, n24488, n24487, n24486, n24485, n24484, n24483,
         n24482, n24481, n24480, n24479, n24478, n24477, n24476, n24475,
         n24474, n24473, n24472, n24471, n24470, n24469, n24468, n24467,
         n24466, n24465, n24464, n24463, n24462, n24461, n24460, n24459,
         n24458, n24457, n24456, n24455, n24454, n24453, n24452, n24451,
         n24450, n24449, n24448, n24447, n24446, n24445, n24444, n24443,
         n24442, n24441, n24440, n24439, n24438, n24437, n24436, n24435,
         n24434, n24433, n24432, n24431, n24430, n24429, n24428, n24427,
         n24426, n24425, n24424, n24423, n24422, n24421, n24420, n24419,
         n24418, n24416, n24415, n24414, n24413, n24412, n24411, n24410,
         n24409, n24408, n24407, n24406, n24405, n24404, n24403, n24402,
         n24401, n24400, n24399, n24398, n24397, n24396, n24395, n24394,
         n24393, n24392, n24391, n24390, n24389, n24388, n24387, n24386,
         n24385, n24384, n24383, n24382, n24381, n24380, n24379, n24378,
         n24377, n24376, n24375, n24374, n24373, n24372, n24371, n24370,
         n24369, n24368, n24367, n24366, n24365, n24364, n24363, n24362,
         n24361, n24360, n24359, n24358, n24357, n24356, n24355, n24354,
         n24353, n24352, n24351, n24350, n24349, n24348, n24347, n24346,
         n24345, n24344, n24343, n24342, n24341, n24340, n24339, n24338,
         n24337, n24336, n24335, n24334, n24333, n24332, n24331, n24330,
         n24329, n24328, n24327, n24326, n24325, n24324, n24323, n24322,
         n24321, n24320, n24319, n24318, n24317, n24316, n24315, n24314,
         n24313, n24312, n24311, n24310, n24309, n24308, n24307, n24306,
         n24305, n24304, n24303, n24302, n24301, n24300, n24299, n24298,
         n24297, n24296, n24295, n24294, n24293, n24292, n24291, n24290,
         n24289, n24288, n24287, n24286, n24285, n24284, n24283, n24282,
         n24281, n24280, n24279, n24278, n24277, n24276, n24275, n24274,
         n24273, n24272, n24271, n24270, n24269, n24268, n24267, n24266,
         n24265, n24264, n24263, n24262, n24261, n24260, n24259, n24258,
         n24257, n24256, n24255, n24254, n24253, n24252, n24251, n24250,
         n24249, n24248, n24247, n24245, n24244, n24243, n24242, n24241,
         n24240, n24239, n24238, n24237, n24236, n24235, n24234, n24233,
         n24232, n24231, n24230, n24229, n24228, n24227, n24226, n24225,
         n24224, n24223, n24222, n24221, n24220, n24219, n24218, n24217,
         n24216, n24215, n24214, n24213, n24212, n24211, n24210, n24209,
         n24208, n24207, n24206, n24205, n24204, n24203, n24202, n24201,
         n24200, n24199, n24198, n24197, n24196, n24195, n24194, n24193,
         n24192, n24191, n24190, n24189, n24188, n24187, n24186, n24185,
         n24184, n24183, n24182, n24181, n24180, n24179, n24178, n24177,
         n24176, n24175, n24174, n24173, n24172, n24171, n24170, n24169,
         n24168, n24167, n24166, n24165, n24164, n24163, n24162, n24161,
         n24160, n24159, n24158, n24157, n24156, n24155, n24154, n24153,
         n24152, n24151, n24150, n24149, n24148, n24147, n24146, n24145,
         n24144, n24143, n24142, n24141, n24140, n24139, n24137, n24136,
         n24135, n24134, n24133, n24132, n24131, n24130, n24129, n24128,
         n24127, n24126, n24125, n24124, n24123, n24122, n24121, n24120,
         n24119, n24118, n24117, n24116, n24115, n24114, n24113, n24112,
         n24111, n24110, n24109, n24108, n24107, n24106, n24105, n24104,
         n24103, n24102, n24101, n24100, n24099, n24098, n24097, n24096,
         n24095, n24094, n24093, n24092, n24091, n24090, n24089, n24088,
         n24087, n24086, n24085, n24084, n24083, n24082, n24081, n24080,
         n24079, n24078, n24077, n24076, n24075, n24074, n24073, n24072,
         n24071, n24070, n24069, n24068, n24067, n24066, n24065, n24064,
         n24063, n24062, n24061, n24060, n24059, n24058, n24057, n24056,
         n24055, n24054, n24053, n24052, n24051, n24050, n24049, n24048,
         n24047, n24046, n24045, n24044, n24043, n24042, n24041, n24040,
         n24039, n24038, n24037, n24036, n24035, n24034, n24033, n24032,
         n24031, n24030, n24029, n24028, n24027, n24026, n24025, n24024,
         n24023, n24022, n24021, n24020, n24019, n24018, n24017, n24016,
         n24015, n24014, n24013, n24012, n24011, n24010, n24009, n24008,
         n24007, n24006, n24005, n24004, n24003, n24002, n24001, n24000,
         n23999, n23998, n23997, n23996, n23995, n23994, n23993, n23992,
         n23991, n23990, n23989, n23988, n23987, n23986, n23985, n23984,
         n23983, n23982, n23981, n23980, n23979, n23978, n23977, n23976,
         n23975, n23974, n23973, n23972, n23971, n23970, n23969, n23968,
         n23966, n23965, n23964, n23963, n23962, n23961, n23960, n23959,
         n23958, n23957, n23956, n23955, n23954, n23953, n23952, n23951,
         n23950, n23949, n23948, n23947, n23946, n23945, n23944, n23943,
         n23942, n23941, n23940, n23939, n23938, n23937, n23936, n23935,
         n23934, n23933, n23932, n23931, n23930, n23929, n23928, n23927,
         n23926, n23925, n23924, n23923, n23922, n23921, n23920, n23919,
         n23918, n23917, n23916, n23915, n23914, n23913, n23912, n23911,
         n23910, n23909, n23908, n23907, n23906, n23905, n23904, n23903,
         n23902, n23901, n23900, n23899, n23898, n23897, n23896, n23895,
         n23894, n23893, n23892, n23891, n23890, n23889, n23888, n23887,
         n23886, n23885, n23884, n23883, n23882, n23881, n23880, n23879,
         n23878, n23877, n23876, n23875, n23874, n23873, n23872, n23871,
         n23870, n23869, n23868, n23867, n23866, n23865, n23864, n23863,
         n23862, n23861, n23860, n23858, n23857, n23856, n23855, n23854,
         n23853, n23852, n23851, n23850, n23849, n23848, n23847, n23846,
         n23845, n23844, n23843, n23842, n23841, n23840, n23839, n23838,
         n23837, n23836, n23835, n23834, n23833, n23832, n23831, n23830,
         n23829, n23828, n23827, n23826, n23825, n23824, n23823, n23821,
         n23820, n23819, n23818, n23817, n23816, n23815, n23814, n23813,
         n23812, n23811, n23810, n23809, n23808, n23807, n23806, n23805,
         n23804, n23803, n23802, n23801, n23800, n23799, n23798, n23797,
         n23796, n23795, n23794, n23793, n23792, n23791, n23790, n23789,
         n23788, n23787, n23786, n23785, n23784, n23783, n23782, n23781,
         n23780, n23779, n23778, n23777, n23776, n23775, n23774, n23773,
         n23772, n23771, n23770, n23769, n23768, n23767, n23766, n23765,
         n23764, n23763, n23762, n23761, n23760, n23759, n23758, n23757,
         n23756, n23755, n23754, n23753, n23752, n23751, n23750, n23749,
         n23748, n23747, n23746, n23745, n23744, n23743, n23742, n23741,
         n23740, n23739, n23738, n23737, n23736, n23735, n23734, n23733,
         n23732, n23731, n23730, n23729, n23728, n23727, n23726, n23725,
         n23724, n23723, n23722, n23721, n23720, n23719, n23718, n23717,
         n23716, n23715, n23714, n23713, n23712, n23711, n23710, n23709,
         n23708, n23707, n23706, n23705, n23704, n23703, n23702, n23701,
         n23700, n23699, n23698, n23697, n23696, n23695, n23694, n23693,
         n23692, n23691, n23690, n23689, n23687, n23686, n23685, n23684,
         n23683, n23682, n23681, n23680, n23679, n23678, n23677, n23676,
         n23675, n23674, n23673, n23672, n23671, n23670, n23669, n23668,
         n23667, n23666, n23665, n23664, n23663, n23662, n23661, n23660,
         n23659, n23658, n23657, n23656, n23655, n23654, n23653, n23652,
         n23651, n23650, n23649, n23648, n23647, n23646, n23645, n23644,
         n23643, n23642, n23641, n23640, n23639, n23638, n23637, n23636,
         n23635, n23634, n23633, n23632, n23631, n23630, n23629, n23628,
         n23627, n23626, n23625, n23624, n23623, n23622, n23621, n23620,
         n23619, n23618, n23617, n23616, n23615, n23614, n23613, n23612,
         n23611, n23610, n23609, n23608, n23607, n23606, n23605, n23604,
         n23603, n23602, n23601, n23600, n23599, n23598, n23597, n23596,
         n23595, n23594, n23593, n23592, n23591, n23590, n23589, n23588,
         n23587, n23586, n23585, n23584, n23583, n23582, n23581, n23579,
         n23578, n23577, n23576, n23575, n23574, n23573, n23572, n23571,
         n23570, n23569, n23568, n23567, n23566, n23565, n23564, n23563,
         n23562, n23561, n23560, n23559, n23558, n23557, n23556, n23555,
         n23554, n23553, n23552, n23551, n23550, n23549, n23548, n23547,
         n23546, n23545, n23544, n23543, n23542, n23541, n23540, n23539,
         n23538, n23537, n23536, n23535, n23534, n23533, n23532, n23531,
         n23530, n23529, n23528, n23527, n23526, n23525, n23524, n23523,
         n23522, n23521, n23520, n23519, n23518, n23517, n23516, n23515,
         n23514, n23513, n23512, n23511, n23510, n23509, n23508, n23507,
         n23506, n23505, n23504, n23503, n23502, n23501, n23500, n23499,
         n23498, n23497, n23496, n23495, n23494, n23493, n23492, n23491,
         n23490, n23489, n23488, n23487, n23486, n23485, n23484, n23483,
         n23482, n23481, n23480, n23479, n23478, n23477, n23476, n23475,
         n23474, n23473, n23472, n23471, n23470, n23469, n23468, n23467,
         n23466, n23465, n23464, n23463, n23462, n23461, n23460, n23459,
         n23458, n23457, n23456, n23455, n23454, n23453, n23452, n23451,
         n23450, n23449, n23448, n23447, n23446, n23445, n23444, n23443,
         n23442, n23441, n23440, n23439, n23438, n23437, n23436, n23435,
         n23434, n23433, n23432, n23431, n23430, n23429, n23428, n23427,
         n23426, n23425, n23424, n23423, n23422, n23421, n23420, n23419,
         n23418, n23417, n23416, n23415, n23414, n23413, n23412, n23411,
         n23410, n23409, n23408, n23407, n23406, n23405, n23404, n23403,
         n23402, n23401, n23400, n23399, n23398, n23397, n23396, n23395,
         n23394, n23393, n23392, n23391, n23390, n23389, n23388, n23387,
         n23386, n23385, n23384, n23383, n23382, n23381, n23380, n23379,
         n23378, n23377, n23376, n23375, n23374, n23373, n23372, n23371,
         n23370, n23369, n23368, n23367, n23366, n23365, n23364, n23363,
         n23362, n23361, n23360, n23359, n23358, n23357, n23356, n23355,
         n23354, n23353, n23352, n23351, n23350, n23349, n23348, n23347,
         n23346, n23345, n23344, n23343, n23342, n23341, n23340, n23339,
         n23338, n23337, n23336, n23335, n23334, n23333, n23332, n23331,
         n23330, n23329, n23328, n23327, n23326, n23325, n23324, n23323,
         n23322, n23321, n23320, n23319, n23318, n23317, n23316, n23315,
         n23314, n23313, n23312, n23311, n23310, n23309, n23308, n23307,
         n23306, n23305, n23304, n23303, n23302, n23300, n23299, n23298,
         n23297, n23296, n23295, n23294, n23293, n23292, n23291, n23290,
         n23289, n23288, n23287, n23286, n23285, n23284, n23283, n23282,
         n23281, n23280, n23279, n23278, n23277, n23276, n23275, n23274,
         n23273, n23272, n23271, n23270, n23269, n23268, n23267, n23266,
         n23265, n23264, n23263, n23262, n23261, n23260, n23259, n23258,
         n23257, n23256, n23255, n23254, n23253, n23252, n23251, n23250,
         n23249, n23248, n23247, n23246, n23245, n23244, n23243, n23242,
         n23241, n23240, n23239, n23238, n23237, n23236, n23235, n23234,
         n23233, n23232, n23231, n23230, n23229, n23228, n23227, n23226,
         n23225, n23224, n23223, n23222, n23221, n23220, n23219, n23218,
         n23217, n23216, n23215, n23214, n23213, n23212, n23211, n23210,
         n23209, n23208, n23207, n23206, n23205, n23204, n23203, n23202,
         n23201, n23200, n23199, n23198, n23197, n23196, n23195, n23194,
         n23193, n23192, n23191, n23190, n23189, n23188, n23187, n23186,
         n23185, n23184, n23183, n23182, n23181, n23180, n23179, n23178,
         n23177, n23176, n23175, n23174, n23173, n23172, n23171, n23170,
         n23169, n23168, n23167, n23166, n23165, n23164, n23163, n23162,
         n23161, n23160, n23159, n23158, n23157, n23156, n23155, n23154,
         n23153, n23152, n23151, n23150, n23149, n23148, n23147, n23146,
         n23145, n23144, n23143, n23142, n23141, n23140, n23139, n23138,
         n23137, n23136, n23135, n23134, n23133, n23132, n23131, n23130,
         n23128, n23127, n23126, n23125, n23124, n23123, n23122, n23121,
         n23120, n23119, n23118, n23117, n23116, n23115, n23114, n23113,
         n23112, n23111, n23110, n23109, n23108, n23107, n23106, n23105,
         n23104, n23103, n23102, n23101, n23100, n23099, n23098, n23097,
         n23096, n23095, n23094, n23093, n23092, n23091, n23090, n23089,
         n23088, n23087, n23086, n23085, n23084, n23083, n23082, n23081,
         n23080, n23079, n23078, n23077, n23076, n23075, n23074, n23073,
         n23072, n23071, n23070, n23069, n23068, n23067, n23066, n23065,
         n23064, n23063, n23062, n23061, n23060, n23059, n23058, n23057,
         n23056, n23055, n23054, n23053, n23052, n23051, n23050, n23049,
         n23048, n23047, n23046, n23045, n23044, n23043, n23042, n23041,
         n23040, n23039, n23038, n23037, n23036, n23035, n23034, n23033,
         n23032, n23031, n23030, n23029, n23028, n23027, n23026, n23025,
         n23024, n23023, n23022, n23020, n23019, n23018, n23017, n23016,
         n23015, n23014, n23013, n23012, n23011, n23010, n23009, n23008,
         n23007, n23006, n23005, n23004, n23003, n23002, n23001, n23000,
         n22999, n22998, n22997, n22996, n22995, n22994, n22993, n22992,
         n22991, n22990, n22989, n22988, n22987, n22986, n22985, n22984,
         n22983, n22982, n22981, n22980, n22979, n22978, n22977, n22976,
         n22975, n22974, n22973, n22972, n22971, n22970, n22969, n22968,
         n22967, n22966, n22965, n22964, n22963, n22962, n22961, n22960,
         n22959, n22958, n22957, n22956, n22955, n22954, n22953, n22952,
         n22951, n22950, n22949, n22948, n22947, n22946, n22945, n22944,
         n22943, n22942, n22941, n22940, n22939, n22938, n22937, n22936,
         n22935, n22934, n22933, n22932, n22931, n22930, n22929, n22928,
         n22927, n22926, n22925, n22924, n22923, n22922, n22921, n22920,
         n22919, n22918, n22917, n22916, n22915, n22914, n22913, n22912,
         n22911, n22910, n22909, n22908, n22907, n22906, n22905, n22904,
         n22903, n22902, n22901, n22900, n22899, n22898, n22897, n22896,
         n22895, n22894, n22893, n22892, n22891, n22890, n22889, n22888,
         n22887, n22886, n22885, n22884, n22883, n22882, n22881, n22880,
         n22879, n22878, n22877, n22876, n22875, n22874, n22873, n22872,
         n22871, n22870, n22869, n22868, n22867, n22866, n22865, n22864,
         n22863, n22862, n22861, n22860, n22859, n22858, n22857, n22856,
         n22855, n22854, n22853, n22851, n22850, n22849, n22848, n22847,
         n22846, n22845, n22844, n22843, n22842, n22841, n22840, n22839,
         n22838, n22837, n22836, n22835, n22834, n22833, n22832, n22831,
         n22830, n22829, n22828, n22827, n22826, n22825, n22824, n22823,
         n22822, n22821, n22820, n22819, n22818, n22817, n22816, n22815,
         n22814, n22813, n22812, n22811, n22810, n22809, n22808, n22807,
         n22806, n22805, n22804, n22803, n22802, n22801, n22800, n22799,
         n22798, n22797, n22796, n22795, n22794, n22793, n22792, n22791,
         n22790, n22789, n22788, n22787, n22786, n22785, n22784, n22783,
         n22782, n22781, n22780, n22779, n22778, n22777, n22776, n22775,
         n22774, n22773, n22772, n22771, n22770, n22769, n22768, n22767,
         n22766, n22765, n22764, n22763, n22762, n22761, n22760, n22759,
         n22758, n22757, n22756, n22755, n22754, n22753, n22752, n22751,
         n22750, n22749, n22748, n22747, n22746, n22745, n22744, n22743,
         n22742, n22741, n22740, n22739, n22738, n22737, n22736, n22735,
         n22734, n22733, n22732, n22731, n22730, n22729, n22728, n22727,
         n22726, n22725, n22724, n22723, n22722, n22721, n22720, n22719,
         n22718, n22717, n22716, n22715, n22714, n22713, n22712, n22711,
         n22710, n22709, n22708, n22707, n22706, n22705, n22704, n22703,
         n22702, n22701, n22700, n22699, n22698, n22697, n22696, n22695,
         n22694, n22693, n22692, n22691, n22690, n22689, n22688, n22687,
         n22686, n22685, n22684, n22683, n22682, n22681, n22680, n22679,
         n22678, n22677, n22676, n22675, n22674, n22673, n22672, n22671,
         n22670, n22669, n22668, n22667, n22666, n22665, n22664, n22663,
         n22662, n22661, n22660, n22659, n22658, n22657, n22656, n22655,
         n22654, n22653, n22652, n22651, n22650, n22649, n22648, n22647,
         n22646, n22645, n22644, n22643, n22642, n22641, n22640, n22639,
         n22638, n22637, n22636, n22635, n22634, n22633, n22632, n22631,
         n22630, n22629, n22628, n22627, n22626, n22625, n22624, n22623,
         n22622, n22621, n22620, n22619, n22618, n22617, n22616, n22615,
         n22614, n22613, n22612, n22611, n22610, n22609, n22608, n22607,
         n22606, n22605, n22604, n22603, n22602, n22601, n22600, n22599,
         n22598, n22597, n22596, n22595, n22594, n22593, n22592, n22591,
         n22590, n22589, n22588, n22587, n22586, n22585, n22584, n22583,
         n22582, n22581, n22580, n22579, n22578, n22577, n22576, n22575,
         n22574, n22573, n22572, n22571, n22570, n22569, n22568, n22567,
         n22566, n22565, n22564, n22563, n22562, n22561, n22560, n22559,
         n22558, n22557, n22556, n22555, n22554, n22553, n22552, n22551,
         n22550, n22549, n22548, n22547, n22546, n22545, n22544, n22543,
         n22542, n22541, n22540, n22539, n22538, n22537, n22536, n22535,
         n22534, n22533, n22532, n22531, n22530, n22529, n22528, n22527,
         n22526, n22525, n22524, n22523, n22522, n22521, n22520, n22519,
         n22518, n22517, n22516, n22515, n22514, n22513, n22512, n22511,
         n22510, n22509, n22508, n22507, n22506, n22505, n22504, n22503,
         n22502, n22501, n22500, n22499, n22498, n22497, n22496, n22495,
         n22494, n22493, n22492, n22491, n22490, n22489, n22488, n22487,
         n22486, n22485, n22484, n22483, n22482, n22481, n22480, n22479,
         n22478, n22477, n22476, n22475, n22474, n22473, n22472, n22471,
         n22470, n22469, n22468, n22467, n22466, n22465, n22464, n22463,
         n22462, n22461, n22460, n22459, n22458, n22457, n22456, n22455,
         n22454, n22453, n22452, n22451, n22450, n22449, n22447, n22446,
         n22445, n22444, n22443, n22442, n22441, n22440, n22439, n22438,
         n22437, n22436, n22435, n22434, n22433, n22432, n22431, n22430,
         n22429, n22428, n22427, n22426, n22425, n22424, n22423, n22422,
         n22421, n22420, n22419, n22418, n22417, n22416, n22415, n22414,
         n22413, n22412, n22411, n22410, n22409, n22408, n22407, n22406,
         n22405, n22404, n22403, n22402, n22401, n22400, n22399, n22398,
         n22397, n22396, n22395, n22394, n22393, n22392, n22391, n22390,
         n22389, n22388, n22387, n22386, n22385, n22384, n22383, n22382,
         n22381, n22380, n22379, n22378, n22377, n22376, n22375, n22374,
         n22373, n22372, n22371, n22370, n22369, n22368, n22367, n22366,
         n22365, n22364, n22363, n22362, n22361, n22360, n22359, n22358,
         n22357, n22356, n22355, n22354, n22353, n22352, n22351, n22350,
         n22349, n22348, n22347, n22346, n22345, n22344, n22343, n22342,
         n22341, n22340, n22339, n22338, n22337, n22336, n22335, n22334,
         n22333, n22332, n22331, n22330, n22329, n22328, n22327, n22326,
         n22325, n22324, n22323, n22322, n22321, n22320, n22319, n22318,
         n22317, n22316, n22315, n22314, n22313, n22312, n22311, n22310,
         n22309, n22308, n22307, n22306, n22305, n22304, n22303, n22302,
         n22301, n22300, n22299, n22298, n22297, n22296, n22295, n22294,
         n22293, n22292, n22291, n22290, n22289, n22288, n22287, n22286,
         n22285, n22284, n22283, n22282, n22281, n22280, n22279, n22278,
         n22277, n22276, n22275, n22274, n22273, n22272, n22271, n22270,
         n22269, n22268, n22267, n22266, n22265, n22264, n22263, n22262,
         n22261, n22260, n22259, n22258, n22257, n22256, n22255, n22254,
         n22253, n22252, n22251, n22250, n22249, n22248, n22247, n22246,
         n22245, n22244, n22243, n22242, n22241, n22240, n22239, n22238,
         n22237, n22236, n22235, n22234, n22233, n22232, n22231, n22230,
         n22229, n22228, n22227, n22226, n22225, n22224, n22223, n22222,
         n22221, n22220, n22219, n22218, n22217, n22216, n22215, n22214,
         n22213, n22212, n22211, n22210, n22209, n22208, n22207, n22206,
         n22205, n22204, n22203, n22202, n22201, n22200, n22199, n22198,
         n22197, n22196, n22195, n22194, n22193, n22192, n22191, n22190,
         n22189, n22188, n22187, n22186, n22185, n22184, n22183, n22182,
         n22181, n22180, n22179, n22178, n22177, n22176, n22175, n22174,
         n22173, n22172, n22171, n22170, n22169, n22168, n22167, n22166,
         n22165, n22164, n22163, n22162, n22161, n22160, n22159, n22158,
         n22157, n22156, n22155, n22154, n22153, n22152, n22151, n22150,
         n22149, n22148, n22147, n22146, n22145, n22144, n22143, n22142,
         n22141, n22140, n22139, n22138, n22137, n22136, n22135, n22134,
         n22133, n22132, n22131, n22130, n22129, n22128, n22127, n22126,
         n22125, n22124, n22123, n22122, n22121, n22120, n22119, n22118,
         n22117, n22116, n22115, n22114, n22113, n22112, n22111, n22110,
         n22109, n22108, n22107, n22106, n22105, n22104, n22103, n22102,
         n22101, n22100, n22099, n22098, n22097, n22096, n22095, n22094,
         n22093, n22092, n22091, n22090, n22089, n22088, n22087, n22086,
         n22085, n22084, n22083, n22082, n22081, n22080, n22079, n22078,
         n22077, n22076, n22075, n22074, n22073, n22072, n22071, n22070,
         n22069, n22068, n22067, n22066, n22065, n22064, n22063, n22062,
         n22061, n22060, n22059, n22058, n22057, n22056, n22055, n22054,
         n22053, n22052, n22051, n22050, n22049, n22048, n22047, n22046,
         n22045, n22044, n22043, n22042, n22041, n22040, n22039, n22038,
         n22037, n22036, n22035, n22034, n22033, n22032, n22031, n22030,
         n22029, n22028, n22027, n22026, n22025, n22024, n22023, n22022,
         n22021, n22020, n22019, n22018, n22017, n22016, n22015, n22014,
         n22013, n22012, n22011, n22010, n22009, n22008, n22007, n22006,
         n22005, n22004, n22003, n22002, n22001, n22000, n21999, n21998,
         n21997, n21996, n21995, n21994, n21993, n21992, n21991, n21990,
         n21989, n21988, n21987, n21986, n21985, n21984, n21983, n21982,
         n21981, n21980, n21979, n21978, n21977, n21976, n21975, n21974,
         n21973, n21972, n21971, n21970, n21969, n21968, n21967, n21966,
         n21965, n21964, n21963, n21962, n21961, n21960, n21959, n21958,
         n21957, n21956, n21955, n21954, n21953, n21952, n21951, n21950,
         n21949, n21948, n21947, n21946, n21945, n21944, n21943, n21942,
         n21941, n21940, n21939, n21938, n21937, n21936, n21935, n21934,
         n21933, n21932, n21931, n21930, n21929, n21928, n21927, n21926,
         n21925, n21924, n21923, n21922, n21921, n21920, n21919, n21918,
         n21917, n21916, n21915, n21914, n21913, n21912, n21911, n21910,
         n21909, n21908, n21907, n21906, n21905, n21904, n21903, n21902,
         n21901, n21900, n21899, n21898, n21897, n21896, n21895, n21894,
         n21893, n21892, n21891, n21890, n21889, n21888, n21887, n21886,
         n21885, n21884, n21883, n21882, n21881, n21880, n21879, n21878,
         n21877, n21876, n21875, n21874, n21873, n21872, n21871, n21870,
         n21869, n21868, n21867, n21866, n21865, n21864, n21863, n21862,
         n21861, n21860, n21859, n21858, n21857, n21856, n21855, n21854,
         n21853, n21852, n21851, n21850, n21849, n21848, n21847, n21846,
         n21845, n21844, n21843, n21842, n21841, n21840, n21839, n21838,
         n21837, n21836, n21835, n21834, n21833, n21832, n21831, n21830,
         n21829, n21828, n21827, n21826, n21825, n21824, n21823, n21822,
         n21821, n21820, n21819, n21818, n21817, n21816, n21815, n21814,
         n21813, n21812, n21811, n21810, n21809, n21808, n21807, n21806,
         n21805, n21804, n21803, n21802, n21801, n21800, n21799, n21798,
         n21797, n21796, n21795, n21794, n21793, n21792, n21791, n21790,
         n21789, n21788, n21787, n21786, n21785, n21784, n21783, n21782,
         n21781, n21780, n21779, n21778, n21777, n21776, n21775, n21774,
         n21773, n21772, n21771, n21770, n21769, n21768, n21767, n21766,
         n21765, n21764, n21763, n21762, n21761, n21760, n21759, n21758,
         n21757, n21756, n21755, n21754, n21753, n21752, n21751, n21750,
         n21749, n21748, n21747, n21746, n21745, n21744, n21743, n21742,
         n21741, n21740, n21739, n21738, n21737, n21736, n21735, n21734,
         n21733, n21732, n21731, n21730, n21729, n21728, n21727, n21726,
         n21725, n21724, n21723, n21722, n21721, n21720, n21719, n21718,
         n21717, n21716, n21715, n21714, n21713, n21712, n21711, n21710,
         n21709, n21708, n21707, n21706, n21705, n21704, n21703, n21702,
         n21701, n21700, n21699, n21698, n21697, n21696, n21695, n21694,
         n21693, n21692, n21691, n21690, n21689, n21688, n21687, n21686,
         n21685, n21684, n21683, n21682, n21681, n21680, n21679, n21678,
         n21677, n21676, n21675, n21674, n21673, n21672, n21671, n21670,
         n21669, n21668, n21667, n21666, n21665, n21664, n21663, n21662,
         n21661, n21660, n21659, n21658, n21657, n21656, n21655, n21654,
         n21653, n21652, n21651, n21650, n21649, n21648, n21647, n21646,
         n21645, n21644, n21643, n21642, n21641, n21640, n21639, n21638,
         n21637, n21636, n21635, n21634, n21633, n21632, n21631, n21630,
         n21629, n21628, n21627, n21626, n21625, n21624, n21623, n21622,
         n21621, n21620, n21619, n21618, n21617, n21616, n21615, n21614,
         n21613, n21612, n21611, n21610, n21609, n21608, n21607, n21606,
         n21605, n21604, n21603, n21602, n21601, n21600, n21599, n21598,
         n21597, n21596, n21595, n21594, n21593, n21592, n21591, n21590,
         n21589, n21588, n21587, n21586, n21585, n21584, n21583, n21582,
         n21581, n21580, n21579, n21578, n21577, n21576, n21575, n21574,
         n21573, n21572, n21571, n21570, n21569, n21568, n21567, n21566,
         n21565, n21564, n21563, n21562, n21561, n21560, n21559, n21558,
         n21557, n21556, n21555, n21554, n21553, n21552, n21551, n21550,
         n21549, n21548, n21547, n21546, n21545, n21544, n21543, n21542,
         n21541, n21540, n21539, n21538, n21537, n21536, n21535, n21534,
         n21533, n21532, n21531, n21530, n21529, n21528, n21527, n21526,
         n21525, n21524, n21523, n21522, n21521, n21520, n21519, n21518,
         n21517, n21516, n21515, n21514, n21513, n21512, n21511, n21510,
         n21509, n21508, n21507, n21506, n21505, n21504, n21503, n21502,
         n21501, n21500, n21499, n21498, n21497, n21496, n21495, n21494,
         n21493, n21492, n21491, n21490, n21489, n21488, n21487, n21486,
         n21485, n21484, n21483, n21482, n21481, n21480, n21479, n21478,
         n21477, n21476, n21475, n21474, n21473, n21472, n21471, n21470,
         n21469, n21468, n21467, n21466, n21465, n21464, n21463, n21462,
         n21461, n21460, n21459, n21458, n21457, n21456, n21455, n21454,
         n21453, n21452, n21451, n21450, n21449, n21448, n21447, n21446,
         n21445, n21444, n21443, n21442, n21441, n21440, n21439, n21438,
         n21437, n21436, n21435, n21434, n21433, n21432, n21431, n21430,
         n21429, n21428, n21427, n21426, n21425, n21424, n21423, n21422,
         n21421, n21420, n21419, n21418, n21417, n21416, n21415, n21414,
         n21413, n21412, n21411, n21410, n21409, n21408, n21407, n21406,
         n21405, n21404, n21403, n21402, n21401, n21400, n21399, n21398,
         n21397, n21396, n21395, n21394, n21393, n21392, n21391, n21390,
         n21389, n21388, n21387, n21386, n21385, n21384, n21383, n21382,
         n21381, n21380, n21379, n21378, n21377, n21376, n21375, n21374,
         n21373, n21372, n21371, n21370, n21369, n21368, n21367, n21366,
         n21365, n21364, n21363, n21362, n21361, n21360, n21359, n21358,
         n21357, n21356, n21355, n21354, n21353, n21352, n21351, n21350,
         n21349, n21348, n21347, n21346, n21345, n21344, n21343, n21342,
         n21341, n21340, n21339, n21338, n21337, n21336, n21335, n21334,
         n21333, n21332, n21331, n21330, n21329, n21328, n21327, n21326,
         n21325, n21324, n21323, n21322, n21321, n21320, n21319, n21318,
         n21317, n21316, n21315, n21314, n21313, n21312, n21311, n21310,
         n21309, n21308, n21307, n21306, n21305, n21304, n21303, n21302,
         n21301, n21300, n21299, n21298, n21297, n21296, n21295, n21294,
         n21293, n21292, n21291, n21290, n21289, n21288, n21287, n21286,
         n21285, n21284, n21283, n21282, n21281, n21280, n21279, n21278,
         n21277, n21276, n21275, n21274, n21273, n21272, n21271, n21270,
         n21269, n21268, n21267, n21266, n21265, n21264, n21263, n21262,
         n21261, n21260, n21259, n21258, n21257, n21256, n21255, n21254,
         n21253, n21252, n21251, n21250, n21249, n21248, n21247, n21246,
         n21245, n21244, n21243, n21242, n21241, n21240, n21239, n21238,
         n21237, n21236, n21235, n21234, n21233, n21232, n21231, n21230,
         n21229, n21228, n21227, n21226, n21225, n21224, n21223, n21222,
         n21221, n21220, n21219, n21218, n21217, n21216, n21215, n21214,
         n21213, n21212, n21211, n21210, n21209, n21208, n21207, n21206,
         n21205, n21204, n21203, n21202, n21201, n21200, n21199, n21198,
         n21197, n21196, n21195, n21194, n21193, n21192, n21191, n21190,
         n21189, n21188, n21187, n21186, n21185, n21184, n21183, n21182,
         n21181, n21180, n21179, n21178, n21177, n21176, n21175, n21174,
         n21173, n21172, n21171, n21170, n21169, n21168, n21167, n21166,
         n21165, n21164, n21163, n21162, n21161, n21160, n21159, n21158,
         n21157, n21156, n21155, n21154, n21153, n21152, n21151, n21150,
         n21149, n21148, n21147, n21146, n21145, n21144, n21143, n21142,
         n21141, n21140, n21139, n21138, n21137, n21136, n21135, n21134,
         n21133, n21132, n21131, n21130, n21129, n21128, n21127, n21126,
         n21125, n21124, n21123, n21122, n21121, n21120, n21119, n21118,
         n21117, n21116, n21115, n21114, n21113, n21112, n21111, n21110,
         n21109, n21108, n21107, n21106, n21105, n21104, n21103, n21102,
         n21101, n21100, n21099, n21098, n21097, n21096, n21095, n21094,
         n21093, n21092, n21091, n21090, n21089, n21088, n21087, n21086,
         n21085, n21084, n21083, n21082, n21081, n21080, n21079, n21078,
         n21077, n21076, n21075, n21074, n21073, n21072, n21071, n21070,
         n21069, n21068, n21067, n21066, n21065, n21064, n21063, n21062,
         n21061, n21060, n21059, n21058, n21057, n21056, n21055, n21054,
         n21053, n21052, n21051, n21050, n21049, n21048, n21047, n21046,
         n21045, n21044, n21043, n21042, n21041, n21040, n21039, n21038,
         n21037, n21036, n21035, n21034, n21033, n21032, n21031, n21030,
         n21029, n21028, n21027, n21026, n21025, n21024, n21023, n21022,
         n21021, n21020, n21019, n21018, n21017, n21016, n21015, n21014,
         n21013, n21012, n21011, n21010, n21009, n21008, n21007, n21006,
         n21005, n21004, n21003, n21002, n21001, n21000, n20999, n20998,
         n20997, n20996, n20995, n20994, n20993, n20992, n20991, n20990,
         n20989, n20988, n20987, n20986, n20985, n20984, n20983, n20982,
         n20981, n20980, n20979, n20978, n20977, n20976, n20975, n20974,
         n20973, n20972, n20971, n20970, n20969, n20968, n20967, n20966,
         n20965, n20964, n20963, n20962, n20961, n20960, n20959, n20958,
         n20957, n20956, n20955, n20954, n20953, n20952, n20951, n20950,
         n20949, n20948, n20947, n20946, n20945, n20944, n20943, n20942,
         n20941, n20940, n20939, n20938, n20937, n20936, n20935, n20934,
         n20933, n20932, n20931, n20930, n20929, n20928, n20927, n20926,
         n20925, n20924, n20923, n20922, n20921, n20920, n20919, n20918,
         n20917, n20916, n20915, n20914, n20913, n20912, n20911, n20910,
         n20909, n20908, n20907, n20906, n20905, n20904, n20903, n20902,
         n20901, n20900, n20899, n20898, n20897, n20896, n20895, n20894,
         n20893, n20892, n20891, n20890, n20889, n20888, n20887, n20886,
         n20885, n20884, n20883, n20882, n20881, n20880, n20879, n20878,
         n20877, n20876, n20875, n20874, n20873, n20872, n20871, n20870,
         n20869, n20868, n20867, n20866, n20865, n20864, n20863, n20862,
         n20861, n20860, n20859, n20858, n20857, n20856, n20855, n20854,
         n20853, n20852, n20851, n20850, n20849, n20848, n20847, n20846,
         n20845, n20844, n20843, n20842, n20841, n20840, n20839, n20838,
         n20837, n20836, n20835, n20834, n20833, n20832, n20831, n20830,
         n20829, n20828, n20827, n20826, n20825, n20824, n20823, n20822,
         n20821, n20820, n20819, n20818, n20817, n20816, n20815, n20814,
         n20813, n20812, n20811, n20810, n20809, n20808, n20807, n20806,
         n20805, n20804, n20803, n20802, n20801, n20800, n20799, n20798,
         n20797, n20796, n20795, n20794, n20793, n20792, n20791, n20790,
         n20789, n20788, n20787, n20786, n20785, n20784, n20783, n20782,
         n20781, n20780, n20779, n20778, n20777, n20776, n20775, n20774,
         n20773, n20772, n20771, n20770, n20769, n20768, n20767, n20766,
         n20765, n20764, n20763, n20762, n20761, n20760, n20759, n20758,
         n20757, n20756, n20755, n20754, n20753, n20752, n20751, n20750,
         n20749, n20748, n20747, n20746, n20745, n20744, n20743, n20742,
         n20741, n20740, n20739, n20738, n20737, n20736, n20735, n20734,
         n20733, n20732, n20731, n20730, n20729, n20728, n20727, n20726,
         n20725, n20724, n20723, n20722, n20721, n20720, n20719, n20718,
         n20717, n20716, n20715, n20714, n20713, n20712, n20711, n20710,
         n20709, n20708, n20707, n20706, n20705, n20704, n20703, n20702,
         n20701, n20700, n20699, n20698, n20697, n20696, n20695, n20694,
         n20693, n20692, n20691, n20690, n20689, n20688, n20687, n20686,
         n20685, n20684, n20683, n20682, n20681, n20680, n20679, n20678,
         n20677, n20676, n20675, n20674, n20673, n20672, n20671, n20670,
         n20669, n20668, n20667, n20666, n20665, n20664, n20663, n20662,
         n20661, n20660, n20659, n20658, n20657, n20656, n20655, n20654,
         n20653, n20652, n20651, n20650, n20649, n20648, n20647, n20646,
         n20645, n20644, n20643, n20642, n20641, n20640, n20639, n20638,
         n20637, n20636, n20635, n20634, n20633, n20632, n20631, n20630,
         n20629, n20628, n20627, n20626, n20625, n20624, n20623, n20622,
         n20621, n20620, n20619, n20618, n20617, n20616, n20615, n20614,
         n20613, n20612, n20611, n20610, n20609, n20608, n20607, n20606,
         n20605, n20604, n20603, n20602, n20601, n20600, n20599, n20598,
         n20597, n20596, n20595, n20594, n20593, n20592, n20591, n20590,
         n20589, n20588, n20587, n20586, n20585, n20584, n20583, n20582,
         n20581, n20580, n20579, n20578, n20577, n20576, n20575, n20574,
         n20573, n20572, n20571, n20570, n20569, n20568, n20567, n20566,
         n20565, n20564, n20563, n20562, n20561, n20560, n20559, n20558,
         n20557, n20556, n20555, n20554, n20553, n20552, n20551, n20550,
         n20549, n20548, n20547, n20546, n20545, n20544, n20543, n20542,
         n20541, n20540, n20539, n20538, n20537, n20536, n20535, n20534,
         n20533, n20532, n20531, n20530, n20529, n20528, n20527, n20526,
         n20525, n20524, n20523, n20522, n20521, n20520, n20519, n20518,
         n20517, n20516, n20515, n20514, n20513, n20512, n20511, n20510,
         n20509, n20508, n20507, n20506, n20505, n20504, n20503, n20502,
         n20501, n20500, n20499, n20498, n20497, n20496, n20495, n20494,
         n20493, n20492, n20491, n20490, n20489, n20488, n20487, n20486,
         n20485, n20484, n20483, n20482, n20481, n20480, n20479, n20478,
         n20477, n20476, n20475, n20474, n20473, n20472, n20471, n20470,
         n20469, n20468, n20467, n20466, n20465, n20464, n20463, n20462,
         n20461, n20460, n20459, n20458, n20457, n20456, n20455, n20454,
         n20453, n20452, n20451, n20450, n20449, n20448, n20447, n20446,
         n20445, n20444, n20443, n20442, n20441, n20440, n20439, n20438,
         n20437, n20436, n20435, n20434, n20433, n20432, n20431, n20430,
         n20429, n20428, n20427, n20426, n20425, n20424, n20423, n20422,
         n20421, n20420, n20419, n20418, n20417, n20416, n20415, n20414,
         n20413, n20412, n20411, n20410, n20409, n20408, n20407, n20406,
         n20405, n20404, n20403, n20402, n20401, n20400, n20399, n20398,
         n20397, n20396, n20395, n20394, n20393, n20392, n20391, n20390,
         n20389, n20388, n20387, n20386, n20385, n20384, n20383, n20382,
         n20381, n20380, n20379, n20378, n20377, n20376, n20375, n20374,
         n20373, n20372, n20371, n20370, n20369, n20368, n20367, n20366,
         n20365, n20364, n20363, n20362, n20361, n20360, n20359, n20358,
         n20357, n20356, n20355, n20354, n20353, n20352, n20351, n20350,
         n20349, n20348, n20347, n20346, n20345, n20344, n20343, n20342,
         n20341, n20340, n20339, n20338, n20337, n20336, n20335, n20334,
         n20333, n20332, n20331, n20330, n20329, n20328, n20327, n20326,
         n20325, n20324, n20323, n20322, n20321, n20320, n20319, n20318,
         n20317, n20316, n20315, n20314, n20313, n20312, n20311, n20310,
         n20309, n20308, n20307, n20306, n20305, n20304, n20303, n20302,
         n20301, n20300, n20299, n20298, n20297, n20296, n20295, n20294,
         n20293, n20292, n20291, n20290, n20289, n20288, n20287, n20286,
         n20285, n20284, n20283, n20282, n20281, n20280, n20279, n20278,
         n20277, n20276, n20275, n20274, n20273, n20272, n20271, n20270,
         n20269, n20268, n20267, n20266, n20265, n20264, n20263, n20262,
         n20261, n20260, n20259, n20258, n20257, n20256, n20255, n20254,
         n20253, n20252, n20251, n20250, n20249, n20248, n20247, n20246,
         n20245, n20244, n20243, n20242, n20241, n20240, n20239, n20238,
         n20237, n20236, n20235, n20234, n20233, n20232, n20231, n20230,
         n20229, n20228, n20227, n20226, n20225, n20224, n20223, n20222,
         n20221, n20220, n20219, n20218, n20217, n20216, n20215, n20214,
         n20213, n20212, n20211, n20210, n20209, n20208, n20207, n20206,
         n20205, n20204, n20203, n20202, n20201, n20200, n20199, n20198,
         n20197, n20196, n20195, n20194, n20193, n20192, n20191, n20190,
         n20189, n20188, n20187, n20186, n20185, n20184, n20183, n20182,
         n20181, n20180, n20179, n20178, n20177, n20176, n20175, n20174,
         n20173, n20172, n20171, n20170, n20169, n20168, n20167, n20166,
         n20165, n20164, n20163, n20162, n20161, n20160, n20159, n20158,
         n20157, n20156, n20155, n20154, n20153, n20152, n20151, n20150,
         n20149, n20148, n20147, n20146, n20145, n20144, n20143, n20142,
         n20141, n20140, n20139, n20138, n20137, n20136, n20135, n20134,
         n20133, n20132, n20131, n20130, n20129, n20128, n20127, n20126,
         n20125, n20124, n20123, n20122, n20121, n20120, n20119, n20118,
         n20117, n20116, n20115, n20114, n20113, n20112, n20111, n20110,
         n20109, n20108, n20107, n20106, n20105, n20104, n20103, n20102,
         n20101, n20100, n20099, n20098, n20097, n20096, n20095, n20094,
         n20093, n20092, n20091, n20090, n20089, n20088, n20087, n20086,
         n20085, n20084, n20083, n20082, n20081, n20080, n20079, n20078,
         n20077, n20076, n20075, n20074, n20073, n20072, n20071, n20070,
         n20069, n20068, n20067, n20066, n20065, n20064, n20063, n20062,
         n20061, n20060, n20059, n20058, n20057, n20056, n20055, n20054,
         n20053, n20052, n20051, n20050, n20049, n20048, n20047, n20046,
         n20045, n20044, n20043, n20042, n20041, n20040, n20039, n20038,
         n20037, n20036, n20035, n20034, n20033, n20032, n20031, n20030,
         n20029, n20028, n20027, n20026, n20025, n20024, n20023, n20022,
         n20021, n20020, n20019, n20018, n20017, n20016, n20015, n20014,
         n20013, n20012, n20011, n20010, n20009, n20008, n20007, n20006,
         n20005, n20004, n20003, n20002, n20001, n20000, n19999, n19998,
         n19997, n19996, n19995, n19994, n19993, n19992, n19991, n19990,
         n19989, n19988, n19987, n19986, n19985, n19984, n19983, n19982,
         n19981, n19980, n19979, n19978, n19977, n19976, n19975, n19974,
         n19973, n19972, n19971, n19970, n19969, n19968, n19967, n19966,
         n19965, n19964, n19963, n19962, n19961, n19960, n19959, n19958,
         n19957, n19956, n19955, n19954, n19953, n19952, n19951, n19950,
         n19949, n19948, n19947, n19946, n19945, n19944, n19943, n19942,
         n19941, n19940, n19939, n19938, n19937, n19936, n19935, n19934,
         n19933, n19932, n19931, n19930, n19929, n19928, n19927, n19926,
         n19925, n19924, n19923, n19922, n19921, n19920, n19919, n19918,
         n19917, n19916, n19915, n19914, n19913, n19912, n19911, n19910,
         n19909, n19908, n19907, n19906, n19905, n19904, n19903, n19902,
         n19901, n19900, n19899, n19898, n19897, n19896, n19895, n19894,
         n19893, n19892, n19891, n19890, n19889, n19888, n19887, n19886,
         n19885, n19884, n19883, n19882, n19881, n19880, n19879, n19878,
         n19877, n19876, n19875, n19874, n19873, n19872, n19871, n19870,
         n19869, n19868, n19867, n19866, n19865, n19864, n19863, n19862,
         n19861, n19860, n19859, n19858, n19857, n19856, n19855, n19854,
         n19853, n19852, n19851, n19850, n19849, n19848, n19847, n19846,
         n19845, n19844, n19843, n19842, n19841, n19840, n19839, n19838,
         n19837, n19836, n19835, n19834, n19833, n19832, n19831, n19830,
         n19829, n19828, n19827, n19826, n19825, n19824, n19823, n19822,
         n19821, n19820, n19819, n19818, n19817, n19816, n19815, n19814,
         n19813, n19812, n19811, n19810, n19809, n19808, n19807, n19806,
         n19805, n19804, n19803, n19802, n19801, n19800, n19799, n19798,
         n19797, n19796, n19795, n19794, n19793, n19792, n19791, n19790,
         n19789, n19788, n19787, n19786, n19785, n19784, n19783, n19782,
         n19781, n19780, n19779, n19778, n19777, n19776, n19775, n19774,
         n19773, n19772, n19771, n19770, n19769, n19768, n19767, n19766,
         n19765, n19764, n19763, n19762, n19761, n19760, n19759, n19758,
         n19757, n19756, n19755, n19754, n19753, n19752, n19751, n19750,
         n19749, n19748, n19747, n19746, n19745, n19744, n19743, n19742,
         n19741, n19740, n19739, n19738, n19737, n19736, n19735, n19734,
         n19733, n19732, n19731, n19730, n19729, n19728, n19727, n19726,
         n19725, n19724, n19723, n19722, n19721, n19720, n19719, n19718,
         n19717, n19716, n19715, n19714, n19713, n19712, n19711, n19710,
         n19709, n19708, n19707, n19706, n19705, n19704, n19703, n19702,
         n19701, n19700, n19699, n19698, n19697, n19696, n19695, n19694,
         n19693, n19692, n19691, n19690, n19689, n19688, n19687, n19686,
         n19685, n19684, n19683, n19682, n19681, n19680, n19679, n19678,
         n19677, n19676, n19675, n19674, n19673, n19672, n19671, n19670,
         n19669, n19668, n19667, n19666, n19665, n19664, n19663, n19662,
         n19661, n19660, n19659, n19658, n19657, n19656, n19655, n19654,
         n19653, n19652, n19651, n19650, n19649, n19648, n19647, n19646,
         n19645, n19644, n19643, n19642, n19641, n19640, n19639, n19638,
         n19637, n19636, n19635, n19634, n19633, n19632, n19631, n19630,
         n19629, n19628, n19627, n19626, n19625, n19624, n19623, n19622,
         n19621, n19620, n19619, n19618, n19617, n19616, n19615, n19614,
         n19613, n19612, n19611, n19610, n19609, n19608, n19607, n19606,
         n19605, n19604, n19603, n19602, n19601, n19600, n19599, n19598,
         n19597, n19596, n19595, n19594, n19593, n19592, n19591, n19590,
         n19589, n19588, n19587, n19586, n19585, n19584, n19583, n19582,
         n19581, n19580, n19579, n19578, n19577, n19576, n19575, n19574,
         n19573, n19572, n19571, n19570, n19569, n19568, n19567, n19566,
         n19565, n19564, n19563, n19562, n19561, n19560, n19559, n19558,
         n19557, n19556, n19555, n19554, n19553, n19552, n19551, n19550,
         n19549, n19548, n19547, n19546, n19545, n19544, n19543, n19542,
         n19541, n19540, n19539, n19538, n19537, n19536, n19535, n19534,
         n19533, n19532, n19531, n19530, n19529, n19528, n19527, n19526,
         n19525, n19524, n19523, n19522, n19521, n19520, n19519, n19518,
         n19517, n19516, n19515, n19514, n19513, n19512, n19511, n19510,
         n19509, n19508, n19507, n19506, n19505, n19504, n19503, n19502,
         n19501, n19500, n19499, n19498, n19497, n19496, n19495, n19494,
         n19493, n19492, n19491, n19490, n19489, n19488, n19486, n19485,
         n19484, n19483, n19482, n19481, n19480, n19479, n19478, n19477,
         n19476, n19475, n19474, n19473, n19472, n19471, n19470, n19469,
         n19468, n19467, n19466, n19465, n19464, n19463, n19462, n19461,
         n19460, n19459, n19458, n19457, n19456, n19455, n19454, n19453,
         n19452, n19451, n19450, n19449, n19448, n19447, n19446, n19445,
         n19444, n19443, n19442, n19441, n19440, n19439, n19438, n19437,
         n19436, n19435, n19434, n19433, n19432, n19431, n19430, n19429,
         n19428, n19427, n19426, n19425, n19424, n19423, n19422, n19421,
         n19420, n19419, n19418, n19417, n19416, n19415, n19414, n19413,
         n19412, n19411, n19410, n19409, n19408, n19407, n19406, n19405,
         n19404, n19403, n19402, n19401, n19400, n19399, n19398, n19397,
         n19396, n19395, n19394, n19393, n19392, n19391, n19390, n19389,
         n19388, n19387, n19386, n19385, n19384, n19383, n19382, n19381,
         n19380, n19379, n19378, n19377, n19376, n19375, n19374, n19373,
         n19372, n19371, n19370, n19369, n19368, n19367, n19366, n19365,
         n19364, n19363, n19362, n19361, n19360, n19359, n19358, n19357,
         n19356, n19355, n19354, n19353, n19352, n19351, n19350, n19349,
         n19348, n19347, n19346, n19345, n19344, n19343, n19342, n19341,
         n19340, n19339, n19338, n19337, n19336, n19335, n19334, n19333,
         n19332, n19331, n19330, n19329, n19328, n19327, n19326, n19325,
         n19324, n19323, n19322, n19321, n19320, n19319, n19318, n19317,
         n19316, n19315, n19314, n19313, n19312, n19311, n19310, n19309,
         n19308, n19307, n19306, n19305, n19304, n19303, n19302, n19301,
         n19300, n19299, n19298, n19297, n19296, n19295, n19294, n19293,
         n19292, n19291, n19290, n19289, n19288, n19287, n19286, n19285,
         n19284, n19283, n19282, n19281, n19280, n19279, n19278, n19277,
         n19276, n19275, n19274, n19273, n19272, n19271, n19270, n19269,
         n19268, n19267, n19266, n19265, n19264, n19263, n19262, n19261,
         n19260, n19259, n19258, n19257, n19256, n19255, n19254, n19253,
         n19252, n19251, n19250, n19249, n19248, n19247, n19246, n19245,
         n19244, n19243, n19242, n19241, n19240, n19239, n19238, n19237,
         n19236, n19235, n19234, n19233, n19232, n19231, n19230, n19229,
         n19228, n19227, n19226, n19225, n19224, n19223, n19222, n19221,
         n19220, n19219, n19218, n19217, n19216, n19215, n19214, n19213,
         n19212, n19211, n19210, n19209, n19208, n19207, n19206, n19205,
         n19204, n19203, n19202, n19201, n19200, n19199, n19198, n19197,
         n19196, n19195, n19194, n19193, n19192, n19191, n19190, n19189,
         n19188, n19187, n19186, n19185, n19184, n19183, n19182, n19181,
         n19180, n19179, n19178, n19177, n19176, n19175, n19174, n19173,
         n19172, n19171, n19170, n19169, n19168, n19167, n19166, n19165,
         n19164, n19163, n19162, n19161, n19160, n19159, n19158, n19157,
         n19156, n19155, n19154, n19153, n19152, n19151, n19150, n19149,
         n19148, n19147, n19146, n19145, n19144, n19143, n19142, n19141,
         n19140, n19139, n19138, n19137, n19136, n19135, n19134, n19133,
         n19132, n19131, n19130, n19129, n19128, n19127, n19126, n19125,
         n19124, n19123, n19122, n19121, n19120, n19119, n19118, n19117,
         n19116, n19115, n19114, n19113, n19112, n19111, n19110, n19109,
         n19108, n19107, n19106, n19105, n19104, n19103, n19102, n19101,
         n19100, n19099, n19098, n19097, n19096, n19095, n19094, n19093,
         n19092, n19091, n19090, n19089, n19088, n19087, n19086, n19085,
         n19084, n19083, n19082, n19081, n19080, n19079, n19078, n19077,
         n19076, n19075, n19074, n19073, n19072, n19071, n19070, n19069,
         n19068, n19067, n19066, n19065, n19064, n19063, n19062, n19061,
         n19060, n19059, n19058, n19057, n19056, n19055, n19054, n19053,
         n19052, n19051, n19050, n19049, n19048, n19047, n19046, n19045,
         n19044, n19043, n19042, n19041, n19040, n19039, n19038, n19037,
         n19036, n19035, n19034, n19033, n19032, n19031, n19030, n19029,
         n19028, n19027, n19026, n19025, n19024, n19023, n19022, n19021,
         n19020, n19019, n19018, n19017, n19016, n19015, n19014, n19013,
         n19012, n19011, n19010, n19009, n19008, n19007, n19006, n19005,
         n19004, n19003, n19002, n19001, n19000, n18999, n18998, n18997,
         n18996, n18995, n18994, n18993, n18992, n18991, n18990, n18989,
         n18988, n18987, n18986, n18985, n18984, n18983, n18982, n18981,
         n18980, n18979, n18978, n18977, n18976, n18975, n18974, n18973,
         n18972, n18971, n18970, n18969, n18968, n18967, n18966, n18965,
         n18964, n18963, n18962, n18961, n18960, n18959, n18958, n18957,
         n18956, n18955, n18954, n18953, n18952, n18951, n18950, n18949,
         n18948, n18947, n18946, n18945, n18944, n18943, n18942, n18941,
         n18940, n18939, n18938, n18937, n18936, n18935, n18934, n18933,
         n18932, n18931, n18930, n18929, n18928, n18927, n18926, n18925,
         n18924, n18923, n18922, n18921, n18920, n18919, n18918, n18917,
         n18916, n18915, n18914, n18913, n18911, n18910, n18909, n18908,
         n18907, n18906, n18905, n18904, n18903, n18902, n18901, n18900,
         n18899, n18898, n18897, n18896, n18895, n18894, n18893, n18892,
         n18891, n18890, n18889, n18888, n18887, n18886, n18885, n18884,
         n18883, n18882, n18881, n18880, n18879, n18878, n18877, n18876,
         n18875, n18874, n18873, n18872, n18871, n18870, n18869, n18868,
         n18867, n18866, n18865, n18864, n18863, n18862, n18861, n18860,
         n18859, n18858, n18857, n18856, n18855, n18854, n18853, n18852,
         n18851, n18850, n18849, n18848, n18847, n18846, n18845, n18844,
         n18843, n18842, n18841, n18840, n18839, n18838, n18837, n18836,
         n18835, n18834, n18833, n18832, n18831, n18830, n18829, n18828,
         n18827, n18826, n18825, n18824, n18823, n18822, n18821, n18820,
         n18819, n18818, n18817, n18816, n18815, n18813, n18812, n18811,
         n18810, n18809, n18808, n18807, n18806, n18805, n18804, n18803,
         n18802, n18801, n18800, n18799, n18798, n18797, n18796, n18795,
         n18794, n18793, n18792, n18791, n18790, n18789, n18788, n18787,
         n18786, n18785, n18784, n18783, n18782, n18781, n18780, n18779,
         n18778, n18777, n18776, n18775, n18774, n18773, n18772, n18771,
         n18770, n18769, n18768, n18767, n18766, n18765, n18764, n18763,
         n18762, n18761, n18760, n18759, n18758, n18757, n18756, n18755,
         n18754, n18753, n18752, n18751, n18750, n18749, n18748, n18747,
         n18746, n18745, n18744, n18743, n18742, n18741, n18740, n18739,
         n18738, n18737, n18736, n18735, n18734, n18733, n18732, n18731,
         n18730, n18729, n18728, n18727, n18726, n18725, n18724, n18723,
         n18722, n18721, n18720, n18719, n18718, n18717, n18716, n18715,
         n18714, n18713, n18712, n18711, n18710, n18709, n18708, n18707,
         n18706, n18705, n18704, n18703, n18702, n18701, n18700, n18699,
         n18698, n18697, n18696, n18695, n18694, n18693, n18692, n18691,
         n18690, n18689, n18688, n18687, n18686, n18685, n18684, n18683,
         n18682, n18681, n18680, n18679, n18678, n18677, n18676, n18675,
         n18674, n18673, n18672, n18671, n18670, n18669, n18668, n18667,
         n18666, n18665, n18664, n18663, n18662, n18661, n18660, n18659,
         n18658, n18657, n18656, n18655, n18654, n18653, n18652, n18651,
         n18650, n18649, n18648, n18647, n18646, n18645, n18644, n18643,
         n18642, n18641, n18640, n18639, n18638, n18637, n18636, n18635,
         n18634, n18633, n18632, n18631, n18630, n18629, n18628, n18627,
         n18626, n18625, n18624, n18623, n18622, n18620, n18619, n18618,
         n18617, n18616, n18615, n18614, n18613, n18612, n18611, n18610,
         n18609, n18608, n18607, n18606, n18605, n18604, n18603, n18602,
         n18601, n18600, n18599, n18598, n18597, n18596, n18595, n18594,
         n18593, n18592, n18591, n18590, n18589, n18588, n18587, n18586,
         n18585, n18584, n18583, n18582, n18581, n18580, n18579, n18578,
         n18577, n18576, n18575, n18574, n18573, n18572, n18571, n18570,
         n18569, n18568, n18567, n18566, n18565, n18564, n18563, n18562,
         n18561, n18560, n18559, n18558, n18557, n18556, n18555, n18554,
         n18553, n18552, n18551, n18550, n18549, n18548, n18547, n18546,
         n18545, n18544, n18543, n18542, n18541, n18540, n18539, n18538,
         n18537, n18536, n18535, n18534, n18533, n18532, n18531, n18530,
         n18529, n18528, n18527, n18526, n18525, n18524, n18523, n18522,
         n18521, n18520, n18519, n18518, n18517, n18516, n18515, n18514,
         n18513, n18512, n18511, n18510, n18509, n18508, n18507, n18506,
         n18505, n18504, n18502, n18501, n18500, n18499, n18498, n18497,
         n18496, n18495, n18494, n18493, n18492, n18491, n18490, n18489,
         n18488, n18487, n18486, n18485, n18484, n18483, n18482, n18481,
         n18480, n18479, n18478, n18477, n18476, n18475, n18474, n18473,
         n18472, n18471, n18470, n18469, n18468, n18467, n18466, n18465,
         n18464, n18463, n18462, n18461, n18460, n18459, n18458, n18456,
         n18455, n18454, n18453, n18452, n18451, n18450, n18449, n18448,
         n18447, n18446, n18445, n18444, n18443, n18442, n18441, n18440,
         n18439, n18438, n18436, n18435, n18434, n18433, n18432, n18431,
         n18430, n18429, n18428, n18427, n18426, n18425, n18424, n18423,
         n18422, n18421, n18420, n18419, n18418, n18417, n18416, n18415,
         n18414, n18413, n18411, n18410, n18409, n18408, n18407, n18406,
         n18405, n18404, n18403, n18402, n18401, n18400, n18399, n18398,
         n18397, n18396, n18395, n18394, n18393, n18392, n18391, n18390,
         n18389, n18388, n18387, n18386, n18385, n18384, n18383, n18382,
         n18381, n18380, n18379, n18378, n18377, n18376, n18375, n18374,
         n18373, n18372, n18371, n18370, n18369, n18368, n18367, n18366,
         n18365, n18364, n18363, n18362, n18361, n18360, n18359, n18358,
         n18357, n18356, n18355, n18354, n18353, n18352, n18351, n18350,
         n18349, n18348, n18347, n18346, n18345, n18344, n18343, n18342,
         n18341, n18340, n18339, n18338, n18337, n18336, n18335, n18334,
         n18333, n18332, n18331, n18330, n18329, n18328, n18327, n18326,
         n18325, n18324, n18323, n18322, n18321, n18320, n18319, n18318,
         n18317, n18316, n18315, n18314, n18313, n18312, n18311, n18310,
         n18309, n18308, n18307, n18306, n18305, n18304, n18303, n18302,
         n18301, n18300, n18299, n18298, n18297, n18296, n18295, n18294,
         n18293, n18291, n18290, n18289, n18288, n18287, n18286, n18285,
         n18284, n18283, n18282, n18281, n18280, n18279, n18278, n18277,
         n18276, n18275, n18274, n18273, n18272, n18271, n18270, n18269,
         n18268, n18267, n18266, n18265, n18264, n18263, n18262, n18261,
         n18260, n18259, n18258, n18257, n18256, n18255, n18254, n18253,
         n18252, n18251, n18250, n18249, n18248, n18247, n18246, n18245,
         n18244, n18243, n18242, n18241, n18240, n18239, n18238, n18237,
         n18236, n18235, n18234, n18233, n18232, n18231, n18230, n18229,
         n18228, n18227, n18226, n18225, n18224, n18223, n18222, n18221,
         n18220, n18219, n18218, n18217, n18216, n18215, n18214, n18213,
         n18212, n18211, n18210, n18209, n18208, n18207, n18206, n18205,
         n18204, n18203, n18202, n18201, n18200, n18199, n18198, n18197,
         n18196, n18195, n18194, n18193, n18192, n18191, n18190, n18189,
         n18188, n18187, n18186, n18185, n18184, n18183, n18182, n18181,
         n18180, n18179, n18178, n18177, n18176, n18175, n18174, n18173,
         n18172, n18171, n18170, n18169, n18168, n18167, n18166, n18165,
         n18164, n18163, n18162, n18161, n18160, n18159, n18158, n18157,
         n18156, n18155, n18154, n18153, n18152, n18151, n18150, n18149,
         n18148, n18147, n18146, n18145, n18144, n18143, n18142, n18141,
         n18139, n18138, n18137, n18136, n18135, n18134, n18133, n18132,
         n18131, n18130, n18129, n18128, n18127, n18126, n18125, n18124,
         n18123, n18122, n18121, n18120, n18119, n18118, n18117, n18116,
         n18115, n18114, n18113, n18112, n18111, n18110, n18109, n18108,
         n18107, n18106, n18105, n18104, n18103, n18102, n18101, n18100,
         n18099, n18098, n18097, n18096, n18095, n18094, n18093, n18092,
         n18091, n18090, n18089, n18088, n18087, n18086, n18085, n18084,
         n18083, n18082, n18081, n18080, n18079, n18078, n18077, n18076,
         n18075, n18074, n18073, n18072, n18071, n18070, n18069, n18068,
         n18067, n18066, n18065, n18064, n18063, n18062, n18061, n18060,
         n18059, n18058, n18057, n18056, n18055, n18054, n18053, n18052,
         n18051, n18050, n18049, n18048, n18047, n18046, n18045, n18044,
         n18043, n18042, n18041, n18040, n18039, n18038, n18037, n18036,
         n18035, n18034, n18033, n18032, n18031, n18030, n18029, n18028,
         n18027, n18026, n18025, n18024, n18023, n18022, n18021, n18020,
         n18019, n18018, n18017, n18016, n18015, n18014, n18013, n18012,
         n18011, n18010, n18009, n18008, n18007, n18006, n18005, n18004,
         n18003, n18002, n18001, n18000, n17999, n17998, n17997, n17996,
         n17995, n17994, n17992, n17991, n17990, n17989, n17988, n17987,
         n17986, n17985, n17984, n17983, n17982, n17981, n17980, n17979,
         n17978, n17977, n17976, n17975, n17974, n17973, n17972, n17971,
         n17970, n17969, n17968, n17967, n17966, n17965, n17964, n17963,
         n17962, n17961, n17960, n17959, n17958, n17957, n17956, n17955,
         n17954, n17953, n17952, n17951, n17950, n17949, n17948, n17947,
         n17946, n17945, n17944, n17943, n17942, n17941, n17940, n17939,
         n17938, n17937, n17936, n17935, n17934, n17933, n17932, n17931,
         n17930, n17929, n17928, n17927, n17926, n17925, n17924, n17923,
         n17922, n17921, n17920, n17919, n17918, n17917, n17916, n17915,
         n17914, n17913, n17912, n17911, n17910, n17909, n17908, n17907,
         n17906, n17905, n17904, n17903, n17902, n17901, n17900, n17899,
         n17898, n17897, n17896, n17895, n17894, n17893, n17892, n17891,
         n17890, n17889, n17888, n17887, n17886, n17885, n17884, n17883,
         n17882, n17881, n17880, n17879, n17878, n17877, n17876, n17875,
         n17874, n17873, n17872, n17871, n17870, n17869, n17868, n17867,
         n17866, n17865, n17864, n17863, n17862, n17861, n17860, n17859,
         n17858, n17857, n17856, n17855, n17854, n17853, n17852, n17851,
         n17850, n17849, n17848, n17847, n17846, n17845, n17844, n17843,
         n17842, n17841, n17840, n17839, n17838, n17837, n17836, n17835,
         n17834, n17833, n17832, n17831, n17830, n17829, n17828, n17827,
         n17826, n17825, n17824, n17823, n17822, n17821, n17820, n17819,
         n17818, n17817, n17816, n17815, n17814, n17813, n17812, n17811,
         n17810, n17809, n17808, n17807, n17806, n17805, n17804, n17803,
         n17802, n17801, n17800, n17799, n17798, n17797, n17796, n17795,
         n17794, n17793, n17792, n17791, n17790, n17789, n17788, n17787,
         n17786, n17785, n17784, n17783, n17782, n17781, n17780, n17779,
         n17778, n17777, n17776, n17775, n17774, n17773, n17772, n17771,
         n17770, n17769, n17768, n17767, n17766, n17765, n17764, n17763,
         n17762, n17761, n17760, n17759, n17758, n17757, n17756, n17755,
         n17754, n17753, n17752, n17751, n17750, n17749, n17748, n17747,
         n17746, n17745, n17744, n17743, n17742, n17741, n17740, n17739,
         n17738, n17737, n17736, n17735, n17734, n17733, n17732, n17731,
         n17730, n17729, n17728, n17727, n17726, n17725, n17724, n17723,
         n17722, n17721, n17720, n17719, n17718, n17717, n17716, n17715,
         n17714, n17713, n17712, n17711, n17710, n17709, n17708, n17707,
         n17706, n17705, n17704, n17703, n17702, n17701, n17700, n17699,
         n17698, n17697, n17696, n17695, n17694, n17693, n17692, n17691,
         n17690, n17689, n17688, n17687, n17686, n17685, n17684, n17683,
         n17681, n17680, n17679, n17678, n17677, n17676, n17675, n17674,
         n17673, n17672, n17671, n17670, n17669, n17668, n17667, n17666,
         n17665, n17664, n17663, n17662, n17661, n17660, n17659, n17658,
         n17657, n17656, n17655, n17654, n17653, n17652, n17651, n17650,
         n17649, n17648, n17647, n17646, n17645, n17644, n17643, n17642,
         n17641, n17640, n17639, n17638, n17637, n17636, n17635, n17634,
         n17633, n17632, n17631, n17630, n17629, n17628, n17627, n17626,
         n17625, n17624, n17623, n17622, n17621, n17620, n17619, n17618,
         n17617, n17615, n17614, n17613, n17612, n17611, n17610, n17609,
         n17608, n17607, n17606, n17605, n17604, n17603, n17602, n17601,
         n17600, n17599, n17598, n17597, n17596, n17595, n17594, n17593,
         n17592, n17590, n17589, n17588, n17587, n17586, n17585, n17584,
         n17583, n17582, n17581, n17580, n17579, n17578, n17577, n17576,
         n17575, n17574, n17573, n17572, n17571, n17570, n17569, n17568,
         n17567, n17566, n17565, n17564, n17563, n17562, n17561, n17560,
         n17559, n17558, n17557, n17556, n17555, n17554, n17553, n17552,
         n17551, n17550, n17549, n17548, n17547, n17546, n17545, n17544,
         n17543, n17542, n17541, n17540, n17539, n17538, n17537, n17536,
         n17535, n17534, n17533, n17532, n17531, n17530, n17529, n17528,
         n17527, n17526, n17525, n17524, n17523, n17522, n17521, n17520,
         n17519, n17518, n17517, n17516, n17515, n17514, n17513, n17512,
         n17511, n17510, n17509, n17508, n17507, n17506, n17505, n17504,
         n17503, n17502, n17501, n17500, n17499, n17498, n17497, n17496,
         n17495, n17494, n17493, n17492, n17491, n17490, n17489, n17488,
         n17487, n17486, n17485, n17484, n17483, n17482, n17481, n17480,
         n17479, n17478, n17477, n17476, n17475, n17474, n17472, n17471,
         n17470, n17468, n17467, n17466, n17465, n17464, n17462, n17461,
         n17460, n17459, n17458, n17457, n17456, n17455, n17454, n17453,
         n17452, n17451, n17450, n17449, n17448, n17447, n17446, n17445,
         n17444, n17443, n17442, n17441, n17440, n17439, n17438, n17437,
         n17436, n17435, n17434, n17433, n17432, n17431, n17430, n17429,
         n17428, n17427, n17426, n17425, n17424, n17423, n17422, n17421,
         n17420, n17419, n17418, n17417, n17416, n17415, n17414, n17413,
         n17412, n17411, n17410, n17409, n17408, n17407, n17406, n17405,
         n17404, n17403, n17402, n17401, n17400, n17399, n17398, n17397,
         n17396, n17395, n17394, n17393, n17392, n17391, n17390, n17389,
         n17388, n17387, n17386, n17385, n17384, n17383, n17382, n17381,
         n17380, n17379, n17378, n17377, n17376, n17375, n17374, n17373,
         n17372, n17371, n17370, n17369, n17368, n17367, n17366, n17365,
         n17364, n17363, n17362, n17361, n17360, n17359, n17358, n17357,
         n17356, n17355, n17354, n17353, n17352, n17351, n17350, n17349,
         n17348, n17347, n17346, n17345, n17344, n17343, n17342, n17341,
         n17340, n17339, n17338, n17337, n17336, n17335, n17334, n17333,
         n17332, n17331, n17330, n17329, n17328, n17327, n17326, n17325,
         n17324, n17323, n17322, n17321, n17320, n17319, n17318, n17317,
         n17316, n17315, n17314, n17313, n17312, n17311, n17310, n17309,
         n17308, n17307, n17306, n17305, n17304, n17303, n17302, n17301,
         n17300, n17299, n17298, n17297, n17296, n17295, n17294, n17293,
         n17292, n17291, n17290, n17289, n17288, n17287, n17286, n17285,
         n17284, n17283, n17282, n17281, n17280, n17279, n17278, n17277,
         n17276, n17275, n17274, n17273, n17272, n17271, n17269, n17268,
         n17267, n17266, n17265, n17264, n17263, n17262, n17261, n17260,
         n17259, n17258, n17257, n17256, n17255, n17254, n17253, n17252,
         n17251, n17250, n17249, n17248, n17247, n17246, n17245, n17244,
         n17243, n17242, n17241, n17240, n17239, n17238, n17237, n17236,
         n17235, n17234, n17233, n17232, n17231, n17230, n17229, n17228,
         n17227, n17226, n17225, n17224, n17223, n17222, n17221, n17220,
         n17219, n17218, n17217, n17216, n17215, n17214, n17213, n17212,
         n17211, n17210, n17209, n17208, n17207, n17206, n17205, n17204,
         n17203, n17202, n17201, n17200, n17199, n17198, n17197, n17196,
         n17195, n17194, n17193, n17192, n17191, n17190, n17189, n17188,
         n17187, n17186, n17185, n17184, n17183, n17182, n17181, n17180,
         n17179, n17178, n17177, n17176, n17175, n17174, n17173, n17171,
         n17170, n17169, n17168, n17167, n17166, n17165, n17164, n17163,
         n17162, n17161, n17160, n17159, n17158, n17157, n17156, n17155,
         n17154, n17153, n17152, n17151, n17150, n17149, n17148, n17147,
         n17146, n17145, n17144, n17143, n17142, n17141, n17140, n17139,
         n17138, n17137, n17136, n17135, n17134, n17133, n17132, n17131,
         n17130, n17129, n17128, n17127, n17126, n17125, n17124, n17123,
         n17122, n17121, n17120, n17119, n17118, n17117, n17116, n17115,
         n17114, n17113, n17112, n17111, n17110, n17108, n17107, n17106,
         n17105, n17104, n17103, n17102, n17101, n17100, n17099, n17098,
         n17097, n17096, n17095, n17094, n17093, n17092, n17091, n17090,
         n17089, n17088, n17087, n17085, n17084, n17083, n17082, n17081,
         n17080, n17079, n17078, n17077, n17076, n17075, n17074, n17073,
         n17072, n17071, n17070, n17069, n17068, n17067, n17066, n17065,
         n17064, n17063, n17062, n17061, n17060, n17059, n17058, n17057,
         n17056, n17055, n17054, n17053, n17052, n17051, n17050, n17049,
         n17048, n17047, n17046, n17045, n17044, n17043, n17042, n17041,
         n17040, n17039, n17038, n17037, n17036, n17035, n17034, n17033,
         n17032, n17031, n17030, n17029, n17028, n17027, n17026, n17025,
         n17024, n17023, n17022, n17021, n17020, n17019, n17018, n17017,
         n17016, n17015, n17014, n17013, n17012, n17011, n17010, n17009,
         n17008, n17007, n17006, n17005, n17004, n17003, n17002, n17001,
         n17000, n16999, n16998, n16997, n16996, n16995, n16994, n16993,
         n16992, n16991, n16990, n16989, n16988, n16987, n16986, n16985,
         n16984, n16983, n16982, n16981, n16980, n16979, n16978, n16977,
         n16976, n16975, n16974, n16973, n16972, n16971, n16970, n16969,
         n16968, n16967, n16966, n16965, n16964, n16963, n16962, n16961,
         n16960, n16959, n16958, n16957, n16956, n16955, n16954, n16953,
         n16952, n16951, n16950, n16949, n16948, n16947, n16946, n16945,
         n16944, n16943, n16942, n16941, n16940, n16939, n16938, n16937,
         n16936, n16935, n16934, n16933, n16932, n16931, n16930, n16929,
         n16928, n16927, n16926, n16925, n16924, n16923, n16922, n16921,
         n16920, n16919, n16918, n16917, n16916, n16915, n16914, n16913,
         n16912, n16911, n16910, n16909, n16908, n16907, n16906, n16905,
         n16904, n16903, n16902, n16901, n16900, n16899, n16898, n16897,
         n16896, n16895, n16894, n16893, n16892, n16891, n16890, n16889,
         n16888, n16887, n16886, n16885, n16884, n16883, n16882, n16881,
         n16880, n16879, n16878, n16877, n16876, n16875, n16874, n16873,
         n16872, n16871, n16870, n16869, n16868, n16867, n16866, n16865,
         n16864, n16862, n16861, n16860, n16859, n16858, n16857, n16856,
         n16855, n16854, n16853, n16852, n16851, n16850, n16848, n16847,
         n16846, n16845, n16844, n16843, n16842, n16841, n16840, n16839,
         n16838, n16837, n16836, n16835, n16834, n16833, n16832, n16831,
         n16830, n16829, n16828, n16827, n16826, n16825, n16824, n16823,
         n16822, n16821, n16820, n16819, n16818, n16817, n16816, n16815,
         n16814, n16813, n16812, n16811, n16810, n16809, n16808, n16807,
         n16806, n16805, n16804, n16803, n16802, n16801, n16800, n16799,
         n16798, n16797, n16796, n16794, n16793, n16792, n16791, n16790,
         n16789, n16788, n16787, n16786, n16785, n16784, n16783, n16782,
         n16781, n16780, n16779, n16778, n16777, n16776, n16775, n16774,
         n16773, n16772, n16771, n16769, n16768, n16767, n16766, n16765,
         n16764, n16763, n16762, n16761, n16760, n16759, n16758, n16757,
         n16756, n16755, n16754, n16753, n16752, n16751, n16750, n16749,
         n16748, n16747, n16746, n16745, n16744, n16743, n16742, n16741,
         n16740, n16739, n16738, n16737, n16736, n16735, n16734, n16733,
         n16732, n16731, n16730, n16729, n16728, n16727, n16726, n16725,
         n16724, n16723, n16722, n16721, n16720, n16719, n16718, n16717,
         n16716, n16715, n16714, n16713, n16712, n16711, n16710, n16709,
         n16708, n16707, n16706, n16705, n16704, n16703, n16702, n16701,
         n16700, n16699, n16698, n16697, n16696, n16695, n16694, n16693,
         n16692, n16691, n16690, n16689, n16688, n16687, n16686, n16685,
         n16684, n16683, n16682, n16681, n16680, n16679, n16678, n16677,
         n16676, n16675, n16674, n16673, n16672, n16671, n16670, n16669,
         n16668, n16667, n16666, n16665, n16664, n16663, n16662, n16661,
         n16660, n16659, n16658, n16657, n16656, n16655, n16654, n16653,
         n16652, n16650, n16649, n16648, n16647, n16646, n16645, n16644,
         n16643, n16642, n16641, n16640, n16639, n16638, n16637, n16636,
         n16635, n16634, n16633, n16632, n16631, n16630, n16629, n16628,
         n16627, n16626, n16625, n16624, n16623, n16622, n16621, n16620,
         n16619, n16618, n16617, n16616, n16615, n16614, n16613, n16612,
         n16611, n16610, n16609, n16608, n16607, n16606, n16605, n16604,
         n16603, n16602, n16601, n16600, n16599, n16598, n16597, n16596,
         n16595, n16594, n16593, n16592, n16591, n16590, n16589, n16588,
         n16587, n16586, n16585, n16584, n16583, n16582, n16581, n16580,
         n16579, n16578, n16577, n16576, n16575, n16574, n16573, n16572,
         n16571, n16570, n16569, n16568, n16567, n16566, n16565, n16564,
         n16563, n16562, n16561, n16560, n16559, n16558, n16557, n16556,
         n16555, n16554, n16553, n16552, n16551, n16550, n16549, n16548,
         n16547, n16546, n16545, n16544, n16543, n16542, n16541, n16540,
         n16539, n16538, n16537, n16536, n16535, n16534, n16533, n16532,
         n16531, n16530, n16529, n16528, n16527, n16526, n16525, n16524,
         n16523, n16522, n16521, n16520, n16519, n16518, n16517, n16516,
         n16515, n16514, n16513, n16512, n16511, n16510, n16509, n16508,
         n16507, n16506, n16505, n16504, n16503, n16502, n16501, n16500,
         n16499, n16498, n16497, n16496, n16495, n16494, n16493, n16492,
         n16491, n16490, n16489, n16488, n16487, n16486, n16485, n16484,
         n16483, n16482, n16481, n16480, n16479, n16478, n16477, n16476,
         n16475, n16474, n16473, n16472, n16471, n16470, n16469, n16468,
         n16467, n16466, n16465, n16464, n16463, n16462, n16461, n16460,
         n16459, n16458, n16457, n16456, n16455, n16454, n16452, n16451,
         n16450, n16449, n16448, n16447, n16446, n16445, n16444, n16443,
         n16442, n16441, n16440, n16439, n16438, n16437, n16436, n16435,
         n16434, n16433, n16432, n16431, n16430, n16429, n16428, n16427,
         n16426, n16425, n16424, n16423, n16422, n16421, n16420, n16419,
         n16418, n16417, n16416, n16415, n16414, n16413, n16412, n16411,
         n16410, n16409, n16408, n16407, n16406, n16405, n16404, n16403,
         n16402, n16401, n16400, n16399, n16398, n16397, n16396, n16395,
         n16394, n16393, n16392, n16391, n16390, n16389, n16388, n16387,
         n16386, n16385, n16384, n16383, n16382, n16381, n16380, n16379,
         n16378, n16377, n16376, n16375, n16374, n16373, n16372, n16371,
         n16370, n16369, n16368, n16367, n16366, n16365, n16364, n16363,
         n16362, n16361, n16360, n16359, n16358, n16357, n16356, n16354,
         n16353, n16352, n16351, n16350, n16349, n16348, n16347, n16346,
         n16345, n16344, n16343, n16342, n16341, n16340, n16339, n16338,
         n16337, n16336, n16335, n16334, n16333, n16332, n16331, n16330,
         n16329, n16328, n16327, n16326, n16325, n16324, n16323, n16322,
         n16321, n16320, n16319, n16318, n16317, n16316, n16315, n16314,
         n16313, n16312, n16311, n16310, n16309, n16308, n16307, n16306,
         n16305, n16304, n16303, n16302, n16301, n16300, n16299, n16298,
         n16297, n16296, n16295, n16294, n16293, n16292, n16291, n16290,
         n16289, n16288, n16287, n16286, n16285, n16284, n16283, n16282,
         n16281, n16280, n16279, n16278, n16277, n16276, n16275, n16274,
         n16273, n16272, n16271, n16270, n16269, n16268, n16267, n16266,
         n16265, n16264, n16263, n16262, n16261, n16260, n16259, n16258,
         n16257, n16256, n16255, n16254, n16253, n16252, n16251, n16250,
         n16249, n16248, n16247, n16246, n16245, n16244, n16243, n16242,
         n16241, n16240, n16239, n16238, n16237, n16236, n16235, n16234,
         n16233, n16232, n16231, n16230, n16229, n16228, n16227, n16226,
         n16225, n16224, n16223, n16222, n16221, n16220, n16219, n16218,
         n16217, n16216, n16215, n16214, n16213, n16212, n16211, n16210,
         n16209, n16208, n16207, n16206, n16205, n16204, n16203, n16202,
         n16201, n16200, n16199, n16198, n16197, n16196, n16195, n16194,
         n16193, n16192, n16191, n16190, n16189, n16188, n16187, n16186,
         n16185, n16184, n16183, n16182, n16181, n16180, n16179, n16178,
         n16177, n16176, n16175, n16174, n16173, n16172, n16171, n16170,
         n16169, n16168, n16167, n16166, n16165, n16164, n16163, n16161,
         n16160, n16159, n16158, n16157, n16156, n16155, n16154, n16153,
         n16152, n16151, n16150, n16149, n16148, n16147, n16146, n16145,
         n16144, n16143, n16142, n16141, n16140, n16139, n16138, n16137,
         n16136, n16135, n16134, n16133, n16132, n16131, n16130, n16129,
         n16128, n16127, n16126, n16125, n16124, n16123, n16122, n16121,
         n16120, n16119, n16118, n16117, n16116, n16115, n16114, n16113,
         n16112, n16111, n16110, n16109, n16108, n16107, n16106, n16105,
         n16104, n16103, n16102, n16101, n16100, n16099, n16098, n16097,
         n16096, n16095, n16094, n16093, n16092, n16091, n16090, n16089,
         n16088, n16087, n16086, n16085, n16084, n16083, n16082, n16081,
         n16080, n16079, n16078, n16077, n16076, n16075, n16074, n16073,
         n16072, n16071, n16070, n16069, n16068, n16067, n16066, n16065,
         n16064, n16063, n16062, n16061, n16060, n16059, n16058, n16057,
         n16056, n16055, n16054, n16053, n16052, n16051, n16050, n16049,
         n16048, n16047, n16046, n16045, n16044, n16043, n16042, n16041,
         n16040, n16039, n16038, n16037, n16036, n16035, n16034, n16033,
         n16032, n16031, n16030, n16029, n16028, n16027, n16026, n16025,
         n16024, n16023, n16022, n16021, n16020, n16019, n16018, n16017,
         n16016, n16015, n16014, n16013, n16012, n16011, n16010, n16009,
         n16008, n16007, n16006, n16004, n16003, n16002, n16001, n16000,
         n15999, n15997, n15996, n15995, n15994, n15993, n15992, n15991,
         n15990, n15989, n15988, n15987, n15986, n15985, n15984, n15983,
         n15982, n15981, n15980, n15979, n15977, n15976, n15975, n15974,
         n15973, n15972, n15971, n15970, n15969, n15968, n15967, n15966,
         n15965, n15964, n15963, n15962, n15961, n15960, n15959, n15958,
         n15957, n15956, n15955, n15954, n15952, n15951, n15950, n15949,
         n15948, n15947, n15946, n15945, n15944, n15943, n15942, n15941,
         n15940, n15939, n15938, n15937, n15936, n15935, n15934, n15933,
         n15932, n15931, n15930, n15929, n15928, n15927, n15926, n15925,
         n15924, n15923, n15922, n15921, n15920, n15919, n15918, n15917,
         n15916, n15915, n15914, n15913, n15912, n15911, n15910, n15909,
         n15908, n15907, n15906, n15905, n15904, n15903, n15902, n15901,
         n15900, n15899, n15898, n15897, n15896, n15895, n15894, n15893,
         n15892, n15891, n15890, n15889, n15888, n15887, n15886, n15885,
         n15884, n15883, n15882, n15881, n15880, n15879, n15878, n15877,
         n15876, n15875, n15874, n15873, n15872, n15871, n15870, n15869,
         n15868, n15867, n15866, n15865, n15864, n15863, n15862, n15861,
         n15860, n15859, n15858, n15857, n15856, n15855, n15854, n15853,
         n15852, n15851, n15850, n15849, n15848, n15847, n15846, n15845,
         n15844, n15843, n15842, n15841, n15840, n15839, n15838, n15837,
         n15836, n15835, n15834, n15832, n15831, n15830, n15829, n15828,
         n15827, n15826, n15825, n15824, n15823, n15822, n15821, n15820,
         n15819, n15818, n15817, n15816, n15815, n15814, n15813, n15812,
         n15811, n15810, n15809, n15808, n15807, n15806, n15805, n15804,
         n15803, n15802, n15801, n15800, n15799, n15798, n15797, n15796,
         n15795, n15794, n15793, n15792, n15791, n15790, n15789, n15788,
         n15787, n15786, n15785, n15784, n15783, n15782, n15781, n15780,
         n15779, n15778, n15777, n15776, n15775, n15774, n15773, n15772,
         n15771, n15770, n15769, n15768, n15767, n15766, n15765, n15764,
         n15763, n15762, n15761, n15760, n15759, n15758, n15757, n15756,
         n15755, n15754, n15753, n15752, n15751, n15750, n15749, n15748,
         n15747, n15746, n15745, n15744, n15743, n15742, n15741, n15740,
         n15739, n15738, n15737, n15736, n15735, n15734, n15733, n15732,
         n15731, n15730, n15729, n15728, n15727, n15726, n15725, n15724,
         n15723, n15722, n15721, n15720, n15719, n15718, n15717, n15716,
         n15715, n15714, n15713, n15712, n15711, n15710, n15709, n15708,
         n15707, n15706, n15705, n15704, n15703, n15702, n15701, n15700,
         n15699, n15698, n15697, n15696, n15695, n15694, n15693, n15692,
         n15691, n15690, n15689, n15688, n15687, n15686, n15685, n15684,
         n15683, n15682, n15681, n15680, n15679, n15678, n15677, n15676,
         n15675, n15674, n15673, n15672, n15671, n15670, n15669, n15668,
         n15667, n15666, n15665, n15664, n15663, n15662, n15661, n15660,
         n15659, n15658, n15657, n15656, n15655, n15654, n15653, n15652,
         n15651, n15650, n15649, n15648, n15647, n15646, n15645, n15644,
         n15643, n15642, n15641, n15640, n15639, n15638, n15637, n15636,
         n15635, n15634, n15633, n15632, n15631, n15630, n15629, n15628,
         n15627, n15626, n15625, n15624, n15623, n15622, n15621, n15620,
         n15619, n15618, n15617, n15616, n15615, n15614, n15613, n15612,
         n15611, n15610, n15609, n15608, n15607, n15606, n15605, n15604,
         n15603, n15602, n15601, n15600, n15599, n15598, n15597, n15596,
         n15595, n15594, n15593, n15592, n15591, n15590, n15589, n15588,
         n15587, n15586, n15585, n15584, n15583, n15582, n15581, n15580,
         n15579, n15578, n15577, n15576, n15575, n15574, n15573, n15572,
         n15571, n15570, n15569, n15568, n15567, n15566, n15565, n15564,
         n15563, n15562, n15561, n15560, n15559, n15558, n15557, n15556,
         n15555, n15554, n15553, n15552, n15551, n15550, n15549, n15548,
         n15547, n15546, n15545, n15544, n15543, n15542, n15541, n15540,
         n15539, n15538, n15537, n15535, n15534, n15533, n15532, n15531,
         n15530, n15529, n15528, n15527, n15526, n15525, n15524, n15523,
         n15522, n15521, n15520, n15519, n15518, n15517, n15516, n15515,
         n15514, n15513, n15512, n15511, n15510, n15509, n15508, n15507,
         n15506, n15505, n15504, n15503, n15502, n15501, n15500, n15499,
         n15498, n15497, n15496, n15495, n15494, n15493, n15492, n15491,
         n15490, n15488, n15487, n15486, n15485, n15484, n15483, n15482,
         n15481, n15480, n15479, n15478, n15477, n15476, n15475, n15474,
         n15473, n15472, n15471, n15470, n15469, n15468, n15467, n15466,
         n15465, n15464, n15463, n15462, n15461, n15460, n15459, n15458,
         n15457, n15456, n15455, n15454, n15453, n15452, n15451, n15450,
         n15449, n15448, n15447, n15446, n15445, n15444, n15443, n15442,
         n15441, n15440, n15439, n15438, n15437, n15436, n15435, n15434,
         n15433, n15432, n15431, n15430, n15429, n15428, n15427, n15426,
         n15425, n15424, n15423, n15422, n15421, n15420, n15419, n15418,
         n15417, n15416, n15415, n15414, n15413, n15412, n15411, n15410,
         n15409, n15408, n15407, n15406, n15405, n15404, n15403, n15402,
         n15401, n15400, n15399, n15398, n15397, n15396, n15395, n15394,
         n15393, n15392, n15391, n15390, n15389, n15388, n15387, n15386,
         n15385, n15384, n15383, n15382, n15381, n15380, n15379, n15378,
         n15377, n15376, n15375, n15374, n15373, n15372, n15371, n15370,
         n15369, n15368, n15367, n15366, n15365, n15364, n15363, n15362,
         n15361, n15360, n15359, n15358, n15357, n15356, n15355, n15354,
         n15353, n15352, n15351, n15350, n15349, n15348, n15347, n15346,
         n15345, n15344, n15342, n15341, n15340, n15339, n15338, n15337,
         n15336, n15335, n15334, n15333, n15332, n15331, n15330, n15329,
         n15328, n15327, n15326, n15325, n15324, n15323, n15322, n15321,
         n15320, n15319, n15318, n15317, n15316, n15315, n15314, n15313,
         n15312, n15311, n15310, n15309, n15308, n15307, n15306, n15305,
         n15304, n15303, n15302, n15301, n15300, n15299, n15298, n15297,
         n15296, n15295, n15294, n15293, n15292, n15291, n15290, n15289,
         n15288, n15287, n15286, n15285, n15284, n15283, n15282, n15281,
         n15280, n15279, n15278, n15277, n15276, n15275, n15274, n15273,
         n15271, n15270, n15269, n15268, n15267, n15266, n15265, n15264,
         n15263, n15262, n15261, n15260, n15259, n15258, n15257, n15256,
         n15255, n15254, n15253, n15252, n15251, n15250, n15249, n15248,
         n15247, n15246, n15245, n15244, n15243, n15242, n15241, n15240,
         n15239, n15238, n15237, n15236, n15235, n15234, n15233, n15232,
         n15231, n15230, n15229, n15228, n15227, n15226, n15225, n15224,
         n15223, n15222, n15221, n15220, n15219, n15218, n15217, n15216,
         n15215, n15214, n15213, n15212, n15211, n15210, n15209, n15208,
         n15207, n15206, n15205, n15204, n15203, n15202, n15201, n15200,
         n15199, n15198, n15197, n15196, n15195, n15194, n15193, n15192,
         n15191, n15190, n15189, n15188, n15187, n15185, n15184, n15183,
         n15182, n15181, n15180, n15178, n15177, n15176, n15175, n15174,
         n15173, n15172, n15171, n15170, n15169, n15168, n15167, n15166,
         n15165, n15164, n15163, n15162, n15161, n15160, n15158, n15157,
         n15156, n15155, n15154, n15153, n15152, n15151, n15150, n15149,
         n15148, n15147, n15146, n15145, n15144, n15143, n15142, n15141,
         n15140, n15139, n15138, n15137, n15136, n15135, n15133, n15132,
         n15131, n15130, n15129, n15128, n15127, n15126, n15125, n15124,
         n15123, n15122, n15121, n15120, n15119, n15118, n15117, n15116,
         n15115, n15114, n15113, n15112, n15111, n15110, n15109, n15108,
         n15107, n15106, n15105, n15104, n15103, n15102, n15101, n15100,
         n15099, n15098, n15097, n15096, n15095, n15094, n15093, n15092,
         n15091, n15090, n15089, n15088, n15087, n15086, n15085, n15084,
         n15083, n15082, n15081, n15080, n15079, n15078, n15077, n15076,
         n15075, n15074, n15073, n15072, n15071, n15070, n15069, n15068,
         n15067, n15066, n15065, n15064, n15063, n15062, n15061, n15060,
         n15059, n15058, n15057, n15056, n15055, n15054, n15053, n15052,
         n15051, n15050, n15049, n15048, n15047, n15046, n15045, n15044,
         n15043, n15042, n15041, n15040, n15039, n15038, n15037, n15036,
         n15035, n15034, n15033, n15032, n15031, n15030, n15029, n15028,
         n15027, n15026, n15025, n15024, n15023, n15022, n15021, n15020,
         n15019, n15018, n15017, n15016, n15015, n15013, n15012, n15011,
         n15010, n15009, n15008, n15007, n15006, n15005, n15004, n15003,
         n15002, n15001, n15000, n14999, n14998, n14997, n14996, n14995,
         n14994, n14993, n14992, n14991, n14990, n14989, n14988, n14987,
         n14986, n14985, n14984, n14983, n14982, n14981, n14980, n14979,
         n14978, n14977, n14976, n14975, n14974, n14973, n14972, n14971,
         n14970, n14969, n14968, n14967, n14966, n14965, n14964, n14963,
         n14962, n14961, n14960, n14959, n14958, n14957, n14956, n14955,
         n14954, n14953, n14952, n14951, n14950, n14949, n14948, n14947,
         n14946, n14945, n14944, n14943, n14942, n14941, n14940, n14939,
         n14938, n14937, n14936, n14935, n14934, n14933, n14932, n14931,
         n14930, n14929, n14928, n14927, n14926, n14925, n14924, n14923,
         n14922, n14921, n14920, n14919, n14918, n14917, n14916, n14915,
         n14914, n14913, n14912, n14911, n14910, n14909, n14908, n14907,
         n14906, n14905, n14904, n14903, n14902, n14901, n14900, n14899,
         n14898, n14897, n14896, n14895, n14894, n14893, n14892, n14891,
         n14890, n14889, n14888, n14887, n14886, n14885, n14884, n14883,
         n14882, n14881, n14880, n14879, n14878, n14877, n14876, n14875,
         n14874, n14873, n14872, n14871, n14870, n14869, n14868, n14867,
         n14866, n14865, n14864, n14863, n14862, n14861, n14860, n14859,
         n14858, n14857, n14856, n14855, n14854, n14853, n14852, n14851,
         n14850, n14849, n14848, n14847, n14846, n14845, n14844, n14843,
         n14842, n14841, n14840, n14839, n14838, n14837, n14836, n14835,
         n14834, n14833, n14832, n14831, n14830, n14829, n14828, n14827,
         n14826, n14825, n14824, n14823, n14822, n14821, n14820, n14819,
         n14818, n14817, n14816, n14814, n14813, n14812, n14811, n14810,
         n14809, n14808, n14807, n14806, n14805, n14804, n14803, n14802,
         n14801, n14800, n14799, n14798, n14797, n14796, n14795, n14794,
         n14793, n14792, n14791, n14790, n14789, n14788, n14787, n14786,
         n14785, n14784, n14783, n14782, n14781, n14780, n14779, n14778,
         n14777, n14776, n14775, n14774, n14773, n14772, n14771, n14770,
         n14769, n14768, n14767, n14766, n14765, n14764, n14763, n14762,
         n14761, n14760, n14759, n14758, n14757, n14756, n14755, n14754,
         n14753, n14752, n14751, n14750, n14749, n14748, n14747, n14746,
         n14745, n14744, n14743, n14742, n14741, n14740, n14739, n14738,
         n14737, n14736, n14735, n14734, n14733, n14732, n14731, n14730,
         n14729, n14728, n14727, n14726, n14725, n14724, n14723, n14722,
         n14721, n14720, n14719, n14718, n14716, n14715, n14714, n14713,
         n14712, n14711, n14710, n14709, n14708, n14707, n14706, n14705,
         n14704, n14703, n14702, n14701, n14700, n14699, n14698, n14697,
         n14696, n14695, n14694, n14693, n14692, n14691, n14690, n14689,
         n14688, n14687, n14686, n14685, n14684, n14683, n14682, n14681,
         n14680, n14679, n14678, n14677, n14676, n14675, n14674, n14673,
         n14672, n14671, n14670, n14669, n14668, n14667, n14666, n14665,
         n14664, n14663, n14662, n14661, n14660, n14659, n14658, n14657,
         n14656, n14655, n14654, n14653, n14652, n14651, n14650, n14649,
         n14648, n14647, n14646, n14645, n14644, n14643, n14642, n14641,
         n14640, n14639, n14638, n14637, n14636, n14635, n14634, n14633,
         n14632, n14631, n14630, n14629, n14628, n14627, n14626, n14625,
         n14624, n14623, n14622, n14621, n14620, n14619, n14618, n14617,
         n14616, n14615, n14614, n14613, n14612, n14611, n14610, n14609,
         n14608, n14607, n14606, n14605, n14604, n14603, n14602, n14601,
         n14600, n14599, n14598, n14597, n14596, n14595, n14594, n14593,
         n14592, n14591, n14590, n14589, n14588, n14587, n14586, n14585,
         n14584, n14583, n14582, n14581, n14580, n14579, n14578, n14577,
         n14576, n14575, n14574, n14573, n14572, n14571, n14570, n14569,
         n14568, n14567, n14566, n14565, n14564, n14563, n14562, n14561,
         n14560, n14559, n14558, n14557, n14556, n14555, n14554, n14553,
         n14552, n14551, n14550, n14549, n14548, n14547, n14546, n14545,
         n14544, n14543, n14542, n14541, n14540, n14539, n14538, n14537,
         n14536, n14535, n14534, n14533, n14532, n14531, n14530, n14529,
         n14528, n14527, n14526, n14525, n14523, n14522, n14521, n14520,
         n14519, n14518, n14517, n14516, n14515, n14514, n14513, n14512,
         n14511, n14510, n14509, n14508, n14507, n14506, n14505, n14504,
         n14503, n14502, n14501, n14500, n14499, n14498, n14497, n14496,
         n14495, n14494, n14493, n14492, n14491, n14490, n14489, n14488,
         n14487, n14486, n14485, n14484, n14483, n14482, n14481, n14480,
         n14479, n14478, n14477, n14476, n14475, n14474, n14473, n14472,
         n14471, n14470, n14469, n14468, n14467, n14466, n14465, n14464,
         n14463, n14462, n14461, n14460, n14459, n14458, n14457, n14456,
         n14455, n14454, n14452, n14451, n14450, n14449, n14448, n14447,
         n14446, n14445, n14444, n14443, n14442, n14441, n14440, n14439,
         n14438, n14437, n14436, n14435, n14434, n14433, n14432, n14431,
         n14430, n14429, n14428, n14427, n14426, n14425, n14424, n14423,
         n14422, n14421, n14420, n14419, n14418, n14417, n14416, n14415,
         n14414, n14413, n14412, n14411, n14410, n14409, n14408, n14407,
         n14406, n14405, n14404, n14403, n14402, n14401, n14400, n14399,
         n14398, n14397, n14396, n14395, n14394, n14393, n14392, n14391,
         n14390, n14389, n14388, n14387, n14386, n14385, n14384, n14383,
         n14382, n14381, n14380, n14379, n14378, n14377, n14376, n14375,
         n14374, n14373, n14372, n14371, n14370, n14369, n14368, n14366,
         n14365, n14364, n14363, n14362, n14361, n14359, n14358, n14357,
         n14356, n14355, n14354, n14353, n14352, n14351, n14350, n14349,
         n14348, n14347, n14346, n14345, n14344, n14343, n14342, n14341,
         n14339, n14338, n14337, n14336, n14335, n14334, n14333, n14332,
         n14331, n14330, n14329, n14328, n14327, n14326, n14325, n14324,
         n14323, n14322, n14321, n14320, n14319, n14318, n14317, n14316,
         n14314, n14313, n14312, n14311, n14310, n14309, n14308, n14307,
         n14306, n14305, n14304, n14303, n14302, n14301, n14300, n14299,
         n14298, n14297, n14296, n14295, n14294, n14293, n14292, n14291,
         n14290, n14289, n14288, n14287, n14286, n14285, n14284, n14283,
         n14282, n14281, n14280, n14279, n14278, n14277, n14276, n14275,
         n14274, n14273, n14272, n14271, n14270, n14269, n14268, n14267,
         n14266, n14265, n14264, n14263, n14262, n14261, n14260, n14259,
         n14258, n14257, n14256, n14255, n14254, n14253, n14252, n14251,
         n14250, n14249, n14248, n14247, n14246, n14245, n14244, n14243,
         n14242, n14241, n14240, n14239, n14238, n14237, n14236, n14235,
         n14234, n14233, n14232, n14231, n14230, n14229, n14228, n14227,
         n14226, n14225, n14224, n14223, n14222, n14221, n14220, n14219,
         n14218, n14217, n14216, n14215, n14214, n14213, n14212, n14211,
         n14210, n14209, n14208, n14207, n14206, n14205, n14204, n14203,
         n14202, n14201, n14200, n14199, n14198, n14197, n14196, n14194,
         n14193, n14192, n14191, n14190, n14189, n14188, n14187, n14186,
         n14185, n14184, n14183, n14182, n14181, n14180, n14179, n14178,
         n14177, n14176, n14175, n14174, n14173, n14172, n14171, n14170,
         n14169, n14168, n14167, n14166, n14165, n14164, n14163, n14162,
         n14161, n14160, n14159, n14158, n14157, n14156, n14155, n14154,
         n14153, n14152, n14151, n14150, n14149, n14148, n14147, n14146,
         n14145, n14144, n14143, n14142, n14141, n14140, n14139, n14138,
         n14137, n14136, n14135, n14134, n14133, n14132, n14131, n14130,
         n14129, n14128, n14127, n14126, n14125, n14124, n14123, n14122,
         n14121, n14120, n14119, n14118, n14117, n14116, n14115, n14114,
         n14113, n14112, n14111, n14110, n14109, n14108, n14107, n14106,
         n14105, n14104, n14103, n14102, n14101, n14100, n14099, n14098,
         n14097, n14096, n14095, n14094, n14093, n14092, n14091, n14090,
         n14089, n14088, n14087, n14086, n14085, n14084, n14083, n14082,
         n14081, n14080, n14079, n14078, n14077, n14076, n14075, n14074,
         n14073, n14072, n14071, n14070, n14069, n14068, n14067, n14066,
         n14065, n14064, n14063, n14062, n14061, n14060, n14059, n14058,
         n14057, n14056, n14055, n14054, n14053, n14052, n14051, n14050,
         n14049, n14048, n14047, n14046, n14045, n14044, n14043, n14042,
         n14041, n14040, n14039, n14038, n14037, n14036, n14035, n14034,
         n14033, n14032, n14031, n14030, n14029, n14028, n14027, n14026,
         n14025, n14024, n14023, n14022, n14021, n14020, n14019, n14018,
         n14017, n14016, n14015, n14014, n14013, n14012, n14011, n14010,
         n14009, n14008, n14007, n14006, n14005, n14004, n14003, n14002,
         n14001, n14000, n13999, n13998, n13997, n13996, n13995, n13994,
         n13993, n13992, n13991, n13990, n13989, n13988, n13987, n13986,
         n13985, n13984, n13983, n13982, n13981, n13980, n13979, n13978,
         n13977, n13976, n13975, n13974, n13973, n13972, n13971, n13970,
         n13969, n13968, n13967, n13966, n13965, n13964, n13963, n13962,
         n13961, n13960, n13959, n13958, n13957, n13956, n13955, n13954,
         n13953, n13952, n13951, n13950, n13949, n13948, n13947, n13946,
         n13945, n13944, n13943, n13942, n13941, n13940, n13939, n13938,
         n13937, n13936, n13935, n13934, n13933, n13932, n13931, n13930,
         n13929, n13928, n13927, n13926, n13925, n13924, n13923, n13922,
         n13921, n13920, n13919, n13918, n13917, n13916, n13915, n13914,
         n13913, n13912, n13911, n13910, n13909, n13908, n13907, n13906,
         n13905, n13904, n13903, n13902, n13901, n13900, n13899, n13897,
         n13896, n13895, n13894, n13893, n13892, n13891, n13890, n13889,
         n13888, n13887, n13886, n13885, n13884, n13883, n13882, n13881,
         n13880, n13879, n13878, n13877, n13876, n13875, n13874, n13873,
         n13872, n13871, n13870, n13869, n13868, n13867, n13866, n13865,
         n13864, n13863, n13862, n13861, n13860, n13859, n13858, n13857,
         n13856, n13855, n13854, n13853, n13852, n13851, n13850, n13849,
         n13848, n13847, n13846, n13845, n13844, n13843, n13842, n13841,
         n13840, n13839, n13838, n13837, n13836, n13835, n13834, n13833,
         n13832, n13831, n13830, n13829, n13828, n13827, n13826, n13825,
         n13824, n13823, n13822, n13821, n13820, n13819, n13818, n13817,
         n13816, n13815, n13814, n13813, n13812, n13811, n13810, n13809,
         n13808, n13807, n13806, n13805, n13804, n13803, n13802, n13801,
         n13800, n13799, n13798, n13797, n13796, n13795, n13794, n13793,
         n13792, n13791, n13790, n13789, n13788, n13787, n13786, n13785,
         n13784, n13783, n13782, n13781, n13780, n13779, n13778, n13777,
         n13776, n13775, n13774, n13773, n13772, n13771, n13770, n13769,
         n13768, n13767, n13766, n13765, n13764, n13763, n13762, n13761,
         n13760, n13759, n13758, n13757, n13756, n13755, n13754, n13753,
         n13752, n13751, n13750, n13749, n13748, n13747, n13746, n13745,
         n13744, n13743, n13742, n13741, n13740, n13739, n13738, n13737,
         n13736, n13735, n13734, n13733, n13732, n13731, n13730, n13729,
         n13728, n13727, n13726, n13725, n13724, n13723, n13722, n13721,
         n13720, n13719, n13718, n13717, n13716, n13715, n13714, n13713,
         n13712, n13711, n13710, n13709, n13708, n13707, n13706, n13704,
         n13703, n13702, n13701, n13700, n13699, n13698, n13697, n13696,
         n13695, n13694, n13693, n13692, n13691, n13690, n13689, n13688,
         n13687, n13686, n13685, n13684, n13683, n13682, n13681, n13680,
         n13679, n13678, n13677, n13676, n13675, n13674, n13673, n13672,
         n13671, n13670, n13669, n13668, n13667, n13666, n13665, n13664,
         n13663, n13662, n13661, n13660, n13659, n13658, n13657, n13656,
         n13655, n13654, n13653, n13652, n13651, n13650, n13649, n13648,
         n13647, n13646, n13645, n13644, n13643, n13642, n13641, n13640,
         n13639, n13638, n13637, n13636, n13635, n13634, n13633, n13632,
         n13631, n13630, n13629, n13628, n13627, n13626, n13625, n13624,
         n13623, n13622, n13621, n13620, n13619, n13618, n13617, n13616,
         n13615, n13614, n13613, n13612, n13611, n13610, n13609, n13608,
         n13607, n13606, n13605, n13604, n13603, n13602, n13601, n13600,
         n13599, n13598, n13597, n13596, n13595, n13594, n13593, n13592,
         n13591, n13590, n13589, n13588, n13587, n13586, n13585, n13584,
         n13583, n13582, n13581, n13580, n13579, n13578, n13577, n13576,
         n13575, n13574, n13573, n13572, n13571, n13570, n13569, n13568,
         n13567, n13566, n13565, n13564, n13563, n13562, n13561, n13560,
         n13559, n13558, n13557, n13556, n13555, n13554, n13553, n13552,
         n13551, n13550, n13549, n13548, n13547, n13546, n13545, n13544,
         n13543, n13542, n13540, n13539, n13538, n13537, n13536, n13535,
         n13534, n13533, n13532, n13531, n13530, n13529, n13528, n13527,
         n13526, n13525, n13524, n13523, n13522, n13520, n13519, n13518,
         n13517, n13516, n13515, n13514, n13513, n13512, n13511, n13510,
         n13509, n13508, n13507, n13506, n13505, n13504, n13503, n13502,
         n13501, n13500, n13499, n13498, n13497, n13495, n13494, n13493,
         n13492, n13491, n13490, n13489, n13488, n13487, n13486, n13485,
         n13484, n13483, n13482, n13481, n13480, n13479, n13478, n13477,
         n13476, n13475, n13474, n13473, n13472, n13471, n13470, n13469,
         n13468, n13467, n13466, n13465, n13464, n13463, n13462, n13461,
         n13460, n13459, n13458, n13457, n13456, n13455, n13454, n13453,
         n13452, n13451, n13450, n13449, n13448, n13447, n13446, n13445,
         n13444, n13443, n13442, n13441, n13440, n13439, n13438, n13437,
         n13436, n13435, n13434, n13433, n13432, n13431, n13430, n13429,
         n13428, n13427, n13426, n13425, n13424, n13423, n13422, n13421,
         n13420, n13419, n13418, n13417, n13416, n13415, n13414, n13413,
         n13412, n13411, n13410, n13409, n13408, n13407, n13406, n13405,
         n13404, n13403, n13402, n13401, n13400, n13399, n13398, n13397,
         n13396, n13395, n13394, n13393, n13392, n13391, n13390, n13389,
         n13388, n13387, n13386, n13385, n13384, n13383, n13382, n13381,
         n13380, n13379, n13378, n13377, n13375, n13374, n13373, n13372,
         n13371, n13370, n13369, n13368, n13367, n13366, n13365, n13364,
         n13363, n13362, n13361, n13360, n13359, n13358, n13357, n13356,
         n13355, n13354, n13353, n13352, n13351, n13350, n13349, n13348,
         n13347, n13346, n13345, n13344, n13343, n13342, n13341, n13340,
         n13339, n13338, n13337, n13336, n13335, n13334, n13333, n13332,
         n13331, n13330, n13329, n13328, n13327, n13326, n13325, n13324,
         n13323, n13322, n13321, n13320, n13319, n13318, n13317, n13316,
         n13315, n13314, n13313, n13312, n13311, n13310, n13309, n13308,
         n13307, n13306, n13305, n13304, n13303, n13302, n13301, n13300,
         n13299, n13298, n13297, n13296, n13295, n13294, n13293, n13292,
         n13291, n13290, n13289, n13288, n13287, n13286, n13285, n13284,
         n13283, n13282, n13281, n13280, n13279, n13278, n13277, n13276,
         n13275, n13274, n13273, n13272, n13271, n13270, n13269, n13268,
         n13267, n13266, n13265, n13264, n13263, n13262, n13261, n13260,
         n13259, n13258, n13257, n13256, n13255, n13254, n13253, n13252,
         n13251, n13250, n13249, n13248, n13247, n13246, n13245, n13244,
         n13243, n13242, n13241, n13240, n13239, n13238, n13237, n13236,
         n13235, n13234, n13233, n13232, n13231, n13230, n13229, n13228,
         n13227, n13226, n13225, n13224, n13223, n13222, n13221, n13220,
         n13219, n13218, n13217, n13216, n13215, n13214, n13213, n13212,
         n13211, n13210, n13209, n13208, n13207, n13206, n13205, n13204,
         n13203, n13202, n13201, n13200, n13199, n13198, n13197, n13196,
         n13195, n13194, n13193, n13192, n13191, n13190, n13189, n13188,
         n13187, n13186, n13185, n13184, n13183, n13182, n13181, n13180,
         n13179, n13178, n13176, n13175, n13174, n13173, n13172, n13171,
         n13170, n13169, n13168, n13167, n13166, n13165, n13164, n13163,
         n13162, n13161, n13160, n13159, n13158, n13157, n13156, n13155,
         n13154, n13153, n13152, n13151, n13150, n13149, n13148, n13147,
         n13146, n13145, n13144, n13143, n13142, n13141, n13140, n13139,
         n13138, n13137, n13136, n13135, n13134, n13133, n13132, n13131,
         n13130, n13129, n13128, n13127, n13126, n13125, n13124, n13123,
         n13122, n13121, n13120, n13119, n13118, n13117, n13116, n13115,
         n13114, n13113, n13112, n13111, n13110, n13109, n13108, n13107,
         n13106, n13105, n13104, n13103, n13102, n13101, n13100, n13099,
         n13098, n13097, n13096, n13095, n13094, n13093, n13092, n13091,
         n13090, n13089, n13088, n13087, n13086, n13085, n13084, n13083,
         n13082, n13081, n13080, n13078, n13077, n13076, n13075, n13074,
         n13073, n13072, n13071, n13070, n13069, n13068, n13067, n13066,
         n13065, n13064, n13063, n13062, n13061, n13060, n13059, n13058,
         n13057, n13056, n13055, n13054, n13053, n13052, n13051, n13050,
         n13049, n13048, n13047, n13046, n13045, n13044, n13043, n13042,
         n13041, n13040, n13039, n13038, n13037, n13036, n13035, n13034,
         n13033, n13032, n13031, n13030, n13029, n13028, n13027, n13026,
         n13025, n13024, n13023, n13022, n13021, n13020, n13019, n13018,
         n13017, n13016, n13015, n13014, n13013, n13012, n13011, n13010,
         n13009, n13008, n13007, n13006, n13005, n13004, n13003, n13002,
         n13001, n13000, n12999, n12998, n12997, n12996, n12995, n12994,
         n12993, n12992, n12991, n12990, n12989, n12988, n12987, n12986,
         n12985, n12984, n12983, n12982, n12981, n12980, n12979, n12978,
         n12977, n12976, n12975, n12974, n12973, n12972, n12971, n12970,
         n12969, n12968, n12967, n12966, n12965, n12964, n12963, n12962,
         n12961, n12960, n12959, n12958, n12957, n12956, n12955, n12954,
         n12953, n12952, n12951, n12950, n12949, n12948, n12947, n12946,
         n12945, n12944, n12943, n12942, n12941, n12940, n12939, n12938,
         n12937, n12936, n12935, n12934, n12933, n12932, n12931, n12930,
         n12929, n12928, n12927, n12926, n12925, n12924, n12923, n12922,
         n12921, n12920, n12919, n12918, n12917, n12916, n12915, n12914,
         n12913, n12912, n12911, n12910, n12909, n12908, n12907, n12906,
         n12905, n12904, n12903, n12902, n12901, n12900, n12899, n12898,
         n12897, n12896, n12895, n12894, n12893, n12892, n12891, n12890,
         n12889, n12888, n12887, n12885, n12884, n12883, n12882, n12881,
         n12880, n12879, n12878, n12877, n12876, n12875, n12874, n12873,
         n12872, n12871, n12870, n12869, n12868, n12867, n12866, n12865,
         n12864, n12863, n12862, n12861, n12860, n12859, n12858, n12857,
         n12856, n12855, n12854, n12853, n12852, n12851, n12850, n12849,
         n12848, n12847, n12846, n12845, n12844, n12843, n12842, n12841,
         n12840, n12839, n12838, n12837, n12836, n12835, n12834, n12833,
         n12832, n12831, n12830, n12829, n12828, n12827, n12826, n12825,
         n12824, n12823, n12822, n12821, n12820, n12819, n12818, n12817,
         n12816, n12815, n12814, n12813, n12812, n12811, n12810, n12809,
         n12808, n12807, n12806, n12805, n12804, n12803, n12802, n12801,
         n12800, n12799, n12798, n12797, n12796, n12795, n12794, n12793,
         n12792, n12791, n12790, n12789, n12788, n12787, n12786, n12785,
         n12784, n12783, n12782, n12781, n12780, n12779, n12778, n12777,
         n12776, n12775, n12774, n12773, n12772, n12771, n12770, n12769,
         n12768, n12767, n12766, n12765, n12764, n12763, n12762, n12761,
         n12760, n12759, n12758, n12757, n12756, n12755, n12754, n12753,
         n12752, n12751, n12750, n12749, n12748, n12747, n12746, n12745,
         n12744, n12743, n12742, n12741, n12740, n12739, n12738, n12737,
         n12736, n12735, n12734, n12733, n12732, n12731, n12730, n12728,
         n12727, n12726, n12725, n12724, n12723, n12721, n12720, n12719,
         n12718, n12717, n12716, n12715, n12714, n12713, n12712, n12711,
         n12710, n12709, n12708, n12707, n12706, n12705, n12704, n12703,
         n12701, n12700, n12699, n12698, n12697, n12696, n12695, n12694,
         n12693, n12692, n12691, n12690, n12689, n12688, n12687, n12686,
         n12685, n12684, n12683, n12682, n12681, n12680, n12679, n12678,
         n12676, n12675, n12674, n12673, n12672, n12671, n12670, n12669,
         n12668, n12667, n12666, n12665, n12664, n12663, n12662, n12661,
         n12660, n12659, n12658, n12657, n12656, n12655, n12654, n12653,
         n12652, n12651, n12650, n12649, n12648, n12647, n12646, n12645,
         n12644, n12643, n12642, n12641, n12640, n12639, n12638, n12637,
         n12636, n12635, n12634, n12633, n12632, n12631, n12630, n12629,
         n12628, n12627, n12626, n12625, n12624, n12623, n12622, n12621,
         n12620, n12619, n12618, n12617, n12616, n12615, n12614, n12613,
         n12612, n12611, n12610, n12609, n12608, n12607, n12606, n12605,
         n12604, n12603, n12602, n12601, n12600, n12599, n12598, n12597,
         n12596, n12595, n12594, n12593, n12592, n12591, n12590, n12589,
         n12588, n12587, n12586, n12585, n12584, n12583, n12582, n12581,
         n12580, n12579, n12578, n12577, n12576, n12575, n12574, n12573,
         n12572, n12571, n12570, n12569, n12568, n12567, n12566, n12565,
         n12564, n12563, n12562, n12561, n12560, n12559, n12558, n12556,
         n12555, n12554, n12553, n12552, n12551, n12550, n12549, n12548,
         n12547, n12546, n12545, n12544, n12543, n12542, n12541, n12540,
         n12539, n12538, n12537, n12536, n12535, n12534, n12533, n12532,
         n12531, n12530, n12529, n12528, n12527, n12526, n12525, n12524,
         n12523, n12522, n12521, n12520, n12519, n12518, n12517, n12516,
         n12515, n12514, n12513, n12512, n12511, n12510, n12509, n12508,
         n12507, n12506, n12505, n12504, n12503, n12502, n12501, n12500,
         n12499, n12498, n12497, n12496, n12495, n12494, n12493, n12492,
         n12491, n12490, n12489, n12488, n12487, n12486, n12485, n12484,
         n12483, n12482, n12481, n12480, n12479, n12478, n12477, n12476,
         n12475, n12474, n12473, n12472, n12471, n12470, n12469, n12468,
         n12467, n12466, n12465, n12464, n12463, n12462, n12461, n12460,
         n12459, n12458, n12457, n12456, n12455, n12454, n12453, n12452,
         n12451, n12450, n12449, n12448, n12447, n12446, n12445, n12444,
         n12443, n12442, n12441, n12440, n12439, n12438, n12437, n12436,
         n12435, n12434, n12433, n12432, n12431, n12430, n12429, n12428,
         n12427, n12426, n12425, n12424, n12423, n12422, n12421, n12420,
         n12419, n12418, n12417, n12416, n12415, n12414, n12413, n12412,
         n12411, n12410, n12409, n12408, n12407, n12406, n12405, n12404,
         n12403, n12402, n12401, n12400, n12399, n12398, n12397, n12396,
         n12395, n12394, n12393, n12392, n12391, n12390, n12389, n12388,
         n12387, n12386, n12385, n12384, n12383, n12382, n12381, n12380,
         n12379, n12378, n12377, n12376, n12375, n12374, n12373, n12372,
         n12371, n12370, n12369, n12368, n12367, n12366, n12365, n12364,
         n12363, n12362, n12361, n12360, n12359, n12358, n12357, n12356,
         n12355, n12354, n12353, n12352, n12351, n12350, n12349, n12348,
         n12347, n12346, n12345, n12344, n12343, n12342, n12341, n12340,
         n12339, n12338, n12337, n12336, n12335, n12334, n12333, n12332,
         n12331, n12330, n12329, n12328, n12327, n12326, n12325, n12324,
         n12323, n12322, n12321, n12320, n12319, n12318, n12317, n12316,
         n12315, n12314, n12313, n12312, n12311, n12310, n12309, n12308,
         n12307, n12306, n12305, n12304, n12303, n12302, n12301, n12300,
         n12299, n12298, n12297, n12296, n12295, n12294, n12293, n12292,
         n12291, n12290, n12289, n12288, n12287, n12286, n12285, n12284,
         n12283, n12282, n12281, n12280, n12279, n12278, n12277, n12276,
         n12275, n12274, n12273, n12272, n12271, n12270, n12269, n12268,
         n12267, n12266, n12265, n12264, n12263, n12262, n12261, n12259,
         n12258, n12257, n12256, n12255, n12254, n12253, n12252, n12251,
         n12250, n12249, n12248, n12247, n12246, n12245, n12244, n12243,
         n12242, n12241, n12240, n12239, n12238, n12237, n12236, n12235,
         n12234, n12233, n12232, n12231, n12230, n12229, n12228, n12227,
         n12226, n12225, n12224, n12223, n12222, n12221, n12220, n12219,
         n12218, n12217, n12216, n12215, n12214, n12213, n12212, n12211,
         n12210, n12209, n12208, n12207, n12206, n12205, n12204, n12203,
         n12202, n12201, n12200, n12199, n12198, n12197, n12196, n12195,
         n12194, n12193, n12192, n12191, n12190, n12189, n12188, n12187,
         n12186, n12185, n12184, n12183, n12182, n12181, n12180, n12179,
         n12178, n12177, n12176, n12175, n12174, n12173, n12172, n12171,
         n12170, n12169, n12168, n12167, n12166, n12165, n12164, n12163,
         n12162, n12161, n12160, n12159, n12158, n12157, n12156, n12155,
         n12154, n12153, n12152, n12151, n12150, n12149, n12148, n12147,
         n12146, n12145, n12144, n12143, n12142, n12141, n12140, n12139,
         n12138, n12137, n12136, n12135, n12134, n12133, n12132, n12131,
         n12130, n12129, n12128, n12127, n12126, n12125, n12124, n12123,
         n12122, n12121, n12120, n12119, n12118, n12117, n12116, n12115,
         n12114, n12113, n12112, n12111, n12110, n12109, n12108, n12107,
         n12106, n12105, n12104, n12103, n12102, n12101, n12100, n12099,
         n12098, n12097, n12096, n12095, n12094, n12093, n12092, n12091,
         n12090, n12089, n12088, n12087, n12086, n12085, n12084, n12083,
         n12082, n12081, n12080, n12079, n12078, n12077, n12076, n12075,
         n12074, n12073, n12072, n12071, n12070, n12069, n12068, n12066,
         n12065, n12064, n12063, n12062, n12061, n12060, n12059, n12058,
         n12057, n12056, n12055, n12054, n12053, n12052, n12051, n12050,
         n12049, n12048, n12047, n12046, n12045, n12044, n12043, n12042,
         n12041, n12040, n12039, n12038, n12037, n12036, n12035, n12034,
         n12033, n12032, n12031, n12030, n12029, n12028, n12027, n12026,
         n12025, n12024, n12023, n12022, n12021, n12020, n12019, n12018,
         n12017, n12016, n12015, n12014, n12013, n12012, n12011, n12010,
         n12009, n12008, n12007, n12006, n12005, n12004, n12003, n12002,
         n12001, n12000, n11999, n11998, n11997, n11996, n11995, n11994,
         n11993, n11992, n11991, n11990, n11989, n11988, n11987, n11986,
         n11985, n11984, n11983, n11982, n11981, n11980, n11979, n11978,
         n11977, n11976, n11975, n11974, n11973, n11972, n11971, n11970,
         n11969, n11968, n11967, n11966, n11965, n11964, n11963, n11962,
         n11961, n11960, n11959, n11958, n11957, n11956, n11955, n11954,
         n11953, n11952, n11951, n11950, n11949, n11948, n11947, n11946,
         n11945, n11944, n11943, n11942, n11941, n11940, n11939, n11938,
         n11937, n11936, n11935, n11934, n11933, n11932, n11931, n11930,
         n11929, n11928, n11927, n11926, n11925, n11924, n11923, n11922,
         n11921, n11920, n11919, n11918, n11917, n11916, n11915, n11914,
         n11913, n11912, n11911, n11909, n11908, n11907, n11906, n11905,
         n11904, n11902, n11901, n11900, n11899, n11898, n11897, n11896,
         n11895, n11894, n11893, n11892, n11891, n11890, n11889, n11888,
         n11887, n11886, n11885, n11884, n11882, n11881, n11880, n11879,
         n11878, n11877, n11876, n11875, n11874, n11873, n11872, n11871,
         n11870, n11869, n11868, n11867, n11866, n11865, n11864, n11863,
         n11862, n11861, n11860, n11859, n11857, n11856, n11855, n11854,
         n11853, n11852, n11851, n11850, n11849, n11848, n11847, n11846,
         n11845, n11844, n11843, n11842, n11841, n11840, n11839, n11838,
         n11837, n11836, n11835, n11834, n11833, n11832, n11831, n11830,
         n11829, n11828, n11827, n11826, n11825, n11824, n11823, n11822,
         n11821, n11820, n11819, n11818, n11817, n11816, n11815, n11814,
         n11813, n11812, n11811, n11810, n11809, n11808, n11807, n11806,
         n11805, n11804, n11803, n11802, n11801, n11800, n11799, n11798,
         n11797, n11796, n11795, n11794, n11793, n11792, n11791, n11790,
         n11789, n11788, n11787, n11786, n11785, n11784, n11783, n11782,
         n11781, n11780, n11779, n11778, n11777, n11776, n11775, n11774,
         n11773, n11772, n11771, n11770, n11769, n11768, n11767, n11766,
         n11765, n11764, n11763, n11762, n11761, n11760, n11759, n11758,
         n11757, n11756, n11755, n11754, n11753, n11752, n11751, n11750,
         n11749, n11748, n11747, n11746, n11745, n11744, n11743, n11742,
         n11741, n11740, n11739, n11737, n11736, n11735, n11734, n11733,
         n11732, n11731, n11730, n11729, n11728, n11727, n11726, n11725,
         n11724, n11723, n11722, n11721, n11720, n11719, n11718, n11717,
         n11716, n11715, n11714, n11713, n11712, n11711, n11710, n11709,
         n11708, n11707, n11706, n11705, n11704, n11703, n11702, n11701,
         n11700, n11699, n11698, n11697, n11696, n11695, n11694, n11693,
         n11692, n11691, n11690, n11689, n11688, n11687, n11686, n11685,
         n11684, n11683, n11682, n11681, n11680, n11679, n11678, n11677,
         n11676, n11675, n11674, n11673, n11672, n11671, n11670, n11669,
         n11668, n11667, n11666, n11665, n11664, n11663, n11662, n11661,
         n11660, n11659, n11658, n11657, n11656, n11655, n11654, n11653,
         n11652, n11651, n11650, n11649, n11648, n11647, n11646, n11645,
         n11644, n11643, n11642, n11641, n11640, n11639, n11638, n11637,
         n11636, n11635, n11634, n11633, n11632, n11631, n11630, n11629,
         n11628, n11627, n11626, n11625, n11624, n11623, n11622, n11621,
         n11620, n11619, n11618, n11617, n11616, n11615, n11614, n11613,
         n11612, n11611, n11610, n11609, n11608, n11607, n11606, n11605,
         n11604, n11603, n11602, n11601, n11600, n11599, n11598, n11597,
         n11596, n11595, n11594, n11593, n11592, n11591, n11590, n11589,
         n11588, n11587, n11586, n11585, n11584, n11583, n11582, n11581,
         n11580, n11579, n11578, n11577, n11576, n11575, n11574, n11573,
         n11572, n11571, n11570, n11569, n11568, n11567, n11566, n11565,
         n11564, n11563, n11562, n11561, n11560, n11559, n11558, n11557,
         n11556, n11555, n11554, n11553, n11552, n11551, n11550, n11549,
         n11548, n11547, n11546, n11545, n11544, n11543, n11542, n11541,
         n11540, n11538, n11537, n11536, n11535, n11534, n11533, n11532,
         n11531, n11530, n11529, n11528, n11527, n11526, n11525, n11524,
         n11523, n11522, n11521, n11520, n11519, n11518, n11517, n11516,
         n11515, n11514, n11513, n11512, n11511, n11510, n11509, n11508,
         n11507, n11506, n11505, n11504, n11503, n11502, n11501, n11500,
         n11499, n11498, n11497, n11496, n11495, n11494, n11493, n11492,
         n11491, n11490, n11489, n11488, n11487, n11486, n11485, n11484,
         n11483, n11482, n11481, n11480, n11479, n11478, n11477, n11476,
         n11475, n11474, n11473, n11472, n11471, n11470, n11469, n11468,
         n11467, n11466, n11465, n11464, n11463, n11462, n11461, n11460,
         n11459, n11458, n11457, n11456, n11455, n11454, n11453, n11452,
         n11451, n11450, n11449, n11448, n11447, n11446, n11445, n11444,
         n11443, n11442, n11440, n11439, n11438, n11437, n11436, n11435,
         n11434, n11433, n11432, n11431, n11430, n11429, n11428, n11427,
         n11426, n11425, n11424, n11423, n11422, n11421, n11420, n11419,
         n11418, n11417, n11416, n11415, n11414, n11413, n11412, n11411,
         n11410, n11409, n11408, n11407, n11406, n11405, n11404, n11403,
         n11402, n11401, n11400, n11399, n11398, n11397, n11396, n11395,
         n11394, n11393, n11392, n11391, n11390, n11389, n11388, n11387,
         n11386, n11385, n11384, n11383, n11382, n11381, n11380, n11379,
         n11378, n11377, n11376, n11375, n11374, n11373, n11372, n11371,
         n11370, n11369, n11368, n11367, n11366, n11365, n11364, n11363,
         n11362, n11361, n11360, n11359, n11358, n11357, n11356, n11355,
         n11354, n11353, n11352, n11351, n11350, n11349, n11348, n11347,
         n11346, n11345, n11344, n11343, n11342, n11341, n11340, n11339,
         n11338, n11337, n11336, n11335, n11334, n11333, n11332, n11331,
         n11330, n11329, n11328, n11327, n11326, n11325, n11324, n11323,
         n11322, n11321, n11320, n11319, n11318, n11317, n11316, n11315,
         n11314, n11313, n11312, n11311, n11310, n11309, n11308, n11307,
         n11306, n11305, n11304, n11303, n11302, n11301, n11300, n11299,
         n11298, n11297, n11296, n11295, n11294, n11293, n11292, n11291,
         n11290, n11289, n11288, n11287, n11286, n11285, n11284, n11283,
         n11282, n11281, n11280, n11279, n11278, n11277, n11276, n11275,
         n11274, n11273, n11272, n11271, n11270, n11269, n11268, n11267,
         n11266, n11265, n11264, n11263, n11262, n11261, n11260, n11259,
         n11258, n11257, n11256, n11255, n11254, n11253, n11252, n11251,
         n11250, n11249, n11247, n11246, n11245, n11244, n11243, n11242,
         n11241, n11240, n11239, n11238, n11237, n11236, n11235, n11234,
         n11233, n11232, n11231, n11230, n11229, n11228, n11227, n11226,
         n11225, n11224, n11223, n11222, n11221, n11220, n11219, n11218,
         n11217, n11216, n11215, n11214, n11213, n11212, n11211, n11210,
         n11209, n11208, n11207, n11206, n11205, n11204, n11203, n11202,
         n11201, n11200, n11199, n11198, n11197, n11196, n11195, n11194,
         n11193, n11192, n11191, n11190, n11189, n11188, n11187, n11186,
         n11185, n11184, n11183, n11182, n11181, n11180, n11179, n11178,
         n11176, n11175, n11174, n11173, n11172, n11171, n11170, n11169,
         n11168, n11167, n11166, n11165, n11164, n11163, n11162, n11161,
         n11160, n11159, n11158, n11157, n11156, n11155, n11154, n11153,
         n11152, n11151, n11150, n11149, n11148, n11147, n11146, n11145,
         n11144, n11143, n11142, n11141, n11140, n11139, n11138, n11137,
         n11136, n11135, n11134, n11133, n11132, n11131, n11130, n11129,
         n11128, n11127, n11126, n11125, n11124, n11123, n11122, n11121,
         n11120, n11119, n11118, n11117, n11116, n11115, n11114, n11113,
         n11112, n11111, n11110, n11109, n11108, n11107, n11106, n11105,
         n11104, n11103, n11102, n11101, n11100, n11099, n11098, n11097,
         n11096, n11095, n11094, n11093, n11092, n11090, n11089, n11088,
         n11087, n11086, n11085, n11083, n11082, n11081, n11080, n11079,
         n11078, n11077, n11076, n11075, n11074, n11073, n11072, n11071,
         n11070, n11069, n11068, n11067, n11066, n11065, n11063, n11062,
         n11061, n11060, n11059, n11058, n11057, n11056, n11055, n11054,
         n11053, n11052, n11051, n11050, n11049, n11048, n11047, n11046,
         n11045, n11044, n11043, n11042, n11041, n11040, n11038, n11037,
         n11036, n11035, n11034, n11033, n11032, n11031, n11030, n11029,
         n11028, n11027, n11026, n11025, n11024, n11023, n11022, n11021,
         n11020, n11019, n11018, n11017, n11016, n11015, n11014, n11013,
         n11012, n11011, n11010, n11009, n11008, n11007, n11006, n11005,
         n11004, n11003, n11002, n11001, n11000, n10999, n10998, n10997,
         n10996, n10995, n10994, n10993, n10992, n10991, n10990, n10989,
         n10988, n10987, n10986, n10985, n10984, n10983, n10982, n10981,
         n10980, n10979, n10978, n10977, n10976, n10975, n10974, n10973,
         n10972, n10971, n10970, n10969, n10968, n10967, n10966, n10965,
         n10964, n10963, n10962, n10961, n10960, n10959, n10958, n10957,
         n10956, n10955, n10954, n10953, n10952, n10951, n10950, n10949,
         n10948, n10947, n10946, n10945, n10944, n10943, n10942, n10941,
         n10940, n10939, n10938, n10937, n10936, n10935, n10934, n10933,
         n10932, n10931, n10930, n10929, n10928, n10927, n10926, n10925,
         n10924, n10923, n10922, n10921, n10920, n10918, n10917, n10916,
         n10915, n10914, n10913, n10912, n10911, n10910, n10909, n10908,
         n10907, n10906, n10905, n10904, n10903, n10902, n10901, n10900,
         n10899, n10898, n10897, n10896, n10895, n10894, n10893, n10892,
         n10891, n10890, n10889, n10888, n10887, n10886, n10885, n10884,
         n10883, n10882, n10881, n10880, n10879, n10878, n10877, n10876,
         n10875, n10874, n10873, n10872, n10871, n10870, n10869, n10868,
         n10867, n10866, n10865, n10864, n10863, n10862, n10861, n10860,
         n10859, n10858, n10857, n10856, n10855, n10854, n10853, n10852,
         n10851, n10850, n10849, n10848, n10847, n10846, n10845, n10844,
         n10843, n10842, n10841, n10840, n10839, n10838, n10837, n10836,
         n10835, n10834, n10833, n10832, n10831, n10830, n10829, n10828,
         n10827, n10826, n10825, n10824, n10823, n10822, n10821, n10820,
         n10819, n10818, n10817, n10816, n10815, n10814, n10813, n10812,
         n10811, n10810, n10809, n10808, n10807, n10806, n10805, n10804,
         n10803, n10802, n10801, n10800, n10799, n10798, n10797, n10796,
         n10795, n10794, n10793, n10792, n10791, n10790, n10789, n10788,
         n10787, n10786, n10785, n10784, n10783, n10782, n10781, n10780,
         n10779, n10778, n10777, n10776, n10775, n10774, n10773, n10772,
         n10771, n10770, n10769, n10768, n10767, n10766, n10765, n10764,
         n10763, n10762, n10761, n10760, n10759, n10758, n10757, n10756,
         n10755, n10754, n10753, n10752, n10751, n10750, n10749, n10748,
         n10747, n10746, n10745, n10744, n10743, n10742, n10741, n10740,
         n10739, n10738, n10737, n10736, n10735, n10734, n10733, n10732,
         n10731, n10730, n10729, n10728, n10727, n10726, n10725, n10724,
         n10723, n10722, n10721, n10720, n10719, n10718, n10717, n10716,
         n10715, n10714, n10713, n10712, n10711, n10710, n10709, n10708,
         n10707, n10706, n10705, n10704, n10703, n10702, n10701, n10700,
         n10699, n10698, n10697, n10696, n10695, n10694, n10693, n10692,
         n10691, n10690, n10689, n10688, n10687, n10686, n10685, n10684,
         n10683, n10682, n10681, n10680, n10679, n10678, n10677, n10676,
         n10675, n10674, n10673, n10672, n10671, n10670, n10669, n10668,
         n10667, n10666, n10665, n10664, n10663, n10662, n10661, n10660,
         n10659, n10658, n10657, n10656, n10655, n10654, n10653, n10652,
         n10651, n10650, n10649, n10648, n10647, n10646, n10645, n10644,
         n10643, n10642, n10641, n10640, n10639, n10638, n10637, n10636,
         n10635, n10634, n10633, n10632, n10631, n10630, n10629, n10628,
         n10627, n10626, n10625, n10624, n10623, n10621, n10620, n10619,
         n10618, n10617, n10616, n10615, n10614, n10613, n10612, n10611,
         n10610, n10609, n10608, n10607, n10606, n10605, n10604, n10603,
         n10602, n10601, n10600, n10599, n10598, n10597, n10596, n10595,
         n10594, n10593, n10592, n10591, n10590, n10589, n10588, n10587,
         n10586, n10585, n10584, n10583, n10582, n10581, n10580, n10579,
         n10578, n10577, n10576, n10575, n10574, n10573, n10572, n10571,
         n10570, n10569, n10568, n10567, n10566, n10565, n10564, n10563,
         n10562, n10561, n10560, n10559, n10558, n10557, n10556, n10555,
         n10554, n10553, n10552, n10551, n10550, n10549, n10548, n10547,
         n10546, n10545, n10544, n10543, n10542, n10541, n10540, n10539,
         n10538, n10537, n10536, n10535, n10534, n10533, n10532, n10531,
         n10530, n10529, n10528, n10527, n10526, n10525, n10524, n10523,
         n10522, n10521, n10520, n10519, n10518, n10517, n10516, n10515,
         n10514, n10513, n10512, n10511, n10510, n10509, n10508, n10507,
         n10506, n10505, n10504, n10503, n10502, n10501, n10500, n10499,
         n10498, n10497, n10496, n10495, n10494, n10493, n10492, n10491,
         n10490, n10489, n10488, n10487, n10486, n10485, n10484, n10483,
         n10482, n10481, n10480, n10479, n10478, n10477, n10476, n10475,
         n10474, n10473, n10472, n10471, n10470, n10469, n10468, n10467,
         n10466, n10465, n10464, n10463, n10462, n10461, n10460, n10459,
         n10458, n10457, n10456, n10455, n10454, n10453, n10452, n10451,
         n10450, n10449, n10448, n10447, n10446, n10445, n10444, n10443,
         n10442, n10441, n10440, n10439, n10438, n10437, n10436, n10435,
         n10434, n10433, n10432, n10431, n10430, n10428, n10427, n10426,
         n10425, n10424, n10423, n10422, n10421, n10420, n10419, n10418,
         n10417, n10416, n10415, n10414, n10413, n10412, n10411, n10410,
         n10409, n10408, n10407, n10406, n10405, n10404, n10403, n10402,
         n10401, n10400, n10399, n10398, n10397, n10396, n10395, n10394,
         n10393, n10392, n10391, n10390, n10389, n10388, n10387, n10386,
         n10385, n10384, n10383, n10382, n10381, n10380, n10379, n10378,
         n10377, n10376, n10375, n10374, n10373, n10372, n10371, n10370,
         n10369, n10368, n10367, n10366, n10365, n10364, n10363, n10362,
         n10361, n10360, n10359, n10358, n10357, n10356, n10355, n10354,
         n10353, n10352, n10351, n10350, n10349, n10348, n10347, n10346,
         n10345, n10344, n10343, n10342, n10341, n10340, n10339, n10338,
         n10337, n10336, n10335, n10334, n10333, n10332, n10331, n10330,
         n10329, n10328, n10327, n10326, n10325, n10324, n10323, n10322,
         n10321, n10320, n10319, n10318, n10317, n10316, n10315, n10314,
         n10313, n10312, n10311, n10310, n10309, n10308, n10307, n10306,
         n10305, n10304, n10303, n10302, n10301, n10300, n10299, n10298,
         n10297, n10296, n10295, n10294, n10293, n10292, n10291, n10290,
         n10289, n10288, n10287, n10286, n10285, n10284, n10283, n10282,
         n10281, n10280, n10279, n10278, n10277, n10276, n10275, n10274,
         n10273, n10272, n10271, n10270, n10269, n10268, n10267, n10266,
         n10264, n10263, n10262, n10261, n10260, n10259, n10258, n10257,
         n10256, n10255, n10254, n10253, n10252, n10251, n10250, n10249,
         n10248, n10247, n10246, n10244, n10243, n10242, n10241, n10240,
         n10239, n10238, n10237, n10236, n10235, n10234, n10233, n10232,
         n10231, n10230, n10229, n10228, n10227, n10226, n10225, n10224,
         n10223, n10222, n10221, n10219, n10218, n10217, n10216, n10215,
         n10214, n10213, n10212, n10211, n10210, n10209, n10208, n10207,
         n10206, n10205, n10204, n10203, n10202, n10201, n10200, n10199,
         n10198, n10197, n10196, n10195, n10194, n10193, n10192, n10191,
         n10190, n10189, n10188, n10187, n10186, n10185, n10184, n10183,
         n10182, n10181, n10180, n10179, n10178, n10177, n10176, n10175,
         n10174, n10173, n10172, n10171, n10170, n10169, n10168, n10167,
         n10166, n10165, n10164, n10163, n10162, n10161, n10160, n10159,
         n10158, n10157, n10156, n10155, n10154, n10153, n10152, n10151,
         n10150, n10149, n10148, n10147, n10146, n10145, n10144, n10143,
         n10142, n10141, n10140, n10139, n10138, n10137, n10136, n10135,
         n10134, n10133, n10132, n10131, n10130, n10129, n10128, n10127,
         n10126, n10125, n10124, n10123, n10122, n10121, n10120, n10119,
         n10118, n10117, n10116, n10115, n10114, n10113, n10112, n10111,
         n10110, n10109, n10108, n10107, n10106, n10105, n10104, n10103,
         n10102, n10101, n10099, n10098, n10097, n10096, n10095, n10094,
         n10093, n10092, n10091, n10090, n10089, n10088, n10087, n10086,
         n10085, n10084, n10083, n10082, n10081, n10080, n10079, n10078,
         n10077, n10076, n10075, n10074, n10073, n10072, n10071, n10070,
         n10069, n10068, n10067, n10066, n10065, n10064, n10063, n10062,
         n10061, n10060, n10059, n10058, n10057, n10056, n10055, n10054,
         n10053, n10052, n10051, n10050, n10049, n10048, n10047, n10046,
         n10045, n10044, n10043, n10042, n10041, n10040, n10039, n10038,
         n10037, n10036, n10035, n10034, n10033, n10032, n10031, n10030,
         n10029, n10028, n10027, n10026, n10025, n10024, n10023, n10022,
         n10021, n10020, n10019, n10018, n10017, n10016, n10015, n10014,
         n10013, n10012, n10011, n10010, n10009, n10008, n10007, n10006,
         n10005, n10004, n10003, n10002, n10001, n10000, \L2_0/n3608 ,
         \L2_0/n3604 , \L2_0/n3600 , \L2_0/n3596 , \L2_0/n3592 , \L2_0/n3588 ,
         \L2_0/n3584 , \L2_0/n3580 , \L2_0/n3576 , \L2_0/n3572 , \L2_0/n3568 ,
         \L2_0/n3564 , \L2_0/n3560 , \L2_0/n3556 , \L2_0/n3552 , \L2_0/n3548 ,
         \L2_0/n3544 , \L2_0/n3540 , \L2_0/n3536 , \L2_0/n3532 , \L2_0/n3531 ,
         \L2_0/n3524 , \L2_0/n3523 , \L2_0/n3520 , \L2_0/n3519 , \L2_0/n3516 ,
         \L2_0/n3515 , \L2_0/n3512 , \L2_0/n3511 , \L2_0/n3508 , \L2_0/n3507 ,
         \L2_0/n3504 , \L2_0/n3503 , \L2_0/n3500 , \L2_0/n3499 , \L2_0/n3496 ,
         \L2_0/n3495 , \L2_0/n3492 , \L2_0/n3491 , \L2_0/n3488 , \L2_0/n3487 ,
         \L2_0/n3484 , \L2_0/n3483 , \L2_0/n3480 , \L2_0/n3479 , \L2_0/n3476 ,
         \L2_0/n3475 , \L2_0/n3472 , \L2_0/n3471 , \L2_0/n3468 , \L2_0/n3467 ,
         \L2_0/n3464 , \L2_0/n3463 , \L2_0/n3460 , \L2_0/n3459 , \L2_0/n3456 ,
         \L2_0/n3455 , \L2_0/n3452 , \L2_0/n3451 , \L2_0/n3447 , \L2_0/n3444 ,
         \L2_0/n3443 , \L2_0/n3440 , \L2_0/n3439 , \L2_0/n3436 , \L2_0/n3435 ,
         \L2_0/n3432 , \L2_0/n3431 , \L2_0/n3428 , \L2_0/n3427 , \L2_0/n3424 ,
         \L2_0/n3423 , \L2_0/n3420 , \L2_0/n3419 , \L2_0/n3416 , \L2_0/n3415 ,
         \L2_0/n3412 , \L2_0/n3411 , \L2_0/n3408 , \L2_0/n3407 , \L2_0/n3404 ,
         \L2_0/n3403 , \L2_0/n3400 , \L2_0/n3399 , \L2_0/n3396 , \L2_0/n3395 ,
         \L2_0/n3392 , \L2_0/n3391 , \L2_0/n3388 , \L2_0/n3387 , \L2_0/n3384 ,
         \L2_0/n3383 , \L2_0/n3380 , \L2_0/n3379 , \L2_0/n3376 , \L2_0/n3375 ,
         \L2_0/n3372 , \L2_0/n3371 , \L2_0/n3367 , \L2_0/n3364 , \L2_0/n3363 ,
         \L2_0/n3360 , \L2_0/n3359 , \L2_0/n3356 , \L2_0/n3355 , \L2_0/n3352 ,
         \L2_0/n3351 , \L2_0/n3348 , \L2_0/n3347 , \L2_0/n3344 , \L2_0/n3343 ,
         \L2_0/n3340 , \L2_0/n3339 , \L2_0/n3336 , \L2_0/n3335 , \L2_0/n3332 ,
         \L2_0/n3331 , \L2_0/n3328 , \L2_0/n3327 , \L2_0/n3324 , \L2_0/n3323 ,
         \L2_0/n3320 , \L2_0/n3319 , \L2_0/n3316 , \L2_0/n3315 , \L2_0/n3312 ,
         \L2_0/n3311 , \L2_0/n3308 , \L2_0/n3307 , \L2_0/n3304 , \L2_0/n3303 ,
         \L2_0/n3300 , \L2_0/n3299 , \L2_0/n3296 , \L2_0/n3295 , \L2_0/n3292 ,
         \L2_0/n3291 , \L2_0/n3284 , \L2_0/n3283 , \L2_0/n3280 , \L2_0/n3279 ,
         \L2_0/n3276 , \L2_0/n3275 , \L2_0/n3272 , \L2_0/n3271 , \L2_0/n3268 ,
         \L2_0/n3267 , \L2_0/n3264 , \L2_0/n3263 , \L2_0/n3260 , \L2_0/n3259 ,
         \L2_0/n3256 , \L2_0/n3255 , \L2_0/n3252 , \L2_0/n3251 , \L2_0/n3248 ,
         \L2_0/n3247 , \L2_0/n3244 , \L2_0/n3243 , \L2_0/n3240 , \L2_0/n3239 ,
         \L2_0/n3236 , \L2_0/n3235 , \L2_0/n3232 , \L2_0/n3231 , \L2_0/n3228 ,
         \L2_0/n3227 , \L2_0/n3224 , \L2_0/n3223 , \L2_0/n3220 , \L2_0/n3219 ,
         \L2_0/n3216 , \L2_0/n3215 , \L2_0/n3212 , \L2_0/n3211 , \L2_0/n3204 ,
         \L2_0/n3203 , \L2_0/n3200 , \L2_0/n3199 , \L2_0/n3196 , \L2_0/n3195 ,
         \L2_0/n3192 , \L2_0/n3191 , \L2_0/n3188 , \L2_0/n3187 , \L2_0/n3184 ,
         \L2_0/n3183 , \L2_0/n3180 , \L2_0/n3179 , \L2_0/n3176 , \L2_0/n3175 ,
         \L2_0/n3172 , \L2_0/n3171 , \L2_0/n3168 , \L2_0/n3167 , \L2_0/n3164 ,
         \L2_0/n3163 , \L2_0/n3160 , \L2_0/n3159 , \L2_0/n3156 , \L2_0/n3155 ,
         \L2_0/n3152 , \L2_0/n3151 , \L2_0/n3148 , \L2_0/n3147 , \L2_0/n3144 ,
         \L2_0/n3143 , \L2_0/n3140 , \L2_0/n3139 , \L2_0/n3136 , \L2_0/n3135 ,
         \L2_0/n3132 , \L2_0/n3131 , \L2_0/n3127 , \L2_0/n3124 , \L2_0/n3123 ,
         \L2_0/n3120 , \L2_0/n3119 , \L2_0/n3116 , \L2_0/n3115 , \L2_0/n3112 ,
         \L2_0/n3111 , \L2_0/n3108 , \L2_0/n3107 , \L2_0/n3104 , \L2_0/n3103 ,
         \L2_0/n3100 , \L2_0/n3099 , \L2_0/n3096 , \L2_0/n3095 , \L2_0/n3092 ,
         \L2_0/n3091 , \L2_0/n3088 , \L2_0/n3087 , \L2_0/n3084 , \L2_0/n3083 ,
         \L2_0/n3080 , \L2_0/n3079 , \L2_0/n3076 , \L2_0/n3075 , \L2_0/n3072 ,
         \L2_0/n3071 , \L2_0/n3068 , \L2_0/n3067 , \L2_0/n3064 , \L2_0/n3063 ,
         \L2_0/n3060 , \L2_0/n3059 , \L2_0/n3056 , \L2_0/n3055 , \L2_0/n3052 ,
         \L2_0/n3051 , \L2_0/n3047 , \L2_0/n3044 , \L2_0/n3043 , \L2_0/n3040 ,
         \L2_0/n3039 , \L2_0/n3036 , \L2_0/n3035 , \L2_0/n3032 , \L2_0/n3031 ,
         \L2_0/n3028 , \L2_0/n3027 , \L2_0/n3024 , \L2_0/n3023 , \L2_0/n3020 ,
         \L2_0/n3019 , \L2_0/n3016 , \L2_0/n3015 , \L2_0/n3012 , \L2_0/n3011 ,
         \L2_0/n3008 , \L2_0/n3007 , \L2_0/n3004 , \L2_0/n3003 , \L2_0/n3000 ,
         \L2_0/n2999 , \L2_0/n2996 , \L2_0/n2995 , \L2_0/n2992 , \L2_0/n2991 ,
         \L2_0/n2988 , \L2_0/n2987 , \L2_0/n2984 , \L2_0/n2983 , \L2_0/n2980 ,
         \L2_0/n2979 , \L2_0/n2976 , \L2_0/n2975 , \L2_0/n2972 , \L2_0/n2971 ,
         \L2_0/n2967 , \L2_0/n2964 , \L2_0/n2963 , \L2_0/n2960 , \L2_0/n2959 ,
         \L2_0/n2956 , \L2_0/n2955 , \L2_0/n2952 , \L2_0/n2951 , \L2_0/n2948 ,
         \L2_0/n2947 , \L2_0/n2944 , \L2_0/n2943 , \L2_0/n2940 , \L2_0/n2939 ,
         \L2_0/n2936 , \L2_0/n2935 , \L2_0/n2932 , \L2_0/n2931 , \L2_0/n2928 ,
         \L2_0/n2927 , \L2_0/n2924 , \L2_0/n2923 , \L2_0/n2920 , \L2_0/n2919 ,
         \L2_0/n2916 , \L2_0/n2915 , \L2_0/n2912 , \L2_0/n2911 , \L2_0/n2908 ,
         \L2_0/n2907 , \L2_0/n2904 , \L2_0/n2903 , \L2_0/n2900 , \L2_0/n2899 ,
         \L2_0/n2896 , \L2_0/n2895 , \L2_0/n2892 , \L2_0/n2891 , \L2_0/n2884 ,
         \L2_0/n2883 , \L2_0/n2880 , \L2_0/n2879 , \L2_0/n2876 , \L2_0/n2875 ,
         \L2_0/n2872 , \L2_0/n2871 , \L2_0/n2868 , \L2_0/n2867 , \L2_0/n2864 ,
         \L2_0/n2863 , \L2_0/n2860 , \L2_0/n2859 , \L2_0/n2856 , \L2_0/n2855 ,
         \L2_0/n2852 , \L2_0/n2851 , \L2_0/n2848 , \L2_0/n2847 , \L2_0/n2844 ,
         \L2_0/n2843 , \L2_0/n2840 , \L2_0/n2839 , \L2_0/n2836 , \L2_0/n2835 ,
         \L2_0/n2832 , \L2_0/n2831 , \L2_0/n2828 , \L2_0/n2827 , \L2_0/n2824 ,
         \L2_0/n2823 , \L2_0/n2820 , \L2_0/n2819 , \L2_0/n2816 , \L2_0/n2815 ,
         \L2_0/n2812 , \L2_0/n2811 , \L2_0/n2804 , \L2_0/n2803 , \L2_0/n2800 ,
         \L2_0/n2799 , \L2_0/n2796 , \L2_0/n2795 , \L2_0/n2792 , \L2_0/n2791 ,
         \L2_0/n2788 , \L2_0/n2787 , \L2_0/n2784 , \L2_0/n2783 , \L2_0/n2780 ,
         \L2_0/n2779 , \L2_0/n2776 , \L2_0/n2775 , \L2_0/n2772 , \L2_0/n2771 ,
         \L2_0/n2768 , \L2_0/n2767 , \L2_0/n2764 , \L2_0/n2763 , \L2_0/n2760 ,
         \L2_0/n2759 , \L2_0/n2756 , \L2_0/n2755 , \L2_0/n2752 , \L2_0/n2751 ,
         \L2_0/n2748 , \L2_0/n2747 , \L2_0/n2744 , \L2_0/n2743 , \L2_0/n2740 ,
         \L2_0/n2739 , \L2_0/n2736 , \L2_0/n2735 , \L2_0/n2732 , \L2_0/n2731 ,
         \L2_0/n2727 , \L2_0/n2724 , \L2_0/n2723 , \L2_0/n2720 , \L2_0/n2719 ,
         \L2_0/n2716 , \L2_0/n2715 , \L2_0/n2712 , \L2_0/n2711 , \L2_0/n2708 ,
         \L2_0/n2707 , \L2_0/n2704 , \L2_0/n2703 , \L2_0/n2700 , \L2_0/n2699 ,
         \L2_0/n2696 , \L2_0/n2695 , \L2_0/n2692 , \L2_0/n2691 , \L2_0/n2688 ,
         \L2_0/n2687 , \L2_0/n2684 , \L2_0/n2683 , \L2_0/n2680 , \L2_0/n2679 ,
         \L2_0/n2676 , \L2_0/n2675 , \L2_0/n2672 , \L2_0/n2671 , \L2_0/n2668 ,
         \L2_0/n2667 , \L2_0/n2664 , \L2_0/n2663 , \L2_0/n2660 , \L2_0/n2659 ,
         \L2_0/n2656 , \L2_0/n2655 , \L2_0/n2652 , \L2_0/n2651 , \L2_0/n2644 ,
         \L2_0/n2643 , \L2_0/n2640 , \L2_0/n2639 , \L2_0/n2636 , \L2_0/n2635 ,
         \L2_0/n2632 , \L2_0/n2631 , \L2_0/n2628 , \L2_0/n2627 , \L2_0/n2624 ,
         \L2_0/n2623 , \L2_0/n2620 , \L2_0/n2619 , \L2_0/n2616 , \L2_0/n2615 ,
         \L2_0/n2612 , \L2_0/n2611 , \L2_0/n2608 , \L2_0/n2607 , \L2_0/n2604 ,
         \L2_0/n2603 , \L2_0/n2600 , \L2_0/n2599 , \L2_0/n2596 , \L2_0/n2595 ,
         \L2_0/n2592 , \L2_0/n2591 , \L2_0/n2588 , \L2_0/n2587 , \L2_0/n2584 ,
         \L2_0/n2583 , \L2_0/n2580 , \L2_0/n2579 , \L2_0/n2576 , \L2_0/n2575 ,
         \L2_0/n2572 , \L2_0/n2571 , \L2_0/n2564 , \L2_0/n2563 , \L2_0/n2560 ,
         \L2_0/n2559 , \L2_0/n2556 , \L2_0/n2555 , \L2_0/n2552 , \L2_0/n2551 ,
         \L2_0/n2548 , \L2_0/n2547 , \L2_0/n2544 , \L2_0/n2543 , \L2_0/n2540 ,
         \L2_0/n2539 , \L2_0/n2536 , \L2_0/n2535 , \L2_0/n2532 , \L2_0/n2531 ,
         \L2_0/n2528 , \L2_0/n2527 , \L2_0/n2524 , \L2_0/n2523 , \L2_0/n2520 ,
         \L2_0/n2519 , \L2_0/n2516 , \L2_0/n2515 , \L2_0/n2512 , \L2_0/n2511 ,
         \L2_0/n2508 , \L2_0/n2507 , \L2_0/n2504 , \L2_0/n2503 , \L2_0/n2500 ,
         \L2_0/n2499 , \L2_0/n2496 , \L2_0/n2495 , \L2_0/n2492 , \L2_0/n2491 ,
         \L2_0/n2484 , \L2_0/n2483 , \L2_0/n2480 , \L2_0/n2479 , \L2_0/n2476 ,
         \L2_0/n2475 , \L2_0/n2472 , \L2_0/n2471 , \L2_0/n2468 , \L2_0/n2467 ,
         \L2_0/n2464 , \L2_0/n2463 , \L2_0/n2460 , \L2_0/n2459 , \L2_0/n2456 ,
         \L2_0/n2455 , \L2_0/n2452 , \L2_0/n2451 , \L2_0/n2448 , \L2_0/n2447 ,
         \L2_0/n2444 , \L2_0/n2443 , \L2_0/n2440 , \L2_0/n2439 , \L2_0/n2436 ,
         \L2_0/n2435 , \L2_0/n2432 , \L2_0/n2431 , \L2_0/n2428 , \L2_0/n2427 ,
         \L2_0/n2424 , \L2_0/n2423 , \L2_0/n2420 , \L2_0/n2419 , \L2_0/n2416 ,
         \L2_0/n2415 , \L2_0/n2412 , \L2_0/n2411 , \L2_0/n2404 , \L2_0/n2403 ,
         \L2_0/n2400 , \L2_0/n2399 , \L2_0/n2396 , \L2_0/n2395 , \L2_0/n2392 ,
         \L2_0/n2391 , \L2_0/n2388 , \L2_0/n2387 , \L2_0/n2384 , \L2_0/n2383 ,
         \L2_0/n2380 , \L2_0/n2379 , \L2_0/n2376 , \L2_0/n2375 , \L2_0/n2372 ,
         \L2_0/n2371 , \L2_0/n2368 , \L2_0/n2367 , \L2_0/n2364 , \L2_0/n2363 ,
         \L2_0/n2360 , \L2_0/n2359 , \L2_0/n2356 , \L2_0/n2355 , \L2_0/n2352 ,
         \L2_0/n2351 , \L2_0/n2348 , \L2_0/n2347 , \L2_0/n2344 , \L2_0/n2343 ,
         \L2_0/n2340 , \L2_0/n2339 , \L2_0/n2336 , \L2_0/n2335 , \L2_0/n2292 ,
         \L1_0/n4511 , \L1_0/n4507 , \L1_0/n4503 , \L1_0/n4499 , \L1_0/n4495 ,
         \L1_0/n4491 , \L1_0/n4487 , \L1_0/n4483 , \L1_0/n4479 , \L1_0/n4475 ,
         \L1_0/n4471 , \L1_0/n4467 , \L1_0/n4463 , \L1_0/n4459 , \L1_0/n4455 ,
         \L1_0/n4451 , \L1_0/n4447 , \L1_0/n4443 , \L1_0/n4439 , \L1_0/n4436 ,
         \L1_0/n4432 , \L1_0/n4428 , \L1_0/n4424 , \L1_0/n4420 , \L1_0/n4416 ,
         \L1_0/n4412 , \L1_0/n4404 , \L1_0/n4400 , \L1_0/n4396 , \L1_0/n4392 ,
         \L1_0/n4388 , \L1_0/n4384 , \L1_0/n4380 , \L1_0/n4376 , \L1_0/n4372 ,
         \L1_0/n4368 , \L1_0/n4364 , \L1_0/n4356 , \L1_0/n4355 , \L1_0/n4352 ,
         \L1_0/n4351 , \L1_0/n4348 , \L1_0/n4347 , \L1_0/n4344 , \L1_0/n4343 ,
         \L1_0/n4340 , \L1_0/n4339 , \L1_0/n4336 , \L1_0/n4335 , \L1_0/n4332 ,
         \L1_0/n4331 , \L1_0/n4328 , \L1_0/n4327 , \L1_0/n4324 , \L1_0/n4323 ,
         \L1_0/n4320 , \L1_0/n4319 , \L1_0/n4316 , \L1_0/n4315 , \L1_0/n4312 ,
         \L1_0/n4311 , \L1_0/n4308 , \L1_0/n4307 , \L1_0/n4304 , \L1_0/n4303 ,
         \L1_0/n4300 , \L1_0/n4299 , \L1_0/n4296 , \L1_0/n4295 , \L1_0/n4292 ,
         \L1_0/n4291 , \L1_0/n4288 , \L1_0/n4287 , \L1_0/n4284 , \L1_0/n4283 ,
         \L1_0/n4280 , \L1_0/n4279 , \L1_0/n4276 , \L1_0/n4275 , \L1_0/n4272 ,
         \L1_0/n4271 , \L1_0/n4268 , \L1_0/n4267 , \L1_0/n4264 , \L1_0/n4263 ,
         \L1_0/n4260 , \L1_0/n4259 , \L1_0/n4256 , \L1_0/n4255 , \L1_0/n4252 ,
         \L1_0/n4251 , \L1_0/n4248 , \L1_0/n4247 , \L1_0/n4244 , \L1_0/n4243 ,
         \L1_0/n4240 , \L1_0/n4239 , \L1_0/n4236 , \L1_0/n4235 , \L1_0/n4232 ,
         \L1_0/n4231 , \L1_0/n4228 , \L1_0/n4227 , \L1_0/n4224 , \L1_0/n4223 ,
         \L1_0/n4220 , \L1_0/n4219 , \L1_0/n4216 , \L1_0/n4215 , \L1_0/n4212 ,
         \L1_0/n4211 , \L1_0/n4208 , \L1_0/n4207 , \L1_0/n4204 , \L1_0/n4203 ,
         \L1_0/n4200 , \L1_0/n4199 , \L1_0/n4196 , \L1_0/n4195 , \L1_0/n4192 ,
         \L1_0/n4191 , \L1_0/n4188 , \L1_0/n4187 , \L1_0/n4184 , \L1_0/n4183 ,
         \L1_0/n4180 , \L1_0/n4179 , \L1_0/n4176 , \L1_0/n4175 , \L1_0/n4172 ,
         \L1_0/n4171 , \L1_0/n4168 , \L1_0/n4167 , \L1_0/n4164 , \L1_0/n4163 ,
         \L1_0/n4160 , \L1_0/n4159 , \L1_0/n4156 , \L1_0/n4155 , \L1_0/n4152 ,
         \L1_0/n4151 , \L1_0/n4148 , \L1_0/n4147 , \L1_0/n4144 , \L1_0/n4143 ,
         \L1_0/n4140 , \L1_0/n4139 , \L1_0/n4136 , \L1_0/n4135 , \L1_0/n4132 ,
         \L1_0/n4131 , \L1_0/n4128 , \L1_0/n4127 , \L1_0/n4124 , \L1_0/n4123 ,
         \L1_0/n4120 , \L1_0/n4119 , \L1_0/n4116 , \L1_0/n4115 , \L1_0/n4112 ,
         \L1_0/n4111 , \L1_0/n4108 , \L1_0/n4107 , \L1_0/n4104 , \L1_0/n4103 ,
         \L1_0/n4100 , \L1_0/n4099 , \L1_0/n4096 , \L1_0/n4095 , \L1_0/n4092 ,
         \L1_0/n4091 , \L1_0/n4088 , \L1_0/n4087 , \L1_0/n4084 , \L1_0/n4083 ,
         \L1_0/n4080 , \L1_0/n4079 , \L1_0/n4076 , \L1_0/n4075 , \L1_0/n4072 ,
         \L1_0/n4071 , \L1_0/n4068 , \L1_0/n4067 , \L1_0/n4064 , \L1_0/n4063 ,
         \L1_0/n4060 , \L1_0/n4059 , \L1_0/n4056 , \L1_0/n4055 , \L1_0/n4052 ,
         \L1_0/n4051 , \L1_0/n4048 , \L1_0/n4047 , \L1_0/n4044 , \L1_0/n4043 ,
         \L1_0/n4040 , \L1_0/n4039 , \L1_0/n4036 , \L1_0/n4035 , \L1_0/n4032 ,
         \L1_0/n4031 , \L1_0/n4028 , \L1_0/n4027 , \L1_0/n4024 , \L1_0/n4023 ,
         \L1_0/n4020 , \L1_0/n4019 , \L1_0/n4016 , \L1_0/n4015 , \L1_0/n4012 ,
         \L1_0/n4011 , \L1_0/n4008 , \L1_0/n4007 , \L1_0/n4004 , \L1_0/n4003 ,
         \L1_0/n4000 , \L1_0/n3999 , \L1_0/n3996 , \L1_0/n3995 , \L1_0/n3992 ,
         \L1_0/n3991 , \L1_0/n3988 , \L1_0/n3987 , \L1_0/n3984 , \L1_0/n3983 ,
         \L1_0/n3980 , \L1_0/n3979 , \L1_0/n3976 , \L1_0/n3975 , \L1_0/n3972 ,
         \L1_0/n3971 , \L1_0/n3968 , \L1_0/n3967 , \L1_0/n3964 , \L1_0/n3963 ,
         \L1_0/n3960 , \L1_0/n3959 , \L1_0/n3956 , \L1_0/n3955 , \L1_0/n3952 ,
         \L1_0/n3951 , \L1_0/n3948 , \L1_0/n3947 , \L1_0/n3944 , \L1_0/n3943 ,
         \L1_0/n3940 , \L1_0/n3939 , \L1_0/n3936 , \L1_0/n3935 , \L1_0/n3932 ,
         \L1_0/n3931 , \L1_0/n3928 , \L1_0/n3927 , \L1_0/n3924 , \L1_0/n3923 ,
         \L1_0/n3920 , \L1_0/n3919 , \L1_0/n3916 , \L1_0/n3915 , \L1_0/n3912 ,
         \L1_0/n3911 , \L1_0/n3908 , \L1_0/n3907 , \L1_0/n3904 , \L1_0/n3903 ,
         \L1_0/n3900 , \L1_0/n3899 , \L1_0/n3896 , \L1_0/n3895 , \L1_0/n3892 ,
         \L1_0/n3891 , \L1_0/n3888 , \L1_0/n3887 , \L1_0/n3884 , \L1_0/n3883 ,
         \L1_0/n3880 , \L1_0/n3879 , \L1_0/n3876 , \L1_0/n3875 , \L1_0/n3872 ,
         \L1_0/n3871 , \L1_0/n3868 , \L1_0/n3867 , \L1_0/n3864 , \L1_0/n3863 ,
         \L1_0/n3860 , \L1_0/n3859 , \L1_0/n3856 , \L1_0/n3855 , \L1_0/n3852 ,
         \L1_0/n3851 , \L1_0/n3848 , \L1_0/n3847 , \L1_0/n3844 , \L1_0/n3843 ,
         \L1_0/n3840 , \L1_0/n3839 , \L1_0/n3836 , \L1_0/n3835 , \L1_0/n3832 ,
         \L1_0/n3831 , \L1_0/n3828 , \L1_0/n3827 , \L1_0/n3824 , \L1_0/n3823 ,
         \L1_0/n3820 , \L1_0/n3819 , \L1_0/n3816 , \L1_0/n3815 , \L1_0/n3812 ,
         \L1_0/n3811 , \L1_0/n3808 , \L1_0/n3807 , \L1_0/n3804 , \L1_0/n3803 ,
         \L1_0/n3800 , \L1_0/n3799 , \L1_0/n3796 , \L1_0/n3795 , \L1_0/n3792 ,
         \L1_0/n3791 , \L1_0/n3788 , \L1_0/n3787 , \L1_0/n3784 , \L1_0/n3783 ,
         \L1_0/n3780 , \L1_0/n3779 , \L1_0/n3776 , \L1_0/n3775 , \L1_0/n3772 ,
         \L1_0/n3771 , \L1_0/n3768 , \L1_0/n3767 , \L1_0/n3764 , \L1_0/n3763 ,
         \L1_0/n3760 , \L1_0/n3759 , \L1_0/n3756 , \L1_0/n3755 , \L1_0/n3752 ,
         \L1_0/n3751 , \L1_0/n3748 , \L1_0/n3747 , \L1_0/n3744 , \L1_0/n3743 ,
         \L1_0/n3740 , \L1_0/n3739 , \L1_0/n3736 , \L1_0/n3735 , \L1_0/n3732 ,
         \L1_0/n3731 , \L1_0/n3728 , \L1_0/n3727 , \L1_0/n3724 , \L1_0/n3723 ,
         \L1_0/n3720 , \L1_0/n3719 , \L1_0/n3716 , \L1_0/n3715 , \L1_0/n3712 ,
         \L1_0/n3711 , \L1_0/n3708 , \L1_0/n3707 , \L1_0/n3704 , \L1_0/n3703 ,
         \L1_0/n3700 , \L1_0/n3699 , \L1_0/n3696 , \L1_0/n3695 , \L1_0/n3692 ,
         \L1_0/n3691 , \L1_0/n3688 , \L1_0/n3687 , \L1_0/n3684 , \L1_0/n3683 ,
         \L1_0/n3680 , \L1_0/n3679 , \L1_0/n3676 , \L1_0/n3675 , \L1_0/n3672 ,
         \L1_0/n3671 , \L1_0/n3668 , \L1_0/n3667 , \L1_0/n3664 , \L1_0/n3663 ,
         \L1_0/n3660 , \L1_0/n3659 , \L1_0/n3656 , \L1_0/n3655 , \L1_0/n3652 ,
         \L1_0/n3651 , \L1_0/n3648 , \L1_0/n3647 , \L1_0/n3644 , \L1_0/n3643 ,
         \L1_0/n3640 , \L1_0/n3639 , \L1_0/n3636 , \L1_0/n3635 , \L1_0/n3632 ,
         \L1_0/n3631 , \L1_0/n3628 , \L1_0/n3627 , \L1_0/n3624 , \L1_0/n3623 ,
         \L1_0/n3620 , \L1_0/n3619 , \L1_0/n3616 , \L1_0/n3615 , \L1_0/n3612 ,
         \L1_0/n3611 , \L1_0/n3608 , \L1_0/n3607 , \L1_0/n3604 , \L1_0/n3603 ,
         \L1_0/n3600 , \L1_0/n3599 , \L1_0/n3596 , \L1_0/n3595 , \L1_0/n3592 ,
         \L1_0/n3591 , \L1_0/n3588 , \L1_0/n3587 , \L1_0/n3584 , \L1_0/n3583 ,
         \L1_0/n3580 , \L1_0/n3579 , \L1_0/n3576 , \L1_0/n3575 , \L1_0/n3572 ,
         \L1_0/n3571 , \L1_0/n3568 , \L1_0/n3567 , \L1_0/n3564 , \L1_0/n3563 ,
         \L1_0/n3560 , \L1_0/n3559 , \L1_0/n3556 , \L1_0/n3555 , \L1_0/n3552 ,
         \L1_0/n3551 , \L1_0/n3548 , \L1_0/n3547 , \L1_0/n3544 , \L1_0/n3543 ,
         \L1_0/n3540 , \L1_0/n3539 , \L1_0/n3536 , \L1_0/n3535 , \L1_0/n3532 ,
         \L1_0/n3531 , \L1_0/n3528 , \L1_0/n3527 , \L1_0/n3524 , \L1_0/n3523 ,
         \L1_0/n3520 , \L1_0/n3519 , \L1_0/n3516 , \L1_0/n3515 , \L1_0/n3512 ,
         \L1_0/n3511 , \L1_0/n3508 , \L1_0/n3507 , \L1_0/n3504 , \L1_0/n3503 ,
         \L1_0/n3500 , \L1_0/n3499 , \L1_0/n3496 , \L1_0/n3495 , \L1_0/n3492 ,
         \L1_0/n3491 , \L1_0/n3488 , \L1_0/n3487 , \L1_0/n3484 , \L1_0/n3483 ,
         \L1_0/n3480 , \L1_0/n3479 , \L1_0/n3476 , \L1_0/n3472 , \L1_0/n3468 ,
         \L1_0/n3464 , \L1_0/n3460 , \L1_0/n3456 , \L1_0/n3452 , \L1_0/n3440 ,
         \L1_0/n3432 , \L1_0/n3424 , \L1_0/n3416 , \L1_0/n3412 , \L1_0/n3408 ,
         \L1_0/n3404 , \L1_0/n3400 , \L1_0/n3396 , \L1_0/n3395 , \L1_0/n3392 ,
         \L1_0/n3388 , \L1_0/n3384 , \L1_0/n3380 , \L1_0/n3376 , \L1_0/n3372 ,
         \L1_0/n3367 , \L1_0/n3363 , \L1_0/n3360 , \L1_0/n3355 , \L1_0/n3352 ,
         \L1_0/n3347 , \L1_0/n3344 , \L1_0/n3339 , \L1_0/n3336 , \L1_0/n3332 ,
         \L1_0/n3328 , \L1_0/n3324 , \L1_0/n3320 , \L1_0/n3319 , \L1_0/n3316 ,
         \L1_0/n3315 , \L1_0/n3312 , \L1_0/n3311 , \L1_0/n3308 , \L1_0/n3307 ,
         \L1_0/n3304 , \L1_0/n3303 , \L1_0/n3300 , \L1_0/n3299 , \L1_0/n3296 ,
         \L1_0/n3295 , \L1_0/n3292 , \L1_0/n3291 , \L1_0/n3288 , \L1_0/n3287 ,
         \L1_0/n3284 , \L1_0/n3283 , \L1_0/n3280 , \L1_0/n3279 , \L1_0/n3276 ,
         \L1_0/n3275 , \L1_0/n3272 , \L1_0/n3271 , \L1_0/n3268 , \L1_0/n3267 ,
         \L1_0/n3264 , \L1_0/n3263 , \L1_0/n3260 , \L1_0/n3259 , \L1_0/n3256 ,
         \L1_0/n3255 , \L1_0/n3252 , \L1_0/n3251 , \L1_0/n3248 , \L1_0/n3247 ,
         \L1_0/n3244 , \L1_0/n3243 , \L1_0/n3240 , \L1_0/n3239 , \L1_0/n3195 ,
         n38121, n38122, n38123, n38124, n38125, n38126, n38127, n38128,
         n38129, n38130, n38131, n38132, n38133, n38134, n38135, n38136,
         n38137, n38138, n38139, n38140, n38141, n38142, n38143, n38144,
         n38145, n38146, n38147, n38148, n38149, n38150, n38151, n38152,
         n38153, n38154, n38155, n38156, n38157, n38158, n38159, n38160,
         n38161, n38162, n38163, n38164, n38165, n38166, n38167, n38168,
         n38169, n38170, n38171, n38172, n38173, n38174, n38175, n38176,
         n38177, n38178, n38179, n38180, n38181, n38182, n38183, n38184,
         n38185, n38186, n38187, n38188, n38189, n38190, n38191, n38192,
         n38193, n38194, n38195, n38196, n38197, n38198, n38199, n38200,
         n38201, n38202, n38203, n38204, n38205, n38206, n38207, n38208,
         n38209, n38210, n38211, n38212, n38213, n38214, n38215, n38216,
         n38217, n38218, n38219, n38220, n38221, n38222, n38223, n38224,
         n38225, n38226, n38227, n38228, n38229, n38230, n38231, n38232,
         n38233, n38234, n38235, n38236, n38237, n38238, n38239, n38240,
         n38241, n38242, n38243, n38244, n38245, n38246, n38247, n38248,
         n38249, n38250, n38251, n38252, n38253, n38254, n38255, n38256,
         n38257, n38258, n38259, n38260, n38261, n38262, n38263, n38264,
         n38265, n38266, n38267, n38268, n38269, n38270, n38271, n38272,
         n38273, n38274, n38275, n38276, n38277, n38278, n38279, n38280,
         n38281, n38282, n38283, n38284, n38285, n38286, n38287, n38288,
         n38289, n38290, n38291, n38292, n38293, n38294, n38295, n38296,
         n38297, n38298, n38299, n38300, n38301, n38302, n38303, n38304,
         n38305, n38306, n38307, n38308, n38309, n38310, n38311, n38312,
         n38313, n38314, n38315, n38316, n38317, n38318, n38319, n38320,
         n38321, n38322, n38323, n38324, n38325, n38326, n38327, n38328,
         n38329, n38330, n38331, n38332, n38333, n38334, n38335, n38336,
         n38337, n38338, n38339, n38340, n38341, n38342, n38343, n38344,
         n38345, n38346, n38347, n38348, n38349, n38350, n38351, n38352,
         n38353, n38354, n38355, n38356, n38357, n38358, n38359, n38360,
         n38361, n38362, n38363, n38364, n38365, n38366, n38367, n38368,
         n38369, n38370, n38371, n38372, n38373, n38374, n38375, n38376,
         n38377, n38378, n38379, n38380, n38381, n38382, n38383, n38384,
         n38385, n38386, n38387, n38388, n38389, n38390, n38391, n38392,
         n38393, n38394, n38395, n38396, n38397, n38398, n38399, n38400,
         n38401, n38402, n38403, n38404, n38405, n38406, n38407, n38408,
         n38409, n38410, n38411, n38412, n38413, n38414, n38415, n38416,
         n38417, n38418, n38419, n38420, n38421, n38422, n38423, n38424,
         n38425, n38426, n38427, n38428, n38429, n38430, n38431, n38432,
         n38433, n38434, n38435, n38436, n38437, n38438, n38439, n38440,
         n38441, n38442, n38443, n38444, n38445, n38446, n38447, n38448,
         n38449, n38450, n38451, n38452, n38453, n38454, n38455, n38456,
         n38457, n38458, n38459, n38460, n38461, n38462, n38463, n38464,
         n38465, n38466, n38467, n38468, n38469, n38470, n38471, n38472,
         n38473, n38474, n38475, n38476, n38477, n38478, n38479, n38480,
         n38481, n38482, n38483, n38484, n38485, n38486, n38487, n38488,
         n38489, n38490, n38491, n38492, n38493, n38494, n38495, n38496,
         n38497, n38498, n38499, n38500, n38501, n38502, n38503, n38504,
         n38505, n38506, n38507, n38508, n38509, n38510, n38511, n38512,
         n38513, n38514, n38515, n38516, n38517, n38518, n38519, n38520,
         n38521, n38522, n38523, n38524, n38525, n38526, n38527, n38528,
         n38529, n38530, n38531, n38532, n38533, n38534, n38535, n38536,
         n38537, n38538, n38539, n38540, n38541, n38542, n38543, n38544,
         n38545, n38546, n38547, n38548, n38549, n38550, n38551, n38552,
         n38553, n38554, n38555, n38556, n38557, n38558, n38559, n38560,
         n38561, n38562, n38563, n38564, n38565, n38566, n38567, n38568,
         n38569, n38570, n38571, n38572, n38573, n38574, n38575, n38576,
         n38577, n38578, n38579, n38580, n38581, n38582, n38583, n38584,
         n38585, n38586, n38587, n38588, n38589, n38590, n38591, n38592,
         n38593, n38594, n38595, n38596, n38597, n38598, n38599, n38600,
         n38601, n38602, n38603, n38604, n38605, n38606, n38607, n38608,
         n38609, n38610, n38611, n38612, n38613, n38614, n38615, n38616,
         n38617, n38618, n38619, n38620, n38621, n38622, n38623, n38624,
         n38625, n38626, n38627, n38628, n38629, n38630, n38631, n38632,
         n38633, n38634, n38635, n38636, n38637, n38638, n38639, n38640,
         n38641, n38642, n38643, n38644, n38645, n38646, n38647, n38648,
         n38649, n38650, n38651, n38652, n38653, n38654, n38655, n38656,
         n38657, n38658, n38659, n38660, n38661, n38662, n38663, n38664,
         n38665, n38666, n38667, n38668, n38669, n38670, n38671, n38672,
         n38673, n38674, n38675, n38676, n38677, n38678, n38679, n38680,
         n38681, n38682, n38683, n38684, n38685, n38686, n38687, n38688,
         n38689, n38690, n38691, n38692, n38693, n38694, n38695, n38696,
         n38697, n38698, n38699, n38700, n38701, n38702, n38703, n38704,
         n38705, n38706, n38707, n38708, n38709, n38710, n38711, n38712,
         n38713, n38714, n38715, n38716, n38717, n38718, n38719, n38720,
         n38721, n38722, n38723, n38724, n38725, n38726, n38727, n38728,
         n38729, n38730, n38731, n38732, n38733, n38734, n38735, n38736,
         n38737, n38738, n38739, n38740, n38741, n38742, n38743, n38744,
         n38745, n38746, n38747, n38748, n38749, n38750, n38751, n38752,
         n38753, n38754, n38755, n38756, n38757, n38758, n38759, n38760,
         n38761, n38762, n38763, n38764, n38765, n38766, n38767, n38768,
         n38769, n38770, n38771, n38772, n38773, n38774, n38775, n38776,
         n38777, n38778, n38779, n38780, n38781, n38782, n38783, n38784,
         n38785, n38786, n38787, n38788, n38789, n38790, n38791, n38792,
         n38793, n38794, n38795, n38796, n38797, n38798, n38799, n38800,
         n38801, n38802, n38803, n38804, n38805, n38806, n38807, n38808,
         n38809, n38810, n38811, n38812, n38813, n38814, n38815, n38816,
         n38817, n38818, n38819, n38820, n38821, n38822, n38823, n38824,
         n38825, n38826, n38827, n38828, n38829, n38830, n38831, n38832,
         n38833, n38834, n38835, n38836, n38837, n38838, n38839, n38840,
         n38841, n38842, n38843, n38844, n38845, n38846, n38847, n38848,
         n38849, n38850, n38851, n38852, n38853, n38854, n38855, n38856,
         n38857, n38858, n38859, n38860, n38861, n38862, n38863, n38864,
         n38865, n38866, n38867, n38868, n38869, n38870, n38871, n38872,
         n38873, n38874, n38875, n38876, n38877, n38878, n38879, n38880,
         n38881, n38882, n38883, n38884, n38885, n38886, n38887, n38888,
         n38889, n38890, n38891, n38892, n38893, n38894, n38895, n38896,
         n38897, n38898, n38899, n38900, n38901, n38902, n38903, n38904,
         n38905, n38906, n38907, n38908, n38909, n38910, n38911, n38912,
         n38913, n38914, n38915, n38916, n38917, n38918, n38919, n38920,
         n38921, n38922, n38923, n38924, n38925, n38926, n38927, n38928,
         n38929, n38930, n38931, n38932, n38933, n38934, n38935, n38936,
         n38937, n38938, n38939, n38940, n38941, n38942, n38943, n38944,
         n38945, n38946, n38947, n38948, n38949, n38950, n38951, n38952,
         n38953, n38954, n38955, n38956, n38957, n38958, n38959, n38960,
         n38961, n38962, n38963, n38964, n38965, n38966, n38967, n38968,
         n38969, n38970, n38971, n38972, n38973, n38974, n38975, n38976,
         n38977, n38978, n38979, n38980, n38981, n38982, n38983, n38984,
         n38985, n38986, n38987, n38988, n38989, n38990, n38991, n38992,
         n38993, n38994, n38995, n38996, n38997, n38998, n38999, n39000,
         n39001, n39002, n39003, n39004, n39005, n39006, n39007, n39008,
         n39009, n39010, n39011, n39012, n39013, n39014, n39015, n39016,
         n39017, n39018, n39019, n39020, n39021, n39022, n39023, n39024,
         n39025, n39026, n39027, n39028, n39029, n39030, n39031, n39032,
         n39033, n39034, n39035, n39036, n39037, n39038, n39039, n39040,
         n39041, n39042, n39043, n39044, n39045, n39046, n39047, n39048,
         n39049, n39050, n39051, n39052, n39053, n39054, n39055, n39056,
         n39057, n39058, n39059, n39060, n39061, n39062, n39063, n39064,
         n39065, n39066, n39067, n39068, n39069, n39070, n39071, n39072,
         n39073, n39074, n39075, n39076, n39077, n39078, n39079, n39080,
         n39081, n39082, n39083, n39084, n39085, n39086, n39087, n39088,
         n39089, n39090, n39091, n39092, n39093, n39094, n39095, n39096,
         n39097, n39098, n39099, n39100, n39101, n39102, n39103, n39104,
         n39105, n39106, n39107, n39108, n39109, n39110, n39111, n39112,
         n39113, n39114, n39115, n39116, n39117, n39118, n39119, n39120,
         n39121, n39122, n39123, n39124, n39125, n39126, n39127, n39128,
         n39129, n39130, n39131, n39132, n39133, n39134, n39135, n39136,
         n39137, n39138, n39139, n39140, n39141, n39142, n39143, n39144,
         n39145, n39146, n39147, n39148, n39149, n39150, n39151, n39152,
         n39153, n39154, n39155, n39156, n39157, n39158, n39159, n39160,
         n39161, n39162, n39163, n39164, n39165, n39166, n39167, n39168,
         n39169, n39170, n39171, n39172, n39173, n39174, n39175, n39176,
         n39177, n39178, n39179, n39180, n39181, n39182, n39183, n39184,
         n39185, n39186, n39187, n39188, n39189, n39190, n39191, n39192,
         n39193, n39194, n39195, n39196, n39197, n39198, n39199, n39200,
         n39201, n39202, n39203, n39204, n39205, n39206, n39207, n39208,
         n39209, n39210, n39211, n39212, n39213, n39214, n39215, n39216,
         n39217, n39218, n39219, n39220, n39221, n39222, n39223, n39224,
         n39225, n39226, n39227, n39228, n39229, n39230, n39231, n39232,
         n39233, n39234, n39235, n39236, n39237, n39238, n39239, n39240,
         n39241, n39242, n39243, n39244, n39245, n39246, n39247, n39248,
         n39249, n39250, n39251, n39252, n39253, n39254, n39255, n39256,
         n39257, n39258, n39259, n39260, n39261, n39262, n39263, n39264,
         n39265, n39266, n39267, n39268, n39269, n39270, n39271, n39272,
         n39273, n39274, n39275, n39276, n39277, n39278, n39279, n39280,
         n39281, n39282, n39283, n39284, n39285, n39286, n39287, n39288,
         n39289, n39290, n39291, n39292, n39293, n39294, n39295, n39296,
         n39297, n39298, n39299, n39300, n39301, n39302, n39303, n39304,
         n39305, n39306, n39307, n39308, n39309, n39310, n39311, n39312,
         n39313, n39314, n39315, n39316, n39317, n39318, n39319, n39320,
         n39321, n39322, n39323, n39324, n39325, n39326, n39327, n39328,
         n39329, n39330, n39331, n39332, n39333, n39334, n39335, n39336,
         n39337, n39338, n39339, n39340, n39341, n39342, n39343, n39344,
         n39345, n39346, n39347, n39348, n39349, n39350, n39351, n39352,
         n39353, n39354, n39355, n39356, n39357, n39358, n39359, n39360,
         n39361, n39362, n39363, n39364, n39365, n39366, n39367, n39368,
         n39369, n39370, n39371, n39372, n39373, n39374, n39375, n39376,
         n39377, n39378, n39379, n39380, n39381, n39382, n39383, n39384,
         n39385, n39386, n39387, n39388, n39389, n39390, n39391, n39392,
         n39393, n39394, n39395, n39396, n39397, n39398, n39399, n39400,
         n39401, n39402, n39403, n39404, n39405, n39406, n39407, n39408,
         n39409, n39410, n39411, n39412, n39413, n39414, n39415, n39416,
         n39417, n39418, n39419, n39420, n39421, n39422, n39423, n39424,
         n39425, n39426, n39427, n39428, n39429, n39430, n39431, n39432,
         n39433, n39434, n39435, n39436, n39437, n39438, n39439, n39440,
         n39441, n39442, n39443, n39444, n39445, n39446, n39447, n39448,
         n39449, n39450, n39451, n39452, n39453, n39454, n39455, n39456,
         n39457, n39458, n39459, n39460, n39461, n39462, n39463, n39464,
         n39465, n39466, n39467, n39468, n39469, n39470, n39471, n39472,
         n39473, n39474, n39475, n39476, n39477, n39478, n39479, n39480,
         n39481, n39482, n39483, n39484, n39485, n39486, n39487, n39488,
         n39489, n39490, n39491, n39492, n39493, n39494, n39495, n39496,
         n39497, n39498, n39499, n39500, n39501, n39502, n39503, n39504,
         n39505, n39506, n39507, n39508, n39509, n39510, n39511, n39512,
         n39513, n39514, n39515, n39516, n39517, n39518, n39519, n39520,
         n39521, n39522, n39523, n39524, n39525, n39526, n39527, n39528,
         n39529, n39530, n39531, n39532, n39533, n39534, n39535, n39536,
         n39537, n39538, n39539, n39540, n39541, n39542, n39543, n39544,
         n39545, n39546, n39547, n39548, n39549, n39550, n39551, n39552,
         n39553, n39554, n39555, n39556, n39557, n39558, n39559, n39560,
         n39561, n39562, n39563, n39564, n39565, n39566, n39567, n39568,
         n39569, n39570, n39571, n39572, n39573, n39574, n39575, n39576,
         n39577, n39578, n39579, n39580, n39581, n39582, n39583, n39584,
         n39585, n39586, n39587, n39588, n39589, n39590, n39591, n39592,
         n39593, n39594, n39595, n39596, n39597, n39598, n39599, n39600,
         n39601, n39602, n39603, n39604, n39605, n39606, n39607, n39608,
         n39609, n39610, n39611, n39612, n39613, n39614, n39615, n39616,
         n39617, n39618, n39619, n39620, n39621, n39622, n39623, n39624,
         n39625, n39626, n39627, n39628, n39629, n39630, n39631, n39632,
         n39633, n39634, n39635, n39636, n39637, n39638, n39639, n39640,
         n39641, n39642, n39643, n39644, n39645, n39646, n39647, n39648,
         n39649, n39650, n39651, n39652, n39653, n39654, n39655, n39656,
         n39657, n39658, n39659, n39660, n39661, n39662, n39663, n39664,
         n39665, n39666, n39667, n39668, n39669, n39670, n39671, n39672,
         n39673, n39674, n39675, n39676, n39677, n39678, n39679, n39680,
         n39681, n39682, n39683, n39684, n39685, n39686, n39687, n39688,
         n39689, n39690, n39691, n39692, n39693, n39694, n39695, n39696,
         n39697, n39698, n39699, n39700, n39701, n39702, n39703, n39704,
         n39705, n39706, n39707, n39708, n39709, n39710, n39711, n39712,
         n39713, n39714, n39715, n39716, n39717, n39718, n39719, n39720,
         n39721, n39722, n39723, n39724, n39725, n39726, n39727, n39728,
         n39729, n39730, n39731, n39732, n39733, n39734, n39735, n39736,
         n39737, n39738, n39739, n39740, n39741, n39742, n39743, n39744,
         n39745, n39746, n39747, n39748, n39749, n39750, n39751, n39752,
         n39753, n39754, n39755, n39756, n39757, n39758, n39759, n39760,
         n39761, n39762, n39763, n39764, n39765, n39766, n39767, n39768,
         n39769, n39770, n39771, n39772, n39773, n39774, n39775, n39776,
         n39777, n39778, n39779, n39780, n39781, n39782, n39783, n39784,
         n39785, n39786, n39787, n39788, n39789, n39790, n39791, n39792,
         n39793, n39794, n39795, n39796, n39797, n39798, n39799, n39800,
         n39801, n39802, n39803, n39804, n39805, n39806, n39807, n39808,
         n39809, n39810, n39811, n39812, n39813, n39814, n39815, n39816,
         n39817, n39818, n39819, n39820, n39821, n39822, n39823, n39824,
         n39825, n39826, n39827, n39828, n39829, n39830, n39831, n39832,
         n39833, n39834, n39835, n39836, n39837, n39838, n39839, n39840,
         n39841, n39842, n39843, n39844, n39845, n39846, n39847, n39848,
         n39849, n39850, n39851, n39852, n39853, n39854, n39855, n39856,
         n39857, n39858, n39859, n39860, n39861, n39862, n39863, n39864,
         n39865, n39866, n39867, n39868, n39869, n39870, n39871, n39872,
         n39873, n39874, n39875, n39876, n39877, n39878, n39879, n39880,
         n39881, n39882, n39883, n39884, n39885, n39886, n39887, n39888,
         n39889, n39890, n39891, n39892, n39893, n39894, n39895, n39896,
         n39897, n39898, n39899, n39900, n39901, n39902, n39903, n39904,
         n39905, n39906, n39907, n39908, n39909, n39910, n39911, n39912,
         n39913, n39914, n39915, n39916, n39917, n39918, n39919, n39920,
         n39921, n39922, n39923, n39924, n39925, n39926, n39927, n39928,
         n39929, n39930, n39931, n39932, n39933, n39934, n39935, n39936,
         n39937, n39938, n39939, n39940, n39941, n39942, n39943, n39944,
         n39945, n39946, n39947, n39948, n39949, n39950, n39951, n39952,
         n39953, n39954, n39955, n39956, n39957, n39958, n39959, n39960,
         n39961, n39962, n39963, n39964, n39965, n39966, n39967, n39968,
         n39969, n39970, n39971, n39972, n39973, n39974, n39975, n39976,
         n39977, n39978, n39979, n39980, n39981, n39982, n39983, n39984,
         n39985, n39986, n39987, n39988, n39989, n39990, n39991, n39992,
         n39993, n39994, n39995, n39996, n39997, n39998, n39999, n40000,
         n40001, n40002, n40003, n40004, n40005, n40006, n40007, n40008,
         n40009, n40010, n40011, n40012, n40013, n40014, n40015, n40016,
         n40017, n40018, n40019, n40020, n40021, n40022, n40023, n40024,
         n40025, n40026, n40027, n40028, n40029, n40030, n40031, n40032,
         n40033, n40034, n40035, n40036, n40037, n40038, n40039, n40040,
         n40041, n40042, n40043, n40044, n40045, n40046, n40047, n40048,
         n40049, n40050, n40051, n40052, n40053, n40054, n40055, n40056,
         n40057, n40058, n40059, n40060, n40061, n40062, n40063, n40064,
         n40065, n40066, n40067, n40068, n40069, n40070, n40071, n40072,
         n40073, n40074, n40075, n40076, n40077, n40078, n40079, n40080,
         n40081, n40082, n40083, n40084, n40085, n40086, n40087, n40088,
         n40089, n40090, n40091, n40092, n40093, n40094, n40095, n40096,
         n40097, n40098, n40099, n40100, n40101, n40102, n40103, n40104,
         n40105, n40106, n40107, n40108, n40109, n40110, n40111, n40112,
         n40113, n40114, n40115, n40116, n40117, n40118, n40119, n40120,
         n40121, n40122, n40123, n40124, n40125, n40126, n40127, n40128,
         n40129, n40130, n40131, n40132, n40133, n40134, n40135, n40136,
         n40137, n40138, n40139, n40140, n40141, n40142, n40143, n40144,
         n40145, n40146, n40147, n40148, n40149, n40150, n40151, n40152,
         n40153, n40154, n40155, n40156, n40157, n40158, n40159, n40160,
         n40161, n40162, n40163, n40164, n40165, n40166, n40167, n40168,
         n40169, n40170, n40171, n40172, n40173, n40174, n40175, n40176,
         n40177, n40178, n40179, n40180, n40181, n40182, n40183, n40184,
         n40185, n40186, n40187, n40188, n40189, n40190, n40191, n40192,
         n40193, n40194, n40195, n40196, n40197, n40198, n40199, n40200,
         n40201, n40202, n40203, n40204, n40205, n40206, n40207, n40208,
         n40209, n40210, n40211, n40212, n40213, n40214, n40215, n40216,
         n40217, n40218, n40219, n40220, n40221, n40222, n40223, n40224,
         n40225, n40226, n40227, n40228, n40229, n40230, n40231, n40232,
         n40233, n40234, n40235, n40236, n40237, n40238, n40239, n40240,
         n40241, n40242, n40243, n40244, n40245, n40246, n40247, n40248,
         n40249, n40250, n40251, n40252, n40253, n40254, n40255, n40256,
         n40257, n40258, n40259, n40260, n40261, n40262, n40263, n40264,
         n40265, n40266, n40267, n40268, n40269, n40270, n40271, n40272,
         n40273, n40274, n40275, n40276, n40277, n40278, n40279, n40280,
         n40281, n40282, n40283, n40284, n40285, n40286, n40287, n40288,
         n40289, n40290, n40291, n40292, n40293, n40294, n40295, n40296,
         n40297, n40298, n40299, n40300, n40301, n40302, n40303, n40304,
         n40305, n40306, n40307, n40308, n40309, n40310, n40311, n40312,
         n40313, n40314, n40315, n40316, n40317, n40318, n40319, n40320,
         n40321, n40322, n40323, n40324, n40325, n40326, n40327, n40328,
         n40329, n40330, n40331, n40332, n40333, n40334, n40335, n40336,
         n40337, n40338, n40339, n40340, n40341, n40342, n40343, n40344,
         n40345, n40346, n40347, n40348, n40349, n40350, n40351, n40352,
         n40353, n40354, n40355, n40356, n40357, n40358, n40359, n40360,
         n40361, n40362, n40363, n40364, n40365, n40366, n40367, n40368,
         n40369, n40370, n40371, n40372, n40373, n40374, n40375, n40376,
         n40377, n40378, n40379, n40380, n40381, n40382, n40383, n40384,
         n40385, n40386, n40387, n40388, n40389, n40390, n40391, n40392,
         n40393, n40394, n40395, n40396, n40397, n40398, n40399, n40400,
         n40401, n40402, n40403, n40404, n40405, n40406, n40407, n40408,
         n40409, n40410, n40411, n40412, n40413, n40414, n40415, n40416,
         n40417, n40418, n40419, n40420, n40421, n40422, n40423, n40424,
         n40425, n40426, n40427, n40428, n40429, n40430, n40431, n40432,
         n40433, n40434, n40435, n40436, n40437, n40438, n40439, n40440,
         n40441, n40442, n40443, n40444, n40445, n40446, n40447, n40448,
         n40449, n40450, n40451, n40452, n40453, n40454, n40455, n40456,
         n40457, n40458, n40459, n40460, n40461, n40462, n40463, n40464,
         n40465, n40466, n40467, n40468, n40469, n40470, n40471, n40472,
         n40473, n40474, n40475, n40476, n40477, n40478, n40479, n40480,
         n40481, n40482, n40483, n40484, n40485, n40486, n40487, n40488,
         n40489, n40490, n40491, n40492, n40493, n40494, n40495, n40496,
         n40497, n40498, n40499, n40500, n40501, n40502, n40503, n40504,
         n40505, n40506, n40507, n40508, n40509, n40510, n40511, n40512,
         n40513, n40514, n40515, n40516, n40517, n40518, n40519, n40520,
         n40521, n40522, n40523, n40524, n40525, n40526, n40527, n40528,
         n40529, n40530, n40531, n40532, n40533, n40534, n40535, n40536,
         n40537, n40538, n40539, n40540, n40541, n40542, n40543, n40544,
         n40545, n40546, n40547, n40548, n40549, n40550, n40551, n40552,
         n40553, n40554, n40555, n40556, n40557, n40558, n40559, n40560,
         n40561, n40562, n40563, n40564, n40565, n40566, n40567, n40568,
         n40569, n40570, n40571, n40572, n40573, n40574, n40575, n40576,
         n40577, n40578, n40579, n40580, n40581, n40582, n40583, n40584,
         n40585, n40586, n40587, n40588, n40589, n40590, n40591, n40592,
         n40593, n40594, n40595, n40596, n40597, n40598, n40599, n40600,
         n40601, n40602, n40603, n40604, n40605, n40606, n40607, n40608,
         n40609, n40610, n40611, n40612, n40613, n40614, n40615, n40616,
         n40617, n40618, n40619, n40620, n40621, n40622, n40623, n40624,
         n40625, n40626, n40627, n40628, n40629, n40630, n40631, n40632,
         n40633, n40634, n40635, n40636, n40637, n40638, n40639, n40640,
         n40641, n40642, n40643, n40644, n40645, n40646, n40647, n40648,
         n40649, n40650, n40651, n40652, n40653, n40654, n40655, n40656,
         n40657, n40658, n40659, n40660, n40661, n40662, n40663, n40664,
         n40665, n40666, n40667, n40668, n40669, n40670, n40671, n40672,
         n40673, n40674, n40675, n40676, n40677, n40678, n40679, n40680,
         n40681, n40682, n40683, n40684, n40685, n40686, n40687, n40688,
         n40689, n40690, n40691, n40692, n40693, n40694, n40695, n40696,
         n40697, n40698, n40699, n40700, n40701, n40702, n40703, n40704,
         n40705, n40706, n40707, n40708, n40709, n40710, n40711, n40712,
         n40713, n40714, n40715, n40716, n40717, n40718, n40719, n40720,
         n40721, n40722, n40723, n40724, n40725, n40726, n40727, n40728,
         n40729, n40730, n40731, n40732, n40733, n40734, n40735, n40736,
         n40737, n40738, n40739, n40740, n40741, n40742, n40743, n40744,
         n40745, n40746, n40747, n40748, n40749, n40750, n40751, n40752,
         n40753, n40754, n40755, n40756, n40757, n40758, n40759, n40760,
         n40761, n40762, n40763, n40764, n40765, n40766, n40767, n40768,
         n40769, n40770, n40771, n40772, n40773, n40774, n40775, n40776,
         n40777, n40778, n40779, n40780, n40781, n40782, n40783, n40784,
         n40785, n40786, n40787, n40788, n40789, n40790, n40791, n40792,
         n40793, n40794, n40795, n40796, n40797, n40798, n40799, n40800,
         n40801, n40802, n40803, n40804, n40805, n40806, n40807, n40808,
         n40809, n40810, n40811, n40812, n40813, n40814, n40815, n40816,
         n40817, n40818, n40819, n40820, n40821, n40822, n40823, n40824,
         n40825, n40826, n40827, n40828, n40829, n40830, n40831, n40832,
         n40833, n40834, n40835, n40836, n40837, n40838, n40839, n40840,
         n40841, n40842, n40843, n40844, n40845, n40846, n40847, n40848,
         n40849, n40850, n40851, n40852, n40853, n40854, n40855, n40856,
         n40857, n40858, n40859, n40860, n40861, n40862, n40863, n40864,
         n40865, n40866, n40867, n40868, n40869, n40870, n40871, n40872,
         n40873, n40874, n40875, n40876, n40877, n40878, n40879, n40880,
         n40881, n40882, n40883, n40884, n40885, n40886, n40887, n40888,
         n40889, n40890, n40891, n40892, n40893, n40894, n40895, n40896,
         n40897, n40898, n40899, n40900, n40901, n40902, n40903, n40904,
         n40905, n40906, n40907, n40908, n40909, n40910, n40911, n40912,
         n40913, n40914, n40915, n40916, n40917, n40918, n40919, n40920,
         n40921, n40922, n40923, n40924, n40925, n40926, n40927, n40928,
         n40929, n40930, n40931, n40932, n40933, n40934, n40935, n40936,
         n40937, n40938, n40939, n40940, n40941, n40942, n40943, n40944,
         n40945, n40946, n40947, n40948, n40949, n40950, n40951, n40952,
         n40953, n40954, n40955, n40956, n40957, n40958, n40959, n40960,
         n40961, n40962, n40963, n40964, n40965, n40966, n40967, n40968,
         n40969, n40970, n40971, n40972, n40973, n40974, n40975, n40976,
         n40977, n40978, n40979, n40980, n40981, n40982, n40983, n40984,
         n40985, n40986, n40987, n40988, n40989, n40990, n40991, n40992,
         n40993, n40994, n40995, n40996, n40997, n40998, n40999, n41000,
         n41001, n41002, n41003, n41004, n41005, n41006, n41007, n41008,
         n41009, n41010, n41011, n41012, n41013, n41014, n41015, n41016,
         n41017, n41018, n41019, n41020, n41021, n41022, n41023, n41024,
         n41025, n41026, n41027, n41028, n41029, n41030, n41031, n41032,
         n41033, n41034, n41035, n41036, n41037, n41038, n41039, n41040,
         n41041, n41042, n41043, n41044, n41045, n41046, n41047, n41048,
         n41049, n41050, n41051, n41052, n41053, n41054, n41055, n41056,
         n41057, n41058, n41059, n41060, n41061, n41062, n41063, n41064,
         n41065, n41066, n41067, n41068, n41069, n41070, n41071, n41072,
         n41073, n41074, n41075, n41076, n41077, n41078, n41079, n41080,
         n41081, n41082, n41083, n41084, n41085, n41086, n41087, n41088,
         n41089, n41090, n41091, n41092, n41093, n41094, n41095, n41096,
         n41097, n41098, n41099, n41100, n41101, n41102, n41103, n41104,
         n41105, n41106, n41107, n41108, n41109, n41110, n41111, n41112,
         n41113, n41114, n41115, n41116, n41117, n41118, n41119, n41120,
         n41121, n41122, n41123, n41124, n41125, n41126, n41127, n41128,
         n41129, n41130, n41131, n41132, n41133, n41134, n41135, n41136,
         n41137, n41138, n41139, n41140, n41141, n41142, n41143, n41144,
         n41145, n41146, n41147, n41148, n41149, n41150, n41151, n41152,
         n41153, n41154, n41155, n41156, n41157, n41158, n41159, n41160,
         n41161, n41162, n41163, n41164, n41165, n41166, n41167, n41168,
         n41169, n41170, n41171, n41172, n41173, n41174, n41175, n41176,
         n41177, n41178, n41179, n41180, n41181, n41182, n41183, n41184,
         n41185, n41186, n41187, n41188, n41189, n41190, n41191, n41192,
         n41193, n41194, n41195, n41196, n41197, n41198, n41199, n41200,
         n41201, n41202, n41203, n41204, n41205, n41206, n41207, n41208,
         n41209, n41210, n41211, n41212, n41213, n41214, n41215, n41216,
         n41217, n41218, n41219, n41220, n41221, n41222, n41223, n41224,
         n41225, n41226, n41227, n41228, n41229, n41230, n41231, n41232,
         n41233, n41234, n41235, n41236, n41237, n41238, n41239, n41240,
         n41241, n41242, n41243, n41244, n41245, n41246, n41247, n41248,
         n41249, n41250, n41251, n41252, n41253, n41254, n41255, n41256,
         n41257, n41258, n41259, n41260, n41261, n41262, n41263, n41264,
         n41265, n41266, n41267, n41268, n41269, n41270, n41271, n41272,
         n41273, n41274, n41275, n41276, n41277, n41278, n41279, n41280,
         n41281, n41282, n41283, n41284, n41285, n41286, n41287, n41288,
         n41289, n41290, n41291, n41292, n41293, n41294, n41295, n41296,
         n41297, n41298, n41299, n41300, n41301, n41302, n41303, n41304,
         n41305, n41306, n41307, n41308, n41309, n41310, n41311, n41312,
         n41313, n41314, n41315, n41316, n41317, n41318, n41319, n41320,
         n41321, n41322, n41323, n41324, n41325, n41326, n41327, n41328,
         n41329, n41330, n41331, n41332, n41333, n41334, n41335, n41336,
         n41337, n41338, n41339, n41340, n41341, n41342, n41343, n41344,
         n41345, n41346, n41347, n41348, n41349, n41350, n41351, n41352,
         n41353, n41354, n41355, n41356, n41357, n41358, n41359, n41360,
         n41361, n41362, n41363, n41364, n41365, n41366, n41367, n41368,
         n41369, n41370, n41371, n41372, n41373, n41374, n41375, n41376,
         n41377, n41378, n41379, n41380, n41381, n41382, n41383, n41384,
         n41385, n41386, n41387, n41388, n41389, n41390, n41391, n41392,
         n41393, n41394, n41395, n41396, n41397, n41398, n41399, n41400,
         n41401, n41402, n41403, n41404, n41405, n41406, n41407, n41408,
         n41409, n41410, n41411, n41412, n41413, n41414, n41415, n41416,
         n41417, n41418, n41419, n41420, n41421, n41422, n41423, n41424,
         n41425, n41426, n41427, n41428, n41429, n41430, n41431, n41432,
         n41433, n41434, n41435, n41436, n41437, n41438, n41439, n41440,
         n41441, n41442, n41443, n41444, n41445, n41446, n41447, n41448,
         n41449, n41450, n41451, n41452, n41453, n41454, n41455, n41456,
         n41457, n41458, n41459, n41460, n41461, n41462, n41463, n41464,
         n41465, n41466, n41467, n41468, n41469, n41470, n41471, n41472,
         n41473, n41474, n41475, n41476, n41477, n41478, n41479, n41480,
         n41481, n41482, n41483, n41484, n41485, n41486, n41487, n41488,
         n41489, n41490, n41491, n41492, n41493, n41494, n41495, n41496,
         n41497, n41498, n41499, n41500, n41501, n41502, n41503, n41504,
         n41505, n41506, n41507, n41508, n41509, n41510, n41511, n41512,
         n41513, n41514, n41515, n41516, n41517, n41518, n41519, n41520,
         n41521, n41522, n41523, n41524, n41525, n41526, n41527, n41528,
         n41529, n41530, n41531, n41532, n41533, n41534, n41535, n41536,
         n41537, n41538, n41539, n41540, n41541, n41542, n41543, n41544,
         n41545, n41546, n41547, n41548, n41549, n41550, n41551, n41552,
         n41553, n41554, n41555, n41556, n41557, n41558, n41559, n41560,
         n41561, n41562, n41563, n41564, n41565, n41566, n41567, n41568,
         n41569, n41570, n41571, n41572, n41573, n41574, n41575, n41576,
         n41577, n41578, n41579, n41580, n41581, n41582, n41583, n41584,
         n41585, n41586, n41587, n41588, n41589, n41590, n41591, n41592,
         n41593, n41594, n41595, n41596, n41597, n41598, n41599, n41600,
         n41601, n41602, n41603, n41604, n41605, n41606, n41607, n41608,
         n41609, n41610, n41611, n41612, n41613, n41614, n41615, n41616,
         n41617, n41618, n41619, n41620, n41621, n41622, n41623, n41624,
         n41625, n41626, n41627, n41628, n41629, n41630, n41631, n41632,
         n41633, n41634, n41635, n41636, n41637, n41638, n41639, n41640,
         n41641, n41642, n41643, n41644, n41645, n41646, n41647, n41648,
         n41649, n41650, n41651, n41652, n41653, n41654, n41655, n41656,
         n41657, n41658, n41659, n41660, n41661, n41662, n41663, n41664,
         n41665, n41666, n41667, n41668, n41669, n41670, n41671, n41672,
         n41673, n41674, n41675, n41676, n41677, n41678, n41679, n41680,
         n41681, n41682, n41683, n41684, n41685, n41686, n41687, n41688,
         n41689, n41690, n41691, n41692, n41693, n41694, n41695, n41696,
         n41697, n41698, n41699, n41700, n41701, n41702, n41703, n41704,
         n41705, n41706, n41707, n41708, n41709, n41710, n41711, n41712,
         n41713, n41714, n41715, n41716, n41717, n41718, n41719, n41720,
         n41721, n41722, n41723, n41724, n41725, n41726, n41727, n41728,
         n41729, n41730, n41731, n41732, n41733, n41734, n41735, n41736,
         n41737, n41738, n41739, n41740, n41741, n41742, n41743, n41744,
         n41745, n41746, n41747, n41748, n41749, n41750, n41751, n41752,
         n41753, n41754, n41755, n41756, n41757, n41758, n41759, n41760,
         n41761, n41762, n41763, n41764, n41765, n41766, n41767, n41768,
         n41769, n41770, n41771, n41772, n41773, n41774, n41775, n41776,
         n41777, n41778, n41779, n41780, n41781, n41782, n41783, n41784,
         n41785, n41786, n41787, n41788, n41789, n41790, n41791, n41792,
         n41793, n41794, n41795, n41796, n41797, n41798, n41799, n41800,
         n41801, n41802, n41803, n41804, n41805, n41806, n41807, n41808,
         n41809, n41810, n41811, n41812, n41813, n41814, n41815, n41816,
         n41817, n41818, n41819, n41820, n41821, n41822, n41823, n41824,
         n41825, n41826, n41827, n41828, n41829, n41830, n41831, n41832,
         n41833, n41834, n41835, n41836, n41837, n41838, n41839, n41840,
         n41841, n41842, n41843, n41844, n41845, n41846, n41847, n41848,
         n41849, n41850, n41851, n41852, n41853, n41854, n41855, n41856,
         n41857, n41858, n41859, n41860, n41861, n41862, n41863, n41864,
         n41865, n41866, n41867, n41868, n41869, n41870, n41871, n41872,
         n41873, n41874, n41875, n41876, n41877, n41878, n41879, n41880,
         n41881, n41882, n41883, n41884, n41885, n41886, n41887, n41888,
         n41889, n41890, n41891, n41892, n41893, n41894, n41895, n41896,
         n41897, n41898, n41899, n41900, n41901, n41902, n41903, n41904,
         n41905, n41906, n41907, n41908, n41909, n41910, n41911, n41912,
         n41913, n41914, n41915, n41916, n41917, n41918, n41919, n41920,
         n41921, n41922, n41923, n41924, n41925, n41926, n41927, n41928,
         n41929, n41930, n41931, n41932, n41933, n41934, n41935, n41936,
         n41937, n41938, n41939, n41940, n41941, n41942, n41943, n41944,
         n41945, n41946, n41947, n41948, n41949, n41950, n41951, n41952,
         n41953, n41954, n41955, n41956, n41957, n41958, n41959, n41960,
         n41961, n41962, n41963, n41964, n41965, n41966, n41967, n41968,
         n41969, n41970, n41971, n41972, n41973, n41974, n41975, n41976,
         n41977, n41978, n41979, n41980, n41981, n41982, n41983, n41984,
         n41985, n41986, n41987, n41988, n41989, n41990, n41991, n41992,
         n41993, n41994, n41995, n41996, n41997, n41998, n41999, n42000,
         n42001, n42002, n42003, n42004, n42005, n42006, n42007, n42008,
         n42009, n42010, n42011, n42012, n42013, n42014, n42015, n42016,
         n42017, n42018, n42019, n42020, n42021, n42022, n42023, n42024,
         n42025, n42026, n42027, n42028, n42029, n42030, n42031, n42032,
         n42033, n42034, n42035, n42036, n42037, n42038, n42039, n42040,
         n42041, n42042, n42043, n42044, n42045, n42046, n42047, n42048,
         n42049, n42050, n42051, n42052, n42053, n42054, n42055, n42056,
         n42057, n42058, n42059, n42060, n42061, n42062, n42063, n42064,
         n42065, n42066, n42067, n42068, n42069, n42070, n42071, n42072,
         n42073, n42074, n42075, n42076, n42077, n42078, n42079, n42080,
         n42081, n42082, n42083, n42084, n42085, n42086, n42087, n42088,
         n42089, n42090, n42091, n42092, n42093, n42094, n42095, n42096,
         n42097, n42098, n42099, n42100, n42101, n42102, n42103, n42104,
         n42105, n42106, n42107, n42108, n42109, n42110, n42111, n42112,
         n42113, n42114, n42115, n42116, n42117, n42118, n42119, n42120,
         n42121, n42122, n42123, n42124, n42125, n42126, n42127, n42128,
         n42129, n42130, n42131, n42132, n42133, n42134, n42135, n42136,
         n42137, n42138, n42139, n42140, n42141, n42142, n42143, n42144,
         n42145, n42146, n42147, n42148, n42149, n42150, n42151, n42152,
         n42153, n42154, n42155, n42156, n42157, n42158, n42159, n42160,
         n42161, n42162, n42163, n42164, n42165, n42166, n42167, n42168,
         n42169, n42170, n42171, n42172, n42173, n42174, n42175, n42176,
         n42177, n42178, n42179, n42180, n42181, n42182, n42183, n42184,
         n42185, n42186, n42187, n42188, n42189, n42190, n42191, n42192,
         n42193, n42194, n42195, n42196, n42197, n42198, n42199, n42200,
         n42201, n42202, n42203, n42204, n42205, n42206, n42207, n42208,
         n42209, n42210, n42211, n42212, n42213, n42214, n42215, n42216,
         n42217, n42218, n42219, n42220, n42221, n42222, n42223, n42224,
         n42225, n42226, n42227, n42228, n42229, n42230, n42231, n42232,
         n42233, n42234, n42235, n42236, n42237, n42238, n42239, n42240,
         n42241, n42242, n42243, n42244, n42245, n42246, n42247, n42248,
         n42249, n42250, n42251, n42252, n42253, n42254, n42255, n42256,
         n42257, n42258, n42259, n42260, n42261, n42262, n42263, n42264,
         n42265, n42266, n42267, n42268, n42269, n42270, n42271, n42272,
         n42273, n42274, n42275, n42276, n42277, n42278, n42279, n42280,
         n42281, n42282, n42283, n42284, n42285, n42286, n42287, n42288,
         n42289, n42290, n42291, n42292, n42293, n42294, n42295, n42296,
         n42297, n42298, n42299, n42300, n42301, n42302, n42303, n42304,
         n42305, n42306, n42307, n42308, n42309, n42310, n42311, n42312,
         n42313, n42314, n42315, n42316, n42317, n42318, n42319, n42320,
         n42321, n42322, n42323, n42324, n42325, n42326, n42327, n42328,
         n42329, n42330, n42331, n42332, n42333, n42334, n42335, n42336,
         n42337, n42338, n42339, n42340, n42341, n42342, n42343, n42344,
         n42345, n42346, n42347, n42348, n42349, n42350, n42351, n42352,
         n42353, n42354, n42355, n42356, n42357, n42358, n42359, n42360,
         n42361, n42362, n42363, n42364, n42365, n42366, n42367, n42368,
         n42369, n42370, n42371, n42372, n42373, n42374, n42375, n42376,
         n42377, n42378, n42379, n42380, n42381, n42382, n42383, n42384,
         n42385, n42386, n42387, n42388, n44964, n44965, n44966, n44967,
         n44968, n44969, n44970, n44971, n44972, n44973, n44974, n44975,
         n44976, n44977, n44978, n44979, n44980, n44981, n44982, n44983,
         n44984, n44985, n44986, n44987, n44988, n44989, n44990, n44991,
         n44992, n44993, n44994, n44995, n44996, n44997, n44998, n44999,
         n45000, n45001, n45002, n45003, n45004, n45005, n45006, n45007,
         n45008, n45009, n45010, n45011, n45012, n45013, n45014, n45015,
         n45016, n45017, n45018, n45019, n45020, n45021, n45022, n45023,
         n45024, n45025, n45026, n45027, n45028, n45029, n45030, n45031,
         n45032, n45033, n45034, n45035, n45036, n45037, n45038, n45039,
         n45040, n45041, n45042, n45043, n45044, n45045, n45046, n45047,
         n45048, n45049, n45050, n45051, n45052, n45053, n45054, n45055,
         n45056, n45057, n45058, n45059, n45060, n45061, n45062, n45063,
         n45064, n45065, n45066, n45067, n45068, n45069, n45070, n45071,
         n45072, n45073, n45074, n45075, n45076, n45077, n45078, n45079,
         n45080, n45081, n45082, n45083, n45084, n45085, n45086, n45087,
         n45088, n45089, n45090, n45091, n45092, n45093, n45094, n45095,
         n45096, n45097, n45098, n45099, n45100, n45101, n45102, n45103,
         n45104, n45105, n45106, n45107, n45108, n45109, n45110, n45111,
         n45112, n45113, n45114, n45115, n45116, n45117, n45118, n45119,
         n45120, n45121, n45122, n45123, n45124, n45125, n45126, n45127,
         n45128, n45129, n45130, n45131, n45132, n45133, n45134, n45135,
         n45136, n45137, n45138, n45139, n45140, n45141, n45142, n45143,
         n45144, n45145, n45146, n45147, n45148, n45149, n45150, n45151,
         n45152, n45153, n45154, n45155, n45156, n45157, n45158, n45159,
         n45160, n45161, n45162, n45163, n45164, n45165, n45166, n45167,
         n45168, n45169, n45170, n45171, n45172, n45173, n45174, n45175,
         n45176, n45177, n45178, n45179, n45180, n45181, n45182, n45183,
         n45184, n45185, n45186, n45187, n45188, n45189, n45190, n45191,
         n45192, n45193, n45194, n45195, n45196, n45197, n45198, n45199,
         n45200, n45201, n45202, n45203, n45204, n45205, n45206, n45207,
         n45208, n45209, n45210, n45211, n45212, n45213, n45214, n45215,
         n45216, n45217, n45218, n45219, n45220, n45221, n45222, n45223,
         n45224, n45225, n45226, n45227, n45228, n45229, n45230, n45231,
         n45232, n45233, n45234, n45235, n45236, n45237, n45238, n45239,
         n45240, n45241, n45242, n45243, n45244, n45245, n45246, n45247,
         n45248, n45249, n45250, n45251, n45252, n45253, n45254, n45255,
         n45256, n45257, n45258, n45259, n45260, n45261, n45262, n45263,
         n45264, n45265, n45266, n45267, n45268, n45269, n45270, n45271,
         n45272, n45273, n45274, n45275, n45276, n45277, n45278, n45279,
         n45280, n45281, n45282, n45283, n45284, n45285, n45286, n45287,
         n45288, n45289, n45290, n45291, n45292, n45293, n45294, n45295,
         n45296, n45297, n45298, n45299, n45300, n45301, n45302, n45303,
         n45304, n45305, n45306, n45307, n45308, n45309, n45310, n45311,
         n45312, n45313, n45314, n45315, n45316, n45317, n45318, n45319,
         n45320, n45321, n45322, n45323, n45324, n45325, n45326, n45327,
         n45328, n45329, n45330, n45331, n45332, n45333, n45334, n45335,
         n45336, n45337, n45338, n45339, n45340, n45341, n45342, n45343,
         n45344, n45345, n45346, n45347, n45348, n45349, n45350, n45351,
         n45352, n45353, n45354, n45355, n45356, n45357, n45358, n45359,
         n45360, n45361, n45362, n45363, n45364, n45365, n45366, n45367,
         n45368, n45369, n45370, n45371, n45372, n45373, n45374, n45375,
         n45376, n45377, n45378, n45379, n45380, n45381, n45382, n45383,
         n45384, n45385, n45386, n45387, n45388, n45389, n45390, n45391,
         n45392, n45393, n45394, n45395, n45396, n45397, n45398, n45399,
         n45400, n45401, n45402, n45403, n45404, n45405, n45406, n45407,
         n45408, n45409, n45410, n45411, n45412, n45413, n45414, n45415,
         n45416, n45417, n45418, n45419, n45420, n45421, n45422, n45423,
         n45424, n45425, n45426, n45427, n45428, n45429, n45430, n45431,
         n45432, n45433, n45434, n45435, n45436, n45437, n45438, n45439,
         n45440, n45441, n45442, n45443, n45444, n45445, n45446, n45447,
         n45448, n45449, n45450, n45451, n45452, n45453, n45454, n45455,
         n45456, n45457, n45458, n45459, n45460, n45461, n45462, n45463,
         n45464, n45465, n45466, n45467, n45468, n45469, n45470, n45471,
         n45472, n45473, n45474, n45475, n45476, n45477, n45478, n45479,
         n45480, n45481, n45482, n45483, n45484, n45485, n45486, n45487,
         n45488, n45489, n45490, n45491, n45492, n45493, n45494, n45495,
         n45496, n45497, n45498, n45499, n45500, n45501, n45502, n45503,
         n45504, n45505, n45506, n45507, n45508, n45509, n45510, n45511,
         n45512, n45513, n45514, n45515, n45516, n45517, n45518, n45519,
         n45520, n45521, n45522, n45523, n45524, n45525, n45526, n45527,
         n45528, n45529, n45530, n45531, n45532, n45533, n45534, n45535,
         n45536, n45537, n45538, n45539, n45540, n45541, n45542, n45543,
         n45544, n45545, n45546, n45547, n45548, n45549, n45550, n45551,
         n45552, n45553, n45554, n45555, n45556, n45557, n45558, n45559,
         n45560, n45561, n45562, n45563, n45564, n45565, n45566, n45567,
         n45568, n45569, n45570, n45571, n45572, n45573, n45574, n45575,
         n45576, n45577, n45578, n45579, n45580, n45581, n45582, n45583,
         n45584, n45585, n45586, n45587, n45588, n45589, n45590, n45591,
         n45592, n45593, n45594, n45595, n45596, n45597, n45598, n45599,
         n45600, n45601, n45602, n45603, n45604, n45605, n45606, n45607,
         n45608, n45609, n45610, n45611, n45612, n45613, n45614, n45615,
         n45616, n45617, n45618, n45619, n45620, n45621, n45622, n45623,
         n45624, n45625, n45626, n45627, n45628, n45629, n45630, n45631,
         n45632, n45633, n45634, n45635, n45636, n45637, n45638, n45639,
         n45640, n45641, n45642, n45643, n45644, n45645, n45646, n45647,
         n45648, n45649, n45650, n45651, n45652, n45653, n45654, n45655,
         n45656, n45657, n45658, n45659, n45660, n45661, n45662, n45663,
         n45664, n45665, n45666, n45667, n45668, n45669, n45670, n45671,
         n45672, n45673, n45674, n45675, n45676, n45677, n45678, n45679,
         n45680, n45681, n45682, n45683, n45684, n45685, n45686, n45687,
         n45688, n45689, n45690, n45691, n45692, n45693, n45694, n45695,
         n45696, n45697, n45698, n45699, n45700, n45701, n45702, n45703,
         n45704, n45705, n45706, n45707, n45708, n45709, n45710, n45711,
         n45712, n45713, n45714, n45715, n45716, n45717, n45718, n45719,
         n45720, n45721, n45722, n45723, n45724, n45725, n45726, n45727,
         n45728, n45729, n45730, n45731, n45732, n45733, n45734, n45735,
         n45736, n45737, n45738, n45739, n45740, n45741, n45742, n45743,
         n45744, n45745, n45746, n45747, n45748, n45749, n45750, n45751,
         n45752, n45753, n45754, n45755, n45756, n45757, n45758, n45759,
         n45760, n45761, n45762, n45763, n45764, n45765, n45766, n45767,
         n45768, n45769, n45770, n45771, n45772, n45773, n45774, n45775,
         n45776, n45777, n45778, n45779, n45780, n45781, n45782, n45783,
         n45784, n45785, n45786, n45787, n45788, n45789, n45790, n45791,
         n45792, n45793, n45794, n45795, n45796, n45797, n45798, n45799,
         n45800, n45801, n45802, n45803, n45804, n45805, n45806, n45807,
         n45808, n45809, n45810, n45811, n45812, n45813, n45814, n45815,
         n45816, n45817, n45818, n45819, n45820, n45821, n45822, n45823,
         n45824, n45825, n45826, n45827, n45828, n45829, n45830, n45831,
         n45832, n45833, n45834, n45835, n45836, n45837, n45838, n45839,
         n45840, n45841, n45842, n45843, n45844, n45845, n45846, n45847,
         n45848, n45849, n45850, n45851, n45852, n45853, n45854, n45855,
         n45856, n45857, n45858, n45859, n45860, n45861, n45862, n45863,
         n45864, n45865, n45866, n45867, n45868, n45869, n45870, n45871,
         n45872, n45873, n45874, n45875, n45876, n45877, n45878, n45879,
         n45880, n45881, n45882, n45883, n45884, n45885, n45886, n45887,
         n45888, n45889, n45890, n45891, n45892, n45893, n45894, n45895,
         n45896, n45897, n45898, n45899, n45900, n45901, n45902, n45903,
         n45904, n45905, n45906, n45907, n45908, n45909, n45910, n45911,
         n45912, n45913, n45914, n45915, n45916, n45917, n45918, n45919,
         n45920, n45921, n45922, n45923, n45924, n45925, n45926, n45927,
         n45928, n45929, n45930, n45931, n45932, n45933, n45934, n45935,
         n45936, n45937, n45938, n45939, n45940, n45941, n45942, n45943,
         n45944, n45945, n45946, n45947, n45948, n45949, n45950, n45951,
         n45952, n45953, n45954, n45955, n45956, n45957, n45958, n45959,
         n45960, n45961, n45962, n45963, n45964, n45965, n45966, n45967,
         n45968, n45969, n45970, n45971, n45972, n45973, n45974, n45975,
         n45976, n45977, n45978, n45979, n45980, n45981, n45982, n45983,
         n45984, n45985, n45986, n45987, n45988, n45989, n45990, n45991,
         n45992, n45993, n45994, n45995, n45996, n45997, n45998, n45999,
         n46000, n46001, n46002, n46003, n46004, n46005, n46006, n46007,
         n46008, n46009, n46010, n46011, n46012, n46013, n46014, n46015,
         n46016, n46017, n46018, n46019, n46020, n46021, n46022, n46023,
         n46024, n46025, n46026, n46027, n46028, n46029, n46030, n46031,
         n46032, n46033, n46034, n46035, n46036, n46037, n46038, n46039,
         n46040, n46041, n46042, n46043, n46044, n46045, n46046, n46047,
         n46048, n46049, n46050, n46051, n46052, n46053, n46054, n46055,
         n46056, n46057, n46058, n46059, n46060, n46061, n46062, n46063,
         n46064, n46065, n46066, n46067, n46068, n46069, n46070, n46071,
         n46072, n46073, n46074, n46075, n46076, n46077, n46078, n46079,
         n46080, n46081, n46082, n46083, n46084, n46085, n46086, n46087,
         n46088, n46089, n46090, n46091, n46092, n46093, n46094, n46095,
         n46096, n46097, n46098, n46099, n46100, n46101, n46102, n46103,
         n46104, n46105, n46106, n46107, n46108, n46109, n46110, n46111,
         n46112, n46113, n46114, n46115, n46116, n46117, n46118, n46119,
         n46120, n46121, n46122, n46123, n46124, n46125, n46126, n46127,
         n46128, n46129, n46130, n46131, n46132, n46133, n46134, n46135,
         n46136, n46137, n46138, n46139, n46140, n46141, n46142, n46143,
         n46144, n46145, n46146, n46147, n46148, n46149, n46150, n46151,
         n46152, n46153, n46154, n46155, n46156, n46157, n46158, n46159,
         n46160, n46161, n46162, n46163, n46164, n46165, n46166, n46167,
         n46168, n46169, n46170, n46171, n46172, n46173, n46174, n46175,
         n46176, n46177, n46178, n46179, n46180, n46181, n46182, n46183,
         n46184, n46185, n46186, n46187, n46188, n46189, n46190, n46191,
         n46192, n46193, n46194, n46195, n46196, n46197, n46198, n46199,
         n46200, n46201, n46202, n46203, n46204, n46205, n46206, n46207,
         n46208, n46209, n46210, n46211, n46212, n46213, n46214, n46215,
         n46216, n46217, n46218, n46219, n46220, n46221, n46222, n46223,
         n46224, n46225, n46226, n46227, n46228, n46229, n46230, n46231,
         n46232, n46233, n46234, n46235, n46236, n46237, n46238, n46239,
         n46240, n46241, n46242, n46243, n46244, n46245, n46246, n46247,
         n46248, n46249, n46250, n46251, n46252, n46253, n46254, n46255,
         n46256, n46257, n46258, n46259, n46260, n46261, n46262, n46263,
         n46264, n46265, n46266, n46267, n46268, n46269, n46270, n46271,
         n46272, n46273, n46274, n46275, n46276, n46277, n46278, n46279,
         n46280, n46281, n46282, n46283, n46284, n46285, n46286, n46287,
         n46288, n46289, n46290, n46291, n46292, n46293, n46294, n46295,
         n46296, n46297, n46298, n46299, n46300, n46301, n46302, n46303,
         n46304, n46305, n46306, n46307, n46308, n46309, n46310, n46311,
         n46312, n46313, n46314, n46315, n46316, n46317, n46318, n46319,
         n46320, n46321, n46322, n46323, n46324, n46325, n46326, n46327,
         n46328, n46329, n46330, n46331, n46332, n46333, n46334, n46335,
         n46336, n46337, n46338, n46339, n46340, n46341, n46342, n46343,
         n46344, n46345, n46346, n46347, n46348, n46349, n46350, n46351,
         n46352, n46353, n46354, n46355, n46356, n46357, n46358, n46359,
         n46360, n46361, n46362, n46363, n46364, n46365, n46366, n46367,
         n46368, n46369, n46370, n46371, n46372, n46373, n46374, n46375,
         n46376, n46377, n46378, n46379, n46380, n46381, n46382, n46383,
         n46384, n46385, n46386, n46387, n46388, n46389, n46390, n46391,
         n46392, n46393, n46394, n46395, n46396, n46397, n46398, n46399,
         n46400, n46401, n46402, n46403, n46404, n46405, n46406, n46407,
         n46408, n46409, n46410, n46411, n46412, n46413, n46414, n46415,
         n46416, n46417, n46418, n46419, n46420, n46421, n46422, n46423,
         n46424, n46425, n46426, n46427, n46428, n46429, n46430, n46431,
         n46432, n46433, n46434, n46435, n46436, n46437, n46438, n46439,
         n46440, n46441, n46442, n46443, n46444, n46445, n46446, n46447,
         n46448, n46449, n46450, n46451, n46452, n46453, n46454, n46455,
         n46456, n46457, n46458, n46459, n46460, n46461, n46462, n46463,
         n46464, n46465, n46466, n46467, n46468, n46469, n46470, n46471,
         n46472, n46473, n46474, n46475, n46476, n46477, n46478, n46479,
         n46480, n46481, n46482, n46483, n46484, n46485, n46486, n46487,
         n46488, n46489, n46490, n46491, n46492, n46493, n46494, n46495,
         n46496, n46497, n46498, n46499, n46500, n46501, n46502, n46503,
         n46504, n46505, n46506, n46507, n46508, n46509, n46510, n46511,
         n46512, n46513, n46514, n46515, n46516, n46517, n46518, n46519,
         n46520, n46521, n46522, n46523, n46524, n46525, n46526, n46527,
         n46528, n46529, n46530, n46531, n46532, n46533, n46534, n46535,
         n46536, n46537, n46538, n46539, n46540, n46541, n46542, n46543,
         n46544, n46545, n46546, n46547, n46548, n46549, n46550, n46551,
         n46552, n46553, n46554, n46555, n46556, n46557, n46558, n46559,
         n46560, n46561, n46562, n46563, n46564, n46565, n46566, n46567,
         n46568, n46569, n46570, n46571, n46572, n46573, n46574, n46575,
         n46576, n46577, n46578, n46579, n46580, n46581, n46582, n46583,
         n46584, n46585, n46586, n46587, n46588, n46589, n46590, n46591,
         n46592, n46593, n46594, n46595, n46596, n46597, n46598, n46599,
         n46600, n46601, n46602, n46603, n46604, n46605, n46606, n46607,
         n46608, n46609, n46610, n46611, n46612, n46613, n46614, n46615,
         n46616, n46617, n46618, n46619, n46620, n46621, n46622, n46623,
         n46624, n46625, n46626, n46627, n46628, n46629, n46630, n46631,
         n46632, n46633, n46634, n46635, n46636, n46637, n46638, n46639,
         n46640, n46641, n46642, n46643, n46644, n46645, n46646, n46647,
         n46648, n46649, n46650, n46651, n46652, n46653, n46654, n46655,
         n46656, n46657, n46658, n46659, n46660, n46661, n46662, n46663,
         n46664, n46665, n46666, n46667, n46668, n46669, n46670, n46671,
         n46672, n46673, n46674, n46675, n46676, n46677, n46678, n46679,
         n46680, n46681, n46682, n46683, n46684, n46685, n46686, n46687,
         n46688, n46689, n46690, n46691, n46692, n46693, n46694, n46695,
         n46696, n46697, n46698, n46699, n46700, n46701, n46702, n46703,
         n46704, n46705, n46706, n46707, n46708, n46709, n46710, n46711,
         n46712, n46713, n46714, n46715, n46716, n46717, n46718, n46719,
         n46720, n46721, n46722, n46723, n46724, n46725, n46726, n46727,
         n46728, n46729, n46730, n46731, n46732, n46733, n46734, n46735,
         n46736, n46737, n46738, n46739, n46740, n46741, n46742, n46743,
         n46744, n46745, n46746, n46747, n46748, n46749, n46750, n46751,
         n46752, n46753, n46754, n46755, n46756, n46757, n46758, n46759,
         n46760, n46761, n46762, n46763, n46764, n46765, n46766, n46767,
         n46768, n46769, n46770, n46771, n46772, n46773, n46774, n46775,
         n46776, n46777, n46778, n46779, n46780, n46781, n46782, n46783,
         n46784, n46785, n46786, n46787, n46788, n46789, n46790, n46791,
         n46792, n46793, n46794, n46795, n46796, n46797, n46798, n46799,
         n46800, n46801, n46802, n46803, n46804, n46805, n46806, n46807,
         n46808, n46809, n46810, n46811, n46812, n46813, n46814, n46815,
         n46816, n46817, n46818, n46819, n46820, n46821, n46822, n46823,
         n46824, n46825, n46826, n46827, n46828, n46829, n46830, n46831,
         n46832, n46833, n46834, n46835, n46836, n46837, n46838, n46839,
         n46840, n46841, n46842, n46843, n46844, n46845, n46846, n46847,
         n46848, n46849, n46850, n46851, n46852, n46853, n46854, n46855,
         n46856, n46857, n46858, n46859, n46860, n46861, n46862, n46863,
         n46864, n46865, n46866, n46867, n46868, n46869, n46870, n46871,
         n46872, n46873, n46874, n46875, n46876, n46877, n46878, n46879,
         n46880, n46881, n46882, n46883, n46884, n46885, n46886, n46887,
         n46888, n46889, n46890, n46891, n46892, n46893, n46894, n46895,
         n46896, n46897, n46898, n46899, n46900, n46901, n46902, n46903,
         n46904, n46905, n46906, n46907, n46908, n46909, n46910, n46911,
         n46912, n46913, n46914, n46915, n46916, n46917, n46918, n46919,
         n46920, n46921, n46922, n46923, n46924, n46925, n46926, n46927,
         n46928, n46929, n46930, n46931, n46932, n46933, n46934, n46935,
         n46936, n46937, n46938, n46939, n46940, n46941, n46942, n46943,
         n46944, n46945, n46946, n46947, n46948, n46949, n46950, n46951,
         n46952, n46953, n46954, n46955, n46956, n46957, n46958, n46959,
         n46960, n46961, n46962, n46963, n46964, n46965, n46966, n46967,
         n46968, n46969, n46970, n46971, n46972, n46973, n46974, n46975,
         n46976, n46977, n46978, n46979, n46980, n46981, n46982, n46983,
         n46984, n46985, n46986, n46987, n46988, n46989, n46990, n46991,
         n46992, n46993, n46994, n46995, n46996, n46997, n46998, n46999,
         n47000, n47001, n47002, n47003, n47004, n47005, n47006, n47007,
         n47008, n47009, n47010, n47011, n47012, n47013, n47014, n47015,
         n47016, n47017, n47018, n47019, n47020, n47021, n47022, n47023,
         n47024, n47025, n47026, n47027, n47028, n47029, n47030, n47031,
         n47032, n47033, n47034, n47035, n47036, n47037, n47038, n47039,
         n47040, n47041, n47042, n47043, n47044, n47045, n47046, n47047,
         n47048, n47049, n47050, n47051, n47052, n47053, n47054, n47055,
         n47056, n47057, n47058, n47059, n47060, n47061, n47062, n47063,
         n47064, n47065, n47066, n47067, n47068, n47069, n47070, n47071,
         n47072, n47073, n47074, n47075, n47076, n47077, n47078, n47079,
         n47080, n47081, n47082, n47083, n47084, n47085, n47086, n47087,
         n47088, n47089, n47090, n47091, n47092, n47093, n47094, n47095,
         n47096, n47097, n47098, n47099, n47100, n47101, n47102, n47103,
         n47104, n47105, n47106, n47107, n47108, n47109, n47110, n47111,
         n47112, n47113, n47114, n47115, n47116, n47117, n47118, n47119,
         n47120, n47121, n47122, n47123, n47124, n47125, n47126, n47127,
         n47128, n47129, n47130, n47131, n47132, n47133, n47134, n47135,
         n47136, n47137, n47138, n47139, n47140, n47141, n47142, n47143,
         n47144, n47145, n47146, n47147, n47148, n47149, n47150, n47151,
         n47152, n47153, n47154, n47155, n47156, n47157, n47158, n47159,
         n47160, n47161, n47162, n47163, n47164, n47165, n47166, n47167,
         n47168, n47169, n47170, n47171, n47172, n47173, n47174, n47175,
         n47176, n47177, n47178, n47179, n47180, n47181, n47182, n47183,
         n47184, n47185, n47186, n47187, n47188, n47189, n47190, n47191,
         n47192, n47193, n47194, n47195, n47196, n47197, n47198, n47199,
         n47200, n47201, n47202, n47203, n47204, n47205, n47206, n47207,
         n47208, n47209, n47210, n47211, n47212, n47213, n47214, n47215,
         n47216, n47217, n47218, n47219, n47220, n47221, n47222, n47223,
         n47224, n47225, n47226, n47227, n47228, n47229, n47230, n47231,
         n47232, n47233, n47234, n47235, n47236, n47237, n47238, n47239,
         n47240, n47241, n47242, n47243, n47244, n47245, n47246, n47247,
         n47248, n47249, n47250, n47251, n47252, n47253, n47254, n47255,
         n47256, n47257, n47258, n47259, n47260, n47261, n47262, n47263,
         n47264, n47265, n47266, n47267, n47268, n47269, n47270, n47271,
         n47272, n47273, n47274, n47275, n47276, n47277, n47278, n47279,
         n47280, n47281, n47282, n47283, n47284, n47285, n47286, n47287,
         n47288, n47289, n47290, n47291, n47292, n47293, n47294, n47295,
         n47296, n47297, n47298, n47299, n47300, n47301, n47302, n47303,
         n47304, n47305, n47306, n47307, n47308, n47309, n47310, n47311,
         n47312, n47313, n47314, n47315, n47316, n47317, n47318, n47319,
         n47320, n47321, n47322, n47323, n47324, n47325, n47326, n47327,
         n47328, n47329, n47330, n47331, n47332, n47333, n47334, n47335,
         n47336, n47337, n47338, n47339, n47340, n47341, n47342, n47343,
         n47344, n47345, n47346, n47347, n47348, n47349, n47350, n47351,
         n47352, n47353, n47354, n47355, n47356, n47357, n47358, n47359,
         n47360, n47361, n47362, n47363, n47364, n47365, n47366, n47367,
         n47368, n47369, n47370, n47371, n47372, n47373, n47374, n47375,
         n47376, n47377, n47378, n47379, n47380, n47381, n47382, n47383,
         n47384, n47385, n47386, n47387, n47388, n47389, n47390, n47391,
         n47392, n47393, n47394, n47395, n47396, n47397, n47398, n47399,
         n47400, n47401, n47402, n47403, n47404, n47405, n47406, n47407,
         n47408, n47409, n47410, n47411, n47412, n47413, n47414, n47415,
         n47416, n47417, n47418, n47419, n47420, n47421, n47422, n47423,
         n47424, n47425, n47426, n47427, n47428, n47429, n47430, n47431,
         n47432, n47433, n47434, n47435, n47436, n47437, n47438, n47439,
         n47440, n47441, n47442, n47443, n47444, n47445, n47446, n47447,
         n47448, n47449, n47450, n47451, n47452, n47453, n47454, n47455,
         n47456, n47457, n47458, n47459, n47460, n47461, n47462, n47463,
         n47464, n47465, n47466, n47467, n47468, n47469, n47470, n47471,
         n47472, n47473, n47474, n47475, n47476, n47477, n47478, n47479,
         n47480, n47481, n47482, n47483, n47484, n47485, n47486, n47487,
         n47488, n47489, n47490, n47491, n47492, n47493, n47494, n47495,
         n47496, n47497, n47498, n47499, n47500, n47501, n47502, n47503,
         n47504, n47505, n47506, n47507, n47508, n47509, n47510, n47511,
         n47512, n47513, n47514, n47515, n47516, n47517, n47518, n47519,
         n47520, n47521, n47522, n47523, n47524, n47525, n47526, n47527,
         n47528, n47529, n47530, n47531, n47532, n47533, n47534, n47535,
         n47536, n47537, n47538, n47539, n47540, n47541, n47542, n47543,
         n47544, n47545, n47546, n47547, n47548, n47549, n47550, n47551,
         n47552, n47553, n47554, n47555, n47556, n47557, n47558, n47559,
         n47560, n47561, n47562, n47563, n47564, n47565, n47566, n47567,
         n47568, n47569, n47570, n47571, n47572, n47573, n47574, n47575,
         n47576, n47577, n47578, n47579, n47580, n47581, n47582, n47583,
         n47584, n47585, n47586, n47587, n47588, n47589, n47590, n47591,
         n47592, n47593, n47594, n47595, n47596, n47597, n47598, n47599,
         n47600, n47601, n47602, n47603, n47604, n47605, n47606, n47607,
         n47608, n47609, n47610, n47611, n47612, n47613, n47614, n47615,
         n47616, n47617, n47618, n47619, n47620, n47621, n47622, n47623,
         n47624, n47625, n47626, n47627, n47628, n47629, n47630, n47631,
         n47632, n47633, n47634, n47635, n47636, n47637, n47638, n47639,
         n47640, n47641, n47642, n47643, n47644, n47645, n47646, n47647,
         n47648, n47649, n47650, n47651, n47652, n47653, n47654, n47655,
         n47656, n47657, n47658, n47659, n47660, n47661, n47662, n47663,
         n47664, n47665, n47666, n47667, n47668, n47669, n47670, n47671,
         n47672, n47673, n47674, n47675, n47676, n47677, n47678, n47679,
         n47680, n47681, n47682, n47683, n47684, n47685, n47686, n47687,
         n47688, n47689, n47690, n47691, n47692, n47693, n47694, n47695,
         n47696, n47697, n47698, n47699, n47700, n47701, n47702, n47703,
         n47704, n47705, n47706, n47707, n47708, n47709, n47710, n47711,
         n47712, n47713, n47714, n47715, n47716, n47717, n47718, n47719,
         n47720, n47721, n47722, n47723, n47724, n47725, n47726, n47727,
         n47728, n47729, n47730, n47731, n47732, n47733, n47734, n47735,
         n47736, n47737, n47738, n47739, n47740, n47741, n47742, n47743,
         n47744, n47745, n47746, n47747, n47748, n47749, n47750, n47751,
         n47752, n47753, n47754, n47755, n47756, n47757, n47758, n47759,
         n47760, n47761, n47762, n47763, n47764, n47765, n47766, n47767,
         n47768, n47769, n47770, n47771, n47772, n47773, n47774, n47775,
         n47776, n47777, n47778, n47779, n47780, n47781, n47782, n47783,
         n47784, n47785, n47786, n47787, n47788, n47789, n47790, n47791,
         n47792, n47793, n47794, n47795, n47796, n47797, n47798, n47799,
         n47800, n47801, n47802, n47803, n47804, n47805, n47806, n47807,
         n47808, n47809, n47810, n47811, n47812, n47813, n47814, n47815,
         n47816, n47817, n47818, n47819, n47820, n47821, n47822, n47823,
         n47824, n47825, n47826, n47827, n47828, n47829, n47830, n47831,
         n47832, n47833, n47834, n47835, n47836, n47837, n47838, n47839,
         n47840, n47841, n47842, n47843, n47844, n47845, n47846, n47847,
         n47848, n47849, n47850, n47851, n47852, n47853, n47854, n47855,
         n47856, n47857, n47858, n47859, n47860, n47861, n47862, n47863,
         n47864, n47865, n47866, n47867, n47868, n47869, n47870, n47871,
         n47872, n47873, n47874, n47875, n47876, n47877, n47878, n47879,
         n47880, n47881, n47882, n47883, n47884, n47885, n47886, n47887,
         n47888, n47889, n47890, n47891, n47892, n47893, n47894, n47895,
         n47896, n47897, n47898, n47899, n47900, n47901, n47902, n47903,
         n47904, n47905, n47906, n47907, n47908, n47909, n47910, n47911,
         n47912, n47913, n47914, n47915, n47916, n47917, n47918, n47919,
         n47920, n47921, n47922, n47923, n47924, n47925, n47926, n47927,
         n47928, n47929, n47930, n47931, n47932, n47933, n47934, n47935,
         n47936, n47937, n47938, n47939, n47940, n47941, n47942, n47943,
         n47944, n47945, n47946, n47947, n47948, n47949, n47950, n47951,
         n47952, n47953, n47954, n47955, n47956, n47957, n47958, n47959,
         n47960, n47961, n47962, n47963, n47964, n47965, n47966, n47967,
         n47968, n47969, n47970, n47971, n47972, n47973, n47974, n47975,
         n47976, n47977, n47978, n47979, n47980, n47981, n47982, n47983,
         n47984, n47985, n47986, n47987, n47988, n47989, n47990, n47991,
         n47992, n47993, n47994, n47995, n47996, n47997, n47998, n47999,
         n48000, n48001, n48002, n48003, n48004, n48005, n48006, n48007,
         n48008, n48009, n48010, n48011, n48012, n48013, n48014, n48015,
         n48016, n48017, n48018, n48019, n48020, n48021, n48022, n48023,
         n48024, n48025, n48026, n48027, n48028, n48029, n48030, n48031,
         n48032, n48033, n48034, n48035, n48036, n48037, n48038, n48039,
         n48040, n48041, n48042, n48043, n48044, n48045, n48046, n48047,
         n48048, n48049, n48050, n48051, n48052, n48053, n48054, n48055,
         n48056, n48057, n48058, n48059, n48060, n48061, n48062, n48063,
         n48064, n48065, n48066, n48067, n48068, n48069, n48070, n48071,
         n48072, n48073, n48074, n48075, n48076, n48077, n48078, n48079,
         n48080, n48081, n48082, n48083, n48084, n48085, n48086, n48087,
         n48088, n48089, n48090, n48091, n48092, n48093, n48094, n48095,
         n48096, n48097, n48098, n48099, n48100, n48101, n48102, n48103,
         n48104, n48105, n48106, n48107, n48108, n48109, n48110, n48111,
         n48112, n48113, n48114, n48115, n48116, n48117, n48118, n48119,
         n48120, n48121, n48122, n48123, n48124, n48125, n48126, n48127,
         n48128, n48129, n48130, n48131, n48132, n48133, n48134, n48135,
         n48136, n48137, n48138, n48139, n48140, n48141, n48142, n48143,
         n48144, n48145, n48146, n48147, n48148, n48149, n48150, n48151,
         n48152, n48153, n48154, n48155, n48156, n48157, n48158, n48159,
         n48160, n48161, n48162, n48163, n48164, n48165, n48166, n48167,
         n48168, n48169, n48170, n48171, n48172, n48173, n48174, n48175,
         n48176, n48177, n48178, n48179, n48180, n48181, n48182, n48183,
         n48184, n48185, n48186, n48187, n48188, n48189, n48190, n48191,
         n48192, n48193, n48194, n48195, n48196, n48197, n48198, n48199,
         n48200, n48201, n48202, n48203, n48204, n48205, n48206, n48207,
         n48208, n48209, n48210, n48211, n48212, n48213, n48214, n48215,
         n48216, n48217, n48218, n48219, n48220, n48221, n48222, n48223,
         n48224, n48225, n48226, n48227, n48228, n48229, n48230, n48231,
         n48232, n48233, n48234, n48235, n48236, n48237, n48238, n48239,
         n48240, n48241, n48242, n48243, n48244, n48245, n48246, n48247,
         n48248, n48249, n48250, n48251, n48252, n48253, n48254, n48255,
         n48256, n48257, n48258, n48259, n48260, n48261, n48262, n48263,
         n48264, n48265, n48266, n48267, n48268, n48269, n48270, n48271,
         n48272, n48273, n48274, n48275, n48276, n48277, n48278, n48279,
         n48280, n48281, n48282, n48283, n48284, n48285, n48286, n48287,
         n48288, n48289, n48290, n48291, n48292, n48293, n48294, n48295,
         n48296, n48297, n48298, n48299, n48300, n48301, n48302, n48303,
         n48304, n48305, n48306, n48307, n48308, n48309, n48310, n48311,
         n48312, n48313, n48314, n48315, n48316, n48317, n48318, n48319,
         n48320, n48321, n48322, n48323, n48324, n48325, n48326, n48327,
         n48328, n48329, n48330, n48331, n48332, n48333, n48334, n48335,
         n48336, n48337, n48338, n48339, n48340, n48341, n48342, n48343,
         n48344, n48345, n48346, n48347, n48348, n48349, n48350, n48351,
         n48352, n48353, n48354, n48355, n48356, n48357, n48358, n48359,
         n48360, n48361, n48362, n48363, n48364, n48365, n48366, n48367,
         n48368, n48369, n48370, n48371, n48372, n48373, n48374, n48375,
         n48376, n48377, n48378, n48379, n48380, n48381, n48382, n48383,
         n48384, n48385, n48386, n48387, n48388, n48389, n48390, n48391,
         n48392, n48393, n48394, n48395, n48396, n48397, n48398, n48399,
         n48400, n48401, n48402, n48403, n48404, n48405, n48406, n48407,
         n48408, n48409, n48410, n48411, n48412, n48413, n48414, n48415,
         n48416, n48417, n48418, n48419, n48420, n48421, n48422, n48423,
         n48424, n48425, n48426, n48427, n48428, n48429, n48430, n48431,
         n48432, n48433, n48434, n48435, n48436, n48437, n48438, n48439,
         n48440, n48441, n48442, n48443, n48444, n48445, n48446, n48447,
         n48448, n48449, n48450, n48451, n48452, n48453, n48454, n48455,
         n48456, n48457, n48458, n48459, n48460, n48461, n48462, n48463,
         n48464, n48465, n48466, n48467, n48468, n48469, n48470, n48471,
         n48472, n48473, n48474, n48475, n48476, n48477, n48478, n48479,
         n48480, n48481, n48482, n48483, n48484, n48485, n48486, n48487,
         n48488, n48489, n48490, n48491, n48492, n48493, n48494, n48495,
         n48496, n48497, n48498, n48499, n48500, n48501, n48502, n48503,
         n48504, n48505, n48506, n48507, n48508, n48509, n48510, n48511,
         n48512, n48513, n48514, n48515, n48516, n48517, n48518, n48519,
         n48520, n48521, n48522, n48523, n48524, n48525, n48526, n48527,
         n48528, n48529, n48530, n48531, n48532, n48533, n48534, n48535,
         n48536, n48537, n48538, n48539, n48540, n48541, n48542, n48543,
         n48544, n48545, n48546, n48547, n48548, n48549, n48550, n48551,
         n48552, n48553, n48554, n48555, n48556, n48557, n48558, n48559,
         n48560, n48561, n48562, n48563, n48564, n48565, n48566, n48567,
         n48568, n48569, n48570, n48571, n48572, n48573, n48574, n48575,
         n48576, n48577, n48578, n48579, n48580, n48581, n48582, n48583,
         n48584, n48585, n48586, n48587, n48588, n48589, n48590, n48591,
         n48592, n48593, n48594, n48595, n48596, n48597, n48598, n48599,
         n48600, n48601, n48602, n48603, n48604, n48605, n48606, n48607,
         n48608, n48609, n48610, n48611, n48612, n48613, n48614, n48615,
         n48616, n48617, n48618, n48619, n48620, n48621, n48622, n48623,
         n48624, n48625, n48626, n48627, n48628, n48629, n48630, n48631,
         n48632, n48633, n48634, n48635, n48636, n48637, n48638, n48639,
         n48640, n48641, n48642, n48643, n48644, n48645, n48646, n48647,
         n48648, n48649, n48650, n48651, n48652, n48653, n48654, n48655,
         n48656, n48657, n48658, n48659, n48660, n48661, n48662, n48663,
         n48664, n48665, n48666, n48667, n48668, n48669, n48670, n48671,
         n48672, n48673, n48674, n48675, n48676, n48677, n48678, n48679,
         n48680, n48681, n48682, n48683, n48684, n48685, n48686, n48687,
         n48688, n48689, n48690, n48691, n48692, n48693, n48694, n48695,
         n48696, n48697, n48698, n48699, n48700, n48701, n48702, n48703,
         n48704, n48705, n48706, n48707, n48708, n48709, n48710, n48711,
         n48712, n48713, n48714, n48715, n48716, n48717, n48718, n48719,
         n48720, n48721, n48722, n48723, n48724, n48725, n48726, n48727,
         n48728, n48729, n48730, n48731, n48732, n48733, n48734, n48735,
         n48736, n48737, n48738, n48739, n48740, n48741, n48742, n48743,
         n48744, n48745, n48746, n48747, n48748, n48749, n48750, n48751,
         n48752, n48753, n48754, n48755, n48756, n48757, n48758, n48759,
         n48760, n48761, n48762, n48763, n48764, n48765, n48766, n48767,
         n48768, n48769, n48770, n48771, n48772, n48773, n48774, n48775,
         n48776, n48777, n48778, n48779, n48780, n48781, n48782, n48783,
         n48784, n48785, n48786, n48787, n48788, n48789, n48790, n48791,
         n48792, n48793, n48794, n48795, n48796, n48797, n48798, n48799,
         n48800, n48801, n48802, n48803, n48804, n48805, n48806, n48807,
         n48808, n48809, n48810, n48811, n48812, n48813, n48814, n48815,
         n48816, n48817, n48818, n48819, n48820, n48821, n48822, n48823,
         n48824, n48825, n48826, n48827, n48828, n48829, n48830, n48831,
         n48832, n48833, n48834, n48835, n48836, n48837, n48838, n48839,
         n48840, n48841, n48842, n48843, n48844, n48845, n48846, n48847,
         n48848, n48849, n48850, n48851, n48852, n48853, n48854, n48855,
         n48856, n48857, n48858, n48859, n48860, n48861, n48862, n48863,
         n48864, n48865, n48866, n48867, n48868, n48869, n48870, n48871,
         n48872, n48873, n48874, n48875, n48876, n48877, n48878, n48879,
         n48880, n48881, n48882, n48883, n48884, n48885, n48886, n48887,
         n48888, n48889, n48890, n48891, n48892, n48893, n48894, n48895,
         n48896, n48897, n48898, n48899, n48900, n48901, n48902, n48903,
         n48904, n48905, n48906, n48907, n48908, n48909, n48910, n48911,
         n48912, n48913, n48914, n48915, n48916, n48917, n48918, n48919,
         n48920, n48921, n48922, n48923, n48924, n48925, n48926, n48927,
         n48928, n48929, n48930, n48931, n48932, n48933, n48934, n48935,
         n48936, n48937, n48938, n48939, n48940, n48941, n48942, n48943,
         n48944, n48945, n48946, n48947, n48948, n48949, n48950, n48951,
         n48952, n48953, n48954, n48955, n48956, n48957, n48958, n48959,
         n48960, n48961, n48962, n48963, n48964, n48965, n48966, n48967,
         n48968, n48969, n48970, n48971, n48972, n48973, n48974, n48975,
         n48976, n48977, n48978, n48979, n48980, n48981, n48982, n48983,
         n48984, n48985, n48986, n48987, n48988, n48989, n48990, n48991,
         n48992, n48993, n48994, n48995, n48996, n48997, n48998, n48999,
         n49000, n49001, n49002, n49003, n49004, n49005, n49006, n49007,
         n49008, n49009, n49010, n49011, n49012, n49013, n49014, n49015,
         n49016, n49017, n49018, n49019, n49020, n49021, n49022, n49023,
         n49024, n49025, n49026, n49027, n49028, n49029, n49030, n49031,
         n49032, n49033, n49034, n49035, n49036, n49037, n49038, n49039,
         n49040, n49041, n49042, n49043, n49044, n49045, n49046, n49047,
         n49048, n49049, n49050, n49051, n49052, n49053, n49054, n49055,
         n49056, n49057, n49058, n49059, n49060, n49061, n49062, n49063,
         n49064, n49065, n49066, n49067, n49068, n49069, n49070, n49071,
         n49072, n49073, n49074, n49075, n49076, n49077, n49078, n49079,
         n49080, n49081, n49082, n49083, n49084, n49085, n49086, n49087,
         n49088, n49089, n49090, n49091, n49092, n49093, n49094, n49095,
         n49096, n49097, n49098, n49099, n49100, n49101, n49102, n49103,
         n49104, n49105, n49106, n49107, n49108, n49109, n49110, n49111,
         n49112, n49113, n49114, n49115, n49116, n49117, n49118, n49119,
         n49120, n49121, n49122, n49123, n49124, n49125, n49126, n49127,
         n49128, n49129, n49130, n49131, n49132, n49133, n49134, n49135,
         n49136, n49137, n49138, n49139, n49140, n49141, n49142, n49143,
         n49144, n49145, n49146, n49147, n49148, n49149, n49150, n49151,
         n49152, n49153, n49154, n49155, n49156, n49157, n49158, n49159,
         n49160, n49161, n49162, n49163, n49164, n49165, n49166, n49167,
         n49168, n49169, n49170, n49171, n49172, n49173, n49174, n49175,
         n49176, n49177, n49178, n49179, n49180, n49181, n49182, n49183,
         n49184, n49185, n49186, n49187, n49188, n49189, n49190, n49191,
         n49192, n49193, n49194, n49195, n49196, n49197, n49198, n49199,
         n49200, n49201, n49202, n49203, n49204, n49205, n49206, n49207,
         n49208, n49209, n49210, n49211, n49212, n49213, n49214, n49215,
         n49216, n49217, n49218, n49219, n49220, n49221, n49222, n49223,
         n49224, n49225, n49226, n49227, n49228, n49229, n49230, n49231,
         n49232, n49233, n49234, n49235, n49236, n49237, n49238, n49239,
         n49240, n49241, n49242, n49243, n49244, n49245, n49246, n49247,
         n49248, n49249, n49250, n49251, n49252, n49253, n49254, n49255,
         n49256, n49257, n49258, n49259, n49260, n49261, n49262, n49263,
         n49264, n49265, n49266, n49267, n49268, n49269, n49270, n49271,
         n49272, n49273, n49274, n49275, n49276, n49277, n49278, n49279,
         n49280, n49281, n49282, n49283, n49284, n49285, n49286, n49287,
         n49288, n49289, n49290, n49291, n49292, n49293, n49294, n49295,
         n49296, n49297, n49298, n49299, n49300, n49301, n49302, n49303,
         n49304, n49305, n49306, n49307, n49308, n49309, n49310, n49311,
         n49312, n49313, n49314, n49315, n49316, n49317, n49318, n49319,
         n49320, n49321, n49322, n49323, n49324, n49325, n49326, n49327,
         n49328, n49329, n49330, n49331, n49332, n49333, n49334, n49335,
         n49336, n49337, n49338, n49339, n49340, n49341, n49342, n49343,
         n49344, n49345, n49346, n49347, n49348, n49349, n49350, n49351,
         n49352, n49353, n49354, n49355, n49356, n49357, n49358, n49359,
         n49360, n49361, n49362, n49363, n49364, n49365, n49366, n49367,
         n49368, n49369, n49370, n49371, n49372, n49373, n49374, n49375,
         n49376, n49377, n49378, n49379, n49380, n49381, n49382, n49383,
         n49384, n49385, n49386, n49387, n49388, n49389, n49390, n49391,
         n49392, n49393, n49394, n49395, n49396, n49397, n49398, n49399,
         n49400, n49401, n49402, n49403, n49404, n49405, n49406, n49407,
         n49408, n49409, n49410, n49411, n49412, n49413, n49414, n49415,
         n49416, n49417, n49418, n49419, n49420, n49421, n49422, n49423,
         n49424, n49425, n49426, n49427, n49428, n49429, n49430, n49431,
         n49432, n49433, n49434, n49435, n49436, n49437, n49438, n49439,
         n49440, n49441, n49442, n49443, n49444, n49445, n49446, n49447,
         n49448, n49449, n49450, n49451, n49452, n49453, n49454, n49455,
         n49456, n49457, n49458, n49459, n49460, n49461, n49462, n49463,
         n49464, n49465, n49466, n49467, n49468, n49469, n49470, n49471,
         n49472, n49473, n49474, n49475, n49476, n49477, n49478, n49479,
         n49480, n49481, n49482, n49483, n49484, n49485, n49486, n49487,
         n49488, n49489, n49490, n49491, n49492, n49493, n49494, n49495,
         n49496, n49497, n49498, n49499, n49500, n49501, n49502, n49503,
         n49504, n49505, n49506, n49507, n49508, n49509, n49510, n49511,
         n49512, n49513, n49514, n49515, n49516, n49517, n49518, n49519,
         n49520, n49521, n49522, n49523, n49524, n49525, n49526, n49527,
         n49528, n49529, n49530, n49531, n49532, n49533, n49534, n49535,
         n49536, n49537, n49538, n49539, n49540, n49541, n49542, n49543,
         n49544, n49545, n49546, n49547, n49548, n49549, n49550, n49551,
         n49552, n49553, n49554, n49555, n49556, n49557, n49558, n49559,
         n49560, n49561, n49562, n49563, n49564, n49565, n49566, n49567,
         n49568, n49569, n49570, n49571, n49572, n49573, n49574, n49575,
         n49576, n49577, n49578, n49579, n49580, n49581, n49582, n49583,
         n49584, n49585, n49586, n49587, n49588, n49589, n49590, n49591,
         n49592, n49593, n49594, n49595, n49596, n49597, n49598, n49599,
         n49600, n49601, n49602, n49603, n49604, n49605, n49606, n49607,
         n49608, n49609, n49610, n49611, n49612, n49613, n49614, n49615,
         n49616, n49617, n49618, n49619, n49620, n49621, n49622, n49623,
         n49624, n49625, n49626, n49627, n49628, n49629, n49630, n49631,
         n49632, n49633, n49634, n49635, n49636, n49637, n49638, n49639,
         n49640, n49641, n49642, n49643, n49644, n49645, n49646, n49647,
         n49648, n49649, n49650, n49651, n49652, n49653, n49654, n49655,
         n49656, n49657, n49658, n49659, n49660, n49661, n49662, n49663,
         n49664, n49665, n49666, n49667, n49668, n49669, n49670, n49671,
         n49672, n49673, n49674, n49675, n49676, n49677, n49678, n49679,
         n49680, n49681, n49682, n49683, n49684, n49685, n49686, n49687,
         n49688, n49689, n49690, n49691, n49692, n49693, n49694, n49695,
         n49696, n49697, n49698, n49699, n49700, n49701, n49702, n49703,
         n49704, n49705, n49706, n49707, n49708, n49709, n49710, n49711,
         n49712, n49713, n49714, n49715, n49716, n49717, n49718, n49719,
         n49720, n49721, n49722, n49723, n49724, n49725, n49726, n49727,
         n49728, n49729, n49730, n49731, n49732, n49733, n49734, n49735,
         n49736, n49737, n49738, n49739, n49740, n49741, n49742, n49743,
         n49744, n49745, n49746, n49747, n49748, n49749, n49750, n49751,
         n49752, n49753, n49754, n49755, n49756, n49757, n49758, n49759,
         n49760, n49761, n49762, n49763, n49764, n49765, n49766, n49767,
         n49768, n49769, n49770, n49771, n49772, n49773, n49774, n49775,
         n49776, n49777, n49778, n49779, n49780, n49781, n49782, n49783,
         n49784, n49785, n49786, n49787, n49788, n49789, n49790, n49791,
         n49792, n49793, n49794, n49795, n49796, n49797, n49798, n49799,
         n49800, n49801, n49802, n49803, n49804, n49805, n49806, n49807,
         n49808, n49809, n49810, n49811, n49812, n49813, n49814, n49815,
         n49816, n49817, n49818, n49819, n49820, n49821, n49822, n49823,
         n49824, n49825, n49826, n49827, n49828, n49829, n49830, n49831,
         n49832, n49833, n49834, n49835, n49836, n49837, n49838, n49839,
         n49840, n49841, n49842, n49843, n49844, n49845, n49846, n49847,
         n49848, n49849, n49850, n49851, n49852, n49853, n49854, n49855,
         n49856, n49857, n49858, n49859, n49860, n49861, n49862, n49863,
         n49864, n49865, n49866, n49867, n49868, n49869, n49870, n49871,
         n49872, n49873, n49874, n49875, n49876, n49877, n49878, n49879,
         n49880, n49881, n49882, n49883, n49884, n49885, n49886, n49887,
         n49888, n49889, n49890, n49891, n49892, n49893, n49894, n49895,
         n49896, n49897, n49898, n49899, n49900, n49901, n49902, n49903,
         n49904, n49905, n49906, n49907, n49908, n49909, n49910, n49911,
         n49912, n49913, n49914, n49915, n49916, n49917, n49918, n49919,
         n49920, n49921, n49922, n49923, n49924, n49925, n49926, n49927,
         n49928, n49929, n49930, n49931, n49932, n49933, n49934, n49935,
         n49936, n49937, n49938, n49939, n49940, n49941, n49942, n49943,
         n49944, n49945, n49946, n49947, n49948, n49949, n49950, n49951,
         n49952, n49953, n49954, n49955, n49956, n49957, n49958, n49959,
         n49960, n49961, n49962, n49963, n49964, n49965, n49966, n49967,
         n49968, n49969, n49970, n49971, n49972, n49973, n49974, n49975,
         n49976, n49977, n49978, n49979, n49980, n49981, n49982, n49983,
         n49984, n49985, n49986, n49987, n49988, n49989, n49990, n49991,
         n49992, n49993, n49994, n49995, n49996, n49997, n49998, n49999,
         n50000, n50001, n50002, n50003, n50004, n50005, n50006, n50007,
         n50008, n50009, n50010, n50011, n50012, n50013, n50014, n50015,
         n50016, n50017, n50018, n50019, n50020, n50021, n50022, n50023,
         n50024, n50025, n50026, n50027, n50028, n50029, n50030, n50031,
         n50032, n50033, n50034, n50035, n50036, n50037, n50038, n50039,
         n50040, n50041, n50042, n50043, n50044, n50045, n50046, n50047,
         n50048, n50049, n50050, n50051, n50052, n50053, n50054, n50055,
         n50056, n50057, n50058, n50059, n50060, n50061, n50062, n50063,
         n50064, n50065, n50066, n50067, n50068, n50069, n50070, n50071,
         n50072, n50073, n50074, n50075, n50076, n50077, n50078, n50079,
         n50080, n50081, n50082, n50083, n50084, n50085, n50086, n50087,
         n50088, n50089, n50090, n50091, n50092, n50093, n50094, n50095,
         n50096, n50097, n50098, n50099, n50100, n50101, n50102, n50103,
         n50104, n50105, n50106, n50107, n50108, n50109, n50110, n50111,
         n50112, n50113, n50114, n50115, n50116, n50117, n50118, n50119,
         n50120, n50121, n50122, n50123, n50124, n50125, n50126, n50127,
         n50128, n50129, n50130, n50131, n50132, n50133, n50134, n50135,
         n50136, n50137, n50138, n50139, n50140, n50141, n50142, n50143,
         n50144, n50145, n50146, n50147, n50148, n50149, n50150, n50151,
         n50152, n50153, n50154, n50155, n50156, n50157, n50158, n50159,
         n50160, n50161, n50162, n50163, n50164, n50165, n50166, n50167,
         n50168, n50169, n50170, n50171, n50172, n50173, n50174, n50175,
         n50176, n50177, n50178, n50179, n50180, n50181, n50182, n50183,
         n50184, n50185, n50186, n50187, n50188, n50189, n50190, n50191,
         n50192, n50193, n50194, n50195, n50196, n50197, n50198, n50199,
         n50200, n50201, n50202, n50203, n50204, n50205, n50206, n50207,
         n50208, n50209, n50210, n50211, n50212, n50213, n50214, n50215,
         n50216, n50217, n50218, n50219, n50220, n50221, n50222, n50223,
         n50224, n50225, n50226, n50227, n50228, n50229, n50230, n50231,
         n50232, n50233, n50234, n50235, n50236, n50237, n50238, n50239,
         n50240, n50241, n50242, n50243, n50244, n50245, n50246, n50247,
         n50248, n50249, n50250, n50251, n50252, n50253, n50254, n50255,
         n50256, n50257, n50258, n50259, n50260, n50261, n50262, n50263,
         n50264, n50265, n50266, n50267, n50268, n50269, n50270, n50271,
         n50272, n50273, n50274, n50275, n50276, n50277, n50278, n50279,
         n50280, n50281, n50282, n50283, n50284, n50285, n50286, n50287,
         n50288, n50289, n50290, n50291, n50292, n50293, n50294, n50295,
         n50296, n50297, n50298, n50299, n50300, n50301, n50302, n50303,
         n50304, n50305, n50306, n50307, n50308, n50309, n50310, n50311,
         n50312, n50313, n50314, n50315, n50316, n50317, n50318, n50319,
         n50320, n50321, n50322, n50323, n50324, n50325, n50326, n50327,
         n50328, n50329, n50330, n50331, n50332, n50333, n50334, n50335,
         n50336, n50337, n50338, n50339, n50340, n50341, n50342, n50343,
         n50344, n50345, n50346, n50347, n50348, n50349, n50350, n50351,
         n50352, n50353, n50354, n50355, n50356, n50357, n50358, n50359,
         n50360, n50361, n50362, n50363, n50364, n50365, n50366, n50367,
         n50368, n50369, n50370, n50371, n50372, n50373, n50374, n50375,
         n50376, n50377, n50378, n50379, n50380, n50381, n50382, n50383,
         n50384, n50385, n50386, n50387, n50388, n50389, n50390, n50391,
         n50392, n50393, n50394, n50395, n50396, n50397, n50398, n50399,
         n50400, n50401, n50402, n50403, n50404, n50405, n50406, n50407,
         n50408, n50409, n50410, n50411, n50412, n50413, n50414, n50415,
         n50416, n50417, n50418, n50419, n50420, n50421, n50422, n50423,
         n50424, n50425, n50426, n50427, n50428, n50429, n50430, n50431,
         n50432, n50433, n50434, n50435, n50436, n50437, n50438, n50439,
         n50440, n50441, n50442, n50443, n50444, n50445, n50446, n50447,
         n50448, n50449, n50450, n50451, n50452, n50453, n50454, n50455,
         n50456, n50457, n50458, n50459, n50460, n50461, n50462, n50463,
         n50464, n50465, n50466, n50467, n50468, n50469, n50470, n50471,
         n50472, n50473, n50474, n50475, n50476, n50477, n50478, n50479,
         n50480, n50481, n50482, n50483, n50484, n50485, n50486, n50487,
         n50488, n50489, n50490, n50491, n50492, n50493, n50494, n50495,
         n50496, n50497, n50498, n50499, n50500, n50501, n50502, n50503,
         n50504, n50505, n50506, n50507, n50508, n50509, n50510, n50511,
         n50512, n50513, n50514, n50515, n50516, n50517, n50518, n50519,
         n50520, n50521, n50522, n50523, n50524, n50525, n50526, n50527,
         n50528, n50529, n50530, n50531, n50532, n50533, n50534, n50535,
         n50536, n50537, n50538, n50539, n50540, n50541, n50542, n50543,
         n50544, n50545, n50546, n50547, n50548, n50549, n50550, n50551,
         n50552, n50553, n50554, n50555, n50556, n50557, n50558, n50559,
         n50560, n50561, n50562, n50563, n50564, n50565, n50566, n50567,
         n50568, n50569, n50570, n50571, n50572, n50573, n50574, n50575,
         n50576, n50577, n50578, n50579, n50580, n50581, n50582, n50583,
         n50584, n50585, n50586, n50587, n50588, n50589, n50590, n50591,
         n50592, n50593, n50594, n50595, n50596, n50597, n50598, n50599,
         n50600, n50601, n50602, n50603, n50604, n50605, n50606, n50607,
         n50608, n50609, n50610, n50611, n50612, n50613, n50614, n50615,
         n50616, n50617, n50618, n50619, n50620, n50621, n50622, n50623,
         n50624, n50625, n50626, n50627, n50628, n50629, n50630, n50631,
         n50632, n50633, n50634, n50635, n50636, n50637, n50638, n50639,
         n50640, n50641, n50642, n50643, n50644, n50645, n50646, n50647,
         n50648, n50649, n50650, n50651, n50652, n50653, n50654, n50655,
         n50656, n50657, n50658, n50659, n50660, n50661, n50662, n50663,
         n50664, n50665, n50666, n50667, n50668, n50669, n50670, n50671,
         n50672, n50673, n50674, n50675, n50676, n50677, n50678, n50679,
         n50680, n50681, n50682, n50683, n50684, n50685, n50686, n50687,
         n50688, n50689, n50690, n50691, n50692, n50693, n50694, n50695,
         n50696, n50697, n50698, n50699, n50700, n50701, n50702, n50703,
         n50704, n50705, n50706, n50707, n50708, n50709, n50710, n50711,
         n50712, n50713, n50714, n50715, n50716, n50717, n50718, n50719,
         n50720, n50721, n50722, n50723, n50724, n50725, n50726, n50727,
         n50728, n50729, n50730, n50731, n50732, n50733, n50734, n50735,
         n50736, n50737, n50738, n50739, n50740, n50741, n50742, n50743,
         n50744, n50745, n50746, n50747, n50748, n50749, n50750, n50751,
         n50752, n50753, n50754, n50755, n50756, n50757, n50758, n50759,
         n50760, n50761, n50762, n50763, n50764, n50765, n50766, n50767,
         n50768, n50769, n50770, n50771, n50772, n50773, n50774, n50775,
         n50776, n50777, n50778, n50779, n50780, n50781, n50782, n50783,
         n50784, n50785, n50786, n50787, n50788, n50789, n50790, n50791,
         n50792, n50793, n50794, n50795, n50796, n50797, n50798, n50799,
         n50800, n50801, n50802, n50803, n50804, n50805, n50806, n50807,
         n50808, n50809, n50810, n50811, n50812, n50813, n50814, n50815,
         n50816, n50817, n50818, n50819, n50820, n50821, n50822, n50823,
         n50824, n50825, n50826, n50827, n50828, n50829, n50830, n50831,
         n50832, n50833, n50834, n50835, n50836, n50837, n50838, n50839,
         n50840, n50841, n50842, n50843, n50844, n50845, n50846, n50847,
         n50848, n50849, n50850, n50851, n50852, n50853, n50854, n50855,
         n50856, n50857, n50858, n50859, n50860, n50861, n50862, n50863,
         n50864, n50865, n50866, n50867, n50868, n50869, n50870, n50871,
         n50872, n50873, n50874, n50875, n50876, n50877, n50878, n50879,
         n50880, n50881, n50882, n50883, n50884, n50885, n50886, n50887,
         n50888, n50889, n50890, n50891, n50892, n50893, n50894, n50895,
         n50896, n50897, n50898, n50899, n50900, n50901, n50902, n50903,
         n50904, n50905, n50906, n50907, n50908, n50909, n50910, n50911,
         n50912, n50913, n50914, n50915, n50916, n50917, n50918, n50919,
         n50920, n50921, n50922, n50923, n50924, n50925, n50926, n50927,
         n50928, n50929, n50930, n50931, n50932, n50933, n50934, n50935,
         n50936, n50937, n50938, n50939, n50940, n50941, n50942, n50943,
         n50944, n50945, n50946, n50947, n50948, n50949, n50950, n50951,
         n50952, n50953, n50954, n50955, n50956, n50957, n50958, n50959,
         n50960, n50961, n50962, n50963, n50964, n50965, n50966, n50967,
         n50968, n50969, n50970, n50971, n50972, n50973, n50974, n50975,
         n50976, n50977, n50978, n50979, n50980, n50981, n50982, n50983,
         n50984, n50985, n50986, n50987, n50988, n50989, n50990, n50991,
         n50992, n50993, n50994, n50995, n50996, n50997, n50998, n50999,
         n51000, n51001, n51002, n51003, n51004, n51005, n51006, n51007,
         n51008, n51009, n51010, n51011, n51012, n51013, n51014, n51015,
         n51016, n51017, n51018, n51019, n51020, n51021, n51022, n51023,
         n51024, n51025, n51026, n51027, n51028, n51029, n51030, n51031,
         n51032, n51033, n51034, n51035, n51036, n51037, n51038, n51039,
         n51040, n51041, n51042, n51043, n51044, n51045, n51046, n51047,
         n51048, n51049, n51050, n51051, n51052, n51053, n51054, n51055,
         n51056, n51057, n51058, n51059, n51060, n51061, n51062, n51063,
         n51064, n51065, n51066, n51067, n51068, n51069, n51070, n51071,
         n51072, n51073, n51074, n51075, n51076, n51077, n51078, n51079,
         n51080, n51081, n51082, n51083, n51084, n51085, n51086, n51087,
         n51088, n51089, n51090, n51091, n51092, n51093, n51094, n51095,
         n51096, n51097, n51098, n51099, n51100, n51101, n51102, n51103,
         n51104, n51105, n51106, n51107, n51108, n51109, n51110, n51111,
         n51112, n51113, n51114, n51115, n51116, n51117, n51118, n51119,
         n51120, n51121, n51122, n51123, n51124, n51125, n51126, n51127,
         n51128, n51129, n51130, n51131, n51132, n51133, n51134, n51135,
         n51136, n51137, n51138, n51139, n51140, n51141, n51142, n51143,
         n51144, n51145, n51146, n51147, n51148, n51149, n51150, n51151,
         n51152, n51153, n51154, n51155, n51156, n51157, n51158, n51159,
         n51160, n51161, n51162, n51163, n51164, n51165, n51166, n51167,
         n51168, n51169, n51170, n51171, n51172, n51173, n51174, n51175,
         n51176, n51177, n51178, n51179, n51180, n51181, n51182, n51183,
         n51184, n51185, n51186, n51187, n51188, n51189, n51190, n51191,
         n51192, n51193, n51194, n51195, n51196, n51197, n51198, n51199,
         n51200, n51201, n51202, n51203, n51204, n51205, n51206, n51207,
         n51208, n51209, n51210, n51211, n51212, n51213, n51214, n51215,
         n51216, n51217, n51218, n51219, n51220, n51221, n51222, n51223,
         n51224, n51225, n51226, n51227, n51228, n51229, n51230, n51231,
         n51232, n51233, n51234, n51235, n51236, n51237, n51238, n51239,
         n51240, n51241, n51242, n51243, n51244, n51245, n51246, n51247,
         n51248, n51249, n51250, n51251, n51252, n51253, n51254, n51255,
         n51256, n51257, n51258, n51259, n51260, n51261, n51262, n51263,
         n51264, n51265, n51266, n51267, n51268, n51269, n51270, n51271,
         n51272, n51273, n51274, n51275, n51276, n51277, n51278, n51279,
         n51280, n51281, n51282, n51283, n51284, n51285, n51286, n51287,
         n51288, n51289, n51290, n51291, n51292, n51293, n51294, n51295,
         n51296, n51297, n51298, n51299, n51300, n51301, n51302, n51303,
         n51304, n51305, n51306, n51307, n51308, n51309, n51310, n51311,
         n51312, n51313, n51314, n51315, n51316, n51317, n51318, n51319,
         n51320, n51321, n51322, n51323, n51324, n51325, n51326, n51327,
         n51328, n51329, n51330, n51331, n51332, n51333, n51334, n51335,
         n51336, n51337, n51338, n51339, n51340, n51341, n51342, n51343,
         n51344, n51345, n51346, n51347, n51348, n51349, n51350, n51351,
         n51352, n51353, n51354, n51355, n51356, n51357, n51358, n51359,
         n51360, n51361, n51362, n51363, n51364, n51365, n51366, n51367,
         n51368, n51369, n51370, n51371, n51372, n51373, n51374, n51375,
         n51376, n51377, n51378, n51379, n51380, n51381, n51382, n51383,
         n51384, n51385, n51386, n51387, n51388, n51389, n51390, n51391,
         n51392, n51393, n51394, n51395, n51396, n51397, n51398, n51399,
         n51400, n51401, n51402, n51403, n51404, n51405, n51406, n51407,
         n51408, n51409, n51410, n51411, n51412, n51413, n51414, n51415,
         n51416, n51417, n51418, n51419, n51420, n51421, n51422, n51423,
         n51424, n51425, n51426, n51427, n51428, n51429, n51430, n51431,
         n51432, n51433, n51434, n51435, n51436, n51437, n51438, n51439,
         n51440, n51441, n51442, n51443, n51444, n51445, n51446, n51447,
         n51448, n51449, n51450, n51451, n51452, n51453, n51454, n51455,
         n51456, n51457, n51458, n51459, n51460, n51461, n51462, n51463,
         n51464, n51465, n51466, n51467, n51468, n51469, n51470, n51471,
         n51472, n51473, n51474, n51475, n51476, n51477, n51478, n51479,
         n51480, n51481, n51482, n51483, n51484, n51485, n51486, n51487,
         n51488, n51489, n51490, n51491, n51492, n51493, n51494, n51495,
         n51496, n51497, n51498, n51499, n51500, n51501, n51502, n51503,
         n51504, n51505, n51506, n51507, n51508, n51509, n51510, n51511,
         n51512, n51513, n51514, n51515, n51516, n51517, n51518, n51519,
         n51520, n51521, n51522, n51523, n51524, n51525, n51526, n51527,
         n51528, n51529, n51530;
  wire   [3:0] reg_num;
  wire   [19:0] out_L1;
  wire   [19:0] out_L2;

  dff_sg done_reg ( .D(n51529), .CP(clk), .Q(done) );
  dff_sg \state_reg[1]  ( .D(n1999), .CP(clk), .Q(state[1]) );
  dff_sg \state_reg[0]  ( .D(n1998), .CP(clk), .Q(state[0]) );
  dff_sg \reg_num_reg[3]  ( .D(n1353), .CP(clk), .Q(reg_num[3]) );
  dff_sg \reg_num_reg[2]  ( .D(n1354), .CP(clk), .Q(reg_num[2]) );
  dff_sg \reg_num_reg[1]  ( .D(n1355), .CP(clk), .Q(reg_num[1]) );
  dff_sg \reg_num_reg[0]  ( .D(n1356), .CP(clk), .Q(reg_num[0]) );
  dff_sg \reg_y_reg[14][19]  ( .D(n1377), .CP(clk), .Q(\reg_y[14][19] ) );
  dff_sg \reg_y_reg[14][18]  ( .D(n1378), .CP(clk), .Q(\reg_y[14][18] ) );
  dff_sg \reg_y_reg[14][17]  ( .D(n1379), .CP(clk), .Q(\reg_y[14][17] ) );
  dff_sg \reg_y_reg[14][16]  ( .D(n1380), .CP(clk), .Q(\reg_y[14][16] ) );
  dff_sg \reg_y_reg[14][15]  ( .D(n1381), .CP(clk), .Q(\reg_y[14][15] ) );
  dff_sg \reg_y_reg[14][14]  ( .D(n1382), .CP(clk), .Q(\reg_y[14][14] ) );
  dff_sg \reg_y_reg[14][13]  ( .D(n1383), .CP(clk), .Q(\reg_y[14][13] ) );
  dff_sg \reg_y_reg[14][12]  ( .D(n1384), .CP(clk), .Q(\reg_y[14][12] ) );
  dff_sg \reg_y_reg[14][11]  ( .D(n1385), .CP(clk), .Q(\reg_y[14][11] ) );
  dff_sg \reg_y_reg[14][10]  ( .D(n1386), .CP(clk), .Q(\reg_y[14][10] ) );
  dff_sg \reg_y_reg[14][9]  ( .D(n1387), .CP(clk), .Q(\reg_y[14][9] ) );
  dff_sg \reg_y_reg[14][8]  ( .D(n1388), .CP(clk), .Q(\reg_y[14][8] ) );
  dff_sg \reg_y_reg[14][7]  ( .D(n1389), .CP(clk), .Q(\reg_y[14][7] ) );
  dff_sg \reg_y_reg[14][6]  ( .D(n1390), .CP(clk), .Q(\reg_y[14][6] ) );
  dff_sg \reg_y_reg[14][5]  ( .D(n1391), .CP(clk), .Q(\reg_y[14][5] ) );
  dff_sg \reg_y_reg[14][4]  ( .D(n1392), .CP(clk), .Q(\reg_y[14][4] ) );
  dff_sg \reg_y_reg[14][3]  ( .D(n1393), .CP(clk), .Q(\reg_y[14][3] ) );
  dff_sg \reg_y_reg[14][2]  ( .D(n1394), .CP(clk), .Q(\reg_y[14][2] ) );
  dff_sg \reg_y_reg[14][1]  ( .D(n1395), .CP(clk), .Q(\reg_y[14][1] ) );
  dff_sg \reg_y_reg[14][0]  ( .D(n1396), .CP(clk), .Q(\reg_y[14][0] ) );
  dff_sg \reg_y_reg[13][19]  ( .D(n1397), .CP(clk), .Q(\reg_y[13][19] ) );
  dff_sg \reg_y_reg[13][18]  ( .D(n1398), .CP(clk), .Q(\reg_y[13][18] ) );
  dff_sg \reg_y_reg[13][17]  ( .D(n1399), .CP(clk), .Q(\reg_y[13][17] ) );
  dff_sg \reg_y_reg[13][16]  ( .D(n1400), .CP(clk), .Q(\reg_y[13][16] ) );
  dff_sg \reg_y_reg[13][15]  ( .D(n1401), .CP(clk), .Q(\reg_y[13][15] ) );
  dff_sg \reg_y_reg[13][14]  ( .D(n1402), .CP(clk), .Q(\reg_y[13][14] ) );
  dff_sg \reg_y_reg[13][13]  ( .D(n1403), .CP(clk), .Q(\reg_y[13][13] ) );
  dff_sg \reg_y_reg[13][12]  ( .D(n1404), .CP(clk), .Q(\reg_y[13][12] ) );
  dff_sg \reg_y_reg[13][11]  ( .D(n1405), .CP(clk), .Q(\reg_y[13][11] ) );
  dff_sg \reg_y_reg[13][10]  ( .D(n1406), .CP(clk), .Q(\reg_y[13][10] ) );
  dff_sg \reg_y_reg[13][9]  ( .D(n1407), .CP(clk), .Q(\reg_y[13][9] ) );
  dff_sg \reg_y_reg[13][8]  ( .D(n1408), .CP(clk), .Q(\reg_y[13][8] ) );
  dff_sg \reg_y_reg[13][7]  ( .D(n1409), .CP(clk), .Q(\reg_y[13][7] ) );
  dff_sg \reg_y_reg[13][6]  ( .D(n1410), .CP(clk), .Q(\reg_y[13][6] ) );
  dff_sg \reg_y_reg[13][5]  ( .D(n1411), .CP(clk), .Q(\reg_y[13][5] ) );
  dff_sg \reg_y_reg[13][4]  ( .D(n1412), .CP(clk), .Q(\reg_y[13][4] ) );
  dff_sg \reg_y_reg[13][3]  ( .D(n1413), .CP(clk), .Q(\reg_y[13][3] ) );
  dff_sg \reg_y_reg[13][2]  ( .D(n1414), .CP(clk), .Q(\reg_y[13][2] ) );
  dff_sg \reg_y_reg[13][1]  ( .D(n1415), .CP(clk), .Q(\reg_y[13][1] ) );
  dff_sg \reg_y_reg[13][0]  ( .D(n1416), .CP(clk), .Q(\reg_y[13][0] ) );
  dff_sg \reg_y_reg[12][19]  ( .D(n1417), .CP(clk), .Q(\reg_y[12][19] ) );
  dff_sg \reg_y_reg[12][18]  ( .D(n1418), .CP(clk), .Q(\reg_y[12][18] ) );
  dff_sg \reg_y_reg[12][17]  ( .D(n1419), .CP(clk), .Q(\reg_y[12][17] ) );
  dff_sg \reg_y_reg[12][16]  ( .D(n1420), .CP(clk), .Q(\reg_y[12][16] ) );
  dff_sg \reg_y_reg[12][15]  ( .D(n1421), .CP(clk), .Q(\reg_y[12][15] ) );
  dff_sg \reg_y_reg[12][14]  ( .D(n1422), .CP(clk), .Q(\reg_y[12][14] ) );
  dff_sg \reg_y_reg[12][13]  ( .D(n1423), .CP(clk), .Q(\reg_y[12][13] ) );
  dff_sg \reg_y_reg[12][12]  ( .D(n1424), .CP(clk), .Q(\reg_y[12][12] ) );
  dff_sg \reg_y_reg[12][11]  ( .D(n1425), .CP(clk), .Q(\reg_y[12][11] ) );
  dff_sg \reg_y_reg[12][10]  ( .D(n1426), .CP(clk), .Q(\reg_y[12][10] ) );
  dff_sg \reg_y_reg[12][9]  ( .D(n1427), .CP(clk), .Q(\reg_y[12][9] ) );
  dff_sg \reg_y_reg[12][8]  ( .D(n1428), .CP(clk), .Q(\reg_y[12][8] ) );
  dff_sg \reg_y_reg[12][7]  ( .D(n1429), .CP(clk), .Q(\reg_y[12][7] ) );
  dff_sg \reg_y_reg[12][6]  ( .D(n1430), .CP(clk), .Q(\reg_y[12][6] ) );
  dff_sg \reg_y_reg[12][5]  ( .D(n1431), .CP(clk), .Q(\reg_y[12][5] ) );
  dff_sg \reg_y_reg[12][4]  ( .D(n1432), .CP(clk), .Q(\reg_y[12][4] ) );
  dff_sg \reg_y_reg[12][3]  ( .D(n1433), .CP(clk), .Q(\reg_y[12][3] ) );
  dff_sg \reg_y_reg[12][2]  ( .D(n1434), .CP(clk), .Q(\reg_y[12][2] ) );
  dff_sg \reg_y_reg[12][1]  ( .D(n1435), .CP(clk), .Q(\reg_y[12][1] ) );
  dff_sg \reg_y_reg[12][0]  ( .D(n1436), .CP(clk), .Q(\reg_y[12][0] ) );
  dff_sg \reg_y_reg[11][19]  ( .D(n1437), .CP(clk), .Q(\reg_y[11][19] ) );
  dff_sg \reg_y_reg[11][18]  ( .D(n1438), .CP(clk), .Q(\reg_y[11][18] ) );
  dff_sg \reg_y_reg[11][17]  ( .D(n1439), .CP(clk), .Q(\reg_y[11][17] ) );
  dff_sg \reg_y_reg[11][16]  ( .D(n1440), .CP(clk), .Q(\reg_y[11][16] ) );
  dff_sg \reg_y_reg[11][15]  ( .D(n1441), .CP(clk), .Q(\reg_y[11][15] ) );
  dff_sg \reg_y_reg[11][14]  ( .D(n1442), .CP(clk), .Q(\reg_y[11][14] ) );
  dff_sg \reg_y_reg[11][13]  ( .D(n1443), .CP(clk), .Q(\reg_y[11][13] ) );
  dff_sg \reg_y_reg[11][12]  ( .D(n1444), .CP(clk), .Q(\reg_y[11][12] ) );
  dff_sg \reg_y_reg[11][11]  ( .D(n1445), .CP(clk), .Q(\reg_y[11][11] ) );
  dff_sg \reg_y_reg[11][10]  ( .D(n1446), .CP(clk), .Q(\reg_y[11][10] ) );
  dff_sg \reg_y_reg[11][9]  ( .D(n1447), .CP(clk), .Q(\reg_y[11][9] ) );
  dff_sg \reg_y_reg[11][8]  ( .D(n1448), .CP(clk), .Q(\reg_y[11][8] ) );
  dff_sg \reg_y_reg[11][7]  ( .D(n1449), .CP(clk), .Q(\reg_y[11][7] ) );
  dff_sg \reg_y_reg[11][6]  ( .D(n1450), .CP(clk), .Q(\reg_y[11][6] ) );
  dff_sg \reg_y_reg[11][5]  ( .D(n1451), .CP(clk), .Q(\reg_y[11][5] ) );
  dff_sg \reg_y_reg[11][4]  ( .D(n1452), .CP(clk), .Q(\reg_y[11][4] ) );
  dff_sg \reg_y_reg[11][3]  ( .D(n1453), .CP(clk), .Q(\reg_y[11][3] ) );
  dff_sg \reg_y_reg[11][2]  ( .D(n1454), .CP(clk), .Q(\reg_y[11][2] ) );
  dff_sg \reg_y_reg[11][1]  ( .D(n1455), .CP(clk), .Q(\reg_y[11][1] ) );
  dff_sg \reg_y_reg[11][0]  ( .D(n1456), .CP(clk), .Q(\reg_y[11][0] ) );
  dff_sg \reg_y_reg[10][19]  ( .D(n1457), .CP(clk), .Q(\reg_y[10][19] ) );
  dff_sg \reg_y_reg[10][18]  ( .D(n1458), .CP(clk), .Q(\reg_y[10][18] ) );
  dff_sg \reg_y_reg[10][17]  ( .D(n1459), .CP(clk), .Q(\reg_y[10][17] ) );
  dff_sg \reg_y_reg[10][16]  ( .D(n1460), .CP(clk), .Q(\reg_y[10][16] ) );
  dff_sg \reg_y_reg[10][15]  ( .D(n1461), .CP(clk), .Q(\reg_y[10][15] ) );
  dff_sg \reg_y_reg[10][14]  ( .D(n1462), .CP(clk), .Q(\reg_y[10][14] ) );
  dff_sg \reg_y_reg[10][13]  ( .D(n1463), .CP(clk), .Q(\reg_y[10][13] ) );
  dff_sg \reg_y_reg[10][12]  ( .D(n1464), .CP(clk), .Q(\reg_y[10][12] ) );
  dff_sg \reg_y_reg[10][11]  ( .D(n1465), .CP(clk), .Q(\reg_y[10][11] ) );
  dff_sg \reg_y_reg[10][10]  ( .D(n1466), .CP(clk), .Q(\reg_y[10][10] ) );
  dff_sg \reg_y_reg[10][9]  ( .D(n1467), .CP(clk), .Q(\reg_y[10][9] ) );
  dff_sg \reg_y_reg[10][8]  ( .D(n1468), .CP(clk), .Q(\reg_y[10][8] ) );
  dff_sg \reg_y_reg[10][7]  ( .D(n1469), .CP(clk), .Q(\reg_y[10][7] ) );
  dff_sg \reg_y_reg[10][6]  ( .D(n1470), .CP(clk), .Q(\reg_y[10][6] ) );
  dff_sg \reg_y_reg[10][5]  ( .D(n1471), .CP(clk), .Q(\reg_y[10][5] ) );
  dff_sg \reg_y_reg[10][4]  ( .D(n1472), .CP(clk), .Q(\reg_y[10][4] ) );
  dff_sg \reg_y_reg[10][3]  ( .D(n1473), .CP(clk), .Q(\reg_y[10][3] ) );
  dff_sg \reg_y_reg[10][2]  ( .D(n1474), .CP(clk), .Q(\reg_y[10][2] ) );
  dff_sg \reg_y_reg[10][1]  ( .D(n1475), .CP(clk), .Q(\reg_y[10][1] ) );
  dff_sg \reg_y_reg[10][0]  ( .D(n1476), .CP(clk), .Q(\reg_y[10][0] ) );
  dff_sg \reg_y_reg[9][19]  ( .D(n1477), .CP(clk), .Q(\reg_y[9][19] ) );
  dff_sg \reg_y_reg[9][18]  ( .D(n1478), .CP(clk), .Q(\reg_y[9][18] ) );
  dff_sg \reg_y_reg[9][17]  ( .D(n1479), .CP(clk), .Q(\reg_y[9][17] ) );
  dff_sg \reg_y_reg[9][16]  ( .D(n1480), .CP(clk), .Q(\reg_y[9][16] ) );
  dff_sg \reg_y_reg[9][15]  ( .D(n1481), .CP(clk), .Q(\reg_y[9][15] ) );
  dff_sg \reg_y_reg[9][14]  ( .D(n1482), .CP(clk), .Q(\reg_y[9][14] ) );
  dff_sg \reg_y_reg[9][13]  ( .D(n1483), .CP(clk), .Q(\reg_y[9][13] ) );
  dff_sg \reg_y_reg[9][12]  ( .D(n1484), .CP(clk), .Q(\reg_y[9][12] ) );
  dff_sg \reg_y_reg[9][11]  ( .D(n1485), .CP(clk), .Q(\reg_y[9][11] ) );
  dff_sg \reg_y_reg[9][10]  ( .D(n1486), .CP(clk), .Q(\reg_y[9][10] ) );
  dff_sg \reg_y_reg[9][9]  ( .D(n1487), .CP(clk), .Q(\reg_y[9][9] ) );
  dff_sg \reg_y_reg[9][8]  ( .D(n1488), .CP(clk), .Q(\reg_y[9][8] ) );
  dff_sg \reg_y_reg[9][7]  ( .D(n1489), .CP(clk), .Q(\reg_y[9][7] ) );
  dff_sg \reg_y_reg[9][6]  ( .D(n1490), .CP(clk), .Q(\reg_y[9][6] ) );
  dff_sg \reg_y_reg[9][5]  ( .D(n1491), .CP(clk), .Q(\reg_y[9][5] ) );
  dff_sg \reg_y_reg[9][4]  ( .D(n1492), .CP(clk), .Q(\reg_y[9][4] ) );
  dff_sg \reg_y_reg[9][3]  ( .D(n1493), .CP(clk), .Q(\reg_y[9][3] ) );
  dff_sg \reg_y_reg[9][2]  ( .D(n1494), .CP(clk), .Q(\reg_y[9][2] ) );
  dff_sg \reg_y_reg[9][1]  ( .D(n1495), .CP(clk), .Q(\reg_y[9][1] ) );
  dff_sg \reg_y_reg[9][0]  ( .D(n1496), .CP(clk), .Q(\reg_y[9][0] ) );
  dff_sg \reg_y_reg[8][19]  ( .D(n1497), .CP(clk), .Q(\reg_y[8][19] ) );
  dff_sg \reg_y_reg[8][18]  ( .D(n1498), .CP(clk), .Q(\reg_y[8][18] ) );
  dff_sg \reg_y_reg[8][17]  ( .D(n1499), .CP(clk), .Q(\reg_y[8][17] ) );
  dff_sg \reg_y_reg[8][16]  ( .D(n1500), .CP(clk), .Q(\reg_y[8][16] ) );
  dff_sg \reg_y_reg[8][15]  ( .D(n1501), .CP(clk), .Q(\reg_y[8][15] ) );
  dff_sg \reg_y_reg[8][14]  ( .D(n1502), .CP(clk), .Q(\reg_y[8][14] ) );
  dff_sg \reg_y_reg[8][13]  ( .D(n1503), .CP(clk), .Q(\reg_y[8][13] ) );
  dff_sg \reg_y_reg[8][12]  ( .D(n1504), .CP(clk), .Q(\reg_y[8][12] ) );
  dff_sg \reg_y_reg[8][11]  ( .D(n1505), .CP(clk), .Q(\reg_y[8][11] ) );
  dff_sg \reg_y_reg[8][10]  ( .D(n1506), .CP(clk), .Q(\reg_y[8][10] ) );
  dff_sg \reg_y_reg[8][9]  ( .D(n1507), .CP(clk), .Q(\reg_y[8][9] ) );
  dff_sg \reg_y_reg[8][8]  ( .D(n1508), .CP(clk), .Q(\reg_y[8][8] ) );
  dff_sg \reg_y_reg[8][7]  ( .D(n1509), .CP(clk), .Q(\reg_y[8][7] ) );
  dff_sg \reg_y_reg[8][6]  ( .D(n1510), .CP(clk), .Q(\reg_y[8][6] ) );
  dff_sg \reg_y_reg[8][5]  ( .D(n1511), .CP(clk), .Q(\reg_y[8][5] ) );
  dff_sg \reg_y_reg[8][4]  ( .D(n1512), .CP(clk), .Q(\reg_y[8][4] ) );
  dff_sg \reg_y_reg[8][3]  ( .D(n1513), .CP(clk), .Q(\reg_y[8][3] ) );
  dff_sg \reg_y_reg[8][2]  ( .D(n1514), .CP(clk), .Q(\reg_y[8][2] ) );
  dff_sg \reg_y_reg[8][1]  ( .D(n1515), .CP(clk), .Q(\reg_y[8][1] ) );
  dff_sg \reg_y_reg[8][0]  ( .D(n1516), .CP(clk), .Q(\reg_y[8][0] ) );
  dff_sg \reg_y_reg[7][19]  ( .D(n1517), .CP(clk), .Q(\reg_y[7][19] ) );
  dff_sg \reg_y_reg[7][18]  ( .D(n1518), .CP(clk), .Q(\reg_y[7][18] ) );
  dff_sg \reg_y_reg[7][17]  ( .D(n1519), .CP(clk), .Q(\reg_y[7][17] ) );
  dff_sg \reg_y_reg[7][16]  ( .D(n1520), .CP(clk), .Q(\reg_y[7][16] ) );
  dff_sg \reg_y_reg[7][15]  ( .D(n1521), .CP(clk), .Q(\reg_y[7][15] ) );
  dff_sg \reg_y_reg[7][14]  ( .D(n1522), .CP(clk), .Q(\reg_y[7][14] ) );
  dff_sg \reg_y_reg[7][13]  ( .D(n1523), .CP(clk), .Q(\reg_y[7][13] ) );
  dff_sg \reg_y_reg[7][12]  ( .D(n1524), .CP(clk), .Q(\reg_y[7][12] ) );
  dff_sg \reg_y_reg[7][11]  ( .D(n1525), .CP(clk), .Q(\reg_y[7][11] ) );
  dff_sg \reg_y_reg[7][10]  ( .D(n1526), .CP(clk), .Q(\reg_y[7][10] ) );
  dff_sg \reg_y_reg[7][9]  ( .D(n1527), .CP(clk), .Q(\reg_y[7][9] ) );
  dff_sg \reg_y_reg[7][8]  ( .D(n1528), .CP(clk), .Q(\reg_y[7][8] ) );
  dff_sg \reg_y_reg[7][7]  ( .D(n1529), .CP(clk), .Q(\reg_y[7][7] ) );
  dff_sg \reg_y_reg[7][6]  ( .D(n1530), .CP(clk), .Q(\reg_y[7][6] ) );
  dff_sg \reg_y_reg[7][5]  ( .D(n1531), .CP(clk), .Q(\reg_y[7][5] ) );
  dff_sg \reg_y_reg[7][4]  ( .D(n1532), .CP(clk), .Q(\reg_y[7][4] ) );
  dff_sg \reg_y_reg[7][3]  ( .D(n1533), .CP(clk), .Q(\reg_y[7][3] ) );
  dff_sg \reg_y_reg[7][2]  ( .D(n1534), .CP(clk), .Q(\reg_y[7][2] ) );
  dff_sg \reg_y_reg[7][1]  ( .D(n1535), .CP(clk), .Q(\reg_y[7][1] ) );
  dff_sg \reg_y_reg[7][0]  ( .D(n1536), .CP(clk), .Q(\reg_y[7][0] ) );
  dff_sg \reg_y_reg[6][19]  ( .D(n1537), .CP(clk), .Q(\reg_y[6][19] ) );
  dff_sg \reg_y_reg[6][18]  ( .D(n1538), .CP(clk), .Q(\reg_y[6][18] ) );
  dff_sg \reg_y_reg[6][17]  ( .D(n1539), .CP(clk), .Q(\reg_y[6][17] ) );
  dff_sg \reg_y_reg[6][16]  ( .D(n1540), .CP(clk), .Q(\reg_y[6][16] ) );
  dff_sg \reg_y_reg[6][15]  ( .D(n1541), .CP(clk), .Q(\reg_y[6][15] ) );
  dff_sg \reg_y_reg[6][14]  ( .D(n1542), .CP(clk), .Q(\reg_y[6][14] ) );
  dff_sg \reg_y_reg[6][13]  ( .D(n1543), .CP(clk), .Q(\reg_y[6][13] ) );
  dff_sg \reg_y_reg[6][12]  ( .D(n1544), .CP(clk), .Q(\reg_y[6][12] ) );
  dff_sg \reg_y_reg[6][11]  ( .D(n1545), .CP(clk), .Q(\reg_y[6][11] ) );
  dff_sg \reg_y_reg[6][10]  ( .D(n1546), .CP(clk), .Q(\reg_y[6][10] ) );
  dff_sg \reg_y_reg[6][9]  ( .D(n1547), .CP(clk), .Q(\reg_y[6][9] ) );
  dff_sg \reg_y_reg[6][8]  ( .D(n1548), .CP(clk), .Q(\reg_y[6][8] ) );
  dff_sg \reg_y_reg[6][7]  ( .D(n1549), .CP(clk), .Q(\reg_y[6][7] ) );
  dff_sg \reg_y_reg[6][6]  ( .D(n1550), .CP(clk), .Q(\reg_y[6][6] ) );
  dff_sg \reg_y_reg[6][5]  ( .D(n1551), .CP(clk), .Q(\reg_y[6][5] ) );
  dff_sg \reg_y_reg[6][4]  ( .D(n1552), .CP(clk), .Q(\reg_y[6][4] ) );
  dff_sg \reg_y_reg[6][3]  ( .D(n1553), .CP(clk), .Q(\reg_y[6][3] ) );
  dff_sg \reg_y_reg[6][2]  ( .D(n1554), .CP(clk), .Q(\reg_y[6][2] ) );
  dff_sg \reg_y_reg[6][1]  ( .D(n1555), .CP(clk), .Q(\reg_y[6][1] ) );
  dff_sg \reg_y_reg[6][0]  ( .D(n1556), .CP(clk), .Q(\reg_y[6][0] ) );
  dff_sg \reg_y_reg[5][19]  ( .D(n1557), .CP(clk), .Q(\reg_y[5][19] ) );
  dff_sg \reg_y_reg[5][18]  ( .D(n1558), .CP(clk), .Q(\reg_y[5][18] ) );
  dff_sg \reg_y_reg[5][17]  ( .D(n1559), .CP(clk), .Q(\reg_y[5][17] ) );
  dff_sg \reg_y_reg[5][16]  ( .D(n1560), .CP(clk), .Q(\reg_y[5][16] ) );
  dff_sg \reg_y_reg[5][15]  ( .D(n1561), .CP(clk), .Q(\reg_y[5][15] ) );
  dff_sg \reg_y_reg[5][14]  ( .D(n1562), .CP(clk), .Q(\reg_y[5][14] ) );
  dff_sg \reg_y_reg[5][13]  ( .D(n1563), .CP(clk), .Q(\reg_y[5][13] ) );
  dff_sg \reg_y_reg[5][12]  ( .D(n1564), .CP(clk), .Q(\reg_y[5][12] ) );
  dff_sg \reg_y_reg[5][11]  ( .D(n1565), .CP(clk), .Q(\reg_y[5][11] ) );
  dff_sg \reg_y_reg[5][10]  ( .D(n1566), .CP(clk), .Q(\reg_y[5][10] ) );
  dff_sg \reg_y_reg[5][9]  ( .D(n1567), .CP(clk), .Q(\reg_y[5][9] ) );
  dff_sg \reg_y_reg[5][8]  ( .D(n1568), .CP(clk), .Q(\reg_y[5][8] ) );
  dff_sg \reg_y_reg[5][7]  ( .D(n1569), .CP(clk), .Q(\reg_y[5][7] ) );
  dff_sg \reg_y_reg[5][6]  ( .D(n1570), .CP(clk), .Q(\reg_y[5][6] ) );
  dff_sg \reg_y_reg[5][5]  ( .D(n1571), .CP(clk), .Q(\reg_y[5][5] ) );
  dff_sg \reg_y_reg[5][4]  ( .D(n1572), .CP(clk), .Q(\reg_y[5][4] ) );
  dff_sg \reg_y_reg[5][3]  ( .D(n1573), .CP(clk), .Q(\reg_y[5][3] ) );
  dff_sg \reg_y_reg[5][2]  ( .D(n1574), .CP(clk), .Q(\reg_y[5][2] ) );
  dff_sg \reg_y_reg[5][1]  ( .D(n1575), .CP(clk), .Q(\reg_y[5][1] ) );
  dff_sg \reg_y_reg[5][0]  ( .D(n1576), .CP(clk), .Q(\reg_y[5][0] ) );
  dff_sg \reg_y_reg[4][19]  ( .D(n1577), .CP(clk), .Q(\reg_y[4][19] ) );
  dff_sg \reg_y_reg[4][18]  ( .D(n1578), .CP(clk), .Q(\reg_y[4][18] ) );
  dff_sg \reg_y_reg[4][17]  ( .D(n1579), .CP(clk), .Q(\reg_y[4][17] ) );
  dff_sg \reg_y_reg[4][16]  ( .D(n1580), .CP(clk), .Q(\reg_y[4][16] ) );
  dff_sg \reg_y_reg[4][15]  ( .D(n1581), .CP(clk), .Q(\reg_y[4][15] ) );
  dff_sg \reg_y_reg[4][14]  ( .D(n1582), .CP(clk), .Q(\reg_y[4][14] ) );
  dff_sg \reg_y_reg[4][13]  ( .D(n1583), .CP(clk), .Q(\reg_y[4][13] ) );
  dff_sg \reg_y_reg[4][12]  ( .D(n1584), .CP(clk), .Q(\reg_y[4][12] ) );
  dff_sg \reg_y_reg[4][11]  ( .D(n1585), .CP(clk), .Q(\reg_y[4][11] ) );
  dff_sg \reg_y_reg[4][10]  ( .D(n1586), .CP(clk), .Q(\reg_y[4][10] ) );
  dff_sg \reg_y_reg[4][9]  ( .D(n1587), .CP(clk), .Q(\reg_y[4][9] ) );
  dff_sg \reg_y_reg[4][8]  ( .D(n1588), .CP(clk), .Q(\reg_y[4][8] ) );
  dff_sg \reg_y_reg[4][7]  ( .D(n1589), .CP(clk), .Q(\reg_y[4][7] ) );
  dff_sg \reg_y_reg[4][6]  ( .D(n1590), .CP(clk), .Q(\reg_y[4][6] ) );
  dff_sg \reg_y_reg[4][5]  ( .D(n1591), .CP(clk), .Q(\reg_y[4][5] ) );
  dff_sg \reg_y_reg[4][4]  ( .D(n1592), .CP(clk), .Q(\reg_y[4][4] ) );
  dff_sg \reg_y_reg[4][3]  ( .D(n1593), .CP(clk), .Q(\reg_y[4][3] ) );
  dff_sg \reg_y_reg[4][2]  ( .D(n1594), .CP(clk), .Q(\reg_y[4][2] ) );
  dff_sg \reg_y_reg[4][1]  ( .D(n1595), .CP(clk), .Q(\reg_y[4][1] ) );
  dff_sg \reg_y_reg[4][0]  ( .D(n1596), .CP(clk), .Q(\reg_y[4][0] ) );
  dff_sg \reg_y_reg[3][19]  ( .D(n1597), .CP(clk), .Q(\reg_y[3][19] ) );
  dff_sg \reg_y_reg[3][18]  ( .D(n1598), .CP(clk), .Q(\reg_y[3][18] ) );
  dff_sg \reg_y_reg[3][17]  ( .D(n1599), .CP(clk), .Q(\reg_y[3][17] ) );
  dff_sg \reg_y_reg[3][16]  ( .D(n1600), .CP(clk), .Q(\reg_y[3][16] ) );
  dff_sg \reg_y_reg[3][15]  ( .D(n1601), .CP(clk), .Q(\reg_y[3][15] ) );
  dff_sg \reg_y_reg[3][14]  ( .D(n1602), .CP(clk), .Q(\reg_y[3][14] ) );
  dff_sg \reg_y_reg[3][13]  ( .D(n1603), .CP(clk), .Q(\reg_y[3][13] ) );
  dff_sg \reg_y_reg[3][12]  ( .D(n1604), .CP(clk), .Q(\reg_y[3][12] ) );
  dff_sg \reg_y_reg[3][11]  ( .D(n1605), .CP(clk), .Q(\reg_y[3][11] ) );
  dff_sg \reg_y_reg[3][10]  ( .D(n1606), .CP(clk), .Q(\reg_y[3][10] ) );
  dff_sg \reg_y_reg[3][9]  ( .D(n1607), .CP(clk), .Q(\reg_y[3][9] ) );
  dff_sg \reg_y_reg[3][8]  ( .D(n1608), .CP(clk), .Q(\reg_y[3][8] ) );
  dff_sg \reg_y_reg[3][7]  ( .D(n1609), .CP(clk), .Q(\reg_y[3][7] ) );
  dff_sg \reg_y_reg[3][6]  ( .D(n1610), .CP(clk), .Q(\reg_y[3][6] ) );
  dff_sg \reg_y_reg[3][5]  ( .D(n1611), .CP(clk), .Q(\reg_y[3][5] ) );
  dff_sg \reg_y_reg[3][4]  ( .D(n1612), .CP(clk), .Q(\reg_y[3][4] ) );
  dff_sg \reg_y_reg[3][3]  ( .D(n1613), .CP(clk), .Q(\reg_y[3][3] ) );
  dff_sg \reg_y_reg[3][2]  ( .D(n1614), .CP(clk), .Q(\reg_y[3][2] ) );
  dff_sg \reg_y_reg[3][1]  ( .D(n1615), .CP(clk), .Q(\reg_y[3][1] ) );
  dff_sg \reg_y_reg[3][0]  ( .D(n1616), .CP(clk), .Q(\reg_y[3][0] ) );
  dff_sg \reg_y_reg[2][19]  ( .D(n1617), .CP(clk), .Q(\reg_y[2][19] ) );
  dff_sg \reg_y_reg[2][18]  ( .D(n1618), .CP(clk), .Q(\reg_y[2][18] ) );
  dff_sg \reg_y_reg[2][17]  ( .D(n1619), .CP(clk), .Q(\reg_y[2][17] ) );
  dff_sg \reg_y_reg[2][16]  ( .D(n1620), .CP(clk), .Q(\reg_y[2][16] ) );
  dff_sg \reg_y_reg[2][15]  ( .D(n1621), .CP(clk), .Q(\reg_y[2][15] ) );
  dff_sg \reg_y_reg[2][14]  ( .D(n1622), .CP(clk), .Q(\reg_y[2][14] ) );
  dff_sg \reg_y_reg[2][13]  ( .D(n1623), .CP(clk), .Q(\reg_y[2][13] ) );
  dff_sg \reg_y_reg[2][12]  ( .D(n1624), .CP(clk), .Q(\reg_y[2][12] ) );
  dff_sg \reg_y_reg[2][11]  ( .D(n1625), .CP(clk), .Q(\reg_y[2][11] ) );
  dff_sg \reg_y_reg[2][10]  ( .D(n1626), .CP(clk), .Q(\reg_y[2][10] ) );
  dff_sg \reg_y_reg[2][9]  ( .D(n1627), .CP(clk), .Q(\reg_y[2][9] ) );
  dff_sg \reg_y_reg[2][8]  ( .D(n1628), .CP(clk), .Q(\reg_y[2][8] ) );
  dff_sg \reg_y_reg[2][7]  ( .D(n1629), .CP(clk), .Q(\reg_y[2][7] ) );
  dff_sg \reg_y_reg[2][6]  ( .D(n1630), .CP(clk), .Q(\reg_y[2][6] ) );
  dff_sg \reg_y_reg[2][5]  ( .D(n1631), .CP(clk), .Q(\reg_y[2][5] ) );
  dff_sg \reg_y_reg[2][4]  ( .D(n1632), .CP(clk), .Q(\reg_y[2][4] ) );
  dff_sg \reg_y_reg[2][3]  ( .D(n1633), .CP(clk), .Q(\reg_y[2][3] ) );
  dff_sg \reg_y_reg[2][2]  ( .D(n1634), .CP(clk), .Q(\reg_y[2][2] ) );
  dff_sg \reg_y_reg[2][1]  ( .D(n1635), .CP(clk), .Q(\reg_y[2][1] ) );
  dff_sg \reg_y_reg[2][0]  ( .D(n1636), .CP(clk), .Q(\reg_y[2][0] ) );
  dff_sg \reg_y_reg[1][19]  ( .D(n1637), .CP(clk), .Q(\reg_y[1][19] ) );
  dff_sg \reg_y_reg[1][18]  ( .D(n1638), .CP(clk), .Q(\reg_y[1][18] ) );
  dff_sg \reg_y_reg[1][17]  ( .D(n1639), .CP(clk), .Q(\reg_y[1][17] ) );
  dff_sg \reg_y_reg[1][16]  ( .D(n1640), .CP(clk), .Q(\reg_y[1][16] ) );
  dff_sg \reg_y_reg[1][15]  ( .D(n1641), .CP(clk), .Q(\reg_y[1][15] ) );
  dff_sg \reg_y_reg[1][14]  ( .D(n1642), .CP(clk), .Q(\reg_y[1][14] ) );
  dff_sg \reg_y_reg[1][13]  ( .D(n1643), .CP(clk), .Q(\reg_y[1][13] ) );
  dff_sg \reg_y_reg[1][12]  ( .D(n1644), .CP(clk), .Q(\reg_y[1][12] ) );
  dff_sg \reg_y_reg[1][11]  ( .D(n1645), .CP(clk), .Q(\reg_y[1][11] ) );
  dff_sg \reg_y_reg[1][10]  ( .D(n1646), .CP(clk), .Q(\reg_y[1][10] ) );
  dff_sg \reg_y_reg[1][9]  ( .D(n1647), .CP(clk), .Q(\reg_y[1][9] ) );
  dff_sg \reg_y_reg[1][8]  ( .D(n1648), .CP(clk), .Q(\reg_y[1][8] ) );
  dff_sg \reg_y_reg[1][7]  ( .D(n1649), .CP(clk), .Q(\reg_y[1][7] ) );
  dff_sg \reg_y_reg[1][6]  ( .D(n1650), .CP(clk), .Q(\reg_y[1][6] ) );
  dff_sg \reg_y_reg[1][5]  ( .D(n1651), .CP(clk), .Q(\reg_y[1][5] ) );
  dff_sg \reg_y_reg[1][4]  ( .D(n1652), .CP(clk), .Q(\reg_y[1][4] ) );
  dff_sg \reg_y_reg[1][3]  ( .D(n1653), .CP(clk), .Q(\reg_y[1][3] ) );
  dff_sg \reg_y_reg[1][2]  ( .D(n1654), .CP(clk), .Q(\reg_y[1][2] ) );
  dff_sg \reg_y_reg[1][1]  ( .D(n1655), .CP(clk), .Q(\reg_y[1][1] ) );
  dff_sg \reg_y_reg[1][0]  ( .D(n1656), .CP(clk), .Q(\reg_y[1][0] ) );
  dff_sg \reg_y_reg[0][19]  ( .D(n1657), .CP(clk), .Q(\reg_y[0][19] ) );
  dff_sg \reg_y_reg[0][18]  ( .D(n1658), .CP(clk), .Q(\reg_y[0][18] ) );
  dff_sg \reg_y_reg[0][17]  ( .D(n1659), .CP(clk), .Q(\reg_y[0][17] ) );
  dff_sg \reg_y_reg[0][16]  ( .D(n1660), .CP(clk), .Q(\reg_y[0][16] ) );
  dff_sg \reg_y_reg[0][15]  ( .D(n1661), .CP(clk), .Q(\reg_y[0][15] ) );
  dff_sg \reg_y_reg[0][14]  ( .D(n1662), .CP(clk), .Q(\reg_y[0][14] ) );
  dff_sg \reg_y_reg[0][13]  ( .D(n1663), .CP(clk), .Q(\reg_y[0][13] ) );
  dff_sg \reg_y_reg[0][12]  ( .D(n1664), .CP(clk), .Q(\reg_y[0][12] ) );
  dff_sg \reg_y_reg[0][11]  ( .D(n1665), .CP(clk), .Q(\reg_y[0][11] ) );
  dff_sg \reg_y_reg[0][10]  ( .D(n1666), .CP(clk), .Q(\reg_y[0][10] ) );
  dff_sg \reg_y_reg[0][9]  ( .D(n1667), .CP(clk), .Q(\reg_y[0][9] ) );
  dff_sg \reg_y_reg[0][8]  ( .D(n1668), .CP(clk), .Q(\reg_y[0][8] ) );
  dff_sg \reg_y_reg[0][7]  ( .D(n1669), .CP(clk), .Q(\reg_y[0][7] ) );
  dff_sg \reg_y_reg[0][6]  ( .D(n1670), .CP(clk), .Q(\reg_y[0][6] ) );
  dff_sg \reg_y_reg[0][5]  ( .D(n1671), .CP(clk), .Q(\reg_y[0][5] ) );
  dff_sg \reg_y_reg[0][4]  ( .D(n1672), .CP(clk), .Q(\reg_y[0][4] ) );
  dff_sg \reg_y_reg[0][3]  ( .D(n1673), .CP(clk), .Q(\reg_y[0][3] ) );
  dff_sg \reg_y_reg[0][2]  ( .D(n1674), .CP(clk), .Q(\reg_y[0][2] ) );
  dff_sg \reg_y_reg[0][1]  ( .D(n1675), .CP(clk), .Q(\reg_y[0][1] ) );
  dff_sg \reg_y_reg[0][0]  ( .D(n1676), .CP(clk), .Q(\reg_y[0][0] ) );
  dff_sg \reg_yHat_reg[14][19]  ( .D(n1697), .CP(clk), .Q(\reg_yHat[14][19] )
         );
  dff_sg \reg_yHat_reg[14][18]  ( .D(n1698), .CP(clk), .Q(\reg_yHat[14][18] )
         );
  dff_sg \reg_yHat_reg[14][17]  ( .D(n1699), .CP(clk), .Q(\reg_yHat[14][17] )
         );
  dff_sg \reg_yHat_reg[14][16]  ( .D(n1700), .CP(clk), .Q(\reg_yHat[14][16] )
         );
  dff_sg \reg_yHat_reg[14][15]  ( .D(n1701), .CP(clk), .Q(\reg_yHat[14][15] )
         );
  dff_sg \reg_yHat_reg[14][14]  ( .D(n1702), .CP(clk), .Q(\reg_yHat[14][14] )
         );
  dff_sg \reg_yHat_reg[14][13]  ( .D(n1703), .CP(clk), .Q(\reg_yHat[14][13] )
         );
  dff_sg \reg_yHat_reg[14][12]  ( .D(n1704), .CP(clk), .Q(\reg_yHat[14][12] )
         );
  dff_sg \reg_yHat_reg[14][11]  ( .D(n1705), .CP(clk), .Q(\reg_yHat[14][11] )
         );
  dff_sg \reg_yHat_reg[14][10]  ( .D(n1706), .CP(clk), .Q(\reg_yHat[14][10] )
         );
  dff_sg \reg_yHat_reg[14][9]  ( .D(n1707), .CP(clk), .Q(\reg_yHat[14][9] ) );
  dff_sg \reg_yHat_reg[14][8]  ( .D(n1708), .CP(clk), .Q(\reg_yHat[14][8] ) );
  dff_sg \reg_yHat_reg[14][7]  ( .D(n1709), .CP(clk), .Q(\reg_yHat[14][7] ) );
  dff_sg \reg_yHat_reg[14][6]  ( .D(n1710), .CP(clk), .Q(\reg_yHat[14][6] ) );
  dff_sg \reg_yHat_reg[14][5]  ( .D(n1711), .CP(clk), .Q(\reg_yHat[14][5] ) );
  dff_sg \reg_yHat_reg[14][4]  ( .D(n1712), .CP(clk), .Q(\reg_yHat[14][4] ) );
  dff_sg \reg_yHat_reg[14][3]  ( .D(n1713), .CP(clk), .Q(\reg_yHat[14][3] ) );
  dff_sg \reg_yHat_reg[14][2]  ( .D(n1714), .CP(clk), .Q(\reg_yHat[14][2] ) );
  dff_sg \reg_yHat_reg[14][1]  ( .D(n1715), .CP(clk), .Q(\reg_yHat[14][1] ) );
  dff_sg \reg_yHat_reg[14][0]  ( .D(n1716), .CP(clk), .Q(\reg_yHat[14][0] ) );
  dff_sg \reg_yHat_reg[13][19]  ( .D(n1717), .CP(clk), .Q(\reg_yHat[13][19] )
         );
  dff_sg \reg_yHat_reg[13][18]  ( .D(n1718), .CP(clk), .Q(\reg_yHat[13][18] )
         );
  dff_sg \reg_yHat_reg[13][17]  ( .D(n1719), .CP(clk), .Q(\reg_yHat[13][17] )
         );
  dff_sg \reg_yHat_reg[13][16]  ( .D(n1720), .CP(clk), .Q(\reg_yHat[13][16] )
         );
  dff_sg \reg_yHat_reg[13][15]  ( .D(n1721), .CP(clk), .Q(\reg_yHat[13][15] )
         );
  dff_sg \reg_yHat_reg[13][14]  ( .D(n1722), .CP(clk), .Q(\reg_yHat[13][14] )
         );
  dff_sg \reg_yHat_reg[13][13]  ( .D(n1723), .CP(clk), .Q(\reg_yHat[13][13] )
         );
  dff_sg \reg_yHat_reg[13][12]  ( .D(n1724), .CP(clk), .Q(\reg_yHat[13][12] )
         );
  dff_sg \reg_yHat_reg[13][11]  ( .D(n1725), .CP(clk), .Q(\reg_yHat[13][11] )
         );
  dff_sg \reg_yHat_reg[13][10]  ( .D(n1726), .CP(clk), .Q(\reg_yHat[13][10] )
         );
  dff_sg \reg_yHat_reg[13][9]  ( .D(n1727), .CP(clk), .Q(\reg_yHat[13][9] ) );
  dff_sg \reg_yHat_reg[13][8]  ( .D(n1728), .CP(clk), .Q(\reg_yHat[13][8] ) );
  dff_sg \reg_yHat_reg[13][7]  ( .D(n1729), .CP(clk), .Q(\reg_yHat[13][7] ) );
  dff_sg \reg_yHat_reg[13][6]  ( .D(n1730), .CP(clk), .Q(\reg_yHat[13][6] ) );
  dff_sg \reg_yHat_reg[13][5]  ( .D(n1731), .CP(clk), .Q(\reg_yHat[13][5] ) );
  dff_sg \reg_yHat_reg[13][4]  ( .D(n1732), .CP(clk), .Q(\reg_yHat[13][4] ) );
  dff_sg \reg_yHat_reg[13][3]  ( .D(n1733), .CP(clk), .Q(\reg_yHat[13][3] ) );
  dff_sg \reg_yHat_reg[13][2]  ( .D(n1734), .CP(clk), .Q(\reg_yHat[13][2] ) );
  dff_sg \reg_yHat_reg[13][1]  ( .D(n1735), .CP(clk), .Q(\reg_yHat[13][1] ) );
  dff_sg \reg_yHat_reg[13][0]  ( .D(n1736), .CP(clk), .Q(\reg_yHat[13][0] ) );
  dff_sg \reg_yHat_reg[12][19]  ( .D(n1737), .CP(clk), .Q(\reg_yHat[12][19] )
         );
  dff_sg \reg_yHat_reg[12][18]  ( .D(n1738), .CP(clk), .Q(\reg_yHat[12][18] )
         );
  dff_sg \reg_yHat_reg[12][17]  ( .D(n1739), .CP(clk), .Q(\reg_yHat[12][17] )
         );
  dff_sg \reg_yHat_reg[12][16]  ( .D(n1740), .CP(clk), .Q(\reg_yHat[12][16] )
         );
  dff_sg \reg_yHat_reg[12][15]  ( .D(n1741), .CP(clk), .Q(\reg_yHat[12][15] )
         );
  dff_sg \reg_yHat_reg[12][14]  ( .D(n1742), .CP(clk), .Q(\reg_yHat[12][14] )
         );
  dff_sg \reg_yHat_reg[12][13]  ( .D(n1743), .CP(clk), .Q(\reg_yHat[12][13] )
         );
  dff_sg \reg_yHat_reg[12][12]  ( .D(n1744), .CP(clk), .Q(\reg_yHat[12][12] )
         );
  dff_sg \reg_yHat_reg[12][11]  ( .D(n1745), .CP(clk), .Q(\reg_yHat[12][11] )
         );
  dff_sg \reg_yHat_reg[12][10]  ( .D(n1746), .CP(clk), .Q(\reg_yHat[12][10] )
         );
  dff_sg \reg_yHat_reg[12][9]  ( .D(n1747), .CP(clk), .Q(\reg_yHat[12][9] ) );
  dff_sg \reg_yHat_reg[12][8]  ( .D(n1748), .CP(clk), .Q(\reg_yHat[12][8] ) );
  dff_sg \reg_yHat_reg[12][7]  ( .D(n1749), .CP(clk), .Q(\reg_yHat[12][7] ) );
  dff_sg \reg_yHat_reg[12][6]  ( .D(n1750), .CP(clk), .Q(\reg_yHat[12][6] ) );
  dff_sg \reg_yHat_reg[12][5]  ( .D(n1751), .CP(clk), .Q(\reg_yHat[12][5] ) );
  dff_sg \reg_yHat_reg[12][4]  ( .D(n1752), .CP(clk), .Q(\reg_yHat[12][4] ) );
  dff_sg \reg_yHat_reg[12][3]  ( .D(n1753), .CP(clk), .Q(\reg_yHat[12][3] ) );
  dff_sg \reg_yHat_reg[12][2]  ( .D(n1754), .CP(clk), .Q(\reg_yHat[12][2] ) );
  dff_sg \reg_yHat_reg[12][1]  ( .D(n1755), .CP(clk), .Q(\reg_yHat[12][1] ) );
  dff_sg \reg_yHat_reg[12][0]  ( .D(n1756), .CP(clk), .Q(\reg_yHat[12][0] ) );
  dff_sg \reg_yHat_reg[11][19]  ( .D(n1757), .CP(clk), .Q(\reg_yHat[11][19] )
         );
  dff_sg \reg_yHat_reg[11][18]  ( .D(n1758), .CP(clk), .Q(\reg_yHat[11][18] )
         );
  dff_sg \reg_yHat_reg[11][17]  ( .D(n1759), .CP(clk), .Q(\reg_yHat[11][17] )
         );
  dff_sg \reg_yHat_reg[11][16]  ( .D(n1760), .CP(clk), .Q(\reg_yHat[11][16] )
         );
  dff_sg \reg_yHat_reg[11][15]  ( .D(n1761), .CP(clk), .Q(\reg_yHat[11][15] )
         );
  dff_sg \reg_yHat_reg[11][14]  ( .D(n1762), .CP(clk), .Q(\reg_yHat[11][14] )
         );
  dff_sg \reg_yHat_reg[11][13]  ( .D(n1763), .CP(clk), .Q(\reg_yHat[11][13] )
         );
  dff_sg \reg_yHat_reg[11][12]  ( .D(n1764), .CP(clk), .Q(\reg_yHat[11][12] )
         );
  dff_sg \reg_yHat_reg[11][11]  ( .D(n1765), .CP(clk), .Q(\reg_yHat[11][11] )
         );
  dff_sg \reg_yHat_reg[11][10]  ( .D(n1766), .CP(clk), .Q(\reg_yHat[11][10] )
         );
  dff_sg \reg_yHat_reg[11][9]  ( .D(n1767), .CP(clk), .Q(\reg_yHat[11][9] ) );
  dff_sg \reg_yHat_reg[11][8]  ( .D(n1768), .CP(clk), .Q(\reg_yHat[11][8] ) );
  dff_sg \reg_yHat_reg[11][7]  ( .D(n1769), .CP(clk), .Q(\reg_yHat[11][7] ) );
  dff_sg \reg_yHat_reg[11][6]  ( .D(n1770), .CP(clk), .Q(\reg_yHat[11][6] ) );
  dff_sg \reg_yHat_reg[11][5]  ( .D(n1771), .CP(clk), .Q(\reg_yHat[11][5] ) );
  dff_sg \reg_yHat_reg[11][4]  ( .D(n1772), .CP(clk), .Q(\reg_yHat[11][4] ) );
  dff_sg \reg_yHat_reg[11][3]  ( .D(n1773), .CP(clk), .Q(\reg_yHat[11][3] ) );
  dff_sg \reg_yHat_reg[11][2]  ( .D(n1774), .CP(clk), .Q(\reg_yHat[11][2] ) );
  dff_sg \reg_yHat_reg[11][1]  ( .D(n1775), .CP(clk), .Q(\reg_yHat[11][1] ) );
  dff_sg \reg_yHat_reg[11][0]  ( .D(n1776), .CP(clk), .Q(\reg_yHat[11][0] ) );
  dff_sg \reg_yHat_reg[10][19]  ( .D(n1777), .CP(clk), .Q(\reg_yHat[10][19] )
         );
  dff_sg \reg_yHat_reg[10][18]  ( .D(n1778), .CP(clk), .Q(\reg_yHat[10][18] )
         );
  dff_sg \reg_yHat_reg[10][17]  ( .D(n1779), .CP(clk), .Q(\reg_yHat[10][17] )
         );
  dff_sg \reg_yHat_reg[10][16]  ( .D(n1780), .CP(clk), .Q(\reg_yHat[10][16] )
         );
  dff_sg \reg_yHat_reg[10][15]  ( .D(n1781), .CP(clk), .Q(\reg_yHat[10][15] )
         );
  dff_sg \reg_yHat_reg[10][14]  ( .D(n1782), .CP(clk), .Q(\reg_yHat[10][14] )
         );
  dff_sg \reg_yHat_reg[10][13]  ( .D(n1783), .CP(clk), .Q(\reg_yHat[10][13] )
         );
  dff_sg \reg_yHat_reg[10][12]  ( .D(n1784), .CP(clk), .Q(\reg_yHat[10][12] )
         );
  dff_sg \reg_yHat_reg[10][11]  ( .D(n1785), .CP(clk), .Q(\reg_yHat[10][11] )
         );
  dff_sg \reg_yHat_reg[10][10]  ( .D(n1786), .CP(clk), .Q(\reg_yHat[10][10] )
         );
  dff_sg \reg_yHat_reg[10][9]  ( .D(n1787), .CP(clk), .Q(\reg_yHat[10][9] ) );
  dff_sg \reg_yHat_reg[10][8]  ( .D(n1788), .CP(clk), .Q(\reg_yHat[10][8] ) );
  dff_sg \reg_yHat_reg[10][7]  ( .D(n1789), .CP(clk), .Q(\reg_yHat[10][7] ) );
  dff_sg \reg_yHat_reg[10][6]  ( .D(n1790), .CP(clk), .Q(\reg_yHat[10][6] ) );
  dff_sg \reg_yHat_reg[10][5]  ( .D(n1791), .CP(clk), .Q(\reg_yHat[10][5] ) );
  dff_sg \reg_yHat_reg[10][4]  ( .D(n1792), .CP(clk), .Q(\reg_yHat[10][4] ) );
  dff_sg \reg_yHat_reg[10][3]  ( .D(n1793), .CP(clk), .Q(\reg_yHat[10][3] ) );
  dff_sg \reg_yHat_reg[10][2]  ( .D(n1794), .CP(clk), .Q(\reg_yHat[10][2] ) );
  dff_sg \reg_yHat_reg[10][1]  ( .D(n1795), .CP(clk), .Q(\reg_yHat[10][1] ) );
  dff_sg \reg_yHat_reg[10][0]  ( .D(n1796), .CP(clk), .Q(\reg_yHat[10][0] ) );
  dff_sg \reg_yHat_reg[9][19]  ( .D(n1797), .CP(clk), .Q(\reg_yHat[9][19] ) );
  dff_sg \reg_yHat_reg[9][18]  ( .D(n1798), .CP(clk), .Q(\reg_yHat[9][18] ) );
  dff_sg \reg_yHat_reg[9][17]  ( .D(n1799), .CP(clk), .Q(\reg_yHat[9][17] ) );
  dff_sg \reg_yHat_reg[9][16]  ( .D(n1800), .CP(clk), .Q(\reg_yHat[9][16] ) );
  dff_sg \reg_yHat_reg[9][15]  ( .D(n1801), .CP(clk), .Q(\reg_yHat[9][15] ) );
  dff_sg \reg_yHat_reg[9][14]  ( .D(n1802), .CP(clk), .Q(\reg_yHat[9][14] ) );
  dff_sg \reg_yHat_reg[9][13]  ( .D(n1803), .CP(clk), .Q(\reg_yHat[9][13] ) );
  dff_sg \reg_yHat_reg[9][12]  ( .D(n1804), .CP(clk), .Q(\reg_yHat[9][12] ) );
  dff_sg \reg_yHat_reg[9][11]  ( .D(n1805), .CP(clk), .Q(\reg_yHat[9][11] ) );
  dff_sg \reg_yHat_reg[9][10]  ( .D(n1806), .CP(clk), .Q(\reg_yHat[9][10] ) );
  dff_sg \reg_yHat_reg[9][9]  ( .D(n1807), .CP(clk), .Q(\reg_yHat[9][9] ) );
  dff_sg \reg_yHat_reg[9][8]  ( .D(n1808), .CP(clk), .Q(\reg_yHat[9][8] ) );
  dff_sg \reg_yHat_reg[9][7]  ( .D(n1809), .CP(clk), .Q(\reg_yHat[9][7] ) );
  dff_sg \reg_yHat_reg[9][6]  ( .D(n1810), .CP(clk), .Q(\reg_yHat[9][6] ) );
  dff_sg \reg_yHat_reg[9][5]  ( .D(n1811), .CP(clk), .Q(\reg_yHat[9][5] ) );
  dff_sg \reg_yHat_reg[9][4]  ( .D(n1812), .CP(clk), .Q(\reg_yHat[9][4] ) );
  dff_sg \reg_yHat_reg[9][3]  ( .D(n1813), .CP(clk), .Q(\reg_yHat[9][3] ) );
  dff_sg \reg_yHat_reg[9][2]  ( .D(n1814), .CP(clk), .Q(\reg_yHat[9][2] ) );
  dff_sg \reg_yHat_reg[9][1]  ( .D(n1815), .CP(clk), .Q(\reg_yHat[9][1] ) );
  dff_sg \reg_yHat_reg[9][0]  ( .D(n1816), .CP(clk), .Q(\reg_yHat[9][0] ) );
  dff_sg \reg_yHat_reg[8][19]  ( .D(n1817), .CP(clk), .Q(\reg_yHat[8][19] ) );
  dff_sg \reg_yHat_reg[8][18]  ( .D(n1818), .CP(clk), .Q(\reg_yHat[8][18] ) );
  dff_sg \reg_yHat_reg[8][17]  ( .D(n1819), .CP(clk), .Q(\reg_yHat[8][17] ) );
  dff_sg \reg_yHat_reg[8][16]  ( .D(n1820), .CP(clk), .Q(\reg_yHat[8][16] ) );
  dff_sg \reg_yHat_reg[8][15]  ( .D(n1821), .CP(clk), .Q(\reg_yHat[8][15] ) );
  dff_sg \reg_yHat_reg[8][14]  ( .D(n1822), .CP(clk), .Q(\reg_yHat[8][14] ) );
  dff_sg \reg_yHat_reg[8][13]  ( .D(n1823), .CP(clk), .Q(\reg_yHat[8][13] ) );
  dff_sg \reg_yHat_reg[8][12]  ( .D(n1824), .CP(clk), .Q(\reg_yHat[8][12] ) );
  dff_sg \reg_yHat_reg[8][11]  ( .D(n1825), .CP(clk), .Q(\reg_yHat[8][11] ) );
  dff_sg \reg_yHat_reg[8][10]  ( .D(n1826), .CP(clk), .Q(\reg_yHat[8][10] ) );
  dff_sg \reg_yHat_reg[8][9]  ( .D(n1827), .CP(clk), .Q(\reg_yHat[8][9] ) );
  dff_sg \reg_yHat_reg[8][8]  ( .D(n1828), .CP(clk), .Q(\reg_yHat[8][8] ) );
  dff_sg \reg_yHat_reg[8][7]  ( .D(n1829), .CP(clk), .Q(\reg_yHat[8][7] ) );
  dff_sg \reg_yHat_reg[8][6]  ( .D(n1830), .CP(clk), .Q(\reg_yHat[8][6] ) );
  dff_sg \reg_yHat_reg[8][5]  ( .D(n1831), .CP(clk), .Q(\reg_yHat[8][5] ) );
  dff_sg \reg_yHat_reg[8][4]  ( .D(n1832), .CP(clk), .Q(\reg_yHat[8][4] ) );
  dff_sg \reg_yHat_reg[8][3]  ( .D(n1833), .CP(clk), .Q(\reg_yHat[8][3] ) );
  dff_sg \reg_yHat_reg[8][2]  ( .D(n1834), .CP(clk), .Q(\reg_yHat[8][2] ) );
  dff_sg \reg_yHat_reg[8][1]  ( .D(n1835), .CP(clk), .Q(\reg_yHat[8][1] ) );
  dff_sg \reg_yHat_reg[8][0]  ( .D(n1836), .CP(clk), .Q(\reg_yHat[8][0] ) );
  dff_sg \reg_yHat_reg[7][19]  ( .D(n1837), .CP(clk), .Q(\reg_yHat[7][19] ) );
  dff_sg \reg_yHat_reg[7][18]  ( .D(n1838), .CP(clk), .Q(\reg_yHat[7][18] ) );
  dff_sg \reg_yHat_reg[7][17]  ( .D(n1839), .CP(clk), .Q(\reg_yHat[7][17] ) );
  dff_sg \reg_yHat_reg[7][16]  ( .D(n1840), .CP(clk), .Q(\reg_yHat[7][16] ) );
  dff_sg \reg_yHat_reg[7][15]  ( .D(n1841), .CP(clk), .Q(\reg_yHat[7][15] ) );
  dff_sg \reg_yHat_reg[7][14]  ( .D(n1842), .CP(clk), .Q(\reg_yHat[7][14] ) );
  dff_sg \reg_yHat_reg[7][13]  ( .D(n1843), .CP(clk), .Q(\reg_yHat[7][13] ) );
  dff_sg \reg_yHat_reg[7][12]  ( .D(n1844), .CP(clk), .Q(\reg_yHat[7][12] ) );
  dff_sg \reg_yHat_reg[7][11]  ( .D(n1845), .CP(clk), .Q(\reg_yHat[7][11] ) );
  dff_sg \reg_yHat_reg[7][10]  ( .D(n1846), .CP(clk), .Q(\reg_yHat[7][10] ) );
  dff_sg \reg_yHat_reg[7][9]  ( .D(n1847), .CP(clk), .Q(\reg_yHat[7][9] ) );
  dff_sg \reg_yHat_reg[7][8]  ( .D(n1848), .CP(clk), .Q(\reg_yHat[7][8] ) );
  dff_sg \reg_yHat_reg[7][7]  ( .D(n1849), .CP(clk), .Q(\reg_yHat[7][7] ) );
  dff_sg \reg_yHat_reg[7][6]  ( .D(n1850), .CP(clk), .Q(\reg_yHat[7][6] ) );
  dff_sg \reg_yHat_reg[7][5]  ( .D(n1851), .CP(clk), .Q(\reg_yHat[7][5] ) );
  dff_sg \reg_yHat_reg[7][4]  ( .D(n1852), .CP(clk), .Q(\reg_yHat[7][4] ) );
  dff_sg \reg_yHat_reg[7][3]  ( .D(n1853), .CP(clk), .Q(\reg_yHat[7][3] ) );
  dff_sg \reg_yHat_reg[7][2]  ( .D(n1854), .CP(clk), .Q(\reg_yHat[7][2] ) );
  dff_sg \reg_yHat_reg[7][1]  ( .D(n1855), .CP(clk), .Q(\reg_yHat[7][1] ) );
  dff_sg \reg_yHat_reg[7][0]  ( .D(n1856), .CP(clk), .Q(\reg_yHat[7][0] ) );
  dff_sg \reg_yHat_reg[6][19]  ( .D(n1857), .CP(clk), .Q(\reg_yHat[6][19] ) );
  dff_sg \reg_yHat_reg[6][18]  ( .D(n1858), .CP(clk), .Q(\reg_yHat[6][18] ) );
  dff_sg \reg_yHat_reg[6][17]  ( .D(n1859), .CP(clk), .Q(\reg_yHat[6][17] ) );
  dff_sg \reg_yHat_reg[6][16]  ( .D(n1860), .CP(clk), .Q(\reg_yHat[6][16] ) );
  dff_sg \reg_yHat_reg[6][15]  ( .D(n1861), .CP(clk), .Q(\reg_yHat[6][15] ) );
  dff_sg \reg_yHat_reg[6][14]  ( .D(n1862), .CP(clk), .Q(\reg_yHat[6][14] ) );
  dff_sg \reg_yHat_reg[6][13]  ( .D(n1863), .CP(clk), .Q(\reg_yHat[6][13] ) );
  dff_sg \reg_yHat_reg[6][12]  ( .D(n1864), .CP(clk), .Q(\reg_yHat[6][12] ) );
  dff_sg \reg_yHat_reg[6][11]  ( .D(n1865), .CP(clk), .Q(\reg_yHat[6][11] ) );
  dff_sg \reg_yHat_reg[6][10]  ( .D(n1866), .CP(clk), .Q(\reg_yHat[6][10] ) );
  dff_sg \reg_yHat_reg[6][9]  ( .D(n1867), .CP(clk), .Q(\reg_yHat[6][9] ) );
  dff_sg \reg_yHat_reg[6][8]  ( .D(n1868), .CP(clk), .Q(\reg_yHat[6][8] ) );
  dff_sg \reg_yHat_reg[6][7]  ( .D(n1869), .CP(clk), .Q(\reg_yHat[6][7] ) );
  dff_sg \reg_yHat_reg[6][6]  ( .D(n1870), .CP(clk), .Q(\reg_yHat[6][6] ) );
  dff_sg \reg_yHat_reg[6][5]  ( .D(n1871), .CP(clk), .Q(\reg_yHat[6][5] ) );
  dff_sg \reg_yHat_reg[6][4]  ( .D(n1872), .CP(clk), .Q(\reg_yHat[6][4] ) );
  dff_sg \reg_yHat_reg[6][3]  ( .D(n1873), .CP(clk), .Q(\reg_yHat[6][3] ) );
  dff_sg \reg_yHat_reg[6][2]  ( .D(n1874), .CP(clk), .Q(\reg_yHat[6][2] ) );
  dff_sg \reg_yHat_reg[6][1]  ( .D(n1875), .CP(clk), .Q(\reg_yHat[6][1] ) );
  dff_sg \reg_yHat_reg[6][0]  ( .D(n1876), .CP(clk), .Q(\reg_yHat[6][0] ) );
  dff_sg \reg_yHat_reg[5][19]  ( .D(n1877), .CP(clk), .Q(\reg_yHat[5][19] ) );
  dff_sg \reg_yHat_reg[5][18]  ( .D(n1878), .CP(clk), .Q(\reg_yHat[5][18] ) );
  dff_sg \reg_yHat_reg[5][17]  ( .D(n1879), .CP(clk), .Q(\reg_yHat[5][17] ) );
  dff_sg \reg_yHat_reg[5][16]  ( .D(n1880), .CP(clk), .Q(\reg_yHat[5][16] ) );
  dff_sg \reg_yHat_reg[5][15]  ( .D(n1881), .CP(clk), .Q(\reg_yHat[5][15] ) );
  dff_sg \reg_yHat_reg[5][14]  ( .D(n1882), .CP(clk), .Q(\reg_yHat[5][14] ) );
  dff_sg \reg_yHat_reg[5][13]  ( .D(n1883), .CP(clk), .Q(\reg_yHat[5][13] ) );
  dff_sg \reg_yHat_reg[5][12]  ( .D(n1884), .CP(clk), .Q(\reg_yHat[5][12] ) );
  dff_sg \reg_yHat_reg[5][11]  ( .D(n1885), .CP(clk), .Q(\reg_yHat[5][11] ) );
  dff_sg \reg_yHat_reg[5][10]  ( .D(n1886), .CP(clk), .Q(\reg_yHat[5][10] ) );
  dff_sg \reg_yHat_reg[5][9]  ( .D(n1887), .CP(clk), .Q(\reg_yHat[5][9] ) );
  dff_sg \reg_yHat_reg[5][8]  ( .D(n1888), .CP(clk), .Q(\reg_yHat[5][8] ) );
  dff_sg \reg_yHat_reg[5][7]  ( .D(n1889), .CP(clk), .Q(\reg_yHat[5][7] ) );
  dff_sg \reg_yHat_reg[5][6]  ( .D(n1890), .CP(clk), .Q(\reg_yHat[5][6] ) );
  dff_sg \reg_yHat_reg[5][5]  ( .D(n1891), .CP(clk), .Q(\reg_yHat[5][5] ) );
  dff_sg \reg_yHat_reg[5][4]  ( .D(n1892), .CP(clk), .Q(\reg_yHat[5][4] ) );
  dff_sg \reg_yHat_reg[5][3]  ( .D(n1893), .CP(clk), .Q(\reg_yHat[5][3] ) );
  dff_sg \reg_yHat_reg[5][2]  ( .D(n1894), .CP(clk), .Q(\reg_yHat[5][2] ) );
  dff_sg \reg_yHat_reg[5][1]  ( .D(n1895), .CP(clk), .Q(\reg_yHat[5][1] ) );
  dff_sg \reg_yHat_reg[5][0]  ( .D(n1896), .CP(clk), .Q(\reg_yHat[5][0] ) );
  dff_sg \reg_yHat_reg[4][19]  ( .D(n1897), .CP(clk), .Q(\reg_yHat[4][19] ) );
  dff_sg \reg_yHat_reg[4][18]  ( .D(n1898), .CP(clk), .Q(\reg_yHat[4][18] ) );
  dff_sg \reg_yHat_reg[4][17]  ( .D(n1899), .CP(clk), .Q(\reg_yHat[4][17] ) );
  dff_sg \reg_yHat_reg[4][16]  ( .D(n1900), .CP(clk), .Q(\reg_yHat[4][16] ) );
  dff_sg \reg_yHat_reg[4][15]  ( .D(n1901), .CP(clk), .Q(\reg_yHat[4][15] ) );
  dff_sg \reg_yHat_reg[4][14]  ( .D(n1902), .CP(clk), .Q(\reg_yHat[4][14] ) );
  dff_sg \reg_yHat_reg[4][13]  ( .D(n1903), .CP(clk), .Q(\reg_yHat[4][13] ) );
  dff_sg \reg_yHat_reg[4][12]  ( .D(n1904), .CP(clk), .Q(\reg_yHat[4][12] ) );
  dff_sg \reg_yHat_reg[4][11]  ( .D(n1905), .CP(clk), .Q(\reg_yHat[4][11] ) );
  dff_sg \reg_yHat_reg[4][10]  ( .D(n1906), .CP(clk), .Q(\reg_yHat[4][10] ) );
  dff_sg \reg_yHat_reg[4][9]  ( .D(n1907), .CP(clk), .Q(\reg_yHat[4][9] ) );
  dff_sg \reg_yHat_reg[4][8]  ( .D(n1908), .CP(clk), .Q(\reg_yHat[4][8] ) );
  dff_sg \reg_yHat_reg[4][7]  ( .D(n1909), .CP(clk), .Q(\reg_yHat[4][7] ) );
  dff_sg \reg_yHat_reg[4][6]  ( .D(n1910), .CP(clk), .Q(\reg_yHat[4][6] ) );
  dff_sg \reg_yHat_reg[4][5]  ( .D(n1911), .CP(clk), .Q(\reg_yHat[4][5] ) );
  dff_sg \reg_yHat_reg[4][4]  ( .D(n1912), .CP(clk), .Q(\reg_yHat[4][4] ) );
  dff_sg \reg_yHat_reg[4][3]  ( .D(n1913), .CP(clk), .Q(\reg_yHat[4][3] ) );
  dff_sg \reg_yHat_reg[4][2]  ( .D(n1914), .CP(clk), .Q(\reg_yHat[4][2] ) );
  dff_sg \reg_yHat_reg[4][1]  ( .D(n1915), .CP(clk), .Q(\reg_yHat[4][1] ) );
  dff_sg \reg_yHat_reg[4][0]  ( .D(n1916), .CP(clk), .Q(\reg_yHat[4][0] ) );
  dff_sg \reg_yHat_reg[3][19]  ( .D(n1917), .CP(clk), .Q(\reg_yHat[3][19] ) );
  dff_sg \reg_yHat_reg[3][18]  ( .D(n1918), .CP(clk), .Q(\reg_yHat[3][18] ) );
  dff_sg \reg_yHat_reg[3][17]  ( .D(n1919), .CP(clk), .Q(\reg_yHat[3][17] ) );
  dff_sg \reg_yHat_reg[3][16]  ( .D(n1920), .CP(clk), .Q(\reg_yHat[3][16] ) );
  dff_sg \reg_yHat_reg[3][15]  ( .D(n1921), .CP(clk), .Q(\reg_yHat[3][15] ) );
  dff_sg \reg_yHat_reg[3][14]  ( .D(n1922), .CP(clk), .Q(\reg_yHat[3][14] ) );
  dff_sg \reg_yHat_reg[3][13]  ( .D(n1923), .CP(clk), .Q(\reg_yHat[3][13] ) );
  dff_sg \reg_yHat_reg[3][12]  ( .D(n1924), .CP(clk), .Q(\reg_yHat[3][12] ) );
  dff_sg \reg_yHat_reg[3][11]  ( .D(n1925), .CP(clk), .Q(\reg_yHat[3][11] ) );
  dff_sg \reg_yHat_reg[3][10]  ( .D(n1926), .CP(clk), .Q(\reg_yHat[3][10] ) );
  dff_sg \reg_yHat_reg[3][9]  ( .D(n1927), .CP(clk), .Q(\reg_yHat[3][9] ) );
  dff_sg \reg_yHat_reg[3][8]  ( .D(n1928), .CP(clk), .Q(\reg_yHat[3][8] ) );
  dff_sg \reg_yHat_reg[3][7]  ( .D(n1929), .CP(clk), .Q(\reg_yHat[3][7] ) );
  dff_sg \reg_yHat_reg[3][6]  ( .D(n1930), .CP(clk), .Q(\reg_yHat[3][6] ) );
  dff_sg \reg_yHat_reg[3][5]  ( .D(n1931), .CP(clk), .Q(\reg_yHat[3][5] ) );
  dff_sg \reg_yHat_reg[3][4]  ( .D(n1932), .CP(clk), .Q(\reg_yHat[3][4] ) );
  dff_sg \reg_yHat_reg[3][3]  ( .D(n1933), .CP(clk), .Q(\reg_yHat[3][3] ) );
  dff_sg \reg_yHat_reg[3][2]  ( .D(n1934), .CP(clk), .Q(\reg_yHat[3][2] ) );
  dff_sg \reg_yHat_reg[3][1]  ( .D(n1935), .CP(clk), .Q(\reg_yHat[3][1] ) );
  dff_sg \reg_yHat_reg[3][0]  ( .D(n1936), .CP(clk), .Q(\reg_yHat[3][0] ) );
  dff_sg \reg_yHat_reg[2][19]  ( .D(n1937), .CP(clk), .Q(\reg_yHat[2][19] ) );
  dff_sg \reg_yHat_reg[2][18]  ( .D(n1938), .CP(clk), .Q(\reg_yHat[2][18] ) );
  dff_sg \reg_yHat_reg[2][17]  ( .D(n1939), .CP(clk), .Q(\reg_yHat[2][17] ) );
  dff_sg \reg_yHat_reg[2][16]  ( .D(n1940), .CP(clk), .Q(\reg_yHat[2][16] ) );
  dff_sg \reg_yHat_reg[2][15]  ( .D(n1941), .CP(clk), .Q(\reg_yHat[2][15] ) );
  dff_sg \reg_yHat_reg[2][14]  ( .D(n1942), .CP(clk), .Q(\reg_yHat[2][14] ) );
  dff_sg \reg_yHat_reg[2][13]  ( .D(n1943), .CP(clk), .Q(\reg_yHat[2][13] ) );
  dff_sg \reg_yHat_reg[2][12]  ( .D(n1944), .CP(clk), .Q(\reg_yHat[2][12] ) );
  dff_sg \reg_yHat_reg[2][11]  ( .D(n1945), .CP(clk), .Q(\reg_yHat[2][11] ) );
  dff_sg \reg_yHat_reg[2][10]  ( .D(n1946), .CP(clk), .Q(\reg_yHat[2][10] ) );
  dff_sg \reg_yHat_reg[2][9]  ( .D(n1947), .CP(clk), .Q(\reg_yHat[2][9] ) );
  dff_sg \reg_yHat_reg[2][8]  ( .D(n1948), .CP(clk), .Q(\reg_yHat[2][8] ) );
  dff_sg \reg_yHat_reg[2][7]  ( .D(n1949), .CP(clk), .Q(\reg_yHat[2][7] ) );
  dff_sg \reg_yHat_reg[2][6]  ( .D(n1950), .CP(clk), .Q(\reg_yHat[2][6] ) );
  dff_sg \reg_yHat_reg[2][5]  ( .D(n1951), .CP(clk), .Q(\reg_yHat[2][5] ) );
  dff_sg \reg_yHat_reg[2][4]  ( .D(n1952), .CP(clk), .Q(\reg_yHat[2][4] ) );
  dff_sg \reg_yHat_reg[2][3]  ( .D(n1953), .CP(clk), .Q(\reg_yHat[2][3] ) );
  dff_sg \reg_yHat_reg[2][2]  ( .D(n1954), .CP(clk), .Q(\reg_yHat[2][2] ) );
  dff_sg \reg_yHat_reg[2][1]  ( .D(n1955), .CP(clk), .Q(\reg_yHat[2][1] ) );
  dff_sg \reg_yHat_reg[2][0]  ( .D(n1956), .CP(clk), .Q(\reg_yHat[2][0] ) );
  dff_sg \reg_yHat_reg[1][19]  ( .D(n1957), .CP(clk), .Q(\reg_yHat[1][19] ) );
  dff_sg \reg_yHat_reg[1][18]  ( .D(n1958), .CP(clk), .Q(\reg_yHat[1][18] ) );
  dff_sg \reg_yHat_reg[1][17]  ( .D(n1959), .CP(clk), .Q(\reg_yHat[1][17] ) );
  dff_sg \reg_yHat_reg[1][16]  ( .D(n1960), .CP(clk), .Q(\reg_yHat[1][16] ) );
  dff_sg \reg_yHat_reg[1][15]  ( .D(n1961), .CP(clk), .Q(\reg_yHat[1][15] ) );
  dff_sg \reg_yHat_reg[1][14]  ( .D(n1962), .CP(clk), .Q(\reg_yHat[1][14] ) );
  dff_sg \reg_yHat_reg[1][13]  ( .D(n1963), .CP(clk), .Q(\reg_yHat[1][13] ) );
  dff_sg \reg_yHat_reg[1][12]  ( .D(n1964), .CP(clk), .Q(\reg_yHat[1][12] ) );
  dff_sg \reg_yHat_reg[1][11]  ( .D(n1965), .CP(clk), .Q(\reg_yHat[1][11] ) );
  dff_sg \reg_yHat_reg[1][10]  ( .D(n1966), .CP(clk), .Q(\reg_yHat[1][10] ) );
  dff_sg \reg_yHat_reg[1][9]  ( .D(n1967), .CP(clk), .Q(\reg_yHat[1][9] ) );
  dff_sg \reg_yHat_reg[1][8]  ( .D(n1968), .CP(clk), .Q(\reg_yHat[1][8] ) );
  dff_sg \reg_yHat_reg[1][7]  ( .D(n1969), .CP(clk), .Q(\reg_yHat[1][7] ) );
  dff_sg \reg_yHat_reg[1][6]  ( .D(n1970), .CP(clk), .Q(\reg_yHat[1][6] ) );
  dff_sg \reg_yHat_reg[1][5]  ( .D(n1971), .CP(clk), .Q(\reg_yHat[1][5] ) );
  dff_sg \reg_yHat_reg[1][4]  ( .D(n1972), .CP(clk), .Q(\reg_yHat[1][4] ) );
  dff_sg \reg_yHat_reg[1][3]  ( .D(n1973), .CP(clk), .Q(\reg_yHat[1][3] ) );
  dff_sg \reg_yHat_reg[1][2]  ( .D(n1974), .CP(clk), .Q(\reg_yHat[1][2] ) );
  dff_sg \reg_yHat_reg[1][1]  ( .D(n1975), .CP(clk), .Q(\reg_yHat[1][1] ) );
  dff_sg \reg_yHat_reg[1][0]  ( .D(n1976), .CP(clk), .Q(\reg_yHat[1][0] ) );
  dff_sg \reg_yHat_reg[0][19]  ( .D(n1977), .CP(clk), .Q(\reg_yHat[0][19] ) );
  dff_sg \reg_yHat_reg[0][18]  ( .D(n1978), .CP(clk), .Q(\reg_yHat[0][18] ) );
  dff_sg \reg_yHat_reg[0][17]  ( .D(n1979), .CP(clk), .Q(\reg_yHat[0][17] ) );
  dff_sg \reg_yHat_reg[0][16]  ( .D(n1980), .CP(clk), .Q(\reg_yHat[0][16] ) );
  dff_sg \reg_yHat_reg[0][15]  ( .D(n1981), .CP(clk), .Q(\reg_yHat[0][15] ) );
  dff_sg \reg_yHat_reg[0][14]  ( .D(n1982), .CP(clk), .Q(\reg_yHat[0][14] ) );
  dff_sg \reg_yHat_reg[0][13]  ( .D(n1983), .CP(clk), .Q(\reg_yHat[0][13] ) );
  dff_sg \reg_yHat_reg[0][12]  ( .D(n1984), .CP(clk), .Q(\reg_yHat[0][12] ) );
  dff_sg \reg_yHat_reg[0][11]  ( .D(n1985), .CP(clk), .Q(\reg_yHat[0][11] ) );
  dff_sg \reg_yHat_reg[0][10]  ( .D(n1986), .CP(clk), .Q(\reg_yHat[0][10] ) );
  dff_sg \reg_yHat_reg[0][9]  ( .D(n1987), .CP(clk), .Q(\reg_yHat[0][9] ) );
  dff_sg \reg_yHat_reg[0][8]  ( .D(n1988), .CP(clk), .Q(\reg_yHat[0][8] ) );
  dff_sg \reg_yHat_reg[0][7]  ( .D(n1989), .CP(clk), .Q(\reg_yHat[0][7] ) );
  dff_sg \reg_yHat_reg[0][6]  ( .D(n1990), .CP(clk), .Q(\reg_yHat[0][6] ) );
  dff_sg \reg_yHat_reg[0][5]  ( .D(n1991), .CP(clk), .Q(\reg_yHat[0][5] ) );
  dff_sg \reg_yHat_reg[0][4]  ( .D(n1992), .CP(clk), .Q(\reg_yHat[0][4] ) );
  dff_sg \reg_yHat_reg[0][3]  ( .D(n1993), .CP(clk), .Q(\reg_yHat[0][3] ) );
  dff_sg \reg_yHat_reg[0][2]  ( .D(n1994), .CP(clk), .Q(\reg_yHat[0][2] ) );
  dff_sg \reg_yHat_reg[0][1]  ( .D(n1995), .CP(clk), .Q(\reg_yHat[0][1] ) );
  dff_sg \reg_yHat_reg[0][0]  ( .D(n1996), .CP(clk), .Q(\reg_yHat[0][0] ) );
  dff_sg reg_model_reg ( .D(n1997), .CP(clk), .Q(reg_model) );
  \**FFGEN**  \L1_0/abs_reg[14][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3239 ), .force_10(\L1_0/n3240 ), 
        .force_11(1'b0), .QN(n5132) );
  \**FFGEN**  \L1_0/abs_reg[14][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3243 ), .force_10(\L1_0/n3244 ), 
        .force_11(1'b0), .Q(n38455), .QN(n5133) );
  \**FFGEN**  \L1_0/abs_reg[14][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3247 ), .force_10(\L1_0/n3248 ), 
        .force_11(1'b0), .Q(n38459), .QN(n5134) );
  \**FFGEN**  \L1_0/abs_reg[14][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3251 ), .force_10(\L1_0/n3252 ), 
        .force_11(1'b0), .Q(n38463), .QN(n5135) );
  \**FFGEN**  \L1_0/abs_reg[14][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3255 ), .force_10(\L1_0/n3256 ), 
        .force_11(1'b0), .Q(n38467), .QN(n5136) );
  \**FFGEN**  \L1_0/abs_reg[14][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3259 ), .force_10(\L1_0/n3260 ), 
        .force_11(1'b0), .Q(n38471), .QN(n5137) );
  \**FFGEN**  \L1_0/abs_reg[14][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3263 ), .force_10(\L1_0/n3264 ), 
        .force_11(1'b0), .Q(n38475), .QN(n5138) );
  \**FFGEN**  \L1_0/abs_reg[14][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3267 ), .force_10(\L1_0/n3268 ), 
        .force_11(1'b0), .Q(n38479), .QN(n5139) );
  \**FFGEN**  \L1_0/abs_reg[14][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3271 ), .force_10(\L1_0/n3272 ), 
        .force_11(1'b0), .Q(n38483), .QN(n5140) );
  \**FFGEN**  \L1_0/abs_reg[14][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3275 ), .force_10(\L1_0/n3276 ), 
        .force_11(1'b0), .Q(n38487), .QN(n5141) );
  \**FFGEN**  \L1_0/abs_reg[14][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3279 ), .force_10(\L1_0/n3280 ), 
        .force_11(1'b0), .Q(n38491), .QN(n5142) );
  \**FFGEN**  \L1_0/abs_reg[14][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3283 ), .force_10(\L1_0/n3284 ), 
        .force_11(1'b0), .Q(n38495), .QN(n5143) );
  \**FFGEN**  \L1_0/abs_reg[14][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3287 ), .force_10(\L1_0/n3288 ), 
        .force_11(1'b0), .Q(n38499), .QN(n5144) );
  \**FFGEN**  \L1_0/abs_reg[14][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3291 ), .force_10(\L1_0/n3292 ), 
        .force_11(1'b0), .Q(n38503), .QN(n5145) );
  \**FFGEN**  \L1_0/abs_reg[14][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3295 ), .force_10(\L1_0/n3296 ), 
        .force_11(1'b0), .Q(n38507), .QN(n5146) );
  \**FFGEN**  \L1_0/abs_reg[14][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3299 ), .force_10(\L1_0/n3300 ), 
        .force_11(1'b0), .Q(n38511), .QN(n5147) );
  \**FFGEN**  \L1_0/abs_reg[14][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3303 ), .force_10(\L1_0/n3304 ), 
        .force_11(1'b0), .Q(n38515), .QN(n5148) );
  \**FFGEN**  \L1_0/abs_reg[14][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3307 ), .force_10(\L1_0/n3308 ), 
        .force_11(1'b0), .Q(n38280), .QN(n5149) );
  \**FFGEN**  \L1_0/abs_reg[14][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3311 ), .force_10(\L1_0/n3312 ), 
        .force_11(1'b0), .Q(n38559) );
  \**FFGEN**  \L1_0/abs_reg[14][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3315 ), .force_10(\L1_0/n3316 ), 
        .force_11(1'b0), .QN(n5717) );
  \**FFGEN**  \L1_0/abs_reg[13][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3319 ), .force_10(\L1_0/n3320 ), 
        .force_11(1'b0), .QN(n5151) );
  \**FFGEN**  \L1_0/abs_reg[13][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n51487), .force_10(\L1_0/n3324 ), 
        .force_11(1'b0), .Q(n38456), .QN(n5152) );
  \**FFGEN**  \L1_0/abs_reg[13][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n51486), .force_10(\L1_0/n3328 ), 
        .force_11(1'b0), .Q(n38460), .QN(n5153) );
  \**FFGEN**  \L1_0/abs_reg[13][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n51485), .force_10(\L1_0/n3332 ), 
        .force_11(1'b0), .Q(n38464), .QN(n5154) );
  \**FFGEN**  \L1_0/abs_reg[13][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n51484), .force_10(\L1_0/n3336 ), 
        .force_11(1'b0), .Q(n38468), .QN(n5155) );
  \**FFGEN**  \L1_0/abs_reg[13][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3339 ), .force_10(n51483), 
        .force_11(1'b0), .Q(n38472), .QN(n5156) );
  \**FFGEN**  \L1_0/abs_reg[13][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n51482), .force_10(\L1_0/n3344 ), 
        .force_11(1'b0), .Q(n38476), .QN(n5157) );
  \**FFGEN**  \L1_0/abs_reg[13][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3347 ), .force_10(n51481), 
        .force_11(1'b0), .Q(n38480), .QN(n5158) );
  \**FFGEN**  \L1_0/abs_reg[13][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n51480), .force_10(\L1_0/n3352 ), 
        .force_11(1'b0), .Q(n38484), .QN(n5159) );
  \**FFGEN**  \L1_0/abs_reg[13][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3355 ), .force_10(n51479), 
        .force_11(1'b0), .Q(n38488), .QN(n5160) );
  \**FFGEN**  \L1_0/abs_reg[13][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n51478), .force_10(\L1_0/n3360 ), 
        .force_11(1'b0), .Q(n38492), .QN(n5161) );
  \**FFGEN**  \L1_0/abs_reg[13][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3363 ), .force_10(n51477), 
        .force_11(1'b0), .Q(n38496), .QN(n5162) );
  \**FFGEN**  \L1_0/abs_reg[13][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3367 ), .force_10(n51476), 
        .force_11(1'b0), .Q(n38500), .QN(n5163) );
  \**FFGEN**  \L1_0/abs_reg[13][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n51475), .force_10(\L1_0/n3372 ), 
        .force_11(1'b0), .Q(n38504), .QN(n5164) );
  \**FFGEN**  \L1_0/abs_reg[13][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n51474), .force_10(\L1_0/n3376 ), 
        .force_11(1'b0), .Q(n38508), .QN(n5165) );
  \**FFGEN**  \L1_0/abs_reg[13][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n51473), .force_10(\L1_0/n3380 ), 
        .force_11(1'b0), .Q(n38512), .QN(n5166) );
  \**FFGEN**  \L1_0/abs_reg[13][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n51472), .force_10(\L1_0/n3384 ), 
        .force_11(1'b0), .Q(n38516), .QN(n5167) );
  \**FFGEN**  \L1_0/abs_reg[13][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n51471), .force_10(\L1_0/n3388 ), 
        .force_11(1'b0), .Q(n38519), .QN(n5168) );
  \**FFGEN**  \L1_0/abs_reg[13][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n51470), .force_10(\L1_0/n3392 ), 
        .force_11(1'b0), .Q(n38188), .QN(n5169) );
  \**FFGEN**  \L1_0/abs_reg[13][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3395 ), .force_10(\L1_0/n3396 ), 
        .force_11(1'b0), .Q(n38524), .QN(n5731) );
  \**FFGEN**  \L1_0/abs_reg[12][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n5128), .force_10(\L1_0/n3400 ), .force_11(
        1'b0), .QN(n5170) );
  \**FFGEN**  \L1_0/abs_reg[12][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n51463), .force_10(\L1_0/n3404 ), 
        .force_11(1'b0), .Q(n38437), .QN(n5171) );
  \**FFGEN**  \L1_0/abs_reg[12][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n51461), .force_10(\L1_0/n3408 ), 
        .force_11(1'b0), .Q(n38432), .QN(n5172) );
  \**FFGEN**  \L1_0/abs_reg[12][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n51462), .force_10(\L1_0/n3412 ), 
        .force_11(1'b0), .Q(n38425), .QN(n5173) );
  \**FFGEN**  \L1_0/abs_reg[12][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n51457), .force_10(\L1_0/n3416 ), 
        .force_11(1'b0), .Q(n38417), .QN(n5174) );
  \**FFGEN**  \L1_0/abs_reg[12][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n5130), .force_10(n51469), .force_11(1'b0), 
        .Q(n38408), .QN(n5175) );
  \**FFGEN**  \L1_0/abs_reg[12][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n51459), .force_10(\L1_0/n3424 ), 
        .force_11(1'b0), .Q(n38400), .QN(n5176) );
  \**FFGEN**  \L1_0/abs_reg[12][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n5127), .force_10(n51468), .force_11(1'b0), 
        .Q(n38391), .QN(n5177) );
  \**FFGEN**  \L1_0/abs_reg[12][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n51464), .force_10(\L1_0/n3432 ), 
        .force_11(1'b0), .Q(n38382), .QN(n5178) );
  \**FFGEN**  \L1_0/abs_reg[12][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n5129), .force_10(n51467), .force_11(1'b0), 
        .Q(n38373), .QN(n5179) );
  \**FFGEN**  \L1_0/abs_reg[12][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n51455), .force_10(\L1_0/n3440 ), 
        .force_11(1'b0), .Q(n38364), .QN(n5180) );
  \**FFGEN**  \L1_0/abs_reg[12][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n5131), .force_10(n51466), .force_11(1'b0), 
        .Q(n38355), .QN(n5181) );
  \**FFGEN**  \L1_0/abs_reg[12][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n5126), .force_10(n51465), .force_11(1'b0), 
        .Q(n38346), .QN(n5182) );
  \**FFGEN**  \L1_0/abs_reg[12][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n51453), .force_10(\L1_0/n3452 ), 
        .force_11(1'b0), .Q(n38337), .QN(n5183) );
  \**FFGEN**  \L1_0/abs_reg[12][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n51456), .force_10(\L1_0/n3456 ), 
        .force_11(1'b0), .Q(n38328), .QN(n5184) );
  \**FFGEN**  \L1_0/abs_reg[12][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n51454), .force_10(\L1_0/n3460 ), 
        .force_11(1'b0), .Q(n38319), .QN(n5185) );
  \**FFGEN**  \L1_0/abs_reg[12][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n51452), .force_10(\L1_0/n3464 ), 
        .force_11(1'b0), .Q(n38310), .QN(n5186) );
  \**FFGEN**  \L1_0/abs_reg[12][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n51460), .force_10(\L1_0/n3468 ), 
        .force_11(1'b0), .Q(n38301), .QN(n5187) );
  \**FFGEN**  \L1_0/abs_reg[12][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n51458), .force_10(\L1_0/n3472 ), 
        .force_11(1'b0), .Q(n38185), .QN(n5188) );
  \**FFGEN**  \L1_0/abs_reg[12][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n5125), .force_10(\L1_0/n3476 ), .force_11(
        1'b0), .Q(n38127), .QN(n5730) );
  \**FFGEN**  \L1_0/abs_reg[11][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3479 ), .force_10(\L1_0/n3480 ), 
        .force_11(1'b0), .QN(n5189) );
  \**FFGEN**  \L1_0/abs_reg[11][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3483 ), .force_10(\L1_0/n3484 ), 
        .force_11(1'b0), .Q(n38433), .QN(n5190) );
  \**FFGEN**  \L1_0/abs_reg[11][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3487 ), .force_10(\L1_0/n3488 ), 
        .force_11(1'b0), .Q(n38426), .QN(n5191) );
  \**FFGEN**  \L1_0/abs_reg[11][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3491 ), .force_10(\L1_0/n3492 ), 
        .force_11(1'b0), .Q(n38418), .QN(n5192) );
  \**FFGEN**  \L1_0/abs_reg[11][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3495 ), .force_10(\L1_0/n3496 ), 
        .force_11(1'b0), .Q(n38409), .QN(n5193) );
  \**FFGEN**  \L1_0/abs_reg[11][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3499 ), .force_10(\L1_0/n3500 ), 
        .force_11(1'b0), .Q(n38401), .QN(n5194) );
  \**FFGEN**  \L1_0/abs_reg[11][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3503 ), .force_10(\L1_0/n3504 ), 
        .force_11(1'b0), .Q(n38392), .QN(n5195) );
  \**FFGEN**  \L1_0/abs_reg[11][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3507 ), .force_10(\L1_0/n3508 ), 
        .force_11(1'b0), .Q(n38383), .QN(n5196) );
  \**FFGEN**  \L1_0/abs_reg[11][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3511 ), .force_10(\L1_0/n3512 ), 
        .force_11(1'b0), .Q(n38374), .QN(n5197) );
  \**FFGEN**  \L1_0/abs_reg[11][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3515 ), .force_10(\L1_0/n3516 ), 
        .force_11(1'b0), .Q(n38365), .QN(n5198) );
  \**FFGEN**  \L1_0/abs_reg[11][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3519 ), .force_10(\L1_0/n3520 ), 
        .force_11(1'b0), .Q(n38356), .QN(n5199) );
  \**FFGEN**  \L1_0/abs_reg[11][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3523 ), .force_10(\L1_0/n3524 ), 
        .force_11(1'b0), .Q(n38347), .QN(n5200) );
  \**FFGEN**  \L1_0/abs_reg[11][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3527 ), .force_10(\L1_0/n3528 ), 
        .force_11(1'b0), .Q(n38338), .QN(n5201) );
  \**FFGEN**  \L1_0/abs_reg[11][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3531 ), .force_10(\L1_0/n3532 ), 
        .force_11(1'b0), .Q(n38329), .QN(n5202) );
  \**FFGEN**  \L1_0/abs_reg[11][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3535 ), .force_10(\L1_0/n3536 ), 
        .force_11(1'b0), .Q(n38320), .QN(n5203) );
  \**FFGEN**  \L1_0/abs_reg[11][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3539 ), .force_10(\L1_0/n3540 ), 
        .force_11(1'b0), .Q(n38311), .QN(n5204) );
  \**FFGEN**  \L1_0/abs_reg[11][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3543 ), .force_10(\L1_0/n3544 ), 
        .force_11(1'b0), .Q(n38302), .QN(n5205) );
  \**FFGEN**  \L1_0/abs_reg[11][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3547 ), .force_10(\L1_0/n3548 ), 
        .force_11(1'b0), .Q(n38290), .QN(n5206) );
  \**FFGEN**  \L1_0/abs_reg[11][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3551 ), .force_10(\L1_0/n3552 ), 
        .force_11(1'b0), .Q(n38181), .QN(n5207) );
  \**FFGEN**  \L1_0/abs_reg[11][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3555 ), .force_10(\L1_0/n3556 ), 
        .force_11(1'b0), .Q(n38523), .QN(n5729) );
  \**FFGEN**  \L1_0/abs_reg[10][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3559 ), .force_10(\L1_0/n3560 ), 
        .force_11(1'b0), .QN(n5208) );
  \**FFGEN**  \L1_0/abs_reg[10][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3563 ), .force_10(\L1_0/n3564 ), 
        .force_11(1'b0), .Q(n38427), .QN(n5209) );
  \**FFGEN**  \L1_0/abs_reg[10][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3567 ), .force_10(\L1_0/n3568 ), 
        .force_11(1'b0), .Q(n38419), .QN(n5210) );
  \**FFGEN**  \L1_0/abs_reg[10][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3571 ), .force_10(\L1_0/n3572 ), 
        .force_11(1'b0), .Q(n38410), .QN(n5211) );
  \**FFGEN**  \L1_0/abs_reg[10][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3575 ), .force_10(\L1_0/n3576 ), 
        .force_11(1'b0), .Q(n38402), .QN(n5212) );
  \**FFGEN**  \L1_0/abs_reg[10][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3579 ), .force_10(\L1_0/n3580 ), 
        .force_11(1'b0), .Q(n38393), .QN(n5213) );
  \**FFGEN**  \L1_0/abs_reg[10][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3583 ), .force_10(\L1_0/n3584 ), 
        .force_11(1'b0), .Q(n38384), .QN(n5214) );
  \**FFGEN**  \L1_0/abs_reg[10][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3587 ), .force_10(\L1_0/n3588 ), 
        .force_11(1'b0), .Q(n38375), .QN(n5215) );
  \**FFGEN**  \L1_0/abs_reg[10][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3591 ), .force_10(\L1_0/n3592 ), 
        .force_11(1'b0), .Q(n38366), .QN(n5216) );
  \**FFGEN**  \L1_0/abs_reg[10][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3595 ), .force_10(\L1_0/n3596 ), 
        .force_11(1'b0), .Q(n38357), .QN(n5217) );
  \**FFGEN**  \L1_0/abs_reg[10][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3599 ), .force_10(\L1_0/n3600 ), 
        .force_11(1'b0), .Q(n38348), .QN(n5218) );
  \**FFGEN**  \L1_0/abs_reg[10][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3603 ), .force_10(\L1_0/n3604 ), 
        .force_11(1'b0), .Q(n38339), .QN(n5219) );
  \**FFGEN**  \L1_0/abs_reg[10][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3607 ), .force_10(\L1_0/n3608 ), 
        .force_11(1'b0), .Q(n38330), .QN(n5220) );
  \**FFGEN**  \L1_0/abs_reg[10][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3611 ), .force_10(\L1_0/n3612 ), 
        .force_11(1'b0), .Q(n38321), .QN(n5221) );
  \**FFGEN**  \L1_0/abs_reg[10][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3615 ), .force_10(\L1_0/n3616 ), 
        .force_11(1'b0), .Q(n38312), .QN(n5222) );
  \**FFGEN**  \L1_0/abs_reg[10][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3619 ), .force_10(\L1_0/n3620 ), 
        .force_11(1'b0), .Q(n38303), .QN(n5223) );
  \**FFGEN**  \L1_0/abs_reg[10][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3623 ), .force_10(\L1_0/n3624 ), 
        .force_11(1'b0), .Q(n38294), .QN(n5224) );
  \**FFGEN**  \L1_0/abs_reg[10][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3627 ), .force_10(\L1_0/n3628 ), 
        .force_11(1'b0), .Q(n38287), .QN(n5225) );
  \**FFGEN**  \L1_0/abs_reg[10][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3631 ), .force_10(\L1_0/n3632 ), 
        .force_11(1'b0), .Q(n38179), .QN(n5226) );
  \**FFGEN**  \L1_0/abs_reg[10][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3635 ), .force_10(\L1_0/n3636 ), 
        .force_11(1'b0), .Q(n38191), .QN(n5728) );
  \**FFGEN**  \L1_0/abs_reg[9][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3639 ), .force_10(\L1_0/n3640 ), 
        .force_11(1'b0), .QN(n5227) );
  \**FFGEN**  \L1_0/abs_reg[9][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3643 ), .force_10(\L1_0/n3644 ), 
        .force_11(1'b0), .Q(n38420), .QN(n5228) );
  \**FFGEN**  \L1_0/abs_reg[9][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3647 ), .force_10(\L1_0/n3648 ), 
        .force_11(1'b0), .Q(n38411), .QN(n5229) );
  \**FFGEN**  \L1_0/abs_reg[9][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3651 ), .force_10(\L1_0/n3652 ), 
        .force_11(1'b0), .Q(n38403), .QN(n5230) );
  \**FFGEN**  \L1_0/abs_reg[9][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3655 ), .force_10(\L1_0/n3656 ), 
        .force_11(1'b0), .Q(n38394), .QN(n5231) );
  \**FFGEN**  \L1_0/abs_reg[9][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3659 ), .force_10(\L1_0/n3660 ), 
        .force_11(1'b0), .Q(n38385), .QN(n5232) );
  \**FFGEN**  \L1_0/abs_reg[9][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3663 ), .force_10(\L1_0/n3664 ), 
        .force_11(1'b0), .Q(n38376), .QN(n5233) );
  \**FFGEN**  \L1_0/abs_reg[9][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3667 ), .force_10(\L1_0/n3668 ), 
        .force_11(1'b0), .Q(n38367), .QN(n5234) );
  \**FFGEN**  \L1_0/abs_reg[9][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3671 ), .force_10(\L1_0/n3672 ), 
        .force_11(1'b0), .Q(n38358), .QN(n5235) );
  \**FFGEN**  \L1_0/abs_reg[9][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3675 ), .force_10(\L1_0/n3676 ), 
        .force_11(1'b0), .Q(n38349), .QN(n5236) );
  \**FFGEN**  \L1_0/abs_reg[9][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3679 ), .force_10(\L1_0/n3680 ), 
        .force_11(1'b0), .Q(n38340), .QN(n5237) );
  \**FFGEN**  \L1_0/abs_reg[9][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3683 ), .force_10(\L1_0/n3684 ), 
        .force_11(1'b0), .Q(n38331), .QN(n5238) );
  \**FFGEN**  \L1_0/abs_reg[9][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3687 ), .force_10(\L1_0/n3688 ), 
        .force_11(1'b0), .Q(n38322), .QN(n5239) );
  \**FFGEN**  \L1_0/abs_reg[9][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3691 ), .force_10(\L1_0/n3692 ), 
        .force_11(1'b0), .Q(n38313), .QN(n5240) );
  \**FFGEN**  \L1_0/abs_reg[9][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3695 ), .force_10(\L1_0/n3696 ), 
        .force_11(1'b0), .Q(n38304), .QN(n5241) );
  \**FFGEN**  \L1_0/abs_reg[9][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3699 ), .force_10(\L1_0/n3700 ), 
        .force_11(1'b0), .Q(n38295), .QN(n5242) );
  \**FFGEN**  \L1_0/abs_reg[9][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3703 ), .force_10(\L1_0/n3704 ), 
        .force_11(1'b0), .Q(n38288), .QN(n5243) );
  \**FFGEN**  \L1_0/abs_reg[9][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3707 ), .force_10(\L1_0/n3708 ), 
        .force_11(1'b0), .Q(n38285), .QN(n5244) );
  \**FFGEN**  \L1_0/abs_reg[9][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3711 ), .force_10(\L1_0/n3712 ), 
        .force_11(1'b0), .Q(n38178), .QN(n5245) );
  \**FFGEN**  \L1_0/abs_reg[9][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3715 ), .force_10(\L1_0/n3716 ), 
        .force_11(1'b0), .Q(n38520), .QN(n5727) );
  \**FFGEN**  \L1_0/abs_reg[8][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3719 ), .force_10(\L1_0/n3720 ), 
        .force_11(1'b0), .QN(n5246) );
  \**FFGEN**  \L1_0/abs_reg[8][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3723 ), .force_10(\L1_0/n3724 ), 
        .force_11(1'b0), .Q(n38412), .QN(n5247) );
  \**FFGEN**  \L1_0/abs_reg[8][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3727 ), .force_10(\L1_0/n3728 ), 
        .force_11(1'b0), .Q(n38404), .QN(n5248) );
  \**FFGEN**  \L1_0/abs_reg[8][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3731 ), .force_10(\L1_0/n3732 ), 
        .force_11(1'b0), .Q(n38395), .QN(n5249) );
  \**FFGEN**  \L1_0/abs_reg[8][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3735 ), .force_10(\L1_0/n3736 ), 
        .force_11(1'b0), .Q(n38386), .QN(n5250) );
  \**FFGEN**  \L1_0/abs_reg[8][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3739 ), .force_10(\L1_0/n3740 ), 
        .force_11(1'b0), .Q(n38377), .QN(n5251) );
  \**FFGEN**  \L1_0/abs_reg[8][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3743 ), .force_10(\L1_0/n3744 ), 
        .force_11(1'b0), .Q(n38368), .QN(n5252) );
  \**FFGEN**  \L1_0/abs_reg[8][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3747 ), .force_10(\L1_0/n3748 ), 
        .force_11(1'b0), .Q(n38359), .QN(n5253) );
  \**FFGEN**  \L1_0/abs_reg[8][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3751 ), .force_10(\L1_0/n3752 ), 
        .force_11(1'b0), .Q(n38350), .QN(n5254) );
  \**FFGEN**  \L1_0/abs_reg[8][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3755 ), .force_10(\L1_0/n3756 ), 
        .force_11(1'b0), .Q(n38341), .QN(n5255) );
  \**FFGEN**  \L1_0/abs_reg[8][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3759 ), .force_10(\L1_0/n3760 ), 
        .force_11(1'b0), .Q(n38332), .QN(n5256) );
  \**FFGEN**  \L1_0/abs_reg[8][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3763 ), .force_10(\L1_0/n3764 ), 
        .force_11(1'b0), .Q(n38323), .QN(n5257) );
  \**FFGEN**  \L1_0/abs_reg[8][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3767 ), .force_10(\L1_0/n3768 ), 
        .force_11(1'b0), .Q(n38314), .QN(n5258) );
  \**FFGEN**  \L1_0/abs_reg[8][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3771 ), .force_10(\L1_0/n3772 ), 
        .force_11(1'b0), .Q(n38305), .QN(n5259) );
  \**FFGEN**  \L1_0/abs_reg[8][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3775 ), .force_10(\L1_0/n3776 ), 
        .force_11(1'b0), .Q(n38296), .QN(n5260) );
  \**FFGEN**  \L1_0/abs_reg[8][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3779 ), .force_10(\L1_0/n3780 ), 
        .force_11(1'b0), .Q(n38292), .QN(n5261) );
  \**FFGEN**  \L1_0/abs_reg[8][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3783 ), .force_10(\L1_0/n3784 ), 
        .force_11(1'b0), .Q(n38291), .QN(n5262) );
  \**FFGEN**  \L1_0/abs_reg[8][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3787 ), .force_10(\L1_0/n3788 ), 
        .force_11(1'b0), .Q(n38283), .QN(n5263) );
  \**FFGEN**  \L1_0/abs_reg[8][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3791 ), .force_10(\L1_0/n3792 ), 
        .force_11(1'b0), .Q(n38177), .QN(n5264) );
  \**FFGEN**  \L1_0/abs_reg[8][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3795 ), .force_10(\L1_0/n3796 ), 
        .force_11(1'b0), .Q(n38133), .QN(n5726) );
  \**FFGEN**  \L1_0/abs_reg[7][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3799 ), .force_10(\L1_0/n3800 ), 
        .force_11(1'b0), .QN(n5265) );
  \**FFGEN**  \L1_0/abs_reg[7][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3803 ), .force_10(\L1_0/n3804 ), 
        .force_11(1'b0), .Q(n38239), .QN(n5266) );
  \**FFGEN**  \L1_0/abs_reg[7][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3807 ), .force_10(\L1_0/n3808 ), 
        .force_11(1'b0), .QN(n5267) );
  \**FFGEN**  \L1_0/abs_reg[7][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3811 ), .force_10(\L1_0/n3812 ), 
        .force_11(1'b0), .QN(n5268) );
  \**FFGEN**  \L1_0/abs_reg[7][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3815 ), .force_10(\L1_0/n3816 ), 
        .force_11(1'b0), .QN(n5269) );
  \**FFGEN**  \L1_0/abs_reg[7][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3819 ), .force_10(\L1_0/n3820 ), 
        .force_11(1'b0), .QN(n5270) );
  \**FFGEN**  \L1_0/abs_reg[7][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3823 ), .force_10(\L1_0/n3824 ), 
        .force_11(1'b0), .QN(n5271) );
  \**FFGEN**  \L1_0/abs_reg[7][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3827 ), .force_10(\L1_0/n3828 ), 
        .force_11(1'b0), .QN(n5272) );
  \**FFGEN**  \L1_0/abs_reg[7][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3831 ), .force_10(\L1_0/n3832 ), 
        .force_11(1'b0), .QN(n5273) );
  \**FFGEN**  \L1_0/abs_reg[7][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3835 ), .force_10(\L1_0/n3836 ), 
        .force_11(1'b0), .QN(n5274) );
  \**FFGEN**  \L1_0/abs_reg[7][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3839 ), .force_10(\L1_0/n3840 ), 
        .force_11(1'b0), .QN(n5275) );
  \**FFGEN**  \L1_0/abs_reg[7][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3843 ), .force_10(\L1_0/n3844 ), 
        .force_11(1'b0), .QN(n5276) );
  \**FFGEN**  \L1_0/abs_reg[7][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3847 ), .force_10(\L1_0/n3848 ), 
        .force_11(1'b0), .QN(n5277) );
  \**FFGEN**  \L1_0/abs_reg[7][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3851 ), .force_10(\L1_0/n3852 ), 
        .force_11(1'b0), .QN(n5278) );
  \**FFGEN**  \L1_0/abs_reg[7][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3855 ), .force_10(\L1_0/n3856 ), 
        .force_11(1'b0), .QN(n5279) );
  \**FFGEN**  \L1_0/abs_reg[7][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3859 ), .force_10(\L1_0/n3860 ), 
        .force_11(1'b0), .QN(n5280) );
  \**FFGEN**  \L1_0/abs_reg[7][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3863 ), .force_10(\L1_0/n3864 ), 
        .force_11(1'b0), .Q(n38128), .QN(n5281) );
  \**FFGEN**  \L1_0/abs_reg[7][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3867 ), .force_10(\L1_0/n3868 ), 
        .force_11(1'b0), .QN(n5282) );
  \**FFGEN**  \L1_0/abs_reg[7][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3871 ), .force_10(\L1_0/n3872 ), 
        .force_11(1'b0), .Q(n38168), .QN(n5283) );
  \**FFGEN**  \L1_0/abs_reg[7][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3875 ), .force_10(\L1_0/n3876 ), 
        .force_11(1'b0), .Q(n38147), .QN(n5725) );
  \**FFGEN**  \L1_0/abs_reg[6][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3879 ), .force_10(\L1_0/n3880 ), 
        .force_11(1'b0), .QN(n5284) );
  \**FFGEN**  \L1_0/abs_reg[6][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3883 ), .force_10(\L1_0/n3884 ), 
        .force_11(1'b0), .Q(n38396), .QN(n5285) );
  \**FFGEN**  \L1_0/abs_reg[6][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3887 ), .force_10(\L1_0/n3888 ), 
        .force_11(1'b0), .Q(n38387), .QN(n5286) );
  \**FFGEN**  \L1_0/abs_reg[6][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3891 ), .force_10(\L1_0/n3892 ), 
        .force_11(1'b0), .Q(n38378), .QN(n5287) );
  \**FFGEN**  \L1_0/abs_reg[6][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3895 ), .force_10(\L1_0/n3896 ), 
        .force_11(1'b0), .Q(n38369), .QN(n5288) );
  \**FFGEN**  \L1_0/abs_reg[6][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3899 ), .force_10(\L1_0/n3900 ), 
        .force_11(1'b0), .Q(n38360), .QN(n5289) );
  \**FFGEN**  \L1_0/abs_reg[6][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3903 ), .force_10(\L1_0/n3904 ), 
        .force_11(1'b0), .Q(n38351), .QN(n5290) );
  \**FFGEN**  \L1_0/abs_reg[6][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3907 ), .force_10(\L1_0/n3908 ), 
        .force_11(1'b0), .Q(n38342), .QN(n5291) );
  \**FFGEN**  \L1_0/abs_reg[6][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3911 ), .force_10(\L1_0/n3912 ), 
        .force_11(1'b0), .Q(n38333), .QN(n5292) );
  \**FFGEN**  \L1_0/abs_reg[6][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3915 ), .force_10(\L1_0/n3916 ), 
        .force_11(1'b0), .Q(n38324), .QN(n5293) );
  \**FFGEN**  \L1_0/abs_reg[6][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3919 ), .force_10(\L1_0/n3920 ), 
        .force_11(1'b0), .Q(n38315), .QN(n5294) );
  \**FFGEN**  \L1_0/abs_reg[6][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3923 ), .force_10(\L1_0/n3924 ), 
        .force_11(1'b0), .Q(n38306), .QN(n5295) );
  \**FFGEN**  \L1_0/abs_reg[6][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3927 ), .force_10(\L1_0/n3928 ), 
        .force_11(1'b0), .Q(n38297), .QN(n5296) );
  \**FFGEN**  \L1_0/abs_reg[6][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3931 ), .force_10(\L1_0/n3932 ), 
        .force_11(1'b0), .Q(n38293), .QN(n5297) );
  \**FFGEN**  \L1_0/abs_reg[6][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3935 ), .force_10(\L1_0/n3936 ), 
        .force_11(1'b0), .Q(n38286), .QN(n5298) );
  \**FFGEN**  \L1_0/abs_reg[6][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3939 ), .force_10(\L1_0/n3940 ), 
        .force_11(1'b0), .Q(n38284), .QN(n5299) );
  \**FFGEN**  \L1_0/abs_reg[6][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3943 ), .force_10(\L1_0/n3944 ), 
        .force_11(1'b0), .Q(n38282), .QN(n5300) );
  \**FFGEN**  \L1_0/abs_reg[6][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3947 ), .force_10(\L1_0/n3948 ), 
        .force_11(1'b0), .Q(n38281), .QN(n5301) );
  \**FFGEN**  \L1_0/abs_reg[6][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3951 ), .force_10(\L1_0/n3952 ), 
        .force_11(1'b0), .Q(n38176), .QN(n5302) );
  \**FFGEN**  \L1_0/abs_reg[6][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3955 ), .force_10(\L1_0/n3956 ), 
        .force_11(1'b0), .Q(n38193), .QN(n5724) );
  \**FFGEN**  \L1_0/abs_reg[5][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3959 ), .force_10(\L1_0/n3960 ), 
        .force_11(1'b0), .QN(n5303) );
  \**FFGEN**  \L1_0/abs_reg[5][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3963 ), .force_10(\L1_0/n3964 ), 
        .force_11(1'b0), .Q(n38453), .QN(n5304) );
  \**FFGEN**  \L1_0/abs_reg[5][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3967 ), .force_10(\L1_0/n3968 ), 
        .force_11(1'b0), .Q(n38457), .QN(n5305) );
  \**FFGEN**  \L1_0/abs_reg[5][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3971 ), .force_10(\L1_0/n3972 ), 
        .force_11(1'b0), .Q(n38461), .QN(n5306) );
  \**FFGEN**  \L1_0/abs_reg[5][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3975 ), .force_10(\L1_0/n3976 ), 
        .force_11(1'b0), .Q(n38465), .QN(n5307) );
  \**FFGEN**  \L1_0/abs_reg[5][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3979 ), .force_10(\L1_0/n3980 ), 
        .force_11(1'b0), .Q(n38469), .QN(n5308) );
  \**FFGEN**  \L1_0/abs_reg[5][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3983 ), .force_10(\L1_0/n3984 ), 
        .force_11(1'b0), .Q(n38473), .QN(n5309) );
  \**FFGEN**  \L1_0/abs_reg[5][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3987 ), .force_10(\L1_0/n3988 ), 
        .force_11(1'b0), .Q(n38477), .QN(n5310) );
  \**FFGEN**  \L1_0/abs_reg[5][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3991 ), .force_10(\L1_0/n3992 ), 
        .force_11(1'b0), .Q(n38481), .QN(n5311) );
  \**FFGEN**  \L1_0/abs_reg[5][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3995 ), .force_10(\L1_0/n3996 ), 
        .force_11(1'b0), .Q(n38485), .QN(n5312) );
  \**FFGEN**  \L1_0/abs_reg[5][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3999 ), .force_10(\L1_0/n4000 ), 
        .force_11(1'b0), .Q(n38489), .QN(n5313) );
  \**FFGEN**  \L1_0/abs_reg[5][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4003 ), .force_10(\L1_0/n4004 ), 
        .force_11(1'b0), .Q(n38493), .QN(n5314) );
  \**FFGEN**  \L1_0/abs_reg[5][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4007 ), .force_10(\L1_0/n4008 ), 
        .force_11(1'b0), .Q(n38497), .QN(n5315) );
  \**FFGEN**  \L1_0/abs_reg[5][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4011 ), .force_10(\L1_0/n4012 ), 
        .force_11(1'b0), .Q(n38501), .QN(n5316) );
  \**FFGEN**  \L1_0/abs_reg[5][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4015 ), .force_10(\L1_0/n4016 ), 
        .force_11(1'b0), .Q(n38505), .QN(n5317) );
  \**FFGEN**  \L1_0/abs_reg[5][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4019 ), .force_10(\L1_0/n4020 ), 
        .force_11(1'b0), .Q(n38509), .QN(n5318) );
  \**FFGEN**  \L1_0/abs_reg[5][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4023 ), .force_10(\L1_0/n4024 ), 
        .force_11(1'b0), .Q(n38513), .QN(n5319) );
  \**FFGEN**  \L1_0/abs_reg[5][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4027 ), .force_10(\L1_0/n4028 ), 
        .force_11(1'b0), .Q(n38517), .QN(n5320) );
  \**FFGEN**  \L1_0/abs_reg[5][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4031 ), .force_10(\L1_0/n4032 ), 
        .force_11(1'b0), .Q(n38186), .QN(n5321) );
  \**FFGEN**  \L1_0/abs_reg[5][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4035 ), .force_10(\L1_0/n4036 ), 
        .force_11(1'b0), .Q(n38522), .QN(n5723) );
  \**FFGEN**  \L1_0/abs_reg[4][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4039 ), .force_10(\L1_0/n4040 ), 
        .force_11(1'b0), .QN(n5322) );
  \**FFGEN**  \L1_0/abs_reg[4][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4043 ), .force_10(\L1_0/n4044 ), 
        .force_11(1'b0), .Q(n38435), .QN(n5323) );
  \**FFGEN**  \L1_0/abs_reg[4][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4047 ), .force_10(\L1_0/n4048 ), 
        .force_11(1'b0), .Q(n38429), .QN(n5324) );
  \**FFGEN**  \L1_0/abs_reg[4][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4051 ), .force_10(\L1_0/n4052 ), 
        .force_11(1'b0), .Q(n38422), .QN(n5325) );
  \**FFGEN**  \L1_0/abs_reg[4][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4055 ), .force_10(\L1_0/n4056 ), 
        .force_11(1'b0), .Q(n38414), .QN(n5326) );
  \**FFGEN**  \L1_0/abs_reg[4][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4059 ), .force_10(\L1_0/n4060 ), 
        .force_11(1'b0), .Q(n38405), .QN(n5327) );
  \**FFGEN**  \L1_0/abs_reg[4][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4063 ), .force_10(\L1_0/n4064 ), 
        .force_11(1'b0), .Q(n38397), .QN(n5328) );
  \**FFGEN**  \L1_0/abs_reg[4][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4067 ), .force_10(\L1_0/n4068 ), 
        .force_11(1'b0), .Q(n38388), .QN(n5329) );
  \**FFGEN**  \L1_0/abs_reg[4][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4071 ), .force_10(\L1_0/n4072 ), 
        .force_11(1'b0), .Q(n38379), .QN(n5330) );
  \**FFGEN**  \L1_0/abs_reg[4][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4075 ), .force_10(\L1_0/n4076 ), 
        .force_11(1'b0), .Q(n38370), .QN(n5331) );
  \**FFGEN**  \L1_0/abs_reg[4][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4079 ), .force_10(\L1_0/n4080 ), 
        .force_11(1'b0), .Q(n38361), .QN(n5332) );
  \**FFGEN**  \L1_0/abs_reg[4][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4083 ), .force_10(\L1_0/n4084 ), 
        .force_11(1'b0), .Q(n38352), .QN(n5333) );
  \**FFGEN**  \L1_0/abs_reg[4][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4087 ), .force_10(\L1_0/n4088 ), 
        .force_11(1'b0), .Q(n38343), .QN(n5334) );
  \**FFGEN**  \L1_0/abs_reg[4][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4091 ), .force_10(\L1_0/n4092 ), 
        .force_11(1'b0), .Q(n38334), .QN(n5335) );
  \**FFGEN**  \L1_0/abs_reg[4][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4095 ), .force_10(\L1_0/n4096 ), 
        .force_11(1'b0), .Q(n38325), .QN(n5336) );
  \**FFGEN**  \L1_0/abs_reg[4][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4099 ), .force_10(\L1_0/n4100 ), 
        .force_11(1'b0), .Q(n38316), .QN(n5337) );
  \**FFGEN**  \L1_0/abs_reg[4][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4103 ), .force_10(\L1_0/n4104 ), 
        .force_11(1'b0), .Q(n38307), .QN(n5338) );
  \**FFGEN**  \L1_0/abs_reg[4][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4107 ), .force_10(\L1_0/n4108 ), 
        .force_11(1'b0), .Q(n38298), .QN(n5339) );
  \**FFGEN**  \L1_0/abs_reg[4][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4111 ), .force_10(\L1_0/n4112 ), 
        .force_11(1'b0), .Q(n38183), .QN(n5340) );
  \**FFGEN**  \L1_0/abs_reg[4][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4115 ), .force_10(\L1_0/n4116 ), 
        .force_11(1'b0), .Q(n38192), .QN(n5722) );
  \**FFGEN**  \L1_0/abs_reg[3][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4119 ), .force_10(\L1_0/n4120 ), 
        .force_11(1'b0), .QN(n5341) );
  \**FFGEN**  \L1_0/abs_reg[3][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4123 ), .force_10(\L1_0/n4124 ), 
        .force_11(1'b0), .Q(n38430), .QN(n5342) );
  \**FFGEN**  \L1_0/abs_reg[3][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4127 ), .force_10(\L1_0/n4128 ), 
        .force_11(1'b0), .Q(n38423), .QN(n5343) );
  \**FFGEN**  \L1_0/abs_reg[3][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4131 ), .force_10(\L1_0/n4132 ), 
        .force_11(1'b0), .Q(n38415), .QN(n5344) );
  \**FFGEN**  \L1_0/abs_reg[3][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4135 ), .force_10(\L1_0/n4136 ), 
        .force_11(1'b0), .Q(n38406), .QN(n5345) );
  \**FFGEN**  \L1_0/abs_reg[3][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4139 ), .force_10(\L1_0/n4140 ), 
        .force_11(1'b0), .Q(n38398), .QN(n5346) );
  \**FFGEN**  \L1_0/abs_reg[3][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4143 ), .force_10(\L1_0/n4144 ), 
        .force_11(1'b0), .Q(n38389), .QN(n5347) );
  \**FFGEN**  \L1_0/abs_reg[3][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4147 ), .force_10(\L1_0/n4148 ), 
        .force_11(1'b0), .Q(n38380), .QN(n5348) );
  \**FFGEN**  \L1_0/abs_reg[3][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4151 ), .force_10(\L1_0/n4152 ), 
        .force_11(1'b0), .Q(n38371), .QN(n5349) );
  \**FFGEN**  \L1_0/abs_reg[3][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4155 ), .force_10(\L1_0/n4156 ), 
        .force_11(1'b0), .Q(n38362), .QN(n5350) );
  \**FFGEN**  \L1_0/abs_reg[3][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4159 ), .force_10(\L1_0/n4160 ), 
        .force_11(1'b0), .Q(n38353), .QN(n5351) );
  \**FFGEN**  \L1_0/abs_reg[3][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4163 ), .force_10(\L1_0/n4164 ), 
        .force_11(1'b0), .Q(n38344), .QN(n5352) );
  \**FFGEN**  \L1_0/abs_reg[3][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4167 ), .force_10(\L1_0/n4168 ), 
        .force_11(1'b0), .Q(n38335), .QN(n5353) );
  \**FFGEN**  \L1_0/abs_reg[3][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4171 ), .force_10(\L1_0/n4172 ), 
        .force_11(1'b0), .Q(n38326), .QN(n5354) );
  \**FFGEN**  \L1_0/abs_reg[3][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4175 ), .force_10(\L1_0/n4176 ), 
        .force_11(1'b0), .Q(n38317), .QN(n5355) );
  \**FFGEN**  \L1_0/abs_reg[3][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4179 ), .force_10(\L1_0/n4180 ), 
        .force_11(1'b0), .Q(n38308), .QN(n5356) );
  \**FFGEN**  \L1_0/abs_reg[3][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4183 ), .force_10(\L1_0/n4184 ), 
        .force_11(1'b0), .Q(n38299), .QN(n5357) );
  \**FFGEN**  \L1_0/abs_reg[3][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4187 ), .force_10(\L1_0/n4188 ), 
        .force_11(1'b0), .Q(n38289), .QN(n5358) );
  \**FFGEN**  \L1_0/abs_reg[3][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4191 ), .force_10(\L1_0/n4192 ), 
        .force_11(1'b0), .Q(n38180), .QN(n5359) );
  \**FFGEN**  \L1_0/abs_reg[3][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4195 ), .force_10(\L1_0/n4196 ), 
        .force_11(1'b0), .Q(n38521), .QN(n5721) );
  \**FFGEN**  \L1_0/abs_reg[2][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4199 ), .force_10(\L1_0/n4200 ), 
        .force_11(1'b0), .QN(n5360) );
  \**FFGEN**  \L1_0/abs_reg[2][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4203 ), .force_10(\L1_0/n4204 ), 
        .force_11(1'b0), .Q(n38454), .QN(n5361) );
  \**FFGEN**  \L1_0/abs_reg[2][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4207 ), .force_10(\L1_0/n4208 ), 
        .force_11(1'b0), .Q(n38458), .QN(n5362) );
  \**FFGEN**  \L1_0/abs_reg[2][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4211 ), .force_10(\L1_0/n4212 ), 
        .force_11(1'b0), .Q(n38462), .QN(n5363) );
  \**FFGEN**  \L1_0/abs_reg[2][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4215 ), .force_10(\L1_0/n4216 ), 
        .force_11(1'b0), .Q(n38466), .QN(n5364) );
  \**FFGEN**  \L1_0/abs_reg[2][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4219 ), .force_10(\L1_0/n4220 ), 
        .force_11(1'b0), .Q(n38470), .QN(n5365) );
  \**FFGEN**  \L1_0/abs_reg[2][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4223 ), .force_10(\L1_0/n4224 ), 
        .force_11(1'b0), .Q(n38474), .QN(n5366) );
  \**FFGEN**  \L1_0/abs_reg[2][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4227 ), .force_10(\L1_0/n4228 ), 
        .force_11(1'b0), .Q(n38478), .QN(n5367) );
  \**FFGEN**  \L1_0/abs_reg[2][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4231 ), .force_10(\L1_0/n4232 ), 
        .force_11(1'b0), .Q(n38482), .QN(n5368) );
  \**FFGEN**  \L1_0/abs_reg[2][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4235 ), .force_10(\L1_0/n4236 ), 
        .force_11(1'b0), .Q(n38486), .QN(n5369) );
  \**FFGEN**  \L1_0/abs_reg[2][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4239 ), .force_10(\L1_0/n4240 ), 
        .force_11(1'b0), .Q(n38490), .QN(n5370) );
  \**FFGEN**  \L1_0/abs_reg[2][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4243 ), .force_10(\L1_0/n4244 ), 
        .force_11(1'b0), .Q(n38494), .QN(n5371) );
  \**FFGEN**  \L1_0/abs_reg[2][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4247 ), .force_10(\L1_0/n4248 ), 
        .force_11(1'b0), .Q(n38498), .QN(n5372) );
  \**FFGEN**  \L1_0/abs_reg[2][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4251 ), .force_10(\L1_0/n4252 ), 
        .force_11(1'b0), .Q(n38502), .QN(n5373) );
  \**FFGEN**  \L1_0/abs_reg[2][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4255 ), .force_10(\L1_0/n4256 ), 
        .force_11(1'b0), .Q(n38506), .QN(n5374) );
  \**FFGEN**  \L1_0/abs_reg[2][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4259 ), .force_10(\L1_0/n4260 ), 
        .force_11(1'b0), .Q(n38510), .QN(n5375) );
  \**FFGEN**  \L1_0/abs_reg[2][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4263 ), .force_10(\L1_0/n4264 ), 
        .force_11(1'b0), .Q(n38514), .QN(n5376) );
  \**FFGEN**  \L1_0/abs_reg[2][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4267 ), .force_10(\L1_0/n4268 ), 
        .force_11(1'b0), .Q(n38518), .QN(n5377) );
  \**FFGEN**  \L1_0/abs_reg[2][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4271 ), .force_10(\L1_0/n4272 ), 
        .force_11(1'b0), .Q(n38187), .QN(n5378) );
  \**FFGEN**  \L1_0/abs_reg[2][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4275 ), .force_10(\L1_0/n4276 ), 
        .force_11(1'b0), .Q(n38134), .QN(n5720) );
  \**FFGEN**  \L1_0/abs_reg[1][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4279 ), .force_10(\L1_0/n4280 ), 
        .force_11(1'b0), .QN(n5379) );
  \**FFGEN**  \L1_0/abs_reg[1][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4283 ), .force_10(\L1_0/n4284 ), 
        .force_11(1'b0), .Q(n38436), .QN(n5380) );
  \**FFGEN**  \L1_0/abs_reg[1][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4287 ), .force_10(\L1_0/n4288 ), 
        .force_11(1'b0), .Q(n38431), .QN(n5381) );
  \**FFGEN**  \L1_0/abs_reg[1][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4291 ), .force_10(\L1_0/n4292 ), 
        .force_11(1'b0), .Q(n38424), .QN(n5382) );
  \**FFGEN**  \L1_0/abs_reg[1][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4295 ), .force_10(\L1_0/n4296 ), 
        .force_11(1'b0), .Q(n38416), .QN(n5383) );
  \**FFGEN**  \L1_0/abs_reg[1][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4299 ), .force_10(\L1_0/n4300 ), 
        .force_11(1'b0), .Q(n38407), .QN(n5384) );
  \**FFGEN**  \L1_0/abs_reg[1][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4303 ), .force_10(\L1_0/n4304 ), 
        .force_11(1'b0), .Q(n38399), .QN(n5385) );
  \**FFGEN**  \L1_0/abs_reg[1][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4307 ), .force_10(\L1_0/n4308 ), 
        .force_11(1'b0), .Q(n38390), .QN(n5386) );
  \**FFGEN**  \L1_0/abs_reg[1][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4311 ), .force_10(\L1_0/n4312 ), 
        .force_11(1'b0), .Q(n38381), .QN(n5387) );
  \**FFGEN**  \L1_0/abs_reg[1][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4315 ), .force_10(\L1_0/n4316 ), 
        .force_11(1'b0), .Q(n38372), .QN(n5388) );
  \**FFGEN**  \L1_0/abs_reg[1][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4319 ), .force_10(\L1_0/n4320 ), 
        .force_11(1'b0), .Q(n38363), .QN(n5389) );
  \**FFGEN**  \L1_0/abs_reg[1][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4323 ), .force_10(\L1_0/n4324 ), 
        .force_11(1'b0), .Q(n38354), .QN(n5390) );
  \**FFGEN**  \L1_0/abs_reg[1][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4327 ), .force_10(\L1_0/n4328 ), 
        .force_11(1'b0), .Q(n38345), .QN(n5391) );
  \**FFGEN**  \L1_0/abs_reg[1][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4331 ), .force_10(\L1_0/n4332 ), 
        .force_11(1'b0), .Q(n38336), .QN(n5392) );
  \**FFGEN**  \L1_0/abs_reg[1][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4335 ), .force_10(\L1_0/n4336 ), 
        .force_11(1'b0), .Q(n38327), .QN(n5393) );
  \**FFGEN**  \L1_0/abs_reg[1][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4339 ), .force_10(\L1_0/n4340 ), 
        .force_11(1'b0), .Q(n38318), .QN(n5394) );
  \**FFGEN**  \L1_0/abs_reg[1][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4343 ), .force_10(\L1_0/n4344 ), 
        .force_11(1'b0), .Q(n38309), .QN(n5395) );
  \**FFGEN**  \L1_0/abs_reg[1][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4347 ), .force_10(\L1_0/n4348 ), 
        .force_11(1'b0), .Q(n38300), .QN(n5396) );
  \**FFGEN**  \L1_0/abs_reg[1][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4351 ), .force_10(\L1_0/n4352 ), 
        .force_11(1'b0), .Q(n38184), .QN(n5397) );
  \**FFGEN**  \L1_0/abs_reg[1][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4355 ), .force_10(\L1_0/n4356 ), 
        .force_11(1'b0), .Q(n38196), .QN(n5719) );
  \**FFGEN**  \L1_0/abs_reg[0][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n5113), .force_10(n51528), .force_11(1'b0), 
        .QN(n5398) );
  \**FFGEN**  \L1_0/abs_reg[0][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n51518), .force_10(\L1_0/n4364 ), 
        .force_11(1'b0), .Q(n38190), .QN(n5399) );
  \**FFGEN**  \L1_0/abs_reg[0][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n51515), .force_10(\L1_0/n4368 ), 
        .force_11(1'b0), .Q(n42118), .QN(n5400) );
  \**FFGEN**  \L1_0/abs_reg[0][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n51526), .force_10(\L1_0/n4372 ), 
        .force_11(1'b0), .Q(n38126) );
  \**FFGEN**  \L1_0/abs_reg[0][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n51524), .force_10(\L1_0/n4376 ), 
        .force_11(1'b0), .Q(n38166), .QN(n5402) );
  \**FFGEN**  \L1_0/abs_reg[0][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n51519), .force_10(\L1_0/n4380 ), 
        .force_11(1'b0), .Q(n38124) );
  \**FFGEN**  \L1_0/abs_reg[0][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n51512), .force_10(\L1_0/n4384 ), 
        .force_11(1'b0), .Q(n38164), .QN(n5404) );
  \**FFGEN**  \L1_0/abs_reg[0][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n51516), .force_10(\L1_0/n4388 ), 
        .force_11(1'b0), .Q(n38122) );
  \**FFGEN**  \L1_0/abs_reg[0][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n51521), .force_10(\L1_0/n4392 ), 
        .force_11(1'b0), .Q(n38163), .QN(n5406) );
  \**FFGEN**  \L1_0/abs_reg[0][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n51513), .force_10(\L1_0/n4396 ), 
        .force_11(1'b0), .Q(n38121) );
  \**FFGEN**  \L1_0/abs_reg[0][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n51517), .force_10(\L1_0/n4400 ), 
        .force_11(1'b0), .Q(n38162), .QN(n5408) );
  \**FFGEN**  \L1_0/abs_reg[0][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n51523), .force_10(\L1_0/n4404 ), 
        .force_11(1'b0), .Q(n42117), .QN(n5409) );
  \**FFGEN**  \L1_0/abs_reg[0][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n5123), .force_10(n51527), .force_11(1'b0), 
        .Q(n38156), .QN(n5410) );
  \**FFGEN**  \L1_0/abs_reg[0][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n51511), .force_10(\L1_0/n4412 ), 
        .force_11(1'b0), .Q(n42116), .QN(n5411) );
  \**FFGEN**  \L1_0/abs_reg[0][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n51520), .force_10(\L1_0/n4416 ), 
        .force_11(1'b0), .Q(n38155), .QN(n5412) );
  \**FFGEN**  \L1_0/abs_reg[0][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n51522), .force_10(\L1_0/n4420 ), 
        .force_11(1'b0), .Q(n42115), .QN(n5413) );
  \**FFGEN**  \L1_0/abs_reg[0][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n51525), .force_10(\L1_0/n4424 ), 
        .force_11(1'b0), .Q(n38154), .QN(n5414) );
  \**FFGEN**  \L1_0/abs_reg[0][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n51514), .force_10(\L1_0/n4428 ), 
        .force_11(1'b0), .Q(n42114), .QN(n5415) );
  \**FFGEN**  \L1_0/abs_reg[0][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n51510), .force_10(\L1_0/n4432 ), 
        .force_11(1'b0), .Q(n38555) );
  \**FFGEN**  \L1_0/abs_reg[0][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n5114), .force_10(\L1_0/n4436 ), .force_11(
        1'b0), .Q(n38598), .QN(n5718) );
  \**FFGEN**  \L1_0/sum_reg[0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4439 ), .force_10(n5104), .force_11(
        1'b0), .Q(out_L1[0]), .QN(n38562) );
  \**FFGEN**  \L1_0/sum_reg[1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4443 ), .force_10(n5102), .force_11(
        1'b0), .Q(out_L1[1]) );
  \**FFGEN**  \L1_0/sum_reg[2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4447 ), .force_10(n5108), .force_11(
        1'b0), .Q(out_L1[2]) );
  \**FFGEN**  \L1_0/sum_reg[3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4451 ), .force_10(n5118), .force_11(
        1'b0), .Q(out_L1[3]), .QN(n38541) );
  \**FFGEN**  \L1_0/sum_reg[4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4455 ), .force_10(n5121), .force_11(
        1'b0), .Q(out_L1[4]) );
  \**FFGEN**  \L1_0/sum_reg[5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4459 ), .force_10(n5117), .force_11(
        1'b0), .Q(out_L1[5]), .QN(n38542) );
  \**FFGEN**  \L1_0/sum_reg[6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4463 ), .force_10(n5111), .force_11(
        1'b0), .Q(out_L1[6]) );
  \**FFGEN**  \L1_0/sum_reg[7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4467 ), .force_10(n5120), .force_11(
        1'b0), .Q(out_L1[7]), .QN(n38543) );
  \**FFGEN**  \L1_0/sum_reg[8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4471 ), .force_10(n5105), .force_11(
        1'b0), .Q(out_L1[8]) );
  \**FFGEN**  \L1_0/sum_reg[9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4475 ), .force_10(n5119), .force_11(
        1'b0), .Q(out_L1[9]), .QN(n38544) );
  \**FFGEN**  \L1_0/sum_reg[10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4479 ), .force_10(n5122), .force_11(
        1'b0), .Q(out_L1[10]) );
  \**FFGEN**  \L1_0/sum_reg[11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4483 ), .force_10(n5110), .force_11(
        1'b0), .Q(out_L1[11]), .QN(n38545) );
  \**FFGEN**  \L1_0/sum_reg[12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4487 ), .force_10(n5112), .force_11(
        1'b0), .Q(out_L1[12]) );
  \**FFGEN**  \L1_0/sum_reg[13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4491 ), .force_10(n5107), .force_11(
        1'b0), .Q(out_L1[13]), .QN(n38546) );
  \**FFGEN**  \L1_0/sum_reg[14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4495 ), .force_10(n5116), .force_11(
        1'b0), .Q(out_L1[14]) );
  \**FFGEN**  \L1_0/sum_reg[15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4499 ), .force_10(n5115), .force_11(
        1'b0), .Q(out_L1[15]), .QN(n38547) );
  \**FFGEN**  \L1_0/sum_reg[16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4503 ), .force_10(n5124), .force_11(
        1'b0), .Q(out_L1[16]) );
  \**FFGEN**  \L1_0/sum_reg[17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4507 ), .force_10(n5106), .force_11(
        1'b0), .Q(out_L1[17]) );
  \**FFGEN**  \L1_0/sum_reg[18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n4511 ), .force_10(n5109), .force_11(
        1'b0), .Q(out_L1[18]), .QN(n38558) );
  \**FFGEN**  \L1_0/sum_reg[19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L1_0/n3195 ), .force_10(n5103), .force_11(
        1'b0), .Q(out_L1[19]), .QN(n38560) );
  \**FFGEN**  \L2_0/square_reg[14][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2335 ), .force_10(\L2_0/n2336 ), 
        .force_11(1'b0), .QN(n5417) );
  \**FFGEN**  \L2_0/square_reg[14][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2339 ), .force_10(\L2_0/n2340 ), 
        .force_11(1'b0), .Q(n38278), .QN(n5418) );
  \**FFGEN**  \L2_0/square_reg[14][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2343 ), .force_10(\L2_0/n2344 ), 
        .force_11(1'b0), .QN(n5419) );
  \**FFGEN**  \L2_0/square_reg[14][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2347 ), .force_10(\L2_0/n2348 ), 
        .force_11(1'b0), .Q(n38440), .QN(n5420) );
  \**FFGEN**  \L2_0/square_reg[14][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2351 ), .force_10(\L2_0/n2352 ), 
        .force_11(1'b0), .Q(n38198), .QN(n5421) );
  \**FFGEN**  \L2_0/square_reg[14][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2355 ), .force_10(\L2_0/n2356 ), 
        .force_11(1'b0), .QN(n5422) );
  \**FFGEN**  \L2_0/square_reg[14][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2359 ), .force_10(\L2_0/n2360 ), 
        .force_11(1'b0), .Q(n38200), .QN(n5423) );
  \**FFGEN**  \L2_0/square_reg[14][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2363 ), .force_10(\L2_0/n2364 ), 
        .force_11(1'b0), .QN(n5424) );
  \**FFGEN**  \L2_0/square_reg[14][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2367 ), .force_10(\L2_0/n2368 ), 
        .force_11(1'b0), .QN(n5425) );
  \**FFGEN**  \L2_0/square_reg[14][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2371 ), .force_10(\L2_0/n2372 ), 
        .force_11(1'b0), .QN(n5426) );
  \**FFGEN**  \L2_0/square_reg[14][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2375 ), .force_10(\L2_0/n2376 ), 
        .force_11(1'b0), .QN(n5427) );
  \**FFGEN**  \L2_0/square_reg[14][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2379 ), .force_10(\L2_0/n2380 ), 
        .force_11(1'b0), .QN(n5428) );
  \**FFGEN**  \L2_0/square_reg[14][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2383 ), .force_10(\L2_0/n2384 ), 
        .force_11(1'b0), .QN(n5429) );
  \**FFGEN**  \L2_0/square_reg[14][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2387 ), .force_10(\L2_0/n2388 ), 
        .force_11(1'b0), .QN(n5430) );
  \**FFGEN**  \L2_0/square_reg[14][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2391 ), .force_10(\L2_0/n2392 ), 
        .force_11(1'b0), .QN(n5431) );
  \**FFGEN**  \L2_0/square_reg[14][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2395 ), .force_10(\L2_0/n2396 ), 
        .force_11(1'b0), .QN(n5432) );
  \**FFGEN**  \L2_0/square_reg[14][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2399 ), .force_10(\L2_0/n2400 ), 
        .force_11(1'b0), .Q(n38131), .QN(n5433) );
  \**FFGEN**  \L2_0/square_reg[14][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2403 ), .force_10(\L2_0/n2404 ), 
        .force_11(1'b0), .QN(n5434) );
  \**FFGEN**  \L2_0/square_reg[14][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n41261), .force_10(1'b0), .force_11(1'b0), 
        .Q(n38172), .QN(n5435) );
  \**FFGEN**  \L2_0/square_reg[14][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2411 ), .force_10(\L2_0/n2412 ), 
        .force_11(1'b0), .Q(n38597), .QN(n5702) );
  \**FFGEN**  \L2_0/square_reg[13][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2415 ), .force_10(\L2_0/n2416 ), 
        .force_11(1'b0), .QN(n5436) );
  \**FFGEN**  \L2_0/square_reg[13][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2419 ), .force_10(\L2_0/n2420 ), 
        .force_11(1'b0), .Q(n38269), .QN(n5437) );
  \**FFGEN**  \L2_0/square_reg[13][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2423 ), .force_10(\L2_0/n2424 ), 
        .force_11(1'b0), .QN(n5438) );
  \**FFGEN**  \L2_0/square_reg[13][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2427 ), .force_10(\L2_0/n2428 ), 
        .force_11(1'b0), .QN(n5439) );
  \**FFGEN**  \L2_0/square_reg[13][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2431 ), .force_10(\L2_0/n2432 ), 
        .force_11(1'b0), .QN(n5440) );
  \**FFGEN**  \L2_0/square_reg[13][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2435 ), .force_10(\L2_0/n2436 ), 
        .force_11(1'b0), .Q(n38532), .QN(n5441) );
  \**FFGEN**  \L2_0/square_reg[13][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2439 ), .force_10(\L2_0/n2440 ), 
        .force_11(1'b0), .Q(n38535), .QN(n5442) );
  \**FFGEN**  \L2_0/square_reg[13][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2443 ), .force_10(\L2_0/n2444 ), 
        .force_11(1'b0), .Q(n38227), .QN(n5443) );
  \**FFGEN**  \L2_0/square_reg[13][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2447 ), .force_10(\L2_0/n2448 ), 
        .force_11(1'b0), .Q(n38228), .QN(n5444) );
  \**FFGEN**  \L2_0/square_reg[13][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2451 ), .force_10(\L2_0/n2452 ), 
        .force_11(1'b0), .Q(n38229), .QN(n5445) );
  \**FFGEN**  \L2_0/square_reg[13][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2455 ), .force_10(\L2_0/n2456 ), 
        .force_11(1'b0), .Q(n38230), .QN(n5446) );
  \**FFGEN**  \L2_0/square_reg[13][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2459 ), .force_10(\L2_0/n2460 ), 
        .force_11(1'b0), .Q(n38231), .QN(n5447) );
  \**FFGEN**  \L2_0/square_reg[13][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2463 ), .force_10(\L2_0/n2464 ), 
        .force_11(1'b0), .Q(n38232), .QN(n5448) );
  \**FFGEN**  \L2_0/square_reg[13][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2467 ), .force_10(\L2_0/n2468 ), 
        .force_11(1'b0), .Q(n38233), .QN(n5449) );
  \**FFGEN**  \L2_0/square_reg[13][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2471 ), .force_10(\L2_0/n2472 ), 
        .force_11(1'b0), .Q(n38234), .QN(n5450) );
  \**FFGEN**  \L2_0/square_reg[13][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2475 ), .force_10(\L2_0/n2476 ), 
        .force_11(1'b0), .Q(n38235), .QN(n5451) );
  \**FFGEN**  \L2_0/square_reg[13][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2479 ), .force_10(\L2_0/n2480 ), 
        .force_11(1'b0), .Q(n38204), .QN(n5452) );
  \**FFGEN**  \L2_0/square_reg[13][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2483 ), .force_10(\L2_0/n2484 ), 
        .force_11(1'b0), .QN(n5453) );
  \**FFGEN**  \L2_0/square_reg[13][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n41118), .force_10(1'b0), .force_11(1'b0), 
        .Q(n38153), .QN(n5454) );
  \**FFGEN**  \L2_0/square_reg[13][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2491 ), .force_10(\L2_0/n2492 ), 
        .force_11(1'b0), .Q(n38146), .QN(n5716) );
  \**FFGEN**  \L2_0/square_reg[12][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2495 ), .force_10(\L2_0/n2496 ), 
        .force_11(1'b0), .QN(n5455) );
  \**FFGEN**  \L2_0/square_reg[12][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2499 ), .force_10(\L2_0/n2500 ), 
        .force_11(1'b0), .Q(n38271), .QN(n5456) );
  \**FFGEN**  \L2_0/square_reg[12][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2503 ), .force_10(\L2_0/n2504 ), 
        .force_11(1'b0), .Q(n38527), .QN(n5457) );
  \**FFGEN**  \L2_0/square_reg[12][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2507 ), .force_10(\L2_0/n2508 ), 
        .force_11(1'b0), .Q(n38195), .QN(n5458) );
  \**FFGEN**  \L2_0/square_reg[12][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2511 ), .force_10(\L2_0/n2512 ), 
        .force_11(1'b0), .QN(n5459) );
  \**FFGEN**  \L2_0/square_reg[12][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2515 ), .force_10(\L2_0/n2516 ), 
        .force_11(1'b0), .Q(n38438), .QN(n5460) );
  \**FFGEN**  \L2_0/square_reg[12][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2519 ), .force_10(\L2_0/n2520 ), 
        .force_11(1'b0), .QN(n5461) );
  \**FFGEN**  \L2_0/square_reg[12][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2523 ), .force_10(\L2_0/n2524 ), 
        .force_11(1'b0), .Q(n38260), .QN(n5462) );
  \**FFGEN**  \L2_0/square_reg[12][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2527 ), .force_10(\L2_0/n2528 ), 
        .force_11(1'b0), .Q(n38261), .QN(n5463) );
  \**FFGEN**  \L2_0/square_reg[12][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2531 ), .force_10(\L2_0/n2532 ), 
        .force_11(1'b0), .Q(n38262), .QN(n5464) );
  \**FFGEN**  \L2_0/square_reg[12][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2535 ), .force_10(\L2_0/n2536 ), 
        .force_11(1'b0), .Q(n38263), .QN(n5465) );
  \**FFGEN**  \L2_0/square_reg[12][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2539 ), .force_10(\L2_0/n2540 ), 
        .force_11(1'b0), .Q(n38264), .QN(n5466) );
  \**FFGEN**  \L2_0/square_reg[12][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2543 ), .force_10(\L2_0/n2544 ), 
        .force_11(1'b0), .Q(n38265), .QN(n5467) );
  \**FFGEN**  \L2_0/square_reg[12][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2547 ), .force_10(\L2_0/n2548 ), 
        .force_11(1'b0), .Q(n38266), .QN(n5468) );
  \**FFGEN**  \L2_0/square_reg[12][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2551 ), .force_10(\L2_0/n2552 ), 
        .force_11(1'b0), .Q(n38267), .QN(n5469) );
  \**FFGEN**  \L2_0/square_reg[12][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2555 ), .force_10(\L2_0/n2556 ), 
        .force_11(1'b0), .Q(n38238), .QN(n5470) );
  \**FFGEN**  \L2_0/square_reg[12][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2559 ), .force_10(\L2_0/n2560 ), 
        .force_11(1'b0), .QN(n5471) );
  \**FFGEN**  \L2_0/square_reg[12][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2563 ), .force_10(\L2_0/n2564 ), 
        .force_11(1'b0), .Q(n38531), .QN(n5472) );
  \**FFGEN**  \L2_0/square_reg[12][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n41216), .force_10(1'b0), .force_11(1'b0), 
        .Q(n38175), .QN(n5473) );
  \**FFGEN**  \L2_0/square_reg[12][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2571 ), .force_10(\L2_0/n2572 ), 
        .force_11(1'b0), .Q(n38139), .QN(n5715) );
  \**FFGEN**  \L2_0/square_reg[11][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2575 ), .force_10(\L2_0/n2576 ), 
        .force_11(1'b0), .QN(n5474) );
  \**FFGEN**  \L2_0/square_reg[11][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2579 ), .force_10(\L2_0/n2580 ), 
        .force_11(1'b0), .Q(n38277), .QN(n5475) );
  \**FFGEN**  \L2_0/square_reg[11][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2583 ), .force_10(\L2_0/n2584 ), 
        .force_11(1'b0), .QN(n5476) );
  \**FFGEN**  \L2_0/square_reg[11][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2587 ), .force_10(\L2_0/n2588 ), 
        .force_11(1'b0), .Q(n38526), .QN(n5477) );
  \**FFGEN**  \L2_0/square_reg[11][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2591 ), .force_10(\L2_0/n2592 ), 
        .force_11(1'b0), .QN(n5478) );
  \**FFGEN**  \L2_0/square_reg[11][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2595 ), .force_10(\L2_0/n2596 ), 
        .force_11(1'b0), .QN(n5479) );
  \**FFGEN**  \L2_0/square_reg[11][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2599 ), .force_10(\L2_0/n2600 ), 
        .force_11(1'b0), .Q(n38536), .QN(n5480) );
  \**FFGEN**  \L2_0/square_reg[11][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2603 ), .force_10(\L2_0/n2604 ), 
        .force_11(1'b0), .Q(n38583) );
  \**FFGEN**  \L2_0/square_reg[11][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2607 ), .force_10(\L2_0/n2608 ), 
        .force_11(1'b0), .Q(n38584) );
  \**FFGEN**  \L2_0/square_reg[11][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2611 ), .force_10(\L2_0/n2612 ), 
        .force_11(1'b0), .Q(n38585) );
  \**FFGEN**  \L2_0/square_reg[11][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2615 ), .force_10(\L2_0/n2616 ), 
        .force_11(1'b0), .Q(n38586) );
  \**FFGEN**  \L2_0/square_reg[11][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2619 ), .force_10(\L2_0/n2620 ), 
        .force_11(1'b0), .Q(n38587) );
  \**FFGEN**  \L2_0/square_reg[11][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2623 ), .force_10(\L2_0/n2624 ), 
        .force_11(1'b0), .Q(n38588) );
  \**FFGEN**  \L2_0/square_reg[11][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2627 ), .force_10(\L2_0/n2628 ), 
        .force_11(1'b0), .Q(n38589) );
  \**FFGEN**  \L2_0/square_reg[11][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2631 ), .force_10(\L2_0/n2632 ), 
        .force_11(1'b0), .Q(n38590) );
  \**FFGEN**  \L2_0/square_reg[11][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2635 ), .force_10(\L2_0/n2636 ), 
        .force_11(1'b0), .Q(n38593) );
  \**FFGEN**  \L2_0/square_reg[11][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2639 ), .force_10(\L2_0/n2640 ), 
        .force_11(1'b0), .QN(n5490) );
  \**FFGEN**  \L2_0/square_reg[11][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2643 ), .force_10(\L2_0/n2644 ), 
        .force_11(1'b0), .QN(n5491) );
  \**FFGEN**  \L2_0/square_reg[11][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n39132), .force_10(1'b0), .force_11(1'b0), 
        .Q(n38152), .QN(n5492) );
  \**FFGEN**  \L2_0/square_reg[11][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2651 ), .force_10(\L2_0/n2652 ), 
        .force_11(1'b0), .Q(n38144), .QN(n5714) );
  \**FFGEN**  \L2_0/square_reg[10][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2655 ), .force_10(\L2_0/n2656 ), 
        .force_11(1'b0), .QN(n5493) );
  \**FFGEN**  \L2_0/square_reg[10][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2659 ), .force_10(\L2_0/n2660 ), 
        .force_11(1'b0), .Q(n38273), .QN(n5494) );
  \**FFGEN**  \L2_0/square_reg[10][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2663 ), .force_10(\L2_0/n2664 ), 
        .force_11(1'b0), .Q(n38595) );
  \**FFGEN**  \L2_0/square_reg[10][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2667 ), .force_10(\L2_0/n2668 ), 
        .force_11(1'b0), .QN(n5496) );
  \**FFGEN**  \L2_0/square_reg[10][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2671 ), .force_10(\L2_0/n2672 ), 
        .force_11(1'b0), .Q(n38530), .QN(n5497) );
  \**FFGEN**  \L2_0/square_reg[10][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2675 ), .force_10(\L2_0/n2676 ), 
        .force_11(1'b0), .Q(n38194), .QN(n5498) );
  \**FFGEN**  \L2_0/square_reg[10][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2679 ), .force_10(\L2_0/n2680 ), 
        .force_11(1'b0), .Q(n38556), .QN(n5499) );
  \**FFGEN**  \L2_0/square_reg[10][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2683 ), .force_10(\L2_0/n2684 ), 
        .force_11(1'b0), .QN(n5500) );
  \**FFGEN**  \L2_0/square_reg[10][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2687 ), .force_10(\L2_0/n2688 ), 
        .force_11(1'b0), .QN(n5501) );
  \**FFGEN**  \L2_0/square_reg[10][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2691 ), .force_10(\L2_0/n2692 ), 
        .force_11(1'b0), .QN(n5502) );
  \**FFGEN**  \L2_0/square_reg[10][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2695 ), .force_10(\L2_0/n2696 ), 
        .force_11(1'b0), .QN(n5503) );
  \**FFGEN**  \L2_0/square_reg[10][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2699 ), .force_10(\L2_0/n2700 ), 
        .force_11(1'b0), .QN(n5504) );
  \**FFGEN**  \L2_0/square_reg[10][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2703 ), .force_10(\L2_0/n2704 ), 
        .force_11(1'b0), .QN(n5505) );
  \**FFGEN**  \L2_0/square_reg[10][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2707 ), .force_10(\L2_0/n2708 ), 
        .force_11(1'b0), .QN(n5506) );
  \**FFGEN**  \L2_0/square_reg[10][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2711 ), .force_10(\L2_0/n2712 ), 
        .force_11(1'b0), .QN(n5507) );
  \**FFGEN**  \L2_0/square_reg[10][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2715 ), .force_10(\L2_0/n2716 ), 
        .force_11(1'b0), .QN(n5508) );
  \**FFGEN**  \L2_0/square_reg[10][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2719 ), .force_10(\L2_0/n2720 ), 
        .force_11(1'b0), .Q(n38130), .QN(n5509) );
  \**FFGEN**  \L2_0/square_reg[10][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2723 ), .force_10(\L2_0/n2724 ), 
        .force_11(1'b0), .QN(n5510) );
  \**FFGEN**  \L2_0/square_reg[10][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n41231), .force_10(1'b0), .force_11(1'b0), 
        .Q(n38170), .QN(n5511) );
  \**FFGEN**  \L2_0/square_reg[10][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2731 ), .force_10(\L2_0/n2732 ), 
        .force_11(1'b0), .Q(n38138), .QN(n5713) );
  \**FFGEN**  \L2_0/square_reg[9][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2735 ), .force_10(\L2_0/n2736 ), 
        .force_11(1'b0), .QN(n5512) );
  \**FFGEN**  \L2_0/square_reg[9][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2739 ), .force_10(\L2_0/n2740 ), 
        .force_11(1'b0), .Q(n38272), .QN(n5513) );
  \**FFGEN**  \L2_0/square_reg[9][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2743 ), .force_10(\L2_0/n2744 ), 
        .force_11(1'b0), .Q(n38538), .QN(n5514) );
  \**FFGEN**  \L2_0/square_reg[9][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2747 ), .force_10(\L2_0/n2748 ), 
        .force_11(1'b0), .Q(n38594) );
  \**FFGEN**  \L2_0/square_reg[9][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2751 ), .force_10(\L2_0/n2752 ), 
        .force_11(1'b0), .QN(n5516) );
  \**FFGEN**  \L2_0/square_reg[9][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2755 ), .force_10(\L2_0/n2756 ), 
        .force_11(1'b0), .Q(n38525), .QN(n5517) );
  \**FFGEN**  \L2_0/square_reg[9][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2759 ), .force_10(\L2_0/n2760 ), 
        .force_11(1'b0), .QN(n5518) );
  \**FFGEN**  \L2_0/square_reg[9][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2763 ), .force_10(\L2_0/n2764 ), 
        .force_11(1'b0), .Q(n38218), .QN(n5519) );
  \**FFGEN**  \L2_0/square_reg[9][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2767 ), .force_10(\L2_0/n2768 ), 
        .force_11(1'b0), .Q(n38219), .QN(n5520) );
  \**FFGEN**  \L2_0/square_reg[9][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2771 ), .force_10(\L2_0/n2772 ), 
        .force_11(1'b0), .Q(n38220), .QN(n5521) );
  \**FFGEN**  \L2_0/square_reg[9][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2775 ), .force_10(\L2_0/n2776 ), 
        .force_11(1'b0), .Q(n38221), .QN(n5522) );
  \**FFGEN**  \L2_0/square_reg[9][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2779 ), .force_10(\L2_0/n2780 ), 
        .force_11(1'b0), .Q(n38222), .QN(n5523) );
  \**FFGEN**  \L2_0/square_reg[9][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2783 ), .force_10(\L2_0/n2784 ), 
        .force_11(1'b0), .Q(n38223), .QN(n5524) );
  \**FFGEN**  \L2_0/square_reg[9][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2787 ), .force_10(\L2_0/n2788 ), 
        .force_11(1'b0), .Q(n38224), .QN(n5525) );
  \**FFGEN**  \L2_0/square_reg[9][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2791 ), .force_10(\L2_0/n2792 ), 
        .force_11(1'b0), .Q(n38225), .QN(n5526) );
  \**FFGEN**  \L2_0/square_reg[9][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2795 ), .force_10(\L2_0/n2796 ), 
        .force_11(1'b0), .Q(n38226), .QN(n5527) );
  \**FFGEN**  \L2_0/square_reg[9][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2799 ), .force_10(\L2_0/n2800 ), 
        .force_11(1'b0), .Q(n38203), .QN(n5528) );
  \**FFGEN**  \L2_0/square_reg[9][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2803 ), .force_10(\L2_0/n2804 ), 
        .force_11(1'b0), .QN(n5529) );
  \**FFGEN**  \L2_0/square_reg[9][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n41226), .force_10(1'b0), .force_11(1'b0), 
        .Q(n38151), .QN(n5530) );
  \**FFGEN**  \L2_0/square_reg[9][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2811 ), .force_10(\L2_0/n2812 ), 
        .force_11(1'b0), .Q(n38143), .QN(n5712) );
  \**FFGEN**  \L2_0/square_reg[8][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2815 ), .force_10(\L2_0/n2816 ), 
        .force_11(1'b0), .QN(n5531) );
  \**FFGEN**  \L2_0/square_reg[8][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2819 ), .force_10(\L2_0/n2820 ), 
        .force_11(1'b0), .Q(n38275), .QN(n5532) );
  \**FFGEN**  \L2_0/square_reg[8][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2823 ), .force_10(\L2_0/n2824 ), 
        .force_11(1'b0), .Q(n38268), .QN(n5533) );
  \**FFGEN**  \L2_0/square_reg[8][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2827 ), .force_10(\L2_0/n2828 ), 
        .force_11(1'b0), .Q(n38537), .QN(n5534) );
  \**FFGEN**  \L2_0/square_reg[8][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2831 ), .force_10(\L2_0/n2832 ), 
        .force_11(1'b0), .Q(n38596) );
  \**FFGEN**  \L2_0/square_reg[8][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2835 ), .force_10(\L2_0/n2836 ), 
        .force_11(1'b0), .QN(n5536) );
  \**FFGEN**  \L2_0/square_reg[8][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2839 ), .force_10(\L2_0/n2840 ), 
        .force_11(1'b0), .Q(n38534), .QN(n5537) );
  \**FFGEN**  \L2_0/square_reg[8][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2843 ), .force_10(\L2_0/n2844 ), 
        .force_11(1'b0), .Q(n38252), .QN(n5538) );
  \**FFGEN**  \L2_0/square_reg[8][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2847 ), .force_10(\L2_0/n2848 ), 
        .force_11(1'b0), .Q(n38253), .QN(n5539) );
  \**FFGEN**  \L2_0/square_reg[8][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2851 ), .force_10(\L2_0/n2852 ), 
        .force_11(1'b0), .Q(n38254), .QN(n5540) );
  \**FFGEN**  \L2_0/square_reg[8][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2855 ), .force_10(\L2_0/n2856 ), 
        .force_11(1'b0), .Q(n38255), .QN(n5541) );
  \**FFGEN**  \L2_0/square_reg[8][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2859 ), .force_10(\L2_0/n2860 ), 
        .force_11(1'b0), .Q(n38256), .QN(n5542) );
  \**FFGEN**  \L2_0/square_reg[8][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2863 ), .force_10(\L2_0/n2864 ), 
        .force_11(1'b0), .Q(n38257), .QN(n5543) );
  \**FFGEN**  \L2_0/square_reg[8][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2867 ), .force_10(\L2_0/n2868 ), 
        .force_11(1'b0), .Q(n38258), .QN(n5544) );
  \**FFGEN**  \L2_0/square_reg[8][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2871 ), .force_10(\L2_0/n2872 ), 
        .force_11(1'b0), .Q(n38259), .QN(n5545) );
  \**FFGEN**  \L2_0/square_reg[8][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2875 ), .force_10(\L2_0/n2876 ), 
        .force_11(1'b0), .Q(n38237), .QN(n5546) );
  \**FFGEN**  \L2_0/square_reg[8][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2879 ), .force_10(\L2_0/n2880 ), 
        .force_11(1'b0), .QN(n5547) );
  \**FFGEN**  \L2_0/square_reg[8][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2883 ), .force_10(\L2_0/n2884 ), 
        .force_11(1'b0), .Q(n38529), .QN(n5548) );
  \**FFGEN**  \L2_0/square_reg[8][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n41241), .force_10(1'b0), .force_11(1'b0), 
        .Q(n38174), .QN(n5549) );
  \**FFGEN**  \L2_0/square_reg[8][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2891 ), .force_10(\L2_0/n2892 ), 
        .force_11(1'b0), .Q(n38137), .QN(n5711) );
  \**FFGEN**  \L2_0/square_reg[7][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2895 ), .force_10(\L2_0/n2896 ), 
        .force_11(1'b0), .QN(n5550) );
  \**FFGEN**  \L2_0/square_reg[7][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2899 ), .force_10(\L2_0/n2900 ), 
        .force_11(1'b0), .Q(n38276), .QN(n5551) );
  \**FFGEN**  \L2_0/square_reg[7][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2903 ), .force_10(\L2_0/n2904 ), 
        .force_11(1'b0), .Q(n38540), .QN(n5552) );
  \**FFGEN**  \L2_0/square_reg[7][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2907 ), .force_10(\L2_0/n2908 ), 
        .force_11(1'b0), .QN(n5553) );
  \**FFGEN**  \L2_0/square_reg[7][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2911 ), .force_10(\L2_0/n2912 ), 
        .force_11(1'b0), .QN(n5554) );
  \**FFGEN**  \L2_0/square_reg[7][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2915 ), .force_10(\L2_0/n2916 ), 
        .force_11(1'b0), .QN(n5555) );
  \**FFGEN**  \L2_0/square_reg[7][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2919 ), .force_10(\L2_0/n2920 ), 
        .force_11(1'b0), .QN(n5556) );
  \**FFGEN**  \L2_0/square_reg[7][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2923 ), .force_10(\L2_0/n2924 ), 
        .force_11(1'b0), .Q(n38575) );
  \**FFGEN**  \L2_0/square_reg[7][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2927 ), .force_10(\L2_0/n2928 ), 
        .force_11(1'b0), .Q(n38576) );
  \**FFGEN**  \L2_0/square_reg[7][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2931 ), .force_10(\L2_0/n2932 ), 
        .force_11(1'b0), .Q(n38577) );
  \**FFGEN**  \L2_0/square_reg[7][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2935 ), .force_10(\L2_0/n2936 ), 
        .force_11(1'b0), .Q(n38578) );
  \**FFGEN**  \L2_0/square_reg[7][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2939 ), .force_10(\L2_0/n2940 ), 
        .force_11(1'b0), .Q(n38579) );
  \**FFGEN**  \L2_0/square_reg[7][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2943 ), .force_10(\L2_0/n2944 ), 
        .force_11(1'b0), .Q(n38580) );
  \**FFGEN**  \L2_0/square_reg[7][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2947 ), .force_10(\L2_0/n2948 ), 
        .force_11(1'b0), .Q(n38581) );
  \**FFGEN**  \L2_0/square_reg[7][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2951 ), .force_10(\L2_0/n2952 ), 
        .force_11(1'b0), .Q(n38582) );
  \**FFGEN**  \L2_0/square_reg[7][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2955 ), .force_10(\L2_0/n2956 ), 
        .force_11(1'b0), .Q(n38592) );
  \**FFGEN**  \L2_0/square_reg[7][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2959 ), .force_10(\L2_0/n2960 ), 
        .force_11(1'b0), .QN(n5566) );
  \**FFGEN**  \L2_0/square_reg[7][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2963 ), .force_10(\L2_0/n2964 ), 
        .force_11(1'b0), .QN(n5567) );
  \**FFGEN**  \L2_0/square_reg[7][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n41256), .force_10(1'b0), .force_11(1'b0), 
        .Q(n38150), .QN(n5568) );
  \**FFGEN**  \L2_0/square_reg[7][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2971 ), .force_10(\L2_0/n2972 ), 
        .force_11(1'b0), .Q(n38142), .QN(n5710) );
  \**FFGEN**  \L2_0/square_reg[6][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2975 ), .force_10(\L2_0/n2976 ), 
        .force_11(1'b0), .QN(n5569) );
  \**FFGEN**  \L2_0/square_reg[6][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2979 ), .force_10(\L2_0/n2980 ), 
        .force_11(1'b0), .QN(n5570) );
  \**FFGEN**  \L2_0/square_reg[6][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2983 ), .force_10(\L2_0/n2984 ), 
        .force_11(1'b0), .QN(n5571) );
  \**FFGEN**  \L2_0/square_reg[6][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2987 ), .force_10(\L2_0/n2988 ), 
        .force_11(1'b0), .Q(n38199), .QN(n5572) );
  \**FFGEN**  \L2_0/square_reg[6][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2991 ), .force_10(\L2_0/n2992 ), 
        .force_11(1'b0), .QN(n5573) );
  \**FFGEN**  \L2_0/square_reg[6][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2995 ), .force_10(\L2_0/n2996 ), 
        .force_11(1'b0), .QN(n5574) );
  \**FFGEN**  \L2_0/square_reg[6][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n2999 ), .force_10(\L2_0/n3000 ), 
        .force_11(1'b0), .QN(n5575) );
  \**FFGEN**  \L2_0/square_reg[6][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3003 ), .force_10(\L2_0/n3004 ), 
        .force_11(1'b0), .QN(n5576) );
  \**FFGEN**  \L2_0/square_reg[6][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3007 ), .force_10(\L2_0/n3008 ), 
        .force_11(1'b0), .QN(n5577) );
  \**FFGEN**  \L2_0/square_reg[6][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3011 ), .force_10(\L2_0/n3012 ), 
        .force_11(1'b0), .QN(n5578) );
  \**FFGEN**  \L2_0/square_reg[6][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3015 ), .force_10(\L2_0/n3016 ), 
        .force_11(1'b0), .QN(n5579) );
  \**FFGEN**  \L2_0/square_reg[6][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3019 ), .force_10(\L2_0/n3020 ), 
        .force_11(1'b0), .QN(n5580) );
  \**FFGEN**  \L2_0/square_reg[6][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3023 ), .force_10(\L2_0/n3024 ), 
        .force_11(1'b0), .QN(n5581) );
  \**FFGEN**  \L2_0/square_reg[6][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3027 ), .force_10(\L2_0/n3028 ), 
        .force_11(1'b0), .QN(n5582) );
  \**FFGEN**  \L2_0/square_reg[6][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3031 ), .force_10(\L2_0/n3032 ), 
        .force_11(1'b0), .QN(n5583) );
  \**FFGEN**  \L2_0/square_reg[6][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3035 ), .force_10(\L2_0/n3036 ), 
        .force_11(1'b0), .QN(n5584) );
  \**FFGEN**  \L2_0/square_reg[6][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3039 ), .force_10(\L2_0/n3040 ), 
        .force_11(1'b0), .Q(n38129), .QN(n5585) );
  \**FFGEN**  \L2_0/square_reg[6][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3043 ), .force_10(\L2_0/n3044 ), 
        .force_11(1'b0), .QN(n5586) );
  \**FFGEN**  \L2_0/square_reg[6][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n41202), .force_10(1'b0), .force_11(1'b0), 
        .Q(n38169), .QN(n5587) );
  \**FFGEN**  \L2_0/square_reg[6][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3051 ), .force_10(\L2_0/n3052 ), 
        .force_11(1'b0), .Q(n38136), .QN(n5709) );
  \**FFGEN**  \L2_0/square_reg[5][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3055 ), .force_10(\L2_0/n3056 ), 
        .force_11(1'b0), .QN(n5588) );
  \**FFGEN**  \L2_0/square_reg[5][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3059 ), .force_10(\L2_0/n3060 ), 
        .force_11(1'b0), .Q(n38279), .QN(n5589) );
  \**FFGEN**  \L2_0/square_reg[5][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3063 ), .force_10(\L2_0/n3064 ), 
        .force_11(1'b0), .QN(n5590) );
  \**FFGEN**  \L2_0/square_reg[5][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3067 ), .force_10(\L2_0/n3068 ), 
        .force_11(1'b0), .Q(n38217), .QN(n5591) );
  \**FFGEN**  \L2_0/square_reg[5][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3071 ), .force_10(\L2_0/n3072 ), 
        .force_11(1'b0), .Q(n38216), .QN(n5592) );
  \**FFGEN**  \L2_0/square_reg[5][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3075 ), .force_10(\L2_0/n3076 ), 
        .force_11(1'b0), .Q(n38215), .QN(n5593) );
  \**FFGEN**  \L2_0/square_reg[5][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3079 ), .force_10(\L2_0/n3080 ), 
        .force_11(1'b0), .Q(n38205), .QN(n5594) );
  \**FFGEN**  \L2_0/square_reg[5][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3083 ), .force_10(\L2_0/n3084 ), 
        .force_11(1'b0), .Q(n38206), .QN(n5595) );
  \**FFGEN**  \L2_0/square_reg[5][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3087 ), .force_10(\L2_0/n3088 ), 
        .force_11(1'b0), .Q(n38207), .QN(n5596) );
  \**FFGEN**  \L2_0/square_reg[5][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3091 ), .force_10(\L2_0/n3092 ), 
        .force_11(1'b0), .Q(n38208), .QN(n5597) );
  \**FFGEN**  \L2_0/square_reg[5][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3095 ), .force_10(\L2_0/n3096 ), 
        .force_11(1'b0), .Q(n38209), .QN(n5598) );
  \**FFGEN**  \L2_0/square_reg[5][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3099 ), .force_10(\L2_0/n3100 ), 
        .force_11(1'b0), .Q(n38210), .QN(n5599) );
  \**FFGEN**  \L2_0/square_reg[5][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3103 ), .force_10(\L2_0/n3104 ), 
        .force_11(1'b0), .Q(n38211), .QN(n5600) );
  \**FFGEN**  \L2_0/square_reg[5][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3107 ), .force_10(\L2_0/n3108 ), 
        .force_11(1'b0), .Q(n38212), .QN(n5601) );
  \**FFGEN**  \L2_0/square_reg[5][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3111 ), .force_10(\L2_0/n3112 ), 
        .force_11(1'b0), .Q(n38213), .QN(n5602) );
  \**FFGEN**  \L2_0/square_reg[5][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3115 ), .force_10(\L2_0/n3116 ), 
        .force_11(1'b0), .Q(n38214), .QN(n5603) );
  \**FFGEN**  \L2_0/square_reg[5][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3119 ), .force_10(\L2_0/n3120 ), 
        .force_11(1'b0), .Q(n38202), .QN(n5604) );
  \**FFGEN**  \L2_0/square_reg[5][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3123 ), .force_10(\L2_0/n3124 ), 
        .force_11(1'b0), .QN(n5605) );
  \**FFGEN**  \L2_0/square_reg[5][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n41221), .force_10(1'b0), .force_11(1'b0), 
        .Q(n38149), .QN(n5606) );
  \**FFGEN**  \L2_0/square_reg[5][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3131 ), .force_10(\L2_0/n3132 ), 
        .force_11(1'b0), .Q(n38141), .QN(n5708) );
  \**FFGEN**  \L2_0/square_reg[4][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3135 ), .force_10(\L2_0/n3136 ), 
        .force_11(1'b0), .QN(n5607) );
  \**FFGEN**  \L2_0/square_reg[4][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3139 ), .force_10(\L2_0/n3140 ), 
        .force_11(1'b0), .Q(n38274), .QN(n5608) );
  \**FFGEN**  \L2_0/square_reg[4][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3143 ), .force_10(\L2_0/n3144 ), 
        .force_11(1'b0), .Q(n38533), .QN(n5609) );
  \**FFGEN**  \L2_0/square_reg[4][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3147 ), .force_10(\L2_0/n3148 ), 
        .force_11(1'b0), .Q(n38251), .QN(n5610) );
  \**FFGEN**  \L2_0/square_reg[4][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3151 ), .force_10(\L2_0/n3152 ), 
        .force_11(1'b0), .Q(n38250), .QN(n5611) );
  \**FFGEN**  \L2_0/square_reg[4][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3155 ), .force_10(\L2_0/n3156 ), 
        .force_11(1'b0), .Q(n38249), .QN(n5612) );
  \**FFGEN**  \L2_0/square_reg[4][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3159 ), .force_10(\L2_0/n3160 ), 
        .force_11(1'b0), .Q(n38240), .QN(n5613) );
  \**FFGEN**  \L2_0/square_reg[4][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3163 ), .force_10(\L2_0/n3164 ), 
        .force_11(1'b0), .Q(n38241), .QN(n5614) );
  \**FFGEN**  \L2_0/square_reg[4][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3167 ), .force_10(\L2_0/n3168 ), 
        .force_11(1'b0), .Q(n38242), .QN(n5615) );
  \**FFGEN**  \L2_0/square_reg[4][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3171 ), .force_10(\L2_0/n3172 ), 
        .force_11(1'b0), .Q(n38243), .QN(n5616) );
  \**FFGEN**  \L2_0/square_reg[4][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3175 ), .force_10(\L2_0/n3176 ), 
        .force_11(1'b0), .Q(n38244), .QN(n5617) );
  \**FFGEN**  \L2_0/square_reg[4][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3179 ), .force_10(\L2_0/n3180 ), 
        .force_11(1'b0), .Q(n38245), .QN(n5618) );
  \**FFGEN**  \L2_0/square_reg[4][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3183 ), .force_10(\L2_0/n3184 ), 
        .force_11(1'b0), .Q(n38246), .QN(n5619) );
  \**FFGEN**  \L2_0/square_reg[4][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3187 ), .force_10(\L2_0/n3188 ), 
        .force_11(1'b0), .Q(n38247), .QN(n5620) );
  \**FFGEN**  \L2_0/square_reg[4][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3191 ), .force_10(\L2_0/n3192 ), 
        .force_11(1'b0), .Q(n38248), .QN(n5621) );
  \**FFGEN**  \L2_0/square_reg[4][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3195 ), .force_10(\L2_0/n3196 ), 
        .force_11(1'b0), .Q(n38236), .QN(n5622) );
  \**FFGEN**  \L2_0/square_reg[4][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3199 ), .force_10(\L2_0/n3200 ), 
        .force_11(1'b0), .QN(n5623) );
  \**FFGEN**  \L2_0/square_reg[4][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3203 ), .force_10(\L2_0/n3204 ), 
        .force_11(1'b0), .Q(n38528), .QN(n5624) );
  \**FFGEN**  \L2_0/square_reg[4][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n41198), .force_10(1'b0), .force_11(1'b0), 
        .Q(n38173), .QN(n5625) );
  \**FFGEN**  \L2_0/square_reg[4][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3211 ), .force_10(\L2_0/n3212 ), 
        .force_11(1'b0), .Q(n38135), .QN(n5707) );
  \**FFGEN**  \L2_0/square_reg[3][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3215 ), .force_10(\L2_0/n3216 ), 
        .force_11(1'b0), .QN(n5626) );
  \**FFGEN**  \L2_0/square_reg[3][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3219 ), .force_10(\L2_0/n3220 ), 
        .force_11(1'b0), .Q(n38270), .QN(n5627) );
  \**FFGEN**  \L2_0/square_reg[3][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3223 ), .force_10(\L2_0/n3224 ), 
        .force_11(1'b0), .Q(n38539), .QN(n5628) );
  \**FFGEN**  \L2_0/square_reg[3][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3227 ), .force_10(\L2_0/n3228 ), 
        .force_11(1'b0), .Q(n38574) );
  \**FFGEN**  \L2_0/square_reg[3][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3231 ), .force_10(\L2_0/n3232 ), 
        .force_11(1'b0), .Q(n38573) );
  \**FFGEN**  \L2_0/square_reg[3][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3235 ), .force_10(\L2_0/n3236 ), 
        .force_11(1'b0), .Q(n38572) );
  \**FFGEN**  \L2_0/square_reg[3][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3239 ), .force_10(\L2_0/n3240 ), 
        .force_11(1'b0), .Q(n38563) );
  \**FFGEN**  \L2_0/square_reg[3][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3243 ), .force_10(\L2_0/n3244 ), 
        .force_11(1'b0), .Q(n38564) );
  \**FFGEN**  \L2_0/square_reg[3][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3247 ), .force_10(\L2_0/n3248 ), 
        .force_11(1'b0), .Q(n38565) );
  \**FFGEN**  \L2_0/square_reg[3][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3251 ), .force_10(\L2_0/n3252 ), 
        .force_11(1'b0), .Q(n38566) );
  \**FFGEN**  \L2_0/square_reg[3][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3255 ), .force_10(\L2_0/n3256 ), 
        .force_11(1'b0), .Q(n38567) );
  \**FFGEN**  \L2_0/square_reg[3][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3259 ), .force_10(\L2_0/n3260 ), 
        .force_11(1'b0), .Q(n38568) );
  \**FFGEN**  \L2_0/square_reg[3][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3263 ), .force_10(\L2_0/n3264 ), 
        .force_11(1'b0), .Q(n38569) );
  \**FFGEN**  \L2_0/square_reg[3][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3267 ), .force_10(\L2_0/n3268 ), 
        .force_11(1'b0), .Q(n38570) );
  \**FFGEN**  \L2_0/square_reg[3][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3271 ), .force_10(\L2_0/n3272 ), 
        .force_11(1'b0), .Q(n38571) );
  \**FFGEN**  \L2_0/square_reg[3][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3275 ), .force_10(\L2_0/n3276 ), 
        .force_11(1'b0), .Q(n38591) );
  \**FFGEN**  \L2_0/square_reg[3][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3279 ), .force_10(\L2_0/n3280 ), 
        .force_11(1'b0), .QN(n5642) );
  \**FFGEN**  \L2_0/square_reg[3][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3283 ), .force_10(\L2_0/n3284 ), 
        .force_11(1'b0), .QN(n5643) );
  \**FFGEN**  \L2_0/square_reg[3][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n41246), .force_10(1'b0), .force_11(1'b0), 
        .Q(n38148), .QN(n5644) );
  \**FFGEN**  \L2_0/square_reg[3][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3291 ), .force_10(\L2_0/n3292 ), 
        .force_11(1'b0), .Q(n38145), .QN(n5706) );
  \**FFGEN**  \L2_0/square_reg[2][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3295 ), .force_10(\L2_0/n3296 ), 
        .force_11(1'b0), .QN(n5645) );
  \**FFGEN**  \L2_0/square_reg[2][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3299 ), .force_10(\L2_0/n3300 ), 
        .force_11(1'b0), .Q(n38201), .QN(n5646) );
  \**FFGEN**  \L2_0/square_reg[2][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3303 ), .force_10(\L2_0/n3304 ), 
        .force_11(1'b0), .QN(n5647) );
  \**FFGEN**  \L2_0/square_reg[2][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3307 ), .force_10(\L2_0/n3308 ), 
        .force_11(1'b0), .QN(n5648) );
  \**FFGEN**  \L2_0/square_reg[2][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3311 ), .force_10(\L2_0/n3312 ), 
        .force_11(1'b0), .QN(n5649) );
  \**FFGEN**  \L2_0/square_reg[2][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3315 ), .force_10(\L2_0/n3316 ), 
        .force_11(1'b0), .QN(n5650) );
  \**FFGEN**  \L2_0/square_reg[2][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3319 ), .force_10(\L2_0/n3320 ), 
        .force_11(1'b0), .QN(n5651) );
  \**FFGEN**  \L2_0/square_reg[2][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3323 ), .force_10(\L2_0/n3324 ), 
        .force_11(1'b0), .QN(n5652) );
  \**FFGEN**  \L2_0/square_reg[2][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3327 ), .force_10(\L2_0/n3328 ), 
        .force_11(1'b0), .QN(n5653) );
  \**FFGEN**  \L2_0/square_reg[2][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3331 ), .force_10(\L2_0/n3332 ), 
        .force_11(1'b0), .QN(n5654) );
  \**FFGEN**  \L2_0/square_reg[2][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3335 ), .force_10(\L2_0/n3336 ), 
        .force_11(1'b0), .QN(n5655) );
  \**FFGEN**  \L2_0/square_reg[2][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3339 ), .force_10(\L2_0/n3340 ), 
        .force_11(1'b0), .QN(n5656) );
  \**FFGEN**  \L2_0/square_reg[2][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3343 ), .force_10(\L2_0/n3344 ), 
        .force_11(1'b0), .QN(n5657) );
  \**FFGEN**  \L2_0/square_reg[2][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3347 ), .force_10(\L2_0/n3348 ), 
        .force_11(1'b0), .QN(n5658) );
  \**FFGEN**  \L2_0/square_reg[2][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3351 ), .force_10(\L2_0/n3352 ), 
        .force_11(1'b0), .QN(n5659) );
  \**FFGEN**  \L2_0/square_reg[2][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3355 ), .force_10(\L2_0/n3356 ), 
        .force_11(1'b0), .QN(n5660) );
  \**FFGEN**  \L2_0/square_reg[2][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3359 ), .force_10(\L2_0/n3360 ), 
        .force_11(1'b0), .Q(n38132), .QN(n5661) );
  \**FFGEN**  \L2_0/square_reg[2][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3363 ), .force_10(\L2_0/n3364 ), 
        .force_11(1'b0), .QN(n5662) );
  \**FFGEN**  \L2_0/square_reg[2][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n41236), .force_10(1'b0), .force_11(1'b0), 
        .Q(n38171), .QN(n5663) );
  \**FFGEN**  \L2_0/square_reg[2][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3371 ), .force_10(\L2_0/n3372 ), 
        .force_11(1'b0), .Q(n38140), .QN(n5705) );
  \**FFGEN**  \L2_0/square_reg[1][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3375 ), .force_10(\L2_0/n3376 ), 
        .force_11(1'b0), .QN(n5664) );
  \**FFGEN**  \L2_0/square_reg[1][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3379 ), .force_10(\L2_0/n3380 ), 
        .force_11(1'b0), .Q(n38434), .QN(n5665) );
  \**FFGEN**  \L2_0/square_reg[1][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3383 ), .force_10(\L2_0/n3384 ), 
        .force_11(1'b0), .Q(n38421), .QN(n5666) );
  \**FFGEN**  \L2_0/square_reg[1][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3387 ), .force_10(\L2_0/n3388 ), 
        .force_11(1'b0), .Q(n38413), .QN(n5667) );
  \**FFGEN**  \L2_0/square_reg[1][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3391 ), .force_10(\L2_0/n3392 ), 
        .force_11(1'b0), .Q(n38441), .QN(n5668) );
  \**FFGEN**  \L2_0/square_reg[1][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3395 ), .force_10(\L2_0/n3396 ), 
        .force_11(1'b0), .Q(n38442), .QN(n5669) );
  \**FFGEN**  \L2_0/square_reg[1][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3399 ), .force_10(\L2_0/n3400 ), 
        .force_11(1'b0), .Q(n38443), .QN(n5670) );
  \**FFGEN**  \L2_0/square_reg[1][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3403 ), .force_10(\L2_0/n3404 ), 
        .force_11(1'b0), .Q(n38444), .QN(n5671) );
  \**FFGEN**  \L2_0/square_reg[1][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3407 ), .force_10(\L2_0/n3408 ), 
        .force_11(1'b0), .Q(n38445), .QN(n5672) );
  \**FFGEN**  \L2_0/square_reg[1][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3411 ), .force_10(\L2_0/n3412 ), 
        .force_11(1'b0), .Q(n38446), .QN(n5673) );
  \**FFGEN**  \L2_0/square_reg[1][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3415 ), .force_10(\L2_0/n3416 ), 
        .force_11(1'b0), .Q(n38447), .QN(n5674) );
  \**FFGEN**  \L2_0/square_reg[1][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3419 ), .force_10(\L2_0/n3420 ), 
        .force_11(1'b0), .Q(n38448), .QN(n5675) );
  \**FFGEN**  \L2_0/square_reg[1][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3423 ), .force_10(\L2_0/n3424 ), 
        .force_11(1'b0), .Q(n38449), .QN(n5676) );
  \**FFGEN**  \L2_0/square_reg[1][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3427 ), .force_10(\L2_0/n3428 ), 
        .force_11(1'b0), .Q(n38450), .QN(n5677) );
  \**FFGEN**  \L2_0/square_reg[1][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3431 ), .force_10(\L2_0/n3432 ), 
        .force_11(1'b0), .Q(n38451), .QN(n5678) );
  \**FFGEN**  \L2_0/square_reg[1][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3435 ), .force_10(\L2_0/n3436 ), 
        .force_11(1'b0), .Q(n38452), .QN(n5679) );
  \**FFGEN**  \L2_0/square_reg[1][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3439 ), .force_10(\L2_0/n3440 ), 
        .force_11(1'b0), .Q(n38439), .QN(n5680) );
  \**FFGEN**  \L2_0/square_reg[1][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3443 ), .force_10(\L2_0/n3444 ), 
        .force_11(1'b0), .Q(n38428), .QN(n5681) );
  \**FFGEN**  \L2_0/square_reg[1][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n39129), .force_10(1'b0), .force_11(1'b0), 
        .Q(n38182), .QN(n5682) );
  \**FFGEN**  \L2_0/square_reg[1][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3451 ), .force_10(\L2_0/n3452 ), 
        .force_11(1'b0), .Q(n38197), .QN(n5704) );
  \**FFGEN**  \L2_0/square_reg[0][19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3455 ), .force_10(\L2_0/n3456 ), 
        .force_11(1'b0), .QN(n5683) );
  \**FFGEN**  \L2_0/square_reg[0][18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3459 ), .force_10(\L2_0/n3460 ), 
        .force_11(1'b0), .Q(n38189), .QN(n5684) );
  \**FFGEN**  \L2_0/square_reg[0][17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3463 ), .force_10(\L2_0/n3464 ), 
        .force_11(1'b0), .Q(n42113), .QN(n5685) );
  \**FFGEN**  \L2_0/square_reg[0][16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3467 ), .force_10(\L2_0/n3468 ), 
        .force_11(1'b0), .Q(n38125) );
  \**FFGEN**  \L2_0/square_reg[0][15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3471 ), .force_10(\L2_0/n3472 ), 
        .force_11(1'b0), .Q(n38165), .QN(n5687) );
  \**FFGEN**  \L2_0/square_reg[0][14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3475 ), .force_10(\L2_0/n3476 ), 
        .force_11(1'b0), .Q(n38123) );
  \**FFGEN**  \L2_0/square_reg[0][13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3479 ), .force_10(\L2_0/n3480 ), 
        .force_11(1'b0), .Q(n38167), .QN(n5689) );
  \**FFGEN**  \L2_0/square_reg[0][12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3483 ), .force_10(\L2_0/n3484 ), 
        .force_11(1'b0), .Q(n42112), .QN(n5690) );
  \**FFGEN**  \L2_0/square_reg[0][11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3487 ), .force_10(\L2_0/n3488 ), 
        .force_11(1'b0), .Q(n38157), .QN(n5691) );
  \**FFGEN**  \L2_0/square_reg[0][10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3491 ), .force_10(\L2_0/n3492 ), 
        .force_11(1'b0), .Q(n42111), .QN(n5692) );
  \**FFGEN**  \L2_0/square_reg[0][9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3495 ), .force_10(\L2_0/n3496 ), 
        .force_11(1'b0), .Q(n38158), .QN(n5693) );
  \**FFGEN**  \L2_0/square_reg[0][8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3499 ), .force_10(\L2_0/n3500 ), 
        .force_11(1'b0), .Q(n42110), .QN(n5694) );
  \**FFGEN**  \L2_0/square_reg[0][7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3503 ), .force_10(\L2_0/n3504 ), 
        .force_11(1'b0), .Q(n38159), .QN(n5695) );
  \**FFGEN**  \L2_0/square_reg[0][6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3507 ), .force_10(\L2_0/n3508 ), 
        .force_11(1'b0), .Q(n42109), .QN(n5696) );
  \**FFGEN**  \L2_0/square_reg[0][5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3511 ), .force_10(\L2_0/n3512 ), 
        .force_11(1'b0), .Q(n38160), .QN(n5697) );
  \**FFGEN**  \L2_0/square_reg[0][4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3515 ), .force_10(\L2_0/n3516 ), 
        .force_11(1'b0), .Q(n42108), .QN(n5698) );
  \**FFGEN**  \L2_0/square_reg[0][3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3519 ), .force_10(\L2_0/n3520 ), 
        .force_11(1'b0), .Q(n38161), .QN(n5699) );
  \**FFGEN**  \L2_0/square_reg[0][2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3523 ), .force_10(\L2_0/n3524 ), 
        .force_11(1'b0), .Q(n42107), .QN(n5700) );
  \**FFGEN**  \L2_0/square_reg[0][1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n39146), .force_10(1'b0), .force_11(1'b0), 
        .Q(n41950) );
  \**FFGEN**  \L2_0/square_reg[0][0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(\L2_0/n3531 ), .force_10(\L2_0/n3532 ), 
        .force_11(1'b0), .Q(n38599), .QN(n5703) );
  \**FFGEN**  \L2_0/sum_reg[0]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n51440), .force_10(\L2_0/n3536 ), 
        .force_11(1'b0), .Q(out_L2[0]), .QN(n38561) );
  \**FFGEN**  \L2_0/sum_reg[1]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n51439), .force_10(\L2_0/n3540 ), 
        .force_11(1'b0), .Q(out_L2[1]) );
  \**FFGEN**  \L2_0/sum_reg[2]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n51438), .force_10(\L2_0/n3544 ), 
        .force_11(1'b0), .Q(out_L2[2]) );
  \**FFGEN**  \L2_0/sum_reg[3]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n51437), .force_10(\L2_0/n3548 ), 
        .force_11(1'b0), .Q(out_L2[3]), .QN(n38548) );
  \**FFGEN**  \L2_0/sum_reg[4]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n51436), .force_10(\L2_0/n3552 ), 
        .force_11(1'b0), .Q(out_L2[4]) );
  \**FFGEN**  \L2_0/sum_reg[5]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n51435), .force_10(\L2_0/n3556 ), 
        .force_11(1'b0), .Q(out_L2[5]), .QN(n38554) );
  \**FFGEN**  \L2_0/sum_reg[6]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n51434), .force_10(\L2_0/n3560 ), 
        .force_11(1'b0), .Q(out_L2[6]) );
  \**FFGEN**  \L2_0/sum_reg[7]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n51433), .force_10(\L2_0/n3564 ), 
        .force_11(1'b0), .Q(out_L2[7]), .QN(n38553) );
  \**FFGEN**  \L2_0/sum_reg[8]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n51432), .force_10(\L2_0/n3568 ), 
        .force_11(1'b0), .Q(out_L2[8]) );
  \**FFGEN**  \L2_0/sum_reg[9]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n51431), .force_10(\L2_0/n3572 ), 
        .force_11(1'b0), .Q(out_L2[9]), .QN(n38552) );
  \**FFGEN**  \L2_0/sum_reg[10]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n51430), .force_10(\L2_0/n3576 ), 
        .force_11(1'b0), .Q(out_L2[10]) );
  \**FFGEN**  \L2_0/sum_reg[11]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n51429), .force_10(\L2_0/n3580 ), 
        .force_11(1'b0), .Q(out_L2[11]), .QN(n38551) );
  \**FFGEN**  \L2_0/sum_reg[12]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n51428), .force_10(\L2_0/n3584 ), 
        .force_11(1'b0), .Q(out_L2[12]) );
  \**FFGEN**  \L2_0/sum_reg[13]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n51427), .force_10(\L2_0/n3588 ), 
        .force_11(1'b0), .Q(out_L2[13]), .QN(n38550) );
  \**FFGEN**  \L2_0/sum_reg[14]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n51426), .force_10(\L2_0/n3592 ), 
        .force_11(1'b0), .Q(out_L2[14]) );
  \**FFGEN**  \L2_0/sum_reg[15]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n51425), .force_10(\L2_0/n3596 ), 
        .force_11(1'b0), .Q(out_L2[15]), .QN(n38549) );
  \**FFGEN**  \L2_0/sum_reg[16]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n51424), .force_10(\L2_0/n3600 ), 
        .force_11(1'b0), .Q(out_L2[16]) );
  \**FFGEN**  \L2_0/sum_reg[17]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n51423), .force_10(\L2_0/n3604 ), 
        .force_11(1'b0), .Q(out_L2[17]) );
  \**FFGEN**  \L2_0/sum_reg[18]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n51422), .force_10(\L2_0/n3608 ), 
        .force_11(1'b0), .Q(out_L2[18]), .QN(n38557) );
  \**FFGEN**  \L2_0/sum_reg[19]  ( .next_state(1'b0), .clocked_on(1'b0), 
        .force_00(1'b0), .force_01(n51441), .force_10(\L2_0/n2292 ), 
        .force_11(1'b0), .Q(out_L2[19]), .QN(n41954) );
  nand_x8_sg U8642 ( .A(n21712), .B(n21713), .X(n21603) );
  nand_x8_sg U9216 ( .A(out_L2[0]), .B(n38599), .X(n21589) );
  nand_x8_sg U29640 ( .A(n29145), .B(n29266), .X(n29149) );
  nand_x8_sg U29836 ( .A(out_L1[1]), .B(n38555), .X(n29145) );
  nand_x8_sg U29974 ( .A(out_L1[0]), .B(n38598), .X(n29140) );
  inv_x1_sg U38801 ( .A(n7608), .X(n47060) );
  inv_x1_sg U38802 ( .A(n8426), .X(n47346) );
  inv_x1_sg U38803 ( .A(n9244), .X(n47631) );
  inv_x1_sg U38804 ( .A(n10064), .X(n47916) );
  inv_x1_sg U38805 ( .A(n10883), .X(n48201) );
  inv_x1_sg U38806 ( .A(n11702), .X(n48486) );
  inv_x1_sg U38807 ( .A(n12521), .X(n48771) );
  inv_x1_sg U38808 ( .A(n13340), .X(n49058) );
  inv_x1_sg U38809 ( .A(n14159), .X(n49344) );
  inv_x1_sg U38810 ( .A(n14978), .X(n49630) );
  inv_x1_sg U38811 ( .A(n15797), .X(n49916) );
  inv_x1_sg U38812 ( .A(n16616), .X(n50202) );
  inv_x1_sg U38813 ( .A(n17433), .X(n50487) );
  inv_x1_sg U38814 ( .A(n18254), .X(n50776) );
  inv_x1_sg U38815 ( .A(n19075), .X(n51063) );
  nand_x1_sg U38816 ( .A(n5529), .B(n20033), .X(n20032) );
  nand_x1_sg U38817 ( .A(n5491), .B(n19639), .X(n19638) );
  nand_x1_sg U38818 ( .A(n5643), .B(n21081), .X(n21080) );
  nand_x1_sg U38819 ( .A(n5605), .B(n20673), .X(n20672) );
  inv_x1_sg U38820 ( .A(n7396), .X(n46936) );
  inv_x1_sg U38821 ( .A(n7374), .X(n46968) );
  nand_x1_sg U38822 ( .A(n7559), .B(n7509), .X(n7558) );
  inv_x1_sg U38823 ( .A(n8214), .X(n47228) );
  inv_x1_sg U38824 ( .A(n8192), .X(n47258) );
  nand_x1_sg U38825 ( .A(n8377), .B(n8327), .X(n8376) );
  inv_x1_sg U38826 ( .A(n9032), .X(n47513) );
  inv_x1_sg U38827 ( .A(n9010), .X(n47543) );
  nand_x1_sg U38828 ( .A(n9195), .B(n9145), .X(n9194) );
  inv_x1_sg U38829 ( .A(n9852), .X(n47798) );
  inv_x1_sg U38830 ( .A(n9830), .X(n47828) );
  nand_x1_sg U38831 ( .A(n10015), .B(n9965), .X(n10014) );
  inv_x1_sg U38832 ( .A(n10671), .X(n48083) );
  inv_x1_sg U38833 ( .A(n10649), .X(n48113) );
  nand_x1_sg U38834 ( .A(n10834), .B(n10784), .X(n10833) );
  inv_x1_sg U38835 ( .A(n11490), .X(n48368) );
  inv_x1_sg U38836 ( .A(n11468), .X(n48398) );
  nand_x1_sg U38837 ( .A(n11653), .B(n11603), .X(n11652) );
  inv_x1_sg U38838 ( .A(n12309), .X(n48653) );
  inv_x1_sg U38839 ( .A(n12287), .X(n48683) );
  nand_x1_sg U38840 ( .A(n12472), .B(n12422), .X(n12471) );
  inv_x1_sg U38841 ( .A(n13128), .X(n48939) );
  inv_x1_sg U38842 ( .A(n13106), .X(n48969) );
  nand_x1_sg U38843 ( .A(n13291), .B(n13241), .X(n13290) );
  inv_x1_sg U38844 ( .A(n13947), .X(n49226) );
  inv_x1_sg U38845 ( .A(n13925), .X(n49256) );
  nand_x1_sg U38846 ( .A(n14110), .B(n14060), .X(n14109) );
  inv_x1_sg U38847 ( .A(n14766), .X(n49512) );
  inv_x1_sg U38848 ( .A(n14744), .X(n49542) );
  nand_x1_sg U38849 ( .A(n14929), .B(n14879), .X(n14928) );
  inv_x1_sg U38850 ( .A(n15585), .X(n49798) );
  inv_x1_sg U38851 ( .A(n15563), .X(n49828) );
  nand_x1_sg U38852 ( .A(n15748), .B(n15698), .X(n15747) );
  inv_x1_sg U38853 ( .A(n16404), .X(n50084) );
  inv_x1_sg U38854 ( .A(n16382), .X(n50114) );
  nand_x1_sg U38855 ( .A(n16567), .B(n16517), .X(n16566) );
  inv_x1_sg U38856 ( .A(n17221), .X(n50369) );
  inv_x1_sg U38857 ( .A(n17199), .X(n50399) );
  nand_x1_sg U38858 ( .A(n17384), .B(n17334), .X(n17383) );
  inv_x1_sg U38859 ( .A(n18042), .X(n50658) );
  inv_x1_sg U38860 ( .A(n18020), .X(n50688) );
  nand_x1_sg U38861 ( .A(n18205), .B(n18155), .X(n18204) );
  inv_x1_sg U38862 ( .A(n18863), .X(n50945) );
  inv_x1_sg U38863 ( .A(n18841), .X(n50975) );
  nand_x1_sg U38864 ( .A(n19026), .B(n18976), .X(n19025) );
  nand_x1_sg U38865 ( .A(n5459), .B(n19494), .X(n19493) );
  nand_x1_sg U38866 ( .A(n5518), .B(n20108), .X(n20107) );
  nand_x2_sg U38867 ( .A(n21706), .B(n21707), .X(n21615) );
  nand_x1_sg U38868 ( .A(out_L2[4]), .B(n21708), .X(n21707) );
  nand_x1_sg U38869 ( .A(n5698), .B(n45917), .X(n21708) );
  nand_x1_sg U38870 ( .A(n5567), .B(n20372), .X(n20371) );
  nand_x1_sg U38871 ( .A(n5453), .B(n19229), .X(n19228) );
  nand_x1_sg U38872 ( .A(n46937), .B(n7271), .X(n7293) );
  inv_x1_sg U38873 ( .A(n7400), .X(n47020) );
  nand_x1_sg U38874 ( .A(n7427), .B(n7425), .X(n7461) );
  nand_x1_sg U38875 ( .A(n46988), .B(n7468), .X(n7460) );
  nand_x1_sg U38876 ( .A(n7423), .B(n7422), .X(n7418) );
  nand_x1_sg U38877 ( .A(n47229), .B(n8090), .X(n8111) );
  inv_x1_sg U38878 ( .A(n8218), .X(n47308) );
  nand_x1_sg U38879 ( .A(n8245), .B(n8243), .X(n8279) );
  nand_x1_sg U38880 ( .A(n47277), .B(n8286), .X(n8278) );
  nand_x1_sg U38881 ( .A(n8241), .B(n8240), .X(n8236) );
  nand_x1_sg U38882 ( .A(n47514), .B(n8908), .X(n8929) );
  inv_x1_sg U38883 ( .A(n9036), .X(n47593) );
  nand_x1_sg U38884 ( .A(n9063), .B(n9061), .X(n9097) );
  nand_x1_sg U38885 ( .A(n47562), .B(n9104), .X(n9096) );
  nand_x1_sg U38886 ( .A(n9059), .B(n9058), .X(n9054) );
  nand_x1_sg U38887 ( .A(n47799), .B(n9728), .X(n9749) );
  inv_x1_sg U38888 ( .A(n9856), .X(n47878) );
  nand_x1_sg U38889 ( .A(n9883), .B(n9881), .X(n9917) );
  nand_x1_sg U38890 ( .A(n47847), .B(n9924), .X(n9916) );
  nand_x1_sg U38891 ( .A(n9879), .B(n9878), .X(n9874) );
  nand_x1_sg U38892 ( .A(n48084), .B(n10547), .X(n10568) );
  inv_x1_sg U38893 ( .A(n10675), .X(n48163) );
  nand_x1_sg U38894 ( .A(n10702), .B(n10700), .X(n10736) );
  nand_x1_sg U38895 ( .A(n48132), .B(n10743), .X(n10735) );
  nand_x1_sg U38896 ( .A(n10698), .B(n10697), .X(n10693) );
  nand_x1_sg U38897 ( .A(n48369), .B(n11366), .X(n11387) );
  inv_x1_sg U38898 ( .A(n11494), .X(n48448) );
  nand_x1_sg U38899 ( .A(n11521), .B(n11519), .X(n11555) );
  nand_x1_sg U38900 ( .A(n48417), .B(n11562), .X(n11554) );
  nand_x1_sg U38901 ( .A(n11517), .B(n11516), .X(n11512) );
  nand_x1_sg U38902 ( .A(n48654), .B(n12185), .X(n12206) );
  inv_x1_sg U38903 ( .A(n12313), .X(n48733) );
  nand_x1_sg U38904 ( .A(n12340), .B(n12338), .X(n12374) );
  nand_x1_sg U38905 ( .A(n48702), .B(n12381), .X(n12373) );
  nand_x1_sg U38906 ( .A(n12336), .B(n12335), .X(n12331) );
  nand_x1_sg U38907 ( .A(n48940), .B(n13004), .X(n13025) );
  inv_x1_sg U38908 ( .A(n13132), .X(n49019) );
  nand_x1_sg U38909 ( .A(n13159), .B(n13157), .X(n13193) );
  nand_x1_sg U38910 ( .A(n48988), .B(n13200), .X(n13192) );
  nand_x1_sg U38911 ( .A(n13155), .B(n13154), .X(n13150) );
  nand_x1_sg U38912 ( .A(n49227), .B(n13823), .X(n13844) );
  inv_x1_sg U38913 ( .A(n13951), .X(n49306) );
  nand_x1_sg U38914 ( .A(n13978), .B(n13976), .X(n14012) );
  nand_x1_sg U38915 ( .A(n49275), .B(n14019), .X(n14011) );
  nand_x1_sg U38916 ( .A(n13974), .B(n13973), .X(n13969) );
  nand_x1_sg U38917 ( .A(n49513), .B(n14642), .X(n14663) );
  inv_x1_sg U38918 ( .A(n14770), .X(n49592) );
  nand_x1_sg U38919 ( .A(n14797), .B(n14795), .X(n14831) );
  nand_x1_sg U38920 ( .A(n49561), .B(n14838), .X(n14830) );
  nand_x1_sg U38921 ( .A(n14793), .B(n14792), .X(n14788) );
  nand_x1_sg U38922 ( .A(n49799), .B(n15461), .X(n15482) );
  inv_x1_sg U38923 ( .A(n15589), .X(n49878) );
  nand_x1_sg U38924 ( .A(n15616), .B(n15614), .X(n15650) );
  nand_x1_sg U38925 ( .A(n49847), .B(n15657), .X(n15649) );
  nand_x1_sg U38926 ( .A(n15612), .B(n15611), .X(n15607) );
  nand_x1_sg U38927 ( .A(n50085), .B(n16280), .X(n16301) );
  inv_x1_sg U38928 ( .A(n16408), .X(n50164) );
  nand_x1_sg U38929 ( .A(n16435), .B(n16433), .X(n16469) );
  nand_x1_sg U38930 ( .A(n50133), .B(n16476), .X(n16468) );
  nand_x1_sg U38931 ( .A(n16431), .B(n16430), .X(n16426) );
  nand_x1_sg U38932 ( .A(n50370), .B(n17096), .X(n17118) );
  inv_x1_sg U38933 ( .A(n17226), .X(n50465) );
  nand_x1_sg U38934 ( .A(n17252), .B(n17250), .X(n17286) );
  nand_x1_sg U38935 ( .A(n50418), .B(n17293), .X(n17285) );
  nand_x1_sg U38936 ( .A(n17248), .B(n17247), .X(n17243) );
  nand_x1_sg U38937 ( .A(n50659), .B(n17918), .X(n17939) );
  inv_x1_sg U38938 ( .A(n18046), .X(n50738) );
  nand_x1_sg U38939 ( .A(n18073), .B(n18071), .X(n18107) );
  nand_x1_sg U38940 ( .A(n50707), .B(n18114), .X(n18106) );
  nand_x1_sg U38941 ( .A(n18069), .B(n18068), .X(n18064) );
  nand_x1_sg U38942 ( .A(n50946), .B(n18739), .X(n18760) );
  inv_x1_sg U38943 ( .A(n18867), .X(n51025) );
  nand_x1_sg U38944 ( .A(n18894), .B(n18892), .X(n18928) );
  nand_x1_sg U38945 ( .A(n50994), .B(n18935), .X(n18927) );
  nand_x1_sg U38946 ( .A(n18890), .B(n18889), .X(n18885) );
  inv_x1_sg U38947 ( .A(n20982), .X(n46583) );
  nand_x1_sg U38948 ( .A(n5419), .B(n6034), .X(n6033) );
  inv_x1_sg U38949 ( .A(n20947), .X(n46506) );
  inv_x1_sg U38950 ( .A(n20940), .X(n46469) );
  nand_x1_sg U38951 ( .A(n5422), .B(n6175), .X(n6174) );
  inv_x1_sg U38952 ( .A(n20933), .X(n46422) );
  inv_x1_sg U38953 ( .A(n20276), .X(n46336) );
  inv_x1_sg U38954 ( .A(n19470), .X(n46339) );
  inv_x1_sg U38955 ( .A(n20912), .X(n46287) );
  inv_x1_sg U38956 ( .A(n19463), .X(n46293) );
  inv_x1_sg U38957 ( .A(n20905), .X(n46242) );
  inv_x1_sg U38958 ( .A(n20262), .X(n46245) );
  inv_x1_sg U38959 ( .A(n19456), .X(n46248) );
  inv_x1_sg U38960 ( .A(n20898), .X(n46196) );
  inv_x1_sg U38961 ( .A(n20255), .X(n46199) );
  inv_x1_sg U38962 ( .A(n19449), .X(n46202) );
  inv_x1_sg U38963 ( .A(n19442), .X(n46157) );
  inv_x1_sg U38964 ( .A(n20891), .X(n46151) );
  inv_x1_sg U38965 ( .A(n20241), .X(n46108) );
  inv_x1_sg U38966 ( .A(n19435), .X(n46111) );
  inv_x1_sg U38967 ( .A(n20884), .X(n46105) );
  inv_x1_sg U38968 ( .A(n20234), .X(n46063) );
  inv_x1_sg U38969 ( .A(n19428), .X(n46066) );
  inv_x1_sg U38970 ( .A(n20227), .X(n46017) );
  inv_x1_sg U38971 ( .A(n19421), .X(n46020) );
  inv_x1_sg U38972 ( .A(n20870), .X(n46014) );
  inv_x1_sg U38973 ( .A(n20220), .X(n45972) );
  inv_x1_sg U38974 ( .A(n19414), .X(n45975) );
  inv_x1_sg U38975 ( .A(n20863), .X(n45969) );
  nand_x1_sg U38976 ( .A(n21428), .B(n21429), .X(n21258) );
  nand_x1_sg U38977 ( .A(n5704), .B(n45798), .X(n21429) );
  nand_x1_sg U38978 ( .A(n7125), .B(n7126), .X(n7124) );
  nand_x1_sg U38979 ( .A(n46918), .B(n7191), .X(n7203) );
  nand_x1_sg U38980 ( .A(n47061), .B(n6945), .X(n6941) );
  nand_x1_sg U38981 ( .A(n7944), .B(n7947), .X(n7945) );
  nand_x1_sg U38982 ( .A(n47210), .B(n8010), .X(n8022) );
  nand_x1_sg U38983 ( .A(n47347), .B(n7762), .X(n7758) );
  nand_x1_sg U38984 ( .A(n8762), .B(n8765), .X(n8763) );
  nand_x1_sg U38985 ( .A(n47495), .B(n8828), .X(n8840) );
  nand_x1_sg U38986 ( .A(n47632), .B(n8580), .X(n8576) );
  nand_x1_sg U38987 ( .A(n9582), .B(n9585), .X(n9583) );
  nand_x1_sg U38988 ( .A(n47780), .B(n9648), .X(n9660) );
  nand_x1_sg U38989 ( .A(n47917), .B(n9400), .X(n9396) );
  nand_x1_sg U38990 ( .A(n10401), .B(n10404), .X(n10402) );
  nand_x1_sg U38991 ( .A(n48065), .B(n10467), .X(n10479) );
  nand_x1_sg U38992 ( .A(n48202), .B(n10219), .X(n10215) );
  nand_x1_sg U38993 ( .A(n11220), .B(n11223), .X(n11221) );
  nand_x1_sg U38994 ( .A(n48350), .B(n11286), .X(n11298) );
  nand_x1_sg U38995 ( .A(n48487), .B(n11038), .X(n11034) );
  nand_x1_sg U38996 ( .A(n12039), .B(n12042), .X(n12040) );
  nand_x1_sg U38997 ( .A(n48635), .B(n12105), .X(n12117) );
  nand_x1_sg U38998 ( .A(n48772), .B(n11857), .X(n11853) );
  nand_x1_sg U38999 ( .A(n12858), .B(n12861), .X(n12859) );
  nand_x1_sg U39000 ( .A(n48921), .B(n12924), .X(n12936) );
  nand_x1_sg U39001 ( .A(n49059), .B(n12676), .X(n12672) );
  nand_x1_sg U39002 ( .A(n13677), .B(n13680), .X(n13678) );
  nand_x1_sg U39003 ( .A(n49208), .B(n13743), .X(n13755) );
  nand_x1_sg U39004 ( .A(n49345), .B(n13495), .X(n13491) );
  nand_x1_sg U39005 ( .A(n14495), .B(n14496), .X(n14494) );
  nand_x1_sg U39006 ( .A(n49494), .B(n14562), .X(n14574) );
  nand_x1_sg U39007 ( .A(n49631), .B(n14314), .X(n14310) );
  nand_x1_sg U39008 ( .A(n15314), .B(n15315), .X(n15313) );
  nand_x1_sg U39009 ( .A(n49780), .B(n15381), .X(n15393) );
  nand_x1_sg U39010 ( .A(n49917), .B(n15133), .X(n15129) );
  nand_x1_sg U39011 ( .A(n16133), .B(n16134), .X(n16132) );
  nand_x1_sg U39012 ( .A(n50066), .B(n16200), .X(n16212) );
  nand_x1_sg U39013 ( .A(n50203), .B(n15952), .X(n15948) );
  nand_x1_sg U39014 ( .A(n16950), .B(n16951), .X(n16949) );
  nand_x1_sg U39015 ( .A(n50351), .B(n17016), .X(n17028) );
  nand_x1_sg U39016 ( .A(n50488), .B(n16769), .X(n16765) );
  nand_x1_sg U39017 ( .A(n17771), .B(n17772), .X(n17770) );
  nand_x1_sg U39018 ( .A(n50640), .B(n17838), .X(n17850) );
  nand_x1_sg U39019 ( .A(n50777), .B(n17590), .X(n17586) );
  nand_x1_sg U39020 ( .A(n18592), .B(n18593), .X(n18591) );
  nand_x1_sg U39021 ( .A(n50927), .B(n18659), .X(n18671) );
  nand_x1_sg U39022 ( .A(n51064), .B(n18411), .X(n18407) );
  inv_x1_sg U39023 ( .A(n20926), .X(n46374) );
  inv_x1_sg U39024 ( .A(n20919), .X(n46333) );
  inv_x1_sg U39025 ( .A(n20269), .X(n46290) );
  inv_x1_sg U39026 ( .A(n20248), .X(n46154) );
  inv_x1_sg U39027 ( .A(n20877), .X(n46060) );
  nand_x1_sg U39028 ( .A(n23096), .B(n23097), .X(n7929) );
  nand_x1_sg U39029 ( .A(n47151), .B(n23093), .X(n23096) );
  nand_x1_sg U39030 ( .A(n8085), .B(n8086), .X(n8083) );
  nand_x1_sg U39031 ( .A(n23376), .B(n23377), .X(n8747) );
  nand_x1_sg U39032 ( .A(n47436), .B(n23373), .X(n23376) );
  nand_x1_sg U39033 ( .A(n8903), .B(n8904), .X(n8901) );
  nand_x1_sg U39034 ( .A(n23655), .B(n23656), .X(n9567) );
  nand_x1_sg U39035 ( .A(n47721), .B(n23652), .X(n23655) );
  nand_x1_sg U39036 ( .A(n9723), .B(n9724), .X(n9721) );
  nand_x1_sg U39037 ( .A(n23934), .B(n23935), .X(n10386) );
  nand_x1_sg U39038 ( .A(n48006), .B(n23931), .X(n23934) );
  nand_x1_sg U39039 ( .A(n10542), .B(n10543), .X(n10540) );
  nand_x1_sg U39040 ( .A(n24213), .B(n24214), .X(n11205) );
  nand_x1_sg U39041 ( .A(n48291), .B(n24210), .X(n24213) );
  nand_x1_sg U39042 ( .A(n11361), .B(n11362), .X(n11359) );
  nand_x1_sg U39043 ( .A(n24492), .B(n24493), .X(n12024) );
  nand_x1_sg U39044 ( .A(n48576), .B(n24489), .X(n24492) );
  nand_x1_sg U39045 ( .A(n12180), .B(n12181), .X(n12178) );
  nand_x1_sg U39046 ( .A(n24770), .B(n24771), .X(n12843) );
  nand_x1_sg U39047 ( .A(n48862), .B(n24767), .X(n24770) );
  nand_x1_sg U39048 ( .A(n12999), .B(n13000), .X(n12997) );
  nand_x1_sg U39049 ( .A(n25049), .B(n25050), .X(n13662) );
  nand_x1_sg U39050 ( .A(n49149), .B(n25046), .X(n25049) );
  nand_x1_sg U39051 ( .A(n13818), .B(n13819), .X(n13816) );
  nand_x1_sg U39052 ( .A(n25328), .B(n25329), .X(n14481) );
  nand_x1_sg U39053 ( .A(n49435), .B(n25325), .X(n25328) );
  nand_x1_sg U39054 ( .A(n14637), .B(n14638), .X(n14635) );
  nand_x1_sg U39055 ( .A(n25607), .B(n25608), .X(n15300) );
  nand_x1_sg U39056 ( .A(n49720), .B(n25604), .X(n25607) );
  nand_x1_sg U39057 ( .A(n15456), .B(n15457), .X(n15454) );
  nand_x1_sg U39058 ( .A(n25884), .B(n25885), .X(n16119) );
  nand_x1_sg U39059 ( .A(n50007), .B(n25881), .X(n25884) );
  nand_x1_sg U39060 ( .A(n16275), .B(n16276), .X(n16273) );
  nand_x1_sg U39061 ( .A(n26444), .B(n26445), .X(n17757) );
  nand_x1_sg U39062 ( .A(n50581), .B(n26441), .X(n26444) );
  nand_x1_sg U39063 ( .A(n17913), .B(n17914), .X(n17911) );
  nand_x1_sg U39064 ( .A(n26722), .B(n26723), .X(n18578) );
  nand_x1_sg U39065 ( .A(n50868), .B(n26719), .X(n26722) );
  nand_x1_sg U39066 ( .A(n18734), .B(n18735), .X(n18732) );
  inv_x1_sg U39067 ( .A(n21742), .X(n45765) );
  inv_x1_sg U39068 ( .A(n28540), .X(n45739) );
  inv_x1_sg U39069 ( .A(n26851), .X(n45753) );
  inv_x1_sg U39070 ( .A(n21789), .X(n45722) );
  inv_x1_sg U39071 ( .A(n21836), .X(n45679) );
  inv_x1_sg U39072 ( .A(n21883), .X(n45635) );
  inv_x1_sg U39073 ( .A(n21929), .X(n45591) );
  inv_x1_sg U39074 ( .A(n21976), .X(n45546) );
  inv_x1_sg U39075 ( .A(n22022), .X(n45502) );
  inv_x1_sg U39076 ( .A(n22069), .X(n45454) );
  inv_x1_sg U39077 ( .A(n22115), .X(n45410) );
  inv_x1_sg U39078 ( .A(n22163), .X(n45364) );
  inv_x1_sg U39079 ( .A(n22210), .X(n45319) );
  inv_x1_sg U39080 ( .A(n22258), .X(n45274) );
  inv_x1_sg U39081 ( .A(n22305), .X(n45229) );
  inv_x1_sg U39082 ( .A(n22353), .X(n45183) );
  inv_x1_sg U39083 ( .A(n22400), .X(n45138) );
  inv_x1_sg U39084 ( .A(n22447), .X(n45091) );
  inv_x1_sg U39085 ( .A(n22493), .X(n45047) );
  nand_x1_sg U39086 ( .A(n23042), .B(n23043), .X(n42161) );
  nand_x1_sg U39087 ( .A(n40102), .B(n23263), .X(n42376) );
  nand_x1_sg U39088 ( .A(n25553), .B(n25554), .X(n42160) );
  nand_x1_sg U39089 ( .A(n7062), .B(n6869), .X(n6876) );
  nand_x1_sg U39090 ( .A(n7059), .B(n6881), .X(n6888) );
  nand_x1_sg U39091 ( .A(n23126), .B(n47134), .X(n23124) );
  nand_x1_sg U39092 ( .A(n7880), .B(n7686), .X(n7693) );
  nand_x1_sg U39093 ( .A(n7877), .B(n7698), .X(n7705) );
  nand_x1_sg U39094 ( .A(n8698), .B(n8504), .X(n8511) );
  nand_x1_sg U39095 ( .A(n8695), .B(n8516), .X(n8523) );
  nand_x1_sg U39096 ( .A(n9518), .B(n9324), .X(n9331) );
  nand_x1_sg U39097 ( .A(n9515), .B(n9336), .X(n9343) );
  nand_x1_sg U39098 ( .A(n10337), .B(n10143), .X(n10150) );
  nand_x1_sg U39099 ( .A(n10334), .B(n10155), .X(n10162) );
  nand_x1_sg U39100 ( .A(n11156), .B(n10962), .X(n10969) );
  nand_x1_sg U39101 ( .A(n11153), .B(n10974), .X(n10981) );
  nand_x1_sg U39102 ( .A(n11975), .B(n11781), .X(n11788) );
  nand_x1_sg U39103 ( .A(n11972), .B(n11793), .X(n11800) );
  nand_x1_sg U39104 ( .A(n12794), .B(n12600), .X(n12607) );
  nand_x1_sg U39105 ( .A(n12791), .B(n12612), .X(n12619) );
  nand_x1_sg U39106 ( .A(n13613), .B(n13419), .X(n13426) );
  nand_x1_sg U39107 ( .A(n13610), .B(n13431), .X(n13438) );
  nand_x1_sg U39108 ( .A(n14432), .B(n14238), .X(n14245) );
  nand_x1_sg U39109 ( .A(n14429), .B(n14250), .X(n14257) );
  nand_x1_sg U39110 ( .A(n15251), .B(n15057), .X(n15064) );
  nand_x1_sg U39111 ( .A(n15248), .B(n15069), .X(n15076) );
  nand_x1_sg U39112 ( .A(n16070), .B(n15876), .X(n15883) );
  nand_x1_sg U39113 ( .A(n16067), .B(n15888), .X(n15895) );
  nand_x1_sg U39114 ( .A(n16889), .B(n16693), .X(n16700) );
  nand_x1_sg U39115 ( .A(n16886), .B(n16705), .X(n16712) );
  nand_x1_sg U39116 ( .A(n17708), .B(n17514), .X(n17521) );
  nand_x1_sg U39117 ( .A(n17705), .B(n17526), .X(n17533) );
  nand_x1_sg U39118 ( .A(n18529), .B(n18335), .X(n18342) );
  nand_x1_sg U39119 ( .A(n18526), .B(n18347), .X(n18354) );
  nand_x1_sg U39120 ( .A(n44967), .B(n28366), .X(n22584) );
  nand_x1_sg U39121 ( .A(n5723), .B(n22594), .X(n28366) );
  nand_x1_sg U39122 ( .A(n44974), .B(n26950), .X(n22589) );
  nand_x1_sg U39123 ( .A(n5731), .B(n22575), .X(n26950) );
  nand_x1_sg U39124 ( .A(n7365), .B(n7366), .X(n7343) );
  nand_x1_sg U39125 ( .A(n47059), .B(n7610), .X(n7608) );
  nand_x1_sg U39126 ( .A(n7616), .B(n47053), .X(n7027) );
  inv_x1_sg U39127 ( .A(n7571), .X(n47081) );
  nand_x1_sg U39128 ( .A(n8183), .B(n8184), .X(n8161) );
  nand_x1_sg U39129 ( .A(n47345), .B(n8428), .X(n8426) );
  nand_x1_sg U39130 ( .A(n8434), .B(n47340), .X(n7845) );
  inv_x1_sg U39131 ( .A(n8389), .X(n47367) );
  nand_x1_sg U39132 ( .A(n9001), .B(n9002), .X(n8979) );
  nand_x1_sg U39133 ( .A(n47630), .B(n9246), .X(n9244) );
  nand_x1_sg U39134 ( .A(n9252), .B(n47625), .X(n8663) );
  inv_x1_sg U39135 ( .A(n9207), .X(n47652) );
  nand_x1_sg U39136 ( .A(n9821), .B(n9822), .X(n9799) );
  nand_x1_sg U39137 ( .A(n47915), .B(n10066), .X(n10064) );
  nand_x1_sg U39138 ( .A(n10072), .B(n47910), .X(n9483) );
  inv_x1_sg U39139 ( .A(n10027), .X(n47937) );
  nand_x1_sg U39140 ( .A(n10640), .B(n10641), .X(n10618) );
  nand_x1_sg U39141 ( .A(n48200), .B(n10885), .X(n10883) );
  nand_x1_sg U39142 ( .A(n10891), .B(n48195), .X(n10302) );
  inv_x1_sg U39143 ( .A(n10846), .X(n48222) );
  nand_x1_sg U39144 ( .A(n11459), .B(n11460), .X(n11437) );
  nand_x1_sg U39145 ( .A(n48485), .B(n11704), .X(n11702) );
  nand_x1_sg U39146 ( .A(n11710), .B(n48480), .X(n11121) );
  inv_x1_sg U39147 ( .A(n11665), .X(n48507) );
  nand_x1_sg U39148 ( .A(n12278), .B(n12279), .X(n12256) );
  nand_x1_sg U39149 ( .A(n48770), .B(n12523), .X(n12521) );
  nand_x1_sg U39150 ( .A(n12529), .B(n48765), .X(n11940) );
  inv_x1_sg U39151 ( .A(n12484), .X(n48792) );
  nand_x1_sg U39152 ( .A(n13097), .B(n13098), .X(n13075) );
  nand_x1_sg U39153 ( .A(n49057), .B(n13342), .X(n13340) );
  nand_x1_sg U39154 ( .A(n13348), .B(n49051), .X(n12759) );
  inv_x1_sg U39155 ( .A(n13303), .X(n49079) );
  nand_x1_sg U39156 ( .A(n13916), .B(n13917), .X(n13894) );
  nand_x1_sg U39157 ( .A(n49343), .B(n14161), .X(n14159) );
  nand_x1_sg U39158 ( .A(n14167), .B(n49338), .X(n13578) );
  inv_x1_sg U39159 ( .A(n14122), .X(n49365) );
  nand_x1_sg U39160 ( .A(n14735), .B(n14736), .X(n14713) );
  nand_x1_sg U39161 ( .A(n49629), .B(n14980), .X(n14978) );
  nand_x1_sg U39162 ( .A(n14986), .B(n49624), .X(n14397) );
  inv_x1_sg U39163 ( .A(n14941), .X(n49651) );
  nand_x1_sg U39164 ( .A(n15554), .B(n15555), .X(n15532) );
  nand_x1_sg U39165 ( .A(n49915), .B(n15799), .X(n15797) );
  nand_x1_sg U39166 ( .A(n15805), .B(n49910), .X(n15216) );
  inv_x1_sg U39167 ( .A(n15760), .X(n49937) );
  nand_x1_sg U39168 ( .A(n16373), .B(n16374), .X(n16351) );
  nand_x1_sg U39169 ( .A(n50201), .B(n16618), .X(n16616) );
  nand_x1_sg U39170 ( .A(n16624), .B(n50196), .X(n16035) );
  inv_x1_sg U39171 ( .A(n16579), .X(n50223) );
  nand_x1_sg U39172 ( .A(n17190), .B(n17191), .X(n17168) );
  nand_x1_sg U39173 ( .A(n17192), .B(n16815), .X(n17191) );
  nand_x1_sg U39174 ( .A(n50486), .B(n17435), .X(n17433) );
  nand_x1_sg U39175 ( .A(n17441), .B(n50481), .X(n16854) );
  inv_x1_sg U39176 ( .A(n17396), .X(n50508) );
  nand_x1_sg U39177 ( .A(n18011), .B(n18012), .X(n17989) );
  nand_x1_sg U39178 ( .A(n50775), .B(n18256), .X(n18254) );
  nand_x1_sg U39179 ( .A(n18262), .B(n50770), .X(n17673) );
  inv_x1_sg U39180 ( .A(n18217), .X(n50797) );
  nand_x1_sg U39181 ( .A(n18832), .B(n18833), .X(n18810) );
  nand_x1_sg U39182 ( .A(n51062), .B(n19077), .X(n19075) );
  nand_x1_sg U39183 ( .A(n19083), .B(n51057), .X(n18494) );
  inv_x1_sg U39184 ( .A(n19038), .X(n51084) );
  inv_x1_sg U39185 ( .A(n20789), .X(n46578) );
  inv_x1_sg U39186 ( .A(n20957), .X(n46535) );
  nand_x1_sg U39187 ( .A(n20139), .B(n46471), .X(n19944) );
  inv_x1_sg U39188 ( .A(n20944), .X(n46455) );
  nand_x1_sg U39189 ( .A(n21023), .B(n21024), .X(n20944) );
  nand_x1_sg U39190 ( .A(n20448), .B(n46377), .X(n20309) );
  inv_x1_sg U39191 ( .A(n20937), .X(n46407) );
  nand_x1_sg U39192 ( .A(n21026), .B(n21027), .X(n20937) );
  inv_x1_sg U39193 ( .A(n20286), .X(n46351) );
  inv_x1_sg U39194 ( .A(n19704), .X(n46347) );
  inv_x1_sg U39195 ( .A(n20930), .X(n46360) );
  nand_x1_sg U39196 ( .A(n21029), .B(n21030), .X(n20930) );
  inv_x1_sg U39197 ( .A(n20923), .X(n46318) );
  nand_x1_sg U39198 ( .A(n21032), .B(n21033), .X(n20923) );
  inv_x1_sg U39199 ( .A(n20273), .X(n46264) );
  nand_x1_sg U39200 ( .A(n20326), .B(n20327), .X(n20273) );
  inv_x1_sg U39201 ( .A(n20252), .X(n46127) );
  nand_x1_sg U39202 ( .A(n20335), .B(n20336), .X(n20252) );
  inv_x1_sg U39203 ( .A(n20881), .X(n46045) );
  nand_x1_sg U39204 ( .A(n21050), .B(n21051), .X(n20881) );
  nand_x1_sg U39205 ( .A(n20195), .B(n20196), .X(n20033) );
  nand_x1_sg U39206 ( .A(n20015), .B(n20016), .X(n19844) );
  nand_x1_sg U39207 ( .A(n20354), .B(n20355), .X(n20212) );
  nand_x1_sg U39208 ( .A(n19621), .B(n19622), .X(n19406) );
  nand_x1_sg U39209 ( .A(n19828), .B(n19829), .X(n19639) );
  nand_x1_sg U39210 ( .A(n21253), .B(n21254), .X(n21081) );
  nand_x1_sg U39211 ( .A(n21063), .B(n21064), .X(n20855) );
  nand_x1_sg U39212 ( .A(n20838), .B(n20839), .X(n20673) );
  nand_x1_sg U39213 ( .A(n7392), .B(n7391), .X(n7393) );
  nand_x1_sg U39214 ( .A(n46935), .B(n7430), .X(n7396) );
  nand_x1_sg U39215 ( .A(n46987), .B(n7503), .X(n7473) );
  nand_x1_sg U39216 ( .A(n47022), .B(n7493), .X(n7464) );
  nand_x1_sg U39217 ( .A(n7549), .B(n7550), .X(n7529) );
  nand_x1_sg U39218 ( .A(n7532), .B(n7531), .X(n7525) );
  nand_x1_sg U39219 ( .A(n7480), .B(n7481), .X(n7478) );
  nand_x1_sg U39220 ( .A(n7606), .B(n7607), .X(n7540) );
  inv_x1_sg U39221 ( .A(n7541), .X(n47083) );
  nand_x1_sg U39222 ( .A(n46960), .B(n7560), .X(n7509) );
  nand_x1_sg U39223 ( .A(n7622), .B(n7623), .X(n7565) );
  nand_x1_sg U39224 ( .A(n7596), .B(n7597), .X(n7029) );
  nand_x1_sg U39225 ( .A(n7540), .B(n7541), .X(n7597) );
  nand_x1_sg U39226 ( .A(n7027), .B(n47104), .X(n7030) );
  nand_x1_sg U39227 ( .A(n39810), .B(n39350), .X(n7022) );
  inv_x1_sg U39228 ( .A(n7031), .X(n47107) );
  nand_x1_sg U39229 ( .A(n7034), .B(n7035), .X(n7033) );
  inv_x1_sg U39230 ( .A(n6987), .X(n47076) );
  nand_x1_sg U39231 ( .A(n8210), .B(n8209), .X(n8211) );
  nand_x1_sg U39232 ( .A(n47227), .B(n8248), .X(n8214) );
  nand_x1_sg U39233 ( .A(n47276), .B(n8321), .X(n8291) );
  nand_x1_sg U39234 ( .A(n47310), .B(n8311), .X(n8282) );
  nand_x1_sg U39235 ( .A(n8367), .B(n8368), .X(n8347) );
  nand_x1_sg U39236 ( .A(n8350), .B(n8349), .X(n8343) );
  nand_x1_sg U39237 ( .A(n8298), .B(n8299), .X(n8296) );
  nand_x1_sg U39238 ( .A(n8424), .B(n8425), .X(n8358) );
  inv_x1_sg U39239 ( .A(n8359), .X(n47369) );
  nand_x1_sg U39240 ( .A(n47251), .B(n8378), .X(n8327) );
  nand_x1_sg U39241 ( .A(n8440), .B(n8441), .X(n8383) );
  nand_x1_sg U39242 ( .A(n8414), .B(n8415), .X(n7847) );
  nand_x1_sg U39243 ( .A(n8358), .B(n8359), .X(n8415) );
  nand_x1_sg U39244 ( .A(n7845), .B(n47390), .X(n7848) );
  nand_x1_sg U39245 ( .A(n39813), .B(n39352), .X(n7840) );
  inv_x1_sg U39246 ( .A(n7849), .X(n47393) );
  nand_x1_sg U39247 ( .A(n7852), .B(n7853), .X(n7851) );
  inv_x1_sg U39248 ( .A(n7804), .X(n47362) );
  nand_x1_sg U39249 ( .A(n9028), .B(n9027), .X(n9029) );
  nand_x1_sg U39250 ( .A(n47512), .B(n9066), .X(n9032) );
  nand_x1_sg U39251 ( .A(n47561), .B(n9139), .X(n9109) );
  nand_x1_sg U39252 ( .A(n47595), .B(n9129), .X(n9100) );
  nand_x1_sg U39253 ( .A(n9185), .B(n9186), .X(n9165) );
  nand_x1_sg U39254 ( .A(n9168), .B(n9167), .X(n9161) );
  nand_x1_sg U39255 ( .A(n9116), .B(n9117), .X(n9114) );
  nand_x1_sg U39256 ( .A(n9242), .B(n9243), .X(n9176) );
  inv_x1_sg U39257 ( .A(n9177), .X(n47654) );
  nand_x1_sg U39258 ( .A(n47536), .B(n9196), .X(n9145) );
  nand_x1_sg U39259 ( .A(n9258), .B(n9259), .X(n9201) );
  nand_x1_sg U39260 ( .A(n9232), .B(n9233), .X(n8665) );
  nand_x1_sg U39261 ( .A(n9176), .B(n9177), .X(n9233) );
  nand_x1_sg U39262 ( .A(n8663), .B(n47675), .X(n8666) );
  nand_x1_sg U39263 ( .A(n39831), .B(n39351), .X(n8658) );
  inv_x1_sg U39264 ( .A(n8667), .X(n47678) );
  nand_x1_sg U39265 ( .A(n8670), .B(n8671), .X(n8669) );
  inv_x1_sg U39266 ( .A(n8622), .X(n47647) );
  nand_x1_sg U39267 ( .A(n9848), .B(n9847), .X(n9849) );
  nand_x1_sg U39268 ( .A(n47797), .B(n9886), .X(n9852) );
  nand_x1_sg U39269 ( .A(n47846), .B(n9959), .X(n9929) );
  nand_x1_sg U39270 ( .A(n47880), .B(n9949), .X(n9920) );
  nand_x1_sg U39271 ( .A(n10005), .B(n10006), .X(n9985) );
  nand_x1_sg U39272 ( .A(n9988), .B(n9987), .X(n9981) );
  nand_x1_sg U39273 ( .A(n9936), .B(n9937), .X(n9934) );
  nand_x1_sg U39274 ( .A(n10062), .B(n10063), .X(n9996) );
  inv_x1_sg U39275 ( .A(n9997), .X(n47939) );
  nand_x1_sg U39276 ( .A(n47821), .B(n10016), .X(n9965) );
  nand_x1_sg U39277 ( .A(n10078), .B(n10079), .X(n10021) );
  nand_x1_sg U39278 ( .A(n10052), .B(n10053), .X(n9485) );
  nand_x1_sg U39279 ( .A(n9996), .B(n9997), .X(n10053) );
  nand_x1_sg U39280 ( .A(n9483), .B(n47960), .X(n9486) );
  nand_x1_sg U39281 ( .A(n39846), .B(n39353), .X(n9478) );
  inv_x1_sg U39282 ( .A(n9487), .X(n47963) );
  nand_x1_sg U39283 ( .A(n9490), .B(n9491), .X(n9489) );
  inv_x1_sg U39284 ( .A(n9442), .X(n47932) );
  nand_x1_sg U39285 ( .A(n10667), .B(n10666), .X(n10668) );
  nand_x1_sg U39286 ( .A(n48082), .B(n10705), .X(n10671) );
  nand_x1_sg U39287 ( .A(n48131), .B(n10778), .X(n10748) );
  nand_x1_sg U39288 ( .A(n48165), .B(n10768), .X(n10739) );
  nand_x1_sg U39289 ( .A(n10824), .B(n10825), .X(n10804) );
  nand_x1_sg U39290 ( .A(n10807), .B(n10806), .X(n10800) );
  nand_x1_sg U39291 ( .A(n10755), .B(n10756), .X(n10753) );
  nand_x1_sg U39292 ( .A(n10881), .B(n10882), .X(n10815) );
  inv_x1_sg U39293 ( .A(n10816), .X(n48224) );
  nand_x1_sg U39294 ( .A(n48106), .B(n10835), .X(n10784) );
  nand_x1_sg U39295 ( .A(n10897), .B(n10898), .X(n10840) );
  nand_x1_sg U39296 ( .A(n10871), .B(n10872), .X(n10304) );
  nand_x1_sg U39297 ( .A(n10815), .B(n10816), .X(n10872) );
  nand_x1_sg U39298 ( .A(n10302), .B(n48245), .X(n10305) );
  nand_x1_sg U39299 ( .A(n39816), .B(n39355), .X(n10297) );
  inv_x1_sg U39300 ( .A(n10306), .X(n48248) );
  nand_x1_sg U39301 ( .A(n10309), .B(n10310), .X(n10308) );
  inv_x1_sg U39302 ( .A(n10261), .X(n48217) );
  nand_x1_sg U39303 ( .A(n11486), .B(n11485), .X(n11487) );
  nand_x1_sg U39304 ( .A(n48367), .B(n11524), .X(n11490) );
  nand_x1_sg U39305 ( .A(n48416), .B(n11597), .X(n11567) );
  nand_x1_sg U39306 ( .A(n48450), .B(n11587), .X(n11558) );
  nand_x1_sg U39307 ( .A(n11643), .B(n11644), .X(n11623) );
  nand_x1_sg U39308 ( .A(n11626), .B(n11625), .X(n11619) );
  nand_x1_sg U39309 ( .A(n11574), .B(n11575), .X(n11572) );
  nand_x1_sg U39310 ( .A(n11700), .B(n11701), .X(n11634) );
  inv_x1_sg U39311 ( .A(n11635), .X(n48509) );
  nand_x1_sg U39312 ( .A(n48391), .B(n11654), .X(n11603) );
  nand_x1_sg U39313 ( .A(n11716), .B(n11717), .X(n11659) );
  nand_x1_sg U39314 ( .A(n11690), .B(n11691), .X(n11123) );
  nand_x1_sg U39315 ( .A(n11634), .B(n11635), .X(n11691) );
  nand_x1_sg U39316 ( .A(n11121), .B(n48530), .X(n11124) );
  nand_x1_sg U39317 ( .A(n39834), .B(n39354), .X(n11116) );
  inv_x1_sg U39318 ( .A(n11125), .X(n48533) );
  nand_x1_sg U39319 ( .A(n11128), .B(n11129), .X(n11127) );
  inv_x1_sg U39320 ( .A(n11080), .X(n48502) );
  nand_x1_sg U39321 ( .A(n12305), .B(n12304), .X(n12306) );
  nand_x1_sg U39322 ( .A(n48652), .B(n12343), .X(n12309) );
  nand_x1_sg U39323 ( .A(n48701), .B(n12416), .X(n12386) );
  nand_x1_sg U39324 ( .A(n48735), .B(n12406), .X(n12377) );
  nand_x1_sg U39325 ( .A(n12462), .B(n12463), .X(n12442) );
  nand_x1_sg U39326 ( .A(n12445), .B(n12444), .X(n12438) );
  nand_x1_sg U39327 ( .A(n12393), .B(n12394), .X(n12391) );
  nand_x1_sg U39328 ( .A(n12519), .B(n12520), .X(n12453) );
  inv_x1_sg U39329 ( .A(n12454), .X(n48794) );
  nand_x1_sg U39330 ( .A(n48676), .B(n12473), .X(n12422) );
  nand_x1_sg U39331 ( .A(n12535), .B(n12536), .X(n12478) );
  nand_x1_sg U39332 ( .A(n12509), .B(n12510), .X(n11942) );
  nand_x1_sg U39333 ( .A(n12453), .B(n12454), .X(n12510) );
  nand_x1_sg U39334 ( .A(n11940), .B(n48815), .X(n11943) );
  nand_x1_sg U39335 ( .A(n39837), .B(n39356), .X(n11935) );
  inv_x1_sg U39336 ( .A(n11944), .X(n48818) );
  nand_x1_sg U39337 ( .A(n11947), .B(n11948), .X(n11946) );
  inv_x1_sg U39338 ( .A(n11899), .X(n48787) );
  nand_x1_sg U39339 ( .A(n13124), .B(n13123), .X(n13125) );
  nand_x1_sg U39340 ( .A(n48938), .B(n13162), .X(n13128) );
  nand_x1_sg U39341 ( .A(n48987), .B(n13235), .X(n13205) );
  nand_x1_sg U39342 ( .A(n49021), .B(n13225), .X(n13196) );
  nand_x1_sg U39343 ( .A(n13281), .B(n13282), .X(n13261) );
  nand_x1_sg U39344 ( .A(n13264), .B(n13263), .X(n13257) );
  nand_x1_sg U39345 ( .A(n13212), .B(n13213), .X(n13210) );
  nand_x1_sg U39346 ( .A(n13338), .B(n13339), .X(n13272) );
  inv_x1_sg U39347 ( .A(n13273), .X(n49081) );
  nand_x1_sg U39348 ( .A(n48962), .B(n13292), .X(n13241) );
  nand_x1_sg U39349 ( .A(n13354), .B(n13355), .X(n13297) );
  nand_x1_sg U39350 ( .A(n13328), .B(n13329), .X(n12761) );
  nand_x1_sg U39351 ( .A(n13272), .B(n13273), .X(n13329) );
  nand_x1_sg U39352 ( .A(n12759), .B(n49102), .X(n12762) );
  nand_x1_sg U39353 ( .A(n39819), .B(n39358), .X(n12754) );
  inv_x1_sg U39354 ( .A(n12763), .X(n49105) );
  nand_x1_sg U39355 ( .A(n12766), .B(n12767), .X(n12765) );
  inv_x1_sg U39356 ( .A(n12718), .X(n49074) );
  nand_x1_sg U39357 ( .A(n13943), .B(n13942), .X(n13944) );
  nand_x1_sg U39358 ( .A(n49225), .B(n13981), .X(n13947) );
  nand_x1_sg U39359 ( .A(n49274), .B(n14054), .X(n14024) );
  nand_x1_sg U39360 ( .A(n49308), .B(n14044), .X(n14015) );
  nand_x1_sg U39361 ( .A(n14100), .B(n14101), .X(n14080) );
  nand_x1_sg U39362 ( .A(n14083), .B(n14082), .X(n14076) );
  nand_x1_sg U39363 ( .A(n14031), .B(n14032), .X(n14029) );
  nand_x1_sg U39364 ( .A(n14157), .B(n14158), .X(n14091) );
  inv_x1_sg U39365 ( .A(n14092), .X(n49367) );
  nand_x1_sg U39366 ( .A(n49249), .B(n14111), .X(n14060) );
  nand_x1_sg U39367 ( .A(n14173), .B(n14174), .X(n14116) );
  nand_x1_sg U39368 ( .A(n14147), .B(n14148), .X(n13580) );
  nand_x1_sg U39369 ( .A(n14091), .B(n14092), .X(n14148) );
  nand_x1_sg U39370 ( .A(n13578), .B(n49388), .X(n13581) );
  nand_x1_sg U39371 ( .A(n39840), .B(n39357), .X(n13573) );
  inv_x1_sg U39372 ( .A(n13582), .X(n49391) );
  nand_x1_sg U39373 ( .A(n13585), .B(n13586), .X(n13584) );
  inv_x1_sg U39374 ( .A(n13537), .X(n49360) );
  nand_x1_sg U39375 ( .A(n14762), .B(n14761), .X(n14763) );
  nand_x1_sg U39376 ( .A(n49511), .B(n14800), .X(n14766) );
  nand_x1_sg U39377 ( .A(n49560), .B(n14873), .X(n14843) );
  nand_x1_sg U39378 ( .A(n49594), .B(n14863), .X(n14834) );
  nand_x1_sg U39379 ( .A(n14919), .B(n14920), .X(n14899) );
  nand_x1_sg U39380 ( .A(n14902), .B(n14901), .X(n14895) );
  nand_x1_sg U39381 ( .A(n14850), .B(n14851), .X(n14848) );
  nand_x1_sg U39382 ( .A(n14976), .B(n14977), .X(n14910) );
  inv_x1_sg U39383 ( .A(n14911), .X(n49653) );
  nand_x1_sg U39384 ( .A(n49535), .B(n14930), .X(n14879) );
  nand_x1_sg U39385 ( .A(n14992), .B(n14993), .X(n14935) );
  nand_x1_sg U39386 ( .A(n14966), .B(n14967), .X(n14399) );
  nand_x1_sg U39387 ( .A(n14910), .B(n14911), .X(n14967) );
  nand_x1_sg U39388 ( .A(n14397), .B(n49674), .X(n14400) );
  nand_x1_sg U39389 ( .A(n39843), .B(n39359), .X(n14392) );
  inv_x1_sg U39390 ( .A(n14401), .X(n49677) );
  nand_x1_sg U39391 ( .A(n14404), .B(n14405), .X(n14403) );
  inv_x1_sg U39392 ( .A(n14356), .X(n49646) );
  nand_x1_sg U39393 ( .A(n15581), .B(n15580), .X(n15582) );
  nand_x1_sg U39394 ( .A(n49797), .B(n15619), .X(n15585) );
  nand_x1_sg U39395 ( .A(n49846), .B(n15692), .X(n15662) );
  nand_x1_sg U39396 ( .A(n49880), .B(n15682), .X(n15653) );
  nand_x1_sg U39397 ( .A(n15738), .B(n15739), .X(n15718) );
  nand_x1_sg U39398 ( .A(n15721), .B(n15720), .X(n15714) );
  nand_x1_sg U39399 ( .A(n15669), .B(n15670), .X(n15667) );
  nand_x1_sg U39400 ( .A(n15795), .B(n15796), .X(n15729) );
  inv_x1_sg U39401 ( .A(n15730), .X(n49939) );
  nand_x1_sg U39402 ( .A(n49821), .B(n15749), .X(n15698) );
  nand_x1_sg U39403 ( .A(n15811), .B(n15812), .X(n15754) );
  nand_x1_sg U39404 ( .A(n15785), .B(n15786), .X(n15218) );
  nand_x1_sg U39405 ( .A(n15729), .B(n15730), .X(n15786) );
  nand_x1_sg U39406 ( .A(n15216), .B(n49960), .X(n15219) );
  nand_x1_sg U39407 ( .A(n39849), .B(n39361), .X(n15211) );
  inv_x1_sg U39408 ( .A(n15220), .X(n49963) );
  nand_x1_sg U39409 ( .A(n15223), .B(n15224), .X(n15222) );
  inv_x1_sg U39410 ( .A(n15175), .X(n49932) );
  nand_x1_sg U39411 ( .A(n16400), .B(n16399), .X(n16401) );
  nand_x1_sg U39412 ( .A(n50083), .B(n16438), .X(n16404) );
  nand_x1_sg U39413 ( .A(n50132), .B(n16511), .X(n16481) );
  nand_x1_sg U39414 ( .A(n50166), .B(n16501), .X(n16472) );
  nand_x1_sg U39415 ( .A(n16557), .B(n16558), .X(n16537) );
  nand_x1_sg U39416 ( .A(n16540), .B(n16539), .X(n16533) );
  nand_x1_sg U39417 ( .A(n16488), .B(n16489), .X(n16486) );
  nand_x1_sg U39418 ( .A(n16614), .B(n16615), .X(n16548) );
  inv_x1_sg U39419 ( .A(n16549), .X(n50225) );
  nand_x1_sg U39420 ( .A(n50107), .B(n16568), .X(n16517) );
  nand_x1_sg U39421 ( .A(n16630), .B(n16631), .X(n16573) );
  nand_x1_sg U39422 ( .A(n16604), .B(n16605), .X(n16037) );
  nand_x1_sg U39423 ( .A(n16548), .B(n16549), .X(n16605) );
  nand_x1_sg U39424 ( .A(n16035), .B(n50246), .X(n16038) );
  nand_x1_sg U39425 ( .A(n39822), .B(n39360), .X(n16030) );
  inv_x1_sg U39426 ( .A(n16039), .X(n50249) );
  nand_x1_sg U39427 ( .A(n16042), .B(n16043), .X(n16041) );
  inv_x1_sg U39428 ( .A(n15994), .X(n50218) );
  nand_x1_sg U39429 ( .A(n17217), .B(n17216), .X(n17218) );
  nand_x1_sg U39430 ( .A(n50368), .B(n17255), .X(n17221) );
  nand_x1_sg U39431 ( .A(n50417), .B(n17328), .X(n17298) );
  nand_x1_sg U39432 ( .A(n50451), .B(n17318), .X(n17289) );
  nand_x1_sg U39433 ( .A(n17374), .B(n17375), .X(n17354) );
  nand_x1_sg U39434 ( .A(n17357), .B(n17356), .X(n17350) );
  nand_x1_sg U39435 ( .A(n17305), .B(n17306), .X(n17303) );
  nand_x1_sg U39436 ( .A(n17431), .B(n17432), .X(n17365) );
  inv_x1_sg U39437 ( .A(n17366), .X(n50510) );
  nand_x1_sg U39438 ( .A(n50392), .B(n17385), .X(n17334) );
  nand_x1_sg U39439 ( .A(n17447), .B(n17448), .X(n17390) );
  nand_x1_sg U39440 ( .A(n17449), .B(n17299), .X(n17448) );
  nand_x1_sg U39441 ( .A(n17421), .B(n17422), .X(n16856) );
  nand_x1_sg U39442 ( .A(n17365), .B(n17366), .X(n17422) );
  nand_x1_sg U39443 ( .A(n16854), .B(n50531), .X(n16857) );
  nand_x1_sg U39444 ( .A(n40608), .B(n39364), .X(n16847) );
  inv_x1_sg U39445 ( .A(n16858), .X(n50534) );
  nand_x1_sg U39446 ( .A(n16861), .B(n16862), .X(n16860) );
  inv_x1_sg U39447 ( .A(n16811), .X(n50503) );
  nand_x1_sg U39448 ( .A(n18038), .B(n18037), .X(n18039) );
  nand_x1_sg U39449 ( .A(n50657), .B(n18076), .X(n18042) );
  nand_x1_sg U39450 ( .A(n50706), .B(n18149), .X(n18119) );
  nand_x1_sg U39451 ( .A(n50740), .B(n18139), .X(n18110) );
  nand_x1_sg U39452 ( .A(n18195), .B(n18196), .X(n18175) );
  nand_x1_sg U39453 ( .A(n18178), .B(n18177), .X(n18171) );
  nand_x1_sg U39454 ( .A(n18126), .B(n18127), .X(n18124) );
  nand_x1_sg U39455 ( .A(n18252), .B(n18253), .X(n18186) );
  inv_x1_sg U39456 ( .A(n18187), .X(n50799) );
  nand_x1_sg U39457 ( .A(n50681), .B(n18206), .X(n18155) );
  nand_x1_sg U39458 ( .A(n18268), .B(n18269), .X(n18211) );
  nand_x1_sg U39459 ( .A(n18242), .B(n18243), .X(n17675) );
  nand_x1_sg U39460 ( .A(n18186), .B(n18187), .X(n18243) );
  nand_x1_sg U39461 ( .A(n17673), .B(n50820), .X(n17676) );
  nand_x1_sg U39462 ( .A(n39828), .B(n39363), .X(n17668) );
  inv_x1_sg U39463 ( .A(n17677), .X(n50823) );
  nand_x1_sg U39464 ( .A(n17680), .B(n17681), .X(n17679) );
  inv_x1_sg U39465 ( .A(n17632), .X(n50792) );
  nand_x1_sg U39466 ( .A(n18859), .B(n18858), .X(n18860) );
  nand_x1_sg U39467 ( .A(n50944), .B(n18897), .X(n18863) );
  nand_x1_sg U39468 ( .A(n50993), .B(n18970), .X(n18940) );
  nand_x1_sg U39469 ( .A(n51027), .B(n18960), .X(n18931) );
  nand_x1_sg U39470 ( .A(n19016), .B(n19017), .X(n18996) );
  nand_x1_sg U39471 ( .A(n18999), .B(n18998), .X(n18992) );
  nand_x1_sg U39472 ( .A(n18947), .B(n18948), .X(n18945) );
  nand_x1_sg U39473 ( .A(n19073), .B(n19074), .X(n19007) );
  inv_x1_sg U39474 ( .A(n19008), .X(n51086) );
  nand_x1_sg U39475 ( .A(n50968), .B(n19027), .X(n18976) );
  nand_x1_sg U39476 ( .A(n19089), .B(n19090), .X(n19032) );
  nand_x1_sg U39477 ( .A(n19063), .B(n19064), .X(n18496) );
  nand_x1_sg U39478 ( .A(n19007), .B(n19008), .X(n19064) );
  nand_x1_sg U39479 ( .A(n18494), .B(n51107), .X(n18497) );
  nand_x1_sg U39480 ( .A(n39825), .B(n39362), .X(n18489) );
  inv_x1_sg U39481 ( .A(n18498), .X(n51110) );
  nand_x1_sg U39482 ( .A(n18501), .B(n18502), .X(n18500) );
  inv_x1_sg U39483 ( .A(n18453), .X(n51079) );
  nand_x1_sg U39484 ( .A(n28251), .B(n28252), .X(n28135) );
  nand_x1_sg U39485 ( .A(n20595), .B(n46553), .X(n19748) );
  inv_x1_sg U39486 ( .A(n20991), .X(n46582) );
  nand_x1_sg U39487 ( .A(n21191), .B(n21192), .X(n20991) );
  nand_x1_sg U39488 ( .A(n46515), .B(n19954), .X(n19767) );
  nand_x1_sg U39489 ( .A(n19574), .B(n19575), .X(n19507) );
  inv_x1_sg U39490 ( .A(n21194), .X(n46542) );
  nand_x1_sg U39491 ( .A(n21361), .B(n21362), .X(n21194) );
  nand_x1_sg U39492 ( .A(n20598), .B(n20599), .X(n19938) );
  nand_x1_sg U39493 ( .A(n46473), .B(n20146), .X(n19951) );
  inv_x1_sg U39494 ( .A(n21364), .X(n46500) );
  nand_x1_sg U39495 ( .A(n21543), .B(n21544), .X(n21364) );
  inv_x1_sg U39496 ( .A(n20951), .X(n46493) );
  nand_x1_sg U39497 ( .A(n21020), .B(n21021), .X(n20951) );
  inv_x1_sg U39498 ( .A(n20771), .X(n46491) );
  nand_x1_sg U39499 ( .A(n20796), .B(n20797), .X(n20771) );
  nand_x1_sg U39500 ( .A(n19967), .B(n19968), .X(n19916) );
  nand_x1_sg U39501 ( .A(n20306), .B(n46425), .X(n20142) );
  nand_x1_sg U39502 ( .A(n19580), .B(n19581), .X(n19494) );
  inv_x1_sg U39503 ( .A(n20764), .X(n46453) );
  nand_x1_sg U39504 ( .A(n20799), .B(n20800), .X(n20764) );
  inv_x1_sg U39505 ( .A(n20757), .X(n46405) );
  nand_x1_sg U39506 ( .A(n20802), .B(n20803), .X(n20757) );
  nand_x1_sg U39507 ( .A(n20162), .B(n20163), .X(n20108) );
  nand_x1_sg U39508 ( .A(n46352), .B(n20451), .X(n20437) );
  nand_x1_sg U39509 ( .A(n19587), .B(n19588), .X(n19480) );
  inv_x1_sg U39510 ( .A(n20750), .X(n46358) );
  nand_x1_sg U39511 ( .A(n20805), .B(n20806), .X(n20750) );
  inv_x1_sg U39512 ( .A(n20280), .X(n46309) );
  nand_x1_sg U39513 ( .A(n20323), .B(n20324), .X(n20280) );
  inv_x1_sg U39514 ( .A(n20103), .X(n46307) );
  nand_x1_sg U39515 ( .A(n20165), .B(n20166), .X(n20103) );
  inv_x1_sg U39516 ( .A(n19474), .X(n46300) );
  nand_x1_sg U39517 ( .A(n19590), .B(n19591), .X(n19474) );
  inv_x1_sg U39518 ( .A(n19299), .X(n46298) );
  nand_x1_sg U39519 ( .A(n19359), .B(n19360), .X(n19299) );
  inv_x1_sg U39520 ( .A(n20743), .X(n46316) );
  nand_x1_sg U39521 ( .A(n20808), .B(n20809), .X(n20743) );
  inv_x1_sg U39522 ( .A(n20916), .X(n46273) );
  nand_x1_sg U39523 ( .A(n21035), .B(n21036), .X(n20916) );
  inv_x1_sg U39524 ( .A(n20736), .X(n46271) );
  nand_x1_sg U39525 ( .A(n20811), .B(n20812), .X(n20736) );
  inv_x1_sg U39526 ( .A(n20096), .X(n46262) );
  nand_x1_sg U39527 ( .A(n20168), .B(n20169), .X(n20096) );
  inv_x1_sg U39528 ( .A(n19467), .X(n46255) );
  nand_x1_sg U39529 ( .A(n19593), .B(n19594), .X(n19467) );
  inv_x1_sg U39530 ( .A(n19292), .X(n46253) );
  nand_x1_sg U39531 ( .A(n19362), .B(n19363), .X(n19292) );
  inv_x1_sg U39532 ( .A(n20909), .X(n46227) );
  nand_x1_sg U39533 ( .A(n21038), .B(n21039), .X(n20909) );
  inv_x1_sg U39534 ( .A(n20729), .X(n46225) );
  nand_x1_sg U39535 ( .A(n20814), .B(n20815), .X(n20729) );
  inv_x1_sg U39536 ( .A(n20266), .X(n46218) );
  nand_x1_sg U39537 ( .A(n20329), .B(n20330), .X(n20266) );
  inv_x1_sg U39538 ( .A(n20089), .X(n46216) );
  nand_x1_sg U39539 ( .A(n20171), .B(n20172), .X(n20089) );
  inv_x1_sg U39540 ( .A(n19460), .X(n46209) );
  nand_x1_sg U39541 ( .A(n19596), .B(n19597), .X(n19460) );
  inv_x1_sg U39542 ( .A(n19285), .X(n46207) );
  nand_x1_sg U39543 ( .A(n19365), .B(n19366), .X(n19285) );
  inv_x1_sg U39544 ( .A(n20902), .X(n46182) );
  nand_x1_sg U39545 ( .A(n21041), .B(n21042), .X(n20902) );
  inv_x1_sg U39546 ( .A(n20722), .X(n46180) );
  nand_x1_sg U39547 ( .A(n20817), .B(n20818), .X(n20722) );
  inv_x1_sg U39548 ( .A(n20259), .X(n46173) );
  nand_x1_sg U39549 ( .A(n20332), .B(n20333), .X(n20259) );
  inv_x1_sg U39550 ( .A(n20082), .X(n46171) );
  nand_x1_sg U39551 ( .A(n20174), .B(n20175), .X(n20082) );
  inv_x1_sg U39552 ( .A(n19453), .X(n46164) );
  nand_x1_sg U39553 ( .A(n19599), .B(n19600), .X(n19453) );
  inv_x1_sg U39554 ( .A(n19278), .X(n46162) );
  nand_x1_sg U39555 ( .A(n19368), .B(n19369), .X(n19278) );
  inv_x1_sg U39556 ( .A(n20075), .X(n46125) );
  nand_x1_sg U39557 ( .A(n20177), .B(n20178), .X(n20075) );
  inv_x1_sg U39558 ( .A(n19446), .X(n46118) );
  nand_x1_sg U39559 ( .A(n19602), .B(n19603), .X(n19446) );
  inv_x1_sg U39560 ( .A(n19271), .X(n46116) );
  nand_x1_sg U39561 ( .A(n19371), .B(n19372), .X(n19271) );
  inv_x1_sg U39562 ( .A(n20895), .X(n46136) );
  nand_x1_sg U39563 ( .A(n21044), .B(n21045), .X(n20895) );
  inv_x1_sg U39564 ( .A(n20715), .X(n46134) );
  nand_x1_sg U39565 ( .A(n20820), .B(n20821), .X(n20715) );
  inv_x1_sg U39566 ( .A(n20245), .X(n46082) );
  nand_x1_sg U39567 ( .A(n20338), .B(n20339), .X(n20245) );
  inv_x1_sg U39568 ( .A(n20068), .X(n46080) );
  nand_x1_sg U39569 ( .A(n20180), .B(n20181), .X(n20068) );
  inv_x1_sg U39570 ( .A(n19439), .X(n46073) );
  nand_x1_sg U39571 ( .A(n19605), .B(n19606), .X(n19439) );
  inv_x1_sg U39572 ( .A(n19264), .X(n46071) );
  nand_x1_sg U39573 ( .A(n19374), .B(n19375), .X(n19264) );
  inv_x1_sg U39574 ( .A(n20888), .X(n46091) );
  nand_x1_sg U39575 ( .A(n21047), .B(n21048), .X(n20888) );
  inv_x1_sg U39576 ( .A(n20708), .X(n46089) );
  nand_x1_sg U39577 ( .A(n20823), .B(n20824), .X(n20708) );
  inv_x1_sg U39578 ( .A(n20238), .X(n46036) );
  nand_x1_sg U39579 ( .A(n20341), .B(n20342), .X(n20238) );
  inv_x1_sg U39580 ( .A(n20061), .X(n46034) );
  nand_x1_sg U39581 ( .A(n20183), .B(n20184), .X(n20061) );
  inv_x1_sg U39582 ( .A(n19432), .X(n46027) );
  nand_x1_sg U39583 ( .A(n19608), .B(n19609), .X(n19432) );
  inv_x1_sg U39584 ( .A(n19257), .X(n46025) );
  nand_x1_sg U39585 ( .A(n19377), .B(n19378), .X(n19257) );
  inv_x1_sg U39586 ( .A(n20701), .X(n46043) );
  nand_x1_sg U39587 ( .A(n20826), .B(n20827), .X(n20701) );
  inv_x1_sg U39588 ( .A(n20231), .X(n45991) );
  nand_x1_sg U39589 ( .A(n20344), .B(n20345), .X(n20231) );
  inv_x1_sg U39590 ( .A(n20054), .X(n45989) );
  nand_x1_sg U39591 ( .A(n20186), .B(n20187), .X(n20054) );
  inv_x1_sg U39592 ( .A(n19425), .X(n45982) );
  nand_x1_sg U39593 ( .A(n19611), .B(n19612), .X(n19425) );
  inv_x1_sg U39594 ( .A(n19250), .X(n45980) );
  nand_x1_sg U39595 ( .A(n19380), .B(n19381), .X(n19250) );
  inv_x1_sg U39596 ( .A(n20874), .X(n46000) );
  nand_x1_sg U39597 ( .A(n21053), .B(n21054), .X(n20874) );
  inv_x1_sg U39598 ( .A(n20694), .X(n45998) );
  nand_x1_sg U39599 ( .A(n20829), .B(n20830), .X(n20694) );
  inv_x1_sg U39600 ( .A(n20047), .X(n45944) );
  nand_x1_sg U39601 ( .A(n20189), .B(n20190), .X(n20047) );
  inv_x1_sg U39602 ( .A(n19243), .X(n45935) );
  nand_x1_sg U39603 ( .A(n19383), .B(n19384), .X(n19243) );
  inv_x1_sg U39604 ( .A(n20687), .X(n45953) );
  nand_x1_sg U39605 ( .A(n20832), .B(n20833), .X(n20687) );
  nand_x1_sg U39606 ( .A(n20485), .B(n20486), .X(n20372) );
  nand_x1_sg U39607 ( .A(n19389), .B(n19390), .X(n19229) );
  nand_x1_sg U39608 ( .A(n21425), .B(n21426), .X(n21270) );
  nand_x1_sg U39609 ( .A(n5681), .B(n21443), .X(n21442) );
  inv_x1_sg U39610 ( .A(n6723), .X(n45873) );
  nand_x1_sg U39611 ( .A(n20655), .B(n20656), .X(n20501) );
  nand_x1_sg U39612 ( .A(n7280), .B(n7281), .X(n7252) );
  nand_x1_sg U39613 ( .A(n7282), .B(n41902), .X(n7281) );
  nand_x1_sg U39614 ( .A(n46933), .B(n7255), .X(n7249) );
  nand_x1_sg U39615 ( .A(n46944), .B(n7301), .X(n7296) );
  nand_x1_sg U39616 ( .A(n7297), .B(n46974), .X(n7271) );
  inv_x1_sg U39617 ( .A(n7388), .X(n46959) );
  nand_x1_sg U39618 ( .A(n7335), .B(n7336), .X(n7329) );
  nand_x1_sg U39619 ( .A(n7331), .B(n7332), .X(n7309) );
  inv_x1_sg U39620 ( .A(n7333), .X(n46969) );
  nand_x1_sg U39621 ( .A(n7378), .B(n46967), .X(n7374) );
  nand_x1_sg U39622 ( .A(n7375), .B(n7376), .X(n7333) );
  nand_x1_sg U39623 ( .A(n7394), .B(n7395), .X(n7388) );
  nand_x1_sg U39624 ( .A(n7360), .B(n7361), .X(n7362) );
  nand_x1_sg U39625 ( .A(n7428), .B(n7429), .X(n7422) );
  nand_x1_sg U39626 ( .A(n7420), .B(n47019), .X(n7400) );
  nand_x1_sg U39627 ( .A(n47036), .B(n7424), .X(n7401) );
  nand_x1_sg U39628 ( .A(n7462), .B(n47023), .X(n7425) );
  nand_x1_sg U39629 ( .A(n7470), .B(n47033), .X(n7468) );
  nand_x1_sg U39630 ( .A(n7478), .B(n47064), .X(n7477) );
  nand_x1_sg U39631 ( .A(n7499), .B(n7498), .X(n7485) );
  nand_x1_sg U39632 ( .A(n7487), .B(n7488), .X(n7448) );
  nand_x1_sg U39633 ( .A(n7464), .B(n7465), .X(n7487) );
  nand_x1_sg U39634 ( .A(n7485), .B(n47028), .X(n7449) );
  nand_x1_sg U39635 ( .A(n7557), .B(n7558), .X(n7555) );
  nand_x1_sg U39636 ( .A(n7563), .B(n47050), .X(n7556) );
  nand_x1_sg U39637 ( .A(n7520), .B(n7519), .X(n7521) );
  inv_x1_sg U39638 ( .A(n7035), .X(n47082) );
  nand_x1_sg U39639 ( .A(n7594), .B(n47106), .X(n7034) );
  nand_x1_sg U39640 ( .A(n8099), .B(n8100), .X(n8071) );
  nand_x1_sg U39641 ( .A(n8101), .B(n41900), .X(n8100) );
  nand_x1_sg U39642 ( .A(n47225), .B(n8074), .X(n8068) );
  nand_x1_sg U39643 ( .A(n47235), .B(n8119), .X(n8114) );
  nand_x1_sg U39644 ( .A(n8115), .B(n47264), .X(n8090) );
  inv_x1_sg U39645 ( .A(n8206), .X(n47250) );
  nand_x1_sg U39646 ( .A(n8153), .B(n8154), .X(n8147) );
  nand_x1_sg U39647 ( .A(n8149), .B(n8150), .X(n8127) );
  inv_x1_sg U39648 ( .A(n8151), .X(n47259) );
  nand_x1_sg U39649 ( .A(n8196), .B(n47257), .X(n8192) );
  nand_x1_sg U39650 ( .A(n8193), .B(n8194), .X(n8151) );
  nand_x1_sg U39651 ( .A(n8212), .B(n8213), .X(n8206) );
  nand_x1_sg U39652 ( .A(n8178), .B(n8179), .X(n8180) );
  nand_x1_sg U39653 ( .A(n8246), .B(n8247), .X(n8240) );
  nand_x1_sg U39654 ( .A(n8238), .B(n47307), .X(n8218) );
  nand_x1_sg U39655 ( .A(n47323), .B(n8242), .X(n8219) );
  nand_x1_sg U39656 ( .A(n8280), .B(n47311), .X(n8243) );
  nand_x1_sg U39657 ( .A(n8288), .B(n47320), .X(n8286) );
  nand_x1_sg U39658 ( .A(n8296), .B(n47350), .X(n8295) );
  nand_x1_sg U39659 ( .A(n8317), .B(n8316), .X(n8303) );
  nand_x1_sg U39660 ( .A(n8305), .B(n8306), .X(n8266) );
  nand_x1_sg U39661 ( .A(n8282), .B(n8283), .X(n8305) );
  nand_x1_sg U39662 ( .A(n8303), .B(n47315), .X(n8267) );
  nand_x1_sg U39663 ( .A(n8375), .B(n8376), .X(n8373) );
  nand_x1_sg U39664 ( .A(n8381), .B(n47337), .X(n8374) );
  nand_x1_sg U39665 ( .A(n8338), .B(n8337), .X(n8339) );
  inv_x1_sg U39666 ( .A(n7853), .X(n47368) );
  nand_x1_sg U39667 ( .A(n8412), .B(n47392), .X(n7852) );
  nand_x1_sg U39668 ( .A(n8917), .B(n8918), .X(n8889) );
  nand_x1_sg U39669 ( .A(n8919), .B(n41888), .X(n8918) );
  nand_x1_sg U39670 ( .A(n47510), .B(n8892), .X(n8886) );
  nand_x1_sg U39671 ( .A(n47520), .B(n8937), .X(n8932) );
  nand_x1_sg U39672 ( .A(n8933), .B(n47549), .X(n8908) );
  inv_x1_sg U39673 ( .A(n9024), .X(n47535) );
  nand_x1_sg U39674 ( .A(n8971), .B(n8972), .X(n8965) );
  nand_x1_sg U39675 ( .A(n8967), .B(n8968), .X(n8945) );
  inv_x1_sg U39676 ( .A(n8969), .X(n47544) );
  nand_x1_sg U39677 ( .A(n9014), .B(n47542), .X(n9010) );
  nand_x1_sg U39678 ( .A(n9011), .B(n9012), .X(n8969) );
  nand_x1_sg U39679 ( .A(n9030), .B(n9031), .X(n9024) );
  nand_x1_sg U39680 ( .A(n8996), .B(n8997), .X(n8998) );
  nand_x1_sg U39681 ( .A(n9064), .B(n9065), .X(n9058) );
  nand_x1_sg U39682 ( .A(n9056), .B(n47592), .X(n9036) );
  nand_x1_sg U39683 ( .A(n47608), .B(n9060), .X(n9037) );
  nand_x1_sg U39684 ( .A(n9098), .B(n47596), .X(n9061) );
  nand_x1_sg U39685 ( .A(n9106), .B(n47605), .X(n9104) );
  nand_x1_sg U39686 ( .A(n9114), .B(n47635), .X(n9113) );
  nand_x1_sg U39687 ( .A(n9135), .B(n9134), .X(n9121) );
  nand_x1_sg U39688 ( .A(n9123), .B(n9124), .X(n9084) );
  nand_x1_sg U39689 ( .A(n9100), .B(n9101), .X(n9123) );
  nand_x1_sg U39690 ( .A(n9121), .B(n47600), .X(n9085) );
  nand_x1_sg U39691 ( .A(n9193), .B(n9194), .X(n9191) );
  nand_x1_sg U39692 ( .A(n9199), .B(n47622), .X(n9192) );
  nand_x1_sg U39693 ( .A(n9156), .B(n9155), .X(n9157) );
  inv_x1_sg U39694 ( .A(n8671), .X(n47653) );
  nand_x1_sg U39695 ( .A(n9230), .B(n47677), .X(n8670) );
  nand_x1_sg U39696 ( .A(n9737), .B(n9738), .X(n9709) );
  nand_x1_sg U39697 ( .A(n9739), .B(n41878), .X(n9738) );
  nand_x1_sg U39698 ( .A(n47795), .B(n9712), .X(n9706) );
  nand_x1_sg U39699 ( .A(n47805), .B(n9757), .X(n9752) );
  nand_x1_sg U39700 ( .A(n9753), .B(n47834), .X(n9728) );
  inv_x1_sg U39701 ( .A(n9844), .X(n47820) );
  nand_x1_sg U39702 ( .A(n9791), .B(n9792), .X(n9785) );
  nand_x1_sg U39703 ( .A(n9787), .B(n9788), .X(n9765) );
  inv_x1_sg U39704 ( .A(n9789), .X(n47829) );
  nand_x1_sg U39705 ( .A(n9834), .B(n47827), .X(n9830) );
  nand_x1_sg U39706 ( .A(n9831), .B(n9832), .X(n9789) );
  nand_x1_sg U39707 ( .A(n9850), .B(n9851), .X(n9844) );
  nand_x1_sg U39708 ( .A(n9816), .B(n9817), .X(n9818) );
  nand_x1_sg U39709 ( .A(n9884), .B(n9885), .X(n9878) );
  nand_x1_sg U39710 ( .A(n9876), .B(n47877), .X(n9856) );
  nand_x1_sg U39711 ( .A(n47893), .B(n9880), .X(n9857) );
  nand_x1_sg U39712 ( .A(n9918), .B(n47881), .X(n9881) );
  nand_x1_sg U39713 ( .A(n9926), .B(n47890), .X(n9924) );
  nand_x1_sg U39714 ( .A(n9934), .B(n47920), .X(n9933) );
  nand_x1_sg U39715 ( .A(n9955), .B(n9954), .X(n9941) );
  nand_x1_sg U39716 ( .A(n9943), .B(n9944), .X(n9904) );
  nand_x1_sg U39717 ( .A(n9920), .B(n9921), .X(n9943) );
  nand_x1_sg U39718 ( .A(n9941), .B(n47885), .X(n9905) );
  nand_x1_sg U39719 ( .A(n10013), .B(n10014), .X(n10011) );
  nand_x1_sg U39720 ( .A(n10019), .B(n47907), .X(n10012) );
  nand_x1_sg U39721 ( .A(n9976), .B(n9975), .X(n9977) );
  inv_x1_sg U39722 ( .A(n9491), .X(n47938) );
  nand_x1_sg U39723 ( .A(n10050), .B(n47962), .X(n9490) );
  nand_x1_sg U39724 ( .A(n10556), .B(n10557), .X(n10528) );
  nand_x1_sg U39725 ( .A(n10558), .B(n41898), .X(n10557) );
  nand_x1_sg U39726 ( .A(n48080), .B(n10531), .X(n10525) );
  nand_x1_sg U39727 ( .A(n48090), .B(n10576), .X(n10571) );
  nand_x1_sg U39728 ( .A(n10572), .B(n48119), .X(n10547) );
  inv_x1_sg U39729 ( .A(n10663), .X(n48105) );
  nand_x1_sg U39730 ( .A(n10610), .B(n10611), .X(n10604) );
  nand_x1_sg U39731 ( .A(n10606), .B(n10607), .X(n10584) );
  inv_x1_sg U39732 ( .A(n10608), .X(n48114) );
  nand_x1_sg U39733 ( .A(n10653), .B(n48112), .X(n10649) );
  nand_x1_sg U39734 ( .A(n10650), .B(n10651), .X(n10608) );
  nand_x1_sg U39735 ( .A(n10669), .B(n10670), .X(n10663) );
  nand_x1_sg U39736 ( .A(n10635), .B(n10636), .X(n10637) );
  nand_x1_sg U39737 ( .A(n10703), .B(n10704), .X(n10697) );
  nand_x1_sg U39738 ( .A(n10695), .B(n48162), .X(n10675) );
  nand_x1_sg U39739 ( .A(n48178), .B(n10699), .X(n10676) );
  nand_x1_sg U39740 ( .A(n10737), .B(n48166), .X(n10700) );
  nand_x1_sg U39741 ( .A(n10745), .B(n48175), .X(n10743) );
  nand_x1_sg U39742 ( .A(n10753), .B(n48205), .X(n10752) );
  nand_x1_sg U39743 ( .A(n10774), .B(n10773), .X(n10760) );
  nand_x1_sg U39744 ( .A(n10762), .B(n10763), .X(n10723) );
  nand_x1_sg U39745 ( .A(n10739), .B(n10740), .X(n10762) );
  nand_x1_sg U39746 ( .A(n10760), .B(n48170), .X(n10724) );
  nand_x1_sg U39747 ( .A(n10832), .B(n10833), .X(n10830) );
  nand_x1_sg U39748 ( .A(n10838), .B(n48192), .X(n10831) );
  nand_x1_sg U39749 ( .A(n10795), .B(n10794), .X(n10796) );
  inv_x1_sg U39750 ( .A(n10310), .X(n48223) );
  nand_x1_sg U39751 ( .A(n10869), .B(n48247), .X(n10309) );
  nand_x1_sg U39752 ( .A(n11375), .B(n11376), .X(n11347) );
  nand_x1_sg U39753 ( .A(n11377), .B(n41886), .X(n11376) );
  nand_x1_sg U39754 ( .A(n48365), .B(n11350), .X(n11344) );
  nand_x1_sg U39755 ( .A(n48375), .B(n11395), .X(n11390) );
  nand_x1_sg U39756 ( .A(n11391), .B(n48404), .X(n11366) );
  inv_x1_sg U39757 ( .A(n11482), .X(n48390) );
  nand_x1_sg U39758 ( .A(n11429), .B(n11430), .X(n11423) );
  nand_x1_sg U39759 ( .A(n11425), .B(n11426), .X(n11403) );
  inv_x1_sg U39760 ( .A(n11427), .X(n48399) );
  nand_x1_sg U39761 ( .A(n11472), .B(n48397), .X(n11468) );
  nand_x1_sg U39762 ( .A(n11469), .B(n11470), .X(n11427) );
  nand_x1_sg U39763 ( .A(n11488), .B(n11489), .X(n11482) );
  nand_x1_sg U39764 ( .A(n11454), .B(n11455), .X(n11456) );
  nand_x1_sg U39765 ( .A(n11522), .B(n11523), .X(n11516) );
  nand_x1_sg U39766 ( .A(n11514), .B(n48447), .X(n11494) );
  nand_x1_sg U39767 ( .A(n48463), .B(n11518), .X(n11495) );
  nand_x1_sg U39768 ( .A(n11556), .B(n48451), .X(n11519) );
  nand_x1_sg U39769 ( .A(n11564), .B(n48460), .X(n11562) );
  nand_x1_sg U39770 ( .A(n11572), .B(n48490), .X(n11571) );
  nand_x1_sg U39771 ( .A(n11593), .B(n11592), .X(n11579) );
  nand_x1_sg U39772 ( .A(n11581), .B(n11582), .X(n11542) );
  nand_x1_sg U39773 ( .A(n11558), .B(n11559), .X(n11581) );
  nand_x1_sg U39774 ( .A(n11579), .B(n48455), .X(n11543) );
  nand_x1_sg U39775 ( .A(n11651), .B(n11652), .X(n11649) );
  nand_x1_sg U39776 ( .A(n11657), .B(n48477), .X(n11650) );
  nand_x1_sg U39777 ( .A(n11614), .B(n11613), .X(n11615) );
  inv_x1_sg U39778 ( .A(n11129), .X(n48508) );
  nand_x1_sg U39779 ( .A(n11688), .B(n48532), .X(n11128) );
  nand_x1_sg U39780 ( .A(n12194), .B(n12195), .X(n12166) );
  nand_x1_sg U39781 ( .A(n12196), .B(n41884), .X(n12195) );
  nand_x1_sg U39782 ( .A(n48650), .B(n12169), .X(n12163) );
  nand_x1_sg U39783 ( .A(n48660), .B(n12214), .X(n12209) );
  nand_x1_sg U39784 ( .A(n12210), .B(n48689), .X(n12185) );
  inv_x1_sg U39785 ( .A(n12301), .X(n48675) );
  nand_x1_sg U39786 ( .A(n12248), .B(n12249), .X(n12242) );
  nand_x1_sg U39787 ( .A(n12244), .B(n12245), .X(n12222) );
  inv_x1_sg U39788 ( .A(n12246), .X(n48684) );
  nand_x1_sg U39789 ( .A(n12291), .B(n48682), .X(n12287) );
  nand_x1_sg U39790 ( .A(n12288), .B(n12289), .X(n12246) );
  nand_x1_sg U39791 ( .A(n12307), .B(n12308), .X(n12301) );
  nand_x1_sg U39792 ( .A(n12273), .B(n12274), .X(n12275) );
  nand_x1_sg U39793 ( .A(n12341), .B(n12342), .X(n12335) );
  nand_x1_sg U39794 ( .A(n12333), .B(n48732), .X(n12313) );
  nand_x1_sg U39795 ( .A(n48748), .B(n12337), .X(n12314) );
  nand_x1_sg U39796 ( .A(n12375), .B(n48736), .X(n12338) );
  nand_x1_sg U39797 ( .A(n12383), .B(n48745), .X(n12381) );
  nand_x1_sg U39798 ( .A(n12391), .B(n48775), .X(n12390) );
  nand_x1_sg U39799 ( .A(n12412), .B(n12411), .X(n12398) );
  nand_x1_sg U39800 ( .A(n12400), .B(n12401), .X(n12361) );
  nand_x1_sg U39801 ( .A(n12377), .B(n12378), .X(n12400) );
  nand_x1_sg U39802 ( .A(n12398), .B(n48740), .X(n12362) );
  nand_x1_sg U39803 ( .A(n12470), .B(n12471), .X(n12468) );
  nand_x1_sg U39804 ( .A(n12476), .B(n48762), .X(n12469) );
  nand_x1_sg U39805 ( .A(n12433), .B(n12432), .X(n12434) );
  inv_x1_sg U39806 ( .A(n11948), .X(n48793) );
  nand_x1_sg U39807 ( .A(n12507), .B(n48817), .X(n11947) );
  nand_x1_sg U39808 ( .A(n13013), .B(n13014), .X(n12985) );
  nand_x1_sg U39809 ( .A(n13015), .B(n41896), .X(n13014) );
  nand_x1_sg U39810 ( .A(n48936), .B(n12988), .X(n12982) );
  nand_x1_sg U39811 ( .A(n48946), .B(n13033), .X(n13028) );
  nand_x1_sg U39812 ( .A(n13029), .B(n48975), .X(n13004) );
  inv_x1_sg U39813 ( .A(n13120), .X(n48961) );
  nand_x1_sg U39814 ( .A(n13067), .B(n13068), .X(n13061) );
  nand_x1_sg U39815 ( .A(n13063), .B(n13064), .X(n13041) );
  inv_x1_sg U39816 ( .A(n13065), .X(n48970) );
  nand_x1_sg U39817 ( .A(n13110), .B(n48968), .X(n13106) );
  nand_x1_sg U39818 ( .A(n13107), .B(n13108), .X(n13065) );
  nand_x1_sg U39819 ( .A(n13126), .B(n13127), .X(n13120) );
  nand_x1_sg U39820 ( .A(n13092), .B(n13093), .X(n13094) );
  nand_x1_sg U39821 ( .A(n13160), .B(n13161), .X(n13154) );
  nand_x1_sg U39822 ( .A(n13152), .B(n49018), .X(n13132) );
  nand_x1_sg U39823 ( .A(n49034), .B(n13156), .X(n13133) );
  nand_x1_sg U39824 ( .A(n13194), .B(n49022), .X(n13157) );
  nand_x1_sg U39825 ( .A(n13202), .B(n49031), .X(n13200) );
  nand_x1_sg U39826 ( .A(n13210), .B(n49062), .X(n13209) );
  nand_x1_sg U39827 ( .A(n13231), .B(n13230), .X(n13217) );
  nand_x1_sg U39828 ( .A(n13219), .B(n13220), .X(n13180) );
  nand_x1_sg U39829 ( .A(n13196), .B(n13197), .X(n13219) );
  nand_x1_sg U39830 ( .A(n13217), .B(n49026), .X(n13181) );
  nand_x1_sg U39831 ( .A(n13289), .B(n13290), .X(n13287) );
  nand_x1_sg U39832 ( .A(n13295), .B(n49048), .X(n13288) );
  nand_x1_sg U39833 ( .A(n13252), .B(n13251), .X(n13253) );
  inv_x1_sg U39834 ( .A(n12767), .X(n49080) );
  nand_x1_sg U39835 ( .A(n13326), .B(n49104), .X(n12766) );
  nand_x1_sg U39836 ( .A(n13832), .B(n13833), .X(n13804) );
  nand_x1_sg U39837 ( .A(n13834), .B(n41882), .X(n13833) );
  nand_x1_sg U39838 ( .A(n49223), .B(n13807), .X(n13801) );
  nand_x1_sg U39839 ( .A(n49233), .B(n13852), .X(n13847) );
  nand_x1_sg U39840 ( .A(n13848), .B(n49262), .X(n13823) );
  inv_x1_sg U39841 ( .A(n13939), .X(n49248) );
  nand_x1_sg U39842 ( .A(n13886), .B(n13887), .X(n13880) );
  nand_x1_sg U39843 ( .A(n13882), .B(n13883), .X(n13860) );
  inv_x1_sg U39844 ( .A(n13884), .X(n49257) );
  nand_x1_sg U39845 ( .A(n13929), .B(n49255), .X(n13925) );
  nand_x1_sg U39846 ( .A(n13926), .B(n13927), .X(n13884) );
  nand_x1_sg U39847 ( .A(n13945), .B(n13946), .X(n13939) );
  nand_x1_sg U39848 ( .A(n13911), .B(n13912), .X(n13913) );
  nand_x1_sg U39849 ( .A(n13979), .B(n13980), .X(n13973) );
  nand_x1_sg U39850 ( .A(n13971), .B(n49305), .X(n13951) );
  nand_x1_sg U39851 ( .A(n49321), .B(n13975), .X(n13952) );
  nand_x1_sg U39852 ( .A(n14013), .B(n49309), .X(n13976) );
  nand_x1_sg U39853 ( .A(n14021), .B(n49318), .X(n14019) );
  nand_x1_sg U39854 ( .A(n14029), .B(n49348), .X(n14028) );
  nand_x1_sg U39855 ( .A(n14050), .B(n14049), .X(n14036) );
  nand_x1_sg U39856 ( .A(n14038), .B(n14039), .X(n13999) );
  nand_x1_sg U39857 ( .A(n14015), .B(n14016), .X(n14038) );
  nand_x1_sg U39858 ( .A(n14036), .B(n49313), .X(n14000) );
  nand_x1_sg U39859 ( .A(n14108), .B(n14109), .X(n14106) );
  nand_x1_sg U39860 ( .A(n14114), .B(n49335), .X(n14107) );
  nand_x1_sg U39861 ( .A(n14071), .B(n14070), .X(n14072) );
  inv_x1_sg U39862 ( .A(n13586), .X(n49366) );
  nand_x1_sg U39863 ( .A(n14145), .B(n49390), .X(n13585) );
  nand_x1_sg U39864 ( .A(n14651), .B(n14652), .X(n14623) );
  nand_x1_sg U39865 ( .A(n14653), .B(n41880), .X(n14652) );
  nand_x1_sg U39866 ( .A(n49509), .B(n14626), .X(n14620) );
  nand_x1_sg U39867 ( .A(n49519), .B(n14671), .X(n14666) );
  nand_x1_sg U39868 ( .A(n14667), .B(n49548), .X(n14642) );
  inv_x1_sg U39869 ( .A(n14758), .X(n49534) );
  nand_x1_sg U39870 ( .A(n14705), .B(n14706), .X(n14699) );
  nand_x1_sg U39871 ( .A(n14701), .B(n14702), .X(n14679) );
  inv_x1_sg U39872 ( .A(n14703), .X(n49543) );
  nand_x1_sg U39873 ( .A(n14748), .B(n49541), .X(n14744) );
  nand_x1_sg U39874 ( .A(n14745), .B(n14746), .X(n14703) );
  nand_x1_sg U39875 ( .A(n14764), .B(n14765), .X(n14758) );
  nand_x1_sg U39876 ( .A(n14730), .B(n14731), .X(n14732) );
  nand_x1_sg U39877 ( .A(n14798), .B(n14799), .X(n14792) );
  nand_x1_sg U39878 ( .A(n14790), .B(n49591), .X(n14770) );
  nand_x1_sg U39879 ( .A(n49607), .B(n14794), .X(n14771) );
  nand_x1_sg U39880 ( .A(n14832), .B(n49595), .X(n14795) );
  nand_x1_sg U39881 ( .A(n14840), .B(n49604), .X(n14838) );
  nand_x1_sg U39882 ( .A(n14848), .B(n49634), .X(n14847) );
  nand_x1_sg U39883 ( .A(n14869), .B(n14868), .X(n14855) );
  nand_x1_sg U39884 ( .A(n14857), .B(n14858), .X(n14818) );
  nand_x1_sg U39885 ( .A(n14834), .B(n14835), .X(n14857) );
  nand_x1_sg U39886 ( .A(n14855), .B(n49599), .X(n14819) );
  nand_x1_sg U39887 ( .A(n14927), .B(n14928), .X(n14925) );
  nand_x1_sg U39888 ( .A(n14933), .B(n49621), .X(n14926) );
  nand_x1_sg U39889 ( .A(n14890), .B(n14889), .X(n14891) );
  inv_x1_sg U39890 ( .A(n14405), .X(n49652) );
  nand_x1_sg U39891 ( .A(n14964), .B(n49676), .X(n14404) );
  nand_x1_sg U39892 ( .A(n15470), .B(n15471), .X(n15442) );
  nand_x1_sg U39893 ( .A(n15472), .B(n41876), .X(n15471) );
  nand_x1_sg U39894 ( .A(n49795), .B(n15445), .X(n15439) );
  nand_x1_sg U39895 ( .A(n49805), .B(n15490), .X(n15485) );
  nand_x1_sg U39896 ( .A(n15486), .B(n49834), .X(n15461) );
  inv_x1_sg U39897 ( .A(n15577), .X(n49820) );
  nand_x1_sg U39898 ( .A(n15524), .B(n15525), .X(n15518) );
  nand_x1_sg U39899 ( .A(n15520), .B(n15521), .X(n15498) );
  inv_x1_sg U39900 ( .A(n15522), .X(n49829) );
  nand_x1_sg U39901 ( .A(n15567), .B(n49827), .X(n15563) );
  nand_x1_sg U39902 ( .A(n15564), .B(n15565), .X(n15522) );
  nand_x1_sg U39903 ( .A(n15583), .B(n15584), .X(n15577) );
  nand_x1_sg U39904 ( .A(n15549), .B(n15550), .X(n15551) );
  nand_x1_sg U39905 ( .A(n15617), .B(n15618), .X(n15611) );
  nand_x1_sg U39906 ( .A(n15609), .B(n49877), .X(n15589) );
  nand_x1_sg U39907 ( .A(n49893), .B(n15613), .X(n15590) );
  nand_x1_sg U39908 ( .A(n15651), .B(n49881), .X(n15614) );
  nand_x1_sg U39909 ( .A(n15659), .B(n49890), .X(n15657) );
  nand_x1_sg U39910 ( .A(n15667), .B(n49920), .X(n15666) );
  nand_x1_sg U39911 ( .A(n15688), .B(n15687), .X(n15674) );
  nand_x1_sg U39912 ( .A(n15676), .B(n15677), .X(n15637) );
  nand_x1_sg U39913 ( .A(n15653), .B(n15654), .X(n15676) );
  nand_x1_sg U39914 ( .A(n15674), .B(n49885), .X(n15638) );
  nand_x1_sg U39915 ( .A(n15746), .B(n15747), .X(n15744) );
  nand_x1_sg U39916 ( .A(n15752), .B(n49907), .X(n15745) );
  nand_x1_sg U39917 ( .A(n15709), .B(n15708), .X(n15710) );
  inv_x1_sg U39918 ( .A(n15224), .X(n49938) );
  nand_x1_sg U39919 ( .A(n15783), .B(n49962), .X(n15223) );
  nand_x1_sg U39920 ( .A(n16289), .B(n16290), .X(n16261) );
  nand_x1_sg U39921 ( .A(n16291), .B(n41894), .X(n16290) );
  nand_x1_sg U39922 ( .A(n50081), .B(n16264), .X(n16258) );
  nand_x1_sg U39923 ( .A(n50091), .B(n16309), .X(n16304) );
  nand_x1_sg U39924 ( .A(n16305), .B(n50120), .X(n16280) );
  inv_x1_sg U39925 ( .A(n16396), .X(n50106) );
  nand_x1_sg U39926 ( .A(n16343), .B(n16344), .X(n16337) );
  nand_x1_sg U39927 ( .A(n16339), .B(n16340), .X(n16317) );
  inv_x1_sg U39928 ( .A(n16341), .X(n50115) );
  nand_x1_sg U39929 ( .A(n16386), .B(n50113), .X(n16382) );
  nand_x1_sg U39930 ( .A(n16383), .B(n16384), .X(n16341) );
  nand_x1_sg U39931 ( .A(n16402), .B(n16403), .X(n16396) );
  nand_x1_sg U39932 ( .A(n16368), .B(n16369), .X(n16370) );
  nand_x1_sg U39933 ( .A(n16436), .B(n16437), .X(n16430) );
  nand_x1_sg U39934 ( .A(n16428), .B(n50163), .X(n16408) );
  nand_x1_sg U39935 ( .A(n50179), .B(n16432), .X(n16409) );
  nand_x1_sg U39936 ( .A(n16470), .B(n50167), .X(n16433) );
  nand_x1_sg U39937 ( .A(n16478), .B(n50176), .X(n16476) );
  nand_x1_sg U39938 ( .A(n16486), .B(n50206), .X(n16485) );
  nand_x1_sg U39939 ( .A(n16507), .B(n16506), .X(n16493) );
  nand_x1_sg U39940 ( .A(n16495), .B(n16496), .X(n16456) );
  nand_x1_sg U39941 ( .A(n16472), .B(n16473), .X(n16495) );
  nand_x1_sg U39942 ( .A(n16493), .B(n50171), .X(n16457) );
  nand_x1_sg U39943 ( .A(n16565), .B(n16566), .X(n16563) );
  nand_x1_sg U39944 ( .A(n16571), .B(n50193), .X(n16564) );
  nand_x1_sg U39945 ( .A(n16528), .B(n16527), .X(n16529) );
  inv_x1_sg U39946 ( .A(n16043), .X(n50224) );
  nand_x1_sg U39947 ( .A(n16602), .B(n50248), .X(n16042) );
  nand_x1_sg U39948 ( .A(n17105), .B(n17106), .X(n17077) );
  nand_x1_sg U39949 ( .A(n50366), .B(n17080), .X(n17074) );
  nand_x1_sg U39950 ( .A(n50376), .B(n17126), .X(n17121) );
  nand_x1_sg U39951 ( .A(n17122), .B(n50405), .X(n17096) );
  inv_x1_sg U39952 ( .A(n17213), .X(n50391) );
  nand_x1_sg U39953 ( .A(n17160), .B(n17161), .X(n17154) );
  nand_x1_sg U39954 ( .A(n17156), .B(n17157), .X(n17134) );
  inv_x1_sg U39955 ( .A(n17158), .X(n50400) );
  nand_x1_sg U39956 ( .A(n17203), .B(n50398), .X(n17199) );
  nand_x1_sg U39957 ( .A(n17200), .B(n17201), .X(n17158) );
  nand_x1_sg U39958 ( .A(n17219), .B(n17220), .X(n17213) );
  nand_x1_sg U39959 ( .A(n17185), .B(n17186), .X(n17187) );
  inv_x1_sg U39960 ( .A(n17225), .X(n50449) );
  nand_x1_sg U39961 ( .A(n17253), .B(n17254), .X(n17247) );
  nand_x1_sg U39962 ( .A(n50464), .B(n17249), .X(n17226) );
  nand_x1_sg U39963 ( .A(n17245), .B(n50448), .X(n17225) );
  nand_x1_sg U39964 ( .A(n17287), .B(n50452), .X(n17250) );
  nand_x1_sg U39965 ( .A(n17295), .B(n50461), .X(n17293) );
  nand_x1_sg U39966 ( .A(n17303), .B(n50491), .X(n17302) );
  nand_x1_sg U39967 ( .A(n17324), .B(n17323), .X(n17310) );
  nand_x1_sg U39968 ( .A(n17312), .B(n17313), .X(n17273) );
  nand_x1_sg U39969 ( .A(n17289), .B(n17290), .X(n17312) );
  nand_x1_sg U39970 ( .A(n17310), .B(n50456), .X(n17274) );
  nand_x1_sg U39971 ( .A(n17382), .B(n17383), .X(n17380) );
  nand_x1_sg U39972 ( .A(n17388), .B(n50478), .X(n17381) );
  nand_x1_sg U39973 ( .A(n17345), .B(n17344), .X(n17346) );
  inv_x1_sg U39974 ( .A(n16862), .X(n50509) );
  nand_x1_sg U39975 ( .A(n17419), .B(n50533), .X(n16861) );
  nand_x1_sg U39976 ( .A(n17927), .B(n17928), .X(n17899) );
  nand_x1_sg U39977 ( .A(n17929), .B(n41890), .X(n17928) );
  nand_x1_sg U39978 ( .A(n50655), .B(n17902), .X(n17896) );
  nand_x1_sg U39979 ( .A(n50665), .B(n17947), .X(n17942) );
  nand_x1_sg U39980 ( .A(n17943), .B(n50694), .X(n17918) );
  inv_x1_sg U39981 ( .A(n18034), .X(n50680) );
  nand_x1_sg U39982 ( .A(n17981), .B(n17982), .X(n17975) );
  nand_x1_sg U39983 ( .A(n17977), .B(n17978), .X(n17955) );
  inv_x1_sg U39984 ( .A(n17979), .X(n50689) );
  nand_x1_sg U39985 ( .A(n18024), .B(n50687), .X(n18020) );
  nand_x1_sg U39986 ( .A(n18021), .B(n18022), .X(n17979) );
  nand_x1_sg U39987 ( .A(n18040), .B(n18041), .X(n18034) );
  nand_x1_sg U39988 ( .A(n18006), .B(n18007), .X(n18008) );
  nand_x1_sg U39989 ( .A(n18074), .B(n18075), .X(n18068) );
  nand_x1_sg U39990 ( .A(n18066), .B(n50737), .X(n18046) );
  nand_x1_sg U39991 ( .A(n50753), .B(n18070), .X(n18047) );
  nand_x1_sg U39992 ( .A(n18108), .B(n50741), .X(n18071) );
  nand_x1_sg U39993 ( .A(n18116), .B(n50750), .X(n18114) );
  nand_x1_sg U39994 ( .A(n18124), .B(n50780), .X(n18123) );
  nand_x1_sg U39995 ( .A(n18145), .B(n18144), .X(n18131) );
  nand_x1_sg U39996 ( .A(n18133), .B(n18134), .X(n18094) );
  nand_x1_sg U39997 ( .A(n18110), .B(n18111), .X(n18133) );
  nand_x1_sg U39998 ( .A(n18131), .B(n50745), .X(n18095) );
  nand_x1_sg U39999 ( .A(n18203), .B(n18204), .X(n18201) );
  nand_x1_sg U40000 ( .A(n18209), .B(n50767), .X(n18202) );
  nand_x1_sg U40001 ( .A(n18166), .B(n18165), .X(n18167) );
  inv_x1_sg U40002 ( .A(n17681), .X(n50798) );
  nand_x1_sg U40003 ( .A(n18240), .B(n50822), .X(n17680) );
  nand_x1_sg U40004 ( .A(n18748), .B(n18749), .X(n18720) );
  nand_x1_sg U40005 ( .A(n18750), .B(n41892), .X(n18749) );
  nand_x1_sg U40006 ( .A(n50942), .B(n18723), .X(n18717) );
  nand_x1_sg U40007 ( .A(n50952), .B(n18768), .X(n18763) );
  nand_x1_sg U40008 ( .A(n18764), .B(n50981), .X(n18739) );
  inv_x1_sg U40009 ( .A(n18855), .X(n50967) );
  nand_x1_sg U40010 ( .A(n18802), .B(n18803), .X(n18796) );
  nand_x1_sg U40011 ( .A(n18798), .B(n18799), .X(n18776) );
  inv_x1_sg U40012 ( .A(n18800), .X(n50976) );
  nand_x1_sg U40013 ( .A(n18845), .B(n50974), .X(n18841) );
  nand_x1_sg U40014 ( .A(n18842), .B(n18843), .X(n18800) );
  nand_x1_sg U40015 ( .A(n18861), .B(n18862), .X(n18855) );
  nand_x1_sg U40016 ( .A(n18827), .B(n18828), .X(n18829) );
  nand_x1_sg U40017 ( .A(n18895), .B(n18896), .X(n18889) );
  nand_x1_sg U40018 ( .A(n18887), .B(n51024), .X(n18867) );
  nand_x1_sg U40019 ( .A(n51040), .B(n18891), .X(n18868) );
  nand_x1_sg U40020 ( .A(n18929), .B(n51028), .X(n18892) );
  nand_x1_sg U40021 ( .A(n18937), .B(n51037), .X(n18935) );
  nand_x1_sg U40022 ( .A(n18945), .B(n51067), .X(n18944) );
  nand_x1_sg U40023 ( .A(n18966), .B(n18965), .X(n18952) );
  nand_x1_sg U40024 ( .A(n18954), .B(n18955), .X(n18915) );
  nand_x1_sg U40025 ( .A(n18931), .B(n18932), .X(n18954) );
  nand_x1_sg U40026 ( .A(n18952), .B(n51032), .X(n18916) );
  nand_x1_sg U40027 ( .A(n19024), .B(n19025), .X(n19022) );
  nand_x1_sg U40028 ( .A(n19030), .B(n51054), .X(n19023) );
  nand_x1_sg U40029 ( .A(n18987), .B(n18986), .X(n18988) );
  inv_x1_sg U40030 ( .A(n18502), .X(n51085) );
  nand_x1_sg U40031 ( .A(n19061), .B(n51109), .X(n18501) );
  inv_x1_sg U40032 ( .A(n26843), .X(n45733) );
  nand_x1_sg U40033 ( .A(n27096), .B(n27097), .X(n26843) );
  inv_x1_sg U40034 ( .A(n26858), .X(n45732) );
  nand_x1_sg U40035 ( .A(n27109), .B(n27110), .X(n26858) );
  inv_x1_sg U40036 ( .A(n26879), .X(n45729) );
  nand_x1_sg U40037 ( .A(n27127), .B(n27128), .X(n26879) );
  inv_x1_sg U40038 ( .A(n26872), .X(n45730) );
  nand_x1_sg U40039 ( .A(n27121), .B(n27122), .X(n26872) );
  inv_x1_sg U40040 ( .A(n26865), .X(n45731) );
  nand_x1_sg U40041 ( .A(n27115), .B(n27116), .X(n26865) );
  inv_x1_sg U40042 ( .A(n26886), .X(n45728) );
  nand_x1_sg U40043 ( .A(n27133), .B(n27134), .X(n26886) );
  inv_x1_sg U40044 ( .A(n27099), .X(n45690) );
  nand_x1_sg U40045 ( .A(n27326), .B(n27327), .X(n27099) );
  inv_x1_sg U40046 ( .A(n27112), .X(n45689) );
  nand_x1_sg U40047 ( .A(n27339), .B(n27340), .X(n27112) );
  inv_x1_sg U40048 ( .A(n27130), .X(n45686) );
  nand_x1_sg U40049 ( .A(n27357), .B(n27358), .X(n27130) );
  inv_x1_sg U40050 ( .A(n27124), .X(n45687) );
  nand_x1_sg U40051 ( .A(n27351), .B(n27352), .X(n27124) );
  inv_x1_sg U40052 ( .A(n27118), .X(n45688) );
  nand_x1_sg U40053 ( .A(n27345), .B(n27346), .X(n27118) );
  inv_x1_sg U40054 ( .A(n27136), .X(n45685) );
  nand_x1_sg U40055 ( .A(n27363), .B(n27364), .X(n27136) );
  inv_x1_sg U40056 ( .A(n27329), .X(n45646) );
  nand_x1_sg U40057 ( .A(n27539), .B(n27540), .X(n27329) );
  inv_x1_sg U40058 ( .A(n27342), .X(n45645) );
  nand_x1_sg U40059 ( .A(n27552), .B(n27553), .X(n27342) );
  inv_x1_sg U40060 ( .A(n27360), .X(n45642) );
  nand_x1_sg U40061 ( .A(n27570), .B(n27571), .X(n27360) );
  inv_x1_sg U40062 ( .A(n27354), .X(n45643) );
  nand_x1_sg U40063 ( .A(n27564), .B(n27565), .X(n27354) );
  inv_x1_sg U40064 ( .A(n27348), .X(n45644) );
  nand_x1_sg U40065 ( .A(n27558), .B(n27559), .X(n27348) );
  inv_x1_sg U40066 ( .A(n27287), .X(n45641) );
  nand_x1_sg U40067 ( .A(n27366), .B(n27367), .X(n27287) );
  inv_x1_sg U40068 ( .A(n27542), .X(n45602) );
  nand_x1_sg U40069 ( .A(n27733), .B(n27734), .X(n27542) );
  inv_x1_sg U40070 ( .A(n27555), .X(n45601) );
  nand_x1_sg U40071 ( .A(n27746), .B(n27747), .X(n27555) );
  inv_x1_sg U40072 ( .A(n27503), .X(n45598) );
  nand_x1_sg U40073 ( .A(n27573), .B(n27574), .X(n27503) );
  inv_x1_sg U40074 ( .A(n27567), .X(n45599) );
  nand_x1_sg U40075 ( .A(n27758), .B(n27759), .X(n27567) );
  inv_x1_sg U40076 ( .A(n27561), .X(n45600) );
  nand_x1_sg U40077 ( .A(n27752), .B(n27753), .X(n27561) );
  inv_x1_sg U40078 ( .A(n27281), .X(n45597) );
  nand_x1_sg U40079 ( .A(n27369), .B(n27370), .X(n27281) );
  inv_x1_sg U40080 ( .A(n27736), .X(n45557) );
  nand_x1_sg U40081 ( .A(n27910), .B(n27911), .X(n27736) );
  inv_x1_sg U40082 ( .A(n27749), .X(n45556) );
  nand_x1_sg U40083 ( .A(n27923), .B(n27924), .X(n27749) );
  inv_x1_sg U40084 ( .A(n27497), .X(n45553) );
  nand_x1_sg U40085 ( .A(n27576), .B(n27577), .X(n27497) );
  inv_x1_sg U40086 ( .A(n27700), .X(n45554) );
  nand_x1_sg U40087 ( .A(n27761), .B(n27762), .X(n27700) );
  inv_x1_sg U40088 ( .A(n27755), .X(n45555) );
  nand_x1_sg U40089 ( .A(n27929), .B(n27930), .X(n27755) );
  inv_x1_sg U40090 ( .A(n27275), .X(n45552) );
  nand_x1_sg U40091 ( .A(n27372), .B(n27373), .X(n27275) );
  inv_x1_sg U40092 ( .A(n27913), .X(n45513) );
  nand_x1_sg U40093 ( .A(n28072), .B(n28073), .X(n27913) );
  inv_x1_sg U40094 ( .A(n27694), .X(n45510) );
  nand_x1_sg U40095 ( .A(n27764), .B(n27765), .X(n27694) );
  inv_x1_sg U40096 ( .A(n27926), .X(n45512) );
  nand_x1_sg U40097 ( .A(n28085), .B(n28086), .X(n27926) );
  inv_x1_sg U40098 ( .A(n27491), .X(n45509) );
  nand_x1_sg U40099 ( .A(n27579), .B(n27580), .X(n27491) );
  inv_x1_sg U40100 ( .A(n27880), .X(n45511) );
  nand_x1_sg U40101 ( .A(n27932), .B(n27933), .X(n27880) );
  inv_x1_sg U40102 ( .A(n27269), .X(n45508) );
  nand_x1_sg U40103 ( .A(n27375), .B(n27376), .X(n27269) );
  inv_x1_sg U40104 ( .A(n28075), .X(n45468) );
  nand_x1_sg U40105 ( .A(n28207), .B(n28208), .X(n28075) );
  inv_x1_sg U40106 ( .A(n28045), .X(n45464) );
  nand_x1_sg U40107 ( .A(n28088), .B(n28089), .X(n28045) );
  inv_x1_sg U40108 ( .A(n27485), .X(n45461) );
  nand_x1_sg U40109 ( .A(n27582), .B(n27583), .X(n27485) );
  inv_x1_sg U40110 ( .A(n27688), .X(n45462) );
  nand_x1_sg U40111 ( .A(n27767), .B(n27768), .X(n27688) );
  inv_x1_sg U40112 ( .A(n27874), .X(n45463) );
  nand_x1_sg U40113 ( .A(n27935), .B(n27936), .X(n27874) );
  inv_x1_sg U40114 ( .A(n27263), .X(n45460) );
  nand_x1_sg U40115 ( .A(n27378), .B(n27379), .X(n27263) );
  inv_x1_sg U40116 ( .A(n28210), .X(n45424) );
  nand_x1_sg U40117 ( .A(n28336), .B(n28337), .X(n28210) );
  inv_x1_sg U40118 ( .A(n28039), .X(n45420) );
  nand_x1_sg U40119 ( .A(n28091), .B(n28092), .X(n28039) );
  inv_x1_sg U40120 ( .A(n27479), .X(n45417) );
  nand_x1_sg U40121 ( .A(n27585), .B(n27586), .X(n27479) );
  inv_x1_sg U40122 ( .A(n27682), .X(n45418) );
  nand_x1_sg U40123 ( .A(n27770), .B(n27771), .X(n27682) );
  inv_x1_sg U40124 ( .A(n27868), .X(n45419) );
  nand_x1_sg U40125 ( .A(n27938), .B(n27939), .X(n27868) );
  inv_x1_sg U40126 ( .A(n27257), .X(n45416) );
  nand_x1_sg U40127 ( .A(n27381), .B(n27382), .X(n27257) );
  inv_x1_sg U40128 ( .A(n27676), .X(n45372) );
  nand_x1_sg U40129 ( .A(n27773), .B(n27774), .X(n27676) );
  inv_x1_sg U40130 ( .A(n28033), .X(n45374) );
  nand_x1_sg U40131 ( .A(n28094), .B(n28095), .X(n28033) );
  inv_x1_sg U40132 ( .A(n27473), .X(n45371) );
  nand_x1_sg U40133 ( .A(n27588), .B(n27589), .X(n27473) );
  inv_x1_sg U40134 ( .A(n27862), .X(n45373) );
  nand_x1_sg U40135 ( .A(n27941), .B(n27942), .X(n27862) );
  inv_x1_sg U40136 ( .A(n27251), .X(n45370) );
  nand_x1_sg U40137 ( .A(n27384), .B(n27385), .X(n27251) );
  inv_x1_sg U40138 ( .A(n27670), .X(n45327) );
  nand_x1_sg U40139 ( .A(n27776), .B(n27777), .X(n27670) );
  inv_x1_sg U40140 ( .A(n28027), .X(n45329) );
  nand_x1_sg U40141 ( .A(n28097), .B(n28098), .X(n28027) );
  inv_x1_sg U40142 ( .A(n27467), .X(n45326) );
  nand_x1_sg U40143 ( .A(n27591), .B(n27592), .X(n27467) );
  inv_x1_sg U40144 ( .A(n27856), .X(n45328) );
  nand_x1_sg U40145 ( .A(n27944), .B(n27945), .X(n27856) );
  inv_x1_sg U40146 ( .A(n27245), .X(n45325) );
  nand_x1_sg U40147 ( .A(n27387), .B(n27388), .X(n27245) );
  inv_x1_sg U40148 ( .A(n27664), .X(n45282) );
  nand_x1_sg U40149 ( .A(n27779), .B(n27780), .X(n27664) );
  inv_x1_sg U40150 ( .A(n28021), .X(n45284) );
  nand_x1_sg U40151 ( .A(n28100), .B(n28101), .X(n28021) );
  inv_x1_sg U40152 ( .A(n27461), .X(n45281) );
  nand_x1_sg U40153 ( .A(n27594), .B(n27595), .X(n27461) );
  inv_x1_sg U40154 ( .A(n27850), .X(n45283) );
  nand_x1_sg U40155 ( .A(n27947), .B(n27948), .X(n27850) );
  inv_x1_sg U40156 ( .A(n27239), .X(n45280) );
  nand_x1_sg U40157 ( .A(n27390), .B(n27391), .X(n27239) );
  inv_x1_sg U40158 ( .A(n28015), .X(n45239) );
  nand_x1_sg U40159 ( .A(n28103), .B(n28104), .X(n28015) );
  inv_x1_sg U40160 ( .A(n27455), .X(n45236) );
  nand_x1_sg U40161 ( .A(n27597), .B(n27598), .X(n27455) );
  inv_x1_sg U40162 ( .A(n27658), .X(n45237) );
  nand_x1_sg U40163 ( .A(n27782), .B(n27783), .X(n27658) );
  inv_x1_sg U40164 ( .A(n27844), .X(n45238) );
  nand_x1_sg U40165 ( .A(n27950), .B(n27951), .X(n27844) );
  inv_x1_sg U40166 ( .A(n27233), .X(n45235) );
  nand_x1_sg U40167 ( .A(n27393), .B(n27394), .X(n27233) );
  inv_x1_sg U40168 ( .A(n27652), .X(n45191) );
  nand_x1_sg U40169 ( .A(n27785), .B(n27786), .X(n27652) );
  inv_x1_sg U40170 ( .A(n28009), .X(n45193) );
  nand_x1_sg U40171 ( .A(n28106), .B(n28107), .X(n28009) );
  inv_x1_sg U40172 ( .A(n27449), .X(n45190) );
  nand_x1_sg U40173 ( .A(n27600), .B(n27601), .X(n27449) );
  inv_x1_sg U40174 ( .A(n27838), .X(n45192) );
  nand_x1_sg U40175 ( .A(n27953), .B(n27954), .X(n27838) );
  inv_x1_sg U40176 ( .A(n27227), .X(n45189) );
  nand_x1_sg U40177 ( .A(n27396), .B(n27397), .X(n27227) );
  inv_x1_sg U40178 ( .A(n27646), .X(n45146) );
  nand_x1_sg U40179 ( .A(n27788), .B(n27789), .X(n27646) );
  inv_x1_sg U40180 ( .A(n28003), .X(n45148) );
  nand_x1_sg U40181 ( .A(n28109), .B(n28110), .X(n28003) );
  inv_x1_sg U40182 ( .A(n27443), .X(n45145) );
  nand_x1_sg U40183 ( .A(n27603), .B(n27604), .X(n27443) );
  inv_x1_sg U40184 ( .A(n27832), .X(n45147) );
  nand_x1_sg U40185 ( .A(n27956), .B(n27957), .X(n27832) );
  inv_x1_sg U40186 ( .A(n27221), .X(n45144) );
  nand_x1_sg U40187 ( .A(n27399), .B(n27400), .X(n27221) );
  inv_x1_sg U40188 ( .A(n27997), .X(n45101) );
  nand_x1_sg U40189 ( .A(n28112), .B(n28113), .X(n27997) );
  inv_x1_sg U40190 ( .A(n27437), .X(n45098) );
  nand_x1_sg U40191 ( .A(n27606), .B(n27607), .X(n27437) );
  inv_x1_sg U40192 ( .A(n27640), .X(n45099) );
  nand_x1_sg U40193 ( .A(n27791), .B(n27792), .X(n27640) );
  inv_x1_sg U40194 ( .A(n27826), .X(n45100) );
  nand_x1_sg U40195 ( .A(n27959), .B(n27960), .X(n27826) );
  inv_x1_sg U40196 ( .A(n27215), .X(n45097) );
  nand_x1_sg U40197 ( .A(n27402), .B(n27403), .X(n27215) );
  inv_x1_sg U40198 ( .A(n27634), .X(n45055) );
  nand_x1_sg U40199 ( .A(n27794), .B(n27795), .X(n27634) );
  inv_x1_sg U40200 ( .A(n27991), .X(n45057) );
  nand_x1_sg U40201 ( .A(n28115), .B(n28116), .X(n27991) );
  inv_x1_sg U40202 ( .A(n27431), .X(n45054) );
  nand_x1_sg U40203 ( .A(n27609), .B(n27610), .X(n27431) );
  inv_x1_sg U40204 ( .A(n27820), .X(n45056) );
  nand_x1_sg U40205 ( .A(n27962), .B(n27963), .X(n27820) );
  inv_x1_sg U40206 ( .A(n27209), .X(n45053) );
  nand_x1_sg U40207 ( .A(n27405), .B(n27406), .X(n27209) );
  nand_x1_sg U40208 ( .A(n46925), .B(n46903), .X(n22780) );
  nand_x1_sg U40209 ( .A(n5474), .B(n19559), .X(n19558) );
  nand_x1_sg U40210 ( .A(n5512), .B(n19545), .X(n19544) );
  nand_x1_sg U40211 ( .A(n5493), .B(n19552), .X(n19551) );
  nand_x1_sg U40212 ( .A(n5550), .B(n19531), .X(n19530) );
  nand_x1_sg U40213 ( .A(n5664), .B(n20987), .X(n20986) );
  nand_x1_sg U40214 ( .A(n21183), .B(n21184), .X(n20982) );
  nand_x1_sg U40215 ( .A(out_L2[17]), .B(n21185), .X(n21184) );
  nand_x1_sg U40216 ( .A(n5685), .B(n46543), .X(n21185) );
  inv_x1_sg U40217 ( .A(n5995), .X(n46585) );
  nand_x1_sg U40218 ( .A(n19157), .B(n19158), .X(n6034) );
  inv_x1_sg U40219 ( .A(n6043), .X(n46545) );
  nand_x1_sg U40220 ( .A(n20793), .B(n20794), .X(n20777) );
  inv_x1_sg U40221 ( .A(n6084), .X(n46480) );
  nand_x1_sg U40222 ( .A(n19160), .B(n19161), .X(n6084) );
  inv_x1_sg U40223 ( .A(n6093), .X(n46503) );
  nand_x1_sg U40224 ( .A(n21159), .B(n46505), .X(n20947) );
  nand_x1_sg U40225 ( .A(n46477), .B(n20117), .X(n19912) );
  inv_x1_sg U40226 ( .A(n19713), .X(n46444) );
  nand_x1_sg U40227 ( .A(n21676), .B(n21677), .X(n21538) );
  nand_x1_sg U40228 ( .A(out_L2[14]), .B(n46368), .X(n21677) );
  inv_x1_sg U40229 ( .A(n21528), .X(n46462) );
  nand_x1_sg U40230 ( .A(n21546), .B(n21547), .X(n21528) );
  nand_x1_sg U40231 ( .A(n21153), .B(n46468), .X(n20940) );
  nand_x1_sg U40232 ( .A(n20938), .B(n20939), .X(n20761) );
  inv_x1_sg U40233 ( .A(n20941), .X(n46456) );
  nand_x1_sg U40234 ( .A(n19166), .B(n19167), .X(n6175) );
  inv_x1_sg U40235 ( .A(n19707), .X(n46395) );
  inv_x1_sg U40236 ( .A(n20440), .X(n46379) );
  inv_x1_sg U40237 ( .A(n21521), .X(n46414) );
  nand_x1_sg U40238 ( .A(n21549), .B(n21550), .X(n21521) );
  nand_x1_sg U40239 ( .A(n21147), .B(n46421), .X(n20933) );
  nand_x1_sg U40240 ( .A(n20931), .B(n20932), .X(n20754) );
  inv_x1_sg U40241 ( .A(n20934), .X(n46408) );
  inv_x1_sg U40242 ( .A(n19305), .X(n46343) );
  inv_x1_sg U40243 ( .A(n21515), .X(n46367) );
  nand_x1_sg U40244 ( .A(n21552), .B(n21553), .X(n21515) );
  nand_x1_sg U40245 ( .A(n21682), .B(n21683), .X(n21663) );
  nand_x1_sg U40246 ( .A(out_L2[12]), .B(n21684), .X(n21683) );
  nand_x1_sg U40247 ( .A(n5690), .B(n46281), .X(n21684) );
  nand_x1_sg U40248 ( .A(n20924), .B(n20925), .X(n20747) );
  inv_x1_sg U40249 ( .A(n20927), .X(n46361) );
  nand_x1_sg U40250 ( .A(n20426), .B(n46335), .X(n20276) );
  nand_x1_sg U40251 ( .A(n19693), .B(n46338), .X(n19470) );
  nor_x4_sg U40252 ( .A(n42112), .B(out_L2[12]), .X(n21660) );
  inv_x1_sg U40253 ( .A(n21508), .X(n46325) );
  nand_x1_sg U40254 ( .A(n21555), .B(n21556), .X(n21508) );
  nand_x1_sg U40255 ( .A(n20917), .B(n20918), .X(n20740) );
  inv_x1_sg U40256 ( .A(n20920), .X(n46319) );
  nand_x1_sg U40257 ( .A(n21688), .B(n21689), .X(n21651) );
  nand_x1_sg U40258 ( .A(out_L2[10]), .B(n21690), .X(n21689) );
  nand_x1_sg U40259 ( .A(n5692), .B(n46190), .X(n21690) );
  inv_x1_sg U40260 ( .A(n21502), .X(n46280) );
  nand_x1_sg U40261 ( .A(n21558), .B(n21559), .X(n21502) );
  nand_x1_sg U40262 ( .A(n21129), .B(n46286), .X(n20912) );
  nand_x1_sg U40263 ( .A(n20267), .B(n20268), .X(n20093) );
  inv_x1_sg U40264 ( .A(n20270), .X(n46265) );
  nand_x1_sg U40265 ( .A(n19687), .B(n46292), .X(n19463) );
  inv_x1_sg U40266 ( .A(n21495), .X(n46234) );
  nand_x1_sg U40267 ( .A(n21561), .B(n21562), .X(n21495) );
  nor_x4_sg U40268 ( .A(n42111), .B(out_L2[10]), .X(n21648) );
  nand_x1_sg U40269 ( .A(n21123), .B(n46241), .X(n20905) );
  nand_x1_sg U40270 ( .A(n20414), .B(n46244), .X(n20262) );
  nand_x1_sg U40271 ( .A(n19681), .B(n46247), .X(n19456) );
  nand_x1_sg U40272 ( .A(n21694), .B(n21695), .X(n21639) );
  nand_x1_sg U40273 ( .A(out_L2[8]), .B(n21696), .X(n21695) );
  nand_x1_sg U40274 ( .A(n5694), .B(n46099), .X(n21696) );
  inv_x1_sg U40275 ( .A(n21489), .X(n46189) );
  nand_x1_sg U40276 ( .A(n21564), .B(n21565), .X(n21489) );
  nand_x1_sg U40277 ( .A(n21117), .B(n46195), .X(n20898) );
  nand_x1_sg U40278 ( .A(n20408), .B(n46198), .X(n20255) );
  nand_x1_sg U40279 ( .A(n19675), .B(n46201), .X(n19449) );
  nand_x1_sg U40280 ( .A(n20246), .B(n20247), .X(n20072) );
  inv_x1_sg U40281 ( .A(n20249), .X(n46128) );
  nand_x1_sg U40282 ( .A(n19669), .B(n46156), .X(n19442) );
  nor_x4_sg U40283 ( .A(n42110), .B(out_L2[8]), .X(n21636) );
  inv_x1_sg U40284 ( .A(n21482), .X(n46143) );
  nand_x1_sg U40285 ( .A(n21567), .B(n21568), .X(n21482) );
  nand_x1_sg U40286 ( .A(n21111), .B(n46150), .X(n20891) );
  nand_x1_sg U40287 ( .A(n20396), .B(n46107), .X(n20241) );
  nand_x1_sg U40288 ( .A(n19663), .B(n46110), .X(n19435) );
  nand_x1_sg U40289 ( .A(n21700), .B(n21701), .X(n21627) );
  nand_x1_sg U40290 ( .A(out_L2[6]), .B(n21702), .X(n21701) );
  nand_x1_sg U40291 ( .A(n5696), .B(n46008), .X(n21702) );
  inv_x1_sg U40292 ( .A(n21476), .X(n46098) );
  nand_x1_sg U40293 ( .A(n21570), .B(n21571), .X(n21476) );
  nand_x1_sg U40294 ( .A(n21105), .B(n46104), .X(n20884) );
  nand_x1_sg U40295 ( .A(n20390), .B(n46062), .X(n20234) );
  nand_x1_sg U40296 ( .A(n19657), .B(n46065), .X(n19428) );
  nor_x4_sg U40297 ( .A(n42109), .B(out_L2[6]), .X(n21624) );
  inv_x1_sg U40298 ( .A(n21469), .X(n46052) );
  nand_x1_sg U40299 ( .A(n21573), .B(n21574), .X(n21469) );
  nand_x1_sg U40300 ( .A(n20875), .B(n20876), .X(n20698) );
  inv_x1_sg U40301 ( .A(n20878), .X(n46046) );
  nand_x1_sg U40302 ( .A(n20384), .B(n46016), .X(n20227) );
  nand_x1_sg U40303 ( .A(n19651), .B(n46019), .X(n19421) );
  nand_x2_sg U40304 ( .A(n21610), .B(n42108), .X(n21706) );
  inv_x1_sg U40305 ( .A(n21463), .X(n46007) );
  nand_x1_sg U40306 ( .A(n21576), .B(n21577), .X(n21463) );
  nand_x1_sg U40307 ( .A(n21093), .B(n46013), .X(n20870) );
  nand_x1_sg U40308 ( .A(n20378), .B(n45971), .X(n20220) );
  nand_x1_sg U40309 ( .A(n19645), .B(n45974), .X(n19414) );
  inv_x1_sg U40310 ( .A(n21456), .X(n45962) );
  nand_x1_sg U40311 ( .A(n21579), .B(n21580), .X(n21456) );
  nand_x1_sg U40312 ( .A(n21087), .B(n45968), .X(n20863) );
  inv_x1_sg U40313 ( .A(n21450), .X(n45916) );
  nand_x1_sg U40314 ( .A(n21582), .B(n21583), .X(n21450) );
  nand_x1_sg U40315 ( .A(n45880), .B(n20027), .X(n19841) );
  inv_x1_sg U40316 ( .A(n19842), .X(n45851) );
  inv_x1_sg U40317 ( .A(n20209), .X(n45843) );
  nand_x1_sg U40318 ( .A(n19211), .B(n19212), .X(n6715) );
  inv_x1_sg U40319 ( .A(n19403), .X(n45859) );
  nand_x1_sg U40320 ( .A(n45882), .B(n19633), .X(n19402) );
  nor_x4_sg U40321 ( .A(n42107), .B(out_L2[2]), .X(n21600) );
  nand_x1_sg U40322 ( .A(n21438), .B(n45874), .X(n21267) );
  nand_x1_sg U40323 ( .A(n45876), .B(n21075), .X(n20851) );
  inv_x1_sg U40324 ( .A(n20852), .X(n45827) );
  nand_x1_sg U40325 ( .A(n45877), .B(n20667), .X(n20498) );
  nand_x1_sg U40326 ( .A(n46874), .B(n7130), .X(n7126) );
  nand_x1_sg U40327 ( .A(n7138), .B(n7137), .X(n7139) );
  nand_x1_sg U40328 ( .A(n7182), .B(n7183), .X(n7165) );
  nand_x1_sg U40329 ( .A(n7204), .B(n7205), .X(n7191) );
  inv_x1_sg U40330 ( .A(n7207), .X(n46889) );
  nand_x1_sg U40331 ( .A(n46888), .B(n7224), .X(n7207) );
  nand_x1_sg U40332 ( .A(n7229), .B(n7230), .X(n7227) );
  nand_x1_sg U40333 ( .A(n46919), .B(n7286), .X(n7275) );
  nand_x1_sg U40334 ( .A(n7244), .B(n7245), .X(n7243) );
  nand_x2_sg U40335 ( .A(n7293), .B(n7294), .X(n7291) );
  inv_x1_sg U40336 ( .A(n7358), .X(n46970) );
  nand_x1_sg U40337 ( .A(n7372), .B(n7373), .X(n7358) );
  nand_x1_sg U40338 ( .A(n7320), .B(n7321), .X(n7322) );
  nand_x1_sg U40339 ( .A(n7398), .B(n7399), .X(n7384) );
  nand_x1_sg U40340 ( .A(n7401), .B(n47020), .X(n7398) );
  nand_x2_sg U40341 ( .A(n7460), .B(n7461), .X(n7416) );
  nand_x1_sg U40342 ( .A(n7417), .B(n7416), .X(n7414) );
  nand_x1_sg U40343 ( .A(n7524), .B(n7523), .X(n7516) );
  nand_x1_sg U40344 ( .A(n7516), .B(n47085), .X(n7511) );
  nand_x1_sg U40345 ( .A(n7544), .B(n7543), .X(n7041) );
  nand_x1_sg U40346 ( .A(n7590), .B(n7591), .X(n6961) );
  nand_x1_sg U40347 ( .A(n7579), .B(n7578), .X(n6947) );
  nand_x1_sg U40348 ( .A(n7574), .B(n7575), .X(n6950) );
  nand_x1_sg U40349 ( .A(n7634), .B(n47094), .X(n6944) );
  nand_x1_sg U40350 ( .A(n7630), .B(n47100), .X(n6945) );
  nand_x1_sg U40351 ( .A(n23124), .B(n42106), .X(n40158) );
  nand_x1_sg U40352 ( .A(n40631), .B(n40686), .X(n7947) );
  nand_x1_sg U40353 ( .A(n47167), .B(n7948), .X(n7944) );
  nand_x1_sg U40354 ( .A(n7956), .B(n7955), .X(n7957) );
  nand_x1_sg U40355 ( .A(n8001), .B(n8002), .X(n7984) );
  nand_x1_sg U40356 ( .A(n8023), .B(n8024), .X(n8010) );
  inv_x1_sg U40357 ( .A(n8026), .X(n47182) );
  nand_x1_sg U40358 ( .A(n47181), .B(n8043), .X(n8026) );
  nand_x1_sg U40359 ( .A(n8048), .B(n8049), .X(n8046) );
  nand_x1_sg U40360 ( .A(n47211), .B(n8104), .X(n8094) );
  nand_x1_sg U40361 ( .A(n8063), .B(n8064), .X(n8062) );
  nand_x2_sg U40362 ( .A(n8111), .B(n8112), .X(n8109) );
  inv_x1_sg U40363 ( .A(n8176), .X(n47260) );
  nand_x1_sg U40364 ( .A(n8190), .B(n8191), .X(n8176) );
  nand_x1_sg U40365 ( .A(n8138), .B(n8139), .X(n8140) );
  nand_x1_sg U40366 ( .A(n8216), .B(n8217), .X(n8202) );
  nand_x1_sg U40367 ( .A(n8219), .B(n47308), .X(n8216) );
  nand_x2_sg U40368 ( .A(n8278), .B(n8279), .X(n8234) );
  nand_x1_sg U40369 ( .A(n8235), .B(n8234), .X(n8232) );
  nand_x1_sg U40370 ( .A(n8342), .B(n8341), .X(n8334) );
  nand_x1_sg U40371 ( .A(n8334), .B(n47371), .X(n8329) );
  nand_x1_sg U40372 ( .A(n8362), .B(n8361), .X(n7859) );
  nand_x1_sg U40373 ( .A(n8408), .B(n8409), .X(n7778) );
  nand_x1_sg U40374 ( .A(n8397), .B(n8396), .X(n7764) );
  nand_x1_sg U40375 ( .A(n8392), .B(n8393), .X(n7767) );
  nand_x1_sg U40376 ( .A(n8452), .B(n47380), .X(n7761) );
  nand_x1_sg U40377 ( .A(n8448), .B(n47386), .X(n7762) );
  nand_x1_sg U40378 ( .A(n40626), .B(n40691), .X(n8765) );
  nand_x1_sg U40379 ( .A(n47452), .B(n8766), .X(n8762) );
  nand_x1_sg U40380 ( .A(n8774), .B(n8773), .X(n8775) );
  nand_x1_sg U40381 ( .A(n8819), .B(n8820), .X(n8802) );
  nand_x1_sg U40382 ( .A(n8841), .B(n8842), .X(n8828) );
  inv_x1_sg U40383 ( .A(n8844), .X(n47467) );
  nand_x1_sg U40384 ( .A(n47466), .B(n8861), .X(n8844) );
  nand_x1_sg U40385 ( .A(n8866), .B(n8867), .X(n8864) );
  nand_x1_sg U40386 ( .A(n47496), .B(n8922), .X(n8912) );
  nand_x1_sg U40387 ( .A(n8881), .B(n8882), .X(n8880) );
  nand_x2_sg U40388 ( .A(n8929), .B(n8930), .X(n8927) );
  inv_x1_sg U40389 ( .A(n8994), .X(n47545) );
  nand_x1_sg U40390 ( .A(n9008), .B(n9009), .X(n8994) );
  nand_x1_sg U40391 ( .A(n8956), .B(n8957), .X(n8958) );
  nand_x1_sg U40392 ( .A(n9034), .B(n9035), .X(n9020) );
  nand_x1_sg U40393 ( .A(n9037), .B(n47593), .X(n9034) );
  nand_x2_sg U40394 ( .A(n9096), .B(n9097), .X(n9052) );
  nand_x1_sg U40395 ( .A(n9053), .B(n9052), .X(n9050) );
  nand_x1_sg U40396 ( .A(n9160), .B(n9159), .X(n9152) );
  nand_x1_sg U40397 ( .A(n9152), .B(n47656), .X(n9147) );
  nand_x1_sg U40398 ( .A(n9180), .B(n9179), .X(n8677) );
  nand_x1_sg U40399 ( .A(n9226), .B(n9227), .X(n8596) );
  nand_x1_sg U40400 ( .A(n9215), .B(n9214), .X(n8582) );
  nand_x1_sg U40401 ( .A(n9210), .B(n9211), .X(n8585) );
  nand_x1_sg U40402 ( .A(n9270), .B(n47665), .X(n8579) );
  nand_x1_sg U40403 ( .A(n9266), .B(n47671), .X(n8580) );
  nand_x1_sg U40404 ( .A(n40666), .B(n40696), .X(n9585) );
  nand_x1_sg U40405 ( .A(n47737), .B(n9586), .X(n9582) );
  nand_x1_sg U40406 ( .A(n9594), .B(n9593), .X(n9595) );
  nand_x1_sg U40407 ( .A(n9639), .B(n9640), .X(n9622) );
  nand_x1_sg U40408 ( .A(n9661), .B(n9662), .X(n9648) );
  inv_x1_sg U40409 ( .A(n9664), .X(n47752) );
  nand_x1_sg U40410 ( .A(n47751), .B(n9681), .X(n9664) );
  nand_x1_sg U40411 ( .A(n9686), .B(n9687), .X(n9684) );
  nand_x1_sg U40412 ( .A(n47781), .B(n9742), .X(n9732) );
  nand_x1_sg U40413 ( .A(n9701), .B(n9702), .X(n9700) );
  nand_x2_sg U40414 ( .A(n9749), .B(n9750), .X(n9747) );
  inv_x1_sg U40415 ( .A(n9814), .X(n47830) );
  nand_x1_sg U40416 ( .A(n9828), .B(n9829), .X(n9814) );
  nand_x1_sg U40417 ( .A(n9776), .B(n9777), .X(n9778) );
  nand_x1_sg U40418 ( .A(n9854), .B(n9855), .X(n9840) );
  nand_x1_sg U40419 ( .A(n9857), .B(n47878), .X(n9854) );
  nand_x2_sg U40420 ( .A(n9916), .B(n9917), .X(n9872) );
  nand_x1_sg U40421 ( .A(n9873), .B(n9872), .X(n9870) );
  nand_x1_sg U40422 ( .A(n9980), .B(n9979), .X(n9972) );
  nand_x1_sg U40423 ( .A(n9972), .B(n47941), .X(n9967) );
  nand_x1_sg U40424 ( .A(n10000), .B(n9999), .X(n9497) );
  nand_x1_sg U40425 ( .A(n10046), .B(n10047), .X(n9416) );
  nand_x1_sg U40426 ( .A(n10035), .B(n10034), .X(n9402) );
  nand_x1_sg U40427 ( .A(n10030), .B(n10031), .X(n9405) );
  nand_x1_sg U40428 ( .A(n10090), .B(n47950), .X(n9399) );
  nand_x1_sg U40429 ( .A(n10086), .B(n47956), .X(n9400) );
  nand_x1_sg U40430 ( .A(n40656), .B(n40701), .X(n10404) );
  nand_x1_sg U40431 ( .A(n48022), .B(n10405), .X(n10401) );
  nand_x1_sg U40432 ( .A(n10413), .B(n10412), .X(n10414) );
  nand_x1_sg U40433 ( .A(n10458), .B(n10459), .X(n10441) );
  nand_x1_sg U40434 ( .A(n10480), .B(n10481), .X(n10467) );
  inv_x1_sg U40435 ( .A(n10483), .X(n48037) );
  nand_x1_sg U40436 ( .A(n48036), .B(n10500), .X(n10483) );
  nand_x1_sg U40437 ( .A(n10505), .B(n10506), .X(n10503) );
  nand_x1_sg U40438 ( .A(n48066), .B(n10561), .X(n10551) );
  nand_x1_sg U40439 ( .A(n10520), .B(n10521), .X(n10519) );
  nand_x2_sg U40440 ( .A(n10568), .B(n10569), .X(n10566) );
  inv_x1_sg U40441 ( .A(n10633), .X(n48115) );
  nand_x1_sg U40442 ( .A(n10647), .B(n10648), .X(n10633) );
  nand_x1_sg U40443 ( .A(n10595), .B(n10596), .X(n10597) );
  nand_x1_sg U40444 ( .A(n10673), .B(n10674), .X(n10659) );
  nand_x1_sg U40445 ( .A(n10676), .B(n48163), .X(n10673) );
  nand_x2_sg U40446 ( .A(n10735), .B(n10736), .X(n10691) );
  nand_x1_sg U40447 ( .A(n10692), .B(n10691), .X(n10689) );
  nand_x1_sg U40448 ( .A(n10799), .B(n10798), .X(n10791) );
  nand_x1_sg U40449 ( .A(n10791), .B(n48226), .X(n10786) );
  nand_x1_sg U40450 ( .A(n10819), .B(n10818), .X(n10316) );
  nand_x1_sg U40451 ( .A(n10865), .B(n10866), .X(n10235) );
  nand_x1_sg U40452 ( .A(n10854), .B(n10853), .X(n10221) );
  nand_x1_sg U40453 ( .A(n10849), .B(n10850), .X(n10224) );
  nand_x1_sg U40454 ( .A(n10909), .B(n48235), .X(n10218) );
  nand_x1_sg U40455 ( .A(n10905), .B(n48241), .X(n10219) );
  nand_x1_sg U40456 ( .A(n40641), .B(n40706), .X(n11223) );
  nand_x1_sg U40457 ( .A(n48307), .B(n11224), .X(n11220) );
  nand_x1_sg U40458 ( .A(n11232), .B(n11231), .X(n11233) );
  nand_x1_sg U40459 ( .A(n11277), .B(n11278), .X(n11260) );
  nand_x1_sg U40460 ( .A(n11299), .B(n11300), .X(n11286) );
  inv_x1_sg U40461 ( .A(n11302), .X(n48322) );
  nand_x1_sg U40462 ( .A(n48321), .B(n11319), .X(n11302) );
  nand_x1_sg U40463 ( .A(n11324), .B(n11325), .X(n11322) );
  nand_x1_sg U40464 ( .A(n48351), .B(n11380), .X(n11370) );
  nand_x1_sg U40465 ( .A(n11339), .B(n11340), .X(n11338) );
  nand_x2_sg U40466 ( .A(n11387), .B(n11388), .X(n11385) );
  inv_x1_sg U40467 ( .A(n11452), .X(n48400) );
  nand_x1_sg U40468 ( .A(n11466), .B(n11467), .X(n11452) );
  nand_x1_sg U40469 ( .A(n11414), .B(n11415), .X(n11416) );
  nand_x1_sg U40470 ( .A(n11492), .B(n11493), .X(n11478) );
  nand_x1_sg U40471 ( .A(n11495), .B(n48448), .X(n11492) );
  nand_x2_sg U40472 ( .A(n11554), .B(n11555), .X(n11510) );
  nand_x1_sg U40473 ( .A(n11511), .B(n11510), .X(n11508) );
  nand_x1_sg U40474 ( .A(n11618), .B(n11617), .X(n11610) );
  nand_x1_sg U40475 ( .A(n11610), .B(n48511), .X(n11605) );
  nand_x1_sg U40476 ( .A(n11638), .B(n11637), .X(n11135) );
  nand_x1_sg U40477 ( .A(n11684), .B(n11685), .X(n11054) );
  nand_x1_sg U40478 ( .A(n11673), .B(n11672), .X(n11040) );
  nand_x1_sg U40479 ( .A(n11668), .B(n11669), .X(n11043) );
  nand_x1_sg U40480 ( .A(n11728), .B(n48520), .X(n11037) );
  nand_x1_sg U40481 ( .A(n11724), .B(n48526), .X(n11038) );
  nand_x1_sg U40482 ( .A(n40636), .B(n40711), .X(n12042) );
  nand_x1_sg U40483 ( .A(n48592), .B(n12043), .X(n12039) );
  nand_x1_sg U40484 ( .A(n12051), .B(n12050), .X(n12052) );
  nand_x1_sg U40485 ( .A(n12096), .B(n12097), .X(n12079) );
  nand_x1_sg U40486 ( .A(n12118), .B(n12119), .X(n12105) );
  inv_x1_sg U40487 ( .A(n12121), .X(n48607) );
  nand_x1_sg U40488 ( .A(n48606), .B(n12138), .X(n12121) );
  nand_x1_sg U40489 ( .A(n12143), .B(n12144), .X(n12141) );
  nand_x1_sg U40490 ( .A(n48636), .B(n12199), .X(n12189) );
  nand_x1_sg U40491 ( .A(n12158), .B(n12159), .X(n12157) );
  nand_x2_sg U40492 ( .A(n12206), .B(n12207), .X(n12204) );
  inv_x1_sg U40493 ( .A(n12271), .X(n48685) );
  nand_x1_sg U40494 ( .A(n12285), .B(n12286), .X(n12271) );
  nand_x1_sg U40495 ( .A(n12233), .B(n12234), .X(n12235) );
  nand_x1_sg U40496 ( .A(n12311), .B(n12312), .X(n12297) );
  nand_x1_sg U40497 ( .A(n12314), .B(n48733), .X(n12311) );
  nand_x2_sg U40498 ( .A(n12373), .B(n12374), .X(n12329) );
  nand_x1_sg U40499 ( .A(n12330), .B(n12329), .X(n12327) );
  nand_x1_sg U40500 ( .A(n12437), .B(n12436), .X(n12429) );
  nand_x1_sg U40501 ( .A(n12429), .B(n48796), .X(n12424) );
  nand_x1_sg U40502 ( .A(n12457), .B(n12456), .X(n11954) );
  nand_x1_sg U40503 ( .A(n12503), .B(n12504), .X(n11873) );
  nand_x1_sg U40504 ( .A(n12492), .B(n12491), .X(n11859) );
  nand_x1_sg U40505 ( .A(n12487), .B(n12488), .X(n11862) );
  nand_x1_sg U40506 ( .A(n12547), .B(n48805), .X(n11856) );
  nand_x1_sg U40507 ( .A(n12543), .B(n48811), .X(n11857) );
  nand_x1_sg U40508 ( .A(n40661), .B(n40716), .X(n12861) );
  nand_x1_sg U40509 ( .A(n48878), .B(n12862), .X(n12858) );
  nand_x1_sg U40510 ( .A(n12870), .B(n12869), .X(n12871) );
  nand_x1_sg U40511 ( .A(n12915), .B(n12916), .X(n12898) );
  nand_x1_sg U40512 ( .A(n12937), .B(n12938), .X(n12924) );
  inv_x1_sg U40513 ( .A(n12940), .X(n48893) );
  nand_x1_sg U40514 ( .A(n48892), .B(n12957), .X(n12940) );
  nand_x1_sg U40515 ( .A(n12962), .B(n12963), .X(n12960) );
  nand_x1_sg U40516 ( .A(n48922), .B(n13018), .X(n13008) );
  nand_x1_sg U40517 ( .A(n12977), .B(n12978), .X(n12976) );
  nand_x2_sg U40518 ( .A(n13025), .B(n13026), .X(n13023) );
  inv_x1_sg U40519 ( .A(n13090), .X(n48971) );
  nand_x1_sg U40520 ( .A(n13104), .B(n13105), .X(n13090) );
  nand_x1_sg U40521 ( .A(n13052), .B(n13053), .X(n13054) );
  nand_x1_sg U40522 ( .A(n13130), .B(n13131), .X(n13116) );
  nand_x1_sg U40523 ( .A(n13133), .B(n49019), .X(n13130) );
  nand_x2_sg U40524 ( .A(n13192), .B(n13193), .X(n13148) );
  nand_x1_sg U40525 ( .A(n13149), .B(n13148), .X(n13146) );
  nand_x1_sg U40526 ( .A(n13256), .B(n13255), .X(n13248) );
  nand_x1_sg U40527 ( .A(n13248), .B(n49083), .X(n13243) );
  nand_x1_sg U40528 ( .A(n13276), .B(n13275), .X(n12773) );
  nand_x1_sg U40529 ( .A(n13322), .B(n13323), .X(n12692) );
  nand_x1_sg U40530 ( .A(n13311), .B(n13310), .X(n12678) );
  nand_x1_sg U40531 ( .A(n13306), .B(n13307), .X(n12681) );
  nand_x1_sg U40532 ( .A(n13366), .B(n49092), .X(n12675) );
  nand_x1_sg U40533 ( .A(n13362), .B(n49098), .X(n12676) );
  nand_x1_sg U40534 ( .A(n40651), .B(n40721), .X(n13680) );
  nand_x1_sg U40535 ( .A(n49165), .B(n13681), .X(n13677) );
  nand_x1_sg U40536 ( .A(n13689), .B(n13688), .X(n13690) );
  nand_x1_sg U40537 ( .A(n13734), .B(n13735), .X(n13717) );
  nand_x1_sg U40538 ( .A(n13756), .B(n13757), .X(n13743) );
  inv_x1_sg U40539 ( .A(n13759), .X(n49180) );
  nand_x1_sg U40540 ( .A(n49179), .B(n13776), .X(n13759) );
  nand_x1_sg U40541 ( .A(n13781), .B(n13782), .X(n13779) );
  nand_x1_sg U40542 ( .A(n49209), .B(n13837), .X(n13827) );
  nand_x1_sg U40543 ( .A(n13796), .B(n13797), .X(n13795) );
  nand_x2_sg U40544 ( .A(n13844), .B(n13845), .X(n13842) );
  inv_x1_sg U40545 ( .A(n13909), .X(n49258) );
  nand_x1_sg U40546 ( .A(n13923), .B(n13924), .X(n13909) );
  nand_x1_sg U40547 ( .A(n13871), .B(n13872), .X(n13873) );
  nand_x1_sg U40548 ( .A(n13949), .B(n13950), .X(n13935) );
  nand_x1_sg U40549 ( .A(n13952), .B(n49306), .X(n13949) );
  nand_x2_sg U40550 ( .A(n14011), .B(n14012), .X(n13967) );
  nand_x1_sg U40551 ( .A(n13968), .B(n13967), .X(n13965) );
  nand_x1_sg U40552 ( .A(n14075), .B(n14074), .X(n14067) );
  nand_x1_sg U40553 ( .A(n14067), .B(n49369), .X(n14062) );
  nand_x1_sg U40554 ( .A(n14095), .B(n14094), .X(n13592) );
  nand_x1_sg U40555 ( .A(n14141), .B(n14142), .X(n13511) );
  nand_x1_sg U40556 ( .A(n14130), .B(n14129), .X(n13497) );
  nand_x1_sg U40557 ( .A(n14125), .B(n14126), .X(n13500) );
  nand_x1_sg U40558 ( .A(n14185), .B(n49378), .X(n13494) );
  nand_x1_sg U40559 ( .A(n14181), .B(n49384), .X(n13495) );
  nand_x1_sg U40560 ( .A(n40621), .B(n40726), .X(n14499) );
  nand_x1_sg U40561 ( .A(n49451), .B(n14500), .X(n14496) );
  nand_x1_sg U40562 ( .A(n14508), .B(n14507), .X(n14509) );
  nand_x1_sg U40563 ( .A(n14553), .B(n14554), .X(n14536) );
  nand_x1_sg U40564 ( .A(n14575), .B(n14576), .X(n14562) );
  inv_x1_sg U40565 ( .A(n14578), .X(n49466) );
  nand_x1_sg U40566 ( .A(n49465), .B(n14595), .X(n14578) );
  nand_x1_sg U40567 ( .A(n14600), .B(n14601), .X(n14598) );
  nand_x1_sg U40568 ( .A(n49495), .B(n14656), .X(n14646) );
  nand_x1_sg U40569 ( .A(n14615), .B(n14616), .X(n14614) );
  nand_x2_sg U40570 ( .A(n14663), .B(n14664), .X(n14661) );
  inv_x1_sg U40571 ( .A(n14728), .X(n49544) );
  nand_x1_sg U40572 ( .A(n14742), .B(n14743), .X(n14728) );
  nand_x1_sg U40573 ( .A(n14690), .B(n14691), .X(n14692) );
  nand_x1_sg U40574 ( .A(n14768), .B(n14769), .X(n14754) );
  nand_x1_sg U40575 ( .A(n14771), .B(n49592), .X(n14768) );
  nand_x2_sg U40576 ( .A(n14830), .B(n14831), .X(n14786) );
  nand_x1_sg U40577 ( .A(n14787), .B(n14786), .X(n14784) );
  nand_x1_sg U40578 ( .A(n14894), .B(n14893), .X(n14886) );
  nand_x1_sg U40579 ( .A(n14886), .B(n49655), .X(n14881) );
  nand_x1_sg U40580 ( .A(n14914), .B(n14913), .X(n14411) );
  nand_x1_sg U40581 ( .A(n14960), .B(n14961), .X(n14330) );
  nand_x1_sg U40582 ( .A(n14949), .B(n14948), .X(n14316) );
  nand_x1_sg U40583 ( .A(n14944), .B(n14945), .X(n14319) );
  nand_x1_sg U40584 ( .A(n15004), .B(n49664), .X(n14313) );
  nand_x1_sg U40585 ( .A(n15000), .B(n49670), .X(n14314) );
  nand_x1_sg U40586 ( .A(n40681), .B(n40731), .X(n15318) );
  nand_x1_sg U40587 ( .A(n49736), .B(n15319), .X(n15315) );
  nand_x1_sg U40588 ( .A(n15327), .B(n15326), .X(n15328) );
  nand_x1_sg U40589 ( .A(n15372), .B(n15373), .X(n15355) );
  nand_x1_sg U40590 ( .A(n15394), .B(n15395), .X(n15381) );
  inv_x1_sg U40591 ( .A(n15397), .X(n49751) );
  nand_x1_sg U40592 ( .A(n49750), .B(n15414), .X(n15397) );
  nand_x1_sg U40593 ( .A(n15419), .B(n15420), .X(n15417) );
  nand_x1_sg U40594 ( .A(n49781), .B(n15475), .X(n15465) );
  nand_x1_sg U40595 ( .A(n15434), .B(n15435), .X(n15433) );
  nand_x2_sg U40596 ( .A(n15482), .B(n15483), .X(n15480) );
  inv_x1_sg U40597 ( .A(n15547), .X(n49830) );
  nand_x1_sg U40598 ( .A(n15561), .B(n15562), .X(n15547) );
  nand_x1_sg U40599 ( .A(n15509), .B(n15510), .X(n15511) );
  nand_x1_sg U40600 ( .A(n15587), .B(n15588), .X(n15573) );
  nand_x1_sg U40601 ( .A(n15590), .B(n49878), .X(n15587) );
  nand_x2_sg U40602 ( .A(n15649), .B(n15650), .X(n15605) );
  nand_x1_sg U40603 ( .A(n15606), .B(n15605), .X(n15603) );
  nand_x1_sg U40604 ( .A(n15713), .B(n15712), .X(n15705) );
  nand_x1_sg U40605 ( .A(n15705), .B(n49941), .X(n15700) );
  nand_x1_sg U40606 ( .A(n15733), .B(n15732), .X(n15230) );
  nand_x1_sg U40607 ( .A(n15779), .B(n15780), .X(n15149) );
  nand_x1_sg U40608 ( .A(n15768), .B(n15767), .X(n15135) );
  nand_x1_sg U40609 ( .A(n15763), .B(n15764), .X(n15138) );
  nand_x1_sg U40610 ( .A(n15823), .B(n49950), .X(n15132) );
  nand_x1_sg U40611 ( .A(n15819), .B(n49956), .X(n15133) );
  nand_x1_sg U40612 ( .A(n40676), .B(n40736), .X(n16137) );
  nand_x1_sg U40613 ( .A(n50023), .B(n16138), .X(n16134) );
  nand_x1_sg U40614 ( .A(n16146), .B(n16145), .X(n16147) );
  nand_x1_sg U40615 ( .A(n16191), .B(n16192), .X(n16174) );
  nand_x1_sg U40616 ( .A(n16213), .B(n16214), .X(n16200) );
  inv_x1_sg U40617 ( .A(n16216), .X(n50038) );
  nand_x1_sg U40618 ( .A(n50037), .B(n16233), .X(n16216) );
  nand_x1_sg U40619 ( .A(n16238), .B(n16239), .X(n16236) );
  nand_x1_sg U40620 ( .A(n50067), .B(n16294), .X(n16284) );
  nand_x1_sg U40621 ( .A(n16253), .B(n16254), .X(n16252) );
  nand_x2_sg U40622 ( .A(n16301), .B(n16302), .X(n16299) );
  inv_x1_sg U40623 ( .A(n16366), .X(n50116) );
  nand_x1_sg U40624 ( .A(n16380), .B(n16381), .X(n16366) );
  nand_x1_sg U40625 ( .A(n16328), .B(n16329), .X(n16330) );
  nand_x1_sg U40626 ( .A(n16406), .B(n16407), .X(n16392) );
  nand_x1_sg U40627 ( .A(n16409), .B(n50164), .X(n16406) );
  nand_x2_sg U40628 ( .A(n16468), .B(n16469), .X(n16424) );
  nand_x1_sg U40629 ( .A(n16425), .B(n16424), .X(n16422) );
  nand_x1_sg U40630 ( .A(n16532), .B(n16531), .X(n16524) );
  nand_x1_sg U40631 ( .A(n16524), .B(n50227), .X(n16519) );
  nand_x1_sg U40632 ( .A(n16552), .B(n16551), .X(n16049) );
  nand_x1_sg U40633 ( .A(n16598), .B(n16599), .X(n15968) );
  nand_x1_sg U40634 ( .A(n16587), .B(n16586), .X(n15954) );
  nand_x1_sg U40635 ( .A(n16582), .B(n16583), .X(n15957) );
  nand_x1_sg U40636 ( .A(n16642), .B(n50236), .X(n15951) );
  nand_x1_sg U40637 ( .A(n16638), .B(n50242), .X(n15952) );
  nand_x1_sg U40638 ( .A(n50308), .B(n16955), .X(n16951) );
  nand_x1_sg U40639 ( .A(n16963), .B(n16962), .X(n16964) );
  nand_x1_sg U40640 ( .A(n17007), .B(n17008), .X(n16990) );
  nand_x1_sg U40641 ( .A(n17029), .B(n17030), .X(n17016) );
  inv_x1_sg U40642 ( .A(n17032), .X(n50323) );
  nand_x1_sg U40643 ( .A(n50322), .B(n17049), .X(n17032) );
  nand_x1_sg U40644 ( .A(n17054), .B(n17055), .X(n17052) );
  nand_x1_sg U40645 ( .A(n50352), .B(n17111), .X(n17100) );
  nand_x1_sg U40646 ( .A(n17069), .B(n17070), .X(n17068) );
  nand_x2_sg U40647 ( .A(n17118), .B(n17119), .X(n17116) );
  inv_x1_sg U40648 ( .A(n17183), .X(n50401) );
  nand_x1_sg U40649 ( .A(n17197), .B(n17198), .X(n17183) );
  nand_x1_sg U40650 ( .A(n17145), .B(n17146), .X(n17147) );
  nand_x2_sg U40651 ( .A(n17285), .B(n17286), .X(n17241) );
  nand_x1_sg U40652 ( .A(n17242), .B(n17241), .X(n17239) );
  nand_x1_sg U40653 ( .A(n17349), .B(n17348), .X(n17341) );
  nand_x1_sg U40654 ( .A(n17341), .B(n50512), .X(n17336) );
  nand_x1_sg U40655 ( .A(n17369), .B(n17368), .X(n16868) );
  nand_x1_sg U40656 ( .A(n17415), .B(n17416), .X(n16785) );
  nand_x1_sg U40657 ( .A(n17404), .B(n17403), .X(n16771) );
  nand_x1_sg U40658 ( .A(n17399), .B(n17400), .X(n16774) );
  nand_x1_sg U40659 ( .A(n17459), .B(n50521), .X(n16768) );
  nand_x1_sg U40660 ( .A(n17455), .B(n50527), .X(n16769) );
  nand_x1_sg U40661 ( .A(n50597), .B(n17776), .X(n17772) );
  nand_x1_sg U40662 ( .A(n17784), .B(n17783), .X(n17785) );
  nand_x1_sg U40663 ( .A(n17829), .B(n17830), .X(n17812) );
  nand_x1_sg U40664 ( .A(n17851), .B(n17852), .X(n17838) );
  inv_x1_sg U40665 ( .A(n17854), .X(n50612) );
  nand_x1_sg U40666 ( .A(n50611), .B(n17871), .X(n17854) );
  nand_x1_sg U40667 ( .A(n17876), .B(n17877), .X(n17874) );
  nand_x1_sg U40668 ( .A(n50641), .B(n17932), .X(n17922) );
  nand_x1_sg U40669 ( .A(n17891), .B(n17892), .X(n17890) );
  nand_x2_sg U40670 ( .A(n17939), .B(n17940), .X(n17937) );
  inv_x1_sg U40671 ( .A(n18004), .X(n50690) );
  nand_x1_sg U40672 ( .A(n18018), .B(n18019), .X(n18004) );
  nand_x1_sg U40673 ( .A(n17966), .B(n17967), .X(n17968) );
  nand_x1_sg U40674 ( .A(n18044), .B(n18045), .X(n18030) );
  nand_x1_sg U40675 ( .A(n18047), .B(n50738), .X(n18044) );
  nand_x2_sg U40676 ( .A(n18106), .B(n18107), .X(n18062) );
  nand_x1_sg U40677 ( .A(n18063), .B(n18062), .X(n18060) );
  nand_x1_sg U40678 ( .A(n18170), .B(n18169), .X(n18162) );
  nand_x1_sg U40679 ( .A(n18162), .B(n50801), .X(n18157) );
  nand_x1_sg U40680 ( .A(n18190), .B(n18189), .X(n17687) );
  nand_x1_sg U40681 ( .A(n18236), .B(n18237), .X(n17606) );
  nand_x1_sg U40682 ( .A(n18225), .B(n18224), .X(n17592) );
  nand_x1_sg U40683 ( .A(n18220), .B(n18221), .X(n17595) );
  nand_x1_sg U40684 ( .A(n18280), .B(n50810), .X(n17589) );
  nand_x1_sg U40685 ( .A(n18276), .B(n50816), .X(n17590) );
  nand_x1_sg U40686 ( .A(n40671), .B(n40741), .X(n18596) );
  nand_x1_sg U40687 ( .A(n50884), .B(n18597), .X(n18593) );
  nand_x1_sg U40688 ( .A(n18605), .B(n18604), .X(n18606) );
  nand_x1_sg U40689 ( .A(n18650), .B(n18651), .X(n18633) );
  nand_x1_sg U40690 ( .A(n18672), .B(n18673), .X(n18659) );
  inv_x1_sg U40691 ( .A(n18675), .X(n50899) );
  nand_x1_sg U40692 ( .A(n50898), .B(n18692), .X(n18675) );
  nand_x1_sg U40693 ( .A(n18697), .B(n18698), .X(n18695) );
  nand_x1_sg U40694 ( .A(n50928), .B(n18753), .X(n18743) );
  nand_x1_sg U40695 ( .A(n18712), .B(n18713), .X(n18711) );
  nand_x2_sg U40696 ( .A(n18760), .B(n18761), .X(n18758) );
  inv_x1_sg U40697 ( .A(n18825), .X(n50977) );
  nand_x1_sg U40698 ( .A(n18839), .B(n18840), .X(n18825) );
  nand_x1_sg U40699 ( .A(n18787), .B(n18788), .X(n18789) );
  nand_x1_sg U40700 ( .A(n18865), .B(n18866), .X(n18851) );
  nand_x1_sg U40701 ( .A(n18868), .B(n51025), .X(n18865) );
  nand_x2_sg U40702 ( .A(n18927), .B(n18928), .X(n18883) );
  nand_x1_sg U40703 ( .A(n18884), .B(n18883), .X(n18881) );
  nand_x1_sg U40704 ( .A(n18991), .B(n18990), .X(n18983) );
  nand_x1_sg U40705 ( .A(n18983), .B(n51088), .X(n18978) );
  nand_x1_sg U40706 ( .A(n19011), .B(n19010), .X(n18508) );
  nand_x1_sg U40707 ( .A(n19057), .B(n19058), .X(n18427) );
  nand_x1_sg U40708 ( .A(n19046), .B(n19045), .X(n18413) );
  nand_x1_sg U40709 ( .A(n19041), .B(n19042), .X(n18416) );
  nand_x1_sg U40710 ( .A(n19101), .B(n51097), .X(n18410) );
  nand_x1_sg U40711 ( .A(n19097), .B(n51103), .X(n18411) );
  nand_x1_sg U40712 ( .A(n5265), .B(n26845), .X(n26844) );
  nand_x1_sg U40713 ( .A(n5208), .B(n26868), .X(n26867) );
  nand_x1_sg U40714 ( .A(n5246), .B(n26854), .X(n26853) );
  nand_x1_sg U40715 ( .A(n5189), .B(n26875), .X(n26874) );
  nand_x1_sg U40716 ( .A(n5227), .B(n26861), .X(n26860) );
  inv_x1_sg U40717 ( .A(n21752), .X(n45751) );
  inv_x1_sg U40718 ( .A(n21736), .X(n45755) );
  inv_x1_sg U40719 ( .A(n21735), .X(n45761) );
  inv_x1_sg U40720 ( .A(n21741), .X(n45759) );
  inv_x1_sg U40721 ( .A(n21731), .X(n45757) );
  inv_x1_sg U40722 ( .A(n21732), .X(n45763) );
  inv_x1_sg U40723 ( .A(n21799), .X(n45708) );
  inv_x1_sg U40724 ( .A(n21783), .X(n45712) );
  inv_x1_sg U40725 ( .A(n21782), .X(n45718) );
  inv_x1_sg U40726 ( .A(n21788), .X(n45716) );
  inv_x1_sg U40727 ( .A(n21778), .X(n45714) );
  inv_x1_sg U40728 ( .A(n21779), .X(n45720) );
  inv_x1_sg U40729 ( .A(n21846), .X(n45664) );
  inv_x1_sg U40730 ( .A(n21830), .X(n45669) );
  inv_x1_sg U40731 ( .A(n21829), .X(n45675) );
  inv_x1_sg U40732 ( .A(n21835), .X(n45673) );
  inv_x1_sg U40733 ( .A(n21825), .X(n45671) );
  inv_x1_sg U40734 ( .A(n21826), .X(n45677) );
  inv_x1_sg U40735 ( .A(n21892), .X(n45620) );
  inv_x1_sg U40736 ( .A(n21877), .X(n45625) );
  inv_x1_sg U40737 ( .A(n21876), .X(n45631) );
  inv_x1_sg U40738 ( .A(n21882), .X(n45629) );
  inv_x1_sg U40739 ( .A(n21872), .X(n45627) );
  inv_x1_sg U40740 ( .A(n21873), .X(n45633) );
  inv_x1_sg U40741 ( .A(n21939), .X(n45576) );
  inv_x1_sg U40742 ( .A(n21923), .X(n45581) );
  inv_x1_sg U40743 ( .A(n21922), .X(n45587) );
  inv_x1_sg U40744 ( .A(n21928), .X(n45585) );
  inv_x1_sg U40745 ( .A(n21918), .X(n45583) );
  inv_x1_sg U40746 ( .A(n21919), .X(n45589) );
  inv_x1_sg U40747 ( .A(n21985), .X(n45531) );
  inv_x1_sg U40748 ( .A(n21975), .X(n45540) );
  inv_x1_sg U40749 ( .A(n21970), .X(n45536) );
  inv_x1_sg U40750 ( .A(n21969), .X(n45542) );
  inv_x1_sg U40751 ( .A(n21965), .X(n45538) );
  inv_x1_sg U40752 ( .A(n21966), .X(n45544) );
  inv_x1_sg U40753 ( .A(n22032), .X(n45487) );
  inv_x1_sg U40754 ( .A(n22016), .X(n45492) );
  inv_x1_sg U40755 ( .A(n22015), .X(n45498) );
  inv_x1_sg U40756 ( .A(n22021), .X(n45496) );
  inv_x1_sg U40757 ( .A(n22011), .X(n45494) );
  inv_x1_sg U40758 ( .A(n22012), .X(n45500) );
  inv_x1_sg U40759 ( .A(n22078), .X(n45442) );
  inv_x1_sg U40760 ( .A(n22063), .X(n45444) );
  inv_x1_sg U40761 ( .A(n22062), .X(n45450) );
  inv_x1_sg U40762 ( .A(n22068), .X(n45448) );
  inv_x1_sg U40763 ( .A(n22058), .X(n45446) );
  inv_x1_sg U40764 ( .A(n22059), .X(n45452) );
  inv_x1_sg U40765 ( .A(n28315), .X(n45378) );
  nand_x1_sg U40766 ( .A(n28339), .B(n28340), .X(n28315) );
  inv_x1_sg U40767 ( .A(n22114), .X(n45404) );
  inv_x1_sg U40768 ( .A(n22109), .X(n45400) );
  inv_x1_sg U40769 ( .A(n22108), .X(n45406) );
  inv_x1_sg U40770 ( .A(n22104), .X(n45402) );
  inv_x1_sg U40771 ( .A(n22105), .X(n45408) );
  inv_x1_sg U40772 ( .A(n28309), .X(n45333) );
  nand_x1_sg U40773 ( .A(n28342), .B(n28343), .X(n28309) );
  inv_x1_sg U40774 ( .A(n22162), .X(n45358) );
  inv_x1_sg U40775 ( .A(n22157), .X(n45354) );
  inv_x1_sg U40776 ( .A(n22156), .X(n45360) );
  inv_x1_sg U40777 ( .A(n22152), .X(n45356) );
  inv_x1_sg U40778 ( .A(n22153), .X(n45362) );
  inv_x1_sg U40779 ( .A(n28303), .X(n45288) );
  nand_x1_sg U40780 ( .A(n28345), .B(n28346), .X(n28303) );
  inv_x1_sg U40781 ( .A(n22209), .X(n45313) );
  inv_x1_sg U40782 ( .A(n22204), .X(n45309) );
  inv_x1_sg U40783 ( .A(n22203), .X(n45315) );
  inv_x1_sg U40784 ( .A(n22199), .X(n45311) );
  inv_x1_sg U40785 ( .A(n22200), .X(n45317) );
  inv_x1_sg U40786 ( .A(n28297), .X(n45243) );
  nand_x1_sg U40787 ( .A(n28348), .B(n28349), .X(n28297) );
  inv_x1_sg U40788 ( .A(n22252), .X(n45264) );
  inv_x1_sg U40789 ( .A(n22251), .X(n45270) );
  inv_x1_sg U40790 ( .A(n22257), .X(n45268) );
  inv_x1_sg U40791 ( .A(n22247), .X(n45266) );
  inv_x1_sg U40792 ( .A(n22248), .X(n45272) );
  inv_x1_sg U40793 ( .A(n28291), .X(n45197) );
  nand_x1_sg U40794 ( .A(n28351), .B(n28352), .X(n28291) );
  inv_x1_sg U40795 ( .A(n22304), .X(n45223) );
  inv_x1_sg U40796 ( .A(n22299), .X(n45219) );
  inv_x1_sg U40797 ( .A(n22298), .X(n45225) );
  inv_x1_sg U40798 ( .A(n22294), .X(n45221) );
  inv_x1_sg U40799 ( .A(n22295), .X(n45227) );
  inv_x1_sg U40800 ( .A(n28285), .X(n45152) );
  nand_x1_sg U40801 ( .A(n28354), .B(n28355), .X(n28285) );
  inv_x1_sg U40802 ( .A(n22352), .X(n45177) );
  inv_x1_sg U40803 ( .A(n22347), .X(n45173) );
  inv_x1_sg U40804 ( .A(n22346), .X(n45179) );
  inv_x1_sg U40805 ( .A(n22342), .X(n45175) );
  inv_x1_sg U40806 ( .A(n22343), .X(n45181) );
  inv_x1_sg U40807 ( .A(n28279), .X(n45106) );
  nand_x1_sg U40808 ( .A(n28357), .B(n28358), .X(n28279) );
  inv_x1_sg U40809 ( .A(n22394), .X(n45128) );
  inv_x1_sg U40810 ( .A(n22393), .X(n45134) );
  inv_x1_sg U40811 ( .A(n22399), .X(n45132) );
  inv_x1_sg U40812 ( .A(n22389), .X(n45130) );
  inv_x1_sg U40813 ( .A(n22390), .X(n45136) );
  inv_x1_sg U40814 ( .A(n28273), .X(n45060) );
  nand_x1_sg U40815 ( .A(n28360), .B(n28361), .X(n28273) );
  inv_x1_sg U40816 ( .A(n22446), .X(n45085) );
  inv_x1_sg U40817 ( .A(n22441), .X(n45087) );
  inv_x1_sg U40818 ( .A(n22437), .X(n45083) );
  inv_x1_sg U40819 ( .A(n22438), .X(n45089) );
  nand_x1_sg U40820 ( .A(n5301), .B(n28267), .X(n28266) );
  inv_x1_sg U40821 ( .A(n22503), .X(n45035) );
  nand_x1_sg U40822 ( .A(n5225), .B(n27628), .X(n27627) );
  inv_x1_sg U40823 ( .A(n22492), .X(n45041) );
  nand_x1_sg U40824 ( .A(n5263), .B(n27984), .X(n27983) );
  nand_x1_sg U40825 ( .A(n5206), .B(n27425), .X(n27424) );
  inv_x1_sg U40826 ( .A(n22487), .X(n45043) );
  nand_x1_sg U40827 ( .A(n5244), .B(n27814), .X(n27813) );
  inv_x1_sg U40828 ( .A(n22483), .X(n45039) );
  nand_x1_sg U40829 ( .A(n5187), .B(n27203), .X(n27202) );
  inv_x1_sg U40830 ( .A(n22484), .X(n45045) );
  inv_x1_sg U40831 ( .A(n22774), .X(n46924) );
  inv_x1_sg U40832 ( .A(n22760), .X(n46965) );
  inv_x1_sg U40833 ( .A(n22739), .X(n47026) );
  nand_x1_sg U40834 ( .A(n23117), .B(n23118), .X(n23111) );
  inv_x1_sg U40835 ( .A(n23051), .X(n47216) );
  inv_x1_sg U40836 ( .A(n23037), .X(n47255) );
  inv_x1_sg U40837 ( .A(n23023), .X(n47295) );
  inv_x1_sg U40838 ( .A(n23016), .X(n47313) );
  nand_x1_sg U40839 ( .A(n23397), .B(n23398), .X(n23391) );
  inv_x1_sg U40840 ( .A(n23317), .X(n47540) );
  inv_x1_sg U40841 ( .A(n23303), .X(n47580) );
  inv_x1_sg U40842 ( .A(n23296), .X(n47598) );
  nand_x1_sg U40843 ( .A(n23676), .B(n23677), .X(n23670) );
  inv_x1_sg U40844 ( .A(n23610), .X(n47786) );
  inv_x1_sg U40845 ( .A(n23596), .X(n47825) );
  inv_x1_sg U40846 ( .A(n23582), .X(n47865) );
  inv_x1_sg U40847 ( .A(n23575), .X(n47883) );
  nand_x1_sg U40848 ( .A(n23955), .B(n23956), .X(n23949) );
  inv_x1_sg U40849 ( .A(n23875), .X(n48110) );
  inv_x1_sg U40850 ( .A(n23861), .X(n48150) );
  inv_x1_sg U40851 ( .A(n23854), .X(n48168) );
  nand_x1_sg U40852 ( .A(n24234), .B(n24235), .X(n24228) );
  inv_x1_sg U40853 ( .A(n24168), .X(n48356) );
  inv_x1_sg U40854 ( .A(n24154), .X(n48395) );
  inv_x1_sg U40855 ( .A(n24140), .X(n48435) );
  inv_x1_sg U40856 ( .A(n24133), .X(n48453) );
  nand_x1_sg U40857 ( .A(n24513), .B(n24514), .X(n24507) );
  inv_x1_sg U40858 ( .A(n24447), .X(n48641) );
  inv_x1_sg U40859 ( .A(n24433), .X(n48680) );
  inv_x1_sg U40860 ( .A(n24419), .X(n48720) );
  inv_x1_sg U40861 ( .A(n24412), .X(n48738) );
  nand_x1_sg U40862 ( .A(n24791), .B(n24792), .X(n24785) );
  inv_x1_sg U40863 ( .A(n24725), .X(n48927) );
  inv_x1_sg U40864 ( .A(n24711), .X(n48966) );
  inv_x1_sg U40865 ( .A(n24697), .X(n49006) );
  inv_x1_sg U40866 ( .A(n24690), .X(n49024) );
  nand_x1_sg U40867 ( .A(n25070), .B(n25071), .X(n25064) );
  inv_x1_sg U40868 ( .A(n25004), .X(n49214) );
  inv_x1_sg U40869 ( .A(n24990), .X(n49253) );
  inv_x1_sg U40870 ( .A(n24976), .X(n49293) );
  inv_x1_sg U40871 ( .A(n24969), .X(n49311) );
  nand_x1_sg U40872 ( .A(n25349), .B(n25350), .X(n25343) );
  inv_x1_sg U40873 ( .A(n25283), .X(n49500) );
  inv_x1_sg U40874 ( .A(n25269), .X(n49539) );
  inv_x1_sg U40875 ( .A(n25255), .X(n49579) );
  nand_x1_sg U40876 ( .A(n25628), .B(n25629), .X(n25622) );
  inv_x1_sg U40877 ( .A(n25562), .X(n49786) );
  inv_x1_sg U40878 ( .A(n25548), .X(n49825) );
  inv_x1_sg U40879 ( .A(n25534), .X(n49865) );
  inv_x1_sg U40880 ( .A(n25527), .X(n49883) );
  nand_x1_sg U40881 ( .A(n25905), .B(n25906), .X(n25899) );
  inv_x1_sg U40882 ( .A(n25825), .X(n50111) );
  inv_x1_sg U40883 ( .A(n25811), .X(n50151) );
  inv_x1_sg U40884 ( .A(n25804), .X(n50169) );
  nand_x1_sg U40885 ( .A(n26174), .B(n26175), .X(n26120) );
  nand_x1_sg U40886 ( .A(n26165), .B(n26166), .X(n26102) );
  inv_x1_sg U40887 ( .A(n26071), .X(n50373) );
  nand_x1_sg U40888 ( .A(n26465), .B(n26466), .X(n26459) );
  inv_x1_sg U40889 ( .A(n26399), .X(n50646) );
  inv_x1_sg U40890 ( .A(n26385), .X(n50685) );
  inv_x1_sg U40891 ( .A(n26371), .X(n50725) );
  inv_x1_sg U40892 ( .A(n26364), .X(n50743) );
  nand_x1_sg U40893 ( .A(n26743), .B(n26744), .X(n26737) );
  inv_x1_sg U40894 ( .A(n26677), .X(n50933) );
  inv_x1_sg U40895 ( .A(n26663), .X(n50972) );
  inv_x1_sg U40896 ( .A(n26649), .X(n51012) );
  inv_x1_sg U40897 ( .A(n26642), .X(n51030) );
  nand_x1_sg U40898 ( .A(n5417), .B(n19148), .X(n19147) );
  nand_x1_sg U40899 ( .A(n5531), .B(n19538), .X(n19537) );
  nand_x1_sg U40900 ( .A(n20979), .B(n20980), .X(n20977) );
  nand_x1_sg U40901 ( .A(n5645), .B(n20993), .X(n20992) );
  nand_x1_sg U40902 ( .A(n5607), .B(n21008), .X(n21007) );
  inv_x1_sg U40903 ( .A(n19746), .X(n41539) );
  nand_x1_sg U40904 ( .A(n21177), .B(n46586), .X(n20999) );
  nand_x1_sg U40905 ( .A(n21353), .B(n21354), .X(n21186) );
  nand_x1_sg U40906 ( .A(out_L2[16]), .B(n46463), .X(n21354) );
  nand_x1_sg U40907 ( .A(n21535), .B(n21536), .X(n21356) );
  nand_x1_sg U40908 ( .A(out_L2[15]), .B(n21537), .X(n21536) );
  nand_x1_sg U40909 ( .A(n20945), .B(n20946), .X(n20768) );
  inv_x1_sg U40910 ( .A(n20948), .X(n46494) );
  nand_x1_sg U40911 ( .A(n19910), .B(n19911), .X(n19712) );
  inv_x1_sg U40912 ( .A(n19913), .X(n46446) );
  nand_x1_sg U40913 ( .A(n19312), .B(n19313), .X(n6127) );
  inv_x1_sg U40914 ( .A(n19490), .X(n41533) );
  inv_x1_sg U40915 ( .A(n20301), .X(n46452) );
  inv_x1_sg U40916 ( .A(n20288), .X(n41537) );
  inv_x1_sg U40917 ( .A(n6184), .X(n46418) );
  nand_x1_sg U40918 ( .A(n21679), .B(n21680), .X(n21670) );
  nand_x1_sg U40919 ( .A(out_L2[13]), .B(n21681), .X(n21680) );
  nand_x1_sg U40920 ( .A(n20441), .B(n20442), .X(n20310) );
  inv_x1_sg U40921 ( .A(n20443), .X(n46404) );
  inv_x1_sg U40922 ( .A(n19478), .X(n41531) );
  nand_x1_sg U40923 ( .A(n21141), .B(n46373), .X(n20926) );
  nand_x1_sg U40924 ( .A(n20274), .B(n20275), .X(n20100) );
  inv_x1_sg U40925 ( .A(n20277), .X(n46310) );
  nand_x1_sg U40926 ( .A(n19468), .B(n19469), .X(n19296) );
  inv_x1_sg U40927 ( .A(n19471), .X(n46301) );
  nand_x1_sg U40928 ( .A(n21685), .B(n21686), .X(n21658) );
  nand_x1_sg U40929 ( .A(out_L2[11]), .B(n21687), .X(n21686) );
  inv_x1_sg U40930 ( .A(n6275), .X(n46329) );
  nand_x1_sg U40931 ( .A(n21135), .B(n46332), .X(n20919) );
  nand_x1_sg U40932 ( .A(n20910), .B(n20911), .X(n20733) );
  inv_x1_sg U40933 ( .A(n20913), .X(n46274) );
  nand_x1_sg U40934 ( .A(n20420), .B(n46289), .X(n20269) );
  nand_x1_sg U40935 ( .A(n19461), .B(n19462), .X(n19289) );
  inv_x1_sg U40936 ( .A(n19464), .X(n46256) );
  inv_x1_sg U40937 ( .A(n6364), .X(n46238) );
  nand_x1_sg U40938 ( .A(n21691), .B(n21692), .X(n21646) );
  nand_x1_sg U40939 ( .A(out_L2[9]), .B(n21693), .X(n21692) );
  nand_x1_sg U40940 ( .A(n20903), .B(n20904), .X(n20726) );
  inv_x1_sg U40941 ( .A(n20906), .X(n46228) );
  nand_x1_sg U40942 ( .A(n20260), .B(n20261), .X(n20086) );
  inv_x1_sg U40943 ( .A(n20263), .X(n46219) );
  nand_x1_sg U40944 ( .A(n19454), .B(n19455), .X(n19282) );
  inv_x1_sg U40945 ( .A(n19457), .X(n46210) );
  nand_x1_sg U40946 ( .A(n20896), .B(n20897), .X(n20719) );
  inv_x1_sg U40947 ( .A(n20899), .X(n46183) );
  nand_x1_sg U40948 ( .A(n20253), .B(n20254), .X(n20079) );
  inv_x1_sg U40949 ( .A(n20256), .X(n46174) );
  nand_x1_sg U40950 ( .A(n19447), .B(n19448), .X(n19275) );
  inv_x1_sg U40951 ( .A(n19450), .X(n46165) );
  nand_x1_sg U40952 ( .A(n20402), .B(n46153), .X(n20248) );
  nand_x1_sg U40953 ( .A(n19440), .B(n19441), .X(n19268) );
  inv_x1_sg U40954 ( .A(n19443), .X(n46119) );
  nand_x1_sg U40955 ( .A(n21697), .B(n21698), .X(n21634) );
  nand_x1_sg U40956 ( .A(out_L2[7]), .B(n21699), .X(n21698) );
  inv_x1_sg U40957 ( .A(n6453), .X(n46147) );
  nand_x1_sg U40958 ( .A(n20889), .B(n20890), .X(n20712) );
  inv_x1_sg U40959 ( .A(n20892), .X(n46137) );
  nand_x1_sg U40960 ( .A(n20239), .B(n20240), .X(n20065) );
  inv_x1_sg U40961 ( .A(n20242), .X(n46083) );
  nand_x1_sg U40962 ( .A(n19433), .B(n19434), .X(n19261) );
  inv_x1_sg U40963 ( .A(n19436), .X(n46074) );
  nand_x1_sg U40964 ( .A(n20882), .B(n20883), .X(n20705) );
  inv_x1_sg U40965 ( .A(n20885), .X(n46092) );
  nand_x1_sg U40966 ( .A(n20232), .B(n20233), .X(n20058) );
  inv_x1_sg U40967 ( .A(n20235), .X(n46037) );
  nand_x1_sg U40968 ( .A(n19426), .B(n19427), .X(n19254) );
  inv_x1_sg U40969 ( .A(n19429), .X(n46028) );
  nand_x1_sg U40970 ( .A(n21703), .B(n21704), .X(n21622) );
  nand_x1_sg U40971 ( .A(out_L2[5]), .B(n21705), .X(n21704) );
  inv_x1_sg U40972 ( .A(n6542), .X(n46056) );
  nand_x1_sg U40973 ( .A(n21099), .B(n46059), .X(n20877) );
  nand_x1_sg U40974 ( .A(n20225), .B(n20226), .X(n20051) );
  inv_x1_sg U40975 ( .A(n20228), .X(n45992) );
  nand_x1_sg U40976 ( .A(n19419), .B(n19420), .X(n19247) );
  inv_x1_sg U40977 ( .A(n19422), .X(n45983) );
  nand_x1_sg U40978 ( .A(n20868), .B(n20869), .X(n20691) );
  inv_x1_sg U40979 ( .A(n20871), .X(n46001) );
  nand_x1_sg U40980 ( .A(n20218), .B(n20219), .X(n20044) );
  inv_x1_sg U40981 ( .A(n20221), .X(n45947) );
  nand_x1_sg U40982 ( .A(n19412), .B(n19413), .X(n19240) );
  inv_x1_sg U40983 ( .A(n19415), .X(n45938) );
  nand_x1_sg U40984 ( .A(n21709), .B(n21710), .X(n21610) );
  nand_x1_sg U40985 ( .A(out_L2[3]), .B(n21711), .X(n21710) );
  inv_x1_sg U40986 ( .A(n6631), .X(n45965) );
  nand_x1_sg U40987 ( .A(n20861), .B(n20862), .X(n20684) );
  inv_x1_sg U40988 ( .A(n20864), .X(n45956) );
  nand_x1_sg U40989 ( .A(n19407), .B(n19408), .X(n19233) );
  inv_x1_sg U40990 ( .A(n19409), .X(n45890) );
  nand_x1_sg U40991 ( .A(n20213), .B(n20214), .X(n20037) );
  inv_x1_sg U40992 ( .A(n20215), .X(n45900) );
  nand_x1_sg U40993 ( .A(n20856), .B(n20857), .X(n20677) );
  inv_x1_sg U40994 ( .A(n20858), .X(n45910) );
  nand_x1_sg U40995 ( .A(n45879), .B(n20366), .X(n20208) );
  inv_x1_sg U40996 ( .A(n19634), .X(n41534) );
  inv_x1_sg U40997 ( .A(n20028), .X(n41528) );
  inv_x1_sg U40998 ( .A(n19224), .X(n41527) );
  inv_x1_sg U40999 ( .A(n6712), .X(n41530) );
  inv_x1_sg U41000 ( .A(n21268), .X(n45819) );
  inv_x1_sg U41001 ( .A(n20499), .X(n45835) );
  inv_x1_sg U41002 ( .A(n20668), .X(n41529) );
  nand_x1_sg U41003 ( .A(n22840), .B(n22841), .X(n22834) );
  nand_x1_sg U41004 ( .A(n7127), .B(n46881), .X(n7107) );
  nand_x1_sg U41005 ( .A(n46869), .B(n7096), .X(n7086) );
  nand_x1_sg U41006 ( .A(n7145), .B(n7144), .X(n7142) );
  nand_x1_sg U41007 ( .A(n7179), .B(n7178), .X(n7175) );
  nand_x1_sg U41008 ( .A(n7222), .B(n7223), .X(n7220) );
  nand_x1_sg U41009 ( .A(n7227), .B(n46946), .X(n7221) );
  nand_x1_sg U41010 ( .A(n7197), .B(n7196), .X(n7194) );
  nand_x1_sg U41011 ( .A(n7292), .B(n7291), .X(n7266) );
  nand_x1_sg U41012 ( .A(n7266), .B(n46998), .X(n7262) );
  nand_x1_sg U41013 ( .A(n7317), .B(n46995), .X(n7311) );
  nand_x1_sg U41014 ( .A(n7384), .B(n7383), .X(n7352) );
  nand_x1_sg U41015 ( .A(n7352), .B(n47038), .X(n7348) );
  nand_x1_sg U41016 ( .A(n7413), .B(n7412), .X(n7409) );
  nand_x1_sg U41017 ( .A(n7414), .B(n47066), .X(n7403) );
  nand_x1_sg U41018 ( .A(n7484), .B(n7483), .X(n7457) );
  nand_x1_sg U41019 ( .A(n7457), .B(n47088), .X(n7453) );
  nand_x1_sg U41020 ( .A(n7516), .B(n7517), .X(n7043) );
  nand_x1_sg U41021 ( .A(n7041), .B(n47111), .X(n7044) );
  inv_x1_sg U41022 ( .A(n6954), .X(n47009) );
  nand_x1_sg U41023 ( .A(n47162), .B(n7914), .X(n7904) );
  nand_x1_sg U41024 ( .A(n23099), .B(n47142), .X(n23093) );
  nand_x1_sg U41025 ( .A(n7943), .B(n7944), .X(n7942) );
  nand_x1_sg U41026 ( .A(n7963), .B(n7962), .X(n7960) );
  nand_x1_sg U41027 ( .A(n7998), .B(n7997), .X(n7994) );
  nand_x1_sg U41028 ( .A(n8041), .B(n8042), .X(n8039) );
  nand_x1_sg U41029 ( .A(n8046), .B(n47237), .X(n8040) );
  nand_x1_sg U41030 ( .A(n8016), .B(n8015), .X(n8013) );
  nand_x1_sg U41031 ( .A(n8110), .B(n8109), .X(n8085) );
  nand_x1_sg U41032 ( .A(n8087), .B(n8062), .X(n8080) );
  nand_x1_sg U41033 ( .A(n8085), .B(n47287), .X(n8081) );
  nand_x1_sg U41034 ( .A(n8135), .B(n47284), .X(n8129) );
  nand_x1_sg U41035 ( .A(n8202), .B(n8201), .X(n8170) );
  nand_x1_sg U41036 ( .A(n8170), .B(n47325), .X(n8166) );
  nand_x1_sg U41037 ( .A(n8231), .B(n8230), .X(n8227) );
  nand_x1_sg U41038 ( .A(n8232), .B(n47352), .X(n8221) );
  nand_x1_sg U41039 ( .A(n8302), .B(n8301), .X(n8275) );
  nand_x1_sg U41040 ( .A(n8275), .B(n47374), .X(n8271) );
  nand_x1_sg U41041 ( .A(n8334), .B(n8335), .X(n7861) );
  nand_x1_sg U41042 ( .A(n7859), .B(n47397), .X(n7862) );
  inv_x1_sg U41043 ( .A(n7771), .X(n47297) );
  nand_x1_sg U41044 ( .A(n47447), .B(n8732), .X(n8722) );
  nand_x1_sg U41045 ( .A(n23379), .B(n47427), .X(n23373) );
  nand_x1_sg U41046 ( .A(n8761), .B(n8762), .X(n8760) );
  nand_x1_sg U41047 ( .A(n8781), .B(n8780), .X(n8778) );
  nand_x1_sg U41048 ( .A(n8816), .B(n8815), .X(n8812) );
  nand_x1_sg U41049 ( .A(n8859), .B(n8860), .X(n8857) );
  nand_x1_sg U41050 ( .A(n8864), .B(n47522), .X(n8858) );
  nand_x1_sg U41051 ( .A(n8834), .B(n8833), .X(n8831) );
  nand_x1_sg U41052 ( .A(n8928), .B(n8927), .X(n8903) );
  nand_x1_sg U41053 ( .A(n8905), .B(n8880), .X(n8898) );
  nand_x1_sg U41054 ( .A(n8903), .B(n47572), .X(n8899) );
  nand_x1_sg U41055 ( .A(n8953), .B(n47569), .X(n8947) );
  nand_x1_sg U41056 ( .A(n9020), .B(n9019), .X(n8988) );
  nand_x1_sg U41057 ( .A(n8988), .B(n47610), .X(n8984) );
  nand_x1_sg U41058 ( .A(n9049), .B(n9048), .X(n9045) );
  nand_x1_sg U41059 ( .A(n9050), .B(n47637), .X(n9039) );
  nand_x1_sg U41060 ( .A(n9120), .B(n9119), .X(n9093) );
  nand_x1_sg U41061 ( .A(n9093), .B(n47659), .X(n9089) );
  nand_x1_sg U41062 ( .A(n9152), .B(n9153), .X(n8679) );
  nand_x1_sg U41063 ( .A(n8677), .B(n47682), .X(n8680) );
  inv_x1_sg U41064 ( .A(n8589), .X(n47582) );
  nand_x1_sg U41065 ( .A(n47732), .B(n9552), .X(n9542) );
  nand_x1_sg U41066 ( .A(n23658), .B(n47712), .X(n23652) );
  nand_x1_sg U41067 ( .A(n9581), .B(n9582), .X(n9580) );
  nand_x1_sg U41068 ( .A(n9601), .B(n9600), .X(n9598) );
  nand_x1_sg U41069 ( .A(n9636), .B(n9635), .X(n9632) );
  nand_x1_sg U41070 ( .A(n9679), .B(n9680), .X(n9677) );
  nand_x1_sg U41071 ( .A(n9684), .B(n47807), .X(n9678) );
  nand_x1_sg U41072 ( .A(n9654), .B(n9653), .X(n9651) );
  nand_x1_sg U41073 ( .A(n9748), .B(n9747), .X(n9723) );
  nand_x1_sg U41074 ( .A(n9725), .B(n9700), .X(n9718) );
  nand_x1_sg U41075 ( .A(n9723), .B(n47857), .X(n9719) );
  nand_x1_sg U41076 ( .A(n9773), .B(n47854), .X(n9767) );
  nand_x1_sg U41077 ( .A(n9840), .B(n9839), .X(n9808) );
  nand_x1_sg U41078 ( .A(n9808), .B(n47895), .X(n9804) );
  nand_x1_sg U41079 ( .A(n9869), .B(n9868), .X(n9865) );
  nand_x1_sg U41080 ( .A(n9870), .B(n47922), .X(n9859) );
  nand_x1_sg U41081 ( .A(n9940), .B(n9939), .X(n9913) );
  nand_x1_sg U41082 ( .A(n9913), .B(n47944), .X(n9909) );
  nand_x1_sg U41083 ( .A(n9972), .B(n9973), .X(n9499) );
  nand_x1_sg U41084 ( .A(n9497), .B(n47967), .X(n9500) );
  inv_x1_sg U41085 ( .A(n9409), .X(n47867) );
  nand_x1_sg U41086 ( .A(n48017), .B(n10371), .X(n10361) );
  nand_x1_sg U41087 ( .A(n23937), .B(n47997), .X(n23931) );
  nand_x1_sg U41088 ( .A(n10400), .B(n10401), .X(n10399) );
  nand_x1_sg U41089 ( .A(n10420), .B(n10419), .X(n10417) );
  nand_x1_sg U41090 ( .A(n10455), .B(n10454), .X(n10451) );
  nand_x1_sg U41091 ( .A(n10498), .B(n10499), .X(n10496) );
  nand_x1_sg U41092 ( .A(n10503), .B(n48092), .X(n10497) );
  nand_x1_sg U41093 ( .A(n10473), .B(n10472), .X(n10470) );
  nand_x1_sg U41094 ( .A(n10567), .B(n10566), .X(n10542) );
  nand_x1_sg U41095 ( .A(n10544), .B(n10519), .X(n10537) );
  nand_x1_sg U41096 ( .A(n10542), .B(n48142), .X(n10538) );
  nand_x1_sg U41097 ( .A(n10592), .B(n48139), .X(n10586) );
  nand_x1_sg U41098 ( .A(n10659), .B(n10658), .X(n10627) );
  nand_x1_sg U41099 ( .A(n10627), .B(n48180), .X(n10623) );
  nand_x1_sg U41100 ( .A(n10688), .B(n10687), .X(n10684) );
  nand_x1_sg U41101 ( .A(n10689), .B(n48207), .X(n10678) );
  nand_x1_sg U41102 ( .A(n10759), .B(n10758), .X(n10732) );
  nand_x1_sg U41103 ( .A(n10732), .B(n48229), .X(n10728) );
  nand_x1_sg U41104 ( .A(n10791), .B(n10792), .X(n10318) );
  nand_x1_sg U41105 ( .A(n10316), .B(n48252), .X(n10319) );
  inv_x1_sg U41106 ( .A(n10228), .X(n48152) );
  nand_x1_sg U41107 ( .A(n48302), .B(n11190), .X(n11180) );
  nand_x1_sg U41108 ( .A(n24216), .B(n48282), .X(n24210) );
  nand_x1_sg U41109 ( .A(n11219), .B(n11220), .X(n11218) );
  nand_x1_sg U41110 ( .A(n11239), .B(n11238), .X(n11236) );
  nand_x1_sg U41111 ( .A(n11274), .B(n11273), .X(n11270) );
  nand_x1_sg U41112 ( .A(n11317), .B(n11318), .X(n11315) );
  nand_x1_sg U41113 ( .A(n11322), .B(n48377), .X(n11316) );
  nand_x1_sg U41114 ( .A(n11292), .B(n11291), .X(n11289) );
  nand_x1_sg U41115 ( .A(n11386), .B(n11385), .X(n11361) );
  nand_x1_sg U41116 ( .A(n11363), .B(n11338), .X(n11356) );
  nand_x1_sg U41117 ( .A(n11361), .B(n48427), .X(n11357) );
  nand_x1_sg U41118 ( .A(n11411), .B(n48424), .X(n11405) );
  nand_x1_sg U41119 ( .A(n11478), .B(n11477), .X(n11446) );
  nand_x1_sg U41120 ( .A(n11446), .B(n48465), .X(n11442) );
  nand_x1_sg U41121 ( .A(n11507), .B(n11506), .X(n11503) );
  nand_x1_sg U41122 ( .A(n11508), .B(n48492), .X(n11497) );
  nand_x1_sg U41123 ( .A(n11578), .B(n11577), .X(n11551) );
  nand_x1_sg U41124 ( .A(n11551), .B(n48514), .X(n11547) );
  nand_x1_sg U41125 ( .A(n11610), .B(n11611), .X(n11137) );
  nand_x1_sg U41126 ( .A(n11135), .B(n48537), .X(n11138) );
  inv_x1_sg U41127 ( .A(n11047), .X(n48437) );
  nand_x1_sg U41128 ( .A(n48587), .B(n12009), .X(n11999) );
  nand_x1_sg U41129 ( .A(n24495), .B(n48567), .X(n24489) );
  nand_x1_sg U41130 ( .A(n12038), .B(n12039), .X(n12037) );
  nand_x1_sg U41131 ( .A(n12058), .B(n12057), .X(n12055) );
  nand_x1_sg U41132 ( .A(n12093), .B(n12092), .X(n12089) );
  nand_x1_sg U41133 ( .A(n12136), .B(n12137), .X(n12134) );
  nand_x1_sg U41134 ( .A(n12141), .B(n48662), .X(n12135) );
  nand_x1_sg U41135 ( .A(n12111), .B(n12110), .X(n12108) );
  nand_x1_sg U41136 ( .A(n12205), .B(n12204), .X(n12180) );
  nand_x1_sg U41137 ( .A(n12182), .B(n12157), .X(n12175) );
  nand_x1_sg U41138 ( .A(n12180), .B(n48712), .X(n12176) );
  nand_x1_sg U41139 ( .A(n12230), .B(n48709), .X(n12224) );
  nand_x1_sg U41140 ( .A(n12297), .B(n12296), .X(n12265) );
  nand_x1_sg U41141 ( .A(n12265), .B(n48750), .X(n12261) );
  nand_x1_sg U41142 ( .A(n12326), .B(n12325), .X(n12322) );
  nand_x1_sg U41143 ( .A(n12327), .B(n48777), .X(n12316) );
  nand_x1_sg U41144 ( .A(n12397), .B(n12396), .X(n12370) );
  nand_x1_sg U41145 ( .A(n12370), .B(n48799), .X(n12366) );
  nand_x1_sg U41146 ( .A(n12429), .B(n12430), .X(n11956) );
  nand_x1_sg U41147 ( .A(n11954), .B(n48822), .X(n11957) );
  inv_x1_sg U41148 ( .A(n11866), .X(n48722) );
  nand_x1_sg U41149 ( .A(n48873), .B(n12828), .X(n12818) );
  nand_x1_sg U41150 ( .A(n24773), .B(n48852), .X(n24767) );
  nand_x1_sg U41151 ( .A(n12857), .B(n12858), .X(n12856) );
  nand_x1_sg U41152 ( .A(n12877), .B(n12876), .X(n12874) );
  nand_x1_sg U41153 ( .A(n12912), .B(n12911), .X(n12908) );
  nand_x1_sg U41154 ( .A(n12955), .B(n12956), .X(n12953) );
  nand_x1_sg U41155 ( .A(n12960), .B(n48948), .X(n12954) );
  nand_x1_sg U41156 ( .A(n12930), .B(n12929), .X(n12927) );
  nand_x1_sg U41157 ( .A(n13024), .B(n13023), .X(n12999) );
  nand_x1_sg U41158 ( .A(n13001), .B(n12976), .X(n12994) );
  nand_x1_sg U41159 ( .A(n12999), .B(n48998), .X(n12995) );
  nand_x1_sg U41160 ( .A(n13049), .B(n48995), .X(n13043) );
  nand_x1_sg U41161 ( .A(n13116), .B(n13115), .X(n13084) );
  nand_x1_sg U41162 ( .A(n13084), .B(n49036), .X(n13080) );
  nand_x1_sg U41163 ( .A(n13145), .B(n13144), .X(n13141) );
  nand_x1_sg U41164 ( .A(n13146), .B(n49064), .X(n13135) );
  nand_x1_sg U41165 ( .A(n13216), .B(n13215), .X(n13189) );
  nand_x1_sg U41166 ( .A(n13189), .B(n49086), .X(n13185) );
  nand_x1_sg U41167 ( .A(n13248), .B(n13249), .X(n12775) );
  nand_x1_sg U41168 ( .A(n12773), .B(n49109), .X(n12776) );
  inv_x1_sg U41169 ( .A(n12685), .X(n49008) );
  nand_x1_sg U41170 ( .A(n49160), .B(n13647), .X(n13637) );
  nand_x1_sg U41171 ( .A(n25052), .B(n49139), .X(n25046) );
  nand_x1_sg U41172 ( .A(n13676), .B(n13677), .X(n13675) );
  nand_x1_sg U41173 ( .A(n13696), .B(n13695), .X(n13693) );
  nand_x1_sg U41174 ( .A(n13731), .B(n13730), .X(n13727) );
  nand_x1_sg U41175 ( .A(n13774), .B(n13775), .X(n13772) );
  nand_x1_sg U41176 ( .A(n13779), .B(n49235), .X(n13773) );
  nand_x1_sg U41177 ( .A(n13749), .B(n13748), .X(n13746) );
  nand_x1_sg U41178 ( .A(n13843), .B(n13842), .X(n13818) );
  nand_x1_sg U41179 ( .A(n13820), .B(n13795), .X(n13813) );
  nand_x1_sg U41180 ( .A(n13818), .B(n49285), .X(n13814) );
  nand_x1_sg U41181 ( .A(n13868), .B(n49282), .X(n13862) );
  nand_x1_sg U41182 ( .A(n13935), .B(n13934), .X(n13903) );
  nand_x1_sg U41183 ( .A(n13903), .B(n49323), .X(n13899) );
  nand_x1_sg U41184 ( .A(n13964), .B(n13963), .X(n13960) );
  nand_x1_sg U41185 ( .A(n13965), .B(n49350), .X(n13954) );
  nand_x1_sg U41186 ( .A(n14035), .B(n14034), .X(n14008) );
  nand_x1_sg U41187 ( .A(n14008), .B(n49372), .X(n14004) );
  nand_x1_sg U41188 ( .A(n14067), .B(n14068), .X(n13594) );
  nand_x1_sg U41189 ( .A(n13592), .B(n49395), .X(n13595) );
  inv_x1_sg U41190 ( .A(n13504), .X(n49295) );
  nand_x1_sg U41191 ( .A(n14497), .B(n49458), .X(n14477) );
  nand_x1_sg U41192 ( .A(n49446), .B(n14466), .X(n14456) );
  nand_x1_sg U41193 ( .A(n25331), .B(n49425), .X(n25325) );
  nand_x1_sg U41194 ( .A(n14515), .B(n14514), .X(n14512) );
  nand_x1_sg U41195 ( .A(n14550), .B(n14549), .X(n14546) );
  nand_x1_sg U41196 ( .A(n14593), .B(n14594), .X(n14591) );
  nand_x1_sg U41197 ( .A(n14598), .B(n49521), .X(n14592) );
  nand_x1_sg U41198 ( .A(n14568), .B(n14567), .X(n14565) );
  nand_x1_sg U41199 ( .A(n14662), .B(n14661), .X(n14637) );
  nand_x1_sg U41200 ( .A(n14639), .B(n14614), .X(n14632) );
  nand_x1_sg U41201 ( .A(n14637), .B(n49571), .X(n14633) );
  nand_x1_sg U41202 ( .A(n14687), .B(n49568), .X(n14681) );
  nand_x1_sg U41203 ( .A(n14754), .B(n14753), .X(n14722) );
  nand_x1_sg U41204 ( .A(n14722), .B(n49609), .X(n14718) );
  nand_x1_sg U41205 ( .A(n14783), .B(n14782), .X(n14779) );
  nand_x1_sg U41206 ( .A(n14784), .B(n49636), .X(n14773) );
  nand_x1_sg U41207 ( .A(n14854), .B(n14853), .X(n14827) );
  nand_x1_sg U41208 ( .A(n14827), .B(n49658), .X(n14823) );
  nand_x1_sg U41209 ( .A(n14886), .B(n14887), .X(n14413) );
  nand_x1_sg U41210 ( .A(n14411), .B(n49681), .X(n14414) );
  inv_x1_sg U41211 ( .A(n14323), .X(n49581) );
  nand_x1_sg U41212 ( .A(n15316), .B(n49743), .X(n15296) );
  nand_x1_sg U41213 ( .A(n49731), .B(n15285), .X(n15275) );
  nand_x1_sg U41214 ( .A(n25610), .B(n49711), .X(n25604) );
  nand_x1_sg U41215 ( .A(n15334), .B(n15333), .X(n15331) );
  nand_x1_sg U41216 ( .A(n15369), .B(n15368), .X(n15365) );
  nand_x1_sg U41217 ( .A(n15412), .B(n15413), .X(n15410) );
  nand_x1_sg U41218 ( .A(n15417), .B(n49807), .X(n15411) );
  nand_x1_sg U41219 ( .A(n15387), .B(n15386), .X(n15384) );
  nand_x1_sg U41220 ( .A(n15481), .B(n15480), .X(n15456) );
  nand_x1_sg U41221 ( .A(n15458), .B(n15433), .X(n15451) );
  nand_x1_sg U41222 ( .A(n15456), .B(n49857), .X(n15452) );
  nand_x1_sg U41223 ( .A(n15506), .B(n49854), .X(n15500) );
  nand_x1_sg U41224 ( .A(n15573), .B(n15572), .X(n15541) );
  nand_x1_sg U41225 ( .A(n15541), .B(n49895), .X(n15537) );
  nand_x1_sg U41226 ( .A(n15602), .B(n15601), .X(n15598) );
  nand_x1_sg U41227 ( .A(n15603), .B(n49922), .X(n15592) );
  nand_x1_sg U41228 ( .A(n15673), .B(n15672), .X(n15646) );
  nand_x1_sg U41229 ( .A(n15646), .B(n49944), .X(n15642) );
  nand_x1_sg U41230 ( .A(n15705), .B(n15706), .X(n15232) );
  nand_x1_sg U41231 ( .A(n15230), .B(n49967), .X(n15233) );
  inv_x1_sg U41232 ( .A(n15142), .X(n49867) );
  nand_x1_sg U41233 ( .A(n16135), .B(n50030), .X(n16115) );
  nand_x1_sg U41234 ( .A(n50018), .B(n16104), .X(n16094) );
  nand_x1_sg U41235 ( .A(n25887), .B(n49997), .X(n25881) );
  nand_x1_sg U41236 ( .A(n16153), .B(n16152), .X(n16150) );
  nand_x1_sg U41237 ( .A(n16188), .B(n16187), .X(n16184) );
  nand_x1_sg U41238 ( .A(n16231), .B(n16232), .X(n16229) );
  nand_x1_sg U41239 ( .A(n16236), .B(n50093), .X(n16230) );
  nand_x1_sg U41240 ( .A(n16206), .B(n16205), .X(n16203) );
  nand_x1_sg U41241 ( .A(n16300), .B(n16299), .X(n16275) );
  nand_x1_sg U41242 ( .A(n16277), .B(n16252), .X(n16270) );
  nand_x1_sg U41243 ( .A(n16275), .B(n50143), .X(n16271) );
  nand_x1_sg U41244 ( .A(n16325), .B(n50140), .X(n16319) );
  nand_x1_sg U41245 ( .A(n16392), .B(n16391), .X(n16360) );
  nand_x1_sg U41246 ( .A(n16360), .B(n50181), .X(n16356) );
  nand_x1_sg U41247 ( .A(n16421), .B(n16420), .X(n16417) );
  nand_x1_sg U41248 ( .A(n16422), .B(n50208), .X(n16411) );
  nand_x1_sg U41249 ( .A(n16492), .B(n16491), .X(n16465) );
  nand_x1_sg U41250 ( .A(n16465), .B(n50230), .X(n16461) );
  nand_x1_sg U41251 ( .A(n16524), .B(n16525), .X(n16051) );
  nand_x1_sg U41252 ( .A(n16049), .B(n50253), .X(n16052) );
  inv_x1_sg U41253 ( .A(n15961), .X(n50153) );
  nand_x1_sg U41254 ( .A(n16952), .B(n50315), .X(n16932) );
  nand_x1_sg U41255 ( .A(n50303), .B(n16921), .X(n16912) );
  nand_x1_sg U41256 ( .A(n16970), .B(n16969), .X(n16967) );
  nand_x1_sg U41257 ( .A(n17004), .B(n17003), .X(n17000) );
  nand_x1_sg U41258 ( .A(n17047), .B(n17048), .X(n17045) );
  nand_x1_sg U41259 ( .A(n17052), .B(n50378), .X(n17046) );
  nand_x1_sg U41260 ( .A(n17022), .B(n17021), .X(n17019) );
  nand_x1_sg U41261 ( .A(n17117), .B(n17116), .X(n17091) );
  nand_x1_sg U41262 ( .A(n17091), .B(n50428), .X(n17087) );
  nand_x1_sg U41263 ( .A(n17142), .B(n50425), .X(n17136) );
  nand_x1_sg U41264 ( .A(n17209), .B(n17208), .X(n17177) );
  nand_x1_sg U41265 ( .A(n17177), .B(n50466), .X(n17173) );
  nand_x1_sg U41266 ( .A(n17238), .B(n17237), .X(n17234) );
  nand_x1_sg U41267 ( .A(n17239), .B(n50493), .X(n17228) );
  nand_x1_sg U41268 ( .A(n17309), .B(n17308), .X(n17282) );
  nand_x1_sg U41269 ( .A(n17282), .B(n50515), .X(n17278) );
  nand_x1_sg U41270 ( .A(n17341), .B(n17342), .X(n16870) );
  nand_x1_sg U41271 ( .A(n16868), .B(n50538), .X(n16871) );
  inv_x1_sg U41272 ( .A(n16778), .X(n50438) );
  nand_x1_sg U41273 ( .A(n17773), .B(n50604), .X(n17753) );
  nand_x1_sg U41274 ( .A(n50592), .B(n17742), .X(n17732) );
  nand_x1_sg U41275 ( .A(n26447), .B(n50572), .X(n26441) );
  nand_x1_sg U41276 ( .A(n17791), .B(n17790), .X(n17788) );
  nand_x1_sg U41277 ( .A(n17826), .B(n17825), .X(n17822) );
  nand_x1_sg U41278 ( .A(n17869), .B(n17870), .X(n17867) );
  nand_x1_sg U41279 ( .A(n17874), .B(n50667), .X(n17868) );
  nand_x1_sg U41280 ( .A(n17844), .B(n17843), .X(n17841) );
  nand_x1_sg U41281 ( .A(n17938), .B(n17937), .X(n17913) );
  nand_x1_sg U41282 ( .A(n17915), .B(n17890), .X(n17908) );
  nand_x1_sg U41283 ( .A(n17913), .B(n50717), .X(n17909) );
  nand_x1_sg U41284 ( .A(n17963), .B(n50714), .X(n17957) );
  nand_x1_sg U41285 ( .A(n18030), .B(n18029), .X(n17998) );
  nand_x1_sg U41286 ( .A(n17998), .B(n50755), .X(n17994) );
  nand_x1_sg U41287 ( .A(n18059), .B(n18058), .X(n18055) );
  nand_x1_sg U41288 ( .A(n18060), .B(n50782), .X(n18049) );
  nand_x1_sg U41289 ( .A(n18130), .B(n18129), .X(n18103) );
  nand_x1_sg U41290 ( .A(n18103), .B(n50804), .X(n18099) );
  nand_x1_sg U41291 ( .A(n18162), .B(n18163), .X(n17689) );
  nand_x1_sg U41292 ( .A(n17687), .B(n50827), .X(n17690) );
  inv_x1_sg U41293 ( .A(n17599), .X(n50727) );
  nand_x1_sg U41294 ( .A(n18594), .B(n50891), .X(n18574) );
  nand_x1_sg U41295 ( .A(n50879), .B(n18563), .X(n18553) );
  nand_x1_sg U41296 ( .A(n26725), .B(n50858), .X(n26719) );
  nand_x1_sg U41297 ( .A(n18612), .B(n18611), .X(n18609) );
  nand_x1_sg U41298 ( .A(n18647), .B(n18646), .X(n18643) );
  nand_x1_sg U41299 ( .A(n18690), .B(n18691), .X(n18688) );
  nand_x1_sg U41300 ( .A(n18695), .B(n50954), .X(n18689) );
  nand_x1_sg U41301 ( .A(n18665), .B(n18664), .X(n18662) );
  nand_x1_sg U41302 ( .A(n18759), .B(n18758), .X(n18734) );
  nand_x1_sg U41303 ( .A(n18736), .B(n18711), .X(n18729) );
  nand_x1_sg U41304 ( .A(n18734), .B(n51004), .X(n18730) );
  nand_x1_sg U41305 ( .A(n18784), .B(n51001), .X(n18778) );
  nand_x1_sg U41306 ( .A(n18851), .B(n18850), .X(n18819) );
  nand_x1_sg U41307 ( .A(n18819), .B(n51042), .X(n18815) );
  nand_x1_sg U41308 ( .A(n18880), .B(n18879), .X(n18876) );
  nand_x1_sg U41309 ( .A(n18881), .B(n51069), .X(n18870) );
  nand_x1_sg U41310 ( .A(n18951), .B(n18950), .X(n18924) );
  nand_x1_sg U41311 ( .A(n18924), .B(n51091), .X(n18920) );
  nand_x1_sg U41312 ( .A(n18983), .B(n18984), .X(n18510) );
  nand_x1_sg U41313 ( .A(n18508), .B(n51114), .X(n18511) );
  inv_x1_sg U41314 ( .A(n18420), .X(n51014) );
  nand_x1_sg U41315 ( .A(n5170), .B(n26882), .X(n26881) );
  nand_x1_sg U41316 ( .A(n5284), .B(n26839), .X(n26838) );
  nand_x1_sg U41317 ( .A(n26820), .B(n45790), .X(n26771) );
  nand_x1_sg U41318 ( .A(n45793), .B(n26811), .X(n26770) );
  nand_x1_sg U41319 ( .A(n45791), .B(n26817), .X(n26765) );
  nand_x1_sg U41320 ( .A(n45794), .B(n26808), .X(n26766) );
  nand_x1_sg U41321 ( .A(n45792), .B(n26814), .X(n26777) );
  inv_x1_sg U41322 ( .A(n28556), .X(n45737) );
  nand_x1_sg U41323 ( .A(n28752), .B(n28753), .X(n28556) );
  inv_x1_sg U41324 ( .A(n26836), .X(n45734) );
  nand_x1_sg U41325 ( .A(n27090), .B(n27091), .X(n26836) );
  inv_x1_sg U41326 ( .A(n21762), .X(n45726) );
  nand_x1_sg U41327 ( .A(n26900), .B(n26901), .X(n21762) );
  inv_x1_sg U41328 ( .A(n26893), .X(n45727) );
  nand_x1_sg U41329 ( .A(n27139), .B(n27140), .X(n26893) );
  nand_x1_sg U41330 ( .A(n28738), .B(n28739), .X(n28540) );
  nand_x1_sg U41331 ( .A(out_L1[17]), .B(n28740), .X(n28739) );
  nand_x1_sg U41332 ( .A(n5400), .B(n45696), .X(n28740) );
  inv_x1_sg U41333 ( .A(n28563), .X(n45736) );
  nand_x1_sg U41334 ( .A(n28758), .B(n28759), .X(n28563) );
  nand_x1_sg U41335 ( .A(n27076), .B(n45752), .X(n26851) );
  nand_x1_sg U41336 ( .A(n27070), .B(n45756), .X(n21731) );
  nand_x1_sg U41337 ( .A(n27061), .B(n45762), .X(n21732) );
  nand_x1_sg U41338 ( .A(n27073), .B(n27074), .X(n21736) );
  inv_x1_sg U41339 ( .A(n27075), .X(n45711) );
  nand_x1_sg U41340 ( .A(n27064), .B(n45760), .X(n21735) );
  nand_x1_sg U41341 ( .A(n27067), .B(n45758), .X(n21741) );
  nand_x1_sg U41342 ( .A(n27058), .B(n45764), .X(n21742) );
  inv_x1_sg U41343 ( .A(n28549), .X(n45738) );
  nand_x1_sg U41344 ( .A(n28746), .B(n28747), .X(n28549) );
  inv_x1_sg U41345 ( .A(n27087), .X(n45735) );
  nand_x1_sg U41346 ( .A(n28570), .B(n28571), .X(n27087) );
  inv_x1_sg U41347 ( .A(n28755), .X(n45694) );
  nand_x1_sg U41348 ( .A(n28931), .B(n28932), .X(n28755) );
  inv_x1_sg U41349 ( .A(n27093), .X(n45691) );
  nand_x1_sg U41350 ( .A(n27320), .B(n27321), .X(n27093) );
  inv_x1_sg U41351 ( .A(n27054), .X(n45684) );
  nand_x1_sg U41352 ( .A(n27142), .B(n27143), .X(n27054) );
  inv_x1_sg U41353 ( .A(n21809), .X(n45683) );
  nand_x1_sg U41354 ( .A(n26903), .B(n26904), .X(n21809) );
  inv_x1_sg U41355 ( .A(n28725), .X(n45693) );
  nand_x1_sg U41356 ( .A(n28761), .B(n28762), .X(n28725) );
  nand_x1_sg U41357 ( .A(n27306), .B(n45709), .X(n27105) );
  nand_x1_sg U41358 ( .A(n27300), .B(n45713), .X(n21778) );
  nand_x1_sg U41359 ( .A(n27291), .B(n45719), .X(n21779) );
  nand_x1_sg U41360 ( .A(n27303), .B(n27304), .X(n21783) );
  inv_x1_sg U41361 ( .A(n27305), .X(n45668) );
  nand_x1_sg U41362 ( .A(n27294), .B(n45717), .X(n21782) );
  nand_x1_sg U41363 ( .A(n27297), .B(n45715), .X(n21788) );
  nand_x1_sg U41364 ( .A(n27288), .B(n45721), .X(n21789) );
  inv_x1_sg U41365 ( .A(n28749), .X(n45695) );
  nand_x1_sg U41366 ( .A(n28925), .B(n28926), .X(n28749) );
  inv_x1_sg U41367 ( .A(n27317), .X(n45692) );
  nand_x1_sg U41368 ( .A(n28573), .B(n28574), .X(n27317) );
  inv_x1_sg U41369 ( .A(n27323), .X(n45647) );
  nand_x1_sg U41370 ( .A(n27533), .B(n27534), .X(n27323) );
  inv_x1_sg U41371 ( .A(n28907), .X(n45650) );
  nand_x1_sg U41372 ( .A(n28934), .B(n28935), .X(n28907) );
  inv_x1_sg U41373 ( .A(n21856), .X(n45639) );
  nand_x1_sg U41374 ( .A(n26906), .B(n26907), .X(n21856) );
  inv_x1_sg U41375 ( .A(n27048), .X(n45640) );
  nand_x1_sg U41376 ( .A(n27145), .B(n27146), .X(n27048) );
  inv_x1_sg U41377 ( .A(n28719), .X(n45649) );
  nand_x1_sg U41378 ( .A(n28764), .B(n28765), .X(n28719) );
  nand_x1_sg U41379 ( .A(n27519), .B(n45665), .X(n27335) );
  nand_x1_sg U41380 ( .A(n27513), .B(n45670), .X(n21825) );
  nand_x1_sg U41381 ( .A(n27504), .B(n45676), .X(n21826) );
  nand_x1_sg U41382 ( .A(n27516), .B(n27517), .X(n21830) );
  inv_x1_sg U41383 ( .A(n27518), .X(n45624) );
  nand_x1_sg U41384 ( .A(n27507), .B(n45674), .X(n21829) );
  nand_x1_sg U41385 ( .A(n27510), .B(n45672), .X(n21835) );
  nand_x1_sg U41386 ( .A(n27282), .B(n45678), .X(n21836) );
  inv_x1_sg U41387 ( .A(n27530), .X(n45648) );
  nand_x1_sg U41388 ( .A(n28576), .B(n28577), .X(n27530) );
  inv_x1_sg U41389 ( .A(n28928), .X(n45651) );
  nand_x1_sg U41390 ( .A(n29094), .B(n29095), .X(n28928) );
  inv_x1_sg U41391 ( .A(n28901), .X(n45606) );
  nand_x1_sg U41392 ( .A(n28937), .B(n28938), .X(n28901) );
  inv_x1_sg U41393 ( .A(n27536), .X(n45603) );
  nand_x1_sg U41394 ( .A(n27727), .B(n27728), .X(n27536) );
  inv_x1_sg U41395 ( .A(n21902), .X(n45595) );
  nand_x1_sg U41396 ( .A(n26909), .B(n26910), .X(n21902) );
  inv_x1_sg U41397 ( .A(n27042), .X(n45596) );
  nand_x1_sg U41398 ( .A(n27148), .B(n27149), .X(n27042) );
  inv_x1_sg U41399 ( .A(n28713), .X(n45605) );
  nand_x1_sg U41400 ( .A(n28767), .B(n28768), .X(n28713) );
  nand_x1_sg U41401 ( .A(n27713), .B(n45621), .X(n27548) );
  nand_x1_sg U41402 ( .A(n27707), .B(n45626), .X(n21872) );
  nand_x1_sg U41403 ( .A(n27498), .B(n45632), .X(n21873) );
  nand_x1_sg U41404 ( .A(n27710), .B(n27711), .X(n21877) );
  inv_x1_sg U41405 ( .A(n27712), .X(n45580) );
  nand_x1_sg U41406 ( .A(n27701), .B(n45630), .X(n21876) );
  nand_x1_sg U41407 ( .A(n27704), .B(n45628), .X(n21882) );
  nand_x1_sg U41408 ( .A(n27276), .B(n45634), .X(n21883) );
  nand_x1_sg U41409 ( .A(n29227), .B(n29228), .X(n29089) );
  nand_x1_sg U41410 ( .A(out_L1[14]), .B(n45519), .X(n29228) );
  inv_x1_sg U41411 ( .A(n29079), .X(n45607) );
  nand_x1_sg U41412 ( .A(n29097), .B(n29098), .X(n29079) );
  inv_x1_sg U41413 ( .A(n27724), .X(n45604) );
  nand_x1_sg U41414 ( .A(n28579), .B(n28580), .X(n27724) );
  inv_x1_sg U41415 ( .A(n28895), .X(n45561) );
  nand_x1_sg U41416 ( .A(n28940), .B(n28941), .X(n28895) );
  inv_x1_sg U41417 ( .A(n27730), .X(n45558) );
  nand_x1_sg U41418 ( .A(n27904), .B(n27905), .X(n27730) );
  inv_x1_sg U41419 ( .A(n27036), .X(n45551) );
  nand_x1_sg U41420 ( .A(n27151), .B(n27152), .X(n27036) );
  inv_x1_sg U41421 ( .A(n21949), .X(n45550) );
  nand_x1_sg U41422 ( .A(n26912), .B(n26913), .X(n21949) );
  inv_x1_sg U41423 ( .A(n28707), .X(n45560) );
  nand_x1_sg U41424 ( .A(n28770), .B(n28771), .X(n28707) );
  nand_x1_sg U41425 ( .A(n27890), .B(n45577), .X(n27742) );
  nand_x1_sg U41426 ( .A(n27884), .B(n45582), .X(n21918) );
  nand_x1_sg U41427 ( .A(n27492), .B(n45588), .X(n21919) );
  nand_x1_sg U41428 ( .A(n27887), .B(n27888), .X(n21923) );
  inv_x1_sg U41429 ( .A(n27889), .X(n45535) );
  nand_x1_sg U41430 ( .A(n27695), .B(n45586), .X(n21922) );
  nand_x1_sg U41431 ( .A(n27881), .B(n45584), .X(n21928) );
  nand_x1_sg U41432 ( .A(n27270), .B(n45590), .X(n21929) );
  inv_x1_sg U41433 ( .A(n29072), .X(n45562) );
  nand_x1_sg U41434 ( .A(n29100), .B(n29101), .X(n29072) );
  inv_x1_sg U41435 ( .A(n27901), .X(n45559) );
  nand_x1_sg U41436 ( .A(n28582), .B(n28583), .X(n27901) );
  inv_x1_sg U41437 ( .A(n28889), .X(n45517) );
  nand_x1_sg U41438 ( .A(n28943), .B(n28944), .X(n28889) );
  inv_x1_sg U41439 ( .A(n27907), .X(n45514) );
  nand_x1_sg U41440 ( .A(n28066), .B(n28067), .X(n27907) );
  inv_x1_sg U41441 ( .A(n21995), .X(n45506) );
  nand_x1_sg U41442 ( .A(n26915), .B(n26916), .X(n21995) );
  inv_x1_sg U41443 ( .A(n27030), .X(n45507) );
  nand_x1_sg U41444 ( .A(n27154), .B(n27155), .X(n27030) );
  inv_x1_sg U41445 ( .A(n28701), .X(n45516) );
  nand_x1_sg U41446 ( .A(n28773), .B(n28774), .X(n28701) );
  nand_x1_sg U41447 ( .A(n28052), .B(n45532), .X(n27919) );
  nand_x1_sg U41448 ( .A(n28049), .B(n28050), .X(n21970) );
  inv_x1_sg U41449 ( .A(n28051), .X(n45491) );
  nand_x1_sg U41450 ( .A(n27689), .B(n45541), .X(n21969) );
  nand_x1_sg U41451 ( .A(n28046), .B(n45537), .X(n21965) );
  nand_x1_sg U41452 ( .A(n27486), .B(n45543), .X(n21966) );
  nand_x1_sg U41453 ( .A(n27875), .B(n45539), .X(n21975) );
  nand_x1_sg U41454 ( .A(n27264), .B(n45545), .X(n21976) );
  nand_x1_sg U41455 ( .A(n29233), .B(n29234), .X(n29214) );
  nand_x1_sg U41456 ( .A(out_L1[12]), .B(n45430), .X(n29234) );
  inv_x1_sg U41457 ( .A(n29066), .X(n45518) );
  nand_x1_sg U41458 ( .A(n29103), .B(n29104), .X(n29066) );
  inv_x1_sg U41459 ( .A(n28063), .X(n45515) );
  nand_x1_sg U41460 ( .A(n28585), .B(n28586), .X(n28063) );
  inv_x1_sg U41461 ( .A(n28883), .X(n45472) );
  nand_x1_sg U41462 ( .A(n28946), .B(n28947), .X(n28883) );
  inv_x1_sg U41463 ( .A(n28069), .X(n45469) );
  nand_x1_sg U41464 ( .A(n28201), .B(n28202), .X(n28069) );
  inv_x1_sg U41465 ( .A(n22042), .X(n45458) );
  nand_x1_sg U41466 ( .A(n26918), .B(n26919), .X(n22042) );
  inv_x1_sg U41467 ( .A(n27024), .X(n45459) );
  nand_x1_sg U41468 ( .A(n27157), .B(n27158), .X(n27024) );
  inv_x1_sg U41469 ( .A(n28695), .X(n45471) );
  nand_x1_sg U41470 ( .A(n28776), .B(n28777), .X(n28695) );
  nand_x1_sg U41471 ( .A(n28187), .B(n45488), .X(n28081) );
  nand_x1_sg U41472 ( .A(n28040), .B(n45493), .X(n22011) );
  nand_x1_sg U41473 ( .A(n27480), .B(n45499), .X(n22012) );
  nand_x1_sg U41474 ( .A(n28184), .B(n28185), .X(n22016) );
  inv_x1_sg U41475 ( .A(n28186), .X(n45467) );
  nand_x1_sg U41476 ( .A(n27683), .B(n45497), .X(n22015) );
  nand_x1_sg U41477 ( .A(n27869), .B(n45495), .X(n22021) );
  nand_x1_sg U41478 ( .A(n27258), .B(n45501), .X(n22022) );
  inv_x1_sg U41479 ( .A(n29059), .X(n45473) );
  nand_x1_sg U41480 ( .A(n29106), .B(n29107), .X(n29059) );
  inv_x1_sg U41481 ( .A(n28198), .X(n45470) );
  nand_x1_sg U41482 ( .A(n28588), .B(n28589), .X(n28198) );
  inv_x1_sg U41483 ( .A(n28877), .X(n45428) );
  nand_x1_sg U41484 ( .A(n28949), .B(n28950), .X(n28877) );
  inv_x1_sg U41485 ( .A(n28204), .X(n45425) );
  nand_x1_sg U41486 ( .A(n28330), .B(n28331), .X(n28204) );
  inv_x1_sg U41487 ( .A(n27018), .X(n45415) );
  nand_x1_sg U41488 ( .A(n27160), .B(n27161), .X(n27018) );
  inv_x1_sg U41489 ( .A(n22088), .X(n45414) );
  nand_x1_sg U41490 ( .A(n26921), .B(n26922), .X(n22088) );
  inv_x1_sg U41491 ( .A(n28689), .X(n45427) );
  nand_x1_sg U41492 ( .A(n28779), .B(n28780), .X(n28689) );
  nand_x1_sg U41493 ( .A(n28316), .B(n45443), .X(n28180) );
  nand_x1_sg U41494 ( .A(n28034), .B(n45445), .X(n22058) );
  nand_x1_sg U41495 ( .A(n27474), .B(n45451), .X(n22059) );
  nand_x1_sg U41496 ( .A(n28178), .B(n28179), .X(n22063) );
  inv_x1_sg U41497 ( .A(n28181), .X(n45423) );
  nand_x1_sg U41498 ( .A(n27677), .B(n45449), .X(n22062) );
  nand_x1_sg U41499 ( .A(n27863), .B(n45447), .X(n22068) );
  nand_x1_sg U41500 ( .A(n27252), .B(n45453), .X(n22069) );
  nand_x1_sg U41501 ( .A(n29239), .B(n29240), .X(n29202) );
  nand_x1_sg U41502 ( .A(out_L1[10]), .B(n45339), .X(n29240) );
  inv_x1_sg U41503 ( .A(n29053), .X(n45429) );
  nand_x1_sg U41504 ( .A(n29109), .B(n29110), .X(n29053) );
  inv_x1_sg U41505 ( .A(n28327), .X(n45426) );
  nand_x1_sg U41506 ( .A(n28591), .B(n28592), .X(n28327) );
  inv_x1_sg U41507 ( .A(n28333), .X(n45379) );
  nand_x1_sg U41508 ( .A(n28434), .B(n28435), .X(n28333) );
  inv_x1_sg U41509 ( .A(n28871), .X(n45382) );
  nand_x1_sg U41510 ( .A(n28952), .B(n28953), .X(n28871) );
  inv_x1_sg U41511 ( .A(n27012), .X(n45369) );
  nand_x1_sg U41512 ( .A(n27163), .B(n27164), .X(n27012) );
  inv_x1_sg U41513 ( .A(n22136), .X(n45368) );
  nand_x1_sg U41514 ( .A(n26924), .B(n26925), .X(n22136) );
  inv_x1_sg U41515 ( .A(n28683), .X(n45381) );
  nand_x1_sg U41516 ( .A(n28782), .B(n28783), .X(n28683) );
  inv_x1_sg U41517 ( .A(n22126), .X(n45397) );
  nand_x1_sg U41518 ( .A(n28173), .B(n28174), .X(n22109) );
  inv_x1_sg U41519 ( .A(n28175), .X(n45377) );
  nand_x1_sg U41520 ( .A(n27671), .B(n45405), .X(n22108) );
  nand_x1_sg U41521 ( .A(n28028), .B(n45401), .X(n22104) );
  nand_x1_sg U41522 ( .A(n27468), .B(n45407), .X(n22105) );
  nand_x1_sg U41523 ( .A(n27857), .B(n45403), .X(n22114) );
  nand_x1_sg U41524 ( .A(n27246), .B(n45409), .X(n22115) );
  inv_x1_sg U41525 ( .A(n28431), .X(n45380) );
  nand_x1_sg U41526 ( .A(n28594), .B(n28595), .X(n28431) );
  inv_x1_sg U41527 ( .A(n29046), .X(n45383) );
  nand_x1_sg U41528 ( .A(n29112), .B(n29113), .X(n29046) );
  inv_x1_sg U41529 ( .A(n28865), .X(n45337) );
  nand_x1_sg U41530 ( .A(n28955), .B(n28956), .X(n28865) );
  inv_x1_sg U41531 ( .A(n28422), .X(n45334) );
  nand_x1_sg U41532 ( .A(n28437), .B(n28438), .X(n28422) );
  inv_x1_sg U41533 ( .A(n22183), .X(n45323) );
  nand_x1_sg U41534 ( .A(n26927), .B(n26928), .X(n22183) );
  inv_x1_sg U41535 ( .A(n27006), .X(n45324) );
  nand_x1_sg U41536 ( .A(n27166), .B(n27167), .X(n27006) );
  inv_x1_sg U41537 ( .A(n28677), .X(n45336) );
  nand_x1_sg U41538 ( .A(n28785), .B(n28786), .X(n28677) );
  inv_x1_sg U41539 ( .A(n22173), .X(n45351) );
  nand_x1_sg U41540 ( .A(n28168), .B(n28169), .X(n22157) );
  inv_x1_sg U41541 ( .A(n28170), .X(n45332) );
  nand_x1_sg U41542 ( .A(n27665), .B(n45359), .X(n22156) );
  nand_x1_sg U41543 ( .A(n28022), .B(n45355), .X(n22152) );
  nand_x1_sg U41544 ( .A(n27462), .B(n45361), .X(n22153) );
  nand_x1_sg U41545 ( .A(n27851), .B(n45357), .X(n22162) );
  nand_x1_sg U41546 ( .A(n27240), .B(n45363), .X(n22163) );
  nand_x1_sg U41547 ( .A(n29245), .B(n29246), .X(n29190) );
  nand_x1_sg U41548 ( .A(out_L1[8]), .B(n29247), .X(n29246) );
  nand_x1_sg U41549 ( .A(n5409), .B(n45249), .X(n29247) );
  inv_x1_sg U41550 ( .A(n29040), .X(n45338) );
  nand_x1_sg U41551 ( .A(n29115), .B(n29116), .X(n29040) );
  inv_x1_sg U41552 ( .A(n28516), .X(n45335) );
  nand_x1_sg U41553 ( .A(n28597), .B(n28598), .X(n28516) );
  inv_x1_sg U41554 ( .A(n28859), .X(n45292) );
  nand_x1_sg U41555 ( .A(n28958), .B(n28959), .X(n28859) );
  inv_x1_sg U41556 ( .A(n28416), .X(n45289) );
  nand_x1_sg U41557 ( .A(n28440), .B(n28441), .X(n28416) );
  inv_x1_sg U41558 ( .A(n27000), .X(n45279) );
  nand_x1_sg U41559 ( .A(n27169), .B(n27170), .X(n27000) );
  inv_x1_sg U41560 ( .A(n22231), .X(n45278) );
  nand_x1_sg U41561 ( .A(n26930), .B(n26931), .X(n22231) );
  inv_x1_sg U41562 ( .A(n28671), .X(n45291) );
  nand_x1_sg U41563 ( .A(n28788), .B(n28789), .X(n28671) );
  inv_x1_sg U41564 ( .A(n22221), .X(n45306) );
  nand_x1_sg U41565 ( .A(n28163), .B(n28164), .X(n22204) );
  inv_x1_sg U41566 ( .A(n28165), .X(n45287) );
  nand_x1_sg U41567 ( .A(n27659), .B(n45314), .X(n22203) );
  nand_x1_sg U41568 ( .A(n28016), .B(n45310), .X(n22199) );
  nand_x1_sg U41569 ( .A(n27456), .B(n45316), .X(n22200) );
  nand_x1_sg U41570 ( .A(n27845), .B(n45312), .X(n22209) );
  nand_x1_sg U41571 ( .A(n27234), .B(n45318), .X(n22210) );
  inv_x1_sg U41572 ( .A(n29033), .X(n45293) );
  nand_x1_sg U41573 ( .A(n29118), .B(n29119), .X(n29033) );
  inv_x1_sg U41574 ( .A(n28510), .X(n45290) );
  nand_x1_sg U41575 ( .A(n28600), .B(n28601), .X(n28510) );
  inv_x1_sg U41576 ( .A(n28410), .X(n45244) );
  nand_x1_sg U41577 ( .A(n28443), .B(n28444), .X(n28410) );
  inv_x1_sg U41578 ( .A(n28853), .X(n45247) );
  nand_x1_sg U41579 ( .A(n28961), .B(n28962), .X(n28853) );
  inv_x1_sg U41580 ( .A(n22278), .X(n45233) );
  nand_x1_sg U41581 ( .A(n26933), .B(n26934), .X(n22278) );
  inv_x1_sg U41582 ( .A(n26994), .X(n45234) );
  nand_x1_sg U41583 ( .A(n27172), .B(n27173), .X(n26994) );
  inv_x1_sg U41584 ( .A(n28665), .X(n45246) );
  nand_x1_sg U41585 ( .A(n28791), .B(n28792), .X(n28665) );
  inv_x1_sg U41586 ( .A(n22268), .X(n45261) );
  nand_x1_sg U41587 ( .A(n28010), .B(n45265), .X(n22247) );
  nand_x1_sg U41588 ( .A(n27450), .B(n45271), .X(n22248) );
  nand_x1_sg U41589 ( .A(n28158), .B(n28159), .X(n22252) );
  inv_x1_sg U41590 ( .A(n28160), .X(n45242) );
  nand_x1_sg U41591 ( .A(n27653), .B(n45269), .X(n22251) );
  nand_x1_sg U41592 ( .A(n27839), .B(n45267), .X(n22257) );
  nand_x1_sg U41593 ( .A(n27228), .B(n45273), .X(n22258) );
  inv_x1_sg U41594 ( .A(n28504), .X(n45245) );
  nand_x1_sg U41595 ( .A(n28603), .B(n28604), .X(n28504) );
  nand_x1_sg U41596 ( .A(n29251), .B(n29252), .X(n29178) );
  nand_x1_sg U41597 ( .A(out_L1[6]), .B(n29253), .X(n29252) );
  nand_x1_sg U41598 ( .A(n5411), .B(n45158), .X(n29253) );
  inv_x1_sg U41599 ( .A(n29027), .X(n45248) );
  nand_x1_sg U41600 ( .A(n29121), .B(n29122), .X(n29027) );
  inv_x1_sg U41601 ( .A(n28847), .X(n45201) );
  nand_x1_sg U41602 ( .A(n28964), .B(n28965), .X(n28847) );
  inv_x1_sg U41603 ( .A(n28404), .X(n45198) );
  nand_x1_sg U41604 ( .A(n28446), .B(n28447), .X(n28404) );
  inv_x1_sg U41605 ( .A(n26988), .X(n45188) );
  nand_x1_sg U41606 ( .A(n27175), .B(n27176), .X(n26988) );
  inv_x1_sg U41607 ( .A(n22326), .X(n45187) );
  nand_x1_sg U41608 ( .A(n26936), .B(n26937), .X(n22326) );
  nor_x4_sg U41609 ( .A(n42116), .B(out_L1[6]), .X(n29175) );
  inv_x1_sg U41610 ( .A(n28659), .X(n45200) );
  nand_x1_sg U41611 ( .A(n28794), .B(n28795), .X(n28659) );
  inv_x1_sg U41612 ( .A(n22316), .X(n45216) );
  nand_x1_sg U41613 ( .A(n28153), .B(n28154), .X(n22299) );
  inv_x1_sg U41614 ( .A(n28155), .X(n45196) );
  nand_x1_sg U41615 ( .A(n27647), .B(n45224), .X(n22298) );
  nand_x1_sg U41616 ( .A(n28004), .B(n45220), .X(n22294) );
  nand_x1_sg U41617 ( .A(n27444), .B(n45226), .X(n22295) );
  nand_x1_sg U41618 ( .A(n27833), .B(n45222), .X(n22304) );
  nand_x1_sg U41619 ( .A(n27222), .B(n45228), .X(n22305) );
  inv_x1_sg U41620 ( .A(n29020), .X(n45202) );
  nand_x1_sg U41621 ( .A(n29124), .B(n29125), .X(n29020) );
  inv_x1_sg U41622 ( .A(n28498), .X(n45199) );
  nand_x1_sg U41623 ( .A(n28606), .B(n28607), .X(n28498) );
  inv_x1_sg U41624 ( .A(n28841), .X(n45156) );
  nand_x1_sg U41625 ( .A(n28967), .B(n28968), .X(n28841) );
  inv_x1_sg U41626 ( .A(n28398), .X(n45153) );
  nand_x1_sg U41627 ( .A(n28449), .B(n28450), .X(n28398) );
  inv_x1_sg U41628 ( .A(n26982), .X(n45143) );
  nand_x1_sg U41629 ( .A(n27178), .B(n27179), .X(n26982) );
  inv_x1_sg U41630 ( .A(n22373), .X(n45142) );
  nand_x1_sg U41631 ( .A(n26939), .B(n26940), .X(n22373) );
  inv_x1_sg U41632 ( .A(n28653), .X(n45155) );
  nand_x1_sg U41633 ( .A(n28797), .B(n28798), .X(n28653) );
  inv_x1_sg U41634 ( .A(n22363), .X(n45170) );
  nand_x1_sg U41635 ( .A(n28148), .B(n28149), .X(n22347) );
  inv_x1_sg U41636 ( .A(n28150), .X(n45151) );
  nand_x1_sg U41637 ( .A(n27641), .B(n45178), .X(n22346) );
  nand_x1_sg U41638 ( .A(n27998), .B(n45174), .X(n22342) );
  nand_x1_sg U41639 ( .A(n27438), .B(n45180), .X(n22343) );
  nand_x1_sg U41640 ( .A(n27827), .B(n45176), .X(n22352) );
  nand_x1_sg U41641 ( .A(n27216), .B(n45182), .X(n22353) );
  nand_x1_sg U41642 ( .A(n29257), .B(n29258), .X(n29166) );
  nand_x1_sg U41643 ( .A(out_L1[4]), .B(n29259), .X(n29258) );
  nand_x1_sg U41644 ( .A(n5413), .B(n45066), .X(n29259) );
  inv_x1_sg U41645 ( .A(n29014), .X(n45157) );
  nand_x1_sg U41646 ( .A(n29127), .B(n29128), .X(n29014) );
  inv_x1_sg U41647 ( .A(n28492), .X(n45154) );
  nand_x1_sg U41648 ( .A(n28609), .B(n28610), .X(n28492) );
  inv_x1_sg U41649 ( .A(n28835), .X(n45110) );
  nand_x1_sg U41650 ( .A(n28970), .B(n28971), .X(n28835) );
  inv_x1_sg U41651 ( .A(n28392), .X(n45107) );
  nand_x1_sg U41652 ( .A(n28452), .B(n28453), .X(n28392) );
  inv_x1_sg U41653 ( .A(n26976), .X(n45096) );
  nand_x1_sg U41654 ( .A(n27181), .B(n27182), .X(n26976) );
  inv_x1_sg U41655 ( .A(n22421), .X(n45095) );
  nand_x1_sg U41656 ( .A(n26942), .B(n26943), .X(n22421) );
  nor_x4_sg U41657 ( .A(n42115), .B(out_L1[4]), .X(n29163) );
  inv_x1_sg U41658 ( .A(n28647), .X(n45109) );
  nand_x1_sg U41659 ( .A(n28800), .B(n28801), .X(n28647) );
  inv_x1_sg U41660 ( .A(n22411), .X(n45125) );
  nand_x1_sg U41661 ( .A(n27992), .B(n45129), .X(n22389) );
  nand_x1_sg U41662 ( .A(n27432), .B(n45135), .X(n22390) );
  nand_x1_sg U41663 ( .A(n28143), .B(n28144), .X(n22394) );
  inv_x1_sg U41664 ( .A(n28145), .X(n45105) );
  nand_x1_sg U41665 ( .A(n27635), .B(n45133), .X(n22393) );
  nand_x1_sg U41666 ( .A(n27821), .B(n45131), .X(n22399) );
  nand_x1_sg U41667 ( .A(n27210), .B(n45137), .X(n22400) );
  inv_x1_sg U41668 ( .A(n29007), .X(n45111) );
  nand_x1_sg U41669 ( .A(n29130), .B(n29131), .X(n29007) );
  inv_x1_sg U41670 ( .A(n28486), .X(n45108) );
  nand_x1_sg U41671 ( .A(n28612), .B(n28613), .X(n28486) );
  inv_x1_sg U41672 ( .A(n28829), .X(n45064) );
  nand_x1_sg U41673 ( .A(n28973), .B(n28974), .X(n28829) );
  inv_x1_sg U41674 ( .A(n28386), .X(n45061) );
  nand_x1_sg U41675 ( .A(n28455), .B(n28456), .X(n28386) );
  inv_x1_sg U41676 ( .A(n26970), .X(n45052) );
  nand_x1_sg U41677 ( .A(n27184), .B(n27185), .X(n26970) );
  inv_x1_sg U41678 ( .A(n22467), .X(n45051) );
  nand_x1_sg U41679 ( .A(n26945), .B(n26946), .X(n22467) );
  inv_x1_sg U41680 ( .A(n28641), .X(n45063) );
  nand_x1_sg U41681 ( .A(n28803), .B(n28804), .X(n28641) );
  inv_x1_sg U41682 ( .A(n22457), .X(n45078) );
  nand_x1_sg U41683 ( .A(n27629), .B(n45086), .X(n22441) );
  nand_x1_sg U41684 ( .A(n27985), .B(n45082), .X(n22437) );
  nand_x1_sg U41685 ( .A(n27426), .B(n45088), .X(n22438) );
  nand_x1_sg U41686 ( .A(n27815), .B(n45084), .X(n22446) );
  nand_x1_sg U41687 ( .A(n27204), .B(n45090), .X(n22447) );
  nand_x1_sg U41688 ( .A(n29263), .B(n29264), .X(n29154) );
  nand_x1_sg U41689 ( .A(out_L1[2]), .B(n29265), .X(n29264) );
  nand_x1_sg U41690 ( .A(n5415), .B(n45021), .X(n29265) );
  inv_x1_sg U41691 ( .A(n29001), .X(n45065) );
  nand_x1_sg U41692 ( .A(n29133), .B(n29134), .X(n29001) );
  inv_x1_sg U41693 ( .A(n28480), .X(n45062) );
  nand_x1_sg U41694 ( .A(n28615), .B(n28616), .X(n28480) );
  nor_x4_sg U41695 ( .A(n42114), .B(out_L1[2]), .X(n29151) );
  nand_x1_sg U41696 ( .A(n27623), .B(n45042), .X(n22487) );
  nand_x1_sg U41697 ( .A(n27978), .B(n45038), .X(n22483) );
  nand_x1_sg U41698 ( .A(n27420), .B(n45044), .X(n22484) );
  nand_x1_sg U41699 ( .A(n27809), .B(n45040), .X(n22492) );
  nand_x1_sg U41700 ( .A(n27198), .B(n45046), .X(n22493) );
  nand_x1_sg U41701 ( .A(n22552), .B(n38559), .X(n22550) );
  nand_x1_sg U41702 ( .A(n44972), .B(n27411), .X(n22566) );
  nand_x1_sg U41703 ( .A(n46943), .B(n22774), .X(n22773) );
  inv_x1_sg U41704 ( .A(n22767), .X(n46942) );
  nand_x1_sg U41705 ( .A(n46985), .B(n22760), .X(n22759) );
  nand_x1_sg U41706 ( .A(n47008), .B(n46984), .X(n22752) );
  nand_x1_sg U41707 ( .A(n47027), .B(n22746), .X(n22745) );
  nand_x1_sg U41708 ( .A(n47217), .B(n47196), .X(n23057) );
  nand_x1_sg U41709 ( .A(n47234), .B(n23051), .X(n23050) );
  nand_x1_sg U41710 ( .A(n47274), .B(n23037), .X(n23036) );
  nand_x1_sg U41711 ( .A(n47296), .B(n47273), .X(n23029) );
  nand_x1_sg U41712 ( .A(n47314), .B(n23023), .X(n23022) );
  nand_x1_sg U41713 ( .A(n47502), .B(n47481), .X(n23337) );
  nand_x1_sg U41714 ( .A(n47519), .B(n23331), .X(n23330) );
  inv_x1_sg U41715 ( .A(n23331), .X(n47501) );
  nand_x1_sg U41716 ( .A(n47559), .B(n23317), .X(n23316) );
  nand_x1_sg U41717 ( .A(n47581), .B(n47558), .X(n23309) );
  nand_x1_sg U41718 ( .A(n47599), .B(n23303), .X(n23302) );
  nand_x1_sg U41719 ( .A(n47787), .B(n47766), .X(n23616) );
  nand_x1_sg U41720 ( .A(n47804), .B(n23610), .X(n23609) );
  nand_x1_sg U41721 ( .A(n47844), .B(n23596), .X(n23595) );
  nand_x1_sg U41722 ( .A(n47866), .B(n47843), .X(n23588) );
  nand_x1_sg U41723 ( .A(n47884), .B(n23582), .X(n23581) );
  nand_x1_sg U41724 ( .A(n48072), .B(n48051), .X(n23895) );
  nand_x1_sg U41725 ( .A(n48089), .B(n23889), .X(n23888) );
  inv_x1_sg U41726 ( .A(n23889), .X(n48071) );
  nand_x1_sg U41727 ( .A(n48129), .B(n23875), .X(n23874) );
  nand_x1_sg U41728 ( .A(n48151), .B(n48128), .X(n23867) );
  nand_x1_sg U41729 ( .A(n48169), .B(n23861), .X(n23860) );
  nand_x1_sg U41730 ( .A(n23845), .B(n23846), .X(n10272) );
  nand_x1_sg U41731 ( .A(n48357), .B(n48336), .X(n24174) );
  nand_x1_sg U41732 ( .A(n48374), .B(n24168), .X(n24167) );
  nand_x1_sg U41733 ( .A(n48414), .B(n24154), .X(n24153) );
  nand_x1_sg U41734 ( .A(n48454), .B(n24140), .X(n24139) );
  nand_x1_sg U41735 ( .A(n48642), .B(n48621), .X(n24453) );
  nand_x1_sg U41736 ( .A(n48659), .B(n24447), .X(n24446) );
  nand_x1_sg U41737 ( .A(n48699), .B(n24433), .X(n24432) );
  nand_x1_sg U41738 ( .A(n48721), .B(n48698), .X(n24425) );
  nand_x1_sg U41739 ( .A(n48739), .B(n24419), .X(n24418) );
  nand_x1_sg U41740 ( .A(n48928), .B(n48907), .X(n24731) );
  nand_x1_sg U41741 ( .A(n48945), .B(n24725), .X(n24724) );
  nand_x1_sg U41742 ( .A(n48985), .B(n24711), .X(n24710) );
  nand_x1_sg U41743 ( .A(n49007), .B(n48984), .X(n24703) );
  nand_x1_sg U41744 ( .A(n49025), .B(n24697), .X(n24696) );
  nand_x1_sg U41745 ( .A(n49215), .B(n49194), .X(n25010) );
  nand_x1_sg U41746 ( .A(n49232), .B(n25004), .X(n25003) );
  nand_x1_sg U41747 ( .A(n49272), .B(n24990), .X(n24989) );
  nand_x1_sg U41748 ( .A(n49294), .B(n49271), .X(n24982) );
  nand_x1_sg U41749 ( .A(n49312), .B(n24976), .X(n24975) );
  nand_x1_sg U41750 ( .A(n24960), .B(n24961), .X(n13548) );
  nand_x1_sg U41751 ( .A(n49501), .B(n49480), .X(n25289) );
  nand_x1_sg U41752 ( .A(n49518), .B(n25283), .X(n25282) );
  nand_x1_sg U41753 ( .A(n49558), .B(n25269), .X(n25268) );
  nand_x1_sg U41754 ( .A(n49580), .B(n49557), .X(n25261) );
  nand_x1_sg U41755 ( .A(n49598), .B(n25255), .X(n25254) );
  inv_x1_sg U41756 ( .A(n25248), .X(n49597) );
  nand_x1_sg U41757 ( .A(n49804), .B(n25562), .X(n25561) );
  nand_x1_sg U41758 ( .A(n49844), .B(n25548), .X(n25547) );
  nand_x1_sg U41759 ( .A(n49866), .B(n49843), .X(n25540) );
  nand_x1_sg U41760 ( .A(n49884), .B(n25534), .X(n25533) );
  nand_x1_sg U41761 ( .A(n50090), .B(n25839), .X(n25838) );
  inv_x1_sg U41762 ( .A(n25839), .X(n50072) );
  nand_x1_sg U41763 ( .A(n50130), .B(n25825), .X(n25824) );
  nand_x1_sg U41764 ( .A(n50152), .B(n50129), .X(n25817) );
  nand_x1_sg U41765 ( .A(n50170), .B(n25811), .X(n25810) );
  nand_x1_sg U41766 ( .A(n50278), .B(n26171), .X(n26113) );
  nand_x1_sg U41767 ( .A(n50358), .B(n50356), .X(n26076) );
  nand_x1_sg U41768 ( .A(n50375), .B(n26071), .X(n26070) );
  nand_x1_sg U41769 ( .A(n50415), .B(n26059), .X(n26058) );
  nand_x1_sg U41770 ( .A(n50437), .B(n50435), .X(n26052) );
  nand_x1_sg U41771 ( .A(n50455), .B(n26047), .X(n26046) );
  inv_x1_sg U41772 ( .A(n26136), .X(n50500) );
  nand_x1_sg U41773 ( .A(n50647), .B(n50626), .X(n26405) );
  nand_x1_sg U41774 ( .A(n50664), .B(n26399), .X(n26398) );
  nand_x1_sg U41775 ( .A(n50704), .B(n26385), .X(n26384) );
  nand_x1_sg U41776 ( .A(n50726), .B(n50703), .X(n26377) );
  nand_x1_sg U41777 ( .A(n50744), .B(n26371), .X(n26370) );
  nand_x1_sg U41778 ( .A(n26355), .B(n26356), .X(n17643) );
  nand_x1_sg U41779 ( .A(n50934), .B(n50913), .X(n26683) );
  nand_x1_sg U41780 ( .A(n50951), .B(n26677), .X(n26676) );
  nand_x1_sg U41781 ( .A(n50991), .B(n26663), .X(n26662) );
  nand_x1_sg U41782 ( .A(n51013), .B(n50990), .X(n26655) );
  nand_x1_sg U41783 ( .A(n51031), .B(n26649), .X(n26648) );
  nand_x1_sg U41784 ( .A(n26633), .B(n26634), .X(n18464) );
  nand_x1_sg U41785 ( .A(n20975), .B(n46618), .X(n20563) );
  nand_x1_sg U41786 ( .A(n20978), .B(n20977), .X(n20975) );
  nand_x1_sg U41787 ( .A(n46584), .B(n21180), .X(n5995) );
  nand_x1_sg U41788 ( .A(n21350), .B(n46544), .X(n6043) );
  nand_x1_sg U41789 ( .A(n21532), .B(n46502), .X(n6093) );
  inv_x1_sg U41790 ( .A(n20143), .X(n41532) );
  nand_x1_sg U41791 ( .A(n21667), .B(n46417), .X(n6184) );
  inv_x1_sg U41792 ( .A(n19899), .X(n41538) );
  nand_x1_sg U41793 ( .A(n21655), .B(n46328), .X(n6275) );
  nand_x1_sg U41794 ( .A(n21643), .B(n46237), .X(n6364) );
  nand_x1_sg U41795 ( .A(n21631), .B(n46146), .X(n6453) );
  nand_x1_sg U41796 ( .A(n21619), .B(n46055), .X(n6542) );
  nand_x1_sg U41797 ( .A(n21607), .B(n45964), .X(n6631) );
  nand_x1_sg U41798 ( .A(n21595), .B(n45872), .X(n6723) );
  inv_x1_sg U41799 ( .A(n21076), .X(n41536) );
  inv_x1_sg U41800 ( .A(n20367), .X(n41535) );
  nand_x1_sg U41801 ( .A(n7090), .B(n7089), .X(n7064) );
  nand_x1_sg U41802 ( .A(n46895), .B(n7113), .X(n7112) );
  nand_x1_sg U41803 ( .A(n7121), .B(n7122), .X(n7119) );
  nand_x1_sg U41804 ( .A(n7142), .B(n46909), .X(n7120) );
  nand_x1_sg U41805 ( .A(n7148), .B(n7147), .X(n7060) );
  nand_x1_sg U41806 ( .A(n7175), .B(n7176), .X(n7173) );
  nand_x1_sg U41807 ( .A(n7194), .B(n46949), .X(n7174) );
  nand_x1_sg U41808 ( .A(n7200), .B(n7199), .X(n7057) );
  nand_x1_sg U41809 ( .A(n7237), .B(n7236), .X(n7055) );
  nand_x1_sg U41810 ( .A(n7265), .B(n7264), .X(n7053) );
  nand_x1_sg U41811 ( .A(n7316), .B(n7315), .X(n7051) );
  nand_x1_sg U41812 ( .A(n7351), .B(n7350), .X(n7049) );
  nand_x1_sg U41813 ( .A(n7408), .B(n7407), .X(n7047) );
  nand_x1_sg U41814 ( .A(n7456), .B(n7455), .X(n7045) );
  nand_x1_sg U41815 ( .A(n6974), .B(n6975), .X(n6973) );
  nand_x1_sg U41816 ( .A(n23127), .B(n23128), .X(n23126) );
  nand_x1_sg U41817 ( .A(n7908), .B(n7907), .X(n7882) );
  nand_x1_sg U41818 ( .A(n47190), .B(n7931), .X(n7930) );
  nand_x1_sg U41819 ( .A(n7939), .B(n7940), .X(n7937) );
  nand_x1_sg U41820 ( .A(n7960), .B(n47202), .X(n7938) );
  nand_x1_sg U41821 ( .A(n7966), .B(n7965), .X(n7878) );
  nand_x1_sg U41822 ( .A(n7994), .B(n7995), .X(n7992) );
  nand_x1_sg U41823 ( .A(n8013), .B(n47240), .X(n7993) );
  nand_x1_sg U41824 ( .A(n8019), .B(n8018), .X(n7875) );
  nand_x1_sg U41825 ( .A(n8056), .B(n8055), .X(n7873) );
  nand_x1_sg U41826 ( .A(n47288), .B(n8080), .X(n8086) );
  nand_x1_sg U41827 ( .A(n8084), .B(n8083), .X(n7871) );
  nand_x1_sg U41828 ( .A(n8134), .B(n8133), .X(n7869) );
  nand_x1_sg U41829 ( .A(n8169), .B(n8168), .X(n7867) );
  nand_x1_sg U41830 ( .A(n8226), .B(n8225), .X(n7865) );
  nand_x1_sg U41831 ( .A(n8274), .B(n8273), .X(n7863) );
  nand_x1_sg U41832 ( .A(n7791), .B(n7792), .X(n7790) );
  nand_x1_sg U41833 ( .A(n8726), .B(n8725), .X(n8700) );
  nand_x1_sg U41834 ( .A(n47475), .B(n8749), .X(n8748) );
  nand_x1_sg U41835 ( .A(n8757), .B(n8758), .X(n8755) );
  nand_x1_sg U41836 ( .A(n8778), .B(n47487), .X(n8756) );
  nand_x1_sg U41837 ( .A(n8784), .B(n8783), .X(n8696) );
  nand_x1_sg U41838 ( .A(n8812), .B(n8813), .X(n8810) );
  nand_x1_sg U41839 ( .A(n8831), .B(n47525), .X(n8811) );
  nand_x1_sg U41840 ( .A(n8837), .B(n8836), .X(n8693) );
  nand_x1_sg U41841 ( .A(n8874), .B(n8873), .X(n8691) );
  nand_x1_sg U41842 ( .A(n47573), .B(n8898), .X(n8904) );
  nand_x1_sg U41843 ( .A(n8902), .B(n8901), .X(n8689) );
  nand_x1_sg U41844 ( .A(n8952), .B(n8951), .X(n8687) );
  nand_x1_sg U41845 ( .A(n8987), .B(n8986), .X(n8685) );
  nand_x1_sg U41846 ( .A(n9044), .B(n9043), .X(n8683) );
  nand_x1_sg U41847 ( .A(n9092), .B(n9091), .X(n8681) );
  nand_x1_sg U41848 ( .A(n8609), .B(n8610), .X(n8608) );
  nand_x1_sg U41849 ( .A(n9546), .B(n9545), .X(n9520) );
  nand_x1_sg U41850 ( .A(n47760), .B(n9569), .X(n9568) );
  nand_x1_sg U41851 ( .A(n9577), .B(n9578), .X(n9575) );
  nand_x1_sg U41852 ( .A(n9598), .B(n47772), .X(n9576) );
  nand_x1_sg U41853 ( .A(n9604), .B(n9603), .X(n9516) );
  nand_x1_sg U41854 ( .A(n9632), .B(n9633), .X(n9630) );
  nand_x1_sg U41855 ( .A(n9651), .B(n47810), .X(n9631) );
  nand_x1_sg U41856 ( .A(n9657), .B(n9656), .X(n9513) );
  nand_x1_sg U41857 ( .A(n9694), .B(n9693), .X(n9511) );
  nand_x1_sg U41858 ( .A(n47858), .B(n9718), .X(n9724) );
  nand_x1_sg U41859 ( .A(n9722), .B(n9721), .X(n9509) );
  nand_x1_sg U41860 ( .A(n9772), .B(n9771), .X(n9507) );
  nand_x1_sg U41861 ( .A(n9807), .B(n9806), .X(n9505) );
  nand_x1_sg U41862 ( .A(n9864), .B(n9863), .X(n9503) );
  nand_x1_sg U41863 ( .A(n9912), .B(n9911), .X(n9501) );
  nand_x1_sg U41864 ( .A(n9429), .B(n9430), .X(n9428) );
  nand_x1_sg U41865 ( .A(n10365), .B(n10364), .X(n10339) );
  nand_x1_sg U41866 ( .A(n48045), .B(n10388), .X(n10387) );
  nand_x1_sg U41867 ( .A(n10396), .B(n10397), .X(n10394) );
  nand_x1_sg U41868 ( .A(n10417), .B(n48057), .X(n10395) );
  nand_x1_sg U41869 ( .A(n10423), .B(n10422), .X(n10335) );
  nand_x1_sg U41870 ( .A(n10451), .B(n10452), .X(n10449) );
  nand_x1_sg U41871 ( .A(n10470), .B(n48095), .X(n10450) );
  nand_x1_sg U41872 ( .A(n10476), .B(n10475), .X(n10332) );
  nand_x1_sg U41873 ( .A(n10513), .B(n10512), .X(n10330) );
  nand_x1_sg U41874 ( .A(n48143), .B(n10537), .X(n10543) );
  nand_x1_sg U41875 ( .A(n10541), .B(n10540), .X(n10328) );
  nand_x1_sg U41876 ( .A(n10591), .B(n10590), .X(n10326) );
  nand_x1_sg U41877 ( .A(n10626), .B(n10625), .X(n10324) );
  nand_x1_sg U41878 ( .A(n10683), .B(n10682), .X(n10322) );
  nand_x1_sg U41879 ( .A(n10731), .B(n10730), .X(n10320) );
  nand_x1_sg U41880 ( .A(n10248), .B(n10249), .X(n10247) );
  nand_x1_sg U41881 ( .A(n11184), .B(n11183), .X(n11158) );
  nand_x1_sg U41882 ( .A(n48330), .B(n11207), .X(n11206) );
  nand_x1_sg U41883 ( .A(n11215), .B(n11216), .X(n11213) );
  nand_x1_sg U41884 ( .A(n11236), .B(n48342), .X(n11214) );
  nand_x1_sg U41885 ( .A(n11242), .B(n11241), .X(n11154) );
  nand_x1_sg U41886 ( .A(n11270), .B(n11271), .X(n11268) );
  nand_x1_sg U41887 ( .A(n11289), .B(n48380), .X(n11269) );
  nand_x1_sg U41888 ( .A(n11295), .B(n11294), .X(n11151) );
  nand_x1_sg U41889 ( .A(n11332), .B(n11331), .X(n11149) );
  nand_x1_sg U41890 ( .A(n48428), .B(n11356), .X(n11362) );
  nand_x1_sg U41891 ( .A(n11360), .B(n11359), .X(n11147) );
  nand_x1_sg U41892 ( .A(n11410), .B(n11409), .X(n11145) );
  nand_x1_sg U41893 ( .A(n11445), .B(n11444), .X(n11143) );
  nand_x1_sg U41894 ( .A(n11502), .B(n11501), .X(n11141) );
  nand_x1_sg U41895 ( .A(n11550), .B(n11549), .X(n11139) );
  nand_x1_sg U41896 ( .A(n11067), .B(n11068), .X(n11066) );
  nand_x1_sg U41897 ( .A(n12003), .B(n12002), .X(n11977) );
  nand_x1_sg U41898 ( .A(n48615), .B(n12026), .X(n12025) );
  nand_x1_sg U41899 ( .A(n12034), .B(n12035), .X(n12032) );
  nand_x1_sg U41900 ( .A(n12055), .B(n48627), .X(n12033) );
  nand_x1_sg U41901 ( .A(n12061), .B(n12060), .X(n11973) );
  nand_x1_sg U41902 ( .A(n12089), .B(n12090), .X(n12087) );
  nand_x1_sg U41903 ( .A(n12108), .B(n48665), .X(n12088) );
  nand_x1_sg U41904 ( .A(n12114), .B(n12113), .X(n11970) );
  nand_x1_sg U41905 ( .A(n12151), .B(n12150), .X(n11968) );
  nand_x1_sg U41906 ( .A(n48713), .B(n12175), .X(n12181) );
  nand_x1_sg U41907 ( .A(n12179), .B(n12178), .X(n11966) );
  nand_x1_sg U41908 ( .A(n12229), .B(n12228), .X(n11964) );
  nand_x1_sg U41909 ( .A(n12264), .B(n12263), .X(n11962) );
  nand_x1_sg U41910 ( .A(n12321), .B(n12320), .X(n11960) );
  nand_x1_sg U41911 ( .A(n12369), .B(n12368), .X(n11958) );
  nand_x1_sg U41912 ( .A(n11886), .B(n11887), .X(n11885) );
  nand_x1_sg U41913 ( .A(n12822), .B(n12821), .X(n12796) );
  nand_x1_sg U41914 ( .A(n48901), .B(n12845), .X(n12844) );
  nand_x1_sg U41915 ( .A(n12853), .B(n12854), .X(n12851) );
  nand_x1_sg U41916 ( .A(n12874), .B(n48913), .X(n12852) );
  nand_x1_sg U41917 ( .A(n12880), .B(n12879), .X(n12792) );
  nand_x1_sg U41918 ( .A(n12908), .B(n12909), .X(n12906) );
  nand_x1_sg U41919 ( .A(n12927), .B(n48951), .X(n12907) );
  nand_x1_sg U41920 ( .A(n12933), .B(n12932), .X(n12789) );
  nand_x1_sg U41921 ( .A(n12970), .B(n12969), .X(n12787) );
  nand_x1_sg U41922 ( .A(n48999), .B(n12994), .X(n13000) );
  nand_x1_sg U41923 ( .A(n12998), .B(n12997), .X(n12785) );
  nand_x1_sg U41924 ( .A(n13048), .B(n13047), .X(n12783) );
  nand_x1_sg U41925 ( .A(n13083), .B(n13082), .X(n12781) );
  nand_x1_sg U41926 ( .A(n13140), .B(n13139), .X(n12779) );
  nand_x1_sg U41927 ( .A(n13188), .B(n13187), .X(n12777) );
  nand_x1_sg U41928 ( .A(n12705), .B(n12706), .X(n12704) );
  nand_x1_sg U41929 ( .A(n13641), .B(n13640), .X(n13615) );
  nand_x1_sg U41930 ( .A(n49188), .B(n13664), .X(n13663) );
  nand_x1_sg U41931 ( .A(n13672), .B(n13673), .X(n13670) );
  nand_x1_sg U41932 ( .A(n13693), .B(n49200), .X(n13671) );
  nand_x1_sg U41933 ( .A(n13699), .B(n13698), .X(n13611) );
  nand_x1_sg U41934 ( .A(n13727), .B(n13728), .X(n13725) );
  nand_x1_sg U41935 ( .A(n13746), .B(n49238), .X(n13726) );
  nand_x1_sg U41936 ( .A(n13752), .B(n13751), .X(n13608) );
  nand_x1_sg U41937 ( .A(n13789), .B(n13788), .X(n13606) );
  nand_x1_sg U41938 ( .A(n49286), .B(n13813), .X(n13819) );
  nand_x1_sg U41939 ( .A(n13817), .B(n13816), .X(n13604) );
  nand_x1_sg U41940 ( .A(n13867), .B(n13866), .X(n13602) );
  nand_x1_sg U41941 ( .A(n13902), .B(n13901), .X(n13600) );
  nand_x1_sg U41942 ( .A(n13959), .B(n13958), .X(n13598) );
  nand_x1_sg U41943 ( .A(n14007), .B(n14006), .X(n13596) );
  nand_x1_sg U41944 ( .A(n13524), .B(n13525), .X(n13523) );
  nand_x1_sg U41945 ( .A(n14460), .B(n14459), .X(n14434) );
  nand_x1_sg U41946 ( .A(n49474), .B(n14483), .X(n14482) );
  nand_x1_sg U41947 ( .A(n14491), .B(n14492), .X(n14489) );
  nand_x1_sg U41948 ( .A(n14512), .B(n49486), .X(n14490) );
  nand_x1_sg U41949 ( .A(n14518), .B(n14517), .X(n14430) );
  nand_x1_sg U41950 ( .A(n14546), .B(n14547), .X(n14544) );
  nand_x1_sg U41951 ( .A(n14565), .B(n49524), .X(n14545) );
  nand_x1_sg U41952 ( .A(n14571), .B(n14570), .X(n14427) );
  nand_x1_sg U41953 ( .A(n14608), .B(n14607), .X(n14425) );
  nand_x1_sg U41954 ( .A(n49572), .B(n14632), .X(n14638) );
  nand_x1_sg U41955 ( .A(n14636), .B(n14635), .X(n14423) );
  nand_x1_sg U41956 ( .A(n14686), .B(n14685), .X(n14421) );
  nand_x1_sg U41957 ( .A(n14721), .B(n14720), .X(n14419) );
  nand_x1_sg U41958 ( .A(n14778), .B(n14777), .X(n14417) );
  nand_x1_sg U41959 ( .A(n14826), .B(n14825), .X(n14415) );
  nand_x1_sg U41960 ( .A(n14343), .B(n14344), .X(n14342) );
  nand_x1_sg U41961 ( .A(n15279), .B(n15278), .X(n15253) );
  nand_x1_sg U41962 ( .A(n49760), .B(n15302), .X(n15301) );
  nand_x1_sg U41963 ( .A(n15310), .B(n15311), .X(n15308) );
  nand_x1_sg U41964 ( .A(n15331), .B(n49772), .X(n15309) );
  nand_x1_sg U41965 ( .A(n15337), .B(n15336), .X(n15249) );
  nand_x1_sg U41966 ( .A(n15365), .B(n15366), .X(n15363) );
  nand_x1_sg U41967 ( .A(n15384), .B(n49810), .X(n15364) );
  nand_x1_sg U41968 ( .A(n15390), .B(n15389), .X(n15246) );
  nand_x1_sg U41969 ( .A(n15427), .B(n15426), .X(n15244) );
  nand_x1_sg U41970 ( .A(n49858), .B(n15451), .X(n15457) );
  nand_x1_sg U41971 ( .A(n15455), .B(n15454), .X(n15242) );
  nand_x1_sg U41972 ( .A(n15505), .B(n15504), .X(n15240) );
  nand_x1_sg U41973 ( .A(n15540), .B(n15539), .X(n15238) );
  nand_x1_sg U41974 ( .A(n15597), .B(n15596), .X(n15236) );
  nand_x1_sg U41975 ( .A(n15645), .B(n15644), .X(n15234) );
  nand_x1_sg U41976 ( .A(n15162), .B(n15163), .X(n15161) );
  nand_x1_sg U41977 ( .A(n16098), .B(n16097), .X(n16072) );
  nand_x1_sg U41978 ( .A(n50046), .B(n16121), .X(n16120) );
  nand_x1_sg U41979 ( .A(n16129), .B(n16130), .X(n16127) );
  nand_x1_sg U41980 ( .A(n16150), .B(n50058), .X(n16128) );
  nand_x1_sg U41981 ( .A(n16156), .B(n16155), .X(n16068) );
  nand_x1_sg U41982 ( .A(n16184), .B(n16185), .X(n16182) );
  nand_x1_sg U41983 ( .A(n16203), .B(n50096), .X(n16183) );
  nand_x1_sg U41984 ( .A(n16209), .B(n16208), .X(n16065) );
  nand_x1_sg U41985 ( .A(n16246), .B(n16245), .X(n16063) );
  nand_x1_sg U41986 ( .A(n50144), .B(n16270), .X(n16276) );
  nand_x1_sg U41987 ( .A(n16274), .B(n16273), .X(n16061) );
  nand_x1_sg U41988 ( .A(n16324), .B(n16323), .X(n16059) );
  nand_x1_sg U41989 ( .A(n16359), .B(n16358), .X(n16057) );
  nand_x1_sg U41990 ( .A(n16416), .B(n16415), .X(n16055) );
  nand_x1_sg U41991 ( .A(n16464), .B(n16463), .X(n16053) );
  nand_x1_sg U41992 ( .A(n15981), .B(n15982), .X(n15980) );
  nand_x1_sg U41993 ( .A(n16916), .B(n16915), .X(n16891) );
  nand_x1_sg U41994 ( .A(n50328), .B(n16938), .X(n16937) );
  nand_x1_sg U41995 ( .A(n16946), .B(n16947), .X(n16944) );
  nand_x1_sg U41996 ( .A(n16967), .B(n50343), .X(n16945) );
  nand_x1_sg U41997 ( .A(n16973), .B(n16972), .X(n16887) );
  nand_x1_sg U41998 ( .A(n17000), .B(n17001), .X(n16998) );
  nand_x1_sg U41999 ( .A(n17019), .B(n50381), .X(n16999) );
  nand_x1_sg U42000 ( .A(n17025), .B(n17024), .X(n16884) );
  nand_x1_sg U42001 ( .A(n17062), .B(n17061), .X(n16882) );
  nand_x1_sg U42002 ( .A(n17090), .B(n17089), .X(n16880) );
  nand_x1_sg U42003 ( .A(n17141), .B(n17140), .X(n16878) );
  nand_x1_sg U42004 ( .A(n17176), .B(n17175), .X(n16876) );
  nand_x1_sg U42005 ( .A(n17233), .B(n17232), .X(n16874) );
  nand_x1_sg U42006 ( .A(n17281), .B(n17280), .X(n16872) );
  nand_x1_sg U42007 ( .A(n16798), .B(n16799), .X(n16797) );
  nand_x1_sg U42008 ( .A(n17736), .B(n17735), .X(n17710) );
  nand_x1_sg U42009 ( .A(n50620), .B(n17759), .X(n17758) );
  nand_x1_sg U42010 ( .A(n17767), .B(n17768), .X(n17765) );
  nand_x1_sg U42011 ( .A(n17788), .B(n50632), .X(n17766) );
  nand_x1_sg U42012 ( .A(n17794), .B(n17793), .X(n17706) );
  nand_x1_sg U42013 ( .A(n17822), .B(n17823), .X(n17820) );
  nand_x1_sg U42014 ( .A(n17841), .B(n50670), .X(n17821) );
  nand_x1_sg U42015 ( .A(n17847), .B(n17846), .X(n17703) );
  nand_x1_sg U42016 ( .A(n17884), .B(n17883), .X(n17701) );
  nand_x1_sg U42017 ( .A(n50718), .B(n17908), .X(n17914) );
  nand_x1_sg U42018 ( .A(n17912), .B(n17911), .X(n17699) );
  nand_x1_sg U42019 ( .A(n17962), .B(n17961), .X(n17697) );
  nand_x1_sg U42020 ( .A(n17997), .B(n17996), .X(n17695) );
  nand_x1_sg U42021 ( .A(n18054), .B(n18053), .X(n17693) );
  nand_x1_sg U42022 ( .A(n18102), .B(n18101), .X(n17691) );
  nand_x1_sg U42023 ( .A(n17619), .B(n17620), .X(n17618) );
  nand_x1_sg U42024 ( .A(n18557), .B(n18556), .X(n18531) );
  nand_x1_sg U42025 ( .A(n50907), .B(n18580), .X(n18579) );
  nand_x1_sg U42026 ( .A(n18588), .B(n18589), .X(n18586) );
  nand_x1_sg U42027 ( .A(n18609), .B(n50919), .X(n18587) );
  nand_x1_sg U42028 ( .A(n18615), .B(n18614), .X(n18527) );
  nand_x1_sg U42029 ( .A(n18643), .B(n18644), .X(n18641) );
  nand_x1_sg U42030 ( .A(n18662), .B(n50957), .X(n18642) );
  nand_x1_sg U42031 ( .A(n18668), .B(n18667), .X(n18524) );
  nand_x1_sg U42032 ( .A(n18705), .B(n18704), .X(n18522) );
  nand_x1_sg U42033 ( .A(n51005), .B(n18729), .X(n18735) );
  nand_x1_sg U42034 ( .A(n18733), .B(n18732), .X(n18520) );
  nand_x1_sg U42035 ( .A(n18783), .B(n18782), .X(n18518) );
  nand_x1_sg U42036 ( .A(n18818), .B(n18817), .X(n18516) );
  nand_x1_sg U42037 ( .A(n18875), .B(n18874), .X(n18514) );
  nand_x1_sg U42038 ( .A(n18923), .B(n18922), .X(n18512) );
  nand_x1_sg U42039 ( .A(n18440), .B(n18441), .X(n18439) );
  nand_x1_sg U42040 ( .A(n5303), .B(n26832), .X(n26831) );
  nand_x1_sg U42041 ( .A(n5360), .B(n28552), .X(n28551) );
  nand_x1_sg U42042 ( .A(n5132), .B(n26896), .X(n26895) );
  nand_x1_sg U42043 ( .A(n5151), .B(n26889), .X(n26888) );
  nand_x1_sg U42044 ( .A(n45795), .B(n26805), .X(n26780) );
  nand_x1_sg U42045 ( .A(n5341), .B(n28559), .X(n28558) );
  nand_x1_sg U42046 ( .A(n28537), .B(n28538), .X(n28535) );
  nand_x1_sg U42047 ( .A(n38934), .B(n26771), .X(n26768) );
  nand_x1_sg U42048 ( .A(n26763), .B(n26764), .X(n26762) );
  nand_x1_sg U42049 ( .A(n5322), .B(n28566), .X(n28565) );
  nand_x1_sg U42050 ( .A(n5379), .B(n28545), .X(n28544) );
  inv_x1_sg U42051 ( .A(n21767), .X(n45743) );
  inv_x1_sg U42052 ( .A(n21766), .X(n45749) );
  inv_x1_sg U42053 ( .A(n21763), .X(n45767) );
  inv_x1_sg U42054 ( .A(n21751), .X(n45745) );
  inv_x1_sg U42055 ( .A(n21746), .X(n45741) );
  inv_x1_sg U42056 ( .A(n21745), .X(n45747) );
  inv_x1_sg U42057 ( .A(n21814), .X(n45700) );
  inv_x1_sg U42058 ( .A(n21813), .X(n45706) );
  inv_x1_sg U42059 ( .A(n21810), .X(n45724) );
  nand_x1_sg U42060 ( .A(n28917), .B(n28918), .X(n28741) );
  nand_x1_sg U42061 ( .A(out_L1[16]), .B(n45608), .X(n28918) );
  inv_x1_sg U42062 ( .A(n21798), .X(n45702) );
  inv_x1_sg U42063 ( .A(n21793), .X(n45698) );
  inv_x1_sg U42064 ( .A(n21792), .X(n45704) );
  inv_x1_sg U42065 ( .A(n21860), .X(n45662) );
  inv_x1_sg U42066 ( .A(n21861), .X(n45656) );
  inv_x1_sg U42067 ( .A(n21857), .X(n45681) );
  inv_x1_sg U42068 ( .A(n21845), .X(n45658) );
  nand_x1_sg U42069 ( .A(n29086), .B(n29087), .X(n28920) );
  nand_x1_sg U42070 ( .A(out_L1[15]), .B(n29088), .X(n29087) );
  inv_x1_sg U42071 ( .A(n21839), .X(n45660) );
  inv_x1_sg U42072 ( .A(n21840), .X(n45654) );
  inv_x1_sg U42073 ( .A(n21907), .X(n45612) );
  inv_x1_sg U42074 ( .A(n21906), .X(n45618) );
  inv_x1_sg U42075 ( .A(n21903), .X(n45637) );
  inv_x1_sg U42076 ( .A(n21891), .X(n45614) );
  inv_x1_sg U42077 ( .A(n21886), .X(n45616) );
  inv_x1_sg U42078 ( .A(n21954), .X(n45568) );
  inv_x1_sg U42079 ( .A(n21953), .X(n45574) );
  inv_x1_sg U42080 ( .A(n21950), .X(n45593) );
  nand_x1_sg U42081 ( .A(n29230), .B(n29231), .X(n29221) );
  nand_x1_sg U42082 ( .A(out_L1[13]), .B(n29232), .X(n29231) );
  inv_x1_sg U42083 ( .A(n21938), .X(n45570) );
  inv_x1_sg U42084 ( .A(n21933), .X(n45566) );
  inv_x1_sg U42085 ( .A(n21932), .X(n45572) );
  inv_x1_sg U42086 ( .A(n22000), .X(n45523) );
  inv_x1_sg U42087 ( .A(n21999), .X(n45529) );
  inv_x1_sg U42088 ( .A(n21996), .X(n45548) );
  inv_x1_sg U42089 ( .A(n21984), .X(n45525) );
  inv_x1_sg U42090 ( .A(n21979), .X(n45527) );
  inv_x1_sg U42091 ( .A(n22047), .X(n45479) );
  inv_x1_sg U42092 ( .A(n22046), .X(n45485) );
  inv_x1_sg U42093 ( .A(n22043), .X(n45504) );
  nand_x1_sg U42094 ( .A(n29236), .B(n29237), .X(n29209) );
  nand_x1_sg U42095 ( .A(out_L1[11]), .B(n29238), .X(n29237) );
  inv_x1_sg U42096 ( .A(n22031), .X(n45481) );
  inv_x1_sg U42097 ( .A(n22026), .X(n45477) );
  inv_x1_sg U42098 ( .A(n22025), .X(n45483) );
  inv_x1_sg U42099 ( .A(n22093), .X(n45434) );
  inv_x1_sg U42100 ( .A(n22092), .X(n45440) );
  inv_x1_sg U42101 ( .A(n22089), .X(n45456) );
  inv_x1_sg U42102 ( .A(n22077), .X(n45436) );
  inv_x1_sg U42103 ( .A(n22072), .X(n45438) );
  inv_x1_sg U42104 ( .A(n22140), .X(n45395) );
  inv_x1_sg U42105 ( .A(n22141), .X(n45389) );
  inv_x1_sg U42106 ( .A(n22137), .X(n45412) );
  inv_x1_sg U42107 ( .A(n22125), .X(n45391) );
  nand_x1_sg U42108 ( .A(n29242), .B(n29243), .X(n29197) );
  nand_x1_sg U42109 ( .A(out_L1[9]), .B(n29244), .X(n29243) );
  inv_x1_sg U42110 ( .A(n22119), .X(n45393) );
  inv_x1_sg U42111 ( .A(n22120), .X(n45387) );
  inv_x1_sg U42112 ( .A(n22188), .X(n45343) );
  inv_x1_sg U42113 ( .A(n22187), .X(n45349) );
  inv_x1_sg U42114 ( .A(n22184), .X(n45366) );
  inv_x1_sg U42115 ( .A(n22172), .X(n45345) );
  inv_x1_sg U42116 ( .A(n22167), .X(n45347) );
  inv_x1_sg U42117 ( .A(n22236), .X(n45298) );
  inv_x1_sg U42118 ( .A(n22235), .X(n45304) );
  inv_x1_sg U42119 ( .A(n22232), .X(n45321) );
  nand_x1_sg U42120 ( .A(n29248), .B(n29249), .X(n29185) );
  nand_x1_sg U42121 ( .A(out_L1[7]), .B(n29250), .X(n29249) );
  inv_x1_sg U42122 ( .A(n22220), .X(n45300) );
  inv_x1_sg U42123 ( .A(n22215), .X(n45296) );
  inv_x1_sg U42124 ( .A(n22214), .X(n45302) );
  inv_x1_sg U42125 ( .A(n22282), .X(n45259) );
  inv_x1_sg U42126 ( .A(n22283), .X(n45253) );
  inv_x1_sg U42127 ( .A(n22279), .X(n45276) );
  inv_x1_sg U42128 ( .A(n22267), .X(n45255) );
  inv_x1_sg U42129 ( .A(n22262), .X(n45257) );
  inv_x1_sg U42130 ( .A(n22331), .X(n45208) );
  inv_x1_sg U42131 ( .A(n22330), .X(n45214) );
  inv_x1_sg U42132 ( .A(n22327), .X(n45231) );
  nand_x1_sg U42133 ( .A(n29254), .B(n29255), .X(n29173) );
  nand_x1_sg U42134 ( .A(out_L1[5]), .B(n29256), .X(n29255) );
  inv_x1_sg U42135 ( .A(n22315), .X(n45210) );
  inv_x1_sg U42136 ( .A(n22310), .X(n45206) );
  inv_x1_sg U42137 ( .A(n22309), .X(n45212) );
  inv_x1_sg U42138 ( .A(n22378), .X(n45162) );
  inv_x1_sg U42139 ( .A(n22377), .X(n45168) );
  inv_x1_sg U42140 ( .A(n22374), .X(n45185) );
  inv_x1_sg U42141 ( .A(n22362), .X(n45164) );
  inv_x1_sg U42142 ( .A(n22357), .X(n45166) );
  inv_x1_sg U42143 ( .A(n22426), .X(n45117) );
  inv_x1_sg U42144 ( .A(n22425), .X(n45123) );
  inv_x1_sg U42145 ( .A(n22422), .X(n45140) );
  nand_x1_sg U42146 ( .A(n29260), .B(n29261), .X(n29161) );
  nand_x1_sg U42147 ( .A(out_L1[3]), .B(n29262), .X(n29261) );
  inv_x1_sg U42148 ( .A(n22410), .X(n45119) );
  inv_x1_sg U42149 ( .A(n22405), .X(n45115) );
  inv_x1_sg U42150 ( .A(n22404), .X(n45121) );
  inv_x1_sg U42151 ( .A(n22472), .X(n45070) );
  inv_x1_sg U42152 ( .A(n22471), .X(n45076) );
  inv_x1_sg U42153 ( .A(n22468), .X(n45093) );
  inv_x1_sg U42154 ( .A(n22456), .X(n45072) );
  inv_x1_sg U42155 ( .A(n22451), .X(n45074) );
  nand_x1_sg U42156 ( .A(n5377), .B(n28823), .X(n28822) );
  inv_x1_sg U42157 ( .A(n22518), .X(n45027) );
  nand_x1_sg U42158 ( .A(n5320), .B(n28380), .X(n28379) );
  inv_x1_sg U42159 ( .A(n22517), .X(n45033) );
  nand_x1_sg U42160 ( .A(n5149), .B(n22513), .X(n22512) );
  inv_x1_sg U42161 ( .A(n22514), .X(n45049) );
  nand_x1_sg U42162 ( .A(n5168), .B(n26964), .X(n26963) );
  nand_x1_sg U42163 ( .A(n5358), .B(n28635), .X(n28634) );
  inv_x1_sg U42164 ( .A(n22502), .X(n45029) );
  inv_x1_sg U42165 ( .A(n28133), .X(n41540) );
  nand_x1_sg U42166 ( .A(n5396), .B(n28994), .X(n28993) );
  inv_x1_sg U42167 ( .A(n22497), .X(n45025) );
  nand_x1_sg U42168 ( .A(n5339), .B(n28474), .X(n28473) );
  inv_x1_sg U42169 ( .A(n22496), .X(n45031) );
  nand_x1_sg U42170 ( .A(n46891), .B(n22789), .X(n22788) );
  nand_x1_sg U42171 ( .A(n22758), .B(n22759), .X(n6991) );
  nand_x1_sg U42172 ( .A(n22758), .B(n22759), .X(n39664) );
  nand_x1_sg U42173 ( .A(n22744), .B(n22745), .X(n39663) );
  nand_x1_sg U42174 ( .A(n22744), .B(n22745), .X(n7474) );
  nand_x1_sg U42175 ( .A(n47075), .B(n22732), .X(n22731) );
  nand_x1_sg U42176 ( .A(n22730), .B(n22731), .X(n39678) );
  nand_x1_sg U42177 ( .A(n22727), .B(n22728), .X(n7015) );
  nand_x1_sg U42178 ( .A(n22719), .B(n22720), .X(n22714) );
  nand_x1_sg U42179 ( .A(n47256), .B(n47233), .X(n23043) );
  nand_x1_sg U42180 ( .A(n47361), .B(n23009), .X(n23008) );
  nand_x1_sg U42181 ( .A(n23007), .B(n23008), .X(n39677) );
  nand_x1_sg U42182 ( .A(n23004), .B(n23005), .X(n7833) );
  nand_x1_sg U42183 ( .A(n47405), .B(n22999), .X(n7829) );
  nand_x1_sg U42184 ( .A(n22996), .B(n22997), .X(n22992) );
  nand_x1_sg U42185 ( .A(n47646), .B(n23289), .X(n23288) );
  nand_x1_sg U42186 ( .A(n23287), .B(n23288), .X(n39676) );
  nand_x1_sg U42187 ( .A(n23284), .B(n23285), .X(n8651) );
  nand_x1_sg U42188 ( .A(n47690), .B(n23279), .X(n8647) );
  nand_x1_sg U42189 ( .A(n23276), .B(n23277), .X(n23272) );
  nand_x1_sg U42190 ( .A(n38942), .B(n23264), .X(n23263) );
  nand_x1_sg U42191 ( .A(n47931), .B(n23568), .X(n23567) );
  nand_x1_sg U42192 ( .A(n23566), .B(n23567), .X(n39674) );
  nand_x1_sg U42193 ( .A(n23563), .B(n23564), .X(n9471) );
  nand_x1_sg U42194 ( .A(n47975), .B(n23558), .X(n9467) );
  nand_x1_sg U42195 ( .A(n23555), .B(n23556), .X(n23551) );
  nand_x1_sg U42196 ( .A(n48216), .B(n23847), .X(n23846) );
  nand_x1_sg U42197 ( .A(n23842), .B(n23843), .X(n10290) );
  nand_x1_sg U42198 ( .A(n48260), .B(n23837), .X(n10286) );
  nand_x1_sg U42199 ( .A(n23834), .B(n23835), .X(n23830) );
  nand_x1_sg U42200 ( .A(n48436), .B(n48413), .X(n24146) );
  nand_x1_sg U42201 ( .A(n48501), .B(n24126), .X(n24125) );
  nand_x1_sg U42202 ( .A(n24124), .B(n24125), .X(n39673) );
  nand_x1_sg U42203 ( .A(n24121), .B(n24122), .X(n11109) );
  nand_x1_sg U42204 ( .A(n48545), .B(n24116), .X(n11105) );
  nand_x1_sg U42205 ( .A(n24113), .B(n24114), .X(n24109) );
  nand_x1_sg U42206 ( .A(n48786), .B(n24405), .X(n24404) );
  nand_x1_sg U42207 ( .A(n24403), .B(n24404), .X(n39672) );
  nand_x1_sg U42208 ( .A(n24400), .B(n24401), .X(n11928) );
  nand_x1_sg U42209 ( .A(n48830), .B(n24395), .X(n11924) );
  nand_x1_sg U42210 ( .A(n24392), .B(n24393), .X(n24388) );
  nand_x1_sg U42211 ( .A(n49073), .B(n24683), .X(n24682) );
  nand_x1_sg U42212 ( .A(n24681), .B(n24682), .X(n39670) );
  nand_x1_sg U42213 ( .A(n24678), .B(n24679), .X(n12747) );
  nand_x1_sg U42214 ( .A(n49117), .B(n24673), .X(n12743) );
  nand_x1_sg U42215 ( .A(n24670), .B(n24671), .X(n24666) );
  nand_x1_sg U42216 ( .A(n49359), .B(n24962), .X(n24961) );
  nand_x1_sg U42217 ( .A(n24957), .B(n24958), .X(n13566) );
  nand_x1_sg U42218 ( .A(n49403), .B(n24952), .X(n13562) );
  nand_x1_sg U42219 ( .A(n24949), .B(n24950), .X(n24945) );
  nand_x1_sg U42220 ( .A(n49645), .B(n25241), .X(n25240) );
  nand_x1_sg U42221 ( .A(n25239), .B(n25240), .X(n39669) );
  nand_x1_sg U42222 ( .A(n25236), .B(n25237), .X(n14385) );
  nand_x1_sg U42223 ( .A(n49689), .B(n25231), .X(n14381) );
  nand_x1_sg U42224 ( .A(n25228), .B(n25229), .X(n25224) );
  nand_x1_sg U42225 ( .A(n49787), .B(n49766), .X(n25568) );
  nand_x1_sg U42226 ( .A(n49826), .B(n49803), .X(n25554) );
  nand_x1_sg U42227 ( .A(n49931), .B(n25520), .X(n25519) );
  nand_x1_sg U42228 ( .A(n25518), .B(n25519), .X(n39668) );
  nand_x1_sg U42229 ( .A(n25515), .B(n25516), .X(n15204) );
  nand_x1_sg U42230 ( .A(n49975), .B(n25510), .X(n15200) );
  nand_x1_sg U42231 ( .A(n25507), .B(n25508), .X(n25503) );
  nand_x1_sg U42232 ( .A(n50073), .B(n50052), .X(n25845) );
  nand_x1_sg U42233 ( .A(n50217), .B(n25797), .X(n25796) );
  nand_x1_sg U42234 ( .A(n25795), .B(n25796), .X(n39666) );
  nand_x1_sg U42235 ( .A(n25792), .B(n25793), .X(n16023) );
  nand_x1_sg U42236 ( .A(n50261), .B(n25787), .X(n16019) );
  nand_x1_sg U42237 ( .A(n25784), .B(n25785), .X(n25780) );
  nand_x1_sg U42238 ( .A(n50502), .B(n26136), .X(n26135) );
  nand_x1_sg U42239 ( .A(n26139), .B(n26149), .X(n16840) );
  inv_x1_sg U42240 ( .A(n16834), .X(n41526) );
  nand_x1_sg U42241 ( .A(n50791), .B(n26357), .X(n26356) );
  nand_x1_sg U42242 ( .A(n26352), .B(n26353), .X(n17661) );
  nand_x1_sg U42243 ( .A(n50835), .B(n26347), .X(n17657) );
  nand_x1_sg U42244 ( .A(n26344), .B(n26345), .X(n26340) );
  nand_x1_sg U42245 ( .A(n51078), .B(n26635), .X(n26634) );
  nand_x1_sg U42246 ( .A(n26630), .B(n26631), .X(n18482) );
  nand_x1_sg U42247 ( .A(n51122), .B(n26625), .X(n18478) );
  nand_x1_sg U42248 ( .A(n26622), .B(n26623), .X(n26618) );
  inv_x1_sg U42249 ( .A(n6848), .X(n46861) );
  nand_x1_sg U42250 ( .A(n7066), .B(n7067), .X(n6858) );
  nand_x1_sg U42251 ( .A(n6854), .B(n6852), .X(n7067) );
  nand_x1_sg U42252 ( .A(n7064), .B(n46883), .X(n6859) );
  nand_x1_sg U42253 ( .A(n6872), .B(n6871), .X(n6869) );
  nand_x1_sg U42254 ( .A(n46910), .B(n7119), .X(n7062) );
  nand_x1_sg U42255 ( .A(n7060), .B(n46930), .X(n6877) );
  nand_x1_sg U42256 ( .A(n6884), .B(n6883), .X(n6881) );
  nand_x1_sg U42257 ( .A(n46950), .B(n7173), .X(n7059) );
  nand_x1_sg U42258 ( .A(n7057), .B(n46978), .X(n6889) );
  nand_x1_sg U42259 ( .A(n7057), .B(n7058), .X(n6894) );
  nand_x1_sg U42260 ( .A(n46979), .B(n6888), .X(n7058) );
  nand_x1_sg U42261 ( .A(n7055), .B(n47001), .X(n6895) );
  nand_x1_sg U42262 ( .A(n7055), .B(n7056), .X(n6900) );
  nand_x1_sg U42263 ( .A(n47002), .B(n6894), .X(n7056) );
  nand_x1_sg U42264 ( .A(n7053), .B(n47015), .X(n6901) );
  nand_x1_sg U42265 ( .A(n7053), .B(n7054), .X(n6906) );
  nand_x1_sg U42266 ( .A(n47016), .B(n6900), .X(n7054) );
  nand_x1_sg U42267 ( .A(n7051), .B(n47041), .X(n6907) );
  nand_x1_sg U42268 ( .A(n7051), .B(n7052), .X(n6912) );
  nand_x1_sg U42269 ( .A(n47042), .B(n6906), .X(n7052) );
  nand_x1_sg U42270 ( .A(n7049), .B(n47069), .X(n6913) );
  nand_x1_sg U42271 ( .A(n7049), .B(n7050), .X(n6918) );
  nand_x1_sg U42272 ( .A(n47070), .B(n6912), .X(n7050) );
  nand_x1_sg U42273 ( .A(n7047), .B(n47091), .X(n6919) );
  nand_x1_sg U42274 ( .A(n7047), .B(n7048), .X(n6924) );
  nand_x1_sg U42275 ( .A(n47092), .B(n6918), .X(n7048) );
  nand_x1_sg U42276 ( .A(n7045), .B(n47115), .X(n6925) );
  inv_x1_sg U42277 ( .A(n7665), .X(n47154) );
  nand_x1_sg U42278 ( .A(n7884), .B(n7885), .X(n7675) );
  nand_x1_sg U42279 ( .A(n7671), .B(n7669), .X(n7885) );
  nand_x1_sg U42280 ( .A(n7882), .B(n47176), .X(n7676) );
  nand_x1_sg U42281 ( .A(n7689), .B(n7688), .X(n7686) );
  nand_x1_sg U42282 ( .A(n47203), .B(n7937), .X(n7880) );
  nand_x1_sg U42283 ( .A(n7878), .B(n47222), .X(n7694) );
  nand_x1_sg U42284 ( .A(n7701), .B(n7700), .X(n7698) );
  nand_x1_sg U42285 ( .A(n47241), .B(n7992), .X(n7877) );
  nand_x1_sg U42286 ( .A(n7875), .B(n47268), .X(n7706) );
  nand_x1_sg U42287 ( .A(n7875), .B(n7876), .X(n7711) );
  nand_x1_sg U42288 ( .A(n47269), .B(n7705), .X(n7876) );
  nand_x1_sg U42289 ( .A(n7873), .B(n47290), .X(n7712) );
  nand_x1_sg U42290 ( .A(n7873), .B(n7874), .X(n7717) );
  nand_x1_sg U42291 ( .A(n47291), .B(n7711), .X(n7874) );
  nand_x1_sg U42292 ( .A(n7871), .B(n47303), .X(n7718) );
  nand_x1_sg U42293 ( .A(n7871), .B(n7872), .X(n7723) );
  nand_x1_sg U42294 ( .A(n47304), .B(n7717), .X(n7872) );
  nand_x1_sg U42295 ( .A(n7869), .B(n47328), .X(n7724) );
  nand_x1_sg U42296 ( .A(n7869), .B(n7870), .X(n7729) );
  nand_x1_sg U42297 ( .A(n47329), .B(n7723), .X(n7870) );
  nand_x1_sg U42298 ( .A(n7867), .B(n47355), .X(n7730) );
  nand_x1_sg U42299 ( .A(n7867), .B(n7868), .X(n7735) );
  nand_x1_sg U42300 ( .A(n47356), .B(n7729), .X(n7868) );
  nand_x1_sg U42301 ( .A(n7865), .B(n47377), .X(n7736) );
  nand_x1_sg U42302 ( .A(n7865), .B(n7866), .X(n7741) );
  nand_x1_sg U42303 ( .A(n47378), .B(n7735), .X(n7866) );
  nand_x1_sg U42304 ( .A(n7863), .B(n47401), .X(n7742) );
  inv_x1_sg U42305 ( .A(n8483), .X(n47439) );
  nand_x1_sg U42306 ( .A(n8702), .B(n8703), .X(n8493) );
  nand_x1_sg U42307 ( .A(n8489), .B(n8487), .X(n8703) );
  nand_x1_sg U42308 ( .A(n8700), .B(n47461), .X(n8494) );
  nand_x1_sg U42309 ( .A(n8507), .B(n8506), .X(n8504) );
  nand_x1_sg U42310 ( .A(n47488), .B(n8755), .X(n8698) );
  nand_x1_sg U42311 ( .A(n8696), .B(n47507), .X(n8512) );
  nand_x1_sg U42312 ( .A(n8519), .B(n8518), .X(n8516) );
  nand_x1_sg U42313 ( .A(n47526), .B(n8810), .X(n8695) );
  nand_x1_sg U42314 ( .A(n8693), .B(n47553), .X(n8524) );
  nand_x1_sg U42315 ( .A(n8693), .B(n8694), .X(n8529) );
  nand_x1_sg U42316 ( .A(n47554), .B(n8523), .X(n8694) );
  nand_x1_sg U42317 ( .A(n8691), .B(n47575), .X(n8530) );
  nand_x1_sg U42318 ( .A(n8691), .B(n8692), .X(n8535) );
  nand_x1_sg U42319 ( .A(n47576), .B(n8529), .X(n8692) );
  nand_x1_sg U42320 ( .A(n8689), .B(n47588), .X(n8536) );
  nand_x1_sg U42321 ( .A(n8689), .B(n8690), .X(n8541) );
  nand_x1_sg U42322 ( .A(n47589), .B(n8535), .X(n8690) );
  nand_x1_sg U42323 ( .A(n8687), .B(n47613), .X(n8542) );
  nand_x1_sg U42324 ( .A(n8687), .B(n8688), .X(n8547) );
  nand_x1_sg U42325 ( .A(n47614), .B(n8541), .X(n8688) );
  nand_x1_sg U42326 ( .A(n8685), .B(n47640), .X(n8548) );
  nand_x1_sg U42327 ( .A(n8685), .B(n8686), .X(n8553) );
  nand_x1_sg U42328 ( .A(n47641), .B(n8547), .X(n8686) );
  nand_x1_sg U42329 ( .A(n8683), .B(n47662), .X(n8554) );
  nand_x1_sg U42330 ( .A(n8683), .B(n8684), .X(n8559) );
  nand_x1_sg U42331 ( .A(n47663), .B(n8553), .X(n8684) );
  nand_x1_sg U42332 ( .A(n8681), .B(n47686), .X(n8560) );
  inv_x1_sg U42333 ( .A(n9303), .X(n47724) );
  nand_x1_sg U42334 ( .A(n9522), .B(n9523), .X(n9313) );
  nand_x1_sg U42335 ( .A(n9309), .B(n9307), .X(n9523) );
  nand_x1_sg U42336 ( .A(n9520), .B(n47746), .X(n9314) );
  nand_x1_sg U42337 ( .A(n9327), .B(n9326), .X(n9324) );
  nand_x1_sg U42338 ( .A(n47773), .B(n9575), .X(n9518) );
  nand_x1_sg U42339 ( .A(n9516), .B(n47792), .X(n9332) );
  nand_x1_sg U42340 ( .A(n9339), .B(n9338), .X(n9336) );
  nand_x1_sg U42341 ( .A(n47811), .B(n9630), .X(n9515) );
  nand_x1_sg U42342 ( .A(n9513), .B(n47838), .X(n9344) );
  nand_x1_sg U42343 ( .A(n9513), .B(n9514), .X(n9349) );
  nand_x1_sg U42344 ( .A(n47839), .B(n9343), .X(n9514) );
  nand_x1_sg U42345 ( .A(n9511), .B(n47860), .X(n9350) );
  nand_x1_sg U42346 ( .A(n9511), .B(n9512), .X(n9355) );
  nand_x1_sg U42347 ( .A(n47861), .B(n9349), .X(n9512) );
  nand_x1_sg U42348 ( .A(n9509), .B(n47873), .X(n9356) );
  nand_x1_sg U42349 ( .A(n9509), .B(n9510), .X(n9361) );
  nand_x1_sg U42350 ( .A(n47874), .B(n9355), .X(n9510) );
  nand_x1_sg U42351 ( .A(n9507), .B(n47898), .X(n9362) );
  nand_x1_sg U42352 ( .A(n9507), .B(n9508), .X(n9367) );
  nand_x1_sg U42353 ( .A(n47899), .B(n9361), .X(n9508) );
  nand_x1_sg U42354 ( .A(n9505), .B(n47925), .X(n9368) );
  nand_x1_sg U42355 ( .A(n9505), .B(n9506), .X(n9373) );
  nand_x1_sg U42356 ( .A(n47926), .B(n9367), .X(n9506) );
  nand_x1_sg U42357 ( .A(n9503), .B(n47947), .X(n9374) );
  nand_x1_sg U42358 ( .A(n9503), .B(n9504), .X(n9379) );
  nand_x1_sg U42359 ( .A(n47948), .B(n9373), .X(n9504) );
  nand_x1_sg U42360 ( .A(n9501), .B(n47971), .X(n9380) );
  inv_x1_sg U42361 ( .A(n10122), .X(n48009) );
  nand_x1_sg U42362 ( .A(n10341), .B(n10342), .X(n10132) );
  nand_x1_sg U42363 ( .A(n10128), .B(n10126), .X(n10342) );
  nand_x1_sg U42364 ( .A(n10339), .B(n48031), .X(n10133) );
  nand_x1_sg U42365 ( .A(n10146), .B(n10145), .X(n10143) );
  nand_x1_sg U42366 ( .A(n48058), .B(n10394), .X(n10337) );
  nand_x1_sg U42367 ( .A(n10335), .B(n48077), .X(n10151) );
  nand_x1_sg U42368 ( .A(n10158), .B(n10157), .X(n10155) );
  nand_x1_sg U42369 ( .A(n48096), .B(n10449), .X(n10334) );
  nand_x1_sg U42370 ( .A(n10332), .B(n48123), .X(n10163) );
  nand_x1_sg U42371 ( .A(n10332), .B(n10333), .X(n10168) );
  nand_x1_sg U42372 ( .A(n48124), .B(n10162), .X(n10333) );
  nand_x1_sg U42373 ( .A(n10330), .B(n48145), .X(n10169) );
  nand_x1_sg U42374 ( .A(n10330), .B(n10331), .X(n10174) );
  nand_x1_sg U42375 ( .A(n48146), .B(n10168), .X(n10331) );
  nand_x1_sg U42376 ( .A(n10328), .B(n48158), .X(n10175) );
  nand_x1_sg U42377 ( .A(n10328), .B(n10329), .X(n10180) );
  nand_x1_sg U42378 ( .A(n48159), .B(n10174), .X(n10329) );
  nand_x1_sg U42379 ( .A(n10326), .B(n48183), .X(n10181) );
  nand_x1_sg U42380 ( .A(n10326), .B(n10327), .X(n10186) );
  nand_x1_sg U42381 ( .A(n48184), .B(n10180), .X(n10327) );
  nand_x1_sg U42382 ( .A(n10324), .B(n48210), .X(n10187) );
  nand_x1_sg U42383 ( .A(n10324), .B(n10325), .X(n10192) );
  nand_x1_sg U42384 ( .A(n48211), .B(n10186), .X(n10325) );
  nand_x1_sg U42385 ( .A(n10322), .B(n48232), .X(n10193) );
  nand_x1_sg U42386 ( .A(n10322), .B(n10323), .X(n10198) );
  nand_x1_sg U42387 ( .A(n48233), .B(n10192), .X(n10323) );
  nand_x1_sg U42388 ( .A(n10320), .B(n48256), .X(n10199) );
  inv_x1_sg U42389 ( .A(n10941), .X(n48294) );
  nand_x1_sg U42390 ( .A(n11160), .B(n11161), .X(n10951) );
  nand_x1_sg U42391 ( .A(n10947), .B(n10945), .X(n11161) );
  nand_x1_sg U42392 ( .A(n11158), .B(n48316), .X(n10952) );
  nand_x1_sg U42393 ( .A(n10965), .B(n10964), .X(n10962) );
  nand_x1_sg U42394 ( .A(n48343), .B(n11213), .X(n11156) );
  nand_x1_sg U42395 ( .A(n11154), .B(n48362), .X(n10970) );
  nand_x1_sg U42396 ( .A(n10977), .B(n10976), .X(n10974) );
  nand_x1_sg U42397 ( .A(n48381), .B(n11268), .X(n11153) );
  nand_x1_sg U42398 ( .A(n11151), .B(n48408), .X(n10982) );
  nand_x1_sg U42399 ( .A(n11151), .B(n11152), .X(n10987) );
  nand_x1_sg U42400 ( .A(n48409), .B(n10981), .X(n11152) );
  nand_x1_sg U42401 ( .A(n11149), .B(n48430), .X(n10988) );
  nand_x1_sg U42402 ( .A(n11149), .B(n11150), .X(n10993) );
  nand_x1_sg U42403 ( .A(n48431), .B(n10987), .X(n11150) );
  nand_x1_sg U42404 ( .A(n11147), .B(n48443), .X(n10994) );
  nand_x1_sg U42405 ( .A(n11147), .B(n11148), .X(n10999) );
  nand_x1_sg U42406 ( .A(n48444), .B(n10993), .X(n11148) );
  nand_x1_sg U42407 ( .A(n11145), .B(n48468), .X(n11000) );
  nand_x1_sg U42408 ( .A(n11145), .B(n11146), .X(n11005) );
  nand_x1_sg U42409 ( .A(n48469), .B(n10999), .X(n11146) );
  nand_x1_sg U42410 ( .A(n11143), .B(n48495), .X(n11006) );
  nand_x1_sg U42411 ( .A(n11143), .B(n11144), .X(n11011) );
  nand_x1_sg U42412 ( .A(n48496), .B(n11005), .X(n11144) );
  nand_x1_sg U42413 ( .A(n11141), .B(n48517), .X(n11012) );
  nand_x1_sg U42414 ( .A(n11141), .B(n11142), .X(n11017) );
  nand_x1_sg U42415 ( .A(n48518), .B(n11011), .X(n11142) );
  nand_x1_sg U42416 ( .A(n11139), .B(n48541), .X(n11018) );
  inv_x1_sg U42417 ( .A(n11760), .X(n48579) );
  nand_x1_sg U42418 ( .A(n11979), .B(n11980), .X(n11770) );
  nand_x1_sg U42419 ( .A(n11766), .B(n11764), .X(n11980) );
  nand_x1_sg U42420 ( .A(n11977), .B(n48601), .X(n11771) );
  nand_x1_sg U42421 ( .A(n11784), .B(n11783), .X(n11781) );
  nand_x1_sg U42422 ( .A(n48628), .B(n12032), .X(n11975) );
  nand_x1_sg U42423 ( .A(n11973), .B(n48647), .X(n11789) );
  nand_x1_sg U42424 ( .A(n11796), .B(n11795), .X(n11793) );
  nand_x1_sg U42425 ( .A(n48666), .B(n12087), .X(n11972) );
  nand_x1_sg U42426 ( .A(n11970), .B(n48693), .X(n11801) );
  nand_x1_sg U42427 ( .A(n11970), .B(n11971), .X(n11806) );
  nand_x1_sg U42428 ( .A(n48694), .B(n11800), .X(n11971) );
  nand_x1_sg U42429 ( .A(n11968), .B(n48715), .X(n11807) );
  nand_x1_sg U42430 ( .A(n11968), .B(n11969), .X(n11812) );
  nand_x1_sg U42431 ( .A(n48716), .B(n11806), .X(n11969) );
  nand_x1_sg U42432 ( .A(n11966), .B(n48728), .X(n11813) );
  nand_x1_sg U42433 ( .A(n11966), .B(n11967), .X(n11818) );
  nand_x1_sg U42434 ( .A(n48729), .B(n11812), .X(n11967) );
  nand_x1_sg U42435 ( .A(n11964), .B(n48753), .X(n11819) );
  nand_x1_sg U42436 ( .A(n11964), .B(n11965), .X(n11824) );
  nand_x1_sg U42437 ( .A(n48754), .B(n11818), .X(n11965) );
  nand_x1_sg U42438 ( .A(n11962), .B(n48780), .X(n11825) );
  nand_x1_sg U42439 ( .A(n11962), .B(n11963), .X(n11830) );
  nand_x1_sg U42440 ( .A(n48781), .B(n11824), .X(n11963) );
  nand_x1_sg U42441 ( .A(n11960), .B(n48802), .X(n11831) );
  nand_x1_sg U42442 ( .A(n11960), .B(n11961), .X(n11836) );
  nand_x1_sg U42443 ( .A(n48803), .B(n11830), .X(n11961) );
  nand_x1_sg U42444 ( .A(n11958), .B(n48826), .X(n11837) );
  inv_x1_sg U42445 ( .A(n12579), .X(n48865) );
  nand_x1_sg U42446 ( .A(n12798), .B(n12799), .X(n12589) );
  nand_x1_sg U42447 ( .A(n12585), .B(n12583), .X(n12799) );
  nand_x1_sg U42448 ( .A(n12796), .B(n48887), .X(n12590) );
  nand_x1_sg U42449 ( .A(n12603), .B(n12602), .X(n12600) );
  nand_x1_sg U42450 ( .A(n48914), .B(n12851), .X(n12794) );
  nand_x1_sg U42451 ( .A(n12792), .B(n48933), .X(n12608) );
  nand_x1_sg U42452 ( .A(n12615), .B(n12614), .X(n12612) );
  nand_x1_sg U42453 ( .A(n48952), .B(n12906), .X(n12791) );
  nand_x1_sg U42454 ( .A(n12789), .B(n48979), .X(n12620) );
  nand_x1_sg U42455 ( .A(n12789), .B(n12790), .X(n12625) );
  nand_x1_sg U42456 ( .A(n48980), .B(n12619), .X(n12790) );
  nand_x1_sg U42457 ( .A(n12787), .B(n49001), .X(n12626) );
  nand_x1_sg U42458 ( .A(n12787), .B(n12788), .X(n12631) );
  nand_x1_sg U42459 ( .A(n49002), .B(n12625), .X(n12788) );
  nand_x1_sg U42460 ( .A(n12785), .B(n49014), .X(n12632) );
  nand_x1_sg U42461 ( .A(n12785), .B(n12786), .X(n12637) );
  nand_x1_sg U42462 ( .A(n49015), .B(n12631), .X(n12786) );
  nand_x1_sg U42463 ( .A(n12783), .B(n49039), .X(n12638) );
  nand_x1_sg U42464 ( .A(n12783), .B(n12784), .X(n12643) );
  nand_x1_sg U42465 ( .A(n49040), .B(n12637), .X(n12784) );
  nand_x1_sg U42466 ( .A(n12781), .B(n49067), .X(n12644) );
  nand_x1_sg U42467 ( .A(n12781), .B(n12782), .X(n12649) );
  nand_x1_sg U42468 ( .A(n49068), .B(n12643), .X(n12782) );
  nand_x1_sg U42469 ( .A(n12779), .B(n49089), .X(n12650) );
  nand_x1_sg U42470 ( .A(n12779), .B(n12780), .X(n12655) );
  nand_x1_sg U42471 ( .A(n49090), .B(n12649), .X(n12780) );
  nand_x1_sg U42472 ( .A(n12777), .B(n49113), .X(n12656) );
  inv_x1_sg U42473 ( .A(n13398), .X(n49152) );
  nand_x1_sg U42474 ( .A(n13617), .B(n13618), .X(n13408) );
  nand_x1_sg U42475 ( .A(n13404), .B(n13402), .X(n13618) );
  nand_x1_sg U42476 ( .A(n13615), .B(n49174), .X(n13409) );
  nand_x1_sg U42477 ( .A(n13422), .B(n13421), .X(n13419) );
  nand_x1_sg U42478 ( .A(n49201), .B(n13670), .X(n13613) );
  nand_x1_sg U42479 ( .A(n13611), .B(n49220), .X(n13427) );
  nand_x1_sg U42480 ( .A(n13434), .B(n13433), .X(n13431) );
  nand_x1_sg U42481 ( .A(n49239), .B(n13725), .X(n13610) );
  nand_x1_sg U42482 ( .A(n13608), .B(n49266), .X(n13439) );
  nand_x1_sg U42483 ( .A(n13608), .B(n13609), .X(n13444) );
  nand_x1_sg U42484 ( .A(n49267), .B(n13438), .X(n13609) );
  nand_x1_sg U42485 ( .A(n13606), .B(n49288), .X(n13445) );
  nand_x1_sg U42486 ( .A(n13606), .B(n13607), .X(n13450) );
  nand_x1_sg U42487 ( .A(n49289), .B(n13444), .X(n13607) );
  nand_x1_sg U42488 ( .A(n13604), .B(n49301), .X(n13451) );
  nand_x1_sg U42489 ( .A(n13604), .B(n13605), .X(n13456) );
  nand_x1_sg U42490 ( .A(n49302), .B(n13450), .X(n13605) );
  nand_x1_sg U42491 ( .A(n13602), .B(n49326), .X(n13457) );
  nand_x1_sg U42492 ( .A(n13602), .B(n13603), .X(n13462) );
  nand_x1_sg U42493 ( .A(n49327), .B(n13456), .X(n13603) );
  nand_x1_sg U42494 ( .A(n13600), .B(n49353), .X(n13463) );
  nand_x1_sg U42495 ( .A(n13600), .B(n13601), .X(n13468) );
  nand_x1_sg U42496 ( .A(n49354), .B(n13462), .X(n13601) );
  nand_x1_sg U42497 ( .A(n13598), .B(n49375), .X(n13469) );
  nand_x1_sg U42498 ( .A(n13598), .B(n13599), .X(n13474) );
  nand_x1_sg U42499 ( .A(n49376), .B(n13468), .X(n13599) );
  nand_x1_sg U42500 ( .A(n13596), .B(n49399), .X(n13475) );
  inv_x1_sg U42501 ( .A(n14217), .X(n49438) );
  nand_x1_sg U42502 ( .A(n14436), .B(n14437), .X(n14227) );
  nand_x1_sg U42503 ( .A(n14223), .B(n14221), .X(n14437) );
  nand_x1_sg U42504 ( .A(n14434), .B(n49460), .X(n14228) );
  nand_x1_sg U42505 ( .A(n14241), .B(n14240), .X(n14238) );
  nand_x1_sg U42506 ( .A(n49487), .B(n14489), .X(n14432) );
  nand_x1_sg U42507 ( .A(n14430), .B(n49506), .X(n14246) );
  nand_x1_sg U42508 ( .A(n14253), .B(n14252), .X(n14250) );
  nand_x1_sg U42509 ( .A(n49525), .B(n14544), .X(n14429) );
  nand_x1_sg U42510 ( .A(n14427), .B(n49552), .X(n14258) );
  nand_x1_sg U42511 ( .A(n14427), .B(n14428), .X(n14263) );
  nand_x1_sg U42512 ( .A(n49553), .B(n14257), .X(n14428) );
  nand_x1_sg U42513 ( .A(n14425), .B(n49574), .X(n14264) );
  nand_x1_sg U42514 ( .A(n14425), .B(n14426), .X(n14269) );
  nand_x1_sg U42515 ( .A(n49575), .B(n14263), .X(n14426) );
  nand_x1_sg U42516 ( .A(n14423), .B(n49587), .X(n14270) );
  nand_x1_sg U42517 ( .A(n14423), .B(n14424), .X(n14275) );
  nand_x1_sg U42518 ( .A(n49588), .B(n14269), .X(n14424) );
  nand_x1_sg U42519 ( .A(n14421), .B(n49612), .X(n14276) );
  nand_x1_sg U42520 ( .A(n14421), .B(n14422), .X(n14281) );
  nand_x1_sg U42521 ( .A(n49613), .B(n14275), .X(n14422) );
  nand_x1_sg U42522 ( .A(n14419), .B(n49639), .X(n14282) );
  nand_x1_sg U42523 ( .A(n14419), .B(n14420), .X(n14287) );
  nand_x1_sg U42524 ( .A(n49640), .B(n14281), .X(n14420) );
  nand_x1_sg U42525 ( .A(n14417), .B(n49661), .X(n14288) );
  nand_x1_sg U42526 ( .A(n14417), .B(n14418), .X(n14293) );
  nand_x1_sg U42527 ( .A(n49662), .B(n14287), .X(n14418) );
  nand_x1_sg U42528 ( .A(n14415), .B(n49685), .X(n14294) );
  inv_x1_sg U42529 ( .A(n15036), .X(n49723) );
  nand_x1_sg U42530 ( .A(n15255), .B(n15256), .X(n15046) );
  nand_x1_sg U42531 ( .A(n15042), .B(n15040), .X(n15256) );
  nand_x1_sg U42532 ( .A(n15253), .B(n49745), .X(n15047) );
  nand_x1_sg U42533 ( .A(n15060), .B(n15059), .X(n15057) );
  nand_x1_sg U42534 ( .A(n49773), .B(n15308), .X(n15251) );
  nand_x1_sg U42535 ( .A(n15249), .B(n49792), .X(n15065) );
  nand_x1_sg U42536 ( .A(n15072), .B(n15071), .X(n15069) );
  nand_x1_sg U42537 ( .A(n49811), .B(n15363), .X(n15248) );
  nand_x1_sg U42538 ( .A(n15246), .B(n49838), .X(n15077) );
  nand_x1_sg U42539 ( .A(n15246), .B(n15247), .X(n15082) );
  nand_x1_sg U42540 ( .A(n49839), .B(n15076), .X(n15247) );
  nand_x1_sg U42541 ( .A(n15244), .B(n49860), .X(n15083) );
  nand_x1_sg U42542 ( .A(n15244), .B(n15245), .X(n15088) );
  nand_x1_sg U42543 ( .A(n49861), .B(n15082), .X(n15245) );
  nand_x1_sg U42544 ( .A(n15242), .B(n49873), .X(n15089) );
  nand_x1_sg U42545 ( .A(n15242), .B(n15243), .X(n15094) );
  nand_x1_sg U42546 ( .A(n49874), .B(n15088), .X(n15243) );
  nand_x1_sg U42547 ( .A(n15240), .B(n49898), .X(n15095) );
  nand_x1_sg U42548 ( .A(n15240), .B(n15241), .X(n15100) );
  nand_x1_sg U42549 ( .A(n49899), .B(n15094), .X(n15241) );
  nand_x1_sg U42550 ( .A(n15238), .B(n49925), .X(n15101) );
  nand_x1_sg U42551 ( .A(n15238), .B(n15239), .X(n15106) );
  nand_x1_sg U42552 ( .A(n49926), .B(n15100), .X(n15239) );
  nand_x1_sg U42553 ( .A(n15236), .B(n49947), .X(n15107) );
  nand_x1_sg U42554 ( .A(n15236), .B(n15237), .X(n15112) );
  nand_x1_sg U42555 ( .A(n49948), .B(n15106), .X(n15237) );
  nand_x1_sg U42556 ( .A(n15234), .B(n49971), .X(n15113) );
  inv_x1_sg U42557 ( .A(n15855), .X(n50010) );
  nand_x1_sg U42558 ( .A(n16074), .B(n16075), .X(n15865) );
  nand_x1_sg U42559 ( .A(n15861), .B(n15859), .X(n16075) );
  nand_x1_sg U42560 ( .A(n16072), .B(n50032), .X(n15866) );
  nand_x1_sg U42561 ( .A(n15879), .B(n15878), .X(n15876) );
  nand_x1_sg U42562 ( .A(n50059), .B(n16127), .X(n16070) );
  nand_x1_sg U42563 ( .A(n16068), .B(n50078), .X(n15884) );
  nand_x1_sg U42564 ( .A(n15891), .B(n15890), .X(n15888) );
  nand_x1_sg U42565 ( .A(n50097), .B(n16182), .X(n16067) );
  nand_x1_sg U42566 ( .A(n16065), .B(n50124), .X(n15896) );
  nand_x1_sg U42567 ( .A(n16065), .B(n16066), .X(n15901) );
  nand_x1_sg U42568 ( .A(n50125), .B(n15895), .X(n16066) );
  nand_x1_sg U42569 ( .A(n16063), .B(n50146), .X(n15902) );
  nand_x1_sg U42570 ( .A(n16063), .B(n16064), .X(n15907) );
  nand_x1_sg U42571 ( .A(n50147), .B(n15901), .X(n16064) );
  nand_x1_sg U42572 ( .A(n16061), .B(n50159), .X(n15908) );
  nand_x1_sg U42573 ( .A(n16061), .B(n16062), .X(n15913) );
  nand_x1_sg U42574 ( .A(n50160), .B(n15907), .X(n16062) );
  nand_x1_sg U42575 ( .A(n16059), .B(n50184), .X(n15914) );
  nand_x1_sg U42576 ( .A(n16059), .B(n16060), .X(n15919) );
  nand_x1_sg U42577 ( .A(n50185), .B(n15913), .X(n16060) );
  nand_x1_sg U42578 ( .A(n16057), .B(n50211), .X(n15920) );
  nand_x1_sg U42579 ( .A(n16057), .B(n16058), .X(n15925) );
  nand_x1_sg U42580 ( .A(n50212), .B(n15919), .X(n16058) );
  nand_x1_sg U42581 ( .A(n16055), .B(n50233), .X(n15926) );
  nand_x1_sg U42582 ( .A(n16055), .B(n16056), .X(n15931) );
  nand_x1_sg U42583 ( .A(n50234), .B(n15925), .X(n16056) );
  nand_x1_sg U42584 ( .A(n16053), .B(n50257), .X(n15932) );
  inv_x1_sg U42585 ( .A(n16672), .X(n50294) );
  inv_x1_sg U42586 ( .A(n16678), .X(n50306) );
  nand_x1_sg U42587 ( .A(n16893), .B(n16894), .X(n16682) );
  nand_x1_sg U42588 ( .A(n16891), .B(n50317), .X(n16683) );
  nand_x1_sg U42589 ( .A(n16696), .B(n16695), .X(n16693) );
  nand_x1_sg U42590 ( .A(n50344), .B(n16944), .X(n16889) );
  nand_x1_sg U42591 ( .A(n16887), .B(n50363), .X(n16701) );
  nand_x1_sg U42592 ( .A(n16708), .B(n16707), .X(n16705) );
  nand_x1_sg U42593 ( .A(n50382), .B(n16998), .X(n16886) );
  nand_x1_sg U42594 ( .A(n16884), .B(n50409), .X(n16713) );
  nand_x1_sg U42595 ( .A(n16884), .B(n16885), .X(n16718) );
  nand_x1_sg U42596 ( .A(n50410), .B(n16712), .X(n16885) );
  nand_x1_sg U42597 ( .A(n16882), .B(n50431), .X(n16719) );
  nand_x1_sg U42598 ( .A(n16882), .B(n16883), .X(n16724) );
  nand_x1_sg U42599 ( .A(n50432), .B(n16718), .X(n16883) );
  nand_x1_sg U42600 ( .A(n16880), .B(n50444), .X(n16725) );
  nand_x1_sg U42601 ( .A(n16880), .B(n16881), .X(n16730) );
  nand_x1_sg U42602 ( .A(n50445), .B(n16724), .X(n16881) );
  nand_x1_sg U42603 ( .A(n16878), .B(n50469), .X(n16731) );
  nand_x1_sg U42604 ( .A(n16878), .B(n16879), .X(n16736) );
  nand_x1_sg U42605 ( .A(n50470), .B(n16730), .X(n16879) );
  nand_x1_sg U42606 ( .A(n16876), .B(n50496), .X(n16737) );
  nand_x1_sg U42607 ( .A(n16876), .B(n16877), .X(n16742) );
  nand_x1_sg U42608 ( .A(n50497), .B(n16736), .X(n16877) );
  nand_x1_sg U42609 ( .A(n16874), .B(n50518), .X(n16743) );
  nand_x1_sg U42610 ( .A(n16874), .B(n16875), .X(n16748) );
  nand_x1_sg U42611 ( .A(n50519), .B(n16742), .X(n16875) );
  nand_x1_sg U42612 ( .A(n16872), .B(n50542), .X(n16749) );
  inv_x1_sg U42613 ( .A(n17493), .X(n50584) );
  nand_x1_sg U42614 ( .A(n17712), .B(n17713), .X(n17503) );
  nand_x1_sg U42615 ( .A(n17499), .B(n17497), .X(n17713) );
  nand_x1_sg U42616 ( .A(n17710), .B(n50606), .X(n17504) );
  nand_x1_sg U42617 ( .A(n17517), .B(n17516), .X(n17514) );
  nand_x1_sg U42618 ( .A(n50633), .B(n17765), .X(n17708) );
  nand_x1_sg U42619 ( .A(n17706), .B(n50652), .X(n17522) );
  nand_x1_sg U42620 ( .A(n17529), .B(n17528), .X(n17526) );
  nand_x1_sg U42621 ( .A(n50671), .B(n17820), .X(n17705) );
  nand_x1_sg U42622 ( .A(n17703), .B(n50698), .X(n17534) );
  nand_x1_sg U42623 ( .A(n17703), .B(n17704), .X(n17539) );
  nand_x1_sg U42624 ( .A(n50699), .B(n17533), .X(n17704) );
  nand_x1_sg U42625 ( .A(n17701), .B(n50720), .X(n17540) );
  nand_x1_sg U42626 ( .A(n17701), .B(n17702), .X(n17545) );
  nand_x1_sg U42627 ( .A(n50721), .B(n17539), .X(n17702) );
  nand_x1_sg U42628 ( .A(n17699), .B(n50733), .X(n17546) );
  nand_x1_sg U42629 ( .A(n17699), .B(n17700), .X(n17551) );
  nand_x1_sg U42630 ( .A(n50734), .B(n17545), .X(n17700) );
  nand_x1_sg U42631 ( .A(n17697), .B(n50758), .X(n17552) );
  nand_x1_sg U42632 ( .A(n17697), .B(n17698), .X(n17557) );
  nand_x1_sg U42633 ( .A(n50759), .B(n17551), .X(n17698) );
  nand_x1_sg U42634 ( .A(n17695), .B(n50785), .X(n17558) );
  nand_x1_sg U42635 ( .A(n17695), .B(n17696), .X(n17563) );
  nand_x1_sg U42636 ( .A(n50786), .B(n17557), .X(n17696) );
  nand_x1_sg U42637 ( .A(n17693), .B(n50807), .X(n17564) );
  nand_x1_sg U42638 ( .A(n17693), .B(n17694), .X(n17569) );
  nand_x1_sg U42639 ( .A(n50808), .B(n17563), .X(n17694) );
  nand_x1_sg U42640 ( .A(n17691), .B(n50831), .X(n17570) );
  inv_x1_sg U42641 ( .A(n18314), .X(n50871) );
  nand_x1_sg U42642 ( .A(n18533), .B(n18534), .X(n18324) );
  nand_x1_sg U42643 ( .A(n18320), .B(n18318), .X(n18534) );
  nand_x1_sg U42644 ( .A(n18531), .B(n50893), .X(n18325) );
  nand_x1_sg U42645 ( .A(n18338), .B(n18337), .X(n18335) );
  nand_x1_sg U42646 ( .A(n50920), .B(n18586), .X(n18529) );
  nand_x1_sg U42647 ( .A(n18527), .B(n50939), .X(n18343) );
  nand_x1_sg U42648 ( .A(n18350), .B(n18349), .X(n18347) );
  nand_x1_sg U42649 ( .A(n50958), .B(n18641), .X(n18526) );
  nand_x1_sg U42650 ( .A(n18524), .B(n50985), .X(n18355) );
  nand_x1_sg U42651 ( .A(n18524), .B(n18525), .X(n18360) );
  nand_x1_sg U42652 ( .A(n50986), .B(n18354), .X(n18525) );
  nand_x1_sg U42653 ( .A(n18522), .B(n51007), .X(n18361) );
  nand_x1_sg U42654 ( .A(n18522), .B(n18523), .X(n18366) );
  nand_x1_sg U42655 ( .A(n51008), .B(n18360), .X(n18523) );
  nand_x1_sg U42656 ( .A(n18520), .B(n51020), .X(n18367) );
  nand_x1_sg U42657 ( .A(n18520), .B(n18521), .X(n18372) );
  nand_x1_sg U42658 ( .A(n51021), .B(n18366), .X(n18521) );
  nand_x1_sg U42659 ( .A(n18518), .B(n51045), .X(n18373) );
  nand_x1_sg U42660 ( .A(n18518), .B(n18519), .X(n18378) );
  nand_x1_sg U42661 ( .A(n51046), .B(n18372), .X(n18519) );
  nand_x1_sg U42662 ( .A(n18516), .B(n51072), .X(n18379) );
  nand_x1_sg U42663 ( .A(n18516), .B(n18517), .X(n18384) );
  nand_x1_sg U42664 ( .A(n51073), .B(n18378), .X(n18517) );
  nand_x1_sg U42665 ( .A(n18514), .B(n51094), .X(n18385) );
  nand_x1_sg U42666 ( .A(n18514), .B(n18515), .X(n18390) );
  nand_x1_sg U42667 ( .A(n51095), .B(n18384), .X(n18515) );
  nand_x1_sg U42668 ( .A(n18512), .B(n51118), .X(n18391) );
  nand_x1_sg U42669 ( .A(n45788), .B(n26826), .X(n26791) );
  nand_x1_sg U42670 ( .A(n45785), .B(n28527), .X(n26790) );
  nand_x1_sg U42671 ( .A(n45796), .B(n26802), .X(n26796) );
  nand_x1_sg U42672 ( .A(n45786), .B(n28524), .X(n26784) );
  nand_x1_sg U42673 ( .A(n28533), .B(n45783), .X(n26785) );
  nand_x1_sg U42674 ( .A(n28536), .B(n28535), .X(n28533) );
  nand_x2_sg U42675 ( .A(n26759), .B(n26760), .X(n5940) );
  nand_x1_sg U42676 ( .A(n45787), .B(n28521), .X(n26827) );
  nand_x1_sg U42677 ( .A(n45784), .B(n28530), .X(n28519) );
  nand_x1_sg U42678 ( .A(n28729), .B(n45744), .X(n21751) );
  nand_x1_sg U42679 ( .A(n27079), .B(n45750), .X(n21752) );
  nand_x1_sg U42680 ( .A(n27055), .B(n45766), .X(n21763) );
  nand_x1_sg U42681 ( .A(n45740), .B(n28735), .X(n21746) );
  nand_x1_sg U42682 ( .A(n28726), .B(n45746), .X(n21745) );
  nand_x2_sg U42683 ( .A(n21725), .B(n21726), .X(n5896) );
  nand_x1_sg U42684 ( .A(n28732), .B(n45742), .X(n21767) );
  nand_x1_sg U42685 ( .A(n27082), .B(n45748), .X(n21766) );
  nand_x1_sg U42686 ( .A(n28908), .B(n45701), .X(n21798) );
  nand_x1_sg U42687 ( .A(n27309), .B(n45707), .X(n21799) );
  nand_x1_sg U42688 ( .A(n27049), .B(n45723), .X(n21810) );
  nand_x1_sg U42689 ( .A(n28914), .B(n45697), .X(n21793) );
  nand_x1_sg U42690 ( .A(n28720), .B(n45703), .X(n21792) );
  nand_x2_sg U42691 ( .A(n21772), .B(n21773), .X(n5919) );
  nand_x1_sg U42692 ( .A(n28911), .B(n45699), .X(n21814) );
  nand_x1_sg U42693 ( .A(n27312), .B(n45705), .X(n21813) );
  nand_x1_sg U42694 ( .A(n27522), .B(n45663), .X(n21846) );
  nand_x1_sg U42695 ( .A(n28902), .B(n45657), .X(n21845) );
  nand_x1_sg U42696 ( .A(n27043), .B(n45680), .X(n21857) );
  nand_x1_sg U42697 ( .A(n28714), .B(n45659), .X(n21839) );
  nand_x1_sg U42698 ( .A(n29083), .B(n45653), .X(n21840) );
  nand_x2_sg U42699 ( .A(n21819), .B(n21820), .X(n5784) );
  nand_x1_sg U42700 ( .A(n27525), .B(n45661), .X(n21860) );
  nand_x1_sg U42701 ( .A(n29080), .B(n45655), .X(n21861) );
  nand_x1_sg U42702 ( .A(n28896), .B(n45613), .X(n21891) );
  nand_x1_sg U42703 ( .A(n27716), .B(n45619), .X(n21892) );
  nand_x1_sg U42704 ( .A(n27037), .B(n45636), .X(n21903) );
  nand_x1_sg U42705 ( .A(n28708), .B(n45615), .X(n21886) );
  nand_x2_sg U42706 ( .A(n21866), .B(n21867), .X(n5855) );
  nand_x1_sg U42707 ( .A(n29073), .B(n45611), .X(n21907) );
  nand_x1_sg U42708 ( .A(n27719), .B(n45617), .X(n21906) );
  nand_x1_sg U42709 ( .A(n28890), .B(n45569), .X(n21938) );
  nand_x1_sg U42710 ( .A(n27893), .B(n45575), .X(n21939) );
  nand_x1_sg U42711 ( .A(n27031), .B(n45592), .X(n21950) );
  nand_x1_sg U42712 ( .A(n29218), .B(n45565), .X(n21933) );
  nand_x1_sg U42713 ( .A(n28702), .B(n45571), .X(n21932) );
  nand_x2_sg U42714 ( .A(n21912), .B(n21913), .X(n5848) );
  nand_x1_sg U42715 ( .A(n29067), .B(n45567), .X(n21954) );
  nand_x1_sg U42716 ( .A(n27896), .B(n45573), .X(n21953) );
  nand_x1_sg U42717 ( .A(n28884), .B(n45524), .X(n21984) );
  nand_x1_sg U42718 ( .A(n28055), .B(n45530), .X(n21985) );
  nand_x1_sg U42719 ( .A(n27025), .B(n45547), .X(n21996) );
  nand_x1_sg U42720 ( .A(n28696), .B(n45526), .X(n21979) );
  nand_x2_sg U42721 ( .A(n21959), .B(n21960), .X(n5910) );
  nand_x1_sg U42722 ( .A(n29060), .B(n45522), .X(n22000) );
  nand_x1_sg U42723 ( .A(n28058), .B(n45528), .X(n21999) );
  nand_x1_sg U42724 ( .A(n28878), .B(n45480), .X(n22031) );
  nand_x1_sg U42725 ( .A(n28190), .B(n45486), .X(n22032) );
  nand_x1_sg U42726 ( .A(n27019), .B(n45503), .X(n22043) );
  nand_x1_sg U42727 ( .A(n29206), .B(n45476), .X(n22026) );
  nand_x1_sg U42728 ( .A(n28690), .B(n45482), .X(n22025) );
  nand_x2_sg U42729 ( .A(n22005), .B(n22006), .X(n5871) );
  nand_x1_sg U42730 ( .A(n29054), .B(n45478), .X(n22047) );
  nand_x1_sg U42731 ( .A(n28193), .B(n45484), .X(n22046) );
  nand_x1_sg U42732 ( .A(n28872), .B(n45435), .X(n22077) );
  nand_x1_sg U42733 ( .A(n28319), .B(n45441), .X(n22078) );
  nand_x1_sg U42734 ( .A(n27013), .B(n45455), .X(n22089) );
  nand_x1_sg U42735 ( .A(n28684), .B(n45437), .X(n22072) );
  nand_x2_sg U42736 ( .A(n22052), .B(n22053), .X(n5889) );
  nand_x1_sg U42737 ( .A(n29047), .B(n45433), .X(n22093) );
  nand_x1_sg U42738 ( .A(n28322), .B(n45439), .X(n22092) );
  nand_x1_sg U42739 ( .A(n28423), .B(n45396), .X(n22126) );
  nand_x1_sg U42740 ( .A(n28866), .B(n45390), .X(n22125) );
  nand_x1_sg U42741 ( .A(n27007), .B(n45411), .X(n22137) );
  nand_x1_sg U42742 ( .A(n28678), .B(n45392), .X(n22119) );
  nand_x1_sg U42743 ( .A(n29194), .B(n45386), .X(n22120) );
  nand_x2_sg U42744 ( .A(n22098), .B(n22099), .X(n5794) );
  nand_x1_sg U42745 ( .A(n28426), .B(n45394), .X(n22140) );
  nand_x1_sg U42746 ( .A(n29041), .B(n45388), .X(n22141) );
  nand_x1_sg U42747 ( .A(n28860), .B(n45344), .X(n22172) );
  nand_x1_sg U42748 ( .A(n28417), .B(n45350), .X(n22173) );
  nand_x1_sg U42749 ( .A(n27001), .B(n45365), .X(n22184) );
  nand_x1_sg U42750 ( .A(n28672), .B(n45346), .X(n22167) );
  nand_x2_sg U42751 ( .A(n22146), .B(n22147), .X(n5817) );
  nand_x1_sg U42752 ( .A(n29034), .B(n45342), .X(n22188) );
  nand_x1_sg U42753 ( .A(n28511), .B(n45348), .X(n22187) );
  nand_x1_sg U42754 ( .A(n28854), .B(n45299), .X(n22220) );
  nand_x1_sg U42755 ( .A(n28411), .B(n45305), .X(n22221) );
  nand_x1_sg U42756 ( .A(n26995), .B(n45320), .X(n22232) );
  nand_x1_sg U42757 ( .A(n29182), .B(n45295), .X(n22215) );
  nand_x1_sg U42758 ( .A(n28666), .B(n45301), .X(n22214) );
  nand_x2_sg U42759 ( .A(n22193), .B(n22194), .X(n5926) );
  nand_x1_sg U42760 ( .A(n29028), .B(n45297), .X(n22236) );
  nand_x1_sg U42761 ( .A(n28505), .B(n45303), .X(n22235) );
  nand_x1_sg U42762 ( .A(n28405), .B(n45260), .X(n22268) );
  nand_x1_sg U42763 ( .A(n28848), .B(n45254), .X(n22267) );
  nand_x1_sg U42764 ( .A(n26989), .B(n45275), .X(n22279) );
  nand_x1_sg U42765 ( .A(n28660), .B(n45256), .X(n22262) );
  nand_x2_sg U42766 ( .A(n22241), .B(n22242), .X(n5810) );
  nand_x1_sg U42767 ( .A(n28499), .B(n45258), .X(n22282) );
  nand_x1_sg U42768 ( .A(n29021), .B(n45252), .X(n22283) );
  nand_x1_sg U42769 ( .A(n28842), .B(n45209), .X(n22315) );
  nand_x1_sg U42770 ( .A(n28399), .B(n45215), .X(n22316) );
  nand_x1_sg U42771 ( .A(n26983), .B(n45230), .X(n22327) );
  nand_x1_sg U42772 ( .A(n29170), .B(n45205), .X(n22310) );
  nand_x1_sg U42773 ( .A(n28654), .B(n45211), .X(n22309) );
  nand_x2_sg U42774 ( .A(n22288), .B(n22289), .X(n5880) );
  nand_x1_sg U42775 ( .A(n29015), .B(n45207), .X(n22331) );
  nand_x1_sg U42776 ( .A(n28493), .B(n45213), .X(n22330) );
  nand_x1_sg U42777 ( .A(n28836), .B(n45163), .X(n22362) );
  nand_x1_sg U42778 ( .A(n28393), .B(n45169), .X(n22363) );
  nand_x1_sg U42779 ( .A(n26977), .B(n45184), .X(n22374) );
  nand_x1_sg U42780 ( .A(n28648), .B(n45165), .X(n22357) );
  nand_x2_sg U42781 ( .A(n22336), .B(n22337), .X(n5839) );
  nand_x1_sg U42782 ( .A(n29008), .B(n45161), .X(n22378) );
  nand_x1_sg U42783 ( .A(n28487), .B(n45167), .X(n22377) );
  nand_x1_sg U42784 ( .A(n28830), .B(n45118), .X(n22410) );
  nand_x1_sg U42785 ( .A(n28387), .B(n45124), .X(n22411) );
  nand_x1_sg U42786 ( .A(n26971), .B(n45139), .X(n22422) );
  nand_x1_sg U42787 ( .A(n29158), .B(n45114), .X(n22405) );
  nand_x1_sg U42788 ( .A(n28642), .B(n45120), .X(n22404) );
  nand_x2_sg U42789 ( .A(n22383), .B(n22384), .X(n5803) );
  nand_x1_sg U42790 ( .A(n29002), .B(n45116), .X(n22426) );
  nand_x1_sg U42791 ( .A(n28481), .B(n45122), .X(n22425) );
  nand_x1_sg U42792 ( .A(n28824), .B(n45071), .X(n22456) );
  nand_x1_sg U42793 ( .A(n28381), .B(n45077), .X(n22457) );
  nand_x1_sg U42794 ( .A(n26965), .B(n45092), .X(n22468) );
  nand_x1_sg U42795 ( .A(n28636), .B(n45073), .X(n22451) );
  nand_x2_sg U42796 ( .A(n22431), .B(n22432), .X(n5824) );
  nand_x1_sg U42797 ( .A(n28995), .B(n45069), .X(n22472) );
  nand_x1_sg U42798 ( .A(n28475), .B(n45075), .X(n22471) );
  nand_x1_sg U42799 ( .A(n28818), .B(n45028), .X(n22502) );
  nand_x1_sg U42800 ( .A(n28375), .B(n45034), .X(n22503) );
  nand_x1_sg U42801 ( .A(n26959), .B(n45048), .X(n22514) );
  nand_x1_sg U42802 ( .A(n29146), .B(n45024), .X(n22497) );
  nand_x1_sg U42803 ( .A(n28630), .B(n45030), .X(n22496) );
  nand_x2_sg U42804 ( .A(n22477), .B(n22478), .X(n5903) );
  nand_x1_sg U42805 ( .A(n28989), .B(n45026), .X(n22518) );
  nand_x1_sg U42806 ( .A(n28469), .B(n45032), .X(n22517) );
  nand_x1_sg U42807 ( .A(n45017), .B(n26952), .X(n22552) );
  nand_x2_sg U42808 ( .A(n22523), .B(n22524), .X(n5947) );
  nand_x2_sg U42809 ( .A(n22559), .B(n22560), .X(n5933) );
  nand_x1_sg U42810 ( .A(n22730), .B(n22731), .X(n42312) );
  nand_x1_sg U42811 ( .A(n23007), .B(n23008), .X(n42311) );
  nand_x1_sg U42812 ( .A(n7826), .B(n47406), .X(n22978) );
  nand_x1_sg U42813 ( .A(n23287), .B(n23288), .X(n42310) );
  nand_x1_sg U42814 ( .A(n8644), .B(n47691), .X(n23255) );
  nand_x1_sg U42815 ( .A(n23566), .B(n23567), .X(n42309) );
  nand_x1_sg U42816 ( .A(n9464), .B(n47976), .X(n23535) );
  nand_x1_sg U42817 ( .A(n23845), .B(n23846), .X(n39675) );
  nand_x1_sg U42818 ( .A(n10283), .B(n48261), .X(n23814) );
  nand_x1_sg U42819 ( .A(n24124), .B(n24125), .X(n42308) );
  nand_x1_sg U42820 ( .A(n11102), .B(n48546), .X(n24093) );
  nand_x1_sg U42821 ( .A(n24403), .B(n24404), .X(n42307) );
  nand_x1_sg U42822 ( .A(n11921), .B(n48831), .X(n24372) );
  nand_x1_sg U42823 ( .A(n24681), .B(n24682), .X(n42306) );
  nand_x1_sg U42824 ( .A(n12740), .B(n49118), .X(n24651) );
  nand_x1_sg U42825 ( .A(n24960), .B(n24961), .X(n39671) );
  nand_x1_sg U42826 ( .A(n13559), .B(n49404), .X(n24929) );
  nand_x1_sg U42827 ( .A(n25239), .B(n25240), .X(n42305) );
  nand_x1_sg U42828 ( .A(n14378), .B(n49690), .X(n25208) );
  nand_x1_sg U42829 ( .A(n25518), .B(n25519), .X(n42304) );
  nand_x1_sg U42830 ( .A(n15197), .B(n49976), .X(n25487) );
  nand_x1_sg U42831 ( .A(n25795), .B(n25796), .X(n42303) );
  nand_x1_sg U42832 ( .A(n16016), .B(n50262), .X(n25766) );
  nand_x1_sg U42833 ( .A(n26355), .B(n26356), .X(n39667) );
  nand_x1_sg U42834 ( .A(n17654), .B(n50836), .X(n26322) );
  nand_x1_sg U42835 ( .A(n26633), .B(n26634), .X(n39665) );
  nand_x1_sg U42836 ( .A(n18475), .B(n51123), .X(n26603) );
  nand_x1_sg U42837 ( .A(n23124), .B(n42106), .X(n42105) );
  nand_x1_sg U42838 ( .A(n23124), .B(n42106), .X(n40157) );
  inv_x1_sg U42839 ( .A(n26787), .X(n51180) );
  inv_x1_sg U42840 ( .A(n26793), .X(n51159) );
  nand_x1_sg U42841 ( .A(n51159), .B(n51180), .X(n26786) );
  inv_x1_sg U42842 ( .A(n21748), .X(n51161) );
  inv_x1_sg U42843 ( .A(n21753), .X(n51141) );
  nand_x1_sg U42844 ( .A(n51141), .B(n51161), .X(n21747) );
  inv_x1_sg U42845 ( .A(n21795), .X(n51162) );
  inv_x1_sg U42846 ( .A(n21800), .X(n51142) );
  nand_x1_sg U42847 ( .A(n51142), .B(n51162), .X(n21794) );
  inv_x1_sg U42848 ( .A(n21842), .X(n51163) );
  inv_x1_sg U42849 ( .A(n21847), .X(n51143) );
  nand_x1_sg U42850 ( .A(n51143), .B(n51163), .X(n21841) );
  inv_x1_sg U42851 ( .A(n21888), .X(n51164) );
  inv_x1_sg U42852 ( .A(n21893), .X(n51144) );
  nand_x1_sg U42853 ( .A(n51144), .B(n51164), .X(n21887) );
  inv_x1_sg U42854 ( .A(n21935), .X(n51165) );
  inv_x1_sg U42855 ( .A(n21940), .X(n51145) );
  nand_x1_sg U42856 ( .A(n51145), .B(n51165), .X(n21934) );
  inv_x1_sg U42857 ( .A(n21981), .X(n51166) );
  inv_x1_sg U42858 ( .A(n21986), .X(n51146) );
  nand_x1_sg U42859 ( .A(n51146), .B(n51166), .X(n21980) );
  inv_x1_sg U42860 ( .A(n22028), .X(n51167) );
  inv_x1_sg U42861 ( .A(n22033), .X(n51147) );
  nand_x1_sg U42862 ( .A(n51147), .B(n51167), .X(n22027) );
  inv_x1_sg U42863 ( .A(n22074), .X(n51168) );
  inv_x1_sg U42864 ( .A(n22079), .X(n51148) );
  nand_x1_sg U42865 ( .A(n51148), .B(n51168), .X(n22073) );
  inv_x1_sg U42866 ( .A(n22122), .X(n51169) );
  inv_x1_sg U42867 ( .A(n22127), .X(n51149) );
  nand_x1_sg U42868 ( .A(n51149), .B(n51169), .X(n22121) );
  inv_x1_sg U42869 ( .A(n22169), .X(n51170) );
  inv_x1_sg U42870 ( .A(n22174), .X(n51150) );
  nand_x1_sg U42871 ( .A(n51150), .B(n51170), .X(n22168) );
  inv_x1_sg U42872 ( .A(n22217), .X(n51171) );
  inv_x1_sg U42873 ( .A(n22222), .X(n51151) );
  nand_x1_sg U42874 ( .A(n51151), .B(n51171), .X(n22216) );
  inv_x1_sg U42875 ( .A(n22264), .X(n51172) );
  inv_x1_sg U42876 ( .A(n22269), .X(n51152) );
  nand_x1_sg U42877 ( .A(n51152), .B(n51172), .X(n22263) );
  inv_x1_sg U42878 ( .A(n22312), .X(n51173) );
  inv_x1_sg U42879 ( .A(n22317), .X(n51153) );
  nand_x1_sg U42880 ( .A(n51153), .B(n51173), .X(n22311) );
  inv_x1_sg U42881 ( .A(n22359), .X(n51174) );
  inv_x1_sg U42882 ( .A(n22364), .X(n51154) );
  nand_x1_sg U42883 ( .A(n51154), .B(n51174), .X(n22358) );
  inv_x1_sg U42884 ( .A(n22407), .X(n51175) );
  inv_x1_sg U42885 ( .A(n22412), .X(n51155) );
  nand_x1_sg U42886 ( .A(n51155), .B(n51175), .X(n22406) );
  inv_x1_sg U42887 ( .A(n22453), .X(n51176) );
  inv_x1_sg U42888 ( .A(n22458), .X(n51156) );
  nand_x1_sg U42889 ( .A(n51156), .B(n51176), .X(n22452) );
  inv_x1_sg U42890 ( .A(n22499), .X(n51177) );
  inv_x1_sg U42891 ( .A(n22504), .X(n51157) );
  nand_x1_sg U42892 ( .A(n51157), .B(n51177), .X(n22498) );
  inv_x1_sg U42893 ( .A(n22539), .X(n51178) );
  inv_x1_sg U42894 ( .A(n22542), .X(n51158) );
  nand_x1_sg U42895 ( .A(n51158), .B(n51178), .X(n22538) );
  inv_x1_sg U42896 ( .A(n22580), .X(n51179) );
  inv_x1_sg U42897 ( .A(n22585), .X(n51160) );
  nand_x1_sg U42898 ( .A(n51160), .B(n51179), .X(n22579) );
  nand_x1_sg U42899 ( .A(n47385), .B(n22978), .X(n22976) );
  nand_x1_sg U42900 ( .A(n47670), .B(n23255), .X(n23253) );
  nand_x1_sg U42901 ( .A(n47955), .B(n23535), .X(n23533) );
  nand_x1_sg U42902 ( .A(n48240), .B(n23814), .X(n23812) );
  nand_x1_sg U42903 ( .A(n48525), .B(n24093), .X(n24091) );
  nand_x1_sg U42904 ( .A(n48810), .B(n24372), .X(n24370) );
  nand_x1_sg U42905 ( .A(n49097), .B(n24651), .X(n24649) );
  nand_x1_sg U42906 ( .A(n49383), .B(n24929), .X(n24927) );
  nand_x1_sg U42907 ( .A(n49669), .B(n25208), .X(n25206) );
  nand_x1_sg U42908 ( .A(n49955), .B(n25487), .X(n25485) );
  nand_x1_sg U42909 ( .A(n50241), .B(n25766), .X(n25764) );
  nor_x1_sg U42910 ( .A(n25976), .B(n25977), .X(n5743) );
  nand_x1_sg U42911 ( .A(n50815), .B(n26322), .X(n26329) );
  nand_x1_sg U42912 ( .A(n51102), .B(n26603), .X(n26601) );
  nand_x1_sg U42913 ( .A(n23090), .B(n23091), .X(n23084) );
  nand_x1_sg U42914 ( .A(n23370), .B(n23371), .X(n23364) );
  nand_x1_sg U42915 ( .A(n23649), .B(n23650), .X(n23643) );
  nand_x1_sg U42916 ( .A(n23928), .B(n23929), .X(n23922) );
  nand_x1_sg U42917 ( .A(n24207), .B(n24208), .X(n24201) );
  nand_x1_sg U42918 ( .A(n24486), .B(n24487), .X(n24480) );
  nand_x1_sg U42919 ( .A(n24764), .B(n24765), .X(n24758) );
  nand_x1_sg U42920 ( .A(n25043), .B(n25044), .X(n25037) );
  nand_x1_sg U42921 ( .A(n25322), .B(n25323), .X(n25316) );
  nand_x1_sg U42922 ( .A(n25601), .B(n25602), .X(n25595) );
  nand_x1_sg U42923 ( .A(n25878), .B(n25879), .X(n25872) );
  nand_x1_sg U42924 ( .A(n26438), .B(n26439), .X(n26432) );
  nand_x1_sg U42925 ( .A(n26716), .B(n26717), .X(n26710) );
  nand_x1_sg U42926 ( .A(n22813), .B(n22814), .X(n22807) );
  nand_x1_sg U42927 ( .A(n41740), .B(n28520), .X(n23264) );
  inv_x1_sg U42928 ( .A(n23264), .X(n42042) );
  nand_x1_sg U42929 ( .A(n20952), .B(n46550), .X(n38600) );
  inv_x1_sg U42930 ( .A(n22583), .X(n38601) );
  inv_x1_sg U42931 ( .A(n38601), .X(n38602) );
  inv_x1_sg U42932 ( .A(n6226), .X(n38603) );
  inv_x1_sg U42933 ( .A(n38603), .X(n38604) );
  inv_x1_sg U42934 ( .A(n6664), .X(n38605) );
  inv_x1_sg U42935 ( .A(n38605), .X(n38606) );
  inv_x1_sg U42936 ( .A(n6038), .X(n38607) );
  inv_x1_sg U42937 ( .A(n38607), .X(n38608) );
  inv_x1_sg U42938 ( .A(n6374), .X(n38609) );
  inv_x1_sg U42939 ( .A(n38609), .X(n38610) );
  inv_x1_sg U42940 ( .A(n6463), .X(n38611) );
  inv_x1_sg U42941 ( .A(n38611), .X(n38612) );
  inv_x1_sg U42942 ( .A(n6596), .X(n38613) );
  inv_x1_sg U42943 ( .A(n38613), .X(n38614) );
  inv_x1_sg U42944 ( .A(n6507), .X(n38615) );
  inv_x1_sg U42945 ( .A(n38615), .X(n38616) );
  inv_x1_sg U42946 ( .A(n41541), .X(n38617) );
  inv_x1_sg U42947 ( .A(n22575), .X(n38618) );
  inv_x1_sg U42948 ( .A(n38618), .X(n38619) );
  inv_x1_sg U42949 ( .A(n22594), .X(n38620) );
  inv_x1_sg U42950 ( .A(n38620), .X(n38621) );
  inv_x1_sg U42951 ( .A(n22565), .X(n38622) );
  inv_x1_sg U42952 ( .A(n38622), .X(n38623) );
  inv_x1_sg U42953 ( .A(n41542), .X(n38624) );
  inv_x1_sg U42954 ( .A(n6023), .X(n38625) );
  inv_x1_sg U42955 ( .A(n38625), .X(n38626) );
  inv_x1_sg U42956 ( .A(n22569), .X(n38627) );
  inv_x1_sg U42957 ( .A(n38627), .X(n38628) );
  inv_x1_sg U42958 ( .A(n41543), .X(n38629) );
  inv_x1_sg U42959 ( .A(n41544), .X(n38630) );
  inv_x1_sg U42960 ( .A(n6210), .X(n38631) );
  inv_x1_sg U42961 ( .A(n38631), .X(n38632) );
  inv_x1_sg U42962 ( .A(n5998), .X(n38633) );
  inv_x1_sg U42963 ( .A(n38633), .X(n38634) );
  inv_x1_sg U42964 ( .A(n42330), .X(n38635) );
  inv_x1_sg U42965 ( .A(n38635), .X(n38636) );
  inv_x1_sg U42966 ( .A(n6207), .X(n38637) );
  inv_x1_sg U42967 ( .A(n38637), .X(n38638) );
  inv_x1_sg U42968 ( .A(n42331), .X(n38639) );
  inv_x1_sg U42969 ( .A(n38639), .X(n38640) );
  inv_x1_sg U42970 ( .A(n6635), .X(n38641) );
  inv_x1_sg U42971 ( .A(n38641), .X(n38642) );
  inv_x1_sg U42972 ( .A(n6590), .X(n38643) );
  inv_x1_sg U42973 ( .A(n38643), .X(n38644) );
  inv_x1_sg U42974 ( .A(n6546), .X(n38645) );
  inv_x1_sg U42975 ( .A(n38645), .X(n38646) );
  inv_x1_sg U42976 ( .A(n6501), .X(n38647) );
  inv_x1_sg U42977 ( .A(n38647), .X(n38648) );
  inv_x1_sg U42978 ( .A(n6457), .X(n38649) );
  inv_x1_sg U42979 ( .A(n38649), .X(n38650) );
  inv_x1_sg U42980 ( .A(n6412), .X(n38651) );
  inv_x1_sg U42981 ( .A(n38651), .X(n38652) );
  inv_x1_sg U42982 ( .A(n6368), .X(n38653) );
  inv_x1_sg U42983 ( .A(n38653), .X(n38654) );
  inv_x1_sg U42984 ( .A(n6323), .X(n38655) );
  inv_x1_sg U42985 ( .A(n38655), .X(n38656) );
  inv_x1_sg U42986 ( .A(n6279), .X(n38657) );
  inv_x1_sg U42987 ( .A(n38657), .X(n38658) );
  inv_x1_sg U42988 ( .A(n6234), .X(n38659) );
  inv_x1_sg U42989 ( .A(n38659), .X(n38660) );
  inv_x1_sg U42990 ( .A(n6188), .X(n38661) );
  inv_x1_sg U42991 ( .A(n38661), .X(n38662) );
  inv_x1_sg U42992 ( .A(n6142), .X(n38663) );
  inv_x1_sg U42993 ( .A(n38663), .X(n38664) );
  inv_x1_sg U42994 ( .A(n6096), .X(n38665) );
  inv_x1_sg U42995 ( .A(n38665), .X(n38666) );
  inv_x1_sg U42996 ( .A(n41545), .X(n38667) );
  inv_x1_sg U42997 ( .A(n41546), .X(n38668) );
  inv_x1_sg U42998 ( .A(n41547), .X(n38669) );
  inv_x1_sg U42999 ( .A(n41548), .X(n38670) );
  inv_x1_sg U43000 ( .A(n41549), .X(n38671) );
  inv_x1_sg U43001 ( .A(n6655), .X(n38672) );
  inv_x1_sg U43002 ( .A(n38672), .X(n38673) );
  inv_x1_sg U43003 ( .A(n42333), .X(n38674) );
  inv_x1_sg U43004 ( .A(n38674), .X(n38675) );
  inv_x1_sg U43005 ( .A(n6567), .X(n38676) );
  inv_x1_sg U43006 ( .A(n38676), .X(n38677) );
  inv_x1_sg U43007 ( .A(n6522), .X(n38678) );
  inv_x1_sg U43008 ( .A(n38678), .X(n38679) );
  inv_x1_sg U43009 ( .A(n6478), .X(n38680) );
  inv_x1_sg U43010 ( .A(n38680), .X(n38681) );
  inv_x1_sg U43011 ( .A(n6433), .X(n38682) );
  inv_x1_sg U43012 ( .A(n38682), .X(n38683) );
  inv_x1_sg U43013 ( .A(n6389), .X(n38684) );
  inv_x1_sg U43014 ( .A(n38684), .X(n38685) );
  inv_x1_sg U43015 ( .A(n6344), .X(n38686) );
  inv_x1_sg U43016 ( .A(n38686), .X(n38687) );
  inv_x1_sg U43017 ( .A(n6611), .X(n38688) );
  inv_x1_sg U43018 ( .A(n38688), .X(n38689) );
  inv_x1_sg U43019 ( .A(n6300), .X(n38690) );
  inv_x1_sg U43020 ( .A(n38690), .X(n38691) );
  inv_x1_sg U43021 ( .A(n6055), .X(n38692) );
  inv_x1_sg U43022 ( .A(n38692), .X(n38693) );
  inv_x1_sg U43023 ( .A(n42334), .X(n38694) );
  inv_x1_sg U43024 ( .A(n38694), .X(n38695) );
  inv_x1_sg U43025 ( .A(n6255), .X(n38696) );
  inv_x1_sg U43026 ( .A(n38696), .X(n38697) );
  inv_x1_sg U43027 ( .A(n6118), .X(n38698) );
  inv_x1_sg U43028 ( .A(n38698), .X(n38699) );
  inv_x1_sg U43029 ( .A(n6687), .X(n38700) );
  inv_x1_sg U43030 ( .A(n38700), .X(n38701) );
  inv_x1_sg U43031 ( .A(n42335), .X(n38702) );
  inv_x1_sg U43032 ( .A(n38702), .X(n38703) );
  inv_x1_sg U43033 ( .A(n6552), .X(n38704) );
  inv_x1_sg U43034 ( .A(n38704), .X(n38705) );
  inv_x1_sg U43035 ( .A(n6418), .X(n38706) );
  inv_x1_sg U43036 ( .A(n38706), .X(n38707) );
  inv_x1_sg U43037 ( .A(n6285), .X(n38708) );
  inv_x1_sg U43038 ( .A(n38708), .X(n38709) );
  inv_x1_sg U43039 ( .A(n41550), .X(n38710) );
  inv_x1_sg U43040 ( .A(n41551), .X(n38711) );
  inv_x1_sg U43041 ( .A(n41552), .X(n38712) );
  inv_x1_sg U43042 ( .A(n42340), .X(n38713) );
  inv_x1_sg U43043 ( .A(n38713), .X(n38714) );
  inv_x1_sg U43044 ( .A(n42341), .X(n38715) );
  inv_x1_sg U43045 ( .A(n38715), .X(n38716) );
  inv_x1_sg U43046 ( .A(n42342), .X(n38717) );
  inv_x1_sg U43047 ( .A(n38717), .X(n38718) );
  inv_x1_sg U43048 ( .A(n42343), .X(n38719) );
  inv_x1_sg U43049 ( .A(n38719), .X(n38720) );
  inv_x1_sg U43050 ( .A(n6641), .X(n38721) );
  inv_x1_sg U43051 ( .A(n38721), .X(n38722) );
  inv_x1_sg U43052 ( .A(n6329), .X(n38723) );
  inv_x1_sg U43053 ( .A(n38723), .X(n38724) );
  inv_x1_sg U43054 ( .A(n41553), .X(n38725) );
  inv_x1_sg U43055 ( .A(n16929), .X(n38726) );
  inv_x1_sg U43056 ( .A(n38726), .X(n38727) );
  inv_x1_sg U43057 ( .A(n7104), .X(n38728) );
  inv_x1_sg U43058 ( .A(n38728), .X(n38729) );
  inv_x1_sg U43059 ( .A(n7922), .X(n38730) );
  inv_x1_sg U43060 ( .A(n38730), .X(n38731) );
  inv_x1_sg U43061 ( .A(n8740), .X(n38732) );
  inv_x1_sg U43062 ( .A(n38732), .X(n38733) );
  inv_x1_sg U43063 ( .A(n9560), .X(n38734) );
  inv_x1_sg U43064 ( .A(n38734), .X(n38735) );
  inv_x1_sg U43065 ( .A(n10379), .X(n38736) );
  inv_x1_sg U43066 ( .A(n38736), .X(n38737) );
  inv_x1_sg U43067 ( .A(n11198), .X(n38738) );
  inv_x1_sg U43068 ( .A(n38738), .X(n38739) );
  inv_x1_sg U43069 ( .A(n12017), .X(n38740) );
  inv_x1_sg U43070 ( .A(n38740), .X(n38741) );
  inv_x1_sg U43071 ( .A(n12836), .X(n38742) );
  inv_x1_sg U43072 ( .A(n38742), .X(n38743) );
  inv_x1_sg U43073 ( .A(n13655), .X(n38744) );
  inv_x1_sg U43074 ( .A(n38744), .X(n38745) );
  inv_x1_sg U43075 ( .A(n14474), .X(n38746) );
  inv_x1_sg U43076 ( .A(n38746), .X(n38747) );
  inv_x1_sg U43077 ( .A(n15293), .X(n38748) );
  inv_x1_sg U43078 ( .A(n38748), .X(n38749) );
  inv_x1_sg U43079 ( .A(n16112), .X(n38750) );
  inv_x1_sg U43080 ( .A(n38750), .X(n38751) );
  inv_x1_sg U43081 ( .A(n17750), .X(n38752) );
  inv_x1_sg U43082 ( .A(n38752), .X(n38753) );
  inv_x1_sg U43083 ( .A(n18571), .X(n38754) );
  inv_x1_sg U43084 ( .A(n38754), .X(n38755) );
  nand_x4_sg U43085 ( .A(n28979), .B(n28980), .X(n38756) );
  nand_x4_sg U43086 ( .A(n28979), .B(n28980), .X(n22595) );
  inv_x1_sg U43087 ( .A(\reg_yHat[0][2] ), .X(n38757) );
  inv_x1_sg U43088 ( .A(n38757), .X(n38758) );
  inv_x1_sg U43089 ( .A(\reg_yHat[0][3] ), .X(n38759) );
  inv_x1_sg U43090 ( .A(n38759), .X(n38760) );
  inv_x1_sg U43091 ( .A(\reg_yHat[1][2] ), .X(n38761) );
  inv_x1_sg U43092 ( .A(n38761), .X(n38762) );
  inv_x1_sg U43093 ( .A(\reg_yHat[1][3] ), .X(n38763) );
  inv_x1_sg U43094 ( .A(n38763), .X(n38764) );
  inv_x1_sg U43095 ( .A(\reg_yHat[2][2] ), .X(n38765) );
  inv_x1_sg U43096 ( .A(n38765), .X(n38766) );
  inv_x1_sg U43097 ( .A(\reg_yHat[2][3] ), .X(n38767) );
  inv_x1_sg U43098 ( .A(n38767), .X(n38768) );
  inv_x1_sg U43099 ( .A(\reg_yHat[3][2] ), .X(n38769) );
  inv_x1_sg U43100 ( .A(n38769), .X(n38770) );
  inv_x1_sg U43101 ( .A(\reg_yHat[3][3] ), .X(n38771) );
  inv_x1_sg U43102 ( .A(n38771), .X(n38772) );
  inv_x1_sg U43103 ( .A(\reg_yHat[4][2] ), .X(n38773) );
  inv_x1_sg U43104 ( .A(n38773), .X(n38774) );
  inv_x1_sg U43105 ( .A(\reg_yHat[4][3] ), .X(n38775) );
  inv_x1_sg U43106 ( .A(n38775), .X(n38776) );
  inv_x1_sg U43107 ( .A(\reg_yHat[5][2] ), .X(n38777) );
  inv_x1_sg U43108 ( .A(n38777), .X(n38778) );
  inv_x1_sg U43109 ( .A(\reg_yHat[5][3] ), .X(n38779) );
  inv_x1_sg U43110 ( .A(n38779), .X(n38780) );
  inv_x1_sg U43111 ( .A(\reg_yHat[6][2] ), .X(n38781) );
  inv_x1_sg U43112 ( .A(n38781), .X(n38782) );
  inv_x1_sg U43113 ( .A(\reg_yHat[6][3] ), .X(n38783) );
  inv_x1_sg U43114 ( .A(n38783), .X(n38784) );
  inv_x1_sg U43115 ( .A(\reg_yHat[7][2] ), .X(n38785) );
  inv_x1_sg U43116 ( .A(n38785), .X(n38786) );
  inv_x1_sg U43117 ( .A(\reg_yHat[7][3] ), .X(n38787) );
  inv_x1_sg U43118 ( .A(n38787), .X(n38788) );
  inv_x1_sg U43119 ( .A(\reg_yHat[8][2] ), .X(n38789) );
  inv_x1_sg U43120 ( .A(n38789), .X(n38790) );
  inv_x1_sg U43121 ( .A(\reg_yHat[8][3] ), .X(n38791) );
  inv_x1_sg U43122 ( .A(n38791), .X(n38792) );
  inv_x1_sg U43123 ( .A(\reg_yHat[9][2] ), .X(n38793) );
  inv_x1_sg U43124 ( .A(n38793), .X(n38794) );
  inv_x1_sg U43125 ( .A(\reg_yHat[9][3] ), .X(n38795) );
  inv_x1_sg U43126 ( .A(n38795), .X(n38796) );
  inv_x1_sg U43127 ( .A(\reg_yHat[10][2] ), .X(n38797) );
  inv_x1_sg U43128 ( .A(n38797), .X(n38798) );
  inv_x1_sg U43129 ( .A(\reg_yHat[10][3] ), .X(n38799) );
  inv_x1_sg U43130 ( .A(n38799), .X(n38800) );
  inv_x1_sg U43131 ( .A(\reg_yHat[11][2] ), .X(n38801) );
  inv_x1_sg U43132 ( .A(n38801), .X(n38802) );
  inv_x1_sg U43133 ( .A(\reg_yHat[11][3] ), .X(n38803) );
  inv_x1_sg U43134 ( .A(n38803), .X(n38804) );
  inv_x1_sg U43135 ( .A(\reg_yHat[13][2] ), .X(n38805) );
  inv_x1_sg U43136 ( .A(n38805), .X(n38806) );
  inv_x1_sg U43137 ( .A(\reg_yHat[13][3] ), .X(n38807) );
  inv_x1_sg U43138 ( .A(n38807), .X(n38808) );
  inv_x1_sg U43139 ( .A(\reg_yHat[14][2] ), .X(n38809) );
  inv_x1_sg U43140 ( .A(n38809), .X(n38810) );
  inv_x1_sg U43141 ( .A(\reg_yHat[14][3] ), .X(n38811) );
  inv_x1_sg U43142 ( .A(n38811), .X(n38812) );
  inv_x1_sg U43143 ( .A(n39273), .X(n38813) );
  inv_x1_sg U43144 ( .A(n39397), .X(n38814) );
  inv_x1_sg U43145 ( .A(n40018), .X(n38815) );
  inv_x1_sg U43146 ( .A(n38815), .X(n38816) );
  inv_x1_sg U43147 ( .A(n7641), .X(n38817) );
  inv_x1_sg U43148 ( .A(n8459), .X(n38818) );
  inv_x1_sg U43149 ( .A(n9279), .X(n38819) );
  inv_x1_sg U43150 ( .A(n10098), .X(n38820) );
  inv_x1_sg U43151 ( .A(n10917), .X(n38821) );
  inv_x1_sg U43152 ( .A(n11736), .X(n38822) );
  inv_x1_sg U43153 ( .A(n12555), .X(n38823) );
  inv_x1_sg U43154 ( .A(n13374), .X(n38824) );
  inv_x1_sg U43155 ( .A(n14193), .X(n38825) );
  inv_x1_sg U43156 ( .A(n15012), .X(n38826) );
  inv_x1_sg U43157 ( .A(n15831), .X(n38827) );
  inv_x1_sg U43158 ( .A(n18290), .X(n38828) );
  inv_x1_sg U43159 ( .A(n39116), .X(n38829) );
  inv_x1_sg U43160 ( .A(n39270), .X(n38830) );
  inv_x1_sg U43161 ( .A(n38830), .X(n38831) );
  inv_x1_sg U43162 ( .A(n40757), .X(n38832) );
  inv_x1_sg U43163 ( .A(n38832), .X(n38833) );
  inv_x1_sg U43164 ( .A(n38833), .X(n38834) );
  inv_x1_sg U43165 ( .A(n40764), .X(n38835) );
  inv_x1_sg U43166 ( .A(n38835), .X(n38836) );
  inv_x1_sg U43167 ( .A(n38836), .X(n38837) );
  inv_x1_sg U43168 ( .A(n40769), .X(n38838) );
  inv_x1_sg U43169 ( .A(n38838), .X(n38839) );
  inv_x1_sg U43170 ( .A(n38839), .X(n38840) );
  inv_x1_sg U43171 ( .A(n40776), .X(n38841) );
  inv_x1_sg U43172 ( .A(n38841), .X(n38842) );
  inv_x1_sg U43173 ( .A(n38842), .X(n38843) );
  inv_x1_sg U43174 ( .A(n40781), .X(n38844) );
  inv_x1_sg U43175 ( .A(n38844), .X(n38845) );
  inv_x1_sg U43176 ( .A(n38845), .X(n38846) );
  inv_x1_sg U43177 ( .A(n40788), .X(n38847) );
  inv_x1_sg U43178 ( .A(n40793), .X(n38848) );
  inv_x1_sg U43179 ( .A(n40800), .X(n38849) );
  inv_x1_sg U43180 ( .A(n38849), .X(n38850) );
  inv_x1_sg U43181 ( .A(n38850), .X(n38851) );
  inv_x1_sg U43182 ( .A(n40812), .X(n38852) );
  inv_x1_sg U43183 ( .A(n38852), .X(n38853) );
  inv_x1_sg U43184 ( .A(n38853), .X(n38854) );
  inv_x1_sg U43185 ( .A(n40817), .X(n38855) );
  inv_x1_sg U43186 ( .A(n40824), .X(n38856) );
  inv_x1_sg U43187 ( .A(n38856), .X(n38857) );
  inv_x1_sg U43188 ( .A(n38857), .X(n38858) );
  inv_x1_sg U43189 ( .A(n40829), .X(n38859) );
  inv_x1_sg U43190 ( .A(n40836), .X(n38860) );
  inv_x1_sg U43191 ( .A(n40841), .X(n38861) );
  inv_x1_sg U43192 ( .A(n18288), .X(n38862) );
  inv_x1_sg U43193 ( .A(n40845), .X(n38863) );
  inv_x1_sg U43194 ( .A(n15010), .X(n38864) );
  inv_x1_sg U43195 ( .A(n40850), .X(n38865) );
  inv_x1_sg U43196 ( .A(n14191), .X(n38866) );
  inv_x1_sg U43197 ( .A(n40855), .X(n38867) );
  inv_x1_sg U43198 ( .A(n13372), .X(n38868) );
  inv_x1_sg U43199 ( .A(n40860), .X(n38869) );
  inv_x1_sg U43200 ( .A(n12553), .X(n38870) );
  inv_x1_sg U43201 ( .A(n40865), .X(n38871) );
  inv_x1_sg U43202 ( .A(n11734), .X(n38872) );
  inv_x1_sg U43203 ( .A(n40870), .X(n38873) );
  inv_x1_sg U43204 ( .A(n10915), .X(n38874) );
  inv_x1_sg U43205 ( .A(n40875), .X(n38875) );
  inv_x1_sg U43206 ( .A(n10096), .X(n38876) );
  inv_x1_sg U43207 ( .A(n40880), .X(n38877) );
  inv_x1_sg U43208 ( .A(n9277), .X(n38878) );
  inv_x1_sg U43209 ( .A(n40885), .X(n38879) );
  inv_x1_sg U43210 ( .A(n8457), .X(n38880) );
  inv_x1_sg U43211 ( .A(n40890), .X(n38881) );
  inv_x1_sg U43212 ( .A(n15829), .X(n38882) );
  inv_x1_sg U43213 ( .A(n40895), .X(n38883) );
  inv_x1_sg U43214 ( .A(n16647), .X(n38884) );
  inv_x1_sg U43215 ( .A(n40900), .X(n38885) );
  inv_x1_sg U43216 ( .A(n17467), .X(n38886) );
  inv_x1_sg U43217 ( .A(n40905), .X(n38887) );
  inv_x1_sg U43218 ( .A(n6823), .X(n38888) );
  inv_x1_sg U43219 ( .A(n40910), .X(n38889) );
  inv_x1_sg U43220 ( .A(n7639), .X(n38890) );
  inv_x1_sg U43221 ( .A(n40915), .X(n38891) );
  inv_x1_sg U43222 ( .A(n40920), .X(n38892) );
  inv_x1_sg U43223 ( .A(n40924), .X(n38893) );
  inv_x1_sg U43224 ( .A(n40928), .X(n38894) );
  inv_x1_sg U43225 ( .A(n40932), .X(n38895) );
  inv_x1_sg U43226 ( .A(n40936), .X(n38896) );
  inv_x1_sg U43227 ( .A(n40940), .X(n38897) );
  inv_x1_sg U43228 ( .A(n40944), .X(n38898) );
  inv_x1_sg U43229 ( .A(n40948), .X(n38899) );
  inv_x1_sg U43230 ( .A(n40952), .X(n38900) );
  inv_x1_sg U43231 ( .A(n40956), .X(n38901) );
  inv_x1_sg U43232 ( .A(n40960), .X(n38902) );
  inv_x1_sg U43233 ( .A(n40964), .X(n38903) );
  inv_x1_sg U43234 ( .A(n40968), .X(n38904) );
  inv_x1_sg U43235 ( .A(n40972), .X(n38905) );
  inv_x1_sg U43236 ( .A(n5987), .X(n38906) );
  inv_x1_sg U43237 ( .A(n42385), .X(n38907) );
  inv_x1_sg U43238 ( .A(n40571), .X(n38908) );
  inv_x1_sg U43239 ( .A(n41918), .X(n38909) );
  inv_x1_sg U43240 ( .A(n40997), .X(n38910) );
  inv_x1_sg U43241 ( .A(n41042), .X(n38911) );
  inv_x1_sg U43242 ( .A(n39249), .X(n38912) );
  inv_x1_sg U43243 ( .A(n40316), .X(n38913) );
  inv_x1_sg U43244 ( .A(n41062), .X(n38914) );
  inv_x1_sg U43245 ( .A(n38914), .X(n38915) );
  inv_x1_sg U43246 ( .A(n5951), .X(n38916) );
  inv_x1_sg U43247 ( .A(n38919), .X(n38917) );
  inv_x1_sg U43248 ( .A(n41071), .X(n38918) );
  inv_x1_sg U43249 ( .A(n38918), .X(n38919) );
  inv_x1_sg U43250 ( .A(n38922), .X(n38920) );
  inv_x1_sg U43251 ( .A(n41076), .X(n38921) );
  inv_x1_sg U43252 ( .A(n38921), .X(n38922) );
  inv_x1_sg U43253 ( .A(n41081), .X(n38923) );
  inv_x1_sg U43254 ( .A(n38923), .X(n38924) );
  inv_x1_sg U43255 ( .A(n41085), .X(n38925) );
  inv_x1_sg U43256 ( .A(n38925), .X(n38926) );
  inv_x1_sg U43257 ( .A(n41089), .X(n38927) );
  inv_x1_sg U43258 ( .A(n38927), .X(n38928) );
  inv_x1_sg U43259 ( .A(n41093), .X(n38929) );
  inv_x1_sg U43260 ( .A(n38929), .X(n38930) );
  inv_x1_sg U43261 ( .A(n41097), .X(n38931) );
  inv_x1_sg U43262 ( .A(n38931), .X(n38932) );
  inv_x1_sg U43263 ( .A(n41101), .X(n38933) );
  inv_x1_sg U43264 ( .A(n38933), .X(n38934) );
  inv_x1_sg U43265 ( .A(n41105), .X(n38935) );
  inv_x1_sg U43266 ( .A(n38935), .X(n38936) );
  inv_x1_sg U43267 ( .A(n41109), .X(n38937) );
  inv_x1_sg U43268 ( .A(n38937), .X(n38938) );
  inv_x1_sg U43269 ( .A(n41113), .X(n38939) );
  inv_x1_sg U43270 ( .A(n38939), .X(n38940) );
  inv_x1_sg U43271 ( .A(n41294), .X(n38941) );
  inv_x1_sg U43272 ( .A(n41298), .X(n38942) );
  inv_x1_sg U43273 ( .A(n39275), .X(n38943) );
  inv_x1_sg U43274 ( .A(n38981), .X(n38944) );
  inv_x1_sg U43275 ( .A(n41574), .X(n38945) );
  inv_x1_sg U43276 ( .A(n41319), .X(n38946) );
  inv_x1_sg U43277 ( .A(n25082), .X(n38947) );
  inv_x1_sg U43278 ( .A(n38947), .X(n38948) );
  inv_x1_sg U43279 ( .A(n41324), .X(n38949) );
  inv_x1_sg U43280 ( .A(n24803), .X(n38950) );
  inv_x1_sg U43281 ( .A(n38950), .X(n38951) );
  inv_x1_sg U43282 ( .A(n41329), .X(n38952) );
  inv_x1_sg U43283 ( .A(n24525), .X(n38953) );
  inv_x1_sg U43284 ( .A(n38953), .X(n38954) );
  inv_x1_sg U43285 ( .A(n41334), .X(n38955) );
  inv_x1_sg U43286 ( .A(n42375), .X(n38956) );
  inv_x1_sg U43287 ( .A(n38956), .X(n38957) );
  inv_x1_sg U43288 ( .A(n41339), .X(n38958) );
  inv_x1_sg U43289 ( .A(n23409), .X(n38959) );
  inv_x1_sg U43290 ( .A(n38959), .X(n38960) );
  inv_x1_sg U43291 ( .A(n41344), .X(n38961) );
  inv_x1_sg U43292 ( .A(n42371), .X(n38962) );
  inv_x1_sg U43293 ( .A(n38962), .X(n38963) );
  inv_x1_sg U43294 ( .A(n41349), .X(n38964) );
  inv_x1_sg U43295 ( .A(n42373), .X(n38965) );
  inv_x1_sg U43296 ( .A(n38965), .X(n38966) );
  inv_x1_sg U43297 ( .A(n41354), .X(n38967) );
  inv_x1_sg U43298 ( .A(n42374), .X(n38968) );
  inv_x1_sg U43299 ( .A(n38968), .X(n38969) );
  inv_x1_sg U43300 ( .A(n41359), .X(n38970) );
  inv_x1_sg U43301 ( .A(n42386), .X(n38971) );
  inv_x1_sg U43302 ( .A(n38971), .X(n38972) );
  inv_x1_sg U43303 ( .A(n41364), .X(n38973) );
  inv_x1_sg U43304 ( .A(n42327), .X(n38974) );
  inv_x1_sg U43305 ( .A(n38974), .X(n38975) );
  inv_x1_sg U43306 ( .A(n41369), .X(n38976) );
  inv_x1_sg U43307 ( .A(n42376), .X(n38977) );
  inv_x1_sg U43308 ( .A(n38977), .X(n38978) );
  inv_x1_sg U43309 ( .A(n41374), .X(n38979) );
  inv_x1_sg U43310 ( .A(n41410), .X(n38980) );
  inv_x1_sg U43311 ( .A(n38980), .X(n38981) );
  inv_x1_sg U43312 ( .A(n5954), .X(n38982) );
  inv_x1_sg U43313 ( .A(n38982), .X(n38983) );
  inv_x1_sg U43314 ( .A(n41416), .X(n38984) );
  inv_x1_sg U43315 ( .A(n41471), .X(n38985) );
  inv_x1_sg U43316 ( .A(n42388), .X(n38986) );
  inv_x1_sg U43317 ( .A(n39769), .X(n38987) );
  inv_x1_sg U43318 ( .A(n42387), .X(n38988) );
  inv_x1_sg U43319 ( .A(n41489), .X(n38989) );
  inv_x1_sg U43320 ( .A(n38989), .X(n38990) );
  inv_x1_sg U43321 ( .A(n38839), .X(n38991) );
  inv_x1_sg U43322 ( .A(n41496), .X(n38992) );
  inv_x1_sg U43323 ( .A(n38992), .X(n38993) );
  inv_x1_sg U43324 ( .A(n39269), .X(n38994) );
  inv_x1_sg U43325 ( .A(n10749), .X(n38995) );
  inv_x1_sg U43326 ( .A(n9930), .X(n38996) );
  inv_x1_sg U43327 ( .A(n9110), .X(n38997) );
  inv_x1_sg U43328 ( .A(n8292), .X(n38998) );
  inv_x1_sg U43329 ( .A(n14025), .X(n38999) );
  inv_x1_sg U43330 ( .A(n13206), .X(n39000) );
  inv_x1_sg U43331 ( .A(n12387), .X(n39001) );
  inv_x1_sg U43332 ( .A(n11568), .X(n39002) );
  inv_x1_sg U43333 ( .A(n18941), .X(n39003) );
  inv_x1_sg U43334 ( .A(n16482), .X(n39004) );
  inv_x1_sg U43335 ( .A(n15663), .X(n39005) );
  inv_x1_sg U43336 ( .A(n14844), .X(n39006) );
  inv_x1_sg U43337 ( .A(n18120), .X(n39007) );
  inv_x1_sg U43338 ( .A(n18635), .X(n39008) );
  nand_x1_sg U43339 ( .A(n41807), .B(n40671), .X(n18635) );
  inv_x1_sg U43340 ( .A(n16176), .X(n39009) );
  nand_x1_sg U43341 ( .A(n41803), .B(n40676), .X(n16176) );
  inv_x1_sg U43342 ( .A(n14538), .X(n39010) );
  nand_x1_sg U43343 ( .A(n41799), .B(n40621), .X(n14538) );
  inv_x1_sg U43344 ( .A(n13719), .X(n39011) );
  nand_x1_sg U43345 ( .A(n41797), .B(n40651), .X(n13719) );
  inv_x1_sg U43346 ( .A(n12900), .X(n39012) );
  nand_x1_sg U43347 ( .A(n41795), .B(n40661), .X(n12900) );
  inv_x1_sg U43348 ( .A(n12081), .X(n39013) );
  nand_x1_sg U43349 ( .A(n41793), .B(n40636), .X(n12081) );
  inv_x1_sg U43350 ( .A(n11262), .X(n39014) );
  nand_x1_sg U43351 ( .A(n41791), .B(n40641), .X(n11262) );
  inv_x1_sg U43352 ( .A(n10443), .X(n39015) );
  nand_x1_sg U43353 ( .A(n41789), .B(n40656), .X(n10443) );
  inv_x1_sg U43354 ( .A(n9624), .X(n39016) );
  nand_x1_sg U43355 ( .A(n41787), .B(n40666), .X(n9624) );
  inv_x1_sg U43356 ( .A(n8804), .X(n39017) );
  nand_x1_sg U43357 ( .A(n41785), .B(n40626), .X(n8804) );
  inv_x1_sg U43358 ( .A(n16992), .X(n39018) );
  nand_x1_sg U43359 ( .A(n40074), .B(n40581), .X(n16992) );
  inv_x1_sg U43360 ( .A(n7167), .X(n39019) );
  nand_x1_sg U43361 ( .A(n41781), .B(n40576), .X(n7167) );
  inv_x1_sg U43362 ( .A(n17814), .X(n39020) );
  nand_x1_sg U43363 ( .A(n41805), .B(n40649), .X(n17814) );
  inv_x1_sg U43364 ( .A(n15357), .X(n39021) );
  nand_x1_sg U43365 ( .A(n41801), .B(n40681), .X(n15357) );
  inv_x1_sg U43366 ( .A(n7986), .X(n39022) );
  nand_x1_sg U43367 ( .A(n41783), .B(n40631), .X(n7986) );
  inv_x1_sg U43368 ( .A(n39313), .X(n39023) );
  inv_x1_sg U43369 ( .A(n16821), .X(n39024) );
  inv_x1_sg U43370 ( .A(n17642), .X(n39025) );
  inv_x1_sg U43371 ( .A(n18463), .X(n39026) );
  inv_x1_sg U43372 ( .A(n15185), .X(n39027) );
  inv_x1_sg U43373 ( .A(n16004), .X(n39028) );
  inv_x1_sg U43374 ( .A(n14366), .X(n39029) );
  inv_x1_sg U43375 ( .A(n13547), .X(n39030) );
  inv_x1_sg U43376 ( .A(n11909), .X(n39031) );
  inv_x1_sg U43377 ( .A(n10271), .X(n39032) );
  inv_x1_sg U43378 ( .A(n11090), .X(n39033) );
  inv_x1_sg U43379 ( .A(n9452), .X(n39034) );
  inv_x1_sg U43380 ( .A(n7814), .X(n39035) );
  inv_x1_sg U43381 ( .A(n8632), .X(n39036) );
  inv_x1_sg U43382 ( .A(n6997), .X(n39037) );
  inv_x1_sg U43383 ( .A(n7445), .X(n39038) );
  inv_x1_sg U43384 ( .A(n9081), .X(n39039) );
  inv_x1_sg U43385 ( .A(n42319), .X(n39040) );
  inv_x1_sg U43386 ( .A(n10720), .X(n39041) );
  inv_x1_sg U43387 ( .A(n42318), .X(n39042) );
  inv_x1_sg U43388 ( .A(n12358), .X(n39043) );
  inv_x1_sg U43389 ( .A(n42317), .X(n39044) );
  inv_x1_sg U43390 ( .A(n13996), .X(n39045) );
  inv_x1_sg U43391 ( .A(n42316), .X(n39046) );
  inv_x1_sg U43392 ( .A(n15634), .X(n39047) );
  inv_x1_sg U43393 ( .A(n42315), .X(n39048) );
  inv_x1_sg U43394 ( .A(n18091), .X(n39049) );
  inv_x1_sg U43395 ( .A(n42314), .X(n39050) );
  inv_x1_sg U43396 ( .A(n42313), .X(n39051) );
  inv_x1_sg U43397 ( .A(n42235), .X(n39052) );
  inv_x1_sg U43398 ( .A(n40216), .X(n39053) );
  inv_x1_sg U43399 ( .A(n40184), .X(n39054) );
  inv_x1_sg U43400 ( .A(n40168), .X(n39055) );
  inv_x1_sg U43401 ( .A(n40172), .X(n39056) );
  inv_x1_sg U43402 ( .A(n40188), .X(n39057) );
  inv_x1_sg U43403 ( .A(n40176), .X(n39058) );
  inv_x1_sg U43404 ( .A(n40192), .X(n39059) );
  inv_x1_sg U43405 ( .A(n40196), .X(n39060) );
  inv_x1_sg U43406 ( .A(n40200), .X(n39061) );
  inv_x1_sg U43407 ( .A(n40204), .X(n39062) );
  inv_x1_sg U43408 ( .A(n40208), .X(n39063) );
  inv_x1_sg U43409 ( .A(n40212), .X(n39064) );
  inv_x1_sg U43410 ( .A(n40180), .X(n39065) );
  inv_x1_sg U43411 ( .A(n42097), .X(n39066) );
  inv_x1_sg U43412 ( .A(n42094), .X(n39067) );
  inv_x1_sg U43413 ( .A(n42093), .X(n39068) );
  inv_x1_sg U43414 ( .A(n40360), .X(n39069) );
  inv_x1_sg U43415 ( .A(n42095), .X(n39070) );
  inv_x1_sg U43416 ( .A(n42098), .X(n39071) );
  inv_x1_sg U43417 ( .A(n42101), .X(n39072) );
  inv_x1_sg U43418 ( .A(n42103), .X(n39073) );
  inv_x1_sg U43419 ( .A(n42102), .X(n39074) );
  inv_x1_sg U43420 ( .A(n42100), .X(n39075) );
  inv_x1_sg U43421 ( .A(n42099), .X(n39076) );
  inv_x1_sg U43422 ( .A(n40581), .X(n39077) );
  inv_x1_sg U43423 ( .A(n40576), .X(n39078) );
  inv_x1_sg U43424 ( .A(n12728), .X(n39079) );
  inv_x1_sg U43425 ( .A(n51137), .X(n39080) );
  inv_x1_sg U43426 ( .A(n39080), .X(n39081) );
  inv_x1_sg U43427 ( .A(n51136), .X(n39082) );
  inv_x1_sg U43428 ( .A(n39082), .X(n39083) );
  inv_x1_sg U43429 ( .A(n42383), .X(n39084) );
  inv_x1_sg U43430 ( .A(\L2_0/n3047 ), .X(n39085) );
  inv_x1_sg U43431 ( .A(n39085), .X(n39086) );
  inv_x1_sg U43432 ( .A(n41201), .X(n39087) );
  inv_x1_sg U43433 ( .A(n5779), .X(n39088) );
  inv_x1_sg U43434 ( .A(n39088), .X(n39089) );
  inv_x1_sg U43435 ( .A(n41206), .X(n39090) );
  inv_x1_sg U43436 ( .A(n42378), .X(n39091) );
  inv_x1_sg U43437 ( .A(n39091), .X(n39092) );
  inv_x1_sg U43438 ( .A(n41210), .X(n39093) );
  inv_x1_sg U43439 ( .A(n42338), .X(n39094) );
  inv_x1_sg U43440 ( .A(n39094), .X(n39095) );
  inv_x1_sg U43441 ( .A(n41215), .X(n39096) );
  inv_x1_sg U43442 ( .A(\L2_0/n3127 ), .X(n39097) );
  inv_x1_sg U43443 ( .A(n39097), .X(n39098) );
  inv_x1_sg U43444 ( .A(n41220), .X(n39099) );
  inv_x1_sg U43445 ( .A(n42381), .X(n39100) );
  inv_x1_sg U43446 ( .A(n39100), .X(n39101) );
  inv_x1_sg U43447 ( .A(n41225), .X(n39102) );
  inv_x1_sg U43448 ( .A(\L2_0/n2727 ), .X(n39103) );
  inv_x1_sg U43449 ( .A(n39103), .X(n39104) );
  inv_x1_sg U43450 ( .A(n41230), .X(n39105) );
  inv_x1_sg U43451 ( .A(\L2_0/n3367 ), .X(n39106) );
  inv_x1_sg U43452 ( .A(n39106), .X(n39107) );
  inv_x1_sg U43453 ( .A(n41235), .X(n39108) );
  inv_x1_sg U43454 ( .A(n42382), .X(n39109) );
  inv_x1_sg U43455 ( .A(n39109), .X(n39110) );
  inv_x1_sg U43456 ( .A(n41240), .X(n39111) );
  inv_x1_sg U43457 ( .A(n42384), .X(n39112) );
  inv_x1_sg U43458 ( .A(n39112), .X(n39113) );
  inv_x1_sg U43459 ( .A(n41245), .X(n39114) );
  inv_x1_sg U43460 ( .A(n42018), .X(n39115) );
  inv_x1_sg U43461 ( .A(n41250), .X(n39116) );
  inv_x1_sg U43462 ( .A(\L2_0/n2967 ), .X(n39117) );
  inv_x1_sg U43463 ( .A(n39117), .X(n39118) );
  inv_x1_sg U43464 ( .A(n41255), .X(n39119) );
  inv_x1_sg U43465 ( .A(n42379), .X(n39120) );
  inv_x1_sg U43466 ( .A(n39120), .X(n39121) );
  inv_x1_sg U43467 ( .A(n41260), .X(n39122) );
  inv_x1_sg U43468 ( .A(n41275), .X(n39123) );
  inv_x1_sg U43469 ( .A(n41275), .X(n39124) );
  inv_x1_sg U43470 ( .A(n42329), .X(n39125) );
  inv_x1_sg U43471 ( .A(n39125), .X(n39126) );
  inv_x1_sg U43472 ( .A(n41279), .X(n39127) );
  inv_x1_sg U43473 ( .A(\L2_0/n3447 ), .X(n39128) );
  inv_x1_sg U43474 ( .A(n39128), .X(n39129) );
  inv_x1_sg U43475 ( .A(n41284), .X(n39130) );
  inv_x1_sg U43476 ( .A(n42380), .X(n39131) );
  inv_x1_sg U43477 ( .A(n39131), .X(n39132) );
  inv_x1_sg U43478 ( .A(n41289), .X(n39133) );
  inv_x1_sg U43479 ( .A(n40036), .X(n39134) );
  inv_x1_sg U43480 ( .A(n9274), .X(n39135) );
  inv_x1_sg U43481 ( .A(n39348), .X(n39136) );
  inv_x1_sg U43482 ( .A(n41303), .X(n39137) );
  inv_x1_sg U43483 ( .A(n40035), .X(n39138) );
  inv_x1_sg U43484 ( .A(n41379), .X(n39139) );
  inv_x1_sg U43485 ( .A(n41379), .X(n39140) );
  inv_x1_sg U43486 ( .A(n40031), .X(n39141) );
  inv_x1_sg U43487 ( .A(n41384), .X(n39142) );
  inv_x1_sg U43488 ( .A(n41384), .X(n39143) );
  inv_x1_sg U43489 ( .A(n40027), .X(n39144) );
  inv_x1_sg U43490 ( .A(n41389), .X(n39145) );
  inv_x1_sg U43491 ( .A(n41389), .X(n39146) );
  inv_x1_sg U43492 ( .A(n5994), .X(n39147) );
  inv_x1_sg U43493 ( .A(n39147), .X(n39148) );
  inv_x1_sg U43494 ( .A(n41394), .X(n39149) );
  inv_x1_sg U43495 ( .A(n40021), .X(n39150) );
  inv_x1_sg U43496 ( .A(n41401), .X(n39151) );
  inv_x1_sg U43497 ( .A(n41401), .X(n39152) );
  inv_x1_sg U43498 ( .A(n40016), .X(n39153) );
  inv_x1_sg U43499 ( .A(n41406), .X(n39154) );
  inv_x1_sg U43500 ( .A(n41406), .X(n39155) );
  inv_x1_sg U43501 ( .A(n38985), .X(n39156) );
  inv_x1_sg U43502 ( .A(n39156), .X(n39157) );
  inv_x1_sg U43503 ( .A(n41411), .X(n39158) );
  inv_x1_sg U43504 ( .A(n41423), .X(n39159) );
  inv_x1_sg U43505 ( .A(n39159), .X(n39160) );
  inv_x1_sg U43506 ( .A(n39159), .X(n39161) );
  inv_x1_sg U43507 ( .A(n39161), .X(n39162) );
  inv_x1_sg U43508 ( .A(n39161), .X(n39163) );
  inv_x1_sg U43509 ( .A(n41455), .X(n39164) );
  inv_x1_sg U43510 ( .A(n39164), .X(n39165) );
  inv_x1_sg U43511 ( .A(n39164), .X(n39166) );
  inv_x1_sg U43512 ( .A(n39166), .X(n39167) );
  inv_x1_sg U43513 ( .A(n39166), .X(n39168) );
  inv_x1_sg U43514 ( .A(n41432), .X(n39169) );
  inv_x1_sg U43515 ( .A(n39169), .X(n39170) );
  inv_x1_sg U43516 ( .A(n39169), .X(n39171) );
  inv_x1_sg U43517 ( .A(n39171), .X(n39172) );
  inv_x1_sg U43518 ( .A(n39171), .X(n39173) );
  inv_x1_sg U43519 ( .A(n41437), .X(n39174) );
  inv_x1_sg U43520 ( .A(n39174), .X(n39175) );
  inv_x1_sg U43521 ( .A(n39174), .X(n39176) );
  inv_x1_sg U43522 ( .A(n39176), .X(n39177) );
  inv_x1_sg U43523 ( .A(n39176), .X(n39178) );
  inv_x1_sg U43524 ( .A(n41446), .X(n39179) );
  inv_x1_sg U43525 ( .A(n39179), .X(n39180) );
  inv_x1_sg U43526 ( .A(n39179), .X(n39181) );
  inv_x1_sg U43527 ( .A(n39181), .X(n39182) );
  inv_x1_sg U43528 ( .A(n39181), .X(n39183) );
  inv_x1_sg U43529 ( .A(n41446), .X(n39184) );
  inv_x1_sg U43530 ( .A(n39184), .X(n39185) );
  inv_x1_sg U43531 ( .A(n39184), .X(n39186) );
  inv_x1_sg U43532 ( .A(n39186), .X(n39187) );
  inv_x1_sg U43533 ( .A(n39186), .X(n39188) );
  inv_x1_sg U43534 ( .A(n41455), .X(n39189) );
  inv_x1_sg U43535 ( .A(n39189), .X(n39190) );
  inv_x1_sg U43536 ( .A(n39189), .X(n39191) );
  inv_x1_sg U43537 ( .A(n39191), .X(n39192) );
  inv_x1_sg U43538 ( .A(n39190), .X(n39193) );
  inv_x1_sg U43539 ( .A(n41455), .X(n39194) );
  inv_x1_sg U43540 ( .A(n39194), .X(n39195) );
  inv_x1_sg U43541 ( .A(n39194), .X(n39196) );
  inv_x1_sg U43542 ( .A(n39195), .X(n39197) );
  inv_x1_sg U43543 ( .A(n39196), .X(n39198) );
  inv_x1_sg U43544 ( .A(n42377), .X(n39199) );
  inv_x1_sg U43545 ( .A(n41949), .X(n39200) );
  inv_x1_sg U43546 ( .A(n38814), .X(n39201) );
  inv_x1_sg U43547 ( .A(n39399), .X(n39202) );
  inv_x1_sg U43548 ( .A(n39409), .X(n39203) );
  inv_x1_sg U43549 ( .A(n6971), .X(n39204) );
  inv_x1_sg U43550 ( .A(n39723), .X(n39205) );
  inv_x1_sg U43551 ( .A(n39720), .X(n39206) );
  inv_x1_sg U43552 ( .A(n39717), .X(n39207) );
  inv_x1_sg U43553 ( .A(n39714), .X(n39208) );
  inv_x1_sg U43554 ( .A(n39711), .X(n39209) );
  inv_x1_sg U43555 ( .A(n39708), .X(n39210) );
  inv_x1_sg U43556 ( .A(n39705), .X(n39211) );
  inv_x1_sg U43557 ( .A(n39702), .X(n39212) );
  inv_x1_sg U43558 ( .A(n39699), .X(n39213) );
  inv_x1_sg U43559 ( .A(n39696), .X(n39214) );
  inv_x1_sg U43560 ( .A(n39693), .X(n39215) );
  inv_x1_sg U43561 ( .A(n39690), .X(n39216) );
  inv_x1_sg U43562 ( .A(n39687), .X(n39217) );
  inv_x1_sg U43563 ( .A(n39684), .X(n39218) );
  inv_x1_sg U43564 ( .A(n39084), .X(n39219) );
  inv_x1_sg U43565 ( .A(n41196), .X(n39220) );
  inv_x1_sg U43566 ( .A(n41862), .X(n39221) );
  inv_x1_sg U43567 ( .A(n41191), .X(n39222) );
  inv_x1_sg U43568 ( .A(n41863), .X(n39223) );
  inv_x1_sg U43569 ( .A(n41186), .X(n39224) );
  inv_x1_sg U43570 ( .A(n41864), .X(n39225) );
  inv_x1_sg U43571 ( .A(n41181), .X(n39226) );
  inv_x1_sg U43572 ( .A(n41865), .X(n39227) );
  inv_x1_sg U43573 ( .A(n41176), .X(n39228) );
  inv_x1_sg U43574 ( .A(n41866), .X(n39229) );
  inv_x1_sg U43575 ( .A(n41171), .X(n39230) );
  inv_x1_sg U43576 ( .A(n41867), .X(n39231) );
  inv_x1_sg U43577 ( .A(n41166), .X(n39232) );
  inv_x1_sg U43578 ( .A(n41868), .X(n39233) );
  inv_x1_sg U43579 ( .A(n41161), .X(n39234) );
  inv_x1_sg U43580 ( .A(n41869), .X(n39235) );
  inv_x1_sg U43581 ( .A(n41156), .X(n39236) );
  inv_x1_sg U43582 ( .A(n41870), .X(n39237) );
  inv_x1_sg U43583 ( .A(n41151), .X(n39238) );
  inv_x1_sg U43584 ( .A(n41871), .X(n39239) );
  inv_x1_sg U43585 ( .A(n41146), .X(n39240) );
  inv_x1_sg U43586 ( .A(n41872), .X(n39241) );
  inv_x1_sg U43587 ( .A(n41141), .X(n39242) );
  inv_x1_sg U43588 ( .A(n41873), .X(n39243) );
  inv_x1_sg U43589 ( .A(n41136), .X(n39244) );
  inv_x1_sg U43590 ( .A(n41874), .X(n39245) );
  inv_x1_sg U43591 ( .A(n41131), .X(n39246) );
  inv_x1_sg U43592 ( .A(n41930), .X(n39247) );
  inv_x1_sg U43593 ( .A(n39247), .X(n39248) );
  inv_x1_sg U43594 ( .A(n41126), .X(n39249) );
  inv_x1_sg U43595 ( .A(n41946), .X(n39250) );
  inv_x1_sg U43596 ( .A(n39250), .X(n39251) );
  inv_x1_sg U43597 ( .A(n41121), .X(n39252) );
  inv_x1_sg U43598 ( .A(n41116), .X(n39253) );
  inv_x1_sg U43599 ( .A(n41112), .X(n39254) );
  inv_x1_sg U43600 ( .A(n41108), .X(n39255) );
  inv_x1_sg U43601 ( .A(n41104), .X(n39256) );
  inv_x1_sg U43602 ( .A(n41100), .X(n39257) );
  inv_x1_sg U43603 ( .A(n41096), .X(n39258) );
  inv_x1_sg U43604 ( .A(n41092), .X(n39259) );
  inv_x1_sg U43605 ( .A(n41088), .X(n39260) );
  inv_x1_sg U43606 ( .A(n41084), .X(n39261) );
  inv_x1_sg U43607 ( .A(n41080), .X(n39262) );
  inv_x1_sg U43608 ( .A(n38920), .X(n39263) );
  inv_x1_sg U43609 ( .A(n38917), .X(n39264) );
  inv_x1_sg U43610 ( .A(n41065), .X(n39265) );
  inv_x1_sg U43611 ( .A(n41061), .X(n39266) );
  inv_x1_sg U43612 ( .A(n41272), .X(n39267) );
  inv_x1_sg U43613 ( .A(n39286), .X(n39268) );
  inv_x1_sg U43614 ( .A(n40810), .X(n39269) );
  inv_x1_sg U43615 ( .A(n39269), .X(n39270) );
  inv_x1_sg U43616 ( .A(n39408), .X(n39271) );
  inv_x1_sg U43617 ( .A(n41506), .X(n39272) );
  inv_x1_sg U43618 ( .A(n41310), .X(n39273) );
  inv_x1_sg U43619 ( .A(n39273), .X(n39274) );
  inv_x1_sg U43620 ( .A(n39273), .X(n39275) );
  inv_x1_sg U43621 ( .A(n39274), .X(n39276) );
  inv_x1_sg U43622 ( .A(n38813), .X(n39277) );
  inv_x1_sg U43623 ( .A(n39656), .X(n39278) );
  inv_x1_sg U43624 ( .A(n41460), .X(n39279) );
  inv_x1_sg U43625 ( .A(n41460), .X(n39280) );
  inv_x1_sg U43626 ( .A(n39199), .X(n39281) );
  inv_x1_sg U43627 ( .A(n39652), .X(n39282) );
  inv_x1_sg U43628 ( .A(n41465), .X(n39283) );
  inv_x1_sg U43629 ( .A(n39200), .X(n39284) );
  inv_x1_sg U43630 ( .A(n39287), .X(n39285) );
  inv_x1_sg U43631 ( .A(n39430), .X(n39286) );
  inv_x1_sg U43632 ( .A(n39423), .X(n39287) );
  inv_x1_sg U43633 ( .A(n41632), .X(n39288) );
  inv_x1_sg U43634 ( .A(n6996), .X(n39289) );
  inv_x1_sg U43635 ( .A(n39289), .X(n39290) );
  inv_x1_sg U43636 ( .A(n17641), .X(n39291) );
  inv_x1_sg U43637 ( .A(n39291), .X(n39292) );
  inv_x1_sg U43638 ( .A(n18462), .X(n39293) );
  inv_x1_sg U43639 ( .A(n39293), .X(n39294) );
  inv_x1_sg U43640 ( .A(n16003), .X(n39295) );
  inv_x1_sg U43641 ( .A(n39295), .X(n39296) );
  inv_x1_sg U43642 ( .A(n15184), .X(n39297) );
  inv_x1_sg U43643 ( .A(n39297), .X(n39298) );
  inv_x1_sg U43644 ( .A(n14365), .X(n39299) );
  inv_x1_sg U43645 ( .A(n39299), .X(n39300) );
  inv_x1_sg U43646 ( .A(n13546), .X(n39301) );
  inv_x1_sg U43647 ( .A(n39301), .X(n39302) );
  inv_x1_sg U43648 ( .A(n12727), .X(n39303) );
  inv_x1_sg U43649 ( .A(n39303), .X(n39304) );
  inv_x1_sg U43650 ( .A(n11908), .X(n39305) );
  inv_x1_sg U43651 ( .A(n39305), .X(n39306) );
  inv_x1_sg U43652 ( .A(n11089), .X(n39307) );
  inv_x1_sg U43653 ( .A(n39307), .X(n39308) );
  inv_x1_sg U43654 ( .A(n10270), .X(n39309) );
  inv_x1_sg U43655 ( .A(n39309), .X(n39310) );
  inv_x1_sg U43656 ( .A(n9451), .X(n39311) );
  inv_x1_sg U43657 ( .A(n39311), .X(n39312) );
  nand_x1_sg U43658 ( .A(n40250), .B(n40361), .X(n39313) );
  inv_x1_sg U43659 ( .A(n7813), .X(n39314) );
  inv_x1_sg U43660 ( .A(n39314), .X(n39315) );
  inv_x1_sg U43661 ( .A(n16820), .X(n39316) );
  inv_x1_sg U43662 ( .A(n39316), .X(n39317) );
  inv_x1_sg U43663 ( .A(n16966), .X(n39318) );
  inv_x1_sg U43664 ( .A(n39318), .X(n39319) );
  inv_x1_sg U43665 ( .A(n18608), .X(n39320) );
  inv_x1_sg U43666 ( .A(n39320), .X(n39321) );
  inv_x1_sg U43667 ( .A(n17787), .X(n39322) );
  inv_x1_sg U43668 ( .A(n39322), .X(n39323) );
  inv_x1_sg U43669 ( .A(n16149), .X(n39324) );
  inv_x1_sg U43670 ( .A(n39324), .X(n39325) );
  inv_x1_sg U43671 ( .A(n15330), .X(n39326) );
  inv_x1_sg U43672 ( .A(n39326), .X(n39327) );
  inv_x1_sg U43673 ( .A(n14511), .X(n39328) );
  inv_x1_sg U43674 ( .A(n39328), .X(n39329) );
  inv_x1_sg U43675 ( .A(n13692), .X(n39330) );
  inv_x1_sg U43676 ( .A(n39330), .X(n39331) );
  inv_x1_sg U43677 ( .A(n12873), .X(n39332) );
  inv_x1_sg U43678 ( .A(n39332), .X(n39333) );
  inv_x1_sg U43679 ( .A(n12054), .X(n39334) );
  inv_x1_sg U43680 ( .A(n39334), .X(n39335) );
  inv_x1_sg U43681 ( .A(n11235), .X(n39336) );
  inv_x1_sg U43682 ( .A(n39336), .X(n39337) );
  inv_x1_sg U43683 ( .A(n10416), .X(n39338) );
  inv_x1_sg U43684 ( .A(n39338), .X(n39339) );
  inv_x1_sg U43685 ( .A(n9597), .X(n39340) );
  inv_x1_sg U43686 ( .A(n39340), .X(n39341) );
  inv_x1_sg U43687 ( .A(n8777), .X(n39342) );
  inv_x1_sg U43688 ( .A(n39342), .X(n39343) );
  inv_x1_sg U43689 ( .A(n7959), .X(n39344) );
  inv_x1_sg U43690 ( .A(n39344), .X(n39345) );
  inv_x1_sg U43691 ( .A(n7141), .X(n39346) );
  inv_x1_sg U43692 ( .A(n39346), .X(n39347) );
  inv_x1_sg U43693 ( .A(n22638), .X(n39348) );
  inv_x1_sg U43694 ( .A(n39348), .X(n39349) );
  nand_x1_sg U43695 ( .A(n22737), .B(n22738), .X(n39350) );
  nand_x1_sg U43696 ( .A(n23294), .B(n23295), .X(n39351) );
  nand_x1_sg U43697 ( .A(n23014), .B(n23015), .X(n39352) );
  nand_x1_sg U43698 ( .A(n23573), .B(n23574), .X(n39353) );
  nand_x1_sg U43699 ( .A(n24131), .B(n24132), .X(n39354) );
  nand_x1_sg U43700 ( .A(n23852), .B(n23853), .X(n39355) );
  nand_x1_sg U43701 ( .A(n24410), .B(n24411), .X(n39356) );
  nand_x1_sg U43702 ( .A(n24967), .B(n24968), .X(n39357) );
  nand_x1_sg U43703 ( .A(n24688), .B(n24689), .X(n39358) );
  nand_x1_sg U43704 ( .A(n25246), .B(n25247), .X(n39359) );
  nand_x1_sg U43705 ( .A(n25802), .B(n25803), .X(n39360) );
  nand_x1_sg U43706 ( .A(n25525), .B(n25526), .X(n39361) );
  nand_x1_sg U43707 ( .A(n26640), .B(n26641), .X(n39362) );
  nand_x1_sg U43708 ( .A(n26362), .B(n26363), .X(n39363) );
  nand_x1_sg U43709 ( .A(n26039), .B(n26040), .X(n39364) );
  inv_x1_sg U43710 ( .A(n41777), .X(n39365) );
  inv_x1_sg U43711 ( .A(n39365), .X(n39366) );
  inv_x1_sg U43712 ( .A(n41776), .X(n39367) );
  inv_x1_sg U43713 ( .A(n39367), .X(n39368) );
  inv_x1_sg U43714 ( .A(n41775), .X(n39369) );
  inv_x1_sg U43715 ( .A(n39369), .X(n39370) );
  inv_x1_sg U43716 ( .A(n41774), .X(n39371) );
  inv_x1_sg U43717 ( .A(n39371), .X(n39372) );
  inv_x1_sg U43718 ( .A(n41773), .X(n39373) );
  inv_x1_sg U43719 ( .A(n39373), .X(n39374) );
  inv_x1_sg U43720 ( .A(n41772), .X(n39375) );
  inv_x1_sg U43721 ( .A(n39375), .X(n39376) );
  inv_x1_sg U43722 ( .A(n41771), .X(n39377) );
  inv_x1_sg U43723 ( .A(n39377), .X(n39378) );
  inv_x1_sg U43724 ( .A(n41770), .X(n39379) );
  inv_x1_sg U43725 ( .A(n39379), .X(n39380) );
  inv_x1_sg U43726 ( .A(n41769), .X(n39381) );
  inv_x1_sg U43727 ( .A(n39381), .X(n39382) );
  inv_x1_sg U43728 ( .A(n41768), .X(n39383) );
  inv_x1_sg U43729 ( .A(n39383), .X(n39384) );
  inv_x1_sg U43730 ( .A(n41767), .X(n39385) );
  inv_x1_sg U43731 ( .A(n39385), .X(n39386) );
  inv_x1_sg U43732 ( .A(n41766), .X(n39387) );
  inv_x1_sg U43733 ( .A(n39387), .X(n39388) );
  inv_x1_sg U43734 ( .A(n41755), .X(n39389) );
  inv_x1_sg U43735 ( .A(n39389), .X(n39390) );
  inv_x1_sg U43736 ( .A(n39288), .X(n39391) );
  inv_x1_sg U43737 ( .A(n41507), .X(n39392) );
  inv_x1_sg U43738 ( .A(n39400), .X(n39393) );
  inv_x1_sg U43739 ( .A(n41504), .X(n39394) );
  inv_x1_sg U43740 ( .A(n39201), .X(n39395) );
  inv_x1_sg U43741 ( .A(n41505), .X(n39396) );
  inv_x1_sg U43742 ( .A(n42387), .X(n39397) );
  inv_x1_sg U43743 ( .A(n39397), .X(n39398) );
  inv_x1_sg U43744 ( .A(n39397), .X(n39399) );
  inv_x1_sg U43745 ( .A(n39398), .X(n39400) );
  inv_x1_sg U43746 ( .A(n39398), .X(n39401) );
  inv_x1_sg U43747 ( .A(n41504), .X(n39402) );
  inv_x1_sg U43748 ( .A(n41507), .X(n39403) );
  inv_x1_sg U43749 ( .A(n39408), .X(n39404) );
  inv_x1_sg U43750 ( .A(n41506), .X(n39405) );
  inv_x1_sg U43751 ( .A(n39401), .X(n39406) );
  inv_x1_sg U43752 ( .A(n41506), .X(n39407) );
  inv_x1_sg U43753 ( .A(n39399), .X(n39408) );
  inv_x1_sg U43754 ( .A(n38814), .X(n39409) );
  inv_x1_sg U43755 ( .A(n39201), .X(n39410) );
  inv_x1_sg U43756 ( .A(n39201), .X(n39411) );
  inv_x1_sg U43757 ( .A(n39287), .X(n39412) );
  inv_x1_sg U43758 ( .A(n39427), .X(n39413) );
  inv_x1_sg U43759 ( .A(n39424), .X(n39414) );
  inv_x1_sg U43760 ( .A(n41485), .X(n39415) );
  inv_x1_sg U43761 ( .A(n39286), .X(n39416) );
  inv_x1_sg U43762 ( .A(n39427), .X(n39417) );
  inv_x1_sg U43763 ( .A(n41484), .X(n39418) );
  inv_x1_sg U43764 ( .A(n41487), .X(n39419) );
  inv_x1_sg U43765 ( .A(n41487), .X(n39420) );
  inv_x1_sg U43766 ( .A(n39428), .X(n39421) );
  inv_x1_sg U43767 ( .A(n41483), .X(n39422) );
  inv_x1_sg U43768 ( .A(n39422), .X(n39423) );
  inv_x1_sg U43769 ( .A(n39423), .X(n39424) );
  inv_x1_sg U43770 ( .A(n41486), .X(n39425) );
  inv_x1_sg U43771 ( .A(n41485), .X(n39426) );
  inv_x1_sg U43772 ( .A(n39285), .X(n39427) );
  inv_x1_sg U43773 ( .A(n41483), .X(n39428) );
  inv_x1_sg U43774 ( .A(n41486), .X(n39429) );
  inv_x1_sg U43775 ( .A(n39287), .X(n39430) );
  inv_x1_sg U43776 ( .A(n39768), .X(n39431) );
  inv_x1_sg U43777 ( .A(n41477), .X(n39432) );
  inv_x1_sg U43778 ( .A(n5954), .X(n39433) );
  inv_x1_sg U43779 ( .A(n41416), .X(n39434) );
  inv_x1_sg U43780 ( .A(n39433), .X(n39435) );
  inv_x1_sg U43781 ( .A(n39200), .X(n39436) );
  inv_x1_sg U43782 ( .A(n39651), .X(n39437) );
  inv_x1_sg U43783 ( .A(n42376), .X(n39438) );
  inv_x1_sg U43784 ( .A(n41374), .X(n39439) );
  inv_x1_sg U43785 ( .A(n39438), .X(n39440) );
  inv_x1_sg U43786 ( .A(n42327), .X(n39441) );
  inv_x1_sg U43787 ( .A(n41369), .X(n39442) );
  inv_x1_sg U43788 ( .A(n39441), .X(n39443) );
  inv_x1_sg U43789 ( .A(n42386), .X(n39444) );
  inv_x1_sg U43790 ( .A(n41364), .X(n39445) );
  inv_x1_sg U43791 ( .A(n39444), .X(n39446) );
  inv_x1_sg U43792 ( .A(n42374), .X(n39447) );
  inv_x1_sg U43793 ( .A(n41359), .X(n39448) );
  inv_x1_sg U43794 ( .A(n39447), .X(n39449) );
  inv_x1_sg U43795 ( .A(n42373), .X(n39450) );
  inv_x1_sg U43796 ( .A(n41354), .X(n39451) );
  inv_x1_sg U43797 ( .A(n39450), .X(n39452) );
  inv_x1_sg U43798 ( .A(n42371), .X(n39453) );
  inv_x1_sg U43799 ( .A(n41349), .X(n39454) );
  inv_x1_sg U43800 ( .A(n39453), .X(n39455) );
  inv_x1_sg U43801 ( .A(n23409), .X(n39456) );
  inv_x1_sg U43802 ( .A(n41344), .X(n39457) );
  inv_x1_sg U43803 ( .A(n39456), .X(n39458) );
  inv_x1_sg U43804 ( .A(n42375), .X(n39459) );
  inv_x1_sg U43805 ( .A(n41339), .X(n39460) );
  inv_x1_sg U43806 ( .A(n39459), .X(n39461) );
  inv_x1_sg U43807 ( .A(n24525), .X(n39462) );
  inv_x1_sg U43808 ( .A(n41334), .X(n39463) );
  inv_x1_sg U43809 ( .A(n39462), .X(n39464) );
  inv_x1_sg U43810 ( .A(n24803), .X(n39465) );
  inv_x1_sg U43811 ( .A(n41329), .X(n39466) );
  inv_x1_sg U43812 ( .A(n39465), .X(n39467) );
  inv_x1_sg U43813 ( .A(n25082), .X(n39468) );
  inv_x1_sg U43814 ( .A(n41324), .X(n39469) );
  inv_x1_sg U43815 ( .A(n39468), .X(n39470) );
  inv_x1_sg U43816 ( .A(n41574), .X(n39471) );
  inv_x1_sg U43817 ( .A(n41319), .X(n39472) );
  inv_x1_sg U43818 ( .A(n39471), .X(n39473) );
  inv_x1_sg U43819 ( .A(n38980), .X(n39474) );
  inv_x1_sg U43820 ( .A(n41314), .X(n39475) );
  inv_x1_sg U43821 ( .A(n41314), .X(n39476) );
  inv_x1_sg U43822 ( .A(n39199), .X(n39477) );
  inv_x1_sg U43823 ( .A(n39655), .X(n39478) );
  inv_x1_sg U43824 ( .A(n41298), .X(n39479) );
  inv_x1_sg U43825 ( .A(n39135), .X(n39480) );
  inv_x1_sg U43826 ( .A(n41294), .X(n39481) );
  inv_x1_sg U43827 ( .A(n41294), .X(n39482) );
  inv_x1_sg U43828 ( .A(n39769), .X(n39483) );
  inv_x1_sg U43829 ( .A(n38986), .X(n39484) );
  inv_x1_sg U43830 ( .A(reg_num[1]), .X(n39485) );
  inv_x1_sg U43831 ( .A(n39485), .X(n39486) );
  inv_x1_sg U43832 ( .A(n39683), .X(n39487) );
  inv_x1_sg U43833 ( .A(n39686), .X(n39488) );
  inv_x1_sg U43834 ( .A(n39689), .X(n39489) );
  inv_x1_sg U43835 ( .A(n39692), .X(n39490) );
  inv_x1_sg U43836 ( .A(n39695), .X(n39491) );
  inv_x1_sg U43837 ( .A(n39698), .X(n39492) );
  inv_x1_sg U43838 ( .A(n39701), .X(n39493) );
  inv_x1_sg U43839 ( .A(n39704), .X(n39494) );
  inv_x1_sg U43840 ( .A(n39707), .X(n39495) );
  inv_x1_sg U43841 ( .A(n39710), .X(n39496) );
  inv_x1_sg U43842 ( .A(n39713), .X(n39497) );
  inv_x1_sg U43843 ( .A(n39716), .X(n39498) );
  inv_x1_sg U43844 ( .A(n39719), .X(n39499) );
  inv_x1_sg U43845 ( .A(n39722), .X(n39500) );
  inv_x1_sg U43846 ( .A(n42369), .X(n39501) );
  inv_x1_sg U43847 ( .A(n39501), .X(n39502) );
  inv_x1_sg U43848 ( .A(n42337), .X(n39503) );
  inv_x1_sg U43849 ( .A(n39503), .X(n39504) );
  nand_x1_sg U43850 ( .A(n41988), .B(n23302), .X(n39505) );
  nand_x1_sg U43851 ( .A(n41988), .B(n23302), .X(n9110) );
  nand_x1_sg U43852 ( .A(n41987), .B(n23022), .X(n39506) );
  nand_x1_sg U43853 ( .A(n41987), .B(n23022), .X(n8292) );
  nand_x1_sg U43854 ( .A(n41989), .B(n23581), .X(n39507) );
  nand_x1_sg U43855 ( .A(n41989), .B(n23581), .X(n9930) );
  nand_x1_sg U43856 ( .A(n41991), .B(n24139), .X(n39508) );
  nand_x1_sg U43857 ( .A(n41991), .B(n24139), .X(n11568) );
  nand_x1_sg U43858 ( .A(n41990), .B(n23860), .X(n39509) );
  nand_x1_sg U43859 ( .A(n41990), .B(n23860), .X(n10749) );
  nand_x1_sg U43860 ( .A(n41993), .B(n24696), .X(n39510) );
  nand_x1_sg U43861 ( .A(n41993), .B(n24696), .X(n13206) );
  nand_x1_sg U43862 ( .A(n41992), .B(n24418), .X(n39511) );
  nand_x1_sg U43863 ( .A(n41992), .B(n24418), .X(n12387) );
  nand_x1_sg U43864 ( .A(n41995), .B(n25254), .X(n39512) );
  nand_x1_sg U43865 ( .A(n41995), .B(n25254), .X(n14844) );
  nand_x1_sg U43866 ( .A(n41994), .B(n24975), .X(n39513) );
  nand_x1_sg U43867 ( .A(n41994), .B(n24975), .X(n14025) );
  nand_x1_sg U43868 ( .A(n41997), .B(n25810), .X(n39514) );
  nand_x1_sg U43869 ( .A(n41997), .B(n25810), .X(n16482) );
  nand_x1_sg U43870 ( .A(n41996), .B(n25533), .X(n39515) );
  nand_x1_sg U43871 ( .A(n41996), .B(n25533), .X(n15663) );
  nand_x1_sg U43872 ( .A(n41999), .B(n26370), .X(n39516) );
  nand_x1_sg U43873 ( .A(n41999), .B(n26370), .X(n18120) );
  nand_x1_sg U43874 ( .A(n41998), .B(n26648), .X(n39517) );
  nand_x1_sg U43875 ( .A(n41998), .B(n26648), .X(n18941) );
  nand_x1_sg U43876 ( .A(n23329), .B(n23330), .X(n39518) );
  nand_x1_sg U43877 ( .A(n23329), .B(n23330), .X(n42344) );
  nand_x1_sg U43878 ( .A(n23049), .B(n23050), .X(n39519) );
  nand_x1_sg U43879 ( .A(n23049), .B(n23050), .X(n42345) );
  nand_x1_sg U43880 ( .A(n26069), .B(n26070), .X(n39520) );
  nand_x1_sg U43881 ( .A(n26069), .B(n26070), .X(n42336) );
  nand_x1_sg U43882 ( .A(n24445), .B(n24446), .X(n39521) );
  nand_x1_sg U43883 ( .A(n24445), .B(n24446), .X(n42352) );
  nand_x1_sg U43884 ( .A(n24166), .B(n24167), .X(n39522) );
  nand_x1_sg U43885 ( .A(n24166), .B(n24167), .X(n42353) );
  nand_x1_sg U43886 ( .A(n23887), .B(n23888), .X(n39523) );
  nand_x1_sg U43887 ( .A(n23887), .B(n23888), .X(n42354) );
  nand_x1_sg U43888 ( .A(n23608), .B(n23609), .X(n39524) );
  nand_x1_sg U43889 ( .A(n23608), .B(n23609), .X(n42355) );
  nand_x1_sg U43890 ( .A(n25560), .B(n25561), .X(n39525) );
  nand_x1_sg U43891 ( .A(n25560), .B(n25561), .X(n42348) );
  nand_x1_sg U43892 ( .A(n25281), .B(n25282), .X(n39526) );
  nand_x1_sg U43893 ( .A(n25281), .B(n25282), .X(n42349) );
  nand_x1_sg U43894 ( .A(n25002), .B(n25003), .X(n39527) );
  nand_x1_sg U43895 ( .A(n25002), .B(n25003), .X(n42350) );
  nand_x1_sg U43896 ( .A(n24723), .B(n24724), .X(n39528) );
  nand_x1_sg U43897 ( .A(n24723), .B(n24724), .X(n42351) );
  nand_x1_sg U43898 ( .A(n26675), .B(n26676), .X(n39529) );
  nand_x1_sg U43899 ( .A(n26675), .B(n26676), .X(n42346) );
  nand_x1_sg U43900 ( .A(n26397), .B(n26398), .X(n39530) );
  nand_x1_sg U43901 ( .A(n26397), .B(n26398), .X(n42356) );
  nand_x1_sg U43902 ( .A(n25837), .B(n25838), .X(n39531) );
  nand_x1_sg U43903 ( .A(n25837), .B(n25838), .X(n42347) );
  nand_x1_sg U43904 ( .A(n23035), .B(n23036), .X(n39532) );
  nand_x1_sg U43905 ( .A(n23035), .B(n23036), .X(n42358) );
  nand_x1_sg U43906 ( .A(n23315), .B(n23316), .X(n39533) );
  nand_x1_sg U43907 ( .A(n23315), .B(n23316), .X(n42357) );
  nand_x1_sg U43908 ( .A(n23594), .B(n23595), .X(n39534) );
  nand_x1_sg U43909 ( .A(n23594), .B(n23595), .X(n42368) );
  nand_x1_sg U43910 ( .A(n23873), .B(n23874), .X(n39535) );
  nand_x1_sg U43911 ( .A(n23873), .B(n23874), .X(n42367) );
  nand_x1_sg U43912 ( .A(n24152), .B(n24153), .X(n39536) );
  nand_x1_sg U43913 ( .A(n24152), .B(n24153), .X(n42366) );
  nand_x1_sg U43914 ( .A(n24431), .B(n24432), .X(n39537) );
  nand_x1_sg U43915 ( .A(n24431), .B(n24432), .X(n42365) );
  nand_x1_sg U43916 ( .A(n24709), .B(n24710), .X(n39538) );
  nand_x1_sg U43917 ( .A(n24709), .B(n24710), .X(n42364) );
  nand_x1_sg U43918 ( .A(n24988), .B(n24989), .X(n39539) );
  nand_x1_sg U43919 ( .A(n24988), .B(n24989), .X(n42363) );
  nand_x1_sg U43920 ( .A(n25267), .B(n25268), .X(n39540) );
  nand_x1_sg U43921 ( .A(n25267), .B(n25268), .X(n42362) );
  nand_x1_sg U43922 ( .A(n25546), .B(n25547), .X(n39541) );
  nand_x1_sg U43923 ( .A(n25546), .B(n25547), .X(n42361) );
  nand_x1_sg U43924 ( .A(n25823), .B(n25824), .X(n39542) );
  nand_x1_sg U43925 ( .A(n25823), .B(n25824), .X(n42360) );
  nand_x1_sg U43926 ( .A(n26383), .B(n26384), .X(n39543) );
  nand_x1_sg U43927 ( .A(n26383), .B(n26384), .X(n17636) );
  nand_x1_sg U43928 ( .A(n26661), .B(n26662), .X(n39544) );
  nand_x1_sg U43929 ( .A(n26661), .B(n26662), .X(n42359) );
  inv_x1_sg U43930 ( .A(n42236), .X(n39545) );
  inv_x1_sg U43931 ( .A(n42321), .X(n39546) );
  inv_x1_sg U43932 ( .A(n42320), .X(n39547) );
  inv_x1_sg U43933 ( .A(n42324), .X(n39548) );
  inv_x1_sg U43934 ( .A(n42323), .X(n39549) );
  inv_x1_sg U43935 ( .A(n42322), .X(n39550) );
  inv_x1_sg U43936 ( .A(n15225), .X(n39551) );
  inv_x1_sg U43937 ( .A(n16044), .X(n39552) );
  inv_x1_sg U43938 ( .A(n14406), .X(n39553) );
  inv_x1_sg U43939 ( .A(n11949), .X(n39554) );
  inv_x1_sg U43940 ( .A(n12768), .X(n39555) );
  inv_x1_sg U43941 ( .A(n13587), .X(n39556) );
  inv_x1_sg U43942 ( .A(n10311), .X(n39557) );
  inv_x1_sg U43943 ( .A(n11130), .X(n39558) );
  inv_x1_sg U43944 ( .A(n41708), .X(n39559) );
  inv_x1_sg U43945 ( .A(n39559), .X(n39560) );
  inv_x1_sg U43946 ( .A(n39559), .X(n39561) );
  inv_x1_sg U43947 ( .A(n41707), .X(n39562) );
  inv_x1_sg U43948 ( .A(n39562), .X(n39563) );
  inv_x1_sg U43949 ( .A(n39562), .X(n39564) );
  inv_x1_sg U43950 ( .A(n41706), .X(n39565) );
  inv_x1_sg U43951 ( .A(n39565), .X(n39566) );
  inv_x1_sg U43952 ( .A(n39565), .X(n39567) );
  inv_x1_sg U43953 ( .A(n41705), .X(n39568) );
  inv_x1_sg U43954 ( .A(n39568), .X(n39569) );
  inv_x1_sg U43955 ( .A(n39568), .X(n39570) );
  inv_x1_sg U43956 ( .A(n41704), .X(n39571) );
  inv_x1_sg U43957 ( .A(n39571), .X(n39572) );
  inv_x1_sg U43958 ( .A(n39571), .X(n39573) );
  inv_x1_sg U43959 ( .A(n41703), .X(n39574) );
  inv_x1_sg U43960 ( .A(n39574), .X(n39575) );
  inv_x1_sg U43961 ( .A(n39574), .X(n39576) );
  inv_x1_sg U43962 ( .A(n41702), .X(n39577) );
  inv_x1_sg U43963 ( .A(n39577), .X(n39578) );
  inv_x1_sg U43964 ( .A(n39577), .X(n39579) );
  inv_x1_sg U43965 ( .A(n41701), .X(n39580) );
  inv_x1_sg U43966 ( .A(n39580), .X(n39581) );
  inv_x1_sg U43967 ( .A(n39580), .X(n39582) );
  inv_x1_sg U43968 ( .A(n41700), .X(n39583) );
  inv_x1_sg U43969 ( .A(n39583), .X(n39584) );
  inv_x1_sg U43970 ( .A(n39583), .X(n39585) );
  inv_x1_sg U43971 ( .A(n41699), .X(n39586) );
  inv_x1_sg U43972 ( .A(n39586), .X(n39587) );
  inv_x1_sg U43973 ( .A(n39586), .X(n39588) );
  inv_x1_sg U43974 ( .A(n41698), .X(n39589) );
  inv_x1_sg U43975 ( .A(n39589), .X(n39590) );
  inv_x1_sg U43976 ( .A(n39589), .X(n39591) );
  inv_x1_sg U43977 ( .A(n41697), .X(n39592) );
  inv_x1_sg U43978 ( .A(n39592), .X(n39593) );
  inv_x1_sg U43979 ( .A(n39592), .X(n39594) );
  inv_x1_sg U43980 ( .A(n41696), .X(n39595) );
  inv_x1_sg U43981 ( .A(n39595), .X(n39596) );
  inv_x1_sg U43982 ( .A(n39595), .X(n39597) );
  inv_x1_sg U43983 ( .A(n41695), .X(n39598) );
  inv_x1_sg U43984 ( .A(n39598), .X(n39599) );
  inv_x1_sg U43985 ( .A(n39598), .X(n39600) );
  inv_x1_sg U43986 ( .A(n41694), .X(n39601) );
  inv_x1_sg U43987 ( .A(n39601), .X(n39602) );
  inv_x1_sg U43988 ( .A(n39601), .X(n39603) );
  inv_x1_sg U43989 ( .A(n41661), .X(n39604) );
  inv_x1_sg U43990 ( .A(n39604), .X(n39605) );
  inv_x1_sg U43991 ( .A(n39604), .X(n39606) );
  inv_x1_sg U43992 ( .A(n41646), .X(n39607) );
  inv_x1_sg U43993 ( .A(n39607), .X(n39608) );
  inv_x1_sg U43994 ( .A(n39607), .X(n39609) );
  inv_x1_sg U43995 ( .A(n41645), .X(n39610) );
  inv_x1_sg U43996 ( .A(n39610), .X(n39611) );
  inv_x1_sg U43997 ( .A(n39610), .X(n39612) );
  inv_x1_sg U43998 ( .A(n41644), .X(n39613) );
  inv_x1_sg U43999 ( .A(n39613), .X(n39614) );
  inv_x1_sg U44000 ( .A(n39613), .X(n39615) );
  inv_x1_sg U44001 ( .A(n41643), .X(n39616) );
  inv_x1_sg U44002 ( .A(n39616), .X(n39617) );
  inv_x1_sg U44003 ( .A(n39616), .X(n39618) );
  inv_x1_sg U44004 ( .A(n41642), .X(n39619) );
  inv_x1_sg U44005 ( .A(n39619), .X(n39620) );
  inv_x1_sg U44006 ( .A(n39619), .X(n39621) );
  inv_x1_sg U44007 ( .A(n41641), .X(n39622) );
  inv_x1_sg U44008 ( .A(n39622), .X(n39623) );
  inv_x1_sg U44009 ( .A(n39622), .X(n39624) );
  inv_x1_sg U44010 ( .A(n41640), .X(n39625) );
  inv_x1_sg U44011 ( .A(n39625), .X(n39626) );
  inv_x1_sg U44012 ( .A(n39625), .X(n39627) );
  inv_x1_sg U44013 ( .A(n41639), .X(n39628) );
  inv_x1_sg U44014 ( .A(n39628), .X(n39629) );
  inv_x1_sg U44015 ( .A(n39628), .X(n39630) );
  inv_x1_sg U44016 ( .A(n41638), .X(n39631) );
  inv_x1_sg U44017 ( .A(n39631), .X(n39632) );
  inv_x1_sg U44018 ( .A(n39631), .X(n39633) );
  inv_x1_sg U44019 ( .A(n41637), .X(n39634) );
  inv_x1_sg U44020 ( .A(n39634), .X(n39635) );
  inv_x1_sg U44021 ( .A(n39634), .X(n39636) );
  inv_x1_sg U44022 ( .A(n41636), .X(n39637) );
  inv_x1_sg U44023 ( .A(n39637), .X(n39638) );
  inv_x1_sg U44024 ( .A(n39637), .X(n39639) );
  inv_x1_sg U44025 ( .A(n41635), .X(n39640) );
  inv_x1_sg U44026 ( .A(n39640), .X(n39641) );
  inv_x1_sg U44027 ( .A(n39640), .X(n39642) );
  inv_x1_sg U44028 ( .A(n41634), .X(n39643) );
  inv_x1_sg U44029 ( .A(n39643), .X(n39644) );
  inv_x1_sg U44030 ( .A(n39643), .X(n39645) );
  inv_x1_sg U44031 ( .A(n41633), .X(n39646) );
  inv_x1_sg U44032 ( .A(n39646), .X(n39647) );
  inv_x1_sg U44033 ( .A(n39646), .X(n39648) );
  inv_x1_sg U44034 ( .A(n38986), .X(n39649) );
  inv_x1_sg U44035 ( .A(n38986), .X(n39650) );
  inv_x1_sg U44036 ( .A(n41949), .X(n39651) );
  inv_x1_sg U44037 ( .A(n41949), .X(n39652) );
  inv_x1_sg U44038 ( .A(n39200), .X(n39653) );
  inv_x1_sg U44039 ( .A(n39651), .X(n39654) );
  inv_x1_sg U44040 ( .A(n42377), .X(n39655) );
  inv_x1_sg U44041 ( .A(n42377), .X(n39656) );
  inv_x1_sg U44042 ( .A(n39199), .X(n39657) );
  inv_x1_sg U44043 ( .A(n39655), .X(n39658) );
  inv_x1_sg U44044 ( .A(n41303), .X(n39659) );
  inv_x1_sg U44045 ( .A(n41303), .X(n39660) );
  nand_x1_sg U44046 ( .A(n26057), .B(n26058), .X(n39661) );
  nand_x1_sg U44047 ( .A(n26045), .B(n26046), .X(n39662) );
  inv_x1_sg U44048 ( .A(n16850), .X(n39679) );
  inv_x1_sg U44049 ( .A(n40611), .X(n39680) );
  inv_x1_sg U44050 ( .A(n16850), .X(n39681) );
  inv_x1_sg U44051 ( .A(n41806), .X(n39682) );
  inv_x1_sg U44052 ( .A(n39682), .X(n39683) );
  inv_x1_sg U44053 ( .A(n39682), .X(n39684) );
  inv_x1_sg U44054 ( .A(n41804), .X(n39685) );
  inv_x1_sg U44055 ( .A(n39685), .X(n39686) );
  inv_x1_sg U44056 ( .A(n39685), .X(n39687) );
  inv_x1_sg U44057 ( .A(n41802), .X(n39688) );
  inv_x1_sg U44058 ( .A(n39688), .X(n39689) );
  inv_x1_sg U44059 ( .A(n39688), .X(n39690) );
  inv_x1_sg U44060 ( .A(n41800), .X(n39691) );
  inv_x1_sg U44061 ( .A(n39691), .X(n39692) );
  inv_x1_sg U44062 ( .A(n39691), .X(n39693) );
  inv_x1_sg U44063 ( .A(n41798), .X(n39694) );
  inv_x1_sg U44064 ( .A(n39694), .X(n39695) );
  inv_x1_sg U44065 ( .A(n39694), .X(n39696) );
  inv_x1_sg U44066 ( .A(n41796), .X(n39697) );
  inv_x1_sg U44067 ( .A(n39697), .X(n39698) );
  inv_x1_sg U44068 ( .A(n39697), .X(n39699) );
  inv_x1_sg U44069 ( .A(n41794), .X(n39700) );
  inv_x1_sg U44070 ( .A(n39700), .X(n39701) );
  inv_x1_sg U44071 ( .A(n39700), .X(n39702) );
  inv_x1_sg U44072 ( .A(n41792), .X(n39703) );
  inv_x1_sg U44073 ( .A(n39703), .X(n39704) );
  inv_x1_sg U44074 ( .A(n39703), .X(n39705) );
  inv_x1_sg U44075 ( .A(n41790), .X(n39706) );
  inv_x1_sg U44076 ( .A(n39706), .X(n39707) );
  inv_x1_sg U44077 ( .A(n39706), .X(n39708) );
  inv_x1_sg U44078 ( .A(n41788), .X(n39709) );
  inv_x1_sg U44079 ( .A(n39709), .X(n39710) );
  inv_x1_sg U44080 ( .A(n39709), .X(n39711) );
  inv_x1_sg U44081 ( .A(n41786), .X(n39712) );
  inv_x1_sg U44082 ( .A(n39712), .X(n39713) );
  inv_x1_sg U44083 ( .A(n39712), .X(n39714) );
  inv_x1_sg U44084 ( .A(n41784), .X(n39715) );
  inv_x1_sg U44085 ( .A(n39715), .X(n39716) );
  inv_x1_sg U44086 ( .A(n39715), .X(n39717) );
  inv_x1_sg U44087 ( .A(n41782), .X(n39718) );
  inv_x1_sg U44088 ( .A(n39718), .X(n39719) );
  inv_x1_sg U44089 ( .A(n39718), .X(n39720) );
  inv_x1_sg U44090 ( .A(n41780), .X(n39721) );
  inv_x1_sg U44091 ( .A(n39721), .X(n39722) );
  inv_x1_sg U44092 ( .A(n39721), .X(n39723) );
  inv_x1_sg U44093 ( .A(n41709), .X(n39724) );
  inv_x1_sg U44094 ( .A(n39724), .X(n39725) );
  inv_x1_sg U44095 ( .A(n39724), .X(n39726) );
  inv_x1_sg U44096 ( .A(n39479), .X(n39727) );
  inv_x1_sg U44097 ( .A(n41299), .X(n39728) );
  inv_x1_sg U44098 ( .A(n41657), .X(n39729) );
  inv_x1_sg U44099 ( .A(n39729), .X(n39730) );
  inv_x1_sg U44100 ( .A(n39729), .X(n39731) );
  inv_x1_sg U44101 ( .A(n41656), .X(n39732) );
  inv_x1_sg U44102 ( .A(n39732), .X(n39733) );
  inv_x1_sg U44103 ( .A(n39732), .X(n39734) );
  inv_x1_sg U44104 ( .A(n41651), .X(n39735) );
  inv_x1_sg U44105 ( .A(n39735), .X(n39736) );
  inv_x1_sg U44106 ( .A(n39735), .X(n39737) );
  inv_x1_sg U44107 ( .A(n41650), .X(n39738) );
  inv_x1_sg U44108 ( .A(n39738), .X(n39739) );
  inv_x1_sg U44109 ( .A(n39738), .X(n39740) );
  inv_x1_sg U44110 ( .A(n41649), .X(n39741) );
  inv_x1_sg U44111 ( .A(n39741), .X(n39742) );
  inv_x1_sg U44112 ( .A(n39741), .X(n39743) );
  inv_x1_sg U44113 ( .A(n41648), .X(n39744) );
  inv_x1_sg U44114 ( .A(n39744), .X(n39745) );
  inv_x1_sg U44115 ( .A(n39744), .X(n39746) );
  inv_x1_sg U44116 ( .A(n41655), .X(n39747) );
  inv_x1_sg U44117 ( .A(n39747), .X(n39748) );
  inv_x1_sg U44118 ( .A(n39747), .X(n39749) );
  inv_x1_sg U44119 ( .A(n41654), .X(n39750) );
  inv_x1_sg U44120 ( .A(n39750), .X(n39751) );
  inv_x1_sg U44121 ( .A(n39750), .X(n39752) );
  inv_x1_sg U44122 ( .A(n41653), .X(n39753) );
  inv_x1_sg U44123 ( .A(n39753), .X(n39754) );
  inv_x1_sg U44124 ( .A(n39753), .X(n39755) );
  inv_x1_sg U44125 ( .A(n41652), .X(n39756) );
  inv_x1_sg U44126 ( .A(n39756), .X(n39757) );
  inv_x1_sg U44127 ( .A(n39756), .X(n39758) );
  inv_x1_sg U44128 ( .A(n41659), .X(n39759) );
  inv_x1_sg U44129 ( .A(n39759), .X(n39760) );
  inv_x1_sg U44130 ( .A(n39759), .X(n39761) );
  inv_x1_sg U44131 ( .A(n41647), .X(n39762) );
  inv_x1_sg U44132 ( .A(n39762), .X(n39763) );
  inv_x1_sg U44133 ( .A(n39762), .X(n39764) );
  inv_x1_sg U44134 ( .A(n41658), .X(n39765) );
  inv_x1_sg U44135 ( .A(n39765), .X(n39766) );
  inv_x1_sg U44136 ( .A(n39765), .X(n39767) );
  inv_x1_sg U44137 ( .A(n42388), .X(n39768) );
  inv_x1_sg U44138 ( .A(n42388), .X(n39769) );
  nand_x1_sg U44139 ( .A(n26099), .B(n42120), .X(n39770) );
  nand_x1_sg U44140 ( .A(n26099), .B(n42120), .X(n39771) );
  nand_x1_sg U44141 ( .A(n22772), .B(n22773), .X(n39772) );
  nand_x1_sg U44142 ( .A(n22772), .B(n22773), .X(n39773) );
  nand_x1_sg U44143 ( .A(n22772), .B(n22773), .X(n6971) );
  nand_x1_sg U44144 ( .A(n26051), .B(n26052), .X(n39774) );
  nand_x1_sg U44145 ( .A(n26051), .B(n26052), .X(n39775) );
  nand_x1_sg U44146 ( .A(n26051), .B(n26052), .X(n42235) );
  nand_x1_sg U44147 ( .A(n26654), .B(n26655), .X(n39776) );
  nand_x1_sg U44148 ( .A(n26654), .B(n26655), .X(n39777) );
  nand_x1_sg U44149 ( .A(n26654), .B(n26655), .X(n42313) );
  nand_x1_sg U44150 ( .A(n25816), .B(n25817), .X(n39778) );
  nand_x1_sg U44151 ( .A(n25816), .B(n25817), .X(n39779) );
  nand_x1_sg U44152 ( .A(n25816), .B(n25817), .X(n42314) );
  nand_x1_sg U44153 ( .A(n26376), .B(n26377), .X(n39780) );
  nand_x1_sg U44154 ( .A(n26376), .B(n26377), .X(n39781) );
  nand_x1_sg U44155 ( .A(n26376), .B(n26377), .X(n18091) );
  nand_x1_sg U44156 ( .A(n25260), .B(n25261), .X(n39782) );
  nand_x1_sg U44157 ( .A(n25260), .B(n25261), .X(n39783) );
  nand_x1_sg U44158 ( .A(n25260), .B(n25261), .X(n42315) );
  nand_x1_sg U44159 ( .A(n25539), .B(n25540), .X(n39784) );
  nand_x1_sg U44160 ( .A(n25539), .B(n25540), .X(n39785) );
  nand_x1_sg U44161 ( .A(n25539), .B(n25540), .X(n15634) );
  nand_x1_sg U44162 ( .A(n24702), .B(n24703), .X(n39786) );
  nand_x1_sg U44163 ( .A(n24702), .B(n24703), .X(n39787) );
  nand_x1_sg U44164 ( .A(n24702), .B(n24703), .X(n42316) );
  nand_x1_sg U44165 ( .A(n24981), .B(n24982), .X(n39788) );
  nand_x1_sg U44166 ( .A(n24981), .B(n24982), .X(n39789) );
  nand_x1_sg U44167 ( .A(n24981), .B(n24982), .X(n13996) );
  nand_x1_sg U44168 ( .A(n24145), .B(n24146), .X(n39790) );
  nand_x1_sg U44169 ( .A(n24145), .B(n24146), .X(n39791) );
  nand_x1_sg U44170 ( .A(n24145), .B(n24146), .X(n42317) );
  nand_x1_sg U44171 ( .A(n24424), .B(n24425), .X(n39792) );
  nand_x1_sg U44172 ( .A(n24424), .B(n24425), .X(n39793) );
  nand_x1_sg U44173 ( .A(n24424), .B(n24425), .X(n12358) );
  nand_x1_sg U44174 ( .A(n23587), .B(n23588), .X(n39794) );
  nand_x1_sg U44175 ( .A(n23587), .B(n23588), .X(n39795) );
  nand_x1_sg U44176 ( .A(n23587), .B(n23588), .X(n42318) );
  nand_x1_sg U44177 ( .A(n23866), .B(n23867), .X(n39796) );
  nand_x1_sg U44178 ( .A(n23866), .B(n23867), .X(n39797) );
  nand_x1_sg U44179 ( .A(n23866), .B(n23867), .X(n10720) );
  nand_x1_sg U44180 ( .A(n23028), .B(n23029), .X(n39798) );
  nand_x1_sg U44181 ( .A(n23028), .B(n23029), .X(n39799) );
  nand_x1_sg U44182 ( .A(n23028), .B(n23029), .X(n42319) );
  nand_x1_sg U44183 ( .A(n23308), .B(n23309), .X(n39800) );
  nand_x1_sg U44184 ( .A(n23308), .B(n23309), .X(n39801) );
  nand_x1_sg U44185 ( .A(n23308), .B(n23309), .X(n9081) );
  nand_x1_sg U44186 ( .A(n22751), .B(n22752), .X(n39802) );
  nand_x1_sg U44187 ( .A(n22751), .B(n22752), .X(n39803) );
  nand_x1_sg U44188 ( .A(n22751), .B(n22752), .X(n7445) );
  nand_x1_sg U44189 ( .A(n22779), .B(n22780), .X(n39804) );
  nand_x1_sg U44190 ( .A(n22779), .B(n22780), .X(n39805) );
  nand_x1_sg U44191 ( .A(n26134), .B(n26135), .X(n39806) );
  nand_x1_sg U44192 ( .A(n26134), .B(n26135), .X(n39807) );
  nand_x1_sg U44193 ( .A(n26134), .B(n26135), .X(n16822) );
  inv_x1_sg U44194 ( .A(n41901), .X(n39808) );
  inv_x1_sg U44195 ( .A(n39808), .X(n39809) );
  inv_x1_sg U44196 ( .A(n39808), .X(n39810) );
  inv_x1_sg U44197 ( .A(n41899), .X(n39811) );
  inv_x1_sg U44198 ( .A(n39811), .X(n39812) );
  inv_x1_sg U44199 ( .A(n39811), .X(n39813) );
  inv_x1_sg U44200 ( .A(n41897), .X(n39814) );
  inv_x1_sg U44201 ( .A(n39814), .X(n39815) );
  inv_x1_sg U44202 ( .A(n39814), .X(n39816) );
  inv_x1_sg U44203 ( .A(n41895), .X(n39817) );
  inv_x1_sg U44204 ( .A(n39817), .X(n39818) );
  inv_x1_sg U44205 ( .A(n39817), .X(n39819) );
  inv_x1_sg U44206 ( .A(n41893), .X(n39820) );
  inv_x1_sg U44207 ( .A(n39820), .X(n39821) );
  inv_x1_sg U44208 ( .A(n39820), .X(n39822) );
  inv_x1_sg U44209 ( .A(n41891), .X(n39823) );
  inv_x1_sg U44210 ( .A(n39823), .X(n39824) );
  inv_x1_sg U44211 ( .A(n39823), .X(n39825) );
  inv_x1_sg U44212 ( .A(n41889), .X(n39826) );
  inv_x1_sg U44213 ( .A(n39826), .X(n39827) );
  inv_x1_sg U44214 ( .A(n39826), .X(n39828) );
  inv_x1_sg U44215 ( .A(n41887), .X(n39829) );
  inv_x1_sg U44216 ( .A(n39829), .X(n39830) );
  inv_x1_sg U44217 ( .A(n39829), .X(n39831) );
  inv_x1_sg U44218 ( .A(n41885), .X(n39832) );
  inv_x1_sg U44219 ( .A(n39832), .X(n39833) );
  inv_x1_sg U44220 ( .A(n39832), .X(n39834) );
  inv_x1_sg U44221 ( .A(n41883), .X(n39835) );
  inv_x1_sg U44222 ( .A(n39835), .X(n39836) );
  inv_x1_sg U44223 ( .A(n39835), .X(n39837) );
  inv_x1_sg U44224 ( .A(n41881), .X(n39838) );
  inv_x1_sg U44225 ( .A(n39838), .X(n39839) );
  inv_x1_sg U44226 ( .A(n39838), .X(n39840) );
  inv_x1_sg U44227 ( .A(n41879), .X(n39841) );
  inv_x1_sg U44228 ( .A(n39841), .X(n39842) );
  inv_x1_sg U44229 ( .A(n39841), .X(n39843) );
  inv_x1_sg U44230 ( .A(n41877), .X(n39844) );
  inv_x1_sg U44231 ( .A(n39844), .X(n39845) );
  inv_x1_sg U44232 ( .A(n39844), .X(n39846) );
  inv_x1_sg U44233 ( .A(n41875), .X(n39847) );
  inv_x1_sg U44234 ( .A(n39847), .X(n39848) );
  inv_x1_sg U44235 ( .A(n39847), .X(n39849) );
  inv_x1_sg U44236 ( .A(n42163), .X(n39850) );
  inv_x1_sg U44237 ( .A(n39931), .X(n39851) );
  inv_x1_sg U44238 ( .A(n39931), .X(n39852) );
  inv_x1_sg U44239 ( .A(n41691), .X(n39853) );
  inv_x1_sg U44240 ( .A(n39853), .X(n39854) );
  inv_x1_sg U44241 ( .A(n39853), .X(n39855) );
  inv_x1_sg U44242 ( .A(n41689), .X(n39856) );
  inv_x1_sg U44243 ( .A(n39856), .X(n39857) );
  inv_x1_sg U44244 ( .A(n39856), .X(n39858) );
  inv_x1_sg U44245 ( .A(n41687), .X(n39859) );
  inv_x1_sg U44246 ( .A(n39859), .X(n39860) );
  inv_x1_sg U44247 ( .A(n39859), .X(n39861) );
  inv_x1_sg U44248 ( .A(n41685), .X(n39862) );
  inv_x1_sg U44249 ( .A(n39862), .X(n39863) );
  inv_x1_sg U44250 ( .A(n39862), .X(n39864) );
  inv_x1_sg U44251 ( .A(n41683), .X(n39865) );
  inv_x1_sg U44252 ( .A(n39865), .X(n39866) );
  inv_x1_sg U44253 ( .A(n39865), .X(n39867) );
  inv_x1_sg U44254 ( .A(n41681), .X(n39868) );
  inv_x1_sg U44255 ( .A(n39868), .X(n39869) );
  inv_x1_sg U44256 ( .A(n39868), .X(n39870) );
  inv_x1_sg U44257 ( .A(n41679), .X(n39871) );
  inv_x1_sg U44258 ( .A(n39871), .X(n39872) );
  inv_x1_sg U44259 ( .A(n39871), .X(n39873) );
  inv_x1_sg U44260 ( .A(n41677), .X(n39874) );
  inv_x1_sg U44261 ( .A(n39874), .X(n39875) );
  inv_x1_sg U44262 ( .A(n39874), .X(n39876) );
  inv_x1_sg U44263 ( .A(n41675), .X(n39877) );
  inv_x1_sg U44264 ( .A(n39877), .X(n39878) );
  inv_x1_sg U44265 ( .A(n39877), .X(n39879) );
  inv_x1_sg U44266 ( .A(n41673), .X(n39880) );
  inv_x1_sg U44267 ( .A(n39880), .X(n39881) );
  inv_x1_sg U44268 ( .A(n39880), .X(n39882) );
  inv_x1_sg U44269 ( .A(n41671), .X(n39883) );
  inv_x1_sg U44270 ( .A(n39883), .X(n39884) );
  inv_x1_sg U44271 ( .A(n39883), .X(n39885) );
  inv_x1_sg U44272 ( .A(n41669), .X(n39886) );
  inv_x1_sg U44273 ( .A(n39886), .X(n39887) );
  inv_x1_sg U44274 ( .A(n39886), .X(n39888) );
  inv_x1_sg U44275 ( .A(n41667), .X(n39889) );
  inv_x1_sg U44276 ( .A(n39889), .X(n39890) );
  inv_x1_sg U44277 ( .A(n39889), .X(n39891) );
  inv_x1_sg U44278 ( .A(n41664), .X(n39892) );
  inv_x1_sg U44279 ( .A(n39892), .X(n39893) );
  inv_x1_sg U44280 ( .A(n39892), .X(n39894) );
  inv_x1_sg U44281 ( .A(n41662), .X(n39895) );
  inv_x1_sg U44282 ( .A(n39895), .X(n39896) );
  inv_x1_sg U44283 ( .A(n39895), .X(n39897) );
  inv_x1_sg U44284 ( .A(n39768), .X(n39898) );
  inv_x1_sg U44285 ( .A(n41477), .X(n39899) );
  inv_x1_sg U44286 ( .A(n41384), .X(n39900) );
  inv_x1_sg U44287 ( .A(n41379), .X(n39901) );
  inv_x1_sg U44288 ( .A(n38977), .X(n39902) );
  inv_x1_sg U44289 ( .A(n38977), .X(n39903) );
  inv_x1_sg U44290 ( .A(n38974), .X(n39904) );
  inv_x1_sg U44291 ( .A(n38974), .X(n39905) );
  inv_x1_sg U44292 ( .A(n38971), .X(n39906) );
  inv_x1_sg U44293 ( .A(n38971), .X(n39907) );
  inv_x1_sg U44294 ( .A(n38968), .X(n39908) );
  inv_x1_sg U44295 ( .A(n38968), .X(n39909) );
  inv_x1_sg U44296 ( .A(n38965), .X(n39910) );
  inv_x1_sg U44297 ( .A(n38965), .X(n39911) );
  inv_x1_sg U44298 ( .A(n38962), .X(n39912) );
  inv_x1_sg U44299 ( .A(n38962), .X(n39913) );
  inv_x1_sg U44300 ( .A(n38959), .X(n39914) );
  inv_x1_sg U44301 ( .A(n38959), .X(n39915) );
  inv_x1_sg U44302 ( .A(n38956), .X(n39916) );
  inv_x1_sg U44303 ( .A(n38956), .X(n39917) );
  inv_x1_sg U44304 ( .A(n38953), .X(n39918) );
  inv_x1_sg U44305 ( .A(n38953), .X(n39919) );
  inv_x1_sg U44306 ( .A(n38950), .X(n39920) );
  inv_x1_sg U44307 ( .A(n38950), .X(n39921) );
  inv_x1_sg U44308 ( .A(n38947), .X(n39922) );
  inv_x1_sg U44309 ( .A(n38947), .X(n39923) );
  inv_x1_sg U44310 ( .A(n38945), .X(n39924) );
  inv_x1_sg U44311 ( .A(n38945), .X(n39925) );
  inv_x1_sg U44312 ( .A(n41314), .X(n39926) );
  inv_x1_sg U44313 ( .A(n41314), .X(n39927) );
  inv_x1_sg U44314 ( .A(n39275), .X(n39928) );
  inv_x1_sg U44315 ( .A(n39274), .X(n39929) );
  nand_x1_sg U44316 ( .A(n22787), .B(n22788), .X(n39930) );
  nand_x1_sg U44317 ( .A(n22787), .B(n22788), .X(n39931) );
  nand_x1_sg U44318 ( .A(n22787), .B(n22788), .X(n42163) );
  nand_x1_sg U44319 ( .A(n26075), .B(n26076), .X(n39932) );
  nand_x1_sg U44320 ( .A(n26075), .B(n26076), .X(n39933) );
  nand_x1_sg U44321 ( .A(n26075), .B(n26076), .X(n42236) );
  nand_x1_sg U44322 ( .A(n26404), .B(n26405), .X(n39934) );
  nand_x1_sg U44323 ( .A(n26404), .B(n26405), .X(n39935) );
  nand_x1_sg U44324 ( .A(n26404), .B(n26405), .X(n42321) );
  nand_x1_sg U44325 ( .A(n26682), .B(n26683), .X(n39936) );
  nand_x1_sg U44326 ( .A(n26682), .B(n26683), .X(n39937) );
  nand_x1_sg U44327 ( .A(n26682), .B(n26683), .X(n42320) );
  nand_x1_sg U44328 ( .A(n23056), .B(n23057), .X(n39938) );
  nand_x1_sg U44329 ( .A(n23056), .B(n23057), .X(n39939) );
  nand_x1_sg U44330 ( .A(n23056), .B(n23057), .X(n42324) );
  nand_x1_sg U44331 ( .A(n23336), .B(n23337), .X(n39940) );
  nand_x1_sg U44332 ( .A(n23336), .B(n23337), .X(n39941) );
  nand_x1_sg U44333 ( .A(n23336), .B(n23337), .X(n42323) );
  nand_x1_sg U44334 ( .A(n23615), .B(n23616), .X(n39942) );
  nand_x1_sg U44335 ( .A(n23615), .B(n23616), .X(n39943) );
  nand_x1_sg U44336 ( .A(n23615), .B(n23616), .X(n42322) );
  nand_x1_sg U44337 ( .A(n25567), .B(n25568), .X(n39944) );
  nand_x1_sg U44338 ( .A(n25567), .B(n25568), .X(n39945) );
  nand_x1_sg U44339 ( .A(n25567), .B(n25568), .X(n15225) );
  nand_x1_sg U44340 ( .A(n25844), .B(n25845), .X(n39946) );
  nand_x1_sg U44341 ( .A(n25844), .B(n25845), .X(n39947) );
  nand_x1_sg U44342 ( .A(n25844), .B(n25845), .X(n16044) );
  nand_x1_sg U44343 ( .A(n25288), .B(n25289), .X(n39948) );
  nand_x1_sg U44344 ( .A(n25288), .B(n25289), .X(n39949) );
  nand_x1_sg U44345 ( .A(n25288), .B(n25289), .X(n14406) );
  nand_x1_sg U44346 ( .A(n24452), .B(n24453), .X(n39950) );
  nand_x1_sg U44347 ( .A(n24452), .B(n24453), .X(n39951) );
  nand_x1_sg U44348 ( .A(n24452), .B(n24453), .X(n11949) );
  nand_x1_sg U44349 ( .A(n24730), .B(n24731), .X(n39952) );
  nand_x1_sg U44350 ( .A(n24730), .B(n24731), .X(n39953) );
  nand_x1_sg U44351 ( .A(n24730), .B(n24731), .X(n12768) );
  nand_x1_sg U44352 ( .A(n25009), .B(n25010), .X(n39954) );
  nand_x1_sg U44353 ( .A(n25009), .B(n25010), .X(n39955) );
  nand_x1_sg U44354 ( .A(n25009), .B(n25010), .X(n13587) );
  nand_x1_sg U44355 ( .A(n22846), .B(n46844), .X(n39956) );
  nand_x1_sg U44356 ( .A(n22846), .B(n46844), .X(n39957) );
  nand_x1_sg U44357 ( .A(n22846), .B(n46844), .X(n6827) );
  nand_x1_sg U44358 ( .A(n22848), .B(n42046), .X(n22846) );
  nand_x1_sg U44359 ( .A(n23894), .B(n23895), .X(n39958) );
  nand_x1_sg U44360 ( .A(n23894), .B(n23895), .X(n39959) );
  nand_x1_sg U44361 ( .A(n23894), .B(n23895), .X(n10311) );
  nand_x1_sg U44362 ( .A(n24173), .B(n24174), .X(n39960) );
  nand_x1_sg U44363 ( .A(n24173), .B(n24174), .X(n39961) );
  nand_x1_sg U44364 ( .A(n24173), .B(n24174), .X(n11130) );
  inv_x1_sg U44365 ( .A(n41929), .X(n39962) );
  inv_x1_sg U44366 ( .A(n39962), .X(n39963) );
  inv_x1_sg U44367 ( .A(n39962), .X(n39964) );
  inv_x1_sg U44368 ( .A(n39962), .X(n39965) );
  inv_x1_sg U44369 ( .A(n41928), .X(n39966) );
  inv_x1_sg U44370 ( .A(n39966), .X(n39967) );
  inv_x1_sg U44371 ( .A(n39966), .X(n39968) );
  inv_x1_sg U44372 ( .A(n39966), .X(n39969) );
  inv_x1_sg U44373 ( .A(n41927), .X(n39970) );
  inv_x1_sg U44374 ( .A(n39970), .X(n39971) );
  inv_x1_sg U44375 ( .A(n39970), .X(n39972) );
  inv_x1_sg U44376 ( .A(n39970), .X(n39973) );
  inv_x1_sg U44377 ( .A(n41926), .X(n39974) );
  inv_x1_sg U44378 ( .A(n39974), .X(n39975) );
  inv_x1_sg U44379 ( .A(n39974), .X(n39976) );
  inv_x1_sg U44380 ( .A(n39974), .X(n39977) );
  inv_x1_sg U44381 ( .A(n41925), .X(n39978) );
  inv_x1_sg U44382 ( .A(n39978), .X(n39979) );
  inv_x1_sg U44383 ( .A(n39978), .X(n39980) );
  inv_x1_sg U44384 ( .A(n39978), .X(n39981) );
  inv_x1_sg U44385 ( .A(n41924), .X(n39982) );
  inv_x1_sg U44386 ( .A(n39982), .X(n39983) );
  inv_x1_sg U44387 ( .A(n39982), .X(n39984) );
  inv_x1_sg U44388 ( .A(n39982), .X(n39985) );
  inv_x1_sg U44389 ( .A(n41923), .X(n39986) );
  inv_x1_sg U44390 ( .A(n39986), .X(n39987) );
  inv_x1_sg U44391 ( .A(n39986), .X(n39988) );
  inv_x1_sg U44392 ( .A(n39986), .X(n39989) );
  inv_x1_sg U44393 ( .A(n41922), .X(n39990) );
  inv_x1_sg U44394 ( .A(n39990), .X(n39991) );
  inv_x1_sg U44395 ( .A(n39990), .X(n39992) );
  inv_x1_sg U44396 ( .A(n39990), .X(n39993) );
  inv_x1_sg U44397 ( .A(n41921), .X(n39994) );
  inv_x1_sg U44398 ( .A(n39994), .X(n39995) );
  inv_x1_sg U44399 ( .A(n39994), .X(n39996) );
  inv_x1_sg U44400 ( .A(n39994), .X(n39997) );
  inv_x1_sg U44401 ( .A(n41920), .X(n39998) );
  inv_x1_sg U44402 ( .A(n39998), .X(n39999) );
  inv_x1_sg U44403 ( .A(n39998), .X(n40000) );
  inv_x1_sg U44404 ( .A(n39998), .X(n40001) );
  inv_x1_sg U44405 ( .A(n41919), .X(n40002) );
  inv_x1_sg U44406 ( .A(n40002), .X(n40003) );
  inv_x1_sg U44407 ( .A(n40002), .X(n40004) );
  inv_x1_sg U44408 ( .A(n40002), .X(n40005) );
  inv_x1_sg U44409 ( .A(n41910), .X(n40006) );
  inv_x1_sg U44410 ( .A(n40006), .X(n40007) );
  inv_x1_sg U44411 ( .A(n40006), .X(n40008) );
  inv_x1_sg U44412 ( .A(n40006), .X(n40009) );
  inv_x1_sg U44413 ( .A(n39156), .X(n40010) );
  inv_x1_sg U44414 ( .A(n41411), .X(n40011) );
  inv_x1_sg U44415 ( .A(n41406), .X(n40012) );
  inv_x1_sg U44416 ( .A(n38816), .X(n40013) );
  inv_x1_sg U44417 ( .A(n40013), .X(n40014) );
  inv_x1_sg U44418 ( .A(n40013), .X(n40015) );
  inv_x1_sg U44419 ( .A(n40013), .X(n40016) );
  inv_x1_sg U44420 ( .A(n39150), .X(n40017) );
  inv_x1_sg U44421 ( .A(n41401), .X(n40018) );
  inv_x1_sg U44422 ( .A(n39280), .X(n40019) );
  inv_x1_sg U44423 ( .A(n39478), .X(n40020) );
  inv_x1_sg U44424 ( .A(n39281), .X(n40021) );
  inv_x1_sg U44425 ( .A(n39144), .X(n40022) );
  inv_x1_sg U44426 ( .A(n41389), .X(n40023) );
  inv_x1_sg U44427 ( .A(n41393), .X(n40024) );
  inv_x1_sg U44428 ( .A(n40024), .X(n40025) );
  inv_x1_sg U44429 ( .A(n40024), .X(n40026) );
  inv_x1_sg U44430 ( .A(n40024), .X(n40027) );
  inv_x1_sg U44431 ( .A(n39142), .X(n40028) );
  inv_x1_sg U44432 ( .A(n40028), .X(n40029) );
  inv_x1_sg U44433 ( .A(n40028), .X(n40030) );
  inv_x1_sg U44434 ( .A(n40028), .X(n40031) );
  inv_x1_sg U44435 ( .A(n39139), .X(n40032) );
  inv_x1_sg U44436 ( .A(n40032), .X(n40033) );
  inv_x1_sg U44437 ( .A(n40032), .X(n40034) );
  inv_x1_sg U44438 ( .A(n40032), .X(n40035) );
  inv_x1_sg U44439 ( .A(n42370), .X(n40036) );
  inv_x1_sg U44440 ( .A(n40036), .X(n40037) );
  inv_x1_sg U44441 ( .A(n40036), .X(n40038) );
  nand_x1_sg U44442 ( .A(n42326), .B(n22828), .X(n40039) );
  nand_x1_sg U44443 ( .A(n42326), .B(n22828), .X(n40040) );
  nand_x1_sg U44444 ( .A(n42131), .B(n23385), .X(n40041) );
  nand_x1_sg U44445 ( .A(n42131), .B(n23385), .X(n40042) );
  nand_x1_sg U44446 ( .A(n42129), .B(n23664), .X(n40043) );
  nand_x1_sg U44447 ( .A(n42129), .B(n23664), .X(n40044) );
  nand_x1_sg U44448 ( .A(n42128), .B(n23943), .X(n40045) );
  nand_x1_sg U44449 ( .A(n42128), .B(n23943), .X(n40046) );
  nand_x1_sg U44450 ( .A(n42127), .B(n24222), .X(n40047) );
  nand_x1_sg U44451 ( .A(n42127), .B(n24222), .X(n40048) );
  nand_x1_sg U44452 ( .A(n42125), .B(n24501), .X(n40049) );
  nand_x1_sg U44453 ( .A(n42125), .B(n24501), .X(n40050) );
  nand_x1_sg U44454 ( .A(n48856), .B(n24779), .X(n40051) );
  nand_x1_sg U44455 ( .A(n48856), .B(n24779), .X(n40052) );
  nand_x1_sg U44456 ( .A(n49429), .B(n25337), .X(n40053) );
  nand_x1_sg U44457 ( .A(n49429), .B(n25337), .X(n40054) );
  nand_x1_sg U44458 ( .A(n42123), .B(n25616), .X(n40055) );
  nand_x1_sg U44459 ( .A(n42123), .B(n25616), .X(n40056) );
  nand_x1_sg U44460 ( .A(n50001), .B(n25893), .X(n40057) );
  nand_x1_sg U44461 ( .A(n50001), .B(n25893), .X(n40058) );
  nand_x1_sg U44462 ( .A(n42121), .B(n26453), .X(n40059) );
  nand_x1_sg U44463 ( .A(n42121), .B(n26453), .X(n40060) );
  nand_x1_sg U44464 ( .A(n50862), .B(n26731), .X(n40061) );
  nand_x1_sg U44465 ( .A(n50862), .B(n26731), .X(n40062) );
  nand_x1_sg U44466 ( .A(n42090), .B(n23105), .X(n40063) );
  nand_x1_sg U44467 ( .A(n42090), .B(n23105), .X(n40064) );
  nand_x1_sg U44468 ( .A(n49143), .B(n25058), .X(n40065) );
  nand_x1_sg U44469 ( .A(n49143), .B(n25058), .X(n40066) );
  nand_x1_sg U44470 ( .A(n26472), .B(n50564), .X(n40067) );
  nand_x1_sg U44471 ( .A(n26472), .B(n50564), .X(n40068) );
  nand_x1_sg U44472 ( .A(n26123), .B(n41959), .X(n40069) );
  nand_x1_sg U44473 ( .A(n26123), .B(n41959), .X(n40070) );
  inv_x1_sg U44474 ( .A(n50301), .X(n40071) );
  inv_x1_sg U44475 ( .A(n40071), .X(n40072) );
  inv_x1_sg U44476 ( .A(n40071), .X(n40073) );
  inv_x1_sg U44477 ( .A(n40071), .X(n40074) );
  inv_x1_sg U44478 ( .A(n39503), .X(n40075) );
  inv_x1_sg U44479 ( .A(n40075), .X(n40076) );
  inv_x1_sg U44480 ( .A(n40075), .X(n40077) );
  inv_x1_sg U44481 ( .A(n40075), .X(n40078) );
  inv_x1_sg U44482 ( .A(n39501), .X(n40079) );
  inv_x1_sg U44483 ( .A(n40079), .X(n40080) );
  inv_x1_sg U44484 ( .A(n40079), .X(n40081) );
  inv_x1_sg U44485 ( .A(n40079), .X(n40082) );
  inv_x1_sg U44486 ( .A(n41779), .X(n40083) );
  inv_x1_sg U44487 ( .A(n40083), .X(n40084) );
  inv_x1_sg U44488 ( .A(n40083), .X(n40085) );
  inv_x1_sg U44489 ( .A(n41778), .X(n40086) );
  inv_x1_sg U44490 ( .A(n40086), .X(n40087) );
  inv_x1_sg U44491 ( .A(n40086), .X(n40088) );
  inv_x1_sg U44492 ( .A(n38982), .X(n40089) );
  inv_x1_sg U44493 ( .A(n38982), .X(n40090) );
  inv_x1_sg U44494 ( .A(n38985), .X(n40091) );
  inv_x1_sg U44495 ( .A(n40091), .X(n40092) );
  inv_x1_sg U44496 ( .A(n40091), .X(n40093) );
  inv_x1_sg U44497 ( .A(n40091), .X(n40094) );
  inv_x1_sg U44498 ( .A(n39147), .X(n40095) );
  inv_x1_sg U44499 ( .A(n41394), .X(n40096) );
  inv_x1_sg U44500 ( .A(n40096), .X(n40097) );
  inv_x1_sg U44501 ( .A(n40097), .X(n40098) );
  inv_x1_sg U44502 ( .A(n40097), .X(n40099) );
  inv_x1_sg U44503 ( .A(n40097), .X(n40100) );
  inv_x1_sg U44504 ( .A(n23262), .X(n40101) );
  inv_x1_sg U44505 ( .A(n40101), .X(n40102) );
  inv_x1_sg U44506 ( .A(n40101), .X(n40103) );
  inv_x1_sg U44507 ( .A(n40101), .X(n40104) );
  nand_x1_sg U44508 ( .A(n23064), .B(n23065), .X(n40105) );
  nand_x1_sg U44509 ( .A(n23064), .B(n23065), .X(n40106) );
  nand_x1_sg U44510 ( .A(n23344), .B(n23345), .X(n40107) );
  nand_x1_sg U44511 ( .A(n23344), .B(n23345), .X(n40108) );
  nand_x1_sg U44512 ( .A(n23623), .B(n23624), .X(n40109) );
  nand_x1_sg U44513 ( .A(n23623), .B(n23624), .X(n40110) );
  nand_x1_sg U44514 ( .A(n23902), .B(n23903), .X(n40111) );
  nand_x1_sg U44515 ( .A(n23902), .B(n23903), .X(n40112) );
  nand_x1_sg U44516 ( .A(n24181), .B(n24182), .X(n40113) );
  nand_x1_sg U44517 ( .A(n24181), .B(n24182), .X(n40114) );
  nand_x1_sg U44518 ( .A(n24460), .B(n24461), .X(n40115) );
  nand_x1_sg U44519 ( .A(n24460), .B(n24461), .X(n40116) );
  nand_x1_sg U44520 ( .A(n24738), .B(n24739), .X(n40117) );
  nand_x1_sg U44521 ( .A(n24738), .B(n24739), .X(n40118) );
  nand_x1_sg U44522 ( .A(n25017), .B(n25018), .X(n40119) );
  nand_x1_sg U44523 ( .A(n25017), .B(n25018), .X(n40120) );
  nand_x1_sg U44524 ( .A(n25296), .B(n25297), .X(n40121) );
  nand_x1_sg U44525 ( .A(n25296), .B(n25297), .X(n40122) );
  nand_x1_sg U44526 ( .A(n25575), .B(n25576), .X(n40123) );
  nand_x1_sg U44527 ( .A(n25575), .B(n25576), .X(n40124) );
  nand_x1_sg U44528 ( .A(n25852), .B(n25853), .X(n40125) );
  nand_x1_sg U44529 ( .A(n25852), .B(n25853), .X(n40126) );
  nand_x1_sg U44530 ( .A(n26690), .B(n26691), .X(n40127) );
  nand_x1_sg U44531 ( .A(n26690), .B(n26691), .X(n40128) );
  nand_x1_sg U44532 ( .A(n26081), .B(n26082), .X(n40129) );
  nand_x1_sg U44533 ( .A(n26081), .B(n26082), .X(n40130) );
  nand_x1_sg U44534 ( .A(n26412), .B(n26413), .X(n40131) );
  nand_x1_sg U44535 ( .A(n26412), .B(n26413), .X(n40132) );
  nand_x1_sg U44536 ( .A(n42186), .B(n23071), .X(n40133) );
  nand_x1_sg U44537 ( .A(n42186), .B(n23071), .X(n40134) );
  nand_x1_sg U44538 ( .A(n42184), .B(n23351), .X(n40135) );
  nand_x1_sg U44539 ( .A(n42184), .B(n23351), .X(n40136) );
  nand_x1_sg U44540 ( .A(n42182), .B(n23630), .X(n40137) );
  nand_x1_sg U44541 ( .A(n42182), .B(n23630), .X(n40138) );
  nand_x1_sg U44542 ( .A(n42180), .B(n23909), .X(n40139) );
  nand_x1_sg U44543 ( .A(n42180), .B(n23909), .X(n40140) );
  nand_x1_sg U44544 ( .A(n42178), .B(n24188), .X(n40141) );
  nand_x1_sg U44545 ( .A(n42178), .B(n24188), .X(n40142) );
  nand_x1_sg U44546 ( .A(n42176), .B(n24467), .X(n40143) );
  nand_x1_sg U44547 ( .A(n42176), .B(n24467), .X(n40144) );
  nand_x1_sg U44548 ( .A(n42174), .B(n24745), .X(n40145) );
  nand_x1_sg U44549 ( .A(n42174), .B(n24745), .X(n40146) );
  nand_x1_sg U44550 ( .A(n42172), .B(n25024), .X(n40147) );
  nand_x1_sg U44551 ( .A(n42172), .B(n25024), .X(n40148) );
  nand_x1_sg U44552 ( .A(n42170), .B(n25303), .X(n40149) );
  nand_x1_sg U44553 ( .A(n42170), .B(n25303), .X(n40150) );
  nand_x1_sg U44554 ( .A(n49754), .B(n25582), .X(n40151) );
  nand_x1_sg U44555 ( .A(n49754), .B(n25582), .X(n40152) );
  nand_x1_sg U44556 ( .A(n42167), .B(n25859), .X(n40153) );
  nand_x1_sg U44557 ( .A(n42167), .B(n25859), .X(n40154) );
  nand_x1_sg U44558 ( .A(n42165), .B(n26697), .X(n40155) );
  nand_x1_sg U44559 ( .A(n42165), .B(n26697), .X(n40156) );
  nand_x1_sg U44560 ( .A(n41986), .B(n26419), .X(n40159) );
  nand_x1_sg U44561 ( .A(n41986), .B(n26419), .X(n40160) );
  inv_x1_sg U44562 ( .A(n41808), .X(n40161) );
  inv_x1_sg U44563 ( .A(n40161), .X(n40162) );
  inv_x1_sg U44564 ( .A(n40161), .X(n40163) );
  inv_x1_sg U44565 ( .A(n40161), .X(n40164) );
  inv_x1_sg U44566 ( .A(n41753), .X(n40165) );
  inv_x1_sg U44567 ( .A(n40165), .X(n40166) );
  inv_x1_sg U44568 ( .A(n40165), .X(n40167) );
  inv_x1_sg U44569 ( .A(n40165), .X(n40168) );
  inv_x1_sg U44570 ( .A(n41752), .X(n40169) );
  inv_x1_sg U44571 ( .A(n40169), .X(n40170) );
  inv_x1_sg U44572 ( .A(n40169), .X(n40171) );
  inv_x1_sg U44573 ( .A(n40169), .X(n40172) );
  inv_x1_sg U44574 ( .A(n41751), .X(n40173) );
  inv_x1_sg U44575 ( .A(n40173), .X(n40174) );
  inv_x1_sg U44576 ( .A(n40173), .X(n40175) );
  inv_x1_sg U44577 ( .A(n40173), .X(n40176) );
  inv_x1_sg U44578 ( .A(n41750), .X(n40177) );
  inv_x1_sg U44579 ( .A(n40177), .X(n40178) );
  inv_x1_sg U44580 ( .A(n40177), .X(n40179) );
  inv_x1_sg U44581 ( .A(n40177), .X(n40180) );
  inv_x1_sg U44582 ( .A(n41749), .X(n40181) );
  inv_x1_sg U44583 ( .A(n40181), .X(n40182) );
  inv_x1_sg U44584 ( .A(n40181), .X(n40183) );
  inv_x1_sg U44585 ( .A(n40181), .X(n40184) );
  inv_x1_sg U44586 ( .A(n41748), .X(n40185) );
  inv_x1_sg U44587 ( .A(n40185), .X(n40186) );
  inv_x1_sg U44588 ( .A(n40185), .X(n40187) );
  inv_x1_sg U44589 ( .A(n40185), .X(n40188) );
  inv_x1_sg U44590 ( .A(n41747), .X(n40189) );
  inv_x1_sg U44591 ( .A(n40189), .X(n40190) );
  inv_x1_sg U44592 ( .A(n40189), .X(n40191) );
  inv_x1_sg U44593 ( .A(n40189), .X(n40192) );
  inv_x1_sg U44594 ( .A(n41746), .X(n40193) );
  inv_x1_sg U44595 ( .A(n40193), .X(n40194) );
  inv_x1_sg U44596 ( .A(n40193), .X(n40195) );
  inv_x1_sg U44597 ( .A(n40193), .X(n40196) );
  inv_x1_sg U44598 ( .A(n41745), .X(n40197) );
  inv_x1_sg U44599 ( .A(n40197), .X(n40198) );
  inv_x1_sg U44600 ( .A(n40197), .X(n40199) );
  inv_x1_sg U44601 ( .A(n40197), .X(n40200) );
  inv_x1_sg U44602 ( .A(n41744), .X(n40201) );
  inv_x1_sg U44603 ( .A(n40201), .X(n40202) );
  inv_x1_sg U44604 ( .A(n40201), .X(n40203) );
  inv_x1_sg U44605 ( .A(n40201), .X(n40204) );
  inv_x1_sg U44606 ( .A(n41743), .X(n40205) );
  inv_x1_sg U44607 ( .A(n40205), .X(n40206) );
  inv_x1_sg U44608 ( .A(n40205), .X(n40207) );
  inv_x1_sg U44609 ( .A(n40205), .X(n40208) );
  inv_x1_sg U44610 ( .A(n41742), .X(n40209) );
  inv_x1_sg U44611 ( .A(n40209), .X(n40210) );
  inv_x1_sg U44612 ( .A(n40209), .X(n40211) );
  inv_x1_sg U44613 ( .A(n40209), .X(n40212) );
  inv_x1_sg U44614 ( .A(n41741), .X(n40213) );
  inv_x1_sg U44615 ( .A(n40213), .X(n40214) );
  inv_x1_sg U44616 ( .A(n40213), .X(n40215) );
  inv_x1_sg U44617 ( .A(n40213), .X(n40216) );
  inv_x1_sg U44618 ( .A(n39199), .X(n40217) );
  inv_x1_sg U44619 ( .A(n39655), .X(n40218) );
  inv_x1_sg U44620 ( .A(n41420), .X(n40219) );
  inv_x1_sg U44621 ( .A(n40219), .X(n40220) );
  inv_x1_sg U44622 ( .A(n40219), .X(n40221) );
  inv_x1_sg U44623 ( .A(n40219), .X(n40222) );
  inv_x1_sg U44624 ( .A(n41463), .X(n40223) );
  inv_x1_sg U44625 ( .A(n40223), .X(n40224) );
  inv_x1_sg U44626 ( .A(n40223), .X(n40225) );
  inv_x1_sg U44627 ( .A(n40223), .X(n40226) );
  inv_x1_sg U44628 ( .A(n40223), .X(n40227) );
  inv_x1_sg U44629 ( .A(n16936), .X(n40228) );
  inv_x1_sg U44630 ( .A(n40228), .X(n40229) );
  inv_x1_sg U44631 ( .A(n40228), .X(n40230) );
  inv_x1_sg U44632 ( .A(n40228), .X(n40231) );
  inv_x1_sg U44633 ( .A(n7111), .X(n40232) );
  inv_x1_sg U44634 ( .A(n40232), .X(n40233) );
  inv_x1_sg U44635 ( .A(n40232), .X(n40234) );
  inv_x1_sg U44636 ( .A(n40232), .X(n40235) );
  inv_x1_sg U44637 ( .A(n40514), .X(n40236) );
  inv_x1_sg U44638 ( .A(n40236), .X(n40237) );
  inv_x1_sg U44639 ( .A(n40236), .X(n40238) );
  inv_x1_sg U44640 ( .A(n40236), .X(n40239) );
  inv_x1_sg U44641 ( .A(n40236), .X(n40240) );
  inv_x1_sg U44642 ( .A(n40558), .X(n40241) );
  inv_x1_sg U44643 ( .A(n40241), .X(n40242) );
  inv_x1_sg U44644 ( .A(n40241), .X(n40243) );
  inv_x1_sg U44645 ( .A(n40241), .X(n40244) );
  inv_x1_sg U44646 ( .A(n40241), .X(n40245) );
  inv_x1_sg U44647 ( .A(n40554), .X(n40246) );
  inv_x1_sg U44648 ( .A(n40246), .X(n40247) );
  inv_x1_sg U44649 ( .A(n40246), .X(n40248) );
  inv_x1_sg U44650 ( .A(n40246), .X(n40249) );
  inv_x1_sg U44651 ( .A(n40246), .X(n40250) );
  inv_x1_sg U44652 ( .A(n40550), .X(n40251) );
  inv_x1_sg U44653 ( .A(n40251), .X(n40252) );
  inv_x1_sg U44654 ( .A(n40251), .X(n40253) );
  inv_x1_sg U44655 ( .A(n40251), .X(n40254) );
  inv_x1_sg U44656 ( .A(n40251), .X(n40255) );
  inv_x1_sg U44657 ( .A(n40546), .X(n40256) );
  inv_x1_sg U44658 ( .A(n40256), .X(n40257) );
  inv_x1_sg U44659 ( .A(n40256), .X(n40258) );
  inv_x1_sg U44660 ( .A(n40256), .X(n40259) );
  inv_x1_sg U44661 ( .A(n40256), .X(n40260) );
  inv_x1_sg U44662 ( .A(n40542), .X(n40261) );
  inv_x1_sg U44663 ( .A(n40261), .X(n40262) );
  inv_x1_sg U44664 ( .A(n40261), .X(n40263) );
  inv_x1_sg U44665 ( .A(n40261), .X(n40264) );
  inv_x1_sg U44666 ( .A(n40261), .X(n40265) );
  inv_x1_sg U44667 ( .A(n40538), .X(n40266) );
  inv_x1_sg U44668 ( .A(n40266), .X(n40267) );
  inv_x1_sg U44669 ( .A(n40266), .X(n40268) );
  inv_x1_sg U44670 ( .A(n40266), .X(n40269) );
  inv_x1_sg U44671 ( .A(n40266), .X(n40270) );
  inv_x1_sg U44672 ( .A(n40534), .X(n40271) );
  inv_x1_sg U44673 ( .A(n40271), .X(n40272) );
  inv_x1_sg U44674 ( .A(n40271), .X(n40273) );
  inv_x1_sg U44675 ( .A(n40271), .X(n40274) );
  inv_x1_sg U44676 ( .A(n40271), .X(n40275) );
  inv_x1_sg U44677 ( .A(n40530), .X(n40276) );
  inv_x1_sg U44678 ( .A(n40276), .X(n40277) );
  inv_x1_sg U44679 ( .A(n40276), .X(n40278) );
  inv_x1_sg U44680 ( .A(n40276), .X(n40279) );
  inv_x1_sg U44681 ( .A(n40276), .X(n40280) );
  inv_x1_sg U44682 ( .A(n40526), .X(n40281) );
  inv_x1_sg U44683 ( .A(n40281), .X(n40282) );
  inv_x1_sg U44684 ( .A(n40281), .X(n40283) );
  inv_x1_sg U44685 ( .A(n40281), .X(n40284) );
  inv_x1_sg U44686 ( .A(n40281), .X(n40285) );
  inv_x1_sg U44687 ( .A(n40522), .X(n40286) );
  inv_x1_sg U44688 ( .A(n40286), .X(n40287) );
  inv_x1_sg U44689 ( .A(n40286), .X(n40288) );
  inv_x1_sg U44690 ( .A(n40286), .X(n40289) );
  inv_x1_sg U44691 ( .A(n40286), .X(n40290) );
  inv_x1_sg U44692 ( .A(n40518), .X(n40291) );
  inv_x1_sg U44693 ( .A(n40291), .X(n40292) );
  inv_x1_sg U44694 ( .A(n40291), .X(n40293) );
  inv_x1_sg U44695 ( .A(n40291), .X(n40294) );
  inv_x1_sg U44696 ( .A(n40291), .X(n40295) );
  inv_x1_sg U44697 ( .A(n40510), .X(n40296) );
  inv_x1_sg U44698 ( .A(n40296), .X(n40297) );
  inv_x1_sg U44699 ( .A(n40296), .X(n40298) );
  inv_x1_sg U44700 ( .A(n40296), .X(n40299) );
  inv_x1_sg U44701 ( .A(n40296), .X(n40300) );
  inv_x1_sg U44702 ( .A(n16658), .X(n40301) );
  inv_x1_sg U44703 ( .A(n40566), .X(n40302) );
  inv_x1_sg U44704 ( .A(n40565), .X(n40303) );
  inv_x1_sg U44705 ( .A(n16658), .X(n40304) );
  inv_x1_sg U44706 ( .A(n41847), .X(n40305) );
  inv_x1_sg U44707 ( .A(n40305), .X(n40306) );
  inv_x1_sg U44708 ( .A(n40305), .X(n40307) );
  inv_x1_sg U44709 ( .A(n40305), .X(n40308) );
  inv_x1_sg U44710 ( .A(n41842), .X(n40309) );
  inv_x1_sg U44711 ( .A(n40309), .X(n40310) );
  inv_x1_sg U44712 ( .A(n40309), .X(n40311) );
  inv_x1_sg U44713 ( .A(n40309), .X(n40312) );
  inv_x1_sg U44714 ( .A(n6831), .X(n40313) );
  inv_x1_sg U44715 ( .A(n40313), .X(n40314) );
  inv_x1_sg U44716 ( .A(n40313), .X(n40315) );
  inv_x1_sg U44717 ( .A(n40313), .X(n40316) );
  inv_x1_sg U44718 ( .A(n42095), .X(n40317) );
  inv_x1_sg U44719 ( .A(n40317), .X(n40318) );
  inv_x1_sg U44720 ( .A(n40317), .X(n40319) );
  inv_x1_sg U44721 ( .A(n40317), .X(n40320) );
  inv_x1_sg U44722 ( .A(n42094), .X(n40321) );
  inv_x1_sg U44723 ( .A(n40321), .X(n40322) );
  inv_x1_sg U44724 ( .A(n40321), .X(n40323) );
  inv_x1_sg U44725 ( .A(n40321), .X(n40324) );
  inv_x1_sg U44726 ( .A(n42100), .X(n40325) );
  inv_x1_sg U44727 ( .A(n40325), .X(n40326) );
  inv_x1_sg U44728 ( .A(n40325), .X(n40327) );
  inv_x1_sg U44729 ( .A(n40325), .X(n40328) );
  inv_x1_sg U44730 ( .A(n42093), .X(n40329) );
  inv_x1_sg U44731 ( .A(n40329), .X(n40330) );
  inv_x1_sg U44732 ( .A(n40329), .X(n40331) );
  inv_x1_sg U44733 ( .A(n40329), .X(n40332) );
  inv_x1_sg U44734 ( .A(n42098), .X(n40333) );
  inv_x1_sg U44735 ( .A(n40333), .X(n40334) );
  inv_x1_sg U44736 ( .A(n40333), .X(n40335) );
  inv_x1_sg U44737 ( .A(n40333), .X(n40336) );
  inv_x1_sg U44738 ( .A(n42099), .X(n40337) );
  inv_x1_sg U44739 ( .A(n40337), .X(n40338) );
  inv_x1_sg U44740 ( .A(n40337), .X(n40339) );
  inv_x1_sg U44741 ( .A(n40337), .X(n40340) );
  inv_x1_sg U44742 ( .A(n42097), .X(n40341) );
  inv_x1_sg U44743 ( .A(n40341), .X(n40342) );
  inv_x1_sg U44744 ( .A(n40341), .X(n40343) );
  inv_x1_sg U44745 ( .A(n40341), .X(n40344) );
  inv_x1_sg U44746 ( .A(n42101), .X(n40345) );
  inv_x1_sg U44747 ( .A(n40345), .X(n40346) );
  inv_x1_sg U44748 ( .A(n40345), .X(n40347) );
  inv_x1_sg U44749 ( .A(n40345), .X(n40348) );
  inv_x1_sg U44750 ( .A(n42102), .X(n40349) );
  inv_x1_sg U44751 ( .A(n40349), .X(n40350) );
  inv_x1_sg U44752 ( .A(n40349), .X(n40351) );
  inv_x1_sg U44753 ( .A(n40349), .X(n40352) );
  inv_x1_sg U44754 ( .A(n42103), .X(n40353) );
  inv_x1_sg U44755 ( .A(n40353), .X(n40354) );
  inv_x1_sg U44756 ( .A(n40353), .X(n40355) );
  inv_x1_sg U44757 ( .A(n40353), .X(n40356) );
  inv_x1_sg U44758 ( .A(n42104), .X(n40357) );
  inv_x1_sg U44759 ( .A(n40357), .X(n40358) );
  inv_x1_sg U44760 ( .A(n40357), .X(n40359) );
  inv_x1_sg U44761 ( .A(n40357), .X(n40360) );
  inv_x1_sg U44762 ( .A(n40357), .X(n40361) );
  inv_x1_sg U44763 ( .A(n50565), .X(n40362) );
  inv_x1_sg U44764 ( .A(n40362), .X(n40363) );
  inv_x1_sg U44765 ( .A(n40362), .X(n40364) );
  inv_x1_sg U44766 ( .A(n40362), .X(n40365) );
  inv_x1_sg U44767 ( .A(n41903), .X(n40366) );
  inv_x1_sg U44768 ( .A(n40366), .X(n40367) );
  inv_x1_sg U44769 ( .A(n40366), .X(n40368) );
  inv_x1_sg U44770 ( .A(n40366), .X(n40369) );
  inv_x1_sg U44771 ( .A(n39200), .X(n40370) );
  inv_x1_sg U44772 ( .A(n39651), .X(n40371) );
  inv_x1_sg U44773 ( .A(n39436), .X(n40372) );
  inv_x1_sg U44774 ( .A(n40372), .X(n40373) );
  inv_x1_sg U44775 ( .A(n40372), .X(n40374) );
  inv_x1_sg U44776 ( .A(n40372), .X(n40375) );
  inv_x1_sg U44777 ( .A(n40372), .X(n40376) );
  inv_x1_sg U44778 ( .A(n39195), .X(n40377) );
  inv_x1_sg U44779 ( .A(n39196), .X(n40378) );
  inv_x1_sg U44780 ( .A(n41457), .X(n40379) );
  inv_x1_sg U44781 ( .A(n40379), .X(n40380) );
  inv_x1_sg U44782 ( .A(n40379), .X(n40381) );
  inv_x1_sg U44783 ( .A(n40379), .X(n40382) );
  inv_x1_sg U44784 ( .A(n40379), .X(n40383) );
  inv_x1_sg U44785 ( .A(n39191), .X(n40384) );
  inv_x1_sg U44786 ( .A(n39190), .X(n40385) );
  inv_x1_sg U44787 ( .A(n41452), .X(n40386) );
  inv_x1_sg U44788 ( .A(n40386), .X(n40387) );
  inv_x1_sg U44789 ( .A(n40386), .X(n40388) );
  inv_x1_sg U44790 ( .A(n40386), .X(n40389) );
  inv_x1_sg U44791 ( .A(n40386), .X(n40390) );
  inv_x1_sg U44792 ( .A(n39185), .X(n40391) );
  inv_x1_sg U44793 ( .A(n39185), .X(n40392) );
  inv_x1_sg U44794 ( .A(n41448), .X(n40393) );
  inv_x1_sg U44795 ( .A(n40393), .X(n40394) );
  inv_x1_sg U44796 ( .A(n40393), .X(n40395) );
  inv_x1_sg U44797 ( .A(n40393), .X(n40396) );
  inv_x1_sg U44798 ( .A(n40393), .X(n40397) );
  inv_x1_sg U44799 ( .A(n39181), .X(n40398) );
  inv_x1_sg U44800 ( .A(n39180), .X(n40399) );
  inv_x1_sg U44801 ( .A(n41443), .X(n40400) );
  inv_x1_sg U44802 ( .A(n40400), .X(n40401) );
  inv_x1_sg U44803 ( .A(n40400), .X(n40402) );
  inv_x1_sg U44804 ( .A(n40400), .X(n40403) );
  inv_x1_sg U44805 ( .A(n40400), .X(n40404) );
  inv_x1_sg U44806 ( .A(n39176), .X(n40405) );
  inv_x1_sg U44807 ( .A(n39175), .X(n40406) );
  inv_x1_sg U44808 ( .A(n41439), .X(n40407) );
  inv_x1_sg U44809 ( .A(n40407), .X(n40408) );
  inv_x1_sg U44810 ( .A(n40407), .X(n40409) );
  inv_x1_sg U44811 ( .A(n40407), .X(n40410) );
  inv_x1_sg U44812 ( .A(n40407), .X(n40411) );
  inv_x1_sg U44813 ( .A(n41438), .X(n40412) );
  inv_x1_sg U44814 ( .A(n40412), .X(n40413) );
  inv_x1_sg U44815 ( .A(n40412), .X(n40414) );
  inv_x1_sg U44816 ( .A(n40412), .X(n40415) );
  inv_x1_sg U44817 ( .A(n40412), .X(n40416) );
  inv_x1_sg U44818 ( .A(n39170), .X(n40417) );
  inv_x1_sg U44819 ( .A(n39170), .X(n40418) );
  inv_x1_sg U44820 ( .A(n41434), .X(n40419) );
  inv_x1_sg U44821 ( .A(n40419), .X(n40420) );
  inv_x1_sg U44822 ( .A(n40419), .X(n40421) );
  inv_x1_sg U44823 ( .A(n40419), .X(n40422) );
  inv_x1_sg U44824 ( .A(n40419), .X(n40423) );
  inv_x1_sg U44825 ( .A(n41433), .X(n40424) );
  inv_x1_sg U44826 ( .A(n40424), .X(n40425) );
  inv_x1_sg U44827 ( .A(n40424), .X(n40426) );
  inv_x1_sg U44828 ( .A(n40424), .X(n40427) );
  inv_x1_sg U44829 ( .A(n40424), .X(n40428) );
  inv_x1_sg U44830 ( .A(n39165), .X(n40429) );
  inv_x1_sg U44831 ( .A(n39165), .X(n40430) );
  inv_x1_sg U44832 ( .A(n41429), .X(n40431) );
  inv_x1_sg U44833 ( .A(n40431), .X(n40432) );
  inv_x1_sg U44834 ( .A(n40431), .X(n40433) );
  inv_x1_sg U44835 ( .A(n40431), .X(n40434) );
  inv_x1_sg U44836 ( .A(n40431), .X(n40435) );
  inv_x1_sg U44837 ( .A(n41428), .X(n40436) );
  inv_x1_sg U44838 ( .A(n40436), .X(n40437) );
  inv_x1_sg U44839 ( .A(n40436), .X(n40438) );
  inv_x1_sg U44840 ( .A(n40436), .X(n40439) );
  inv_x1_sg U44841 ( .A(n40436), .X(n40440) );
  inv_x1_sg U44842 ( .A(n39161), .X(n40441) );
  inv_x1_sg U44843 ( .A(n39160), .X(n40442) );
  inv_x1_sg U44844 ( .A(n41424), .X(n40443) );
  inv_x1_sg U44845 ( .A(n40443), .X(n40444) );
  inv_x1_sg U44846 ( .A(n40443), .X(n40445) );
  inv_x1_sg U44847 ( .A(n40443), .X(n40446) );
  inv_x1_sg U44848 ( .A(n40443), .X(n40447) );
  inv_x1_sg U44849 ( .A(n41425), .X(n40448) );
  inv_x1_sg U44850 ( .A(n40448), .X(n40449) );
  inv_x1_sg U44851 ( .A(n40448), .X(n40450) );
  inv_x1_sg U44852 ( .A(n40448), .X(n40451) );
  inv_x1_sg U44853 ( .A(n40448), .X(n40452) );
  inv_x1_sg U44854 ( .A(n39283), .X(n40453) );
  inv_x1_sg U44855 ( .A(n40453), .X(n40454) );
  inv_x1_sg U44856 ( .A(n40453), .X(n40455) );
  inv_x1_sg U44857 ( .A(n40453), .X(n40456) );
  inv_x1_sg U44858 ( .A(n40453), .X(n40457) );
  inv_x1_sg U44859 ( .A(n26485), .X(n40458) );
  inv_x1_sg U44860 ( .A(n40458), .X(n40459) );
  inv_x1_sg U44861 ( .A(n40458), .X(n40460) );
  inv_x1_sg U44862 ( .A(n40458), .X(n40461) );
  inv_x1_sg U44863 ( .A(n26189), .X(n40462) );
  inv_x1_sg U44864 ( .A(n40462), .X(n40463) );
  inv_x1_sg U44865 ( .A(n40462), .X(n40464) );
  inv_x1_sg U44866 ( .A(n40462), .X(n40465) );
  inv_x1_sg U44867 ( .A(n25648), .X(n40466) );
  inv_x1_sg U44868 ( .A(n40466), .X(n40467) );
  inv_x1_sg U44869 ( .A(n40466), .X(n40468) );
  inv_x1_sg U44870 ( .A(n40466), .X(n40469) );
  inv_x1_sg U44871 ( .A(n25369), .X(n40470) );
  inv_x1_sg U44872 ( .A(n40470), .X(n40471) );
  inv_x1_sg U44873 ( .A(n40470), .X(n40472) );
  inv_x1_sg U44874 ( .A(n40470), .X(n40473) );
  inv_x1_sg U44875 ( .A(n25090), .X(n40474) );
  inv_x1_sg U44876 ( .A(n40474), .X(n40475) );
  inv_x1_sg U44877 ( .A(n40474), .X(n40476) );
  inv_x1_sg U44878 ( .A(n40474), .X(n40477) );
  inv_x1_sg U44879 ( .A(n24811), .X(n40478) );
  inv_x1_sg U44880 ( .A(n40478), .X(n40479) );
  inv_x1_sg U44881 ( .A(n40478), .X(n40480) );
  inv_x1_sg U44882 ( .A(n40478), .X(n40481) );
  inv_x1_sg U44883 ( .A(n24533), .X(n40482) );
  inv_x1_sg U44884 ( .A(n40482), .X(n40483) );
  inv_x1_sg U44885 ( .A(n40482), .X(n40484) );
  inv_x1_sg U44886 ( .A(n40482), .X(n40485) );
  inv_x1_sg U44887 ( .A(n24254), .X(n40486) );
  inv_x1_sg U44888 ( .A(n40486), .X(n40487) );
  inv_x1_sg U44889 ( .A(n40486), .X(n40488) );
  inv_x1_sg U44890 ( .A(n40486), .X(n40489) );
  inv_x1_sg U44891 ( .A(n23975), .X(n40490) );
  inv_x1_sg U44892 ( .A(n40490), .X(n40491) );
  inv_x1_sg U44893 ( .A(n40490), .X(n40492) );
  inv_x1_sg U44894 ( .A(n40490), .X(n40493) );
  inv_x1_sg U44895 ( .A(n23696), .X(n40494) );
  inv_x1_sg U44896 ( .A(n40494), .X(n40495) );
  inv_x1_sg U44897 ( .A(n40494), .X(n40496) );
  inv_x1_sg U44898 ( .A(n40494), .X(n40497) );
  inv_x1_sg U44899 ( .A(n23417), .X(n40498) );
  inv_x1_sg U44900 ( .A(n40498), .X(n40499) );
  inv_x1_sg U44901 ( .A(n40498), .X(n40500) );
  inv_x1_sg U44902 ( .A(n40498), .X(n40501) );
  inv_x1_sg U44903 ( .A(n23137), .X(n40502) );
  inv_x1_sg U44904 ( .A(n40502), .X(n40503) );
  inv_x1_sg U44905 ( .A(n40502), .X(n40504) );
  inv_x1_sg U44906 ( .A(n40502), .X(n40505) );
  inv_x1_sg U44907 ( .A(n22860), .X(n40506) );
  inv_x1_sg U44908 ( .A(n40506), .X(n40507) );
  inv_x1_sg U44909 ( .A(n40506), .X(n40508) );
  inv_x1_sg U44910 ( .A(n40506), .X(n40509) );
  inv_x1_sg U44911 ( .A(n18300), .X(n40510) );
  inv_x1_sg U44912 ( .A(n40510), .X(n40511) );
  inv_x1_sg U44913 ( .A(n40510), .X(n40512) );
  inv_x1_sg U44914 ( .A(n40510), .X(n40513) );
  inv_x1_sg U44915 ( .A(n17479), .X(n40514) );
  inv_x1_sg U44916 ( .A(n40514), .X(n40515) );
  inv_x1_sg U44917 ( .A(n40514), .X(n40516) );
  inv_x1_sg U44918 ( .A(n40514), .X(n40517) );
  inv_x1_sg U44919 ( .A(n15841), .X(n40518) );
  inv_x1_sg U44920 ( .A(n40518), .X(n40519) );
  inv_x1_sg U44921 ( .A(n40518), .X(n40520) );
  inv_x1_sg U44922 ( .A(n40518), .X(n40521) );
  inv_x1_sg U44923 ( .A(n15022), .X(n40522) );
  inv_x1_sg U44924 ( .A(n40522), .X(n40523) );
  inv_x1_sg U44925 ( .A(n40522), .X(n40524) );
  inv_x1_sg U44926 ( .A(n40522), .X(n40525) );
  inv_x1_sg U44927 ( .A(n14203), .X(n40526) );
  inv_x1_sg U44928 ( .A(n40526), .X(n40527) );
  inv_x1_sg U44929 ( .A(n40526), .X(n40528) );
  inv_x1_sg U44930 ( .A(n40526), .X(n40529) );
  inv_x1_sg U44931 ( .A(n13384), .X(n40530) );
  inv_x1_sg U44932 ( .A(n40530), .X(n40531) );
  inv_x1_sg U44933 ( .A(n40530), .X(n40532) );
  inv_x1_sg U44934 ( .A(n40530), .X(n40533) );
  inv_x1_sg U44935 ( .A(n12565), .X(n40534) );
  inv_x1_sg U44936 ( .A(n40534), .X(n40535) );
  inv_x1_sg U44937 ( .A(n40534), .X(n40536) );
  inv_x1_sg U44938 ( .A(n40534), .X(n40537) );
  inv_x1_sg U44939 ( .A(n11746), .X(n40538) );
  inv_x1_sg U44940 ( .A(n40538), .X(n40539) );
  inv_x1_sg U44941 ( .A(n40538), .X(n40540) );
  inv_x1_sg U44942 ( .A(n40538), .X(n40541) );
  inv_x1_sg U44943 ( .A(n10927), .X(n40542) );
  inv_x1_sg U44944 ( .A(n40542), .X(n40543) );
  inv_x1_sg U44945 ( .A(n40542), .X(n40544) );
  inv_x1_sg U44946 ( .A(n40542), .X(n40545) );
  inv_x1_sg U44947 ( .A(n10108), .X(n40546) );
  inv_x1_sg U44948 ( .A(n40546), .X(n40547) );
  inv_x1_sg U44949 ( .A(n40546), .X(n40548) );
  inv_x1_sg U44950 ( .A(n40546), .X(n40549) );
  inv_x1_sg U44951 ( .A(n9289), .X(n40550) );
  inv_x1_sg U44952 ( .A(n40550), .X(n40551) );
  inv_x1_sg U44953 ( .A(n40550), .X(n40552) );
  inv_x1_sg U44954 ( .A(n40550), .X(n40553) );
  inv_x1_sg U44955 ( .A(n8469), .X(n40554) );
  inv_x1_sg U44956 ( .A(n40554), .X(n40555) );
  inv_x1_sg U44957 ( .A(n40554), .X(n40556) );
  inv_x1_sg U44958 ( .A(n40554), .X(n40557) );
  inv_x1_sg U44959 ( .A(n7651), .X(n40558) );
  inv_x1_sg U44960 ( .A(n40558), .X(n40559) );
  inv_x1_sg U44961 ( .A(n40558), .X(n40560) );
  inv_x1_sg U44962 ( .A(n40558), .X(n40561) );
  inv_x1_sg U44963 ( .A(n16658), .X(n40562) );
  inv_x1_sg U44964 ( .A(n40562), .X(n40563) );
  inv_x1_sg U44965 ( .A(n40562), .X(n40564) );
  inv_x1_sg U44966 ( .A(n40562), .X(n40565) );
  inv_x1_sg U44967 ( .A(n40562), .X(n40566) );
  inv_x1_sg U44968 ( .A(n16655), .X(n40567) );
  inv_x1_sg U44969 ( .A(n40567), .X(n40568) );
  inv_x1_sg U44970 ( .A(n40567), .X(n40569) );
  inv_x1_sg U44971 ( .A(n40567), .X(n40570) );
  inv_x1_sg U44972 ( .A(n40567), .X(n40571) );
  inv_x1_sg U44973 ( .A(n6994), .X(n40572) );
  inv_x1_sg U44974 ( .A(n40572), .X(n40573) );
  inv_x1_sg U44975 ( .A(n40572), .X(n40574) );
  inv_x1_sg U44976 ( .A(n40572), .X(n40575) );
  inv_x1_sg U44977 ( .A(n40572), .X(n40576) );
  inv_x1_sg U44978 ( .A(n16818), .X(n40577) );
  inv_x1_sg U44979 ( .A(n40577), .X(n40578) );
  inv_x1_sg U44980 ( .A(n40577), .X(n40579) );
  inv_x1_sg U44981 ( .A(n40577), .X(n40580) );
  inv_x1_sg U44982 ( .A(n40577), .X(n40581) );
  inv_x1_sg U44983 ( .A(n40219), .X(n40582) );
  inv_x1_sg U44984 ( .A(n40582), .X(n40583) );
  inv_x1_sg U44985 ( .A(n40582), .X(n40584) );
  inv_x1_sg U44986 ( .A(n40582), .X(n40585) );
  inv_x1_sg U44987 ( .A(n40582), .X(n40586) );
  inv_x1_sg U44988 ( .A(n41456), .X(n40587) );
  inv_x1_sg U44989 ( .A(n40587), .X(n40588) );
  inv_x1_sg U44990 ( .A(n40587), .X(n40589) );
  inv_x1_sg U44991 ( .A(n40587), .X(n40590) );
  inv_x1_sg U44992 ( .A(n40587), .X(n40591) );
  inv_x1_sg U44993 ( .A(n41451), .X(n40592) );
  inv_x1_sg U44994 ( .A(n40592), .X(n40593) );
  inv_x1_sg U44995 ( .A(n40592), .X(n40594) );
  inv_x1_sg U44996 ( .A(n40592), .X(n40595) );
  inv_x1_sg U44997 ( .A(n40592), .X(n40596) );
  inv_x1_sg U44998 ( .A(n41447), .X(n40597) );
  inv_x1_sg U44999 ( .A(n40597), .X(n40598) );
  inv_x1_sg U45000 ( .A(n40597), .X(n40599) );
  inv_x1_sg U45001 ( .A(n40597), .X(n40600) );
  inv_x1_sg U45002 ( .A(n40597), .X(n40601) );
  inv_x1_sg U45003 ( .A(n41442), .X(n40602) );
  inv_x1_sg U45004 ( .A(n40602), .X(n40603) );
  inv_x1_sg U45005 ( .A(n40602), .X(n40604) );
  inv_x1_sg U45006 ( .A(n40602), .X(n40605) );
  inv_x1_sg U45007 ( .A(n40602), .X(n40606) );
  inv_x1_sg U45008 ( .A(n16850), .X(n40607) );
  inv_x1_sg U45009 ( .A(n40607), .X(n40608) );
  inv_x1_sg U45010 ( .A(n40607), .X(n40609) );
  inv_x1_sg U45011 ( .A(n40607), .X(n40610) );
  inv_x1_sg U45012 ( .A(n40607), .X(n40611) );
  inv_x1_sg U45013 ( .A(n6834), .X(n40612) );
  inv_x1_sg U45014 ( .A(n40612), .X(n40613) );
  inv_x1_sg U45015 ( .A(n40612), .X(n40614) );
  inv_x1_sg U45016 ( .A(n40612), .X(n40615) );
  inv_x1_sg U45017 ( .A(n42044), .X(n40616) );
  inv_x1_sg U45018 ( .A(n40616), .X(n40617) );
  inv_x1_sg U45019 ( .A(n40616), .X(n40618) );
  inv_x1_sg U45020 ( .A(n40616), .X(n40619) );
  inv_x1_sg U45021 ( .A(n14363), .X(n40620) );
  inv_x1_sg U45022 ( .A(n40620), .X(n40621) );
  inv_x1_sg U45023 ( .A(n40620), .X(n40622) );
  inv_x1_sg U45024 ( .A(n40620), .X(n40623) );
  inv_x1_sg U45025 ( .A(n40620), .X(n40624) );
  inv_x1_sg U45026 ( .A(n8629), .X(n40625) );
  inv_x1_sg U45027 ( .A(n40625), .X(n40626) );
  inv_x1_sg U45028 ( .A(n40625), .X(n40627) );
  inv_x1_sg U45029 ( .A(n40625), .X(n40628) );
  inv_x1_sg U45030 ( .A(n40625), .X(n40629) );
  inv_x1_sg U45031 ( .A(n7811), .X(n40630) );
  inv_x1_sg U45032 ( .A(n40630), .X(n40631) );
  inv_x1_sg U45033 ( .A(n40630), .X(n40632) );
  inv_x1_sg U45034 ( .A(n40630), .X(n40633) );
  inv_x1_sg U45035 ( .A(n40630), .X(n40634) );
  inv_x1_sg U45036 ( .A(n11906), .X(n40635) );
  inv_x1_sg U45037 ( .A(n40635), .X(n40636) );
  inv_x1_sg U45038 ( .A(n40635), .X(n40637) );
  inv_x1_sg U45039 ( .A(n40635), .X(n40638) );
  inv_x1_sg U45040 ( .A(n40635), .X(n40639) );
  inv_x1_sg U45041 ( .A(n11087), .X(n40640) );
  inv_x1_sg U45042 ( .A(n40640), .X(n40641) );
  inv_x1_sg U45043 ( .A(n40640), .X(n40642) );
  inv_x1_sg U45044 ( .A(n40640), .X(n40643) );
  inv_x1_sg U45045 ( .A(n40640), .X(n40644) );
  inv_x1_sg U45046 ( .A(n17639), .X(n40645) );
  inv_x1_sg U45047 ( .A(n40645), .X(n40646) );
  inv_x1_sg U45048 ( .A(n40645), .X(n40647) );
  inv_x1_sg U45049 ( .A(n40645), .X(n40648) );
  inv_x1_sg U45050 ( .A(n40645), .X(n40649) );
  inv_x1_sg U45051 ( .A(n13544), .X(n40650) );
  inv_x1_sg U45052 ( .A(n40650), .X(n40651) );
  inv_x1_sg U45053 ( .A(n40650), .X(n40652) );
  inv_x1_sg U45054 ( .A(n40650), .X(n40653) );
  inv_x1_sg U45055 ( .A(n40650), .X(n40654) );
  inv_x1_sg U45056 ( .A(n10268), .X(n40655) );
  inv_x1_sg U45057 ( .A(n40655), .X(n40656) );
  inv_x1_sg U45058 ( .A(n40655), .X(n40657) );
  inv_x1_sg U45059 ( .A(n40655), .X(n40658) );
  inv_x1_sg U45060 ( .A(n40655), .X(n40659) );
  inv_x1_sg U45061 ( .A(n12725), .X(n40660) );
  inv_x1_sg U45062 ( .A(n40660), .X(n40661) );
  inv_x1_sg U45063 ( .A(n40660), .X(n40662) );
  inv_x1_sg U45064 ( .A(n40660), .X(n40663) );
  inv_x1_sg U45065 ( .A(n40660), .X(n40664) );
  inv_x1_sg U45066 ( .A(n9449), .X(n40665) );
  inv_x1_sg U45067 ( .A(n40665), .X(n40666) );
  inv_x1_sg U45068 ( .A(n40665), .X(n40667) );
  inv_x1_sg U45069 ( .A(n40665), .X(n40668) );
  inv_x1_sg U45070 ( .A(n40665), .X(n40669) );
  inv_x1_sg U45071 ( .A(n18460), .X(n40670) );
  inv_x1_sg U45072 ( .A(n40670), .X(n40671) );
  inv_x1_sg U45073 ( .A(n40670), .X(n40672) );
  inv_x1_sg U45074 ( .A(n40670), .X(n40673) );
  inv_x1_sg U45075 ( .A(n40670), .X(n40674) );
  inv_x1_sg U45076 ( .A(n16001), .X(n40675) );
  inv_x1_sg U45077 ( .A(n40675), .X(n40676) );
  inv_x1_sg U45078 ( .A(n40675), .X(n40677) );
  inv_x1_sg U45079 ( .A(n40675), .X(n40678) );
  inv_x1_sg U45080 ( .A(n40675), .X(n40679) );
  inv_x1_sg U45081 ( .A(n15182), .X(n40680) );
  inv_x1_sg U45082 ( .A(n40680), .X(n40681) );
  inv_x1_sg U45083 ( .A(n40680), .X(n40682) );
  inv_x1_sg U45084 ( .A(n40680), .X(n40683) );
  inv_x1_sg U45085 ( .A(n40680), .X(n40684) );
  inv_x1_sg U45086 ( .A(n7641), .X(n40685) );
  inv_x1_sg U45087 ( .A(n40685), .X(n40686) );
  inv_x1_sg U45088 ( .A(n38817), .X(n40687) );
  inv_x1_sg U45089 ( .A(n40685), .X(n40688) );
  inv_x1_sg U45090 ( .A(n38817), .X(n40689) );
  inv_x1_sg U45091 ( .A(n8459), .X(n40690) );
  inv_x1_sg U45092 ( .A(n40690), .X(n40691) );
  inv_x1_sg U45093 ( .A(n38818), .X(n40692) );
  inv_x1_sg U45094 ( .A(n40690), .X(n40693) );
  inv_x1_sg U45095 ( .A(n38818), .X(n40694) );
  inv_x1_sg U45096 ( .A(n9279), .X(n40695) );
  inv_x1_sg U45097 ( .A(n40695), .X(n40696) );
  inv_x1_sg U45098 ( .A(n38819), .X(n40697) );
  inv_x1_sg U45099 ( .A(n40695), .X(n40698) );
  inv_x1_sg U45100 ( .A(n38819), .X(n40699) );
  inv_x1_sg U45101 ( .A(n10098), .X(n40700) );
  inv_x1_sg U45102 ( .A(n40700), .X(n40701) );
  inv_x1_sg U45103 ( .A(n38820), .X(n40702) );
  inv_x1_sg U45104 ( .A(n40700), .X(n40703) );
  inv_x1_sg U45105 ( .A(n38820), .X(n40704) );
  inv_x1_sg U45106 ( .A(n10917), .X(n40705) );
  inv_x1_sg U45107 ( .A(n40705), .X(n40706) );
  inv_x1_sg U45108 ( .A(n38821), .X(n40707) );
  inv_x1_sg U45109 ( .A(n40705), .X(n40708) );
  inv_x1_sg U45110 ( .A(n38821), .X(n40709) );
  inv_x1_sg U45111 ( .A(n11736), .X(n40710) );
  inv_x1_sg U45112 ( .A(n40710), .X(n40711) );
  inv_x1_sg U45113 ( .A(n38822), .X(n40712) );
  inv_x1_sg U45114 ( .A(n40710), .X(n40713) );
  inv_x1_sg U45115 ( .A(n38822), .X(n40714) );
  inv_x1_sg U45116 ( .A(n12555), .X(n40715) );
  inv_x1_sg U45117 ( .A(n40715), .X(n40716) );
  inv_x1_sg U45118 ( .A(n38823), .X(n40717) );
  inv_x1_sg U45119 ( .A(n40715), .X(n40718) );
  inv_x1_sg U45120 ( .A(n38823), .X(n40719) );
  inv_x1_sg U45121 ( .A(n13374), .X(n40720) );
  inv_x1_sg U45122 ( .A(n40720), .X(n40721) );
  inv_x1_sg U45123 ( .A(n38824), .X(n40722) );
  inv_x1_sg U45124 ( .A(n40720), .X(n40723) );
  inv_x1_sg U45125 ( .A(n38824), .X(n40724) );
  inv_x1_sg U45126 ( .A(n14193), .X(n40725) );
  inv_x1_sg U45127 ( .A(n40725), .X(n40726) );
  inv_x1_sg U45128 ( .A(n38825), .X(n40727) );
  inv_x1_sg U45129 ( .A(n40725), .X(n40728) );
  inv_x1_sg U45130 ( .A(n38825), .X(n40729) );
  inv_x1_sg U45131 ( .A(n15012), .X(n40730) );
  inv_x1_sg U45132 ( .A(n40730), .X(n40731) );
  inv_x1_sg U45133 ( .A(n38826), .X(n40732) );
  inv_x1_sg U45134 ( .A(n40730), .X(n40733) );
  inv_x1_sg U45135 ( .A(n38826), .X(n40734) );
  inv_x1_sg U45136 ( .A(n15831), .X(n40735) );
  inv_x1_sg U45137 ( .A(n40735), .X(n40736) );
  inv_x1_sg U45138 ( .A(n38827), .X(n40737) );
  inv_x1_sg U45139 ( .A(n40735), .X(n40738) );
  inv_x1_sg U45140 ( .A(n38827), .X(n40739) );
  inv_x1_sg U45141 ( .A(n18290), .X(n40740) );
  inv_x1_sg U45142 ( .A(n40740), .X(n40741) );
  inv_x1_sg U45143 ( .A(n38828), .X(n40742) );
  inv_x1_sg U45144 ( .A(n40740), .X(n40743) );
  inv_x1_sg U45145 ( .A(n38828), .X(n40744) );
  inv_x1_sg U45146 ( .A(n38829), .X(n40745) );
  inv_x1_sg U45147 ( .A(n40745), .X(n40746) );
  inv_x1_sg U45148 ( .A(n40745), .X(n40747) );
  inv_x1_sg U45149 ( .A(n40745), .X(n40748) );
  inv_x1_sg U45150 ( .A(n40745), .X(n40749) );
  inv_x1_sg U45151 ( .A(n39408), .X(n40750) );
  inv_x1_sg U45152 ( .A(n39202), .X(n40751) );
  inv_x1_sg U45153 ( .A(n41521), .X(n40752) );
  inv_x1_sg U45154 ( .A(n38830), .X(n40753) );
  inv_x1_sg U45155 ( .A(n40752), .X(n40754) );
  inv_x1_sg U45156 ( .A(n40752), .X(n40755) );
  inv_x1_sg U45157 ( .A(n40752), .X(n40756) );
  inv_x1_sg U45158 ( .A(n41520), .X(n40757) );
  inv_x1_sg U45159 ( .A(n38833), .X(n40758) );
  inv_x1_sg U45160 ( .A(n40757), .X(n40759) );
  inv_x1_sg U45161 ( .A(n40757), .X(n40760) );
  inv_x1_sg U45162 ( .A(n40757), .X(n40761) );
  inv_x1_sg U45163 ( .A(n41507), .X(n40762) );
  inv_x1_sg U45164 ( .A(n41504), .X(n40763) );
  inv_x1_sg U45165 ( .A(n41517), .X(n40764) );
  inv_x1_sg U45166 ( .A(n38836), .X(n40765) );
  inv_x1_sg U45167 ( .A(n40764), .X(n40766) );
  inv_x1_sg U45168 ( .A(n40764), .X(n40767) );
  inv_x1_sg U45169 ( .A(n40764), .X(n40768) );
  inv_x1_sg U45170 ( .A(n41516), .X(n40769) );
  inv_x1_sg U45171 ( .A(n38839), .X(n40770) );
  inv_x1_sg U45172 ( .A(n40769), .X(n40771) );
  inv_x1_sg U45173 ( .A(n40769), .X(n40772) );
  inv_x1_sg U45174 ( .A(n40769), .X(n40773) );
  inv_x1_sg U45175 ( .A(n39401), .X(n40774) );
  inv_x1_sg U45176 ( .A(n39201), .X(n40775) );
  inv_x1_sg U45177 ( .A(n41513), .X(n40776) );
  inv_x1_sg U45178 ( .A(n38842), .X(n40777) );
  inv_x1_sg U45179 ( .A(n40776), .X(n40778) );
  inv_x1_sg U45180 ( .A(n40776), .X(n40779) );
  inv_x1_sg U45181 ( .A(n40776), .X(n40780) );
  inv_x1_sg U45182 ( .A(n41512), .X(n40781) );
  inv_x1_sg U45183 ( .A(n38845), .X(n40782) );
  inv_x1_sg U45184 ( .A(n40781), .X(n40783) );
  inv_x1_sg U45185 ( .A(n40781), .X(n40784) );
  inv_x1_sg U45186 ( .A(n40781), .X(n40785) );
  inv_x1_sg U45187 ( .A(n39400), .X(n40786) );
  inv_x1_sg U45188 ( .A(n41505), .X(n40787) );
  inv_x1_sg U45189 ( .A(n41509), .X(n40788) );
  inv_x1_sg U45190 ( .A(n40788), .X(n40789) );
  inv_x1_sg U45191 ( .A(n40788), .X(n40790) );
  inv_x1_sg U45192 ( .A(n40788), .X(n40791) );
  inv_x1_sg U45193 ( .A(n38857), .X(n40792) );
  inv_x1_sg U45194 ( .A(n38994), .X(n40793) );
  inv_x1_sg U45195 ( .A(n40793), .X(n40794) );
  inv_x1_sg U45196 ( .A(n40793), .X(n40795) );
  inv_x1_sg U45197 ( .A(n40793), .X(n40796) );
  inv_x1_sg U45198 ( .A(n38830), .X(n40797) );
  inv_x1_sg U45199 ( .A(n39422), .X(n40798) );
  inv_x1_sg U45200 ( .A(n39424), .X(n40799) );
  inv_x1_sg U45201 ( .A(n41501), .X(n40800) );
  inv_x1_sg U45202 ( .A(n40800), .X(n40801) );
  inv_x1_sg U45203 ( .A(n40800), .X(n40802) );
  inv_x1_sg U45204 ( .A(n40800), .X(n40803) );
  inv_x1_sg U45205 ( .A(n39202), .X(n40804) );
  inv_x1_sg U45206 ( .A(n41500), .X(n40805) );
  inv_x1_sg U45207 ( .A(n38850), .X(n40806) );
  inv_x1_sg U45208 ( .A(n40805), .X(n40807) );
  inv_x1_sg U45209 ( .A(n40805), .X(n40808) );
  inv_x1_sg U45210 ( .A(n40805), .X(n40809) );
  inv_x1_sg U45211 ( .A(n39422), .X(n40810) );
  inv_x1_sg U45212 ( .A(n39428), .X(n40811) );
  inv_x1_sg U45213 ( .A(n41497), .X(n40812) );
  inv_x1_sg U45214 ( .A(n38853), .X(n40813) );
  inv_x1_sg U45215 ( .A(n40812), .X(n40814) );
  inv_x1_sg U45216 ( .A(n40812), .X(n40815) );
  inv_x1_sg U45217 ( .A(n40812), .X(n40816) );
  inv_x1_sg U45218 ( .A(n41496), .X(n40817) );
  inv_x1_sg U45219 ( .A(n38992), .X(n40818) );
  inv_x1_sg U45220 ( .A(n40817), .X(n40819) );
  inv_x1_sg U45221 ( .A(n38992), .X(n40820) );
  inv_x1_sg U45222 ( .A(n40817), .X(n40821) );
  inv_x1_sg U45223 ( .A(n39286), .X(n40822) );
  inv_x1_sg U45224 ( .A(n38988), .X(n40823) );
  inv_x1_sg U45225 ( .A(n41493), .X(n40824) );
  inv_x1_sg U45226 ( .A(n38857), .X(n40825) );
  inv_x1_sg U45227 ( .A(n40824), .X(n40826) );
  inv_x1_sg U45228 ( .A(n40824), .X(n40827) );
  inv_x1_sg U45229 ( .A(n40824), .X(n40828) );
  inv_x1_sg U45230 ( .A(n41492), .X(n40829) );
  inv_x1_sg U45231 ( .A(n40829), .X(n40830) );
  inv_x1_sg U45232 ( .A(n40829), .X(n40831) );
  inv_x1_sg U45233 ( .A(n40829), .X(n40832) );
  inv_x1_sg U45234 ( .A(n40836), .X(n40833) );
  inv_x1_sg U45235 ( .A(n39287), .X(n40834) );
  inv_x1_sg U45236 ( .A(n39286), .X(n40835) );
  inv_x1_sg U45237 ( .A(n41489), .X(n40836) );
  inv_x1_sg U45238 ( .A(n38989), .X(n40837) );
  inv_x1_sg U45239 ( .A(n40836), .X(n40838) );
  inv_x1_sg U45240 ( .A(n38989), .X(n40839) );
  inv_x1_sg U45241 ( .A(n40836), .X(n40840) );
  inv_x1_sg U45242 ( .A(n8456), .X(n40841) );
  inv_x1_sg U45243 ( .A(n40841), .X(n40842) );
  inv_x1_sg U45244 ( .A(n40841), .X(n40843) );
  inv_x1_sg U45245 ( .A(n40841), .X(n40844) );
  inv_x1_sg U45246 ( .A(n18288), .X(n40845) );
  inv_x1_sg U45247 ( .A(n40845), .X(n40846) );
  inv_x1_sg U45248 ( .A(n38862), .X(n40847) );
  inv_x1_sg U45249 ( .A(n40845), .X(n40848) );
  inv_x1_sg U45250 ( .A(n38862), .X(n40849) );
  inv_x1_sg U45251 ( .A(n15010), .X(n40850) );
  inv_x1_sg U45252 ( .A(n40850), .X(n40851) );
  inv_x1_sg U45253 ( .A(n38864), .X(n40852) );
  inv_x1_sg U45254 ( .A(n40850), .X(n40853) );
  inv_x1_sg U45255 ( .A(n38864), .X(n40854) );
  inv_x1_sg U45256 ( .A(n14191), .X(n40855) );
  inv_x1_sg U45257 ( .A(n40855), .X(n40856) );
  inv_x1_sg U45258 ( .A(n38866), .X(n40857) );
  inv_x1_sg U45259 ( .A(n40855), .X(n40858) );
  inv_x1_sg U45260 ( .A(n38866), .X(n40859) );
  inv_x1_sg U45261 ( .A(n13372), .X(n40860) );
  inv_x1_sg U45262 ( .A(n40860), .X(n40861) );
  inv_x1_sg U45263 ( .A(n38868), .X(n40862) );
  inv_x1_sg U45264 ( .A(n40860), .X(n40863) );
  inv_x1_sg U45265 ( .A(n38868), .X(n40864) );
  inv_x1_sg U45266 ( .A(n12553), .X(n40865) );
  inv_x1_sg U45267 ( .A(n40865), .X(n40866) );
  inv_x1_sg U45268 ( .A(n38870), .X(n40867) );
  inv_x1_sg U45269 ( .A(n40865), .X(n40868) );
  inv_x1_sg U45270 ( .A(n38870), .X(n40869) );
  inv_x1_sg U45271 ( .A(n11734), .X(n40870) );
  inv_x1_sg U45272 ( .A(n40870), .X(n40871) );
  inv_x1_sg U45273 ( .A(n38872), .X(n40872) );
  inv_x1_sg U45274 ( .A(n40870), .X(n40873) );
  inv_x1_sg U45275 ( .A(n38872), .X(n40874) );
  inv_x1_sg U45276 ( .A(n10915), .X(n40875) );
  inv_x1_sg U45277 ( .A(n40875), .X(n40876) );
  inv_x1_sg U45278 ( .A(n38874), .X(n40877) );
  inv_x1_sg U45279 ( .A(n40875), .X(n40878) );
  inv_x1_sg U45280 ( .A(n38874), .X(n40879) );
  inv_x1_sg U45281 ( .A(n10096), .X(n40880) );
  inv_x1_sg U45282 ( .A(n40880), .X(n40881) );
  inv_x1_sg U45283 ( .A(n38876), .X(n40882) );
  inv_x1_sg U45284 ( .A(n40880), .X(n40883) );
  inv_x1_sg U45285 ( .A(n38876), .X(n40884) );
  inv_x1_sg U45286 ( .A(n9277), .X(n40885) );
  inv_x1_sg U45287 ( .A(n40885), .X(n40886) );
  inv_x1_sg U45288 ( .A(n38878), .X(n40887) );
  inv_x1_sg U45289 ( .A(n40885), .X(n40888) );
  inv_x1_sg U45290 ( .A(n38878), .X(n40889) );
  inv_x1_sg U45291 ( .A(n8457), .X(n40890) );
  inv_x1_sg U45292 ( .A(n40890), .X(n40891) );
  inv_x1_sg U45293 ( .A(n38880), .X(n40892) );
  inv_x1_sg U45294 ( .A(n40890), .X(n40893) );
  inv_x1_sg U45295 ( .A(n38880), .X(n40894) );
  inv_x1_sg U45296 ( .A(n15829), .X(n40895) );
  inv_x1_sg U45297 ( .A(n40895), .X(n40896) );
  inv_x1_sg U45298 ( .A(n38882), .X(n40897) );
  inv_x1_sg U45299 ( .A(n40895), .X(n40898) );
  inv_x1_sg U45300 ( .A(n38882), .X(n40899) );
  inv_x1_sg U45301 ( .A(n16647), .X(n40900) );
  inv_x1_sg U45302 ( .A(n40900), .X(n40901) );
  inv_x1_sg U45303 ( .A(n38884), .X(n40902) );
  inv_x1_sg U45304 ( .A(n40900), .X(n40903) );
  inv_x1_sg U45305 ( .A(n38884), .X(n40904) );
  inv_x1_sg U45306 ( .A(n17467), .X(n40905) );
  inv_x1_sg U45307 ( .A(n40905), .X(n40906) );
  inv_x1_sg U45308 ( .A(n38886), .X(n40907) );
  inv_x1_sg U45309 ( .A(n40905), .X(n40908) );
  inv_x1_sg U45310 ( .A(n38886), .X(n40909) );
  inv_x1_sg U45311 ( .A(n6823), .X(n40910) );
  inv_x1_sg U45312 ( .A(n40910), .X(n40911) );
  inv_x1_sg U45313 ( .A(n38888), .X(n40912) );
  inv_x1_sg U45314 ( .A(n40910), .X(n40913) );
  inv_x1_sg U45315 ( .A(n38888), .X(n40914) );
  inv_x1_sg U45316 ( .A(n7639), .X(n40915) );
  inv_x1_sg U45317 ( .A(n40915), .X(n40916) );
  inv_x1_sg U45318 ( .A(n38890), .X(n40917) );
  inv_x1_sg U45319 ( .A(n40915), .X(n40918) );
  inv_x1_sg U45320 ( .A(n38890), .X(n40919) );
  inv_x1_sg U45321 ( .A(n6822), .X(n40920) );
  inv_x1_sg U45322 ( .A(n40920), .X(n40921) );
  inv_x1_sg U45323 ( .A(n40920), .X(n40922) );
  inv_x1_sg U45324 ( .A(n40920), .X(n40923) );
  inv_x1_sg U45325 ( .A(n16646), .X(n40924) );
  inv_x1_sg U45326 ( .A(n40924), .X(n40925) );
  inv_x1_sg U45327 ( .A(n40924), .X(n40926) );
  inv_x1_sg U45328 ( .A(n40924), .X(n40927) );
  inv_x1_sg U45329 ( .A(n10914), .X(n40928) );
  inv_x1_sg U45330 ( .A(n40928), .X(n40929) );
  inv_x1_sg U45331 ( .A(n40928), .X(n40930) );
  inv_x1_sg U45332 ( .A(n40928), .X(n40931) );
  inv_x1_sg U45333 ( .A(n11733), .X(n40932) );
  inv_x1_sg U45334 ( .A(n40932), .X(n40933) );
  inv_x1_sg U45335 ( .A(n40932), .X(n40934) );
  inv_x1_sg U45336 ( .A(n40932), .X(n40935) );
  inv_x1_sg U45337 ( .A(n12552), .X(n40936) );
  inv_x1_sg U45338 ( .A(n40936), .X(n40937) );
  inv_x1_sg U45339 ( .A(n40936), .X(n40938) );
  inv_x1_sg U45340 ( .A(n40936), .X(n40939) );
  inv_x1_sg U45341 ( .A(n13371), .X(n40940) );
  inv_x1_sg U45342 ( .A(n40940), .X(n40941) );
  inv_x1_sg U45343 ( .A(n40940), .X(n40942) );
  inv_x1_sg U45344 ( .A(n40940), .X(n40943) );
  inv_x1_sg U45345 ( .A(n14190), .X(n40944) );
  inv_x1_sg U45346 ( .A(n40944), .X(n40945) );
  inv_x1_sg U45347 ( .A(n40944), .X(n40946) );
  inv_x1_sg U45348 ( .A(n40944), .X(n40947) );
  inv_x1_sg U45349 ( .A(n15009), .X(n40948) );
  inv_x1_sg U45350 ( .A(n40948), .X(n40949) );
  inv_x1_sg U45351 ( .A(n40948), .X(n40950) );
  inv_x1_sg U45352 ( .A(n40948), .X(n40951) );
  inv_x1_sg U45353 ( .A(n15828), .X(n40952) );
  inv_x1_sg U45354 ( .A(n40952), .X(n40953) );
  inv_x1_sg U45355 ( .A(n40952), .X(n40954) );
  inv_x1_sg U45356 ( .A(n40952), .X(n40955) );
  inv_x1_sg U45357 ( .A(n18287), .X(n40956) );
  inv_x1_sg U45358 ( .A(n40956), .X(n40957) );
  inv_x1_sg U45359 ( .A(n40956), .X(n40958) );
  inv_x1_sg U45360 ( .A(n40956), .X(n40959) );
  inv_x1_sg U45361 ( .A(n10095), .X(n40960) );
  inv_x1_sg U45362 ( .A(n40960), .X(n40961) );
  inv_x1_sg U45363 ( .A(n40960), .X(n40962) );
  inv_x1_sg U45364 ( .A(n40960), .X(n40963) );
  inv_x1_sg U45365 ( .A(n17466), .X(n40964) );
  inv_x1_sg U45366 ( .A(n40964), .X(n40965) );
  inv_x1_sg U45367 ( .A(n40964), .X(n40966) );
  inv_x1_sg U45368 ( .A(n40964), .X(n40967) );
  inv_x1_sg U45369 ( .A(n9276), .X(n40968) );
  inv_x1_sg U45370 ( .A(n40968), .X(n40969) );
  inv_x1_sg U45371 ( .A(n40968), .X(n40970) );
  inv_x1_sg U45372 ( .A(n40968), .X(n40971) );
  inv_x1_sg U45373 ( .A(n7638), .X(n40972) );
  inv_x1_sg U45374 ( .A(n40972), .X(n40973) );
  inv_x1_sg U45375 ( .A(n40972), .X(n40974) );
  inv_x1_sg U45376 ( .A(n40972), .X(n40975) );
  inv_x1_sg U45377 ( .A(n42332), .X(n40976) );
  inv_x1_sg U45378 ( .A(n40976), .X(n40977) );
  inv_x1_sg U45379 ( .A(n40976), .X(n40978) );
  inv_x1_sg U45380 ( .A(n40976), .X(n40979) );
  inv_x1_sg U45381 ( .A(n40976), .X(n40980) );
  inv_x1_sg U45382 ( .A(n41944), .X(n40981) );
  inv_x1_sg U45383 ( .A(n40981), .X(n40982) );
  inv_x1_sg U45384 ( .A(n40981), .X(n40983) );
  inv_x1_sg U45385 ( .A(n40981), .X(n40984) );
  inv_x1_sg U45386 ( .A(n40981), .X(n40985) );
  inv_x1_sg U45387 ( .A(n5987), .X(n40986) );
  inv_x1_sg U45388 ( .A(n38922), .X(n40987) );
  inv_x1_sg U45389 ( .A(n5987), .X(n40988) );
  inv_x1_sg U45390 ( .A(n42385), .X(n40989) );
  inv_x1_sg U45391 ( .A(n38919), .X(n40990) );
  inv_x1_sg U45392 ( .A(n42385), .X(n40991) );
  inv_x1_sg U45393 ( .A(n41931), .X(n40992) );
  inv_x1_sg U45394 ( .A(n40992), .X(n40993) );
  inv_x1_sg U45395 ( .A(n40992), .X(n40994) );
  inv_x1_sg U45396 ( .A(n40992), .X(n40995) );
  inv_x1_sg U45397 ( .A(n40992), .X(n40996) );
  inv_x1_sg U45398 ( .A(n41918), .X(n40997) );
  inv_x1_sg U45399 ( .A(n40997), .X(n40998) );
  inv_x1_sg U45400 ( .A(n38909), .X(n40999) );
  inv_x1_sg U45401 ( .A(n40997), .X(n41000) );
  inv_x1_sg U45402 ( .A(n38909), .X(n41001) );
  inv_x1_sg U45403 ( .A(n41573), .X(n41002) );
  inv_x1_sg U45404 ( .A(n41002), .X(n41003) );
  inv_x1_sg U45405 ( .A(n41002), .X(n41004) );
  inv_x1_sg U45406 ( .A(n41002), .X(n41005) );
  inv_x1_sg U45407 ( .A(n41002), .X(n41006) );
  inv_x1_sg U45408 ( .A(n41572), .X(n41007) );
  inv_x1_sg U45409 ( .A(n41007), .X(n41008) );
  inv_x1_sg U45410 ( .A(n41007), .X(n41009) );
  inv_x1_sg U45411 ( .A(n41007), .X(n41010) );
  inv_x1_sg U45412 ( .A(n41007), .X(n41011) );
  inv_x1_sg U45413 ( .A(n41571), .X(n41012) );
  inv_x1_sg U45414 ( .A(n41012), .X(n41013) );
  inv_x1_sg U45415 ( .A(n41012), .X(n41014) );
  inv_x1_sg U45416 ( .A(n41012), .X(n41015) );
  inv_x1_sg U45417 ( .A(n41012), .X(n41016) );
  inv_x1_sg U45418 ( .A(n41570), .X(n41017) );
  inv_x1_sg U45419 ( .A(n41017), .X(n41018) );
  inv_x1_sg U45420 ( .A(n41017), .X(n41019) );
  inv_x1_sg U45421 ( .A(n41017), .X(n41020) );
  inv_x1_sg U45422 ( .A(n41017), .X(n41021) );
  inv_x1_sg U45423 ( .A(n41569), .X(n41022) );
  inv_x1_sg U45424 ( .A(n41022), .X(n41023) );
  inv_x1_sg U45425 ( .A(n41022), .X(n41024) );
  inv_x1_sg U45426 ( .A(n41022), .X(n41025) );
  inv_x1_sg U45427 ( .A(n41022), .X(n41026) );
  inv_x1_sg U45428 ( .A(n41568), .X(n41027) );
  inv_x1_sg U45429 ( .A(n41027), .X(n41028) );
  inv_x1_sg U45430 ( .A(n41027), .X(n41029) );
  inv_x1_sg U45431 ( .A(n41027), .X(n41030) );
  inv_x1_sg U45432 ( .A(n41027), .X(n41031) );
  inv_x1_sg U45433 ( .A(n41567), .X(n41032) );
  inv_x1_sg U45434 ( .A(n41032), .X(n41033) );
  inv_x1_sg U45435 ( .A(n41032), .X(n41034) );
  inv_x1_sg U45436 ( .A(n41032), .X(n41035) );
  inv_x1_sg U45437 ( .A(n41032), .X(n41036) );
  inv_x1_sg U45438 ( .A(n41566), .X(n41037) );
  inv_x1_sg U45439 ( .A(n41037), .X(n41038) );
  inv_x1_sg U45440 ( .A(n41037), .X(n41039) );
  inv_x1_sg U45441 ( .A(n41037), .X(n41040) );
  inv_x1_sg U45442 ( .A(n41037), .X(n41041) );
  inv_x1_sg U45443 ( .A(n38990), .X(n41042) );
  inv_x1_sg U45444 ( .A(n41042), .X(n41043) );
  inv_x1_sg U45445 ( .A(n38988), .X(n41044) );
  inv_x1_sg U45446 ( .A(n41042), .X(n41045) );
  inv_x1_sg U45447 ( .A(n41042), .X(n41046) );
  inv_x1_sg U45448 ( .A(n26184), .X(n41047) );
  inv_x1_sg U45449 ( .A(n41047), .X(n41048) );
  inv_x1_sg U45450 ( .A(n41047), .X(n41049) );
  inv_x1_sg U45451 ( .A(n41047), .X(n41050) );
  inv_x1_sg U45452 ( .A(n41047), .X(n41051) );
  inv_x1_sg U45453 ( .A(n41270), .X(n41052) );
  inv_x1_sg U45454 ( .A(n41271), .X(n41053) );
  inv_x1_sg U45455 ( .A(n41273), .X(n41054) );
  inv_x1_sg U45456 ( .A(n41273), .X(n41055) );
  inv_x1_sg U45457 ( .A(n41809), .X(n41056) );
  inv_x1_sg U45458 ( .A(n41056), .X(n41057) );
  inv_x1_sg U45459 ( .A(n41056), .X(n41058) );
  inv_x1_sg U45460 ( .A(n41056), .X(n41059) );
  inv_x1_sg U45461 ( .A(n41056), .X(n41060) );
  inv_x1_sg U45462 ( .A(n20961), .X(n41061) );
  inv_x1_sg U45463 ( .A(n41061), .X(n41062) );
  inv_x1_sg U45464 ( .A(n41061), .X(n41063) );
  inv_x1_sg U45465 ( .A(n41061), .X(n41064) );
  inv_x1_sg U45466 ( .A(n5951), .X(n41065) );
  inv_x1_sg U45467 ( .A(n41065), .X(n41066) );
  inv_x1_sg U45468 ( .A(n38916), .X(n41067) );
  inv_x1_sg U45469 ( .A(n41065), .X(n41068) );
  inv_x1_sg U45470 ( .A(n38916), .X(n41069) );
  inv_x1_sg U45471 ( .A(n42385), .X(n41070) );
  inv_x1_sg U45472 ( .A(n41070), .X(n41071) );
  inv_x1_sg U45473 ( .A(n41070), .X(n41072) );
  inv_x1_sg U45474 ( .A(n41070), .X(n41073) );
  inv_x1_sg U45475 ( .A(n41070), .X(n41074) );
  inv_x1_sg U45476 ( .A(n5987), .X(n41075) );
  inv_x1_sg U45477 ( .A(n41075), .X(n41076) );
  inv_x1_sg U45478 ( .A(n41075), .X(n41077) );
  inv_x1_sg U45479 ( .A(n41075), .X(n41078) );
  inv_x1_sg U45480 ( .A(n41075), .X(n41079) );
  inv_x1_sg U45481 ( .A(n19120), .X(n41080) );
  inv_x1_sg U45482 ( .A(n41080), .X(n41081) );
  inv_x1_sg U45483 ( .A(n41080), .X(n41082) );
  inv_x1_sg U45484 ( .A(n41080), .X(n41083) );
  inv_x1_sg U45485 ( .A(n20575), .X(n41084) );
  inv_x1_sg U45486 ( .A(n41084), .X(n41085) );
  inv_x1_sg U45487 ( .A(n41084), .X(n41086) );
  inv_x1_sg U45488 ( .A(n41084), .X(n41087) );
  inv_x1_sg U45489 ( .A(n19118), .X(n41088) );
  inv_x1_sg U45490 ( .A(n41088), .X(n41089) );
  inv_x1_sg U45491 ( .A(n41088), .X(n41090) );
  inv_x1_sg U45492 ( .A(n41088), .X(n41091) );
  inv_x1_sg U45493 ( .A(n20962), .X(n41092) );
  inv_x1_sg U45494 ( .A(n41092), .X(n41093) );
  inv_x1_sg U45495 ( .A(n41092), .X(n41094) );
  inv_x1_sg U45496 ( .A(n41092), .X(n41095) );
  inv_x1_sg U45497 ( .A(n19126), .X(n41096) );
  inv_x1_sg U45498 ( .A(n41096), .X(n41097) );
  inv_x1_sg U45499 ( .A(n41096), .X(n41098) );
  inv_x1_sg U45500 ( .A(n41096), .X(n41099) );
  inv_x1_sg U45501 ( .A(n19124), .X(n41100) );
  inv_x1_sg U45502 ( .A(n41100), .X(n41101) );
  inv_x1_sg U45503 ( .A(n41100), .X(n41102) );
  inv_x1_sg U45504 ( .A(n41100), .X(n41103) );
  inv_x1_sg U45505 ( .A(n20567), .X(n41104) );
  inv_x1_sg U45506 ( .A(n41104), .X(n41105) );
  inv_x1_sg U45507 ( .A(n41104), .X(n41106) );
  inv_x1_sg U45508 ( .A(n41104), .X(n41107) );
  inv_x1_sg U45509 ( .A(n20569), .X(n41108) );
  inv_x1_sg U45510 ( .A(n41108), .X(n41109) );
  inv_x1_sg U45511 ( .A(n41108), .X(n41110) );
  inv_x1_sg U45512 ( .A(n41108), .X(n41111) );
  inv_x1_sg U45513 ( .A(n42372), .X(n41112) );
  inv_x1_sg U45514 ( .A(n41112), .X(n41113) );
  inv_x1_sg U45515 ( .A(n41112), .X(n41114) );
  inv_x1_sg U45516 ( .A(n41112), .X(n41115) );
  inv_x1_sg U45517 ( .A(n42328), .X(n41116) );
  inv_x1_sg U45518 ( .A(n42059), .X(n41117) );
  inv_x1_sg U45519 ( .A(n41116), .X(n41118) );
  inv_x1_sg U45520 ( .A(n42059), .X(n41119) );
  inv_x1_sg U45521 ( .A(n41116), .X(n41120) );
  inv_x1_sg U45522 ( .A(n41946), .X(n41121) );
  inv_x1_sg U45523 ( .A(n39250), .X(n41122) );
  inv_x1_sg U45524 ( .A(n41121), .X(n41123) );
  inv_x1_sg U45525 ( .A(n39250), .X(n41124) );
  inv_x1_sg U45526 ( .A(n41121), .X(n41125) );
  inv_x1_sg U45527 ( .A(n41930), .X(n41126) );
  inv_x1_sg U45528 ( .A(n39247), .X(n41127) );
  inv_x1_sg U45529 ( .A(n41126), .X(n41128) );
  inv_x1_sg U45530 ( .A(n39247), .X(n41129) );
  inv_x1_sg U45531 ( .A(n41126), .X(n41130) );
  inv_x1_sg U45532 ( .A(n41874), .X(n41131) );
  inv_x1_sg U45533 ( .A(n39245), .X(n41132) );
  inv_x1_sg U45534 ( .A(n41131), .X(n41133) );
  inv_x1_sg U45535 ( .A(n39245), .X(n41134) );
  inv_x1_sg U45536 ( .A(n41131), .X(n41135) );
  inv_x1_sg U45537 ( .A(n41873), .X(n41136) );
  inv_x1_sg U45538 ( .A(n39243), .X(n41137) );
  inv_x1_sg U45539 ( .A(n41136), .X(n41138) );
  inv_x1_sg U45540 ( .A(n39243), .X(n41139) );
  inv_x1_sg U45541 ( .A(n41136), .X(n41140) );
  inv_x1_sg U45542 ( .A(n41872), .X(n41141) );
  inv_x1_sg U45543 ( .A(n39241), .X(n41142) );
  inv_x1_sg U45544 ( .A(n41141), .X(n41143) );
  inv_x1_sg U45545 ( .A(n39241), .X(n41144) );
  inv_x1_sg U45546 ( .A(n41141), .X(n41145) );
  inv_x1_sg U45547 ( .A(n41871), .X(n41146) );
  inv_x1_sg U45548 ( .A(n39239), .X(n41147) );
  inv_x1_sg U45549 ( .A(n41146), .X(n41148) );
  inv_x1_sg U45550 ( .A(n39239), .X(n41149) );
  inv_x1_sg U45551 ( .A(n41146), .X(n41150) );
  inv_x1_sg U45552 ( .A(n41870), .X(n41151) );
  inv_x1_sg U45553 ( .A(n39237), .X(n41152) );
  inv_x1_sg U45554 ( .A(n41151), .X(n41153) );
  inv_x1_sg U45555 ( .A(n39237), .X(n41154) );
  inv_x1_sg U45556 ( .A(n41151), .X(n41155) );
  inv_x1_sg U45557 ( .A(n41869), .X(n41156) );
  inv_x1_sg U45558 ( .A(n39235), .X(n41157) );
  inv_x1_sg U45559 ( .A(n41156), .X(n41158) );
  inv_x1_sg U45560 ( .A(n39235), .X(n41159) );
  inv_x1_sg U45561 ( .A(n41156), .X(n41160) );
  inv_x1_sg U45562 ( .A(n41868), .X(n41161) );
  inv_x1_sg U45563 ( .A(n39233), .X(n41162) );
  inv_x1_sg U45564 ( .A(n41161), .X(n41163) );
  inv_x1_sg U45565 ( .A(n39233), .X(n41164) );
  inv_x1_sg U45566 ( .A(n41161), .X(n41165) );
  inv_x1_sg U45567 ( .A(n41867), .X(n41166) );
  inv_x1_sg U45568 ( .A(n39231), .X(n41167) );
  inv_x1_sg U45569 ( .A(n41166), .X(n41168) );
  inv_x1_sg U45570 ( .A(n39231), .X(n41169) );
  inv_x1_sg U45571 ( .A(n41166), .X(n41170) );
  inv_x1_sg U45572 ( .A(n41866), .X(n41171) );
  inv_x1_sg U45573 ( .A(n39229), .X(n41172) );
  inv_x1_sg U45574 ( .A(n41171), .X(n41173) );
  inv_x1_sg U45575 ( .A(n39229), .X(n41174) );
  inv_x1_sg U45576 ( .A(n41171), .X(n41175) );
  inv_x1_sg U45577 ( .A(n41865), .X(n41176) );
  inv_x1_sg U45578 ( .A(n39227), .X(n41177) );
  inv_x1_sg U45579 ( .A(n41176), .X(n41178) );
  inv_x1_sg U45580 ( .A(n39227), .X(n41179) );
  inv_x1_sg U45581 ( .A(n41176), .X(n41180) );
  inv_x1_sg U45582 ( .A(n41864), .X(n41181) );
  inv_x1_sg U45583 ( .A(n39225), .X(n41182) );
  inv_x1_sg U45584 ( .A(n41181), .X(n41183) );
  inv_x1_sg U45585 ( .A(n39225), .X(n41184) );
  inv_x1_sg U45586 ( .A(n41181), .X(n41185) );
  inv_x1_sg U45587 ( .A(n41863), .X(n41186) );
  inv_x1_sg U45588 ( .A(n39223), .X(n41187) );
  inv_x1_sg U45589 ( .A(n41186), .X(n41188) );
  inv_x1_sg U45590 ( .A(n39223), .X(n41189) );
  inv_x1_sg U45591 ( .A(n41186), .X(n41190) );
  inv_x1_sg U45592 ( .A(n41862), .X(n41191) );
  inv_x1_sg U45593 ( .A(n39221), .X(n41192) );
  inv_x1_sg U45594 ( .A(n41191), .X(n41193) );
  inv_x1_sg U45595 ( .A(n39221), .X(n41194) );
  inv_x1_sg U45596 ( .A(n41191), .X(n41195) );
  inv_x1_sg U45597 ( .A(n42383), .X(n41196) );
  inv_x1_sg U45598 ( .A(n39084), .X(n41197) );
  inv_x1_sg U45599 ( .A(n41196), .X(n41198) );
  inv_x1_sg U45600 ( .A(n39084), .X(n41199) );
  inv_x1_sg U45601 ( .A(n41196), .X(n41200) );
  inv_x1_sg U45602 ( .A(\L2_0/n3047 ), .X(n41201) );
  inv_x1_sg U45603 ( .A(n39085), .X(n41202) );
  inv_x1_sg U45604 ( .A(n41201), .X(n41203) );
  inv_x1_sg U45605 ( .A(n39085), .X(n41204) );
  inv_x1_sg U45606 ( .A(n41201), .X(n41205) );
  inv_x1_sg U45607 ( .A(n5779), .X(n41206) );
  inv_x1_sg U45608 ( .A(n41206), .X(n41207) );
  inv_x1_sg U45609 ( .A(n39088), .X(n41208) );
  inv_x1_sg U45610 ( .A(n41206), .X(n41209) );
  inv_x1_sg U45611 ( .A(n42378), .X(n41210) );
  inv_x1_sg U45612 ( .A(n39091), .X(n41211) );
  inv_x1_sg U45613 ( .A(n41210), .X(n41212) );
  inv_x1_sg U45614 ( .A(n39091), .X(n41213) );
  inv_x1_sg U45615 ( .A(n41210), .X(n41214) );
  inv_x1_sg U45616 ( .A(n42338), .X(n41215) );
  inv_x1_sg U45617 ( .A(n39094), .X(n41216) );
  inv_x1_sg U45618 ( .A(n41215), .X(n41217) );
  inv_x1_sg U45619 ( .A(n39094), .X(n41218) );
  inv_x1_sg U45620 ( .A(n41215), .X(n41219) );
  inv_x1_sg U45621 ( .A(\L2_0/n3127 ), .X(n41220) );
  inv_x1_sg U45622 ( .A(n39097), .X(n41221) );
  inv_x1_sg U45623 ( .A(n41220), .X(n41222) );
  inv_x1_sg U45624 ( .A(n39097), .X(n41223) );
  inv_x1_sg U45625 ( .A(n41220), .X(n41224) );
  inv_x1_sg U45626 ( .A(n42381), .X(n41225) );
  inv_x1_sg U45627 ( .A(n39100), .X(n41226) );
  inv_x1_sg U45628 ( .A(n41225), .X(n41227) );
  inv_x1_sg U45629 ( .A(n39100), .X(n41228) );
  inv_x1_sg U45630 ( .A(n41225), .X(n41229) );
  inv_x1_sg U45631 ( .A(\L2_0/n2727 ), .X(n41230) );
  inv_x1_sg U45632 ( .A(n39103), .X(n41231) );
  inv_x1_sg U45633 ( .A(n41230), .X(n41232) );
  inv_x1_sg U45634 ( .A(n39103), .X(n41233) );
  inv_x1_sg U45635 ( .A(n41230), .X(n41234) );
  inv_x1_sg U45636 ( .A(\L2_0/n3367 ), .X(n41235) );
  inv_x1_sg U45637 ( .A(n39106), .X(n41236) );
  inv_x1_sg U45638 ( .A(n41235), .X(n41237) );
  inv_x1_sg U45639 ( .A(n39106), .X(n41238) );
  inv_x1_sg U45640 ( .A(n41235), .X(n41239) );
  inv_x1_sg U45641 ( .A(n42382), .X(n41240) );
  inv_x1_sg U45642 ( .A(n39109), .X(n41241) );
  inv_x1_sg U45643 ( .A(n41240), .X(n41242) );
  inv_x1_sg U45644 ( .A(n39109), .X(n41243) );
  inv_x1_sg U45645 ( .A(n41240), .X(n41244) );
  inv_x1_sg U45646 ( .A(n42384), .X(n41245) );
  inv_x1_sg U45647 ( .A(n39112), .X(n41246) );
  inv_x1_sg U45648 ( .A(n41245), .X(n41247) );
  inv_x1_sg U45649 ( .A(n39112), .X(n41248) );
  inv_x1_sg U45650 ( .A(n41245), .X(n41249) );
  inv_x1_sg U45651 ( .A(n42018), .X(n41250) );
  inv_x1_sg U45652 ( .A(n39115), .X(n41251) );
  inv_x1_sg U45653 ( .A(n41250), .X(n41252) );
  inv_x1_sg U45654 ( .A(n39115), .X(n41253) );
  inv_x1_sg U45655 ( .A(n41250), .X(n41254) );
  inv_x1_sg U45656 ( .A(\L2_0/n2967 ), .X(n41255) );
  inv_x1_sg U45657 ( .A(n39117), .X(n41256) );
  inv_x1_sg U45658 ( .A(n41255), .X(n41257) );
  inv_x1_sg U45659 ( .A(n39117), .X(n41258) );
  inv_x1_sg U45660 ( .A(n41255), .X(n41259) );
  inv_x1_sg U45661 ( .A(n42379), .X(n41260) );
  inv_x1_sg U45662 ( .A(n39120), .X(n41261) );
  inv_x1_sg U45663 ( .A(n41260), .X(n41262) );
  inv_x1_sg U45664 ( .A(n39120), .X(n41263) );
  inv_x1_sg U45665 ( .A(n41260), .X(n41264) );
  inv_x1_sg U45666 ( .A(reg_model), .X(n41265) );
  inv_x1_sg U45667 ( .A(reg_model), .X(n41266) );
  inv_x1_sg U45668 ( .A(n41265), .X(n41267) );
  inv_x1_sg U45669 ( .A(n41265), .X(n41268) );
  inv_x1_sg U45670 ( .A(n41265), .X(n41269) );
  inv_x1_sg U45671 ( .A(n41266), .X(n41270) );
  inv_x1_sg U45672 ( .A(n41266), .X(n41271) );
  inv_x1_sg U45673 ( .A(n41266), .X(n41272) );
  inv_x1_sg U45674 ( .A(n41945), .X(n41273) );
  inv_x1_sg U45675 ( .A(n41945), .X(n41274) );
  inv_x1_sg U45676 ( .A(n5977), .X(n41275) );
  inv_x1_sg U45677 ( .A(n39251), .X(n41276) );
  inv_x1_sg U45678 ( .A(n39252), .X(n41277) );
  inv_x1_sg U45679 ( .A(n41275), .X(n41278) );
  inv_x1_sg U45680 ( .A(n42329), .X(n41279) );
  inv_x1_sg U45681 ( .A(n39125), .X(n41280) );
  inv_x1_sg U45682 ( .A(n41279), .X(n41281) );
  inv_x1_sg U45683 ( .A(n39125), .X(n41282) );
  inv_x1_sg U45684 ( .A(n41279), .X(n41283) );
  inv_x1_sg U45685 ( .A(\L2_0/n3447 ), .X(n41284) );
  inv_x1_sg U45686 ( .A(n39128), .X(n41285) );
  inv_x1_sg U45687 ( .A(n41284), .X(n41286) );
  inv_x1_sg U45688 ( .A(n39128), .X(n41287) );
  inv_x1_sg U45689 ( .A(n41284), .X(n41288) );
  inv_x1_sg U45690 ( .A(n42380), .X(n41289) );
  inv_x1_sg U45691 ( .A(n39131), .X(n41290) );
  inv_x1_sg U45692 ( .A(n41289), .X(n41291) );
  inv_x1_sg U45693 ( .A(n39131), .X(n41292) );
  inv_x1_sg U45694 ( .A(n41289), .X(n41293) );
  inv_x1_sg U45695 ( .A(n41947), .X(n41294) );
  inv_x1_sg U45696 ( .A(n39134), .X(n41295) );
  inv_x1_sg U45697 ( .A(n39134), .X(n41296) );
  inv_x1_sg U45698 ( .A(n41294), .X(n41297) );
  inv_x1_sg U45699 ( .A(n9274), .X(n41298) );
  inv_x1_sg U45700 ( .A(n41298), .X(n41299) );
  inv_x1_sg U45701 ( .A(n39135), .X(n41300) );
  inv_x1_sg U45702 ( .A(n41298), .X(n41301) );
  inv_x1_sg U45703 ( .A(n39135), .X(n41302) );
  inv_x1_sg U45704 ( .A(n41948), .X(n41303) );
  inv_x1_sg U45705 ( .A(n39136), .X(n41304) );
  inv_x1_sg U45706 ( .A(n39136), .X(n41305) );
  inv_x1_sg U45707 ( .A(n39136), .X(n41306) );
  inv_x1_sg U45708 ( .A(n39136), .X(n41307) );
  inv_x1_sg U45709 ( .A(n39656), .X(n41308) );
  inv_x1_sg U45710 ( .A(n39655), .X(n41309) );
  inv_x1_sg U45711 ( .A(n40217), .X(n41310) );
  inv_x1_sg U45712 ( .A(n38813), .X(n41311) );
  inv_x1_sg U45713 ( .A(n38813), .X(n41312) );
  inv_x1_sg U45714 ( .A(n39275), .X(n41313) );
  inv_x1_sg U45715 ( .A(n40224), .X(n41314) );
  inv_x1_sg U45716 ( .A(n39474), .X(n41315) );
  inv_x1_sg U45717 ( .A(n39474), .X(n41316) );
  inv_x1_sg U45718 ( .A(n39474), .X(n41317) );
  inv_x1_sg U45719 ( .A(n39474), .X(n41318) );
  inv_x1_sg U45720 ( .A(n41574), .X(n41319) );
  inv_x1_sg U45721 ( .A(n41319), .X(n41320) );
  inv_x1_sg U45722 ( .A(n39471), .X(n41321) );
  inv_x1_sg U45723 ( .A(n39471), .X(n41322) );
  inv_x1_sg U45724 ( .A(n41319), .X(n41323) );
  inv_x1_sg U45725 ( .A(n25082), .X(n41324) );
  inv_x1_sg U45726 ( .A(n41324), .X(n41325) );
  inv_x1_sg U45727 ( .A(n39468), .X(n41326) );
  inv_x1_sg U45728 ( .A(n39468), .X(n41327) );
  inv_x1_sg U45729 ( .A(n41324), .X(n41328) );
  inv_x1_sg U45730 ( .A(n24803), .X(n41329) );
  inv_x1_sg U45731 ( .A(n41329), .X(n41330) );
  inv_x1_sg U45732 ( .A(n39465), .X(n41331) );
  inv_x1_sg U45733 ( .A(n39465), .X(n41332) );
  inv_x1_sg U45734 ( .A(n41329), .X(n41333) );
  inv_x1_sg U45735 ( .A(n24525), .X(n41334) );
  inv_x1_sg U45736 ( .A(n41334), .X(n41335) );
  inv_x1_sg U45737 ( .A(n39462), .X(n41336) );
  inv_x1_sg U45738 ( .A(n39462), .X(n41337) );
  inv_x1_sg U45739 ( .A(n41334), .X(n41338) );
  inv_x1_sg U45740 ( .A(n42375), .X(n41339) );
  inv_x1_sg U45741 ( .A(n41339), .X(n41340) );
  inv_x1_sg U45742 ( .A(n39459), .X(n41341) );
  inv_x1_sg U45743 ( .A(n39459), .X(n41342) );
  inv_x1_sg U45744 ( .A(n41339), .X(n41343) );
  inv_x1_sg U45745 ( .A(n23409), .X(n41344) );
  inv_x1_sg U45746 ( .A(n41344), .X(n41345) );
  inv_x1_sg U45747 ( .A(n39456), .X(n41346) );
  inv_x1_sg U45748 ( .A(n39456), .X(n41347) );
  inv_x1_sg U45749 ( .A(n41344), .X(n41348) );
  inv_x1_sg U45750 ( .A(n42371), .X(n41349) );
  inv_x1_sg U45751 ( .A(n41349), .X(n41350) );
  inv_x1_sg U45752 ( .A(n39453), .X(n41351) );
  inv_x1_sg U45753 ( .A(n39453), .X(n41352) );
  inv_x1_sg U45754 ( .A(n41349), .X(n41353) );
  inv_x1_sg U45755 ( .A(n42373), .X(n41354) );
  inv_x1_sg U45756 ( .A(n41354), .X(n41355) );
  inv_x1_sg U45757 ( .A(n39450), .X(n41356) );
  inv_x1_sg U45758 ( .A(n39450), .X(n41357) );
  inv_x1_sg U45759 ( .A(n41354), .X(n41358) );
  inv_x1_sg U45760 ( .A(n42374), .X(n41359) );
  inv_x1_sg U45761 ( .A(n41359), .X(n41360) );
  inv_x1_sg U45762 ( .A(n39447), .X(n41361) );
  inv_x1_sg U45763 ( .A(n39447), .X(n41362) );
  inv_x1_sg U45764 ( .A(n41359), .X(n41363) );
  inv_x1_sg U45765 ( .A(n42386), .X(n41364) );
  inv_x1_sg U45766 ( .A(n41364), .X(n41365) );
  inv_x1_sg U45767 ( .A(n39444), .X(n41366) );
  inv_x1_sg U45768 ( .A(n39444), .X(n41367) );
  inv_x1_sg U45769 ( .A(n41364), .X(n41368) );
  inv_x1_sg U45770 ( .A(n42327), .X(n41369) );
  inv_x1_sg U45771 ( .A(n41369), .X(n41370) );
  inv_x1_sg U45772 ( .A(n39441), .X(n41371) );
  inv_x1_sg U45773 ( .A(n39441), .X(n41372) );
  inv_x1_sg U45774 ( .A(n41369), .X(n41373) );
  inv_x1_sg U45775 ( .A(n42376), .X(n41374) );
  inv_x1_sg U45776 ( .A(n41374), .X(n41375) );
  inv_x1_sg U45777 ( .A(n39438), .X(n41376) );
  inv_x1_sg U45778 ( .A(n39438), .X(n41377) );
  inv_x1_sg U45779 ( .A(n41374), .X(n41378) );
  inv_x1_sg U45780 ( .A(n25640), .X(n41379) );
  inv_x1_sg U45781 ( .A(n39138), .X(n41380) );
  inv_x1_sg U45782 ( .A(n39138), .X(n41381) );
  inv_x1_sg U45783 ( .A(n39138), .X(n41382) );
  inv_x1_sg U45784 ( .A(n39138), .X(n41383) );
  inv_x1_sg U45785 ( .A(n42000), .X(n41384) );
  inv_x1_sg U45786 ( .A(n39141), .X(n41385) );
  inv_x1_sg U45787 ( .A(n39141), .X(n41386) );
  inv_x1_sg U45788 ( .A(n39141), .X(n41387) );
  inv_x1_sg U45789 ( .A(n39141), .X(n41388) );
  inv_x1_sg U45790 ( .A(n38916), .X(n41389) );
  inv_x1_sg U45791 ( .A(n39144), .X(n41390) );
  inv_x1_sg U45792 ( .A(n39144), .X(n41391) );
  inv_x1_sg U45793 ( .A(n39144), .X(n41392) );
  inv_x1_sg U45794 ( .A(n41389), .X(n41393) );
  inv_x1_sg U45795 ( .A(n5994), .X(n41394) );
  inv_x1_sg U45796 ( .A(n39147), .X(n41395) );
  inv_x1_sg U45797 ( .A(n41394), .X(n41396) );
  inv_x1_sg U45798 ( .A(n39147), .X(n41397) );
  inv_x1_sg U45799 ( .A(n41394), .X(n41398) );
  inv_x1_sg U45800 ( .A(n39652), .X(n41399) );
  inv_x1_sg U45801 ( .A(n39651), .X(n41400) );
  inv_x1_sg U45802 ( .A(n41400), .X(n41401) );
  inv_x1_sg U45803 ( .A(n39150), .X(n41402) );
  inv_x1_sg U45804 ( .A(n39150), .X(n41403) );
  inv_x1_sg U45805 ( .A(n39150), .X(n41404) );
  inv_x1_sg U45806 ( .A(n41401), .X(n41405) );
  inv_x1_sg U45807 ( .A(n40375), .X(n41406) );
  inv_x1_sg U45808 ( .A(n39153), .X(n41407) );
  inv_x1_sg U45809 ( .A(n39153), .X(n41408) );
  inv_x1_sg U45810 ( .A(n39153), .X(n41409) );
  inv_x1_sg U45811 ( .A(n39153), .X(n41410) );
  inv_x1_sg U45812 ( .A(n41476), .X(n41411) );
  inv_x1_sg U45813 ( .A(n41411), .X(n41412) );
  inv_x1_sg U45814 ( .A(n39156), .X(n41413) );
  inv_x1_sg U45815 ( .A(n41411), .X(n41414) );
  inv_x1_sg U45816 ( .A(n39156), .X(n41415) );
  inv_x1_sg U45817 ( .A(n5954), .X(n41416) );
  inv_x1_sg U45818 ( .A(n41416), .X(n41417) );
  inv_x1_sg U45819 ( .A(n39433), .X(n41418) );
  inv_x1_sg U45820 ( .A(n39433), .X(n41419) );
  inv_x1_sg U45821 ( .A(n41416), .X(n41420) );
  inv_x1_sg U45822 ( .A(n41477), .X(n41421) );
  inv_x1_sg U45823 ( .A(n39769), .X(n41422) );
  inv_x1_sg U45824 ( .A(n41422), .X(n41423) );
  inv_x1_sg U45825 ( .A(n39161), .X(n41424) );
  inv_x1_sg U45826 ( .A(n39160), .X(n41425) );
  inv_x1_sg U45827 ( .A(n39160), .X(n41426) );
  inv_x1_sg U45828 ( .A(n39160), .X(n41427) );
  inv_x1_sg U45829 ( .A(n39165), .X(n41428) );
  inv_x1_sg U45830 ( .A(n39166), .X(n41429) );
  inv_x1_sg U45831 ( .A(n39166), .X(n41430) );
  inv_x1_sg U45832 ( .A(n39165), .X(n41431) );
  inv_x1_sg U45833 ( .A(n38987), .X(n41432) );
  inv_x1_sg U45834 ( .A(n39171), .X(n41433) );
  inv_x1_sg U45835 ( .A(n39170), .X(n41434) );
  inv_x1_sg U45836 ( .A(n39171), .X(n41435) );
  inv_x1_sg U45837 ( .A(n39170), .X(n41436) );
  inv_x1_sg U45838 ( .A(n41478), .X(n41437) );
  inv_x1_sg U45839 ( .A(n39175), .X(n41438) );
  inv_x1_sg U45840 ( .A(n39176), .X(n41439) );
  inv_x1_sg U45841 ( .A(n39175), .X(n41440) );
  inv_x1_sg U45842 ( .A(n39175), .X(n41441) );
  inv_x1_sg U45843 ( .A(n39180), .X(n41442) );
  inv_x1_sg U45844 ( .A(n39181), .X(n41443) );
  inv_x1_sg U45845 ( .A(n39180), .X(n41444) );
  inv_x1_sg U45846 ( .A(n39180), .X(n41445) );
  inv_x1_sg U45847 ( .A(n41474), .X(n41446) );
  inv_x1_sg U45848 ( .A(n39185), .X(n41447) );
  inv_x1_sg U45849 ( .A(n39186), .X(n41448) );
  inv_x1_sg U45850 ( .A(n39186), .X(n41449) );
  inv_x1_sg U45851 ( .A(n39185), .X(n41450) );
  inv_x1_sg U45852 ( .A(n39190), .X(n41451) );
  inv_x1_sg U45853 ( .A(n39191), .X(n41452) );
  inv_x1_sg U45854 ( .A(n39190), .X(n41453) );
  inv_x1_sg U45855 ( .A(n39191), .X(n41454) );
  inv_x1_sg U45856 ( .A(n41472), .X(n41455) );
  inv_x1_sg U45857 ( .A(n39195), .X(n41456) );
  inv_x1_sg U45858 ( .A(n39196), .X(n41457) );
  inv_x1_sg U45859 ( .A(n39195), .X(n41458) );
  inv_x1_sg U45860 ( .A(n39196), .X(n41459) );
  inv_x1_sg U45861 ( .A(n42377), .X(n41460) );
  inv_x1_sg U45862 ( .A(n39656), .X(n41461) );
  inv_x1_sg U45863 ( .A(n41460), .X(n41462) );
  inv_x1_sg U45864 ( .A(n39656), .X(n41463) );
  inv_x1_sg U45865 ( .A(n41460), .X(n41464) );
  inv_x1_sg U45866 ( .A(n41949), .X(n41465) );
  inv_x1_sg U45867 ( .A(n39652), .X(n41466) );
  inv_x1_sg U45868 ( .A(n41465), .X(n41467) );
  inv_x1_sg U45869 ( .A(n39652), .X(n41468) );
  inv_x1_sg U45870 ( .A(n41465), .X(n41469) );
  nor_x1_sg U45871 ( .A(n39727), .B(n41044), .X(n41470) );
  inv_x1_sg U45872 ( .A(n41470), .X(n41471) );
  inv_x1_sg U45873 ( .A(n41471), .X(n41472) );
  inv_x1_sg U45874 ( .A(n41455), .X(n41473) );
  inv_x1_sg U45875 ( .A(n41471), .X(n41474) );
  inv_x1_sg U45876 ( .A(n41446), .X(n41475) );
  inv_x1_sg U45877 ( .A(n41471), .X(n41476) );
  inv_x1_sg U45878 ( .A(n42388), .X(n41477) );
  inv_x1_sg U45879 ( .A(n39768), .X(n41478) );
  inv_x1_sg U45880 ( .A(n38986), .X(n41479) );
  inv_x1_sg U45881 ( .A(n41477), .X(n41480) );
  inv_x1_sg U45882 ( .A(n39769), .X(n41481) );
  inv_x1_sg U45883 ( .A(n39768), .X(n41482) );
  nor_x1_sg U45884 ( .A(n36902), .B(n39135), .X(n41483) );
  inv_x1_sg U45885 ( .A(n41483), .X(n41484) );
  inv_x1_sg U45886 ( .A(n39423), .X(n41485) );
  inv_x1_sg U45887 ( .A(n39423), .X(n41486) );
  inv_x1_sg U45888 ( .A(n41483), .X(n41487) );
  inv_x1_sg U45889 ( .A(n38988), .X(n41488) );
  inv_x1_sg U45890 ( .A(n39428), .X(n41489) );
  inv_x1_sg U45891 ( .A(n41486), .X(n41490) );
  inv_x1_sg U45892 ( .A(n41484), .X(n41491) );
  inv_x1_sg U45893 ( .A(n39424), .X(n41492) );
  inv_x1_sg U45894 ( .A(n41487), .X(n41493) );
  inv_x1_sg U45895 ( .A(n41487), .X(n41494) );
  inv_x1_sg U45896 ( .A(n39422), .X(n41495) );
  inv_x1_sg U45897 ( .A(n41485), .X(n41496) );
  inv_x1_sg U45898 ( .A(n41486), .X(n41497) );
  inv_x1_sg U45899 ( .A(n39428), .X(n41498) );
  inv_x1_sg U45900 ( .A(n41485), .X(n41499) );
  inv_x1_sg U45901 ( .A(n39427), .X(n41500) );
  inv_x1_sg U45902 ( .A(n41484), .X(n41501) );
  inv_x1_sg U45903 ( .A(n39427), .X(n41502) );
  inv_x1_sg U45904 ( .A(n39424), .X(n41503) );
  inv_x1_sg U45905 ( .A(n39399), .X(n41504) );
  inv_x1_sg U45906 ( .A(n39398), .X(n41505) );
  inv_x1_sg U45907 ( .A(n39399), .X(n41506) );
  inv_x1_sg U45908 ( .A(n38814), .X(n41507) );
  inv_x1_sg U45909 ( .A(n39401), .X(n41508) );
  inv_x1_sg U45910 ( .A(n39409), .X(n41509) );
  inv_x1_sg U45911 ( .A(n39401), .X(n41510) );
  inv_x1_sg U45912 ( .A(n39409), .X(n41511) );
  inv_x1_sg U45913 ( .A(n39408), .X(n41512) );
  inv_x1_sg U45914 ( .A(n39400), .X(n41513) );
  inv_x1_sg U45915 ( .A(n39400), .X(n41514) );
  inv_x1_sg U45916 ( .A(n39409), .X(n41515) );
  inv_x1_sg U45917 ( .A(n41484), .X(n41516) );
  inv_x1_sg U45918 ( .A(n41505), .X(n41517) );
  inv_x1_sg U45919 ( .A(n39202), .X(n41518) );
  inv_x1_sg U45920 ( .A(n41505), .X(n41519) );
  inv_x1_sg U45921 ( .A(n41507), .X(n41520) );
  inv_x1_sg U45922 ( .A(n41506), .X(n41521) );
  inv_x1_sg U45923 ( .A(n39202), .X(n41522) );
  inv_x1_sg U45924 ( .A(n41504), .X(n41523) );
  inv_x1_sg U45925 ( .A(n38756), .X(n41524) );
  inv_x1_sg U45926 ( .A(n42359), .X(n41658) );
  inv_x1_sg U45927 ( .A(n17636), .X(n41647) );
  inv_x1_sg U45928 ( .A(n42360), .X(n41659) );
  inv_x1_sg U45929 ( .A(n42361), .X(n41652) );
  inv_x1_sg U45930 ( .A(n42362), .X(n41653) );
  inv_x1_sg U45931 ( .A(n42363), .X(n41654) );
  inv_x1_sg U45932 ( .A(n42364), .X(n41655) );
  inv_x1_sg U45933 ( .A(n42365), .X(n41648) );
  inv_x1_sg U45934 ( .A(n42366), .X(n41649) );
  inv_x1_sg U45935 ( .A(n42367), .X(n41650) );
  inv_x1_sg U45936 ( .A(n42368), .X(n41651) );
  inv_x1_sg U45937 ( .A(n42357), .X(n41656) );
  inv_x1_sg U45938 ( .A(n42358), .X(n41657) );
  nor_x4_sg U45939 ( .A(n42118), .B(out_L1[17]), .X(n28922) );
  inv_x4_sg U45940 ( .A(n28922), .X(n42086) );
  nor_x4_sg U45941 ( .A(n42113), .B(out_L2[17]), .X(n21358) );
  inv_x4_sg U45942 ( .A(n21358), .X(n42081) );
  nor_x4_sg U45943 ( .A(n42117), .B(out_L1[8]), .X(n29187) );
  inv_x4_sg U45944 ( .A(n29187), .X(n42085) );
  nor_x4_sg U45945 ( .A(n42108), .B(out_L2[4]), .X(n21612) );
  inv_x4_sg U45946 ( .A(n21612), .X(n42076) );
  inv_x1_sg U45947 ( .A(n42339), .X(n41525) );
  nand_x1_sg U45948 ( .A(n19839), .B(n19840), .X(n19634) );
  nand_x1_sg U45949 ( .A(n20496), .B(n20497), .X(n20367) );
  nand_x1_sg U45950 ( .A(n20438), .B(n20439), .X(n20288) );
  nand_x1_sg U45951 ( .A(n21265), .B(n21266), .X(n21076) );
  nand_x1_sg U45952 ( .A(n19400), .B(n19401), .X(n19224) );
  nand_x1_sg U45953 ( .A(n19710), .B(n19711), .X(n19490) );
  nand_x1_sg U45954 ( .A(n20206), .B(n20207), .X(n20028) );
  nand_x1_sg U45955 ( .A(n20849), .B(n20850), .X(n20668) );
  nand_x1_sg U45956 ( .A(n20299), .B(n20300), .X(n20143) );
  nand_x1_sg U45957 ( .A(n19323), .B(n46569), .X(n19156) );
  nand_x1_sg U45958 ( .A(n45883), .B(n19223), .X(n6712) );
  nand_x1_sg U45959 ( .A(n28262), .B(n45036), .X(n28133) );
  nand_x1_sg U45960 ( .A(n19699), .B(n46383), .X(n19478) );
  nand_x1_sg U45961 ( .A(n20778), .B(n46594), .X(n19746) );
  nand_x1_sg U45962 ( .A(n20104), .B(n46381), .X(n19899) );
  nand_x1_sg U45963 ( .A(n20952), .B(n46550), .X(n42339) );
  nand_x1_sg U45964 ( .A(n26133), .B(n26148), .X(n16834) );
  inv_x1_sg U45965 ( .A(n5965), .X(n41541) );
  inv_x1_sg U45966 ( .A(n5969), .X(n41542) );
  inv_x1_sg U45967 ( .A(n5964), .X(n41543) );
  inv_x1_sg U45968 ( .A(n6003), .X(n41544) );
  inv_x1_sg U45969 ( .A(n6077), .X(n41545) );
  inv_x1_sg U45970 ( .A(n6087), .X(n41546) );
  inv_x1_sg U45971 ( .A(n5974), .X(n41547) );
  inv_x1_sg U45972 ( .A(n6161), .X(n41548) );
  inv_x1_sg U45973 ( .A(n5968), .X(n41549) );
  inv_x1_sg U45974 ( .A(n6024), .X(n41550) );
  inv_x1_sg U45975 ( .A(n6211), .X(n41551) );
  inv_x1_sg U45976 ( .A(n6071), .X(n41552) );
  inv_x1_sg U45977 ( .A(n6169), .X(n41553) );
  inv_x1_sg U45978 ( .A(n40973), .X(n41554) );
  inv_x1_sg U45979 ( .A(n40969), .X(n41555) );
  inv_x1_sg U45980 ( .A(n40961), .X(n41556) );
  inv_x1_sg U45981 ( .A(n40957), .X(n41557) );
  inv_x1_sg U45982 ( .A(n40953), .X(n41558) );
  inv_x1_sg U45983 ( .A(n40949), .X(n41559) );
  inv_x1_sg U45984 ( .A(n40945), .X(n41560) );
  inv_x1_sg U45985 ( .A(n40941), .X(n41561) );
  inv_x1_sg U45986 ( .A(n40937), .X(n41562) );
  inv_x1_sg U45987 ( .A(n40933), .X(n41563) );
  inv_x1_sg U45988 ( .A(n40929), .X(n41564) );
  inv_x1_sg U45989 ( .A(n40842), .X(n41565) );
  inv_x1_sg U45990 ( .A(n41081), .X(n41566) );
  inv_x1_sg U45991 ( .A(n41093), .X(n41567) );
  inv_x1_sg U45992 ( .A(n41101), .X(n41568) );
  inv_x1_sg U45993 ( .A(n41109), .X(n41569) );
  inv_x1_sg U45994 ( .A(n41105), .X(n41570) );
  inv_x1_sg U45995 ( .A(n41062), .X(n41571) );
  inv_x1_sg U45996 ( .A(n41097), .X(n41572) );
  inv_x1_sg U45997 ( .A(n41089), .X(n41573) );
  inv_x1_sg U45998 ( .A(n41282), .X(n41574) );
  inv_x1_sg U45999 ( .A(n10749), .X(n41575) );
  inv_x1_sg U46000 ( .A(n9930), .X(n41576) );
  inv_x1_sg U46001 ( .A(n9110), .X(n41577) );
  inv_x1_sg U46002 ( .A(n8292), .X(n41578) );
  inv_x1_sg U46003 ( .A(n14025), .X(n41579) );
  inv_x1_sg U46004 ( .A(n13206), .X(n41580) );
  inv_x1_sg U46005 ( .A(n12387), .X(n41581) );
  inv_x1_sg U46006 ( .A(n11568), .X(n41582) );
  inv_x1_sg U46007 ( .A(n18941), .X(n41583) );
  inv_x1_sg U46008 ( .A(n16482), .X(n41584) );
  inv_x1_sg U46009 ( .A(n15663), .X(n41585) );
  inv_x1_sg U46010 ( .A(n14844), .X(n41586) );
  inv_x1_sg U46011 ( .A(n18120), .X(n41587) );
  inv_x1_sg U46012 ( .A(n18635), .X(n41588) );
  inv_x1_sg U46013 ( .A(n16176), .X(n41589) );
  inv_x1_sg U46014 ( .A(n14538), .X(n41590) );
  inv_x1_sg U46015 ( .A(n13719), .X(n41591) );
  inv_x1_sg U46016 ( .A(n12900), .X(n41592) );
  inv_x1_sg U46017 ( .A(n12081), .X(n41593) );
  inv_x1_sg U46018 ( .A(n11262), .X(n41594) );
  inv_x1_sg U46019 ( .A(n10443), .X(n41595) );
  inv_x1_sg U46020 ( .A(n9624), .X(n41596) );
  inv_x1_sg U46021 ( .A(n8804), .X(n41597) );
  inv_x1_sg U46022 ( .A(n16992), .X(n41598) );
  inv_x1_sg U46023 ( .A(n7167), .X(n41599) );
  inv_x1_sg U46024 ( .A(n17814), .X(n41600) );
  inv_x1_sg U46025 ( .A(n15357), .X(n41601) );
  inv_x1_sg U46026 ( .A(n7986), .X(n41602) );
  inv_x1_sg U46027 ( .A(n39317), .X(n41603) );
  inv_x1_sg U46028 ( .A(n39290), .X(n41604) );
  inv_x1_sg U46029 ( .A(n39315), .X(n41605) );
  inv_x1_sg U46030 ( .A(n39313), .X(n41606) );
  inv_x1_sg U46031 ( .A(n39312), .X(n41607) );
  inv_x1_sg U46032 ( .A(n39310), .X(n41608) );
  inv_x1_sg U46033 ( .A(n39308), .X(n41609) );
  inv_x1_sg U46034 ( .A(n39306), .X(n41610) );
  inv_x1_sg U46035 ( .A(n39304), .X(n41611) );
  inv_x1_sg U46036 ( .A(n39302), .X(n41612) );
  inv_x1_sg U46037 ( .A(n39300), .X(n41613) );
  inv_x1_sg U46038 ( .A(n39298), .X(n41614) );
  inv_x1_sg U46039 ( .A(n39296), .X(n41615) );
  inv_x1_sg U46040 ( .A(n39292), .X(n41616) );
  inv_x1_sg U46041 ( .A(n39294), .X(n41617) );
  inv_x1_sg U46042 ( .A(n39364), .X(n41618) );
  inv_x1_sg U46043 ( .A(n39363), .X(n41619) );
  inv_x1_sg U46044 ( .A(n39362), .X(n41620) );
  inv_x1_sg U46045 ( .A(n39361), .X(n41621) );
  inv_x1_sg U46046 ( .A(n39360), .X(n41622) );
  inv_x1_sg U46047 ( .A(n39359), .X(n41623) );
  inv_x1_sg U46048 ( .A(n39357), .X(n41624) );
  inv_x1_sg U46049 ( .A(n39356), .X(n41625) );
  inv_x1_sg U46050 ( .A(n39355), .X(n41626) );
  inv_x1_sg U46051 ( .A(n39354), .X(n41627) );
  inv_x1_sg U46052 ( .A(n39353), .X(n41628) );
  inv_x1_sg U46053 ( .A(n39352), .X(n41629) );
  inv_x1_sg U46054 ( .A(n39351), .X(n41630) );
  inv_x1_sg U46055 ( .A(n39350), .X(n41631) );
  inv_x1_sg U46056 ( .A(reg_num[3]), .X(n41632) );
  inv_x1_sg U46057 ( .A(n42347), .X(n41633) );
  inv_x1_sg U46058 ( .A(n42356), .X(n41634) );
  inv_x1_sg U46059 ( .A(n42346), .X(n41635) );
  inv_x1_sg U46060 ( .A(n42351), .X(n41636) );
  inv_x1_sg U46061 ( .A(n42350), .X(n41637) );
  inv_x1_sg U46062 ( .A(n42349), .X(n41638) );
  inv_x1_sg U46063 ( .A(n42348), .X(n41639) );
  inv_x1_sg U46064 ( .A(n42355), .X(n41640) );
  inv_x1_sg U46065 ( .A(n42354), .X(n41641) );
  inv_x1_sg U46066 ( .A(n42353), .X(n41642) );
  inv_x1_sg U46067 ( .A(n42352), .X(n41643) );
  inv_x1_sg U46068 ( .A(n42336), .X(n41644) );
  inv_x1_sg U46069 ( .A(n42345), .X(n41645) );
  inv_x1_sg U46070 ( .A(n42344), .X(n41646) );
  inv_x1_sg U46071 ( .A(n39486), .X(n41660) );
  inv_x1_sg U46072 ( .A(n6991), .X(n41661) );
  inv_x1_sg U46073 ( .A(n42160), .X(n41662) );
  inv_x1_sg U46074 ( .A(n39897), .X(n41663) );
  inv_x1_sg U46075 ( .A(n42161), .X(n41664) );
  inv_x1_sg U46076 ( .A(n39894), .X(n41665) );
  inv_x1_sg U46077 ( .A(n7474), .X(n41666) );
  inv_x1_sg U46078 ( .A(n18767), .X(n41667) );
  inv_x1_sg U46079 ( .A(n39891), .X(n41668) );
  inv_x1_sg U46080 ( .A(n17946), .X(n41669) );
  inv_x1_sg U46081 ( .A(n39888), .X(n41670) );
  inv_x1_sg U46082 ( .A(n17125), .X(n41671) );
  inv_x1_sg U46083 ( .A(n39885), .X(n41672) );
  inv_x1_sg U46084 ( .A(n16308), .X(n41673) );
  inv_x1_sg U46085 ( .A(n39882), .X(n41674) );
  inv_x1_sg U46086 ( .A(n14670), .X(n41675) );
  inv_x1_sg U46087 ( .A(n39879), .X(n41676) );
  inv_x1_sg U46088 ( .A(n13851), .X(n41677) );
  inv_x1_sg U46089 ( .A(n39876), .X(n41678) );
  inv_x1_sg U46090 ( .A(n13032), .X(n41679) );
  inv_x1_sg U46091 ( .A(n39873), .X(n41680) );
  inv_x1_sg U46092 ( .A(n12213), .X(n41681) );
  inv_x1_sg U46093 ( .A(n39870), .X(n41682) );
  inv_x1_sg U46094 ( .A(n11394), .X(n41683) );
  inv_x1_sg U46095 ( .A(n39867), .X(n41684) );
  inv_x1_sg U46096 ( .A(n10575), .X(n41685) );
  inv_x1_sg U46097 ( .A(n39864), .X(n41686) );
  inv_x1_sg U46098 ( .A(n8936), .X(n41687) );
  inv_x1_sg U46099 ( .A(n39861), .X(n41688) );
  inv_x1_sg U46100 ( .A(n9756), .X(n41689) );
  inv_x1_sg U46101 ( .A(n39858), .X(n41690) );
  inv_x1_sg U46102 ( .A(n7300), .X(n41691) );
  inv_x1_sg U46103 ( .A(n39855), .X(n41692) );
  inv_x1_sg U46104 ( .A(n39662), .X(n41693) );
  inv_x1_sg U46105 ( .A(n39661), .X(n41694) );
  inv_x1_sg U46106 ( .A(n40132), .X(n41695) );
  inv_x1_sg U46107 ( .A(n40128), .X(n41696) );
  inv_x1_sg U46108 ( .A(n40126), .X(n41697) );
  inv_x1_sg U46109 ( .A(n40124), .X(n41698) );
  inv_x1_sg U46110 ( .A(n40122), .X(n41699) );
  inv_x1_sg U46111 ( .A(n40120), .X(n41700) );
  inv_x1_sg U46112 ( .A(n40118), .X(n41701) );
  inv_x1_sg U46113 ( .A(n40116), .X(n41702) );
  inv_x1_sg U46114 ( .A(n40114), .X(n41703) );
  inv_x1_sg U46115 ( .A(n40112), .X(n41704) );
  inv_x1_sg U46116 ( .A(n40110), .X(n41705) );
  inv_x1_sg U46117 ( .A(n40108), .X(n41706) );
  inv_x1_sg U46118 ( .A(n40106), .X(n41707) );
  inv_x1_sg U46119 ( .A(n40130), .X(n41708) );
  inv_x1_sg U46120 ( .A(n39805), .X(n41709) );
  inv_x1_sg U46121 ( .A(n39802), .X(n41710) );
  inv_x1_sg U46122 ( .A(n39800), .X(n41711) );
  inv_x1_sg U46123 ( .A(n39798), .X(n41712) );
  inv_x1_sg U46124 ( .A(n39796), .X(n41713) );
  inv_x1_sg U46125 ( .A(n39794), .X(n41714) );
  inv_x1_sg U46126 ( .A(n39792), .X(n41715) );
  inv_x1_sg U46127 ( .A(n39790), .X(n41716) );
  inv_x1_sg U46128 ( .A(n39788), .X(n41717) );
  inv_x1_sg U46129 ( .A(n39786), .X(n41718) );
  inv_x1_sg U46130 ( .A(n39784), .X(n41719) );
  inv_x1_sg U46131 ( .A(n39782), .X(n41720) );
  inv_x1_sg U46132 ( .A(n39780), .X(n41721) );
  inv_x1_sg U46133 ( .A(n39778), .X(n41722) );
  inv_x1_sg U46134 ( .A(n39776), .X(n41723) );
  inv_x1_sg U46135 ( .A(n39774), .X(n41724) );
  inv_x1_sg U46136 ( .A(n39772), .X(n41725) );
  inv_x1_sg U46137 ( .A(n39961), .X(n41726) );
  inv_x1_sg U46138 ( .A(n39959), .X(n41727) );
  inv_x1_sg U46139 ( .A(n39955), .X(n41728) );
  inv_x1_sg U46140 ( .A(n39953), .X(n41729) );
  inv_x1_sg U46141 ( .A(n39951), .X(n41730) );
  inv_x1_sg U46142 ( .A(n39949), .X(n41731) );
  inv_x1_sg U46143 ( .A(n39947), .X(n41732) );
  inv_x1_sg U46144 ( .A(n39945), .X(n41733) );
  inv_x1_sg U46145 ( .A(n39943), .X(n41734) );
  inv_x1_sg U46146 ( .A(n39941), .X(n41735) );
  inv_x1_sg U46147 ( .A(n39939), .X(n41736) );
  inv_x1_sg U46148 ( .A(n39937), .X(n41737) );
  inv_x1_sg U46149 ( .A(n39935), .X(n41738) );
  inv_x1_sg U46150 ( .A(n39933), .X(n41739) );
  inv_x1_sg U46151 ( .A(n40095), .X(n41740) );
  inv_x1_sg U46152 ( .A(n17757), .X(n41741) );
  inv_x1_sg U46153 ( .A(n8747), .X(n41742) );
  inv_x1_sg U46154 ( .A(n9567), .X(n41743) );
  inv_x1_sg U46155 ( .A(n10386), .X(n41744) );
  inv_x1_sg U46156 ( .A(n11205), .X(n41745) );
  inv_x1_sg U46157 ( .A(n12024), .X(n41746) );
  inv_x1_sg U46158 ( .A(n12843), .X(n41747) );
  inv_x1_sg U46159 ( .A(n14481), .X(n41748) );
  inv_x1_sg U46160 ( .A(n18578), .X(n41749) );
  inv_x1_sg U46161 ( .A(n7929), .X(n41750) );
  inv_x1_sg U46162 ( .A(n13662), .X(n41751) );
  inv_x1_sg U46163 ( .A(n15300), .X(n41752) );
  inv_x1_sg U46164 ( .A(n16119), .X(n41753) );
  inv_x1_sg U46165 ( .A(n40360), .X(n41754) );
  inv_x1_sg U46166 ( .A(n40159), .X(n41755) );
  inv_x1_sg U46167 ( .A(n40356), .X(n41756) );
  inv_x1_sg U46168 ( .A(n40352), .X(n41757) );
  inv_x1_sg U46169 ( .A(n40348), .X(n41758) );
  inv_x1_sg U46170 ( .A(n40344), .X(n41759) );
  inv_x1_sg U46171 ( .A(n40340), .X(n41760) );
  inv_x1_sg U46172 ( .A(n40336), .X(n41761) );
  inv_x1_sg U46173 ( .A(n40332), .X(n41762) );
  inv_x1_sg U46174 ( .A(n40328), .X(n41763) );
  inv_x1_sg U46175 ( .A(n40324), .X(n41764) );
  inv_x1_sg U46176 ( .A(n40320), .X(n41765) );
  inv_x1_sg U46177 ( .A(n40155), .X(n41766) );
  inv_x1_sg U46178 ( .A(n40153), .X(n41767) );
  inv_x1_sg U46179 ( .A(n40151), .X(n41768) );
  inv_x1_sg U46180 ( .A(n40149), .X(n41769) );
  inv_x1_sg U46181 ( .A(n40147), .X(n41770) );
  inv_x1_sg U46182 ( .A(n40145), .X(n41771) );
  inv_x1_sg U46183 ( .A(n40143), .X(n41772) );
  inv_x1_sg U46184 ( .A(n40141), .X(n41773) );
  inv_x1_sg U46185 ( .A(n40139), .X(n41774) );
  inv_x1_sg U46186 ( .A(n40137), .X(n41775) );
  inv_x1_sg U46187 ( .A(n40135), .X(n41776) );
  inv_x1_sg U46188 ( .A(n40133), .X(n41777) );
  inv_x1_sg U46189 ( .A(n40230), .X(n41778) );
  inv_x1_sg U46190 ( .A(n40234), .X(n41779) );
  inv_x1_sg U46191 ( .A(n7094), .X(n41780) );
  inv_x1_sg U46192 ( .A(n39722), .X(n41781) );
  inv_x1_sg U46193 ( .A(n7912), .X(n41782) );
  inv_x1_sg U46194 ( .A(n39719), .X(n41783) );
  inv_x1_sg U46195 ( .A(n8730), .X(n41784) );
  inv_x1_sg U46196 ( .A(n39716), .X(n41785) );
  inv_x1_sg U46197 ( .A(n9550), .X(n41786) );
  inv_x1_sg U46198 ( .A(n39713), .X(n41787) );
  inv_x1_sg U46199 ( .A(n10369), .X(n41788) );
  inv_x1_sg U46200 ( .A(n39710), .X(n41789) );
  inv_x1_sg U46201 ( .A(n11188), .X(n41790) );
  inv_x1_sg U46202 ( .A(n39707), .X(n41791) );
  inv_x1_sg U46203 ( .A(n12007), .X(n41792) );
  inv_x1_sg U46204 ( .A(n39704), .X(n41793) );
  inv_x1_sg U46205 ( .A(n12826), .X(n41794) );
  inv_x1_sg U46206 ( .A(n39701), .X(n41795) );
  inv_x1_sg U46207 ( .A(n13645), .X(n41796) );
  inv_x1_sg U46208 ( .A(n39698), .X(n41797) );
  inv_x1_sg U46209 ( .A(n14464), .X(n41798) );
  inv_x1_sg U46210 ( .A(n39695), .X(n41799) );
  inv_x1_sg U46211 ( .A(n15283), .X(n41800) );
  inv_x1_sg U46212 ( .A(n39692), .X(n41801) );
  inv_x1_sg U46213 ( .A(n16102), .X(n41802) );
  inv_x1_sg U46214 ( .A(n39689), .X(n41803) );
  inv_x1_sg U46215 ( .A(n17740), .X(n41804) );
  inv_x1_sg U46216 ( .A(n39686), .X(n41805) );
  inv_x1_sg U46217 ( .A(n18561), .X(n41806) );
  inv_x1_sg U46218 ( .A(n39683), .X(n41807) );
  inv_x1_sg U46219 ( .A(n40614), .X(n41808) );
  inv_x1_sg U46220 ( .A(n40315), .X(n41809) );
  inv_x1_sg U46221 ( .A(n40216), .X(n41810) );
  inv_x1_sg U46222 ( .A(n40215), .X(n41811) );
  inv_x1_sg U46223 ( .A(n40184), .X(n41812) );
  inv_x1_sg U46224 ( .A(n40183), .X(n41813) );
  inv_x1_sg U46225 ( .A(n40168), .X(n41814) );
  inv_x1_sg U46226 ( .A(n40167), .X(n41815) );
  inv_x1_sg U46227 ( .A(n40172), .X(n41816) );
  inv_x1_sg U46228 ( .A(n40171), .X(n41817) );
  inv_x1_sg U46229 ( .A(n40188), .X(n41818) );
  inv_x1_sg U46230 ( .A(n40187), .X(n41819) );
  inv_x1_sg U46231 ( .A(n40176), .X(n41820) );
  inv_x1_sg U46232 ( .A(n40175), .X(n41821) );
  inv_x1_sg U46233 ( .A(n40192), .X(n41822) );
  inv_x1_sg U46234 ( .A(n40191), .X(n41823) );
  inv_x1_sg U46235 ( .A(n40196), .X(n41824) );
  inv_x1_sg U46236 ( .A(n40195), .X(n41825) );
  inv_x1_sg U46237 ( .A(n40200), .X(n41826) );
  inv_x1_sg U46238 ( .A(n40199), .X(n41827) );
  inv_x1_sg U46239 ( .A(n40204), .X(n41828) );
  inv_x1_sg U46240 ( .A(n40203), .X(n41829) );
  inv_x1_sg U46241 ( .A(n40208), .X(n41830) );
  inv_x1_sg U46242 ( .A(n40207), .X(n41831) );
  inv_x1_sg U46243 ( .A(n40212), .X(n41832) );
  inv_x1_sg U46244 ( .A(n40211), .X(n41833) );
  inv_x1_sg U46245 ( .A(n40180), .X(n41834) );
  inv_x1_sg U46246 ( .A(n40179), .X(n41835) );
  inv_x1_sg U46247 ( .A(n40342), .X(n41836) );
  inv_x1_sg U46248 ( .A(n40344), .X(n41837) );
  inv_x1_sg U46249 ( .A(n40322), .X(n41838) );
  inv_x1_sg U46250 ( .A(n40324), .X(n41839) );
  inv_x1_sg U46251 ( .A(n40330), .X(n41840) );
  inv_x1_sg U46252 ( .A(n40332), .X(n41841) );
  inv_x1_sg U46253 ( .A(n40070), .X(n41842) );
  inv_x1_sg U46254 ( .A(n40358), .X(n41843) );
  inv_x1_sg U46255 ( .A(n40361), .X(n41844) );
  inv_x1_sg U46256 ( .A(n40318), .X(n41845) );
  inv_x1_sg U46257 ( .A(n40320), .X(n41846) );
  inv_x1_sg U46258 ( .A(n40158), .X(n41847) );
  inv_x1_sg U46259 ( .A(n40334), .X(n41848) );
  inv_x1_sg U46260 ( .A(n40336), .X(n41849) );
  inv_x1_sg U46261 ( .A(n40346), .X(n41850) );
  inv_x1_sg U46262 ( .A(n40348), .X(n41851) );
  inv_x1_sg U46263 ( .A(n40354), .X(n41852) );
  inv_x1_sg U46264 ( .A(n40356), .X(n41853) );
  inv_x1_sg U46265 ( .A(n40350), .X(n41854) );
  inv_x1_sg U46266 ( .A(n40352), .X(n41855) );
  inv_x1_sg U46267 ( .A(n40326), .X(n41856) );
  inv_x1_sg U46268 ( .A(n40328), .X(n41857) );
  inv_x1_sg U46269 ( .A(n40338), .X(n41858) );
  inv_x1_sg U46270 ( .A(n40340), .X(n41859) );
  inv_x1_sg U46271 ( .A(n40578), .X(n41860) );
  inv_x1_sg U46272 ( .A(n40573), .X(n41861) );
  inv_x1_sg U46273 ( .A(n40507), .X(n41862) );
  inv_x1_sg U46274 ( .A(n40503), .X(n41863) );
  inv_x1_sg U46275 ( .A(n40499), .X(n41864) );
  inv_x1_sg U46276 ( .A(n40495), .X(n41865) );
  inv_x1_sg U46277 ( .A(n40491), .X(n41866) );
  inv_x1_sg U46278 ( .A(n40487), .X(n41867) );
  inv_x1_sg U46279 ( .A(n40483), .X(n41868) );
  inv_x1_sg U46280 ( .A(n40479), .X(n41869) );
  inv_x1_sg U46281 ( .A(n40475), .X(n41870) );
  inv_x1_sg U46282 ( .A(n40471), .X(n41871) );
  inv_x1_sg U46283 ( .A(n40467), .X(n41872) );
  inv_x1_sg U46284 ( .A(n40463), .X(n41873) );
  inv_x1_sg U46285 ( .A(n40459), .X(n41874) );
  inv_x1_sg U46286 ( .A(n40055), .X(n41875) );
  inv_x1_sg U46287 ( .A(n42122), .X(n41876) );
  inv_x1_sg U46288 ( .A(n40043), .X(n41877) );
  inv_x1_sg U46289 ( .A(n9539), .X(n41878) );
  inv_x1_sg U46290 ( .A(n40053), .X(n41879) );
  inv_x1_sg U46291 ( .A(n42124), .X(n41880) );
  inv_x1_sg U46292 ( .A(n40065), .X(n41881) );
  inv_x1_sg U46293 ( .A(n13634), .X(n41882) );
  inv_x1_sg U46294 ( .A(n40049), .X(n41883) );
  inv_x1_sg U46295 ( .A(n11996), .X(n41884) );
  inv_x1_sg U46296 ( .A(n40047), .X(n41885) );
  inv_x1_sg U46297 ( .A(n42126), .X(n41886) );
  inv_x1_sg U46298 ( .A(n40041), .X(n41887) );
  inv_x1_sg U46299 ( .A(n42130), .X(n41888) );
  inv_x1_sg U46300 ( .A(n40059), .X(n41889) );
  inv_x1_sg U46301 ( .A(n17729), .X(n41890) );
  inv_x1_sg U46302 ( .A(n40061), .X(n41891) );
  inv_x1_sg U46303 ( .A(n18550), .X(n41892) );
  inv_x1_sg U46304 ( .A(n40057), .X(n41893) );
  inv_x1_sg U46305 ( .A(n16091), .X(n41894) );
  inv_x1_sg U46306 ( .A(n40051), .X(n41895) );
  inv_x1_sg U46307 ( .A(n12815), .X(n41896) );
  inv_x1_sg U46308 ( .A(n40045), .X(n41897) );
  inv_x1_sg U46309 ( .A(n10358), .X(n41898) );
  inv_x1_sg U46310 ( .A(n40063), .X(n41899) );
  inv_x1_sg U46311 ( .A(n42089), .X(n41900) );
  inv_x1_sg U46312 ( .A(n40039), .X(n41901) );
  inv_x1_sg U46313 ( .A(n42325), .X(n41902) );
  inv_x1_sg U46314 ( .A(n39957), .X(n41903) );
  inv_x1_sg U46315 ( .A(n40682), .X(n41904) );
  inv_x1_sg U46316 ( .A(n40677), .X(n41905) );
  inv_x1_sg U46317 ( .A(n40672), .X(n41906) );
  inv_x1_sg U46318 ( .A(n40667), .X(n41907) );
  inv_x1_sg U46319 ( .A(n40662), .X(n41908) );
  inv_x1_sg U46320 ( .A(n40657), .X(n41909) );
  inv_x1_sg U46321 ( .A(n40742), .X(n41910) );
  inv_x1_sg U46322 ( .A(n40652), .X(n41911) );
  inv_x1_sg U46323 ( .A(n40646), .X(n41912) );
  inv_x1_sg U46324 ( .A(n40642), .X(n41913) );
  inv_x1_sg U46325 ( .A(n40637), .X(n41914) );
  inv_x1_sg U46326 ( .A(n40632), .X(n41915) );
  inv_x1_sg U46327 ( .A(n40627), .X(n41916) );
  inv_x1_sg U46328 ( .A(n40622), .X(n41917) );
  inv_x1_sg U46329 ( .A(n40619), .X(n41918) );
  inv_x1_sg U46330 ( .A(n40737), .X(n41919) );
  inv_x1_sg U46331 ( .A(n40732), .X(n41920) );
  inv_x1_sg U46332 ( .A(n40727), .X(n41921) );
  inv_x1_sg U46333 ( .A(n40722), .X(n41922) );
  inv_x1_sg U46334 ( .A(n40717), .X(n41923) );
  inv_x1_sg U46335 ( .A(n40712), .X(n41924) );
  inv_x1_sg U46336 ( .A(n40707), .X(n41925) );
  inv_x1_sg U46337 ( .A(n40702), .X(n41926) );
  inv_x1_sg U46338 ( .A(n40697), .X(n41927) );
  inv_x1_sg U46339 ( .A(n40692), .X(n41928) );
  inv_x1_sg U46340 ( .A(n40687), .X(n41929) );
  inv_x1_sg U46341 ( .A(n41051), .X(n41930) );
  inv_x1_sg U46342 ( .A(n40569), .X(n41931) );
  inv_x1_sg U46343 ( .A(n40729), .X(n41932) );
  inv_x1_sg U46344 ( .A(n40699), .X(n41933) );
  inv_x1_sg U46345 ( .A(n40734), .X(n41934) );
  inv_x1_sg U46346 ( .A(n40719), .X(n41935) );
  inv_x1_sg U46347 ( .A(n40704), .X(n41936) );
  inv_x1_sg U46348 ( .A(n40689), .X(n41937) );
  inv_x1_sg U46349 ( .A(n40724), .X(n41938) );
  inv_x1_sg U46350 ( .A(n40709), .X(n41939) );
  inv_x1_sg U46351 ( .A(n40694), .X(n41940) );
  inv_x1_sg U46352 ( .A(n40744), .X(n41941) );
  inv_x1_sg U46353 ( .A(n40739), .X(n41942) );
  inv_x1_sg U46354 ( .A(n40714), .X(n41943) );
  inv_x1_sg U46355 ( .A(n41113), .X(n41944) );
  inv_x1_sg U46356 ( .A(reg_model), .X(n41945) );
  inv_x1_sg U46357 ( .A(n39124), .X(n41946) );
  inv_x1_sg U46358 ( .A(n40037), .X(n41947) );
  inv_x1_sg U46359 ( .A(n39349), .X(n41948) );
  inv_x1_sg U46360 ( .A(n39927), .X(n41949) );
  nand_x8_sg U46361 ( .A(n38120), .B(input_ready), .X(n36902) );
  inv_x2_sg U46362 ( .A(n21600), .X(n45871) );
  inv_x2_sg U46363 ( .A(n29151), .X(n45023) );
  inv_x2_sg U46364 ( .A(n29163), .X(n45113) );
  inv_x2_sg U46365 ( .A(n29175), .X(n45204) );
  inv_x2_sg U46366 ( .A(n21660), .X(n46327) );
  inv_x2_sg U46367 ( .A(n21648), .X(n46236) );
  inv_x2_sg U46368 ( .A(n21636), .X(n46145) );
  inv_x2_sg U46369 ( .A(n21624), .X(n46054) );
  nand_x16_sg U46370 ( .A(n21594), .B(n21715), .X(n21598) );
  nor_x2_sg U46371 ( .A(n41950), .B(out_L2[1]), .X(n41952) );
  nor_x2_sg U46372 ( .A(n41950), .B(out_L2[1]), .X(n21593) );
  nand_x8_sg U46373 ( .A(n21598), .B(n42107), .X(n21712) );
  nand_x16_sg U46374 ( .A(out_L2[1]), .B(n41950), .X(n21594) );
  nor_x1_sg U46375 ( .A(n19346), .B(n19347), .X(n19322) );
  nor_x1_sg U46376 ( .A(n19783), .B(n19784), .X(n19722) );
  nor_x1_sg U46377 ( .A(n20159), .B(n20160), .X(n20116) );
  nand_x1_sg U46378 ( .A(n44970), .B(n27800), .X(n22574) );
  nand_x1_sg U46379 ( .A(n44965), .B(n28621), .X(n22578) );
  nand_x8_sg U46380 ( .A(n22574), .B(n38191), .X(n27616) );
  nand_x8_sg U46381 ( .A(n22578), .B(n38192), .X(n28462) );
  nand_x8_sg U46382 ( .A(n22584), .B(n38193), .X(n28255) );
  nand_x2_sg U46383 ( .A(n46583), .B(n5684), .X(n20981) );
  nand_x2_sg U46384 ( .A(n45739), .B(n5399), .X(n28539) );
  nor_x1_sg U46385 ( .A(n19948), .B(n19949), .X(n19761) );
  nor_x1_sg U46386 ( .A(n21204), .B(n21205), .X(n21005) );
  nor_x1_sg U46387 ( .A(n19571), .B(n19572), .X(n19337) );
  nand_x8_sg U46388 ( .A(n5719), .B(n44964), .X(n28980) );
  nand_x1_sg U46389 ( .A(n41299), .B(n18285), .X(n42380) );
  nor_x1_sg U46390 ( .A(n21246), .B(n21247), .X(n21092) );
  nor_x1_sg U46391 ( .A(n19960), .B(n19961), .X(n19773) );
  nor_x1_sg U46392 ( .A(n20152), .B(n20153), .X(n19956) );
  nor_x1_sg U46393 ( .A(n20478), .B(n20479), .X(n20383) );
  nor_x1_sg U46394 ( .A(n20313), .B(n20314), .X(n20148) );
  nor_x1_sg U46395 ( .A(n19821), .B(n19822), .X(n19650) );
  nor_x1_sg U46396 ( .A(n19973), .B(n19974), .X(n19903) );
  nand_x1_sg U46397 ( .A(n41300), .B(n19105), .X(n42379) );
  nand_x1_sg U46398 ( .A(n38942), .B(n13370), .X(\L2_0/n2967 ) );
  nor_x1_sg U46399 ( .A(n38555), .B(out_L1[1]), .X(n41951) );
  nand_x1_sg U46400 ( .A(n39133), .B(n18284), .X(n42059) );
  nand_x4_sg U46401 ( .A(n26797), .B(n39486), .X(n42018) );
  nand_x1_sg U46402 ( .A(n38984), .B(n41286), .X(n7638) );
  nand_x1_sg U46403 ( .A(n41301), .B(n21720), .X(\L2_0/n3447 ) );
  inv_x1_sg U46404 ( .A(n19719), .X(n41953) );
  nand_x1_sg U46405 ( .A(n46519), .B(n19917), .X(n19719) );
  nand_x1_sg U46406 ( .A(n26039), .B(n26040), .X(n16821) );
  nand_x1_sg U46407 ( .A(n26362), .B(n26363), .X(n17642) );
  nand_x1_sg U46408 ( .A(n23404), .B(n41964), .X(n42104) );
  nor_x1_sg U46409 ( .A(reset), .B(n29274), .X(n9274) );
  nand_x1_sg U46410 ( .A(n40220), .B(n39114), .X(n9276) );
  nand_x1_sg U46411 ( .A(n41302), .B(n10094), .X(n42384) );
  nand_x1_sg U46412 ( .A(n25589), .B(n25590), .X(n15182) );
  nand_x1_sg U46413 ( .A(n26123), .B(n41959), .X(n42092) );
  nand_x1_sg U46414 ( .A(n41986), .B(n26419), .X(n17800) );
  nand_x1_sg U46415 ( .A(n26093), .B(n26094), .X(n16818) );
  nand_x1_sg U46416 ( .A(n22801), .B(n22802), .X(n6994) );
  nand_x1_sg U46417 ( .A(n25866), .B(n25867), .X(n16001) );
  nand_x1_sg U46418 ( .A(n26704), .B(n26705), .X(n18460) );
  nand_x1_sg U46419 ( .A(n23637), .B(n23638), .X(n9449) );
  nand_x1_sg U46420 ( .A(n26627), .B(n26628), .X(n19100) );
  nand_x1_sg U46421 ( .A(n26349), .B(n26350), .X(n18279) );
  nand_x1_sg U46422 ( .A(n25789), .B(n25790), .X(n16641) );
  nand_x1_sg U46423 ( .A(n25512), .B(n25513), .X(n15822) );
  nand_x1_sg U46424 ( .A(n25233), .B(n25234), .X(n15003) );
  nand_x1_sg U46425 ( .A(n24954), .B(n24955), .X(n14184) );
  nand_x1_sg U46426 ( .A(n24675), .B(n24676), .X(n13365) );
  nand_x1_sg U46427 ( .A(n24397), .B(n24398), .X(n12546) );
  nand_x1_sg U46428 ( .A(n24118), .B(n24119), .X(n11727) );
  nand_x1_sg U46429 ( .A(n23839), .B(n23840), .X(n10908) );
  nand_x1_sg U46430 ( .A(n23560), .B(n23561), .X(n10089) );
  nand_x1_sg U46431 ( .A(n23001), .B(n23002), .X(n8451) );
  nand_x1_sg U46432 ( .A(n23281), .B(n23282), .X(n9269) );
  nand_x1_sg U46433 ( .A(n22724), .B(n22725), .X(n7633) );
  nand_x1_sg U46434 ( .A(n26640), .B(n26641), .X(n18463) );
  nand_x1_sg U46435 ( .A(n25525), .B(n25526), .X(n15185) );
  nand_x1_sg U46436 ( .A(n25802), .B(n25803), .X(n16004) );
  nand_x1_sg U46437 ( .A(n25246), .B(n25247), .X(n14366) );
  nand_x1_sg U46438 ( .A(n24688), .B(n24689), .X(n12728) );
  nand_x1_sg U46439 ( .A(n24967), .B(n24968), .X(n13547) );
  nand_x1_sg U46440 ( .A(n24410), .B(n24411), .X(n11909) );
  nand_x1_sg U46441 ( .A(n23852), .B(n23853), .X(n10271) );
  nand_x1_sg U46442 ( .A(n24131), .B(n24132), .X(n11090) );
  nand_x1_sg U46443 ( .A(n23573), .B(n23574), .X(n9452) );
  nand_x1_sg U46444 ( .A(n23014), .B(n23015), .X(n7814) );
  nand_x1_sg U46445 ( .A(n23294), .B(n23295), .X(n8632) );
  nand_x1_sg U46446 ( .A(n22737), .B(n22738), .X(n6997) );
  nand_x1_sg U46447 ( .A(n26668), .B(n26669), .X(n18767) );
  nand_x1_sg U46448 ( .A(n26390), .B(n26391), .X(n17946) );
  nand_x1_sg U46449 ( .A(n26063), .B(n26064), .X(n17125) );
  nand_x1_sg U46450 ( .A(n25830), .B(n25831), .X(n16308) );
  nand_x1_sg U46451 ( .A(n25274), .B(n25275), .X(n14670) );
  nand_x1_sg U46452 ( .A(n24995), .B(n24996), .X(n13851) );
  nand_x1_sg U46453 ( .A(n24716), .B(n24717), .X(n13032) );
  nand_x1_sg U46454 ( .A(n24438), .B(n24439), .X(n12213) );
  nand_x1_sg U46455 ( .A(n24159), .B(n24160), .X(n11394) );
  nand_x1_sg U46456 ( .A(n23880), .B(n23881), .X(n10575) );
  nand_x1_sg U46457 ( .A(n23322), .B(n23323), .X(n8936) );
  nand_x1_sg U46458 ( .A(n23601), .B(n23602), .X(n9756) );
  nand_x1_sg U46459 ( .A(n22765), .B(n22766), .X(n7300) );
  nand_x1_sg U46460 ( .A(n41300), .B(n14189), .X(n42382) );
  nand_x1_sg U46461 ( .A(n24752), .B(n24753), .X(n12725) );
  inv_x1_sg U46462 ( .A(n17458), .X(n50525) );
  nand_x1_sg U46463 ( .A(n23916), .B(n23917), .X(n10268) );
  nand_x1_sg U46464 ( .A(n26129), .B(n26130), .X(n17458) );
  nand_x1_sg U46465 ( .A(n46428), .B(n20287), .X(n20113) );
  nand_x1_sg U46466 ( .A(n21347), .B(n46546), .X(n21200) );
  nand_x1_sg U46467 ( .A(n46568), .B(n19723), .X(n19504) );
  nand_x1_sg U46468 ( .A(n21529), .B(n46504), .X(n21341) );
  nand_x1_sg U46469 ( .A(n26472), .B(n50564), .X(n42091) );
  nand_x1_sg U46470 ( .A(n39480), .B(n9275), .X(\L2_0/n3367 ) );
  nand_x1_sg U46471 ( .A(n50850), .B(n26749), .X(n18290) );
  nand_x1_sg U46472 ( .A(n23683), .B(n41965), .X(n42103) );
  nand_x1_sg U46473 ( .A(n23962), .B(n41966), .X(n42102) );
  nand_x1_sg U46474 ( .A(n24241), .B(n41967), .X(n42101) );
  nand_x1_sg U46475 ( .A(n25356), .B(n41963), .X(n42097) );
  nand_x1_sg U46476 ( .A(n24798), .B(n41961), .X(n42099) );
  nand_x1_sg U46477 ( .A(n25077), .B(n41962), .X(n42098) );
  nand_x1_sg U46478 ( .A(n26750), .B(n41958), .X(n42093) );
  nand_x1_sg U46479 ( .A(n24520), .B(n41960), .X(n42100) );
  nand_x1_sg U46480 ( .A(n41128), .B(n26140), .X(n42372) );
  nand_x1_sg U46481 ( .A(n40030), .B(n29272), .X(n42329) );
  nand_x1_sg U46482 ( .A(n25912), .B(n41957), .X(n42094) );
  nand_x1_sg U46483 ( .A(n25031), .B(n25032), .X(n13544) );
  nand_x1_sg U46484 ( .A(n26426), .B(n26427), .X(n17639) );
  nand_x1_sg U46485 ( .A(n39480), .B(n15827), .X(\L2_0/n2727 ) );
  nand_x1_sg U46486 ( .A(n41300), .B(n15008), .X(n42381) );
  nand_x1_sg U46487 ( .A(n24195), .B(n24196), .X(n11087) );
  nand_x1_sg U46488 ( .A(n41301), .B(n11732), .X(\L2_0/n3127 ) );
  nand_x1_sg U46489 ( .A(n24474), .B(n24475), .X(n11906) );
  nand_x1_sg U46490 ( .A(n23078), .B(n23079), .X(n7811) );
  nand_x1_sg U46491 ( .A(n23358), .B(n23359), .X(n8629) );
  nand_x1_sg U46492 ( .A(n25310), .B(n25311), .X(n14363) );
  inv_x1_sg U46493 ( .A(n28542), .X(n41955) );
  inv_x1_sg U46494 ( .A(n20984), .X(n41956) );
  nor_x2_sg U46495 ( .A(n38560), .B(n5398), .X(n28542) );
  nor_x2_sg U46496 ( .A(n41954), .B(n5683), .X(n20984) );
  inv_x1_sg U46497 ( .A(n25913), .X(n41957) );
  inv_x1_sg U46498 ( .A(n26751), .X(n41958) );
  inv_x1_sg U46499 ( .A(n26124), .X(n41959) );
  inv_x1_sg U46500 ( .A(n24521), .X(n41960) );
  inv_x1_sg U46501 ( .A(n24799), .X(n41961) );
  inv_x1_sg U46502 ( .A(n25078), .X(n41962) );
  inv_x1_sg U46503 ( .A(n25357), .X(n41963) );
  inv_x1_sg U46504 ( .A(n23405), .X(n41964) );
  inv_x1_sg U46505 ( .A(n23684), .X(n41965) );
  inv_x1_sg U46506 ( .A(n23963), .X(n41966) );
  inv_x1_sg U46507 ( .A(n24242), .X(n41967) );
  inv_x1_sg U46508 ( .A(n21200), .X(n41968) );
  inv_x1_sg U46509 ( .A(n21341), .X(n41969) );
  inv_x1_sg U46510 ( .A(n20113), .X(n41970) );
  inv_x1_sg U46511 ( .A(n19504), .X(n41971) );
  inv_x1_sg U46512 ( .A(n16641), .X(n41972) );
  inv_x1_sg U46513 ( .A(n18279), .X(n41973) );
  inv_x1_sg U46514 ( .A(n19100), .X(n41974) );
  inv_x1_sg U46515 ( .A(n13365), .X(n41975) );
  inv_x1_sg U46516 ( .A(n14184), .X(n41976) );
  inv_x1_sg U46517 ( .A(n15003), .X(n41977) );
  inv_x1_sg U46518 ( .A(n15822), .X(n41978) );
  inv_x1_sg U46519 ( .A(n10089), .X(n41979) );
  inv_x1_sg U46520 ( .A(n10908), .X(n41980) );
  inv_x1_sg U46521 ( .A(n11727), .X(n41981) );
  inv_x1_sg U46522 ( .A(n12546), .X(n41982) );
  inv_x1_sg U46523 ( .A(n7633), .X(n41983) );
  inv_x1_sg U46524 ( .A(n8451), .X(n41984) );
  inv_x1_sg U46525 ( .A(n9269), .X(n41985) );
  inv_x1_sg U46526 ( .A(n26421), .X(n41986) );
  nand_x1_sg U46527 ( .A(n47295), .B(n23024), .X(n41987) );
  nand_x1_sg U46528 ( .A(n47580), .B(n23304), .X(n41988) );
  nand_x1_sg U46529 ( .A(n47865), .B(n23583), .X(n41989) );
  nand_x1_sg U46530 ( .A(n48150), .B(n23862), .X(n41990) );
  nand_x1_sg U46531 ( .A(n48435), .B(n24141), .X(n41991) );
  nand_x1_sg U46532 ( .A(n48720), .B(n24420), .X(n41992) );
  nand_x1_sg U46533 ( .A(n49006), .B(n24698), .X(n41993) );
  nand_x1_sg U46534 ( .A(n49293), .B(n24977), .X(n41994) );
  nand_x1_sg U46535 ( .A(n49579), .B(n25256), .X(n41995) );
  nand_x1_sg U46536 ( .A(n49865), .B(n25535), .X(n41996) );
  nand_x1_sg U46537 ( .A(n50151), .B(n25812), .X(n41997) );
  nand_x1_sg U46538 ( .A(n51012), .B(n26650), .X(n41998) );
  nand_x1_sg U46539 ( .A(n50725), .B(n26372), .X(n41999) );
  nand_x1_sg U46540 ( .A(n40103), .B(n29273), .X(n42000) );
  inv_x1_sg U46541 ( .A(\reg_yHat[14][17] ), .X(n42001) );
  inv_x1_sg U46542 ( .A(\reg_yHat[12][2] ), .X(n42002) );
  inv_x1_sg U46543 ( .A(\reg_yHat[10][17] ), .X(n42003) );
  inv_x1_sg U46544 ( .A(\reg_yHat[11][17] ), .X(n42004) );
  inv_x1_sg U46545 ( .A(\reg_yHat[12][17] ), .X(n42005) );
  inv_x1_sg U46546 ( .A(\reg_yHat[13][17] ), .X(n42006) );
  inv_x1_sg U46547 ( .A(\reg_yHat[6][17] ), .X(n42007) );
  inv_x1_sg U46548 ( .A(\reg_yHat[7][17] ), .X(n42008) );
  inv_x1_sg U46549 ( .A(\reg_yHat[8][17] ), .X(n42009) );
  inv_x1_sg U46550 ( .A(\reg_yHat[9][17] ), .X(n42010) );
  inv_x1_sg U46551 ( .A(\reg_yHat[2][17] ), .X(n42011) );
  inv_x1_sg U46552 ( .A(\reg_yHat[3][17] ), .X(n42012) );
  inv_x1_sg U46553 ( .A(\reg_yHat[4][17] ), .X(n42013) );
  inv_x1_sg U46554 ( .A(\reg_yHat[5][17] ), .X(n42014) );
  inv_x1_sg U46555 ( .A(\reg_yHat[12][3] ), .X(n42015) );
  inv_x1_sg U46556 ( .A(\reg_yHat[0][17] ), .X(n42016) );
  inv_x1_sg U46557 ( .A(\reg_yHat[1][17] ), .X(n42017) );
  nand_x1_sg U46558 ( .A(n39600), .B(n40649), .X(n42019) );
  inv_x1_sg U46559 ( .A(n24101), .X(n42020) );
  inv_x1_sg U46560 ( .A(reg_num[2]), .X(n42021) );
  inv_x1_sg U46561 ( .A(state[1]), .X(n42022) );
  inv_x1_sg U46562 ( .A(n21013), .X(n42023) );
  inv_x1_sg U46563 ( .A(n19583), .X(n42024) );
  inv_x1_sg U46564 ( .A(\reg_yHat[13][6] ), .X(n42025) );
  inv_x1_sg U46565 ( .A(\reg_yHat[14][6] ), .X(n42026) );
  inv_x1_sg U46566 ( .A(\reg_yHat[10][6] ), .X(n42027) );
  inv_x1_sg U46567 ( .A(\reg_yHat[11][6] ), .X(n42028) );
  inv_x1_sg U46568 ( .A(\reg_yHat[12][6] ), .X(n42029) );
  inv_x1_sg U46569 ( .A(\reg_yHat[12][18] ), .X(n42030) );
  inv_x1_sg U46570 ( .A(\reg_yHat[6][6] ), .X(n42031) );
  inv_x1_sg U46571 ( .A(\reg_yHat[7][6] ), .X(n42032) );
  inv_x1_sg U46572 ( .A(\reg_yHat[8][6] ), .X(n42033) );
  inv_x1_sg U46573 ( .A(\reg_yHat[9][6] ), .X(n42034) );
  inv_x1_sg U46574 ( .A(\reg_yHat[2][6] ), .X(n42035) );
  inv_x1_sg U46575 ( .A(\reg_yHat[3][6] ), .X(n42036) );
  inv_x1_sg U46576 ( .A(\reg_yHat[4][6] ), .X(n42037) );
  inv_x1_sg U46577 ( .A(\reg_yHat[5][6] ), .X(n42038) );
  inv_x1_sg U46578 ( .A(\reg_yHat[0][6] ), .X(n42039) );
  inv_x1_sg U46579 ( .A(\reg_yHat[0][18] ), .X(n42040) );
  inv_x1_sg U46580 ( .A(\reg_yHat[1][6] ), .X(n42041) );
  inv_x1_sg U46581 ( .A(n26177), .X(n42043) );
  nand_x1_sg U46582 ( .A(n42047), .B(n26471), .X(n42044) );
  nand_x1_sg U46583 ( .A(n7008), .B(n7009), .X(n42045) );
  inv_x1_sg U46584 ( .A(n22843), .X(n42046) );
  inv_x1_sg U46585 ( .A(n26468), .X(n42047) );
  inv_x1_sg U46586 ( .A(n25908), .X(n42048) );
  inv_x1_sg U46587 ( .A(n25631), .X(n42049) );
  inv_x1_sg U46588 ( .A(n25352), .X(n42050) );
  inv_x1_sg U46589 ( .A(n25073), .X(n42051) );
  inv_x1_sg U46590 ( .A(n24794), .X(n42052) );
  inv_x1_sg U46591 ( .A(n24516), .X(n42053) );
  inv_x1_sg U46592 ( .A(n24237), .X(n42054) );
  inv_x1_sg U46593 ( .A(n23958), .X(n42055) );
  inv_x1_sg U46594 ( .A(n23679), .X(n42056) );
  inv_x1_sg U46595 ( .A(n23400), .X(n42057) );
  nand_x1_sg U46596 ( .A(n39081), .B(n29271), .X(n42058) );
  inv_x1_sg U46597 ( .A(n25595), .X(n42060) );
  nand_x1_sg U46598 ( .A(n19096), .B(n18656), .X(n42061) );
  nand_x1_sg U46599 ( .A(n18275), .B(n17835), .X(n42062) );
  nand_x1_sg U46600 ( .A(n16637), .B(n16197), .X(n42063) );
  nand_x1_sg U46601 ( .A(n14999), .B(n14559), .X(n42064) );
  nand_x1_sg U46602 ( .A(n14180), .B(n13740), .X(n42065) );
  nand_x1_sg U46603 ( .A(n13361), .B(n12921), .X(n42066) );
  nand_x1_sg U46604 ( .A(n12542), .B(n12102), .X(n42067) );
  nand_x1_sg U46605 ( .A(n11723), .B(n11283), .X(n42068) );
  nand_x1_sg U46606 ( .A(n10904), .B(n10464), .X(n42069) );
  nand_x1_sg U46607 ( .A(n10085), .B(n9645), .X(n42070) );
  nand_x1_sg U46608 ( .A(n9265), .B(n8825), .X(n42071) );
  nand_x2_sg U46609 ( .A(n6558), .B(n6559), .X(n6557) );
  nand_x2_sg U46610 ( .A(n6469), .B(n6470), .X(n6468) );
  nand_x2_sg U46611 ( .A(n6335), .B(n6336), .X(n6334) );
  nand_x1_sg U46612 ( .A(n15818), .B(n15378), .X(n42072) );
  nand_x1_sg U46613 ( .A(n8447), .B(n8007), .X(n42073) );
  nand_x1_sg U46614 ( .A(n7629), .B(n7188), .X(n42074) );
  inv_x2_sg U46615 ( .A(n21600), .X(n42075) );
  inv_x2_sg U46616 ( .A(n21624), .X(n42077) );
  inv_x2_sg U46617 ( .A(n21636), .X(n42078) );
  inv_x2_sg U46618 ( .A(n21648), .X(n42079) );
  inv_x2_sg U46619 ( .A(n21660), .X(n42080) );
  inv_x2_sg U46620 ( .A(n29151), .X(n42082) );
  inv_x2_sg U46621 ( .A(n29163), .X(n42083) );
  inv_x2_sg U46622 ( .A(n29175), .X(n42084) );
  nand_x2_sg U46623 ( .A(n6695), .B(n6696), .X(n6694) );
  nand_x2_sg U46624 ( .A(n6647), .B(n6648), .X(n6646) );
  nand_x2_sg U46625 ( .A(n6513), .B(n6514), .X(n6512) );
  nand_x2_sg U46626 ( .A(n6424), .B(n6425), .X(n6423) );
  nand_x2_sg U46627 ( .A(n6291), .B(n6292), .X(n6290) );
  nand_x2_sg U46628 ( .A(n6246), .B(n6247), .X(n6245) );
  nand_x2_sg U46629 ( .A(n6153), .B(n6154), .X(n6152) );
  nand_x1_sg U46630 ( .A(n19584), .B(n46390), .X(n42087) );
  nand_x1_sg U46631 ( .A(n17454), .B(n17013), .X(n42088) );
  nand_x1_sg U46632 ( .A(n26045), .B(n26046), .X(n17299) );
  nand_x1_sg U46633 ( .A(n49143), .B(n25058), .X(n13634) );
  nand_x1_sg U46634 ( .A(n42090), .B(n23105), .X(n42089) );
  inv_x1_sg U46635 ( .A(n23107), .X(n42090) );
  nand_x1_sg U46636 ( .A(n25635), .B(n42096), .X(n42095) );
  inv_x1_sg U46637 ( .A(n25636), .X(n42096) );
  inv_x1_sg U46638 ( .A(n23125), .X(n42106) );
  inv_x1_sg U46639 ( .A(n24380), .X(n42119) );
  inv_x1_sg U46640 ( .A(n26100), .X(n42120) );
  nand_x1_sg U46641 ( .A(n50862), .B(n26731), .X(n18550) );
  inv_x1_sg U46642 ( .A(n26455), .X(n42121) );
  nand_x1_sg U46643 ( .A(n42121), .B(n26453), .X(n17729) );
  nand_x1_sg U46644 ( .A(n50001), .B(n25893), .X(n16091) );
  nand_x1_sg U46645 ( .A(n42123), .B(n25616), .X(n42122) );
  inv_x1_sg U46646 ( .A(n25618), .X(n42123) );
  nand_x1_sg U46647 ( .A(n49429), .B(n25337), .X(n42124) );
  nand_x1_sg U46648 ( .A(n48856), .B(n24779), .X(n12815) );
  inv_x1_sg U46649 ( .A(n24503), .X(n42125) );
  nand_x1_sg U46650 ( .A(n42125), .B(n24501), .X(n11996) );
  nand_x1_sg U46651 ( .A(n42127), .B(n24222), .X(n42126) );
  inv_x1_sg U46652 ( .A(n24224), .X(n42127) );
  inv_x1_sg U46653 ( .A(n23945), .X(n42128) );
  nand_x1_sg U46654 ( .A(n42128), .B(n23943), .X(n10358) );
  inv_x1_sg U46655 ( .A(n23666), .X(n42129) );
  nand_x1_sg U46656 ( .A(n42129), .B(n23664), .X(n9539) );
  nand_x1_sg U46657 ( .A(n42131), .B(n23385), .X(n42130) );
  inv_x1_sg U46658 ( .A(n23387), .X(n42131) );
  nand_x2_sg U46659 ( .A(n5683), .B(n41954), .X(n42132) );
  nand_x2_sg U46660 ( .A(n5683), .B(n41954), .X(n20983) );
  nand_x2_sg U46661 ( .A(n5398), .B(n38560), .X(n42133) );
  nand_x2_sg U46662 ( .A(n5398), .B(n38560), .X(n28541) );
  nand_x2_sg U46663 ( .A(n6786), .B(n6787), .X(n6785) );
  nand_x2_sg U46664 ( .A(n6602), .B(n6603), .X(n6601) );
  nand_x2_sg U46665 ( .A(n6380), .B(n6381), .X(n6379) );
  nand_x2_sg U46666 ( .A(n6199), .B(n6200), .X(n6198) );
  nand_x2_sg U46667 ( .A(n6108), .B(n6109), .X(n6107) );
  nand_x2_sg U46668 ( .A(n6060), .B(n6061), .X(n6059) );
  nand_x2_sg U46669 ( .A(n5956), .B(n5957), .X(n5955) );
  inv_x1_sg U46670 ( .A(n26710), .X(n42134) );
  inv_x1_sg U46671 ( .A(n26432), .X(n42135) );
  inv_x1_sg U46672 ( .A(n25872), .X(n42136) );
  inv_x1_sg U46673 ( .A(n25316), .X(n42137) );
  inv_x1_sg U46674 ( .A(n25037), .X(n42138) );
  inv_x1_sg U46675 ( .A(n24758), .X(n42139) );
  inv_x1_sg U46676 ( .A(n24480), .X(n42140) );
  inv_x1_sg U46677 ( .A(n24201), .X(n42141) );
  inv_x1_sg U46678 ( .A(n23922), .X(n42142) );
  inv_x1_sg U46679 ( .A(n23643), .X(n42143) );
  inv_x1_sg U46680 ( .A(n23364), .X(n42144) );
  inv_x1_sg U46681 ( .A(n23084), .X(n42145) );
  inv_x1_sg U46682 ( .A(n22807), .X(n42146) );
  nand_x1_sg U46683 ( .A(n26038), .B(n26010), .X(n42147) );
  inv_x1_sg U46684 ( .A(n20691), .X(n42148) );
  inv_x1_sg U46685 ( .A(n20058), .X(n42149) );
  inv_x1_sg U46686 ( .A(n20705), .X(n42150) );
  inv_x1_sg U46687 ( .A(n20712), .X(n42151) );
  inv_x1_sg U46688 ( .A(n20726), .X(n42152) );
  inv_x1_sg U46689 ( .A(n28180), .X(n42153) );
  inv_x1_sg U46690 ( .A(n28081), .X(n42154) );
  inv_x1_sg U46691 ( .A(n27919), .X(n42155) );
  inv_x1_sg U46692 ( .A(n27742), .X(n42156) );
  inv_x1_sg U46693 ( .A(n27548), .X(n42157) );
  inv_x1_sg U46694 ( .A(n27335), .X(n42158) );
  inv_x1_sg U46695 ( .A(n27970), .X(n42159) );
  nor_x1_sg U46696 ( .A(n28809), .B(n28810), .X(n22583) );
  nand_x1_sg U46697 ( .A(n40221), .B(n42042), .X(n9275) );
  inv_x1_sg U46698 ( .A(n18286), .X(n42162) );
  nand_x1_sg U46699 ( .A(n42165), .B(n26697), .X(n42164) );
  inv_x1_sg U46700 ( .A(n26699), .X(n42165) );
  nand_x1_sg U46701 ( .A(n42167), .B(n25859), .X(n42166) );
  inv_x1_sg U46702 ( .A(n25861), .X(n42167) );
  nand_x1_sg U46703 ( .A(n49754), .B(n25582), .X(n42168) );
  nand_x1_sg U46704 ( .A(n42170), .B(n25303), .X(n42169) );
  inv_x1_sg U46705 ( .A(n25305), .X(n42170) );
  nand_x1_sg U46706 ( .A(n42172), .B(n25024), .X(n42171) );
  inv_x1_sg U46707 ( .A(n25026), .X(n42172) );
  nand_x1_sg U46708 ( .A(n42174), .B(n24745), .X(n42173) );
  inv_x1_sg U46709 ( .A(n24747), .X(n42174) );
  nand_x1_sg U46710 ( .A(n42176), .B(n24467), .X(n42175) );
  inv_x1_sg U46711 ( .A(n24469), .X(n42176) );
  nand_x1_sg U46712 ( .A(n42178), .B(n24188), .X(n42177) );
  inv_x1_sg U46713 ( .A(n24190), .X(n42178) );
  nand_x1_sg U46714 ( .A(n42180), .B(n23909), .X(n42179) );
  inv_x1_sg U46715 ( .A(n23911), .X(n42180) );
  nand_x1_sg U46716 ( .A(n42182), .B(n23630), .X(n42181) );
  inv_x1_sg U46717 ( .A(n23632), .X(n42182) );
  nand_x1_sg U46718 ( .A(n42184), .B(n23351), .X(n42183) );
  inv_x1_sg U46719 ( .A(n23353), .X(n42184) );
  nand_x1_sg U46720 ( .A(n42186), .B(n23071), .X(n42185) );
  inv_x1_sg U46721 ( .A(n23073), .X(n42186) );
  nand_x1_sg U46722 ( .A(n26412), .B(n26413), .X(n17863) );
  nand_x1_sg U46723 ( .A(n26081), .B(n26082), .X(n17041) );
  nand_x1_sg U46724 ( .A(n22819), .B(n22820), .X(n7111) );
  nand_x1_sg U46725 ( .A(n50291), .B(n26105), .X(n16936) );
  nand_x1_sg U46726 ( .A(n42046), .B(n22851), .X(n6831) );
  nand_x1_sg U46727 ( .A(n42043), .B(n26128), .X(n16655) );
  nand_x1_sg U46728 ( .A(n42075), .B(n21599), .X(n42187) );
  nand_x4_sg U46729 ( .A(out_L2[2]), .B(n42107), .X(n21599) );
  nand_x1_sg U46730 ( .A(n42076), .B(n21611), .X(n42188) );
  nand_x4_sg U46731 ( .A(out_L2[4]), .B(n42108), .X(n21611) );
  nand_x1_sg U46732 ( .A(n42077), .B(n21623), .X(n42189) );
  nand_x4_sg U46733 ( .A(out_L2[6]), .B(n42109), .X(n21623) );
  nand_x1_sg U46734 ( .A(n42078), .B(n21635), .X(n42190) );
  nand_x4_sg U46735 ( .A(out_L2[8]), .B(n42110), .X(n21635) );
  nand_x1_sg U46736 ( .A(n42079), .B(n21647), .X(n42191) );
  nand_x4_sg U46737 ( .A(out_L2[10]), .B(n42111), .X(n21647) );
  nand_x1_sg U46738 ( .A(n42080), .B(n21659), .X(n42192) );
  nand_x4_sg U46739 ( .A(out_L2[12]), .B(n42112), .X(n21659) );
  nand_x1_sg U46740 ( .A(n42081), .B(n21357), .X(n42193) );
  nand_x4_sg U46741 ( .A(out_L2[17]), .B(n42113), .X(n21357) );
  nand_x1_sg U46742 ( .A(n42082), .B(n29150), .X(n42194) );
  nand_x4_sg U46743 ( .A(out_L1[2]), .B(n42114), .X(n29150) );
  nand_x1_sg U46744 ( .A(n42083), .B(n29162), .X(n42195) );
  nand_x4_sg U46745 ( .A(out_L1[4]), .B(n42115), .X(n29162) );
  nand_x1_sg U46746 ( .A(n42084), .B(n29174), .X(n42196) );
  nand_x4_sg U46747 ( .A(out_L1[6]), .B(n42116), .X(n29174) );
  nand_x1_sg U46748 ( .A(n42085), .B(n29186), .X(n42197) );
  nand_x4_sg U46749 ( .A(out_L1[8]), .B(n42117), .X(n29186) );
  nand_x1_sg U46750 ( .A(n42086), .B(n28921), .X(n42198) );
  nand_x4_sg U46751 ( .A(out_L1[17]), .B(n42118), .X(n28921) );
  inv_x1_sg U46752 ( .A(n20677), .X(n42199) );
  inv_x1_sg U46753 ( .A(n20037), .X(n42200) );
  inv_x1_sg U46754 ( .A(n20684), .X(n42201) );
  inv_x1_sg U46755 ( .A(n20044), .X(n42202) );
  inv_x1_sg U46756 ( .A(n20051), .X(n42203) );
  inv_x1_sg U46757 ( .A(n20698), .X(n42204) );
  inv_x1_sg U46758 ( .A(n20065), .X(n42205) );
  inv_x1_sg U46759 ( .A(n20072), .X(n42206) );
  inv_x1_sg U46760 ( .A(n20719), .X(n42207) );
  inv_x1_sg U46761 ( .A(n20079), .X(n42208) );
  inv_x1_sg U46762 ( .A(n20086), .X(n42209) );
  inv_x1_sg U46763 ( .A(n20733), .X(n42210) );
  inv_x1_sg U46764 ( .A(n20093), .X(n42211) );
  inv_x1_sg U46765 ( .A(n20740), .X(n42212) );
  inv_x1_sg U46766 ( .A(n20100), .X(n42213) );
  inv_x1_sg U46767 ( .A(n20747), .X(n42214) );
  inv_x1_sg U46768 ( .A(\reg_y[0][2] ), .X(n42215) );
  inv_x1_sg U46769 ( .A(n19268), .X(n42216) );
  inv_x1_sg U46770 ( .A(n19233), .X(n42217) );
  inv_x1_sg U46771 ( .A(n19240), .X(n42218) );
  inv_x1_sg U46772 ( .A(n19254), .X(n42219) );
  inv_x1_sg U46773 ( .A(n19261), .X(n42220) );
  inv_x1_sg U46774 ( .A(n19275), .X(n42221) );
  inv_x1_sg U46775 ( .A(n19282), .X(n42222) );
  inv_x1_sg U46776 ( .A(n19289), .X(n42223) );
  inv_x1_sg U46777 ( .A(n19296), .X(n42224) );
  inv_x1_sg U46778 ( .A(n19402), .X(n42225) );
  inv_x1_sg U46779 ( .A(n19912), .X(n42226) );
  inv_x1_sg U46780 ( .A(n20208), .X(n42227) );
  inv_x1_sg U46781 ( .A(n27105), .X(n42228) );
  inv_x1_sg U46782 ( .A(n20851), .X(n42229) );
  nor_x1_sg U46783 ( .A(n19244), .B(n19245), .X(n42230) );
  nor_x1_sg U46784 ( .A(n20723), .B(n20724), .X(n42231) );
  nor_x1_sg U46785 ( .A(n20709), .B(n20710), .X(n42232) );
  nor_x1_sg U46786 ( .A(n20688), .B(n20689), .X(n42233) );
  nor_x1_sg U46787 ( .A(n20702), .B(n20703), .X(n42234) );
  nor_x1_sg U46788 ( .A(n19475), .B(n19476), .X(n6226) );
  nor_x1_sg U46789 ( .A(n23264), .B(n51137), .X(n20569) );
  nor_x1_sg U46790 ( .A(n42042), .B(n41398), .X(n20567) );
  nor_x1_sg U46791 ( .A(n41632), .B(n51140), .X(n19124) );
  nand_x1_sg U46792 ( .A(n42048), .B(n25911), .X(n15831) );
  nand_x1_sg U46793 ( .A(n42049), .B(n25634), .X(n15012) );
  nand_x1_sg U46794 ( .A(n42050), .B(n25355), .X(n14193) );
  nand_x1_sg U46795 ( .A(n42051), .B(n25076), .X(n13374) );
  nand_x1_sg U46796 ( .A(n42052), .B(n24797), .X(n12555) );
  nand_x1_sg U46797 ( .A(n42053), .B(n24519), .X(n11736) );
  nand_x1_sg U46798 ( .A(n42054), .B(n24240), .X(n10917) );
  nand_x1_sg U46799 ( .A(n42055), .B(n23961), .X(n10098) );
  nand_x1_sg U46800 ( .A(n42056), .B(n23682), .X(n9279) );
  nand_x1_sg U46801 ( .A(n42057), .B(n23403), .X(n8459) );
  nand_x1_sg U46802 ( .A(n47134), .B(n23123), .X(n7641) );
  nand_x2_sg U46803 ( .A(n6735), .B(n6736), .X(n6734) );
  nand_x2_sg U46804 ( .A(n6011), .B(n6012), .X(n6010) );
  nand_x2_sg U46805 ( .A(n19109), .B(n19110), .X(n19108) );
  nand_x8_sg U46806 ( .A(n45811), .B(n38597), .X(n6757) );
  nand_x1_sg U46807 ( .A(n42132), .B(n41956), .X(n42237) );
  nand_x1_sg U46808 ( .A(n42133), .B(n41955), .X(n42238) );
  nand_x1_sg U46809 ( .A(n18821), .B(n18789), .X(n42239) );
  nand_x1_sg U46810 ( .A(n18000), .B(n17968), .X(n42240) );
  nand_x1_sg U46811 ( .A(n17179), .B(n17147), .X(n42241) );
  nand_x1_sg U46812 ( .A(n17093), .B(n17068), .X(n42242) );
  nand_x1_sg U46813 ( .A(n16362), .B(n16330), .X(n42243) );
  nand_x1_sg U46814 ( .A(n15543), .B(n15511), .X(n42244) );
  nand_x1_sg U46815 ( .A(n14724), .B(n14692), .X(n42245) );
  nand_x1_sg U46816 ( .A(n13905), .B(n13873), .X(n42246) );
  nand_x1_sg U46817 ( .A(n13086), .B(n13054), .X(n42247) );
  nand_x1_sg U46818 ( .A(n12267), .B(n12235), .X(n42248) );
  nand_x1_sg U46819 ( .A(n11448), .B(n11416), .X(n42249) );
  nand_x1_sg U46820 ( .A(n10629), .B(n10597), .X(n42250) );
  nand_x1_sg U46821 ( .A(n9810), .B(n9778), .X(n42251) );
  nand_x1_sg U46822 ( .A(n8990), .B(n8958), .X(n42252) );
  nand_x1_sg U46823 ( .A(n8172), .B(n8140), .X(n42253) );
  nand_x1_sg U46824 ( .A(n7354), .B(n7322), .X(n42254) );
  nand_x1_sg U46825 ( .A(n7268), .B(n7243), .X(n42255) );
  inv_x1_sg U46826 ( .A(n20754), .X(n42256) );
  inv_x1_sg U46827 ( .A(n20761), .X(n42257) );
  inv_x1_sg U46828 ( .A(n6127), .X(n42258) );
  inv_x1_sg U46829 ( .A(n20768), .X(n42259) );
  inv_x1_sg U46830 ( .A(n20999), .X(n42260) );
  inv_x1_sg U46831 ( .A(n19247), .X(n42261) );
  inv_x1_sg U46832 ( .A(n19712), .X(n42262) );
  nand_x2_sg U46833 ( .A(out_L2[14]), .B(n38123), .X(n21671) );
  nand_x2_sg U46834 ( .A(out_L2[16]), .B(n38125), .X(n21539) );
  nand_x2_sg U46835 ( .A(out_L1[10]), .B(n38121), .X(n29198) );
  nand_x2_sg U46836 ( .A(out_L1[12]), .B(n38122), .X(n29210) );
  nand_x2_sg U46837 ( .A(out_L1[14]), .B(n38124), .X(n29222) );
  nand_x2_sg U46838 ( .A(out_L1[16]), .B(n38126), .X(n29090) );
  nor_x1_sg U46839 ( .A(n45966), .B(n21451), .X(n42263) );
  nor_x1_sg U46840 ( .A(n46011), .B(n21457), .X(n42264) );
  nor_x1_sg U46841 ( .A(n46057), .B(n21464), .X(n42265) );
  nor_x1_sg U46842 ( .A(n46102), .B(n21470), .X(n42266) );
  nor_x1_sg U46843 ( .A(n46148), .B(n21477), .X(n42267) );
  nor_x1_sg U46844 ( .A(n19265), .B(n19266), .X(n42268) );
  nor_x1_sg U46845 ( .A(n46193), .B(n21483), .X(n42269) );
  nor_x1_sg U46846 ( .A(n46239), .B(n21490), .X(n42270) );
  nor_x1_sg U46847 ( .A(n46284), .B(n21496), .X(n42271) );
  nor_x1_sg U46848 ( .A(n46330), .B(n21503), .X(n42272) );
  nor_x1_sg U46849 ( .A(n46371), .B(n21509), .X(n42273) );
  nor_x1_sg U46850 ( .A(n46419), .B(n21516), .X(n42274) );
  nor_x1_sg U46851 ( .A(n46466), .B(n21522), .X(n42275) );
  nor_x1_sg U46852 ( .A(n19237), .B(n19238), .X(n42276) );
  nor_x1_sg U46853 ( .A(n19251), .B(n19252), .X(n42277) );
  nor_x1_sg U46854 ( .A(n19258), .B(n19259), .X(n42278) );
  nor_x1_sg U46855 ( .A(n19272), .B(n19273), .X(n42279) );
  nor_x1_sg U46856 ( .A(n19279), .B(n19280), .X(n42280) );
  nor_x1_sg U46857 ( .A(n19286), .B(n19287), .X(n42281) );
  nor_x1_sg U46858 ( .A(n19293), .B(n19294), .X(n42282) );
  nor_x1_sg U46859 ( .A(n46556), .B(n19934), .X(n42283) );
  nor_x1_sg U46860 ( .A(n20744), .B(n20745), .X(n42284) );
  nor_x1_sg U46861 ( .A(n45927), .B(n19846), .X(n42285) );
  nor_x1_sg U46862 ( .A(n20069), .B(n20070), .X(n42286) );
  nor_x1_sg U46863 ( .A(n20041), .B(n20042), .X(n42287) );
  nor_x1_sg U46864 ( .A(n20048), .B(n20049), .X(n42288) );
  nor_x1_sg U46865 ( .A(n20055), .B(n20056), .X(n42289) );
  nor_x1_sg U46866 ( .A(n20062), .B(n20063), .X(n42290) );
  nor_x1_sg U46867 ( .A(n20076), .B(n20077), .X(n42291) );
  nor_x1_sg U46868 ( .A(n20083), .B(n20084), .X(n42292) );
  nor_x1_sg U46869 ( .A(n20090), .B(n20091), .X(n42293) );
  nor_x1_sg U46870 ( .A(n20097), .B(n20098), .X(n42294) );
  nor_x1_sg U46871 ( .A(n21344), .B(n21345), .X(n42295) );
  nor_x1_sg U46872 ( .A(n20737), .B(n20738), .X(n42296) );
  nor_x1_sg U46873 ( .A(n20730), .B(n20731), .X(n42297) );
  nor_x1_sg U46874 ( .A(n45924), .B(n20503), .X(n42298) );
  nor_x1_sg U46875 ( .A(n20716), .B(n20717), .X(n42299) );
  nor_x1_sg U46876 ( .A(n20681), .B(n20682), .X(n42300) );
  nor_x1_sg U46877 ( .A(n20695), .B(n20696), .X(n42301) );
  nor_x1_sg U46878 ( .A(n45921), .B(n21272), .X(n42302) );
  nor_x1_sg U46879 ( .A(n19230), .B(n19231), .X(n6664) );
  nor_x1_sg U46880 ( .A(n19501), .B(n19502), .X(n6038) );
  nor_x1_sg U46881 ( .A(n20539), .B(n20540), .X(n6374) );
  nor_x1_sg U46882 ( .A(n20529), .B(n20530), .X(n6463) );
  nor_x1_sg U46883 ( .A(n20514), .B(n20515), .X(n6596) );
  nor_x1_sg U46884 ( .A(n20524), .B(n20525), .X(n6507) );
  nand_x1_sg U46885 ( .A(n26057), .B(n26058), .X(n16815) );
  nand_x1_sg U46886 ( .A(n42326), .B(n22828), .X(n42325) );
  inv_x1_sg U46887 ( .A(n22830), .X(n42326) );
  nand_x1_sg U46888 ( .A(n26690), .B(n26691), .X(n18684) );
  nand_x1_sg U46889 ( .A(n25852), .B(n25853), .X(n16225) );
  nand_x1_sg U46890 ( .A(n25575), .B(n25576), .X(n15406) );
  nand_x1_sg U46891 ( .A(n25296), .B(n25297), .X(n14587) );
  nand_x1_sg U46892 ( .A(n25017), .B(n25018), .X(n13768) );
  nand_x1_sg U46893 ( .A(n24738), .B(n24739), .X(n12949) );
  nand_x1_sg U46894 ( .A(n24460), .B(n24461), .X(n12130) );
  nand_x1_sg U46895 ( .A(n24181), .B(n24182), .X(n11311) );
  nand_x1_sg U46896 ( .A(n23902), .B(n23903), .X(n10492) );
  nand_x1_sg U46897 ( .A(n23623), .B(n23624), .X(n9673) );
  nand_x1_sg U46898 ( .A(n23344), .B(n23345), .X(n8853) );
  nand_x1_sg U46899 ( .A(n23064), .B(n23065), .X(n8035) );
  nand_x1_sg U46900 ( .A(n40104), .B(n25494), .X(n42327) );
  nand_x1_sg U46901 ( .A(n26117), .B(n50281), .X(n16658) );
  inv_x1_sg U46902 ( .A(n42059), .X(n42328) );
  nor_x1_sg U46903 ( .A(n19780), .B(n19781), .X(n19779) );
  nor_x1_sg U46904 ( .A(n19782), .B(n5477), .X(n19781) );
  nor_x1_sg U46905 ( .A(n19785), .B(n5478), .X(n19784) );
  nor_x1_sg U46906 ( .A(n19787), .B(n19788), .X(n19786) );
  nor_x1_sg U46907 ( .A(n19789), .B(n5479), .X(n19788) );
  nor_x1_sg U46908 ( .A(n19791), .B(n19792), .X(n19790) );
  inv_x1_sg U46909 ( .A(n19793), .X(n46392) );
  nor_x1_sg U46910 ( .A(n20609), .B(n20610), .X(n20608) );
  nor_x1_sg U46911 ( .A(n20611), .B(n5575), .X(n20610) );
  nor_x1_sg U46912 ( .A(n19618), .B(n19619), .X(n19617) );
  nor_x1_sg U46913 ( .A(n19620), .B(n5472), .X(n19619) );
  nor_x1_sg U46914 ( .A(n7572), .B(n7573), .X(n7571) );
  nand_x1_sg U46915 ( .A(n7598), .B(n7599), .X(n7541) );
  nand_x1_sg U46916 ( .A(n7627), .B(n47103), .X(n7616) );
  nand_x1_sg U46917 ( .A(n7533), .B(n7534), .X(n7531) );
  nor_x1_sg U46918 ( .A(n8390), .B(n8391), .X(n8389) );
  nand_x1_sg U46919 ( .A(n8416), .B(n8417), .X(n8359) );
  nand_x1_sg U46920 ( .A(n8445), .B(n47389), .X(n8434) );
  nand_x1_sg U46921 ( .A(n8351), .B(n8352), .X(n8349) );
  nor_x1_sg U46922 ( .A(n9208), .B(n9209), .X(n9207) );
  nand_x1_sg U46923 ( .A(n9234), .B(n9235), .X(n9177) );
  nand_x1_sg U46924 ( .A(n9263), .B(n47674), .X(n9252) );
  nand_x1_sg U46925 ( .A(n9169), .B(n9170), .X(n9167) );
  nor_x1_sg U46926 ( .A(n10028), .B(n10029), .X(n10027) );
  nand_x1_sg U46927 ( .A(n10054), .B(n10055), .X(n9997) );
  nand_x1_sg U46928 ( .A(n10083), .B(n47959), .X(n10072) );
  nand_x1_sg U46929 ( .A(n9989), .B(n9990), .X(n9987) );
  nor_x1_sg U46930 ( .A(n10847), .B(n10848), .X(n10846) );
  nand_x1_sg U46931 ( .A(n10873), .B(n10874), .X(n10816) );
  nand_x1_sg U46932 ( .A(n10902), .B(n48244), .X(n10891) );
  nand_x1_sg U46933 ( .A(n10808), .B(n10809), .X(n10806) );
  nor_x1_sg U46934 ( .A(n11666), .B(n11667), .X(n11665) );
  nand_x1_sg U46935 ( .A(n11692), .B(n11693), .X(n11635) );
  nand_x1_sg U46936 ( .A(n11721), .B(n48529), .X(n11710) );
  nand_x1_sg U46937 ( .A(n11627), .B(n11628), .X(n11625) );
  nor_x1_sg U46938 ( .A(n12485), .B(n12486), .X(n12484) );
  nand_x1_sg U46939 ( .A(n12511), .B(n12512), .X(n12454) );
  nand_x1_sg U46940 ( .A(n12540), .B(n48814), .X(n12529) );
  nand_x1_sg U46941 ( .A(n12446), .B(n12447), .X(n12444) );
  nor_x1_sg U46942 ( .A(n13304), .B(n13305), .X(n13303) );
  nand_x1_sg U46943 ( .A(n13330), .B(n13331), .X(n13273) );
  nand_x1_sg U46944 ( .A(n13359), .B(n49101), .X(n13348) );
  nand_x1_sg U46945 ( .A(n13265), .B(n13266), .X(n13263) );
  nor_x1_sg U46946 ( .A(n14123), .B(n14124), .X(n14122) );
  nand_x1_sg U46947 ( .A(n14149), .B(n14150), .X(n14092) );
  nand_x1_sg U46948 ( .A(n14178), .B(n49387), .X(n14167) );
  nand_x1_sg U46949 ( .A(n14084), .B(n14085), .X(n14082) );
  nor_x1_sg U46950 ( .A(n14942), .B(n14943), .X(n14941) );
  nand_x1_sg U46951 ( .A(n14968), .B(n14969), .X(n14911) );
  nand_x1_sg U46952 ( .A(n14997), .B(n49673), .X(n14986) );
  nand_x1_sg U46953 ( .A(n14903), .B(n14904), .X(n14901) );
  nor_x1_sg U46954 ( .A(n15761), .B(n15762), .X(n15760) );
  nand_x1_sg U46955 ( .A(n15787), .B(n15788), .X(n15730) );
  nand_x1_sg U46956 ( .A(n15816), .B(n49959), .X(n15805) );
  nand_x1_sg U46957 ( .A(n15722), .B(n15723), .X(n15720) );
  nor_x1_sg U46958 ( .A(n16580), .B(n16581), .X(n16579) );
  nand_x1_sg U46959 ( .A(n16606), .B(n16607), .X(n16549) );
  nand_x1_sg U46960 ( .A(n16635), .B(n50245), .X(n16624) );
  nand_x1_sg U46961 ( .A(n16541), .B(n16542), .X(n16539) );
  nor_x1_sg U46962 ( .A(n17397), .B(n17398), .X(n17396) );
  nand_x1_sg U46963 ( .A(n17423), .B(n17424), .X(n17366) );
  nand_x1_sg U46964 ( .A(n17452), .B(n50530), .X(n17441) );
  nand_x1_sg U46965 ( .A(n17358), .B(n17359), .X(n17356) );
  nor_x1_sg U46966 ( .A(n18218), .B(n18219), .X(n18217) );
  nand_x1_sg U46967 ( .A(n18244), .B(n18245), .X(n18187) );
  nand_x1_sg U46968 ( .A(n18273), .B(n50819), .X(n18262) );
  nand_x1_sg U46969 ( .A(n18179), .B(n18180), .X(n18177) );
  nor_x1_sg U46970 ( .A(n19039), .B(n19040), .X(n19038) );
  nand_x1_sg U46971 ( .A(n19065), .B(n19066), .X(n19008) );
  nand_x1_sg U46972 ( .A(n19094), .B(n51106), .X(n19083) );
  nand_x1_sg U46973 ( .A(n19000), .B(n19001), .X(n18998) );
  nor_x1_sg U46974 ( .A(n19770), .B(n46564), .X(n19557) );
  inv_x1_sg U46975 ( .A(n19771), .X(n46564) );
  nor_x1_sg U46976 ( .A(n19764), .B(n19765), .X(n19550) );
  nor_x1_sg U46977 ( .A(n19766), .B(n5514), .X(n19765) );
  nor_x1_sg U46978 ( .A(n19752), .B(n19753), .X(n19536) );
  nor_x1_sg U46979 ( .A(n19754), .B(n5552), .X(n19753) );
  nor_x1_sg U46980 ( .A(n19343), .B(n19344), .X(n19328) );
  inv_x1_sg U46981 ( .A(n19345), .X(n46525) );
  nor_x1_sg U46982 ( .A(n19776), .B(n19777), .X(n19564) );
  nor_x1_sg U46983 ( .A(n19778), .B(n5476), .X(n19777) );
  nor_x1_sg U46984 ( .A(n19573), .B(n5457), .X(n19572) );
  nand_x1_sg U46985 ( .A(n19768), .B(n19769), .X(n19732) );
  nand_x1_sg U46986 ( .A(n19762), .B(n19763), .X(n19735) );
  nand_x1_sg U46987 ( .A(n19750), .B(n19751), .X(n19741) );
  nand_x1_sg U46988 ( .A(n46554), .B(n19747), .X(n19745) );
  nand_x1_sg U46989 ( .A(n20790), .B(n46577), .X(n20789) );
  nor_x1_sg U46990 ( .A(n21206), .B(n5628), .X(n21205) );
  nor_x1_sg U46991 ( .A(n19964), .B(n19965), .X(n19963) );
  nor_x1_sg U46992 ( .A(n19966), .B(n5497), .X(n19965) );
  nor_x1_sg U46993 ( .A(n21367), .B(n21368), .X(n21201) );
  nor_x1_sg U46994 ( .A(n21369), .B(n5648), .X(n21368) );
  nand_x1_sg U46995 ( .A(n21017), .B(n21018), .X(n20957) );
  nand_x1_sg U46996 ( .A(n19720), .B(n19721), .X(n19718) );
  nor_x1_sg U46997 ( .A(n19577), .B(n19578), .X(n19500) );
  nor_x1_sg U46998 ( .A(n19579), .B(n5459), .X(n19578) );
  nor_x1_sg U46999 ( .A(n19348), .B(n5440), .X(n19347) );
  nor_x1_sg U47000 ( .A(n20156), .B(n20157), .X(n20155) );
  nor_x1_sg U47001 ( .A(n20158), .B(n5517), .X(n20157) );
  nor_x1_sg U47002 ( .A(n21371), .B(n21372), .X(n21370) );
  nor_x1_sg U47003 ( .A(n21373), .B(n5649), .X(n21372) );
  nor_x1_sg U47004 ( .A(n20605), .B(n20606), .X(n20604) );
  nor_x1_sg U47005 ( .A(n20607), .B(n5574), .X(n20606) );
  nor_x1_sg U47006 ( .A(n21210), .B(n46495), .X(n21164) );
  inv_x1_sg U47007 ( .A(n21211), .X(n46495) );
  nor_x1_sg U47008 ( .A(n19350), .B(n19351), .X(n19349) );
  inv_x1_sg U47009 ( .A(n19352), .X(n46436) );
  nor_x1_sg U47010 ( .A(n21375), .B(n21376), .X(n21374) );
  nor_x1_sg U47011 ( .A(n21377), .B(n5650), .X(n21376) );
  nor_x1_sg U47012 ( .A(n21213), .B(n46457), .X(n21158) );
  inv_x1_sg U47013 ( .A(n21214), .X(n46457) );
  nor_x1_sg U47014 ( .A(n20161), .B(n5518), .X(n20160) );
  nor_x1_sg U47015 ( .A(n21379), .B(n21380), .X(n21378) );
  nor_x1_sg U47016 ( .A(n21381), .B(n5651), .X(n21380) );
  nor_x1_sg U47017 ( .A(n21216), .B(n46409), .X(n21152) );
  inv_x1_sg U47018 ( .A(n21217), .X(n46409) );
  nand_x1_sg U47019 ( .A(n46346), .B(n19794), .X(n19704) );
  nor_x1_sg U47020 ( .A(n21383), .B(n21384), .X(n21382) );
  nor_x1_sg U47021 ( .A(n21385), .B(n5652), .X(n21384) );
  nor_x1_sg U47022 ( .A(n20613), .B(n20614), .X(n20612) );
  nor_x1_sg U47023 ( .A(n20615), .B(n5576), .X(n20614) );
  nor_x1_sg U47024 ( .A(n21219), .B(n46362), .X(n21146) );
  inv_x1_sg U47025 ( .A(n21220), .X(n46362) );
  nor_x1_sg U47026 ( .A(n19797), .B(n46302), .X(n19698) );
  inv_x1_sg U47027 ( .A(n19798), .X(n46302) );
  nor_x1_sg U47028 ( .A(n19977), .B(n19978), .X(n19976) );
  nor_x1_sg U47029 ( .A(n19979), .B(n5501), .X(n19978) );
  nor_x1_sg U47030 ( .A(n20454), .B(n46311), .X(n20431) );
  inv_x1_sg U47031 ( .A(n20455), .X(n46311) );
  nor_x1_sg U47032 ( .A(n21387), .B(n21388), .X(n21386) );
  nor_x1_sg U47033 ( .A(n21389), .B(n5653), .X(n21388) );
  nor_x1_sg U47034 ( .A(n20617), .B(n20618), .X(n20616) );
  nor_x1_sg U47035 ( .A(n20619), .B(n5577), .X(n20618) );
  nor_x1_sg U47036 ( .A(n21222), .B(n46320), .X(n21140) );
  inv_x1_sg U47037 ( .A(n21223), .X(n46320) );
  nor_x1_sg U47038 ( .A(n19800), .B(n46257), .X(n19692) );
  inv_x1_sg U47039 ( .A(n19801), .X(n46257) );
  nor_x1_sg U47040 ( .A(n19981), .B(n19982), .X(n19980) );
  nor_x1_sg U47041 ( .A(n19983), .B(n5502), .X(n19982) );
  nor_x1_sg U47042 ( .A(n20457), .B(n46266), .X(n20425) );
  inv_x1_sg U47043 ( .A(n20458), .X(n46266) );
  nor_x1_sg U47044 ( .A(n21391), .B(n21392), .X(n21390) );
  nor_x1_sg U47045 ( .A(n21393), .B(n5654), .X(n21392) );
  nor_x1_sg U47046 ( .A(n20621), .B(n20622), .X(n20620) );
  nor_x1_sg U47047 ( .A(n20623), .B(n5578), .X(n20622) );
  nor_x1_sg U47048 ( .A(n21225), .B(n46275), .X(n21134) );
  inv_x1_sg U47049 ( .A(n21226), .X(n46275) );
  nor_x1_sg U47050 ( .A(n19803), .B(n46211), .X(n19686) );
  inv_x1_sg U47051 ( .A(n19804), .X(n46211) );
  nor_x1_sg U47052 ( .A(n19985), .B(n19986), .X(n19984) );
  nor_x1_sg U47053 ( .A(n19987), .B(n5503), .X(n19986) );
  nor_x1_sg U47054 ( .A(n20460), .B(n46220), .X(n20419) );
  inv_x1_sg U47055 ( .A(n20461), .X(n46220) );
  nor_x1_sg U47056 ( .A(n21395), .B(n21396), .X(n21394) );
  nor_x1_sg U47057 ( .A(n21397), .B(n5655), .X(n21396) );
  nor_x1_sg U47058 ( .A(n20625), .B(n20626), .X(n20624) );
  nor_x1_sg U47059 ( .A(n20627), .B(n5579), .X(n20626) );
  nor_x1_sg U47060 ( .A(n21228), .B(n46229), .X(n21128) );
  inv_x1_sg U47061 ( .A(n21229), .X(n46229) );
  nor_x1_sg U47062 ( .A(n19806), .B(n46166), .X(n19680) );
  inv_x1_sg U47063 ( .A(n19807), .X(n46166) );
  nor_x1_sg U47064 ( .A(n19989), .B(n19990), .X(n19988) );
  nor_x1_sg U47065 ( .A(n19991), .B(n5504), .X(n19990) );
  nor_x1_sg U47066 ( .A(n20463), .B(n46175), .X(n20413) );
  inv_x1_sg U47067 ( .A(n20464), .X(n46175) );
  nor_x1_sg U47068 ( .A(n21399), .B(n21400), .X(n21398) );
  nor_x1_sg U47069 ( .A(n21401), .B(n5656), .X(n21400) );
  nor_x1_sg U47070 ( .A(n20629), .B(n20630), .X(n20628) );
  nor_x1_sg U47071 ( .A(n20631), .B(n5580), .X(n20630) );
  nor_x1_sg U47072 ( .A(n21231), .B(n46184), .X(n21122) );
  inv_x1_sg U47073 ( .A(n21232), .X(n46184) );
  nor_x1_sg U47074 ( .A(n19809), .B(n46120), .X(n19674) );
  inv_x1_sg U47075 ( .A(n19810), .X(n46120) );
  nor_x1_sg U47076 ( .A(n19993), .B(n19994), .X(n19992) );
  nor_x1_sg U47077 ( .A(n19995), .B(n5505), .X(n19994) );
  nor_x1_sg U47078 ( .A(n20466), .B(n46129), .X(n20407) );
  inv_x1_sg U47079 ( .A(n20467), .X(n46129) );
  nor_x1_sg U47080 ( .A(n21403), .B(n21404), .X(n21402) );
  nor_x1_sg U47081 ( .A(n21405), .B(n5657), .X(n21404) );
  nor_x1_sg U47082 ( .A(n20633), .B(n20634), .X(n20632) );
  nor_x1_sg U47083 ( .A(n20635), .B(n5581), .X(n20634) );
  nor_x1_sg U47084 ( .A(n21234), .B(n46138), .X(n21116) );
  inv_x1_sg U47085 ( .A(n21235), .X(n46138) );
  nor_x1_sg U47086 ( .A(n19812), .B(n46075), .X(n19668) );
  inv_x1_sg U47087 ( .A(n19813), .X(n46075) );
  nor_x1_sg U47088 ( .A(n19997), .B(n19998), .X(n19996) );
  nor_x1_sg U47089 ( .A(n19999), .B(n5506), .X(n19998) );
  nor_x1_sg U47090 ( .A(n20469), .B(n46084), .X(n20401) );
  inv_x1_sg U47091 ( .A(n20470), .X(n46084) );
  nor_x1_sg U47092 ( .A(n21407), .B(n21408), .X(n21406) );
  nor_x1_sg U47093 ( .A(n21409), .B(n5658), .X(n21408) );
  nor_x1_sg U47094 ( .A(n20637), .B(n20638), .X(n20636) );
  nor_x1_sg U47095 ( .A(n20639), .B(n5582), .X(n20638) );
  nor_x1_sg U47096 ( .A(n21237), .B(n46093), .X(n21110) );
  inv_x1_sg U47097 ( .A(n21238), .X(n46093) );
  nor_x1_sg U47098 ( .A(n19815), .B(n46029), .X(n19662) );
  inv_x1_sg U47099 ( .A(n19816), .X(n46029) );
  nor_x1_sg U47100 ( .A(n20001), .B(n20002), .X(n20000) );
  nor_x1_sg U47101 ( .A(n20003), .B(n5507), .X(n20002) );
  nor_x1_sg U47102 ( .A(n20472), .B(n46038), .X(n20395) );
  inv_x1_sg U47103 ( .A(n20473), .X(n46038) );
  nor_x1_sg U47104 ( .A(n21411), .B(n21412), .X(n21410) );
  nor_x1_sg U47105 ( .A(n21413), .B(n5659), .X(n21412) );
  nor_x1_sg U47106 ( .A(n20641), .B(n20642), .X(n20640) );
  nor_x1_sg U47107 ( .A(n20643), .B(n5583), .X(n20642) );
  nor_x1_sg U47108 ( .A(n21240), .B(n46047), .X(n21104) );
  inv_x1_sg U47109 ( .A(n21241), .X(n46047) );
  nor_x1_sg U47110 ( .A(n19818), .B(n45984), .X(n19656) );
  inv_x1_sg U47111 ( .A(n19819), .X(n45984) );
  nor_x1_sg U47112 ( .A(n20005), .B(n20006), .X(n20004) );
  nor_x1_sg U47113 ( .A(n20007), .B(n5508), .X(n20006) );
  nor_x1_sg U47114 ( .A(n20475), .B(n45993), .X(n20389) );
  inv_x1_sg U47115 ( .A(n20476), .X(n45993) );
  nor_x1_sg U47116 ( .A(n21415), .B(n21416), .X(n21414) );
  nor_x1_sg U47117 ( .A(n21417), .B(n5660), .X(n21416) );
  nor_x1_sg U47118 ( .A(n20645), .B(n20646), .X(n20644) );
  nor_x1_sg U47119 ( .A(n20647), .B(n5584), .X(n20646) );
  nor_x1_sg U47120 ( .A(n21243), .B(n46002), .X(n21098) );
  inv_x1_sg U47121 ( .A(n21244), .X(n46002) );
  nor_x1_sg U47122 ( .A(n19823), .B(n5490), .X(n19822) );
  nor_x1_sg U47123 ( .A(n19614), .B(n19615), .X(n19418) );
  nor_x1_sg U47124 ( .A(n19616), .B(n5471), .X(n19615) );
  nor_x1_sg U47125 ( .A(n20009), .B(n20010), .X(n20008) );
  inv_x1_sg U47126 ( .A(n20011), .X(n45940) );
  nor_x1_sg U47127 ( .A(n20480), .B(n5566), .X(n20479) );
  nor_x1_sg U47128 ( .A(n21419), .B(n21420), .X(n21418) );
  inv_x1_sg U47129 ( .A(n21421), .X(n45958) );
  nor_x1_sg U47130 ( .A(n20649), .B(n20650), .X(n20648) );
  inv_x1_sg U47131 ( .A(n20651), .X(n45949) );
  nor_x1_sg U47132 ( .A(n21248), .B(n5642), .X(n21247) );
  nor_x1_sg U47133 ( .A(n19825), .B(n19826), .X(n19824) );
  nor_x1_sg U47134 ( .A(n19827), .B(n5491), .X(n19826) );
  nor_x1_sg U47135 ( .A(n20351), .B(n20352), .X(n20350) );
  nor_x1_sg U47136 ( .A(n20353), .B(n5548), .X(n20352) );
  nor_x1_sg U47137 ( .A(n20482), .B(n20483), .X(n20481) );
  nor_x1_sg U47138 ( .A(n20484), .B(n5567), .X(n20483) );
  nor_x1_sg U47139 ( .A(n21060), .B(n21061), .X(n21059) );
  nor_x1_sg U47140 ( .A(n21062), .B(n5624), .X(n21061) );
  nor_x1_sg U47141 ( .A(n21250), .B(n21251), .X(n21249) );
  nor_x1_sg U47142 ( .A(n21252), .B(n5643), .X(n21251) );
  nand_x1_sg U47143 ( .A(n7341), .B(n46992), .X(n7330) );
  nand_x1_sg U47144 ( .A(n7441), .B(n7442), .X(n7392) );
  nand_x1_sg U47145 ( .A(n7435), .B(n7436), .X(n7391) );
  inv_x1_sg U47146 ( .A(n7427), .X(n47035) );
  nand_x1_sg U47147 ( .A(n7569), .B(n7570), .X(n7035) );
  nand_x1_sg U47148 ( .A(n7526), .B(n47063), .X(n7481) );
  nand_x1_sg U47149 ( .A(n46955), .B(n7489), .X(n7465) );
  nand_x1_sg U47150 ( .A(n7506), .B(n46981), .X(n7499) );
  nand_x2_sg U47151 ( .A(n7500), .B(n7501), .X(n7498) );
  nand_x1_sg U47152 ( .A(n7027), .B(n7028), .X(n7025) );
  nand_x1_sg U47153 ( .A(n47105), .B(n7029), .X(n7028) );
  nand_x1_sg U47154 ( .A(n7032), .B(n7033), .X(n7031) );
  nand_x1_sg U47155 ( .A(n6999), .B(n7000), .X(n6985) );
  nand_x1_sg U47156 ( .A(n6988), .B(n6989), .X(n6987) );
  nand_x1_sg U47157 ( .A(n7008), .B(n7009), .X(n7007) );
  inv_x1_sg U47158 ( .A(n7603), .X(n46972) );
  nand_x1_sg U47159 ( .A(n8159), .B(n47281), .X(n8148) );
  nand_x1_sg U47160 ( .A(n8253), .B(n8254), .X(n8209) );
  nand_x1_sg U47161 ( .A(n8259), .B(n8260), .X(n8210) );
  inv_x1_sg U47162 ( .A(n8245), .X(n47322) );
  nand_x1_sg U47163 ( .A(n8387), .B(n8388), .X(n7853) );
  nand_x1_sg U47164 ( .A(n8344), .B(n47349), .X(n8299) );
  nand_x1_sg U47165 ( .A(n47246), .B(n8307), .X(n8283) );
  nand_x1_sg U47166 ( .A(n8324), .B(n47271), .X(n8317) );
  nand_x2_sg U47167 ( .A(n8318), .B(n8319), .X(n8316) );
  nand_x1_sg U47168 ( .A(n7845), .B(n7846), .X(n7843) );
  nand_x1_sg U47169 ( .A(n47391), .B(n7847), .X(n7846) );
  nand_x1_sg U47170 ( .A(n7850), .B(n7851), .X(n7849) );
  nand_x1_sg U47171 ( .A(n7816), .B(n7817), .X(n7802) );
  nand_x1_sg U47172 ( .A(n7805), .B(n7806), .X(n7804) );
  nand_x1_sg U47173 ( .A(n7825), .B(n7826), .X(n7824) );
  inv_x1_sg U47174 ( .A(n8421), .X(n47262) );
  nand_x1_sg U47175 ( .A(n8977), .B(n47566), .X(n8966) );
  nand_x1_sg U47176 ( .A(n9071), .B(n9072), .X(n9027) );
  nand_x1_sg U47177 ( .A(n9077), .B(n9078), .X(n9028) );
  inv_x1_sg U47178 ( .A(n9063), .X(n47607) );
  nand_x1_sg U47179 ( .A(n9205), .B(n9206), .X(n8671) );
  nand_x1_sg U47180 ( .A(n9162), .B(n47634), .X(n9117) );
  nand_x1_sg U47181 ( .A(n47531), .B(n9125), .X(n9101) );
  nand_x1_sg U47182 ( .A(n9142), .B(n47556), .X(n9135) );
  nand_x2_sg U47183 ( .A(n9136), .B(n9137), .X(n9134) );
  nand_x1_sg U47184 ( .A(n8663), .B(n8664), .X(n8661) );
  nand_x1_sg U47185 ( .A(n47676), .B(n8665), .X(n8664) );
  nand_x1_sg U47186 ( .A(n8668), .B(n8669), .X(n8667) );
  nand_x1_sg U47187 ( .A(n8634), .B(n8635), .X(n8620) );
  nand_x1_sg U47188 ( .A(n8623), .B(n8624), .X(n8622) );
  nand_x1_sg U47189 ( .A(n8643), .B(n8644), .X(n8642) );
  inv_x1_sg U47190 ( .A(n9239), .X(n47547) );
  nand_x1_sg U47191 ( .A(n9797), .B(n47851), .X(n9786) );
  nand_x1_sg U47192 ( .A(n9891), .B(n9892), .X(n9847) );
  nand_x1_sg U47193 ( .A(n9897), .B(n9898), .X(n9848) );
  inv_x1_sg U47194 ( .A(n9883), .X(n47892) );
  nand_x1_sg U47195 ( .A(n10025), .B(n10026), .X(n9491) );
  nand_x1_sg U47196 ( .A(n9982), .B(n47919), .X(n9937) );
  nand_x1_sg U47197 ( .A(n47816), .B(n9945), .X(n9921) );
  nand_x1_sg U47198 ( .A(n9962), .B(n47841), .X(n9955) );
  nand_x2_sg U47199 ( .A(n9956), .B(n9957), .X(n9954) );
  nand_x1_sg U47200 ( .A(n9483), .B(n9484), .X(n9481) );
  nand_x1_sg U47201 ( .A(n47961), .B(n9485), .X(n9484) );
  nand_x1_sg U47202 ( .A(n9488), .B(n9489), .X(n9487) );
  nand_x1_sg U47203 ( .A(n9454), .B(n9455), .X(n9440) );
  nand_x1_sg U47204 ( .A(n9443), .B(n9444), .X(n9442) );
  nand_x1_sg U47205 ( .A(n9463), .B(n9464), .X(n9462) );
  inv_x1_sg U47206 ( .A(n10059), .X(n47832) );
  nand_x1_sg U47207 ( .A(n10616), .B(n48136), .X(n10605) );
  nand_x1_sg U47208 ( .A(n10710), .B(n10711), .X(n10666) );
  nand_x1_sg U47209 ( .A(n10716), .B(n10717), .X(n10667) );
  inv_x1_sg U47210 ( .A(n10702), .X(n48177) );
  nand_x1_sg U47211 ( .A(n10844), .B(n10845), .X(n10310) );
  nand_x1_sg U47212 ( .A(n10801), .B(n48204), .X(n10756) );
  nand_x1_sg U47213 ( .A(n48101), .B(n10764), .X(n10740) );
  nand_x1_sg U47214 ( .A(n10781), .B(n48126), .X(n10774) );
  nand_x2_sg U47215 ( .A(n10775), .B(n10776), .X(n10773) );
  nand_x1_sg U47216 ( .A(n10302), .B(n10303), .X(n10300) );
  nand_x1_sg U47217 ( .A(n48246), .B(n10304), .X(n10303) );
  nand_x1_sg U47218 ( .A(n10307), .B(n10308), .X(n10306) );
  nand_x1_sg U47219 ( .A(n10273), .B(n10274), .X(n10259) );
  nand_x1_sg U47220 ( .A(n10262), .B(n10263), .X(n10261) );
  nand_x1_sg U47221 ( .A(n10282), .B(n10283), .X(n10281) );
  inv_x1_sg U47222 ( .A(n10878), .X(n48117) );
  nand_x1_sg U47223 ( .A(n11435), .B(n48421), .X(n11424) );
  nand_x1_sg U47224 ( .A(n11529), .B(n11530), .X(n11485) );
  nand_x1_sg U47225 ( .A(n11535), .B(n11536), .X(n11486) );
  inv_x1_sg U47226 ( .A(n11521), .X(n48462) );
  nand_x1_sg U47227 ( .A(n11663), .B(n11664), .X(n11129) );
  nand_x1_sg U47228 ( .A(n11620), .B(n48489), .X(n11575) );
  nand_x1_sg U47229 ( .A(n48386), .B(n11583), .X(n11559) );
  nand_x1_sg U47230 ( .A(n11600), .B(n48411), .X(n11593) );
  nand_x2_sg U47231 ( .A(n11594), .B(n11595), .X(n11592) );
  nand_x1_sg U47232 ( .A(n11121), .B(n11122), .X(n11119) );
  nand_x1_sg U47233 ( .A(n48531), .B(n11123), .X(n11122) );
  nand_x1_sg U47234 ( .A(n11126), .B(n11127), .X(n11125) );
  nand_x1_sg U47235 ( .A(n11092), .B(n11093), .X(n11078) );
  nand_x1_sg U47236 ( .A(n11081), .B(n11082), .X(n11080) );
  nand_x1_sg U47237 ( .A(n11101), .B(n11102), .X(n11100) );
  inv_x1_sg U47238 ( .A(n11697), .X(n48402) );
  nand_x1_sg U47239 ( .A(n12254), .B(n48706), .X(n12243) );
  nand_x1_sg U47240 ( .A(n12348), .B(n12349), .X(n12304) );
  nand_x1_sg U47241 ( .A(n12354), .B(n12355), .X(n12305) );
  inv_x1_sg U47242 ( .A(n12340), .X(n48747) );
  nand_x1_sg U47243 ( .A(n12482), .B(n12483), .X(n11948) );
  nand_x1_sg U47244 ( .A(n12439), .B(n48774), .X(n12394) );
  nand_x1_sg U47245 ( .A(n48671), .B(n12402), .X(n12378) );
  nand_x1_sg U47246 ( .A(n12419), .B(n48696), .X(n12412) );
  nand_x2_sg U47247 ( .A(n12413), .B(n12414), .X(n12411) );
  nand_x1_sg U47248 ( .A(n11940), .B(n11941), .X(n11938) );
  nand_x1_sg U47249 ( .A(n48816), .B(n11942), .X(n11941) );
  nand_x1_sg U47250 ( .A(n11945), .B(n11946), .X(n11944) );
  nand_x1_sg U47251 ( .A(n11911), .B(n11912), .X(n11897) );
  nand_x1_sg U47252 ( .A(n11900), .B(n11901), .X(n11899) );
  nand_x1_sg U47253 ( .A(n11920), .B(n11921), .X(n11919) );
  inv_x1_sg U47254 ( .A(n12516), .X(n48687) );
  nand_x1_sg U47255 ( .A(n13073), .B(n48992), .X(n13062) );
  nand_x1_sg U47256 ( .A(n13167), .B(n13168), .X(n13123) );
  nand_x1_sg U47257 ( .A(n13173), .B(n13174), .X(n13124) );
  inv_x1_sg U47258 ( .A(n13159), .X(n49033) );
  nand_x1_sg U47259 ( .A(n13301), .B(n13302), .X(n12767) );
  nand_x1_sg U47260 ( .A(n13258), .B(n49061), .X(n13213) );
  nand_x1_sg U47261 ( .A(n48957), .B(n13221), .X(n13197) );
  nand_x1_sg U47262 ( .A(n13238), .B(n48982), .X(n13231) );
  nand_x2_sg U47263 ( .A(n13232), .B(n13233), .X(n13230) );
  nand_x1_sg U47264 ( .A(n12759), .B(n12760), .X(n12757) );
  nand_x1_sg U47265 ( .A(n49103), .B(n12761), .X(n12760) );
  nand_x1_sg U47266 ( .A(n12764), .B(n12765), .X(n12763) );
  nand_x1_sg U47267 ( .A(n12730), .B(n12731), .X(n12716) );
  nand_x1_sg U47268 ( .A(n12719), .B(n12720), .X(n12718) );
  nand_x1_sg U47269 ( .A(n12739), .B(n12740), .X(n12738) );
  inv_x1_sg U47270 ( .A(n13335), .X(n48973) );
  nand_x1_sg U47271 ( .A(n13892), .B(n49279), .X(n13881) );
  nand_x1_sg U47272 ( .A(n13986), .B(n13987), .X(n13942) );
  nand_x1_sg U47273 ( .A(n13992), .B(n13993), .X(n13943) );
  inv_x1_sg U47274 ( .A(n13978), .X(n49320) );
  nand_x1_sg U47275 ( .A(n14120), .B(n14121), .X(n13586) );
  nand_x1_sg U47276 ( .A(n14077), .B(n49347), .X(n14032) );
  nand_x1_sg U47277 ( .A(n49244), .B(n14040), .X(n14016) );
  nand_x1_sg U47278 ( .A(n14057), .B(n49269), .X(n14050) );
  nand_x2_sg U47279 ( .A(n14051), .B(n14052), .X(n14049) );
  nand_x1_sg U47280 ( .A(n13578), .B(n13579), .X(n13576) );
  nand_x1_sg U47281 ( .A(n49389), .B(n13580), .X(n13579) );
  nand_x1_sg U47282 ( .A(n13583), .B(n13584), .X(n13582) );
  nand_x1_sg U47283 ( .A(n13549), .B(n13550), .X(n13535) );
  nand_x1_sg U47284 ( .A(n13538), .B(n13539), .X(n13537) );
  nand_x1_sg U47285 ( .A(n13558), .B(n13559), .X(n13557) );
  inv_x1_sg U47286 ( .A(n14154), .X(n49260) );
  nand_x1_sg U47287 ( .A(n14711), .B(n49565), .X(n14700) );
  nand_x1_sg U47288 ( .A(n14805), .B(n14806), .X(n14761) );
  nand_x1_sg U47289 ( .A(n14811), .B(n14812), .X(n14762) );
  inv_x1_sg U47290 ( .A(n14797), .X(n49606) );
  nand_x1_sg U47291 ( .A(n14939), .B(n14940), .X(n14405) );
  nand_x1_sg U47292 ( .A(n14896), .B(n49633), .X(n14851) );
  nand_x1_sg U47293 ( .A(n49530), .B(n14859), .X(n14835) );
  nand_x1_sg U47294 ( .A(n14876), .B(n49555), .X(n14869) );
  nand_x2_sg U47295 ( .A(n14870), .B(n14871), .X(n14868) );
  nand_x1_sg U47296 ( .A(n14397), .B(n14398), .X(n14395) );
  nand_x1_sg U47297 ( .A(n49675), .B(n14399), .X(n14398) );
  nand_x1_sg U47298 ( .A(n14402), .B(n14403), .X(n14401) );
  nand_x1_sg U47299 ( .A(n14368), .B(n14369), .X(n14354) );
  nand_x1_sg U47300 ( .A(n14357), .B(n14358), .X(n14356) );
  nand_x1_sg U47301 ( .A(n14377), .B(n14378), .X(n14376) );
  inv_x1_sg U47302 ( .A(n14973), .X(n49546) );
  nand_x1_sg U47303 ( .A(n15530), .B(n49851), .X(n15519) );
  nand_x1_sg U47304 ( .A(n15624), .B(n15625), .X(n15580) );
  nand_x1_sg U47305 ( .A(n15630), .B(n15631), .X(n15581) );
  inv_x1_sg U47306 ( .A(n15616), .X(n49892) );
  nand_x1_sg U47307 ( .A(n15758), .B(n15759), .X(n15224) );
  nand_x1_sg U47308 ( .A(n15715), .B(n49919), .X(n15670) );
  nand_x1_sg U47309 ( .A(n49816), .B(n15678), .X(n15654) );
  nand_x1_sg U47310 ( .A(n15695), .B(n49841), .X(n15688) );
  nand_x2_sg U47311 ( .A(n15689), .B(n15690), .X(n15687) );
  nand_x1_sg U47312 ( .A(n15216), .B(n15217), .X(n15214) );
  nand_x1_sg U47313 ( .A(n49961), .B(n15218), .X(n15217) );
  nand_x1_sg U47314 ( .A(n15221), .B(n15222), .X(n15220) );
  nand_x1_sg U47315 ( .A(n15187), .B(n15188), .X(n15173) );
  nand_x1_sg U47316 ( .A(n15176), .B(n15177), .X(n15175) );
  nand_x1_sg U47317 ( .A(n15196), .B(n15197), .X(n15195) );
  inv_x1_sg U47318 ( .A(n15792), .X(n49832) );
  nand_x1_sg U47319 ( .A(n16349), .B(n50137), .X(n16338) );
  nand_x1_sg U47320 ( .A(n16443), .B(n16444), .X(n16399) );
  nand_x1_sg U47321 ( .A(n16449), .B(n16450), .X(n16400) );
  inv_x1_sg U47322 ( .A(n16435), .X(n50178) );
  nand_x1_sg U47323 ( .A(n16577), .B(n16578), .X(n16043) );
  nand_x1_sg U47324 ( .A(n16534), .B(n50205), .X(n16489) );
  nand_x1_sg U47325 ( .A(n50102), .B(n16497), .X(n16473) );
  nand_x1_sg U47326 ( .A(n16514), .B(n50127), .X(n16507) );
  nand_x2_sg U47327 ( .A(n16508), .B(n16509), .X(n16506) );
  nand_x1_sg U47328 ( .A(n16035), .B(n16036), .X(n16033) );
  nand_x1_sg U47329 ( .A(n50247), .B(n16037), .X(n16036) );
  nand_x1_sg U47330 ( .A(n16040), .B(n16041), .X(n16039) );
  nand_x1_sg U47331 ( .A(n16006), .B(n16007), .X(n15992) );
  nand_x1_sg U47332 ( .A(n15995), .B(n15996), .X(n15994) );
  nand_x1_sg U47333 ( .A(n16015), .B(n16016), .X(n16014) );
  inv_x1_sg U47334 ( .A(n16611), .X(n50118) );
  nand_x1_sg U47335 ( .A(n17166), .B(n50422), .X(n17155) );
  nand_x1_sg U47336 ( .A(n17266), .B(n17267), .X(n17217) );
  nand_x1_sg U47337 ( .A(n17260), .B(n17261), .X(n17216) );
  inv_x1_sg U47338 ( .A(n17252), .X(n50463) );
  inv_x1_sg U47339 ( .A(n17290), .X(n50388) );
  nand_x1_sg U47340 ( .A(n17394), .B(n17395), .X(n16862) );
  nand_x1_sg U47341 ( .A(n17351), .B(n50490), .X(n17306) );
  nand_x1_sg U47342 ( .A(n50387), .B(n17314), .X(n17290) );
  nand_x2_sg U47343 ( .A(n17325), .B(n17326), .X(n17323) );
  nand_x1_sg U47344 ( .A(n17331), .B(n50412), .X(n17324) );
  nand_x1_sg U47345 ( .A(n16823), .B(n16824), .X(n16809) );
  nand_x1_sg U47346 ( .A(n16812), .B(n16813), .X(n16811) );
  nand_x1_sg U47347 ( .A(n16832), .B(n16833), .X(n16831) );
  nand_x1_sg U47348 ( .A(n16854), .B(n16855), .X(n16852) );
  nand_x1_sg U47349 ( .A(n50532), .B(n16856), .X(n16855) );
  nand_x1_sg U47350 ( .A(n16859), .B(n16860), .X(n16858) );
  inv_x1_sg U47351 ( .A(n17428), .X(n50403) );
  nand_x1_sg U47352 ( .A(n17987), .B(n50711), .X(n17976) );
  nand_x1_sg U47353 ( .A(n18081), .B(n18082), .X(n18037) );
  nand_x1_sg U47354 ( .A(n18087), .B(n18088), .X(n18038) );
  inv_x1_sg U47355 ( .A(n18073), .X(n50752) );
  nand_x1_sg U47356 ( .A(n18215), .B(n18216), .X(n17681) );
  nand_x1_sg U47357 ( .A(n18172), .B(n50779), .X(n18127) );
  nand_x1_sg U47358 ( .A(n50676), .B(n18135), .X(n18111) );
  nand_x1_sg U47359 ( .A(n18152), .B(n50701), .X(n18145) );
  nand_x2_sg U47360 ( .A(n18146), .B(n18147), .X(n18144) );
  nand_x1_sg U47361 ( .A(n17673), .B(n17674), .X(n17671) );
  nand_x1_sg U47362 ( .A(n50821), .B(n17675), .X(n17674) );
  nand_x1_sg U47363 ( .A(n17678), .B(n17679), .X(n17677) );
  nand_x1_sg U47364 ( .A(n17644), .B(n17645), .X(n17630) );
  nand_x1_sg U47365 ( .A(n17633), .B(n17634), .X(n17632) );
  nand_x1_sg U47366 ( .A(n17653), .B(n17654), .X(n17652) );
  inv_x1_sg U47367 ( .A(n18249), .X(n50692) );
  nand_x1_sg U47368 ( .A(n18808), .B(n50998), .X(n18797) );
  nand_x1_sg U47369 ( .A(n18902), .B(n18903), .X(n18858) );
  nand_x1_sg U47370 ( .A(n18908), .B(n18909), .X(n18859) );
  inv_x1_sg U47371 ( .A(n18894), .X(n51039) );
  nand_x1_sg U47372 ( .A(n19036), .B(n19037), .X(n18502) );
  nand_x1_sg U47373 ( .A(n18993), .B(n51066), .X(n18948) );
  nand_x1_sg U47374 ( .A(n50963), .B(n18956), .X(n18932) );
  nand_x1_sg U47375 ( .A(n18973), .B(n50988), .X(n18966) );
  nand_x2_sg U47376 ( .A(n18967), .B(n18968), .X(n18965) );
  nand_x1_sg U47377 ( .A(n18494), .B(n18495), .X(n18492) );
  nand_x1_sg U47378 ( .A(n51108), .B(n18496), .X(n18495) );
  nand_x1_sg U47379 ( .A(n18499), .B(n18500), .X(n18498) );
  nand_x1_sg U47380 ( .A(n18465), .B(n18466), .X(n18451) );
  nand_x1_sg U47381 ( .A(n18454), .B(n18455), .X(n18453) );
  nand_x1_sg U47382 ( .A(n18474), .B(n18475), .X(n18473) );
  inv_x1_sg U47383 ( .A(n19070), .X(n50979) );
  nor_x1_sg U47384 ( .A(n27332), .B(n27333), .X(n27106) );
  nor_x1_sg U47385 ( .A(n27334), .B(n5268), .X(n27333) );
  nor_x1_sg U47386 ( .A(n27545), .B(n27546), .X(n27336) );
  nor_x1_sg U47387 ( .A(n27547), .B(n5269), .X(n27546) );
  nor_x1_sg U47388 ( .A(n27739), .B(n27740), .X(n27549) );
  nor_x1_sg U47389 ( .A(n27741), .B(n5270), .X(n27740) );
  nor_x1_sg U47390 ( .A(n27916), .B(n27917), .X(n27743) );
  nor_x1_sg U47391 ( .A(n27918), .B(n5271), .X(n27917) );
  nor_x1_sg U47392 ( .A(n28078), .B(n28079), .X(n27920) );
  nor_x1_sg U47393 ( .A(n28080), .B(n5272), .X(n28079) );
  nor_x1_sg U47394 ( .A(n28213), .B(n28214), .X(n28082) );
  nor_x1_sg U47395 ( .A(n28215), .B(n5273), .X(n28214) );
  nor_x1_sg U47396 ( .A(n28217), .B(n28218), .X(n28216) );
  nor_x1_sg U47397 ( .A(n28219), .B(n5274), .X(n28218) );
  nor_x1_sg U47398 ( .A(n28221), .B(n28222), .X(n28220) );
  nor_x1_sg U47399 ( .A(n28223), .B(n5275), .X(n28222) );
  nor_x1_sg U47400 ( .A(n28225), .B(n28226), .X(n28224) );
  nor_x1_sg U47401 ( .A(n28227), .B(n5276), .X(n28226) );
  nor_x1_sg U47402 ( .A(n28229), .B(n28230), .X(n28228) );
  nor_x1_sg U47403 ( .A(n28231), .B(n5277), .X(n28230) );
  nor_x1_sg U47404 ( .A(n28233), .B(n28234), .X(n28232) );
  nor_x1_sg U47405 ( .A(n28235), .B(n5278), .X(n28234) );
  nor_x1_sg U47406 ( .A(n28237), .B(n28238), .X(n28236) );
  nor_x1_sg U47407 ( .A(n28239), .B(n5279), .X(n28238) );
  nor_x1_sg U47408 ( .A(n28241), .B(n28242), .X(n28240) );
  nor_x1_sg U47409 ( .A(n28243), .B(n5280), .X(n28242) );
  nor_x1_sg U47410 ( .A(n28245), .B(n28246), .X(n28244) );
  inv_x1_sg U47411 ( .A(n28247), .X(n45102) );
  nor_x1_sg U47412 ( .A(n45058), .B(n28248), .X(n28142) );
  inv_x1_sg U47413 ( .A(n28250), .X(n45058) );
  nand_x1_sg U47414 ( .A(n28363), .B(n28364), .X(n28267) );
  nand_x1_sg U47415 ( .A(n19561), .B(n19562), .X(n19559) );
  nand_x1_sg U47416 ( .A(n46611), .B(n19568), .X(n19566) );
  nor_x1_sg U47417 ( .A(n19758), .B(n46559), .X(n19543) );
  inv_x1_sg U47418 ( .A(n19759), .X(n46559) );
  nand_x1_sg U47419 ( .A(n19554), .B(n19555), .X(n19552) );
  nand_x1_sg U47420 ( .A(n19547), .B(n19548), .X(n19545) );
  nand_x1_sg U47421 ( .A(n19533), .B(n19534), .X(n19531) );
  nand_x1_sg U47422 ( .A(n20995), .B(n20996), .X(n20993) );
  nand_x1_sg U47423 ( .A(n46592), .B(n20586), .X(n20584) );
  nand_x1_sg U47424 ( .A(n46588), .B(n21003), .X(n21001) );
  nor_x1_sg U47425 ( .A(n19340), .B(n19341), .X(n19145) );
  inv_x1_sg U47426 ( .A(n19342), .X(n46573) );
  nand_x1_sg U47427 ( .A(n19774), .B(n19775), .X(n19729) );
  nand_x1_sg U47428 ( .A(n19335), .B(n19336), .X(n19333) );
  nand_x1_sg U47429 ( .A(n5456), .B(n46575), .X(n19336) );
  nand_x1_sg U47430 ( .A(n19756), .B(n19757), .X(n19738) );
  inv_x1_sg U47431 ( .A(n19733), .X(n46602) );
  inv_x1_sg U47432 ( .A(n19736), .X(n46600) );
  inv_x1_sg U47433 ( .A(n19742), .X(n46596) );
  nor_x1_sg U47434 ( .A(n21197), .B(n21198), .X(n20998) );
  nor_x1_sg U47435 ( .A(n21199), .B(n5647), .X(n21198) );
  nor_x1_sg U47436 ( .A(n21014), .B(n21015), .X(n20786) );
  inv_x1_sg U47437 ( .A(n21016), .X(n46579) );
  nand_x1_sg U47438 ( .A(n20787), .B(n20788), .X(n20780) );
  nand_x1_sg U47439 ( .A(n5589), .B(n20789), .X(n20788) );
  nand_x1_sg U47440 ( .A(n21202), .B(n21203), .X(n21173) );
  nand_x1_sg U47441 ( .A(n5627), .B(n46581), .X(n21203) );
  inv_x1_sg U47442 ( .A(n19727), .X(n46531) );
  nand_x1_sg U47443 ( .A(n46527), .B(n19326), .X(n19325) );
  nor_x1_sg U47444 ( .A(n19962), .B(n5496), .X(n19961) );
  nand_x1_sg U47445 ( .A(n19952), .B(n19953), .X(n19926) );
  nor_x1_sg U47446 ( .A(n46509), .B(n19942), .X(n19755) );
  inv_x1_sg U47447 ( .A(n19945), .X(n46509) );
  nand_x1_sg U47448 ( .A(n20955), .B(n20956), .X(n20954) );
  nand_x1_sg U47449 ( .A(n5609), .B(n20957), .X(n20956) );
  nor_x1_sg U47450 ( .A(n21207), .B(n46536), .X(n21170) );
  inv_x1_sg U47451 ( .A(n21208), .X(n46536) );
  nand_x1_sg U47452 ( .A(n19498), .B(n19499), .X(n19496) );
  nand_x1_sg U47453 ( .A(n19500), .B(n38195), .X(n19498) );
  inv_x1_sg U47454 ( .A(n19921), .X(n46487) );
  nor_x1_sg U47455 ( .A(n20154), .B(n5516), .X(n20153) );
  nor_x1_sg U47456 ( .A(n20601), .B(n20602), .X(n20136) );
  nor_x1_sg U47457 ( .A(n20603), .B(n5573), .X(n20602) );
  nand_x1_sg U47458 ( .A(n21162), .B(n46496), .X(n21161) );
  nand_x1_sg U47459 ( .A(n19583), .B(n42087), .X(n19580) );
  nand_x1_sg U47460 ( .A(n46443), .B(n19714), .X(n19713) );
  nor_x1_sg U47461 ( .A(n20317), .B(n20318), .X(n20316) );
  inv_x1_sg U47462 ( .A(n20319), .X(n46399) );
  nand_x1_sg U47463 ( .A(n19914), .B(n19915), .X(n19913) );
  inv_x1_sg U47464 ( .A(n20121), .X(n46448) );
  nand_x1_sg U47465 ( .A(n46451), .B(n20302), .X(n20301) );
  nand_x1_sg U47466 ( .A(n21156), .B(n46458), .X(n21155) );
  nand_x1_sg U47467 ( .A(n46394), .B(n19708), .X(n19707) );
  nand_x1_sg U47468 ( .A(n19485), .B(n19486), .X(n19483) );
  nand_x1_sg U47469 ( .A(n5460), .B(n42087), .X(n19486) );
  nor_x1_sg U47470 ( .A(n19353), .B(n19354), .X(n19311) );
  inv_x1_sg U47471 ( .A(n19355), .X(n46388) );
  nand_x1_sg U47472 ( .A(n20114), .B(n20115), .X(n20112) );
  nor_x1_sg U47473 ( .A(n19970), .B(n19971), .X(n19909) );
  nor_x1_sg U47474 ( .A(n19972), .B(n5499), .X(n19971) );
  nand_x1_sg U47475 ( .A(n46378), .B(n20446), .X(n20440) );
  nand_x1_sg U47476 ( .A(n46403), .B(n20444), .X(n20443) );
  nand_x1_sg U47477 ( .A(n21150), .B(n46410), .X(n21149) );
  nand_x1_sg U47478 ( .A(n19702), .B(n19703), .X(n19701) );
  nand_x1_sg U47479 ( .A(n5480), .B(n19704), .X(n19703) );
  nor_x1_sg U47480 ( .A(n19975), .B(n5500), .X(n19974) );
  nand_x1_sg U47481 ( .A(n46350), .B(n20107), .X(n20106) );
  nand_x1_sg U47482 ( .A(n21144), .B(n46363), .X(n21143) );
  nor_x1_sg U47483 ( .A(n19173), .B(n19174), .X(n19172) );
  nor_x1_sg U47484 ( .A(n19175), .B(n5425), .X(n19174) );
  nand_x1_sg U47485 ( .A(n19696), .B(n46303), .X(n19695) );
  nand_x1_sg U47486 ( .A(n19472), .B(n19473), .X(n19471) );
  nand_x1_sg U47487 ( .A(n5462), .B(n19474), .X(n19473) );
  nand_x1_sg U47488 ( .A(n20429), .B(n46312), .X(n20428) );
  nand_x1_sg U47489 ( .A(n21138), .B(n46321), .X(n21137) );
  nor_x1_sg U47490 ( .A(n19177), .B(n19178), .X(n19176) );
  nor_x1_sg U47491 ( .A(n19179), .B(n5426), .X(n19178) );
  nand_x1_sg U47492 ( .A(n19690), .B(n46258), .X(n19689) );
  nand_x1_sg U47493 ( .A(n19465), .B(n19466), .X(n19464) );
  nand_x1_sg U47494 ( .A(n5463), .B(n19467), .X(n19466) );
  nand_x1_sg U47495 ( .A(n20423), .B(n46267), .X(n20422) );
  nand_x1_sg U47496 ( .A(n21132), .B(n46276), .X(n21131) );
  nor_x1_sg U47497 ( .A(n19181), .B(n19182), .X(n19180) );
  nor_x1_sg U47498 ( .A(n19183), .B(n5427), .X(n19182) );
  nand_x1_sg U47499 ( .A(n19684), .B(n46212), .X(n19683) );
  nand_x1_sg U47500 ( .A(n19458), .B(n19459), .X(n19457) );
  nand_x1_sg U47501 ( .A(n5464), .B(n19460), .X(n19459) );
  nand_x1_sg U47502 ( .A(n20417), .B(n46221), .X(n20416) );
  nand_x1_sg U47503 ( .A(n21126), .B(n46230), .X(n21125) );
  nor_x1_sg U47504 ( .A(n19185), .B(n19186), .X(n19184) );
  nor_x1_sg U47505 ( .A(n19187), .B(n5428), .X(n19186) );
  nand_x1_sg U47506 ( .A(n19678), .B(n46167), .X(n19677) );
  nand_x1_sg U47507 ( .A(n19451), .B(n19452), .X(n19450) );
  nand_x1_sg U47508 ( .A(n5465), .B(n19453), .X(n19452) );
  nand_x1_sg U47509 ( .A(n20411), .B(n46176), .X(n20410) );
  nand_x1_sg U47510 ( .A(n21120), .B(n46185), .X(n21119) );
  nand_x1_sg U47511 ( .A(n19672), .B(n46121), .X(n19671) );
  nor_x1_sg U47512 ( .A(n19189), .B(n19190), .X(n19188) );
  nor_x1_sg U47513 ( .A(n19191), .B(n5429), .X(n19190) );
  nand_x1_sg U47514 ( .A(n20405), .B(n46130), .X(n20404) );
  nand_x1_sg U47515 ( .A(n21114), .B(n46139), .X(n21113) );
  nor_x1_sg U47516 ( .A(n19193), .B(n19194), .X(n19192) );
  nor_x1_sg U47517 ( .A(n19195), .B(n5430), .X(n19194) );
  nand_x1_sg U47518 ( .A(n19666), .B(n46076), .X(n19665) );
  nand_x1_sg U47519 ( .A(n19437), .B(n19438), .X(n19436) );
  nand_x1_sg U47520 ( .A(n5467), .B(n19439), .X(n19438) );
  nand_x1_sg U47521 ( .A(n20399), .B(n46085), .X(n20398) );
  nand_x1_sg U47522 ( .A(n21108), .B(n46094), .X(n21107) );
  nor_x1_sg U47523 ( .A(n19197), .B(n19198), .X(n19196) );
  nor_x1_sg U47524 ( .A(n19199), .B(n5431), .X(n19198) );
  nand_x1_sg U47525 ( .A(n19660), .B(n46030), .X(n19659) );
  nand_x1_sg U47526 ( .A(n19430), .B(n19431), .X(n19429) );
  nand_x1_sg U47527 ( .A(n5468), .B(n19432), .X(n19431) );
  nand_x1_sg U47528 ( .A(n20393), .B(n46039), .X(n20392) );
  nand_x1_sg U47529 ( .A(n21102), .B(n46048), .X(n21101) );
  nor_x1_sg U47530 ( .A(n19201), .B(n19202), .X(n19200) );
  nor_x1_sg U47531 ( .A(n19203), .B(n5432), .X(n19202) );
  nand_x1_sg U47532 ( .A(n19654), .B(n45985), .X(n19653) );
  nand_x1_sg U47533 ( .A(n19423), .B(n19424), .X(n19422) );
  nand_x1_sg U47534 ( .A(n5469), .B(n19425), .X(n19424) );
  nand_x1_sg U47535 ( .A(n20387), .B(n45994), .X(n20386) );
  nand_x1_sg U47536 ( .A(n21096), .B(n46003), .X(n21095) );
  nor_x1_sg U47537 ( .A(n19205), .B(n19206), .X(n19204) );
  inv_x1_sg U47538 ( .A(n19207), .X(n45931) );
  nand_x1_sg U47539 ( .A(n19648), .B(n45939), .X(n19647) );
  nand_x1_sg U47540 ( .A(n19416), .B(n19417), .X(n19415) );
  nor_x1_sg U47541 ( .A(n20347), .B(n20348), .X(n20224) );
  nor_x1_sg U47542 ( .A(n20349), .B(n5547), .X(n20348) );
  nand_x1_sg U47543 ( .A(n20381), .B(n45948), .X(n20380) );
  nor_x1_sg U47544 ( .A(n21056), .B(n21057), .X(n20867) );
  nor_x1_sg U47545 ( .A(n21058), .B(n5623), .X(n21057) );
  nand_x1_sg U47546 ( .A(n21090), .B(n45957), .X(n21089) );
  nor_x1_sg U47547 ( .A(n19386), .B(n19387), .X(n19236) );
  nor_x1_sg U47548 ( .A(n19388), .B(n5453), .X(n19387) );
  nand_x1_sg U47549 ( .A(n45889), .B(n19410), .X(n19409) );
  nor_x1_sg U47550 ( .A(n20192), .B(n20193), .X(n20040) );
  nor_x1_sg U47551 ( .A(n20194), .B(n5529), .X(n20193) );
  nor_x1_sg U47552 ( .A(n45894), .B(n20012), .X(n19851) );
  inv_x1_sg U47553 ( .A(n20014), .X(n45894) );
  nor_x1_sg U47554 ( .A(n45914), .B(n21422), .X(n21277) );
  inv_x1_sg U47555 ( .A(n21424), .X(n45914) );
  nor_x1_sg U47556 ( .A(n45904), .B(n20652), .X(n20508) );
  inv_x1_sg U47557 ( .A(n20654), .X(n45904) );
  nor_x1_sg U47558 ( .A(n20835), .B(n20836), .X(n20680) );
  nor_x1_sg U47559 ( .A(n20837), .B(n5605), .X(n20836) );
  inv_x1_sg U47560 ( .A(n19638), .X(n45855) );
  nand_x1_sg U47561 ( .A(n19404), .B(n19405), .X(n19403) );
  nand_x1_sg U47562 ( .A(n45850), .B(n19843), .X(n19842) );
  inv_x1_sg U47563 ( .A(n20032), .X(n45847) );
  inv_x1_sg U47564 ( .A(n20371), .X(n45839) );
  nand_x1_sg U47565 ( .A(n21585), .B(n21586), .X(n21443) );
  nand_x1_sg U47566 ( .A(n45818), .B(n21269), .X(n21268) );
  nand_x1_sg U47567 ( .A(n45834), .B(n20500), .X(n20499) );
  inv_x1_sg U47568 ( .A(n20672), .X(n45831) );
  inv_x1_sg U47569 ( .A(n21080), .X(n45823) );
  nand_x1_sg U47570 ( .A(n7151), .B(n7152), .X(n7137) );
  nand_x1_sg U47571 ( .A(n46880), .B(n7155), .X(n7138) );
  nor_x1_sg U47572 ( .A(n7212), .B(n46915), .X(n7210) );
  inv_x1_sg U47573 ( .A(n7213), .X(n46915) );
  nor_x1_sg U47574 ( .A(n7277), .B(n7278), .X(n7276) );
  nor_x1_sg U47575 ( .A(n7338), .B(n7339), .X(n7288) );
  nor_x1_sg U47576 ( .A(n7327), .B(n7328), .X(n7308) );
  nand_x1_sg U47577 ( .A(n7386), .B(n7387), .X(n7361) );
  inv_x1_sg U47578 ( .A(n7370), .X(n46986) );
  nand_x1_sg U47579 ( .A(n7393), .B(n7434), .X(n7423) );
  nand_x1_sg U47580 ( .A(n7466), .B(n47034), .X(n7427) );
  nand_x2_sg U47581 ( .A(n7546), .B(n7547), .X(n7519) );
  nand_x1_sg U47582 ( .A(n7538), .B(n47084), .X(n7524) );
  inv_x1_sg U47583 ( .A(n7026), .X(n47108) );
  nand_x1_sg U47584 ( .A(n47062), .B(n7020), .X(n7017) );
  inv_x1_sg U47585 ( .A(n7005), .X(n47121) );
  nand_x1_sg U47586 ( .A(n7580), .B(n7581), .X(n7578) );
  inv_x1_sg U47587 ( .A(n7585), .X(n46990) );
  nand_x1_sg U47588 ( .A(n7969), .B(n7970), .X(n7955) );
  nand_x1_sg U47589 ( .A(n47173), .B(n7974), .X(n7956) );
  nor_x1_sg U47590 ( .A(n8031), .B(n47207), .X(n8029) );
  inv_x1_sg U47591 ( .A(n8032), .X(n47207) );
  nor_x1_sg U47592 ( .A(n8096), .B(n8097), .X(n8095) );
  nor_x1_sg U47593 ( .A(n8156), .B(n8157), .X(n8106) );
  nor_x1_sg U47594 ( .A(n8145), .B(n8146), .X(n8126) );
  nand_x1_sg U47595 ( .A(n8204), .B(n8205), .X(n8179) );
  inv_x1_sg U47596 ( .A(n8188), .X(n47275) );
  nand_x1_sg U47597 ( .A(n8211), .B(n8252), .X(n8241) );
  nand_x1_sg U47598 ( .A(n8284), .B(n47321), .X(n8245) );
  nand_x2_sg U47599 ( .A(n8364), .B(n8365), .X(n8337) );
  nand_x1_sg U47600 ( .A(n8356), .B(n47370), .X(n8342) );
  inv_x1_sg U47601 ( .A(n7844), .X(n47394) );
  nand_x1_sg U47602 ( .A(n47348), .B(n7838), .X(n7835) );
  inv_x1_sg U47603 ( .A(n7822), .X(n47407) );
  nand_x1_sg U47604 ( .A(n8406), .B(n47334), .X(n8397) );
  nand_x1_sg U47605 ( .A(n8398), .B(n8399), .X(n8396) );
  inv_x1_sg U47606 ( .A(n8403), .X(n47279) );
  nand_x1_sg U47607 ( .A(n8787), .B(n8788), .X(n8773) );
  nand_x1_sg U47608 ( .A(n47458), .B(n8792), .X(n8774) );
  nor_x1_sg U47609 ( .A(n8849), .B(n47492), .X(n8847) );
  inv_x1_sg U47610 ( .A(n8850), .X(n47492) );
  nor_x1_sg U47611 ( .A(n8914), .B(n8915), .X(n8913) );
  nor_x1_sg U47612 ( .A(n8974), .B(n8975), .X(n8924) );
  nor_x1_sg U47613 ( .A(n8963), .B(n8964), .X(n8944) );
  nand_x1_sg U47614 ( .A(n9022), .B(n9023), .X(n8997) );
  inv_x1_sg U47615 ( .A(n9006), .X(n47560) );
  nand_x1_sg U47616 ( .A(n9029), .B(n9070), .X(n9059) );
  nand_x1_sg U47617 ( .A(n9102), .B(n47606), .X(n9063) );
  nand_x2_sg U47618 ( .A(n9182), .B(n9183), .X(n9155) );
  nand_x1_sg U47619 ( .A(n9174), .B(n47655), .X(n9160) );
  inv_x1_sg U47620 ( .A(n8662), .X(n47679) );
  nand_x1_sg U47621 ( .A(n47633), .B(n8656), .X(n8653) );
  inv_x1_sg U47622 ( .A(n8640), .X(n47692) );
  nand_x1_sg U47623 ( .A(n9224), .B(n47619), .X(n9215) );
  nand_x1_sg U47624 ( .A(n9216), .B(n9217), .X(n9214) );
  inv_x1_sg U47625 ( .A(n9221), .X(n47564) );
  nand_x1_sg U47626 ( .A(n9607), .B(n9608), .X(n9593) );
  nand_x1_sg U47627 ( .A(n47743), .B(n9612), .X(n9594) );
  nor_x1_sg U47628 ( .A(n9669), .B(n47777), .X(n9667) );
  inv_x1_sg U47629 ( .A(n9670), .X(n47777) );
  nor_x1_sg U47630 ( .A(n9734), .B(n9735), .X(n9733) );
  nor_x1_sg U47631 ( .A(n9794), .B(n9795), .X(n9744) );
  nor_x1_sg U47632 ( .A(n9783), .B(n9784), .X(n9764) );
  nand_x1_sg U47633 ( .A(n9842), .B(n9843), .X(n9817) );
  inv_x1_sg U47634 ( .A(n9826), .X(n47845) );
  nand_x1_sg U47635 ( .A(n9849), .B(n9890), .X(n9879) );
  nand_x1_sg U47636 ( .A(n9922), .B(n47891), .X(n9883) );
  nand_x2_sg U47637 ( .A(n10002), .B(n10003), .X(n9975) );
  nand_x1_sg U47638 ( .A(n9994), .B(n47940), .X(n9980) );
  inv_x1_sg U47639 ( .A(n9482), .X(n47964) );
  nand_x1_sg U47640 ( .A(n47918), .B(n9476), .X(n9473) );
  inv_x1_sg U47641 ( .A(n9460), .X(n47977) );
  nand_x1_sg U47642 ( .A(n10044), .B(n47904), .X(n10035) );
  nand_x1_sg U47643 ( .A(n10036), .B(n10037), .X(n10034) );
  inv_x1_sg U47644 ( .A(n10041), .X(n47849) );
  nand_x1_sg U47645 ( .A(n10426), .B(n10427), .X(n10412) );
  nand_x1_sg U47646 ( .A(n48028), .B(n10431), .X(n10413) );
  nor_x1_sg U47647 ( .A(n10488), .B(n48062), .X(n10486) );
  inv_x1_sg U47648 ( .A(n10489), .X(n48062) );
  nor_x1_sg U47649 ( .A(n10553), .B(n10554), .X(n10552) );
  nor_x1_sg U47650 ( .A(n10613), .B(n10614), .X(n10563) );
  nor_x1_sg U47651 ( .A(n10602), .B(n10603), .X(n10583) );
  nand_x1_sg U47652 ( .A(n10661), .B(n10662), .X(n10636) );
  inv_x1_sg U47653 ( .A(n10645), .X(n48130) );
  nand_x1_sg U47654 ( .A(n10668), .B(n10709), .X(n10698) );
  nand_x1_sg U47655 ( .A(n10741), .B(n48176), .X(n10702) );
  nand_x2_sg U47656 ( .A(n10821), .B(n10822), .X(n10794) );
  nand_x1_sg U47657 ( .A(n10813), .B(n48225), .X(n10799) );
  inv_x1_sg U47658 ( .A(n10301), .X(n48249) );
  nand_x1_sg U47659 ( .A(n48203), .B(n10295), .X(n10292) );
  inv_x1_sg U47660 ( .A(n10279), .X(n48262) );
  nand_x1_sg U47661 ( .A(n10863), .B(n48189), .X(n10854) );
  nand_x1_sg U47662 ( .A(n10855), .B(n10856), .X(n10853) );
  inv_x1_sg U47663 ( .A(n10860), .X(n48134) );
  nand_x1_sg U47664 ( .A(n11245), .B(n11246), .X(n11231) );
  nand_x1_sg U47665 ( .A(n48313), .B(n11250), .X(n11232) );
  nor_x1_sg U47666 ( .A(n11307), .B(n48347), .X(n11305) );
  inv_x1_sg U47667 ( .A(n11308), .X(n48347) );
  nor_x1_sg U47668 ( .A(n11372), .B(n11373), .X(n11371) );
  nor_x1_sg U47669 ( .A(n11432), .B(n11433), .X(n11382) );
  nor_x1_sg U47670 ( .A(n11421), .B(n11422), .X(n11402) );
  nand_x1_sg U47671 ( .A(n11480), .B(n11481), .X(n11455) );
  inv_x1_sg U47672 ( .A(n11464), .X(n48415) );
  nand_x1_sg U47673 ( .A(n11487), .B(n11528), .X(n11517) );
  nand_x1_sg U47674 ( .A(n11560), .B(n48461), .X(n11521) );
  nand_x2_sg U47675 ( .A(n11640), .B(n11641), .X(n11613) );
  nand_x1_sg U47676 ( .A(n11632), .B(n48510), .X(n11618) );
  inv_x1_sg U47677 ( .A(n11120), .X(n48534) );
  nand_x1_sg U47678 ( .A(n48488), .B(n11114), .X(n11111) );
  inv_x1_sg U47679 ( .A(n11098), .X(n48547) );
  nand_x1_sg U47680 ( .A(n11682), .B(n48474), .X(n11673) );
  nand_x1_sg U47681 ( .A(n11674), .B(n11675), .X(n11672) );
  inv_x1_sg U47682 ( .A(n11679), .X(n48419) );
  nand_x1_sg U47683 ( .A(n12064), .B(n12065), .X(n12050) );
  nand_x1_sg U47684 ( .A(n48598), .B(n12069), .X(n12051) );
  nor_x1_sg U47685 ( .A(n12126), .B(n48632), .X(n12124) );
  inv_x1_sg U47686 ( .A(n12127), .X(n48632) );
  nor_x1_sg U47687 ( .A(n12191), .B(n12192), .X(n12190) );
  nor_x1_sg U47688 ( .A(n12251), .B(n12252), .X(n12201) );
  nor_x1_sg U47689 ( .A(n12240), .B(n12241), .X(n12221) );
  nand_x1_sg U47690 ( .A(n12299), .B(n12300), .X(n12274) );
  inv_x1_sg U47691 ( .A(n12283), .X(n48700) );
  nand_x1_sg U47692 ( .A(n12306), .B(n12347), .X(n12336) );
  nand_x1_sg U47693 ( .A(n12379), .B(n48746), .X(n12340) );
  nand_x2_sg U47694 ( .A(n12459), .B(n12460), .X(n12432) );
  nand_x1_sg U47695 ( .A(n12451), .B(n48795), .X(n12437) );
  inv_x1_sg U47696 ( .A(n11939), .X(n48819) );
  nand_x1_sg U47697 ( .A(n48773), .B(n11933), .X(n11930) );
  inv_x1_sg U47698 ( .A(n11917), .X(n48832) );
  nand_x1_sg U47699 ( .A(n12501), .B(n48759), .X(n12492) );
  nand_x1_sg U47700 ( .A(n12493), .B(n12494), .X(n12491) );
  inv_x1_sg U47701 ( .A(n12498), .X(n48704) );
  nand_x1_sg U47702 ( .A(n12883), .B(n12884), .X(n12869) );
  nand_x1_sg U47703 ( .A(n48884), .B(n12888), .X(n12870) );
  nor_x1_sg U47704 ( .A(n12945), .B(n48918), .X(n12943) );
  inv_x1_sg U47705 ( .A(n12946), .X(n48918) );
  nor_x1_sg U47706 ( .A(n13010), .B(n13011), .X(n13009) );
  nor_x1_sg U47707 ( .A(n13070), .B(n13071), .X(n13020) );
  nor_x1_sg U47708 ( .A(n13059), .B(n13060), .X(n13040) );
  nand_x1_sg U47709 ( .A(n13118), .B(n13119), .X(n13093) );
  inv_x1_sg U47710 ( .A(n13102), .X(n48986) );
  nand_x1_sg U47711 ( .A(n13125), .B(n13166), .X(n13155) );
  nand_x1_sg U47712 ( .A(n13198), .B(n49032), .X(n13159) );
  nand_x2_sg U47713 ( .A(n13278), .B(n13279), .X(n13251) );
  nand_x1_sg U47714 ( .A(n13270), .B(n49082), .X(n13256) );
  inv_x1_sg U47715 ( .A(n12758), .X(n49106) );
  nand_x1_sg U47716 ( .A(n49060), .B(n12752), .X(n12749) );
  inv_x1_sg U47717 ( .A(n12736), .X(n49119) );
  nand_x1_sg U47718 ( .A(n13320), .B(n49045), .X(n13311) );
  nand_x1_sg U47719 ( .A(n13312), .B(n13313), .X(n13310) );
  inv_x1_sg U47720 ( .A(n13317), .X(n48990) );
  nand_x1_sg U47721 ( .A(n13702), .B(n13703), .X(n13688) );
  nand_x1_sg U47722 ( .A(n49171), .B(n13707), .X(n13689) );
  nor_x1_sg U47723 ( .A(n13764), .B(n49205), .X(n13762) );
  inv_x1_sg U47724 ( .A(n13765), .X(n49205) );
  nor_x1_sg U47725 ( .A(n13829), .B(n13830), .X(n13828) );
  nor_x1_sg U47726 ( .A(n13889), .B(n13890), .X(n13839) );
  nor_x1_sg U47727 ( .A(n13878), .B(n13879), .X(n13859) );
  nand_x1_sg U47728 ( .A(n13937), .B(n13938), .X(n13912) );
  inv_x1_sg U47729 ( .A(n13921), .X(n49273) );
  nand_x1_sg U47730 ( .A(n13944), .B(n13985), .X(n13974) );
  nand_x1_sg U47731 ( .A(n14017), .B(n49319), .X(n13978) );
  nand_x2_sg U47732 ( .A(n14097), .B(n14098), .X(n14070) );
  nand_x1_sg U47733 ( .A(n14089), .B(n49368), .X(n14075) );
  inv_x1_sg U47734 ( .A(n13577), .X(n49392) );
  nand_x1_sg U47735 ( .A(n49346), .B(n13571), .X(n13568) );
  inv_x1_sg U47736 ( .A(n13555), .X(n49405) );
  nand_x1_sg U47737 ( .A(n14139), .B(n49332), .X(n14130) );
  nand_x1_sg U47738 ( .A(n14131), .B(n14132), .X(n14129) );
  inv_x1_sg U47739 ( .A(n14136), .X(n49277) );
  nand_x1_sg U47740 ( .A(n14521), .B(n14522), .X(n14507) );
  nand_x1_sg U47741 ( .A(n49457), .B(n14526), .X(n14508) );
  nor_x1_sg U47742 ( .A(n14583), .B(n49491), .X(n14581) );
  inv_x1_sg U47743 ( .A(n14584), .X(n49491) );
  nor_x1_sg U47744 ( .A(n14648), .B(n14649), .X(n14647) );
  nor_x1_sg U47745 ( .A(n14708), .B(n14709), .X(n14658) );
  nor_x1_sg U47746 ( .A(n14697), .B(n14698), .X(n14678) );
  nand_x1_sg U47747 ( .A(n14756), .B(n14757), .X(n14731) );
  inv_x1_sg U47748 ( .A(n14740), .X(n49559) );
  nand_x1_sg U47749 ( .A(n14763), .B(n14804), .X(n14793) );
  nand_x1_sg U47750 ( .A(n14836), .B(n49605), .X(n14797) );
  nand_x2_sg U47751 ( .A(n14916), .B(n14917), .X(n14889) );
  nand_x1_sg U47752 ( .A(n14908), .B(n49654), .X(n14894) );
  inv_x1_sg U47753 ( .A(n14396), .X(n49678) );
  nand_x1_sg U47754 ( .A(n49632), .B(n14390), .X(n14387) );
  inv_x1_sg U47755 ( .A(n14374), .X(n49691) );
  nand_x1_sg U47756 ( .A(n14958), .B(n49618), .X(n14949) );
  nand_x1_sg U47757 ( .A(n14950), .B(n14951), .X(n14948) );
  inv_x1_sg U47758 ( .A(n14955), .X(n49563) );
  nand_x1_sg U47759 ( .A(n15340), .B(n15341), .X(n15326) );
  nand_x1_sg U47760 ( .A(n49742), .B(n15345), .X(n15327) );
  nor_x1_sg U47761 ( .A(n15402), .B(n49777), .X(n15400) );
  inv_x1_sg U47762 ( .A(n15403), .X(n49777) );
  nor_x1_sg U47763 ( .A(n15467), .B(n15468), .X(n15466) );
  nor_x1_sg U47764 ( .A(n15527), .B(n15528), .X(n15477) );
  nor_x1_sg U47765 ( .A(n15516), .B(n15517), .X(n15497) );
  nand_x1_sg U47766 ( .A(n15575), .B(n15576), .X(n15550) );
  inv_x1_sg U47767 ( .A(n15559), .X(n49845) );
  nand_x1_sg U47768 ( .A(n15582), .B(n15623), .X(n15612) );
  nand_x1_sg U47769 ( .A(n15655), .B(n49891), .X(n15616) );
  nand_x2_sg U47770 ( .A(n15735), .B(n15736), .X(n15708) );
  nand_x1_sg U47771 ( .A(n15727), .B(n49940), .X(n15713) );
  inv_x1_sg U47772 ( .A(n15215), .X(n49964) );
  nand_x1_sg U47773 ( .A(n49918), .B(n15209), .X(n15206) );
  inv_x1_sg U47774 ( .A(n15193), .X(n49977) );
  nand_x1_sg U47775 ( .A(n15777), .B(n49904), .X(n15768) );
  nand_x1_sg U47776 ( .A(n15769), .B(n15770), .X(n15767) );
  inv_x1_sg U47777 ( .A(n15774), .X(n49849) );
  nand_x1_sg U47778 ( .A(n16159), .B(n16160), .X(n16145) );
  nand_x1_sg U47779 ( .A(n50029), .B(n16164), .X(n16146) );
  nor_x1_sg U47780 ( .A(n16221), .B(n50063), .X(n16219) );
  inv_x1_sg U47781 ( .A(n16222), .X(n50063) );
  nor_x1_sg U47782 ( .A(n16286), .B(n16287), .X(n16285) );
  nor_x1_sg U47783 ( .A(n16346), .B(n16347), .X(n16296) );
  nor_x1_sg U47784 ( .A(n16335), .B(n16336), .X(n16316) );
  nand_x1_sg U47785 ( .A(n16394), .B(n16395), .X(n16369) );
  inv_x1_sg U47786 ( .A(n16378), .X(n50131) );
  nand_x1_sg U47787 ( .A(n16401), .B(n16442), .X(n16431) );
  nand_x1_sg U47788 ( .A(n16474), .B(n50177), .X(n16435) );
  nand_x2_sg U47789 ( .A(n16554), .B(n16555), .X(n16527) );
  nand_x1_sg U47790 ( .A(n16546), .B(n50226), .X(n16532) );
  inv_x1_sg U47791 ( .A(n16034), .X(n50250) );
  nand_x1_sg U47792 ( .A(n50204), .B(n16028), .X(n16025) );
  inv_x1_sg U47793 ( .A(n16012), .X(n50263) );
  nand_x1_sg U47794 ( .A(n16596), .B(n50190), .X(n16587) );
  nand_x1_sg U47795 ( .A(n16588), .B(n16589), .X(n16586) );
  inv_x1_sg U47796 ( .A(n16593), .X(n50135) );
  nand_x1_sg U47797 ( .A(n16976), .B(n16977), .X(n16962) );
  nand_x1_sg U47798 ( .A(n50314), .B(n16980), .X(n16963) );
  nor_x1_sg U47799 ( .A(n17037), .B(n50348), .X(n17035) );
  inv_x1_sg U47800 ( .A(n17038), .X(n50348) );
  nor_x1_sg U47801 ( .A(n17102), .B(n17103), .X(n17101) );
  nor_x1_sg U47802 ( .A(n17163), .B(n17164), .X(n17113) );
  nor_x1_sg U47803 ( .A(n17152), .B(n17153), .X(n17133) );
  nand_x1_sg U47804 ( .A(n17211), .B(n17212), .X(n17186) );
  inv_x1_sg U47805 ( .A(n17195), .X(n50416) );
  nand_x1_sg U47806 ( .A(n17218), .B(n17259), .X(n17248) );
  nand_x1_sg U47807 ( .A(n17291), .B(n50462), .X(n17252) );
  nand_x2_sg U47808 ( .A(n17371), .B(n17372), .X(n17344) );
  nand_x1_sg U47809 ( .A(n17363), .B(n50511), .X(n17349) );
  inv_x1_sg U47810 ( .A(n16829), .X(n50549) );
  inv_x1_sg U47811 ( .A(n16853), .X(n50535) );
  nand_x1_sg U47812 ( .A(n50489), .B(n16845), .X(n16842) );
  nand_x1_sg U47813 ( .A(n17405), .B(n17406), .X(n17403) );
  inv_x1_sg U47814 ( .A(n17410), .X(n50420) );
  nand_x1_sg U47815 ( .A(n17797), .B(n17798), .X(n17783) );
  nand_x1_sg U47816 ( .A(n50603), .B(n17802), .X(n17784) );
  nor_x1_sg U47817 ( .A(n17859), .B(n50637), .X(n17857) );
  inv_x1_sg U47818 ( .A(n17860), .X(n50637) );
  nor_x1_sg U47819 ( .A(n17924), .B(n17925), .X(n17923) );
  nor_x1_sg U47820 ( .A(n17984), .B(n17985), .X(n17934) );
  nor_x1_sg U47821 ( .A(n17973), .B(n17974), .X(n17954) );
  nand_x1_sg U47822 ( .A(n18032), .B(n18033), .X(n18007) );
  inv_x1_sg U47823 ( .A(n18016), .X(n50705) );
  nand_x1_sg U47824 ( .A(n18039), .B(n18080), .X(n18069) );
  nand_x1_sg U47825 ( .A(n18112), .B(n50751), .X(n18073) );
  nand_x2_sg U47826 ( .A(n18192), .B(n18193), .X(n18165) );
  nand_x1_sg U47827 ( .A(n18184), .B(n50800), .X(n18170) );
  inv_x1_sg U47828 ( .A(n17672), .X(n50824) );
  nand_x1_sg U47829 ( .A(n50778), .B(n17666), .X(n17663) );
  inv_x1_sg U47830 ( .A(n17650), .X(n50837) );
  nand_x1_sg U47831 ( .A(n18234), .B(n50764), .X(n18225) );
  nand_x1_sg U47832 ( .A(n18226), .B(n18227), .X(n18224) );
  inv_x1_sg U47833 ( .A(n18231), .X(n50709) );
  nand_x1_sg U47834 ( .A(n18618), .B(n18619), .X(n18604) );
  nand_x1_sg U47835 ( .A(n50890), .B(n18623), .X(n18605) );
  nor_x1_sg U47836 ( .A(n18680), .B(n50924), .X(n18678) );
  inv_x1_sg U47837 ( .A(n18681), .X(n50924) );
  nor_x1_sg U47838 ( .A(n18745), .B(n18746), .X(n18744) );
  nor_x1_sg U47839 ( .A(n18805), .B(n18806), .X(n18755) );
  nor_x1_sg U47840 ( .A(n18794), .B(n18795), .X(n18775) );
  nand_x1_sg U47841 ( .A(n18853), .B(n18854), .X(n18828) );
  inv_x1_sg U47842 ( .A(n18837), .X(n50992) );
  nand_x1_sg U47843 ( .A(n18860), .B(n18901), .X(n18890) );
  nand_x1_sg U47844 ( .A(n18933), .B(n51038), .X(n18894) );
  nand_x2_sg U47845 ( .A(n19013), .B(n19014), .X(n18986) );
  nand_x1_sg U47846 ( .A(n19005), .B(n51087), .X(n18991) );
  inv_x1_sg U47847 ( .A(n18493), .X(n51111) );
  nand_x1_sg U47848 ( .A(n51065), .B(n18487), .X(n18484) );
  inv_x1_sg U47849 ( .A(n18471), .X(n51124) );
  nand_x1_sg U47850 ( .A(n19055), .B(n51051), .X(n19046) );
  nand_x1_sg U47851 ( .A(n19047), .B(n19048), .X(n19045) );
  inv_x1_sg U47852 ( .A(n19052), .X(n50996) );
  nand_x1_sg U47853 ( .A(n26869), .B(n26870), .X(n26868) );
  nand_x1_sg U47854 ( .A(n26847), .B(n26848), .X(n26845) );
  nand_x1_sg U47855 ( .A(n26840), .B(n26841), .X(n26839) );
  nand_x1_sg U47856 ( .A(n26862), .B(n26863), .X(n26861) );
  nand_x1_sg U47857 ( .A(n26855), .B(n26856), .X(n26854) );
  nand_x1_sg U47858 ( .A(n26876), .B(n26877), .X(n26875) );
  nor_x1_sg U47859 ( .A(n27102), .B(n27103), .X(n26850) );
  nor_x1_sg U47860 ( .A(n27104), .B(n5267), .X(n27103) );
  nand_x1_sg U47861 ( .A(n27094), .B(n27095), .X(n27078) );
  nand_x1_sg U47862 ( .A(n5285), .B(n26843), .X(n27095) );
  nand_x1_sg U47863 ( .A(n27324), .B(n27325), .X(n27308) );
  nand_x1_sg U47864 ( .A(n5286), .B(n27099), .X(n27325) );
  nand_x1_sg U47865 ( .A(n27537), .B(n27538), .X(n27521) );
  nand_x1_sg U47866 ( .A(n5287), .B(n27329), .X(n27538) );
  nand_x1_sg U47867 ( .A(n27731), .B(n27732), .X(n27715) );
  nand_x1_sg U47868 ( .A(n5288), .B(n27542), .X(n27732) );
  nand_x1_sg U47869 ( .A(n27908), .B(n27909), .X(n27892) );
  nand_x1_sg U47870 ( .A(n5289), .B(n27736), .X(n27909) );
  nand_x1_sg U47871 ( .A(n28070), .B(n28071), .X(n28054) );
  nand_x1_sg U47872 ( .A(n5290), .B(n27913), .X(n28071) );
  nand_x1_sg U47873 ( .A(n28205), .B(n28206), .X(n28189) );
  nand_x1_sg U47874 ( .A(n5291), .B(n28075), .X(n28206) );
  nand_x1_sg U47875 ( .A(n28334), .B(n28335), .X(n28318) );
  nand_x1_sg U47876 ( .A(n5292), .B(n28210), .X(n28335) );
  nand_x1_sg U47877 ( .A(n28271), .B(n28272), .X(n28269) );
  nand_x1_sg U47878 ( .A(n5300), .B(n28273), .X(n28272) );
  nand_x1_sg U47879 ( .A(n28140), .B(n45059), .X(n28138) );
  nand_x1_sg U47880 ( .A(n27797), .B(n27798), .X(n27628) );
  nand_x1_sg U47881 ( .A(n28265), .B(n28266), .X(n28264) );
  nand_x1_sg U47882 ( .A(n27965), .B(n27966), .X(n27814) );
  nand_x1_sg U47883 ( .A(n27408), .B(n27409), .X(n27203) );
  nand_x1_sg U47884 ( .A(n44997), .B(n28134), .X(n28132) );
  nand_x1_sg U47885 ( .A(n28118), .B(n28119), .X(n27984) );
  nand_x1_sg U47886 ( .A(n27612), .B(n27613), .X(n27425) );
  nand_x1_sg U47887 ( .A(n46606), .B(n19143), .X(n19141) );
  nand_x1_sg U47888 ( .A(n46603), .B(n19558), .X(n19515) );
  nand_x1_sg U47889 ( .A(n46612), .B(n19565), .X(n19512) );
  nand_x1_sg U47890 ( .A(n19150), .B(n19151), .X(n19148) );
  nand_x1_sg U47891 ( .A(n19540), .B(n19541), .X(n19538) );
  nand_x1_sg U47892 ( .A(n46601), .B(n19551), .X(n19518) );
  nand_x1_sg U47893 ( .A(n46599), .B(n19544), .X(n19521) );
  nand_x1_sg U47894 ( .A(n46595), .B(n19530), .X(n19528) );
  nand_x1_sg U47895 ( .A(n20988), .B(n20989), .X(n20987) );
  nand_x1_sg U47896 ( .A(n46587), .B(n20992), .X(n20970) );
  nand_x1_sg U47897 ( .A(n21010), .B(n21011), .X(n21008) );
  nand_x1_sg U47898 ( .A(n46614), .B(n20589), .X(n20577) );
  nand_x1_sg U47899 ( .A(n46593), .B(n20583), .X(n20581) );
  nand_x1_sg U47900 ( .A(n46589), .B(n21000), .X(n20967) );
  nand_x1_sg U47901 ( .A(n19338), .B(n19339), .X(n19330) );
  nand_x1_sg U47902 ( .A(n5437), .B(n46574), .X(n19339) );
  nor_x1_sg U47903 ( .A(n19153), .B(n19154), .X(n5983) );
  nor_x1_sg U47904 ( .A(n19155), .B(n5419), .X(n19154) );
  inv_x1_sg U47905 ( .A(n19739), .X(n46598) );
  nand_x1_sg U47906 ( .A(n21189), .B(n21190), .X(n21179) );
  nand_x1_sg U47907 ( .A(n5665), .B(n20991), .X(n21190) );
  nand_x1_sg U47908 ( .A(n21195), .B(n21196), .X(n21176) );
  nand_x1_sg U47909 ( .A(n20784), .B(n20785), .X(n20782) );
  nand_x1_sg U47910 ( .A(n21171), .B(n46590), .X(n21013) );
  nand_x1_sg U47911 ( .A(n19505), .B(n19506), .X(n19503) );
  nor_x1_sg U47912 ( .A(n19950), .B(n5534), .X(n19949) );
  nand_x1_sg U47913 ( .A(n19958), .B(n46532), .X(n19923) );
  nor_x1_sg U47914 ( .A(n19940), .B(n19941), .X(n19933) );
  nand_x1_sg U47915 ( .A(n21359), .B(n21360), .X(n21349) );
  nand_x1_sg U47916 ( .A(n5666), .B(n21194), .X(n21360) );
  nand_x1_sg U47917 ( .A(n46540), .B(n21365), .X(n21346) );
  nand_x1_sg U47918 ( .A(n46533), .B(n19937), .X(n19935) );
  inv_x1_sg U47919 ( .A(n20776), .X(n46534) );
  nor_x1_sg U47920 ( .A(n21168), .B(n21169), .X(n21167) );
  nand_x1_sg U47921 ( .A(n46482), .B(n19320), .X(n19318) );
  nand_x1_sg U47922 ( .A(n20144), .B(n20145), .X(n20126) );
  nand_x1_sg U47923 ( .A(n20150), .B(n46488), .X(n20123) );
  nand_x1_sg U47924 ( .A(n46472), .B(n20137), .X(n20129) );
  nand_x1_sg U47925 ( .A(n21541), .B(n21542), .X(n21531) );
  nand_x1_sg U47926 ( .A(n5667), .B(n21364), .X(n21542) );
  nand_x1_sg U47927 ( .A(n46498), .B(n21342), .X(n21340) );
  nand_x1_sg U47928 ( .A(n20949), .B(n20950), .X(n20948) );
  nand_x1_sg U47929 ( .A(n5610), .B(n20951), .X(n20950) );
  nand_x1_sg U47930 ( .A(n20134), .B(n20135), .X(n20133) );
  nand_x1_sg U47931 ( .A(n20769), .B(n20770), .X(n20767) );
  nand_x1_sg U47932 ( .A(n5591), .B(n20771), .X(n20770) );
  inv_x1_sg U47933 ( .A(n19493), .X(n46441) );
  inv_x1_sg U47934 ( .A(n19316), .X(n46438) );
  nor_x1_sg U47935 ( .A(n19163), .B(n19164), .X(n6131) );
  nor_x1_sg U47936 ( .A(n19165), .B(n5422), .X(n19164) );
  nor_x1_sg U47937 ( .A(n20315), .B(n5536), .X(n20314) );
  nand_x1_sg U47938 ( .A(n46426), .B(n20304), .X(n20298) );
  nor_x1_sg U47939 ( .A(n21717), .B(n21718), .X(n21675) );
  nand_x1_sg U47940 ( .A(n46460), .B(n21336), .X(n21335) );
  nand_x1_sg U47941 ( .A(n20942), .B(n20943), .X(n20941) );
  nand_x1_sg U47942 ( .A(n5611), .B(n20944), .X(n20943) );
  nand_x1_sg U47943 ( .A(n20762), .B(n20763), .X(n20760) );
  nand_x1_sg U47944 ( .A(n5592), .B(n20764), .X(n20763) );
  nand_x1_sg U47945 ( .A(n19705), .B(n19706), .X(n19583) );
  nand_x1_sg U47946 ( .A(n19309), .B(n19310), .X(n19307) );
  nand_x1_sg U47947 ( .A(n5441), .B(n46389), .X(n19310) );
  inv_x1_sg U47948 ( .A(n20292), .X(n46401) );
  nand_x1_sg U47949 ( .A(n19907), .B(n19908), .X(n19905) );
  nand_x1_sg U47950 ( .A(n19909), .B(n38194), .X(n19907) );
  nand_x1_sg U47951 ( .A(n46412), .B(n21331), .X(n21330) );
  nand_x1_sg U47952 ( .A(n20935), .B(n20936), .X(n20934) );
  nand_x1_sg U47953 ( .A(n5612), .B(n20937), .X(n20936) );
  nand_x1_sg U47954 ( .A(n20755), .B(n20756), .X(n20753) );
  nand_x1_sg U47955 ( .A(n5593), .B(n20757), .X(n20756) );
  nand_x1_sg U47956 ( .A(n19356), .B(n19357), .X(n19305) );
  nand_x1_sg U47957 ( .A(n46344), .B(n19479), .X(n19477) );
  nor_x1_sg U47958 ( .A(n19169), .B(n19170), .X(n6223) );
  nor_x1_sg U47959 ( .A(n19171), .B(n5424), .X(n19170) );
  nand_x1_sg U47960 ( .A(n20320), .B(n20321), .X(n20286) );
  nor_x1_sg U47961 ( .A(n19901), .B(n19902), .X(n19900) );
  inv_x1_sg U47962 ( .A(n20436), .X(n46353) );
  nor_x1_sg U47963 ( .A(n21665), .B(n21666), .X(n21664) );
  nand_x1_sg U47964 ( .A(n46365), .B(n21326), .X(n21325) );
  nand_x1_sg U47965 ( .A(n20928), .B(n20929), .X(n20927) );
  nand_x1_sg U47966 ( .A(n5613), .B(n20930), .X(n20929) );
  nand_x1_sg U47967 ( .A(n46356), .B(n20557), .X(n20556) );
  nand_x1_sg U47968 ( .A(n20748), .B(n20749), .X(n20746) );
  nand_x1_sg U47969 ( .A(n5594), .B(n20750), .X(n20749) );
  nand_x1_sg U47970 ( .A(n19297), .B(n19298), .X(n19295) );
  nand_x1_sg U47971 ( .A(n5443), .B(n19299), .X(n19298) );
  nand_x1_sg U47972 ( .A(n20278), .B(n20279), .X(n20277) );
  nand_x1_sg U47973 ( .A(n5538), .B(n20280), .X(n20279) );
  nand_x1_sg U47974 ( .A(n46305), .B(n19895), .X(n19894) );
  nand_x1_sg U47975 ( .A(n20101), .B(n20102), .X(n20099) );
  nand_x1_sg U47976 ( .A(n5519), .B(n20103), .X(n20102) );
  nand_x1_sg U47977 ( .A(n46323), .B(n21321), .X(n21320) );
  nand_x1_sg U47978 ( .A(n20921), .B(n20922), .X(n20920) );
  nand_x1_sg U47979 ( .A(n5614), .B(n20923), .X(n20922) );
  nand_x1_sg U47980 ( .A(n46314), .B(n20552), .X(n20551) );
  nand_x1_sg U47981 ( .A(n20741), .B(n20742), .X(n20739) );
  nand_x1_sg U47982 ( .A(n5595), .B(n20743), .X(n20742) );
  nand_x1_sg U47983 ( .A(n19290), .B(n19291), .X(n19288) );
  nand_x1_sg U47984 ( .A(n5444), .B(n19292), .X(n19291) );
  nand_x1_sg U47985 ( .A(n20271), .B(n20272), .X(n20270) );
  nand_x1_sg U47986 ( .A(n5539), .B(n20273), .X(n20272) );
  nand_x1_sg U47987 ( .A(n46260), .B(n19890), .X(n19889) );
  nand_x1_sg U47988 ( .A(n20094), .B(n20095), .X(n20092) );
  nand_x1_sg U47989 ( .A(n5520), .B(n20096), .X(n20095) );
  nor_x1_sg U47990 ( .A(n21653), .B(n21654), .X(n21652) );
  nand_x1_sg U47991 ( .A(n46278), .B(n21316), .X(n21315) );
  nand_x1_sg U47992 ( .A(n20914), .B(n20915), .X(n20913) );
  nand_x1_sg U47993 ( .A(n5615), .B(n20916), .X(n20915) );
  nand_x1_sg U47994 ( .A(n46269), .B(n20547), .X(n20546) );
  nand_x1_sg U47995 ( .A(n20734), .B(n20735), .X(n20732) );
  nand_x1_sg U47996 ( .A(n5596), .B(n20736), .X(n20735) );
  nand_x1_sg U47997 ( .A(n19283), .B(n19284), .X(n19281) );
  nand_x1_sg U47998 ( .A(n5445), .B(n19285), .X(n19284) );
  nand_x1_sg U47999 ( .A(n20264), .B(n20265), .X(n20263) );
  nand_x1_sg U48000 ( .A(n5540), .B(n20266), .X(n20265) );
  nand_x1_sg U48001 ( .A(n46214), .B(n19885), .X(n19884) );
  nand_x1_sg U48002 ( .A(n20087), .B(n20088), .X(n20085) );
  nand_x1_sg U48003 ( .A(n5521), .B(n20089), .X(n20088) );
  nand_x1_sg U48004 ( .A(n46232), .B(n21311), .X(n21310) );
  nand_x1_sg U48005 ( .A(n20907), .B(n20908), .X(n20906) );
  nand_x1_sg U48006 ( .A(n5616), .B(n20909), .X(n20908) );
  nand_x1_sg U48007 ( .A(n46223), .B(n20542), .X(n20541) );
  nand_x1_sg U48008 ( .A(n20727), .B(n20728), .X(n20725) );
  nand_x1_sg U48009 ( .A(n5597), .B(n20729), .X(n20728) );
  nand_x1_sg U48010 ( .A(n19276), .B(n19277), .X(n19274) );
  nand_x1_sg U48011 ( .A(n5446), .B(n19278), .X(n19277) );
  nand_x1_sg U48012 ( .A(n20257), .B(n20258), .X(n20256) );
  nand_x1_sg U48013 ( .A(n5541), .B(n20259), .X(n20258) );
  nand_x1_sg U48014 ( .A(n46169), .B(n19880), .X(n19879) );
  nand_x1_sg U48015 ( .A(n20080), .B(n20081), .X(n20078) );
  nand_x1_sg U48016 ( .A(n5522), .B(n20082), .X(n20081) );
  nor_x1_sg U48017 ( .A(n21641), .B(n21642), .X(n21640) );
  nand_x1_sg U48018 ( .A(n46187), .B(n21306), .X(n21305) );
  nand_x1_sg U48019 ( .A(n20900), .B(n20901), .X(n20899) );
  nand_x1_sg U48020 ( .A(n5617), .B(n20902), .X(n20901) );
  nand_x1_sg U48021 ( .A(n46178), .B(n20537), .X(n20536) );
  nand_x1_sg U48022 ( .A(n20720), .B(n20721), .X(n20718) );
  nand_x1_sg U48023 ( .A(n5598), .B(n20722), .X(n20721) );
  nand_x1_sg U48024 ( .A(n19444), .B(n19445), .X(n19443) );
  nand_x1_sg U48025 ( .A(n5466), .B(n19446), .X(n19445) );
  nand_x1_sg U48026 ( .A(n20250), .B(n20251), .X(n20249) );
  nand_x1_sg U48027 ( .A(n5542), .B(n20252), .X(n20251) );
  nand_x1_sg U48028 ( .A(n46123), .B(n19875), .X(n19874) );
  nand_x1_sg U48029 ( .A(n20073), .B(n20074), .X(n20071) );
  nand_x1_sg U48030 ( .A(n5523), .B(n20075), .X(n20074) );
  nand_x1_sg U48031 ( .A(n46141), .B(n21301), .X(n21300) );
  nand_x1_sg U48032 ( .A(n20893), .B(n20894), .X(n20892) );
  nand_x1_sg U48033 ( .A(n5618), .B(n20895), .X(n20894) );
  nand_x1_sg U48034 ( .A(n46132), .B(n20532), .X(n20531) );
  nand_x1_sg U48035 ( .A(n20713), .B(n20714), .X(n20711) );
  nand_x1_sg U48036 ( .A(n5599), .B(n20715), .X(n20714) );
  nand_x1_sg U48037 ( .A(n19262), .B(n19263), .X(n19260) );
  nand_x1_sg U48038 ( .A(n5448), .B(n19264), .X(n19263) );
  nand_x1_sg U48039 ( .A(n20243), .B(n20244), .X(n20242) );
  nand_x1_sg U48040 ( .A(n5543), .B(n20245), .X(n20244) );
  nand_x1_sg U48041 ( .A(n46078), .B(n19870), .X(n19869) );
  nand_x1_sg U48042 ( .A(n20066), .B(n20067), .X(n20064) );
  nand_x1_sg U48043 ( .A(n5524), .B(n20068), .X(n20067) );
  nor_x1_sg U48044 ( .A(n21629), .B(n21630), .X(n21628) );
  nand_x1_sg U48045 ( .A(n46096), .B(n21296), .X(n21295) );
  nand_x1_sg U48046 ( .A(n20886), .B(n20887), .X(n20885) );
  nand_x1_sg U48047 ( .A(n5619), .B(n20888), .X(n20887) );
  nand_x1_sg U48048 ( .A(n46087), .B(n20527), .X(n20526) );
  nand_x1_sg U48049 ( .A(n20706), .B(n20707), .X(n20704) );
  nand_x1_sg U48050 ( .A(n5600), .B(n20708), .X(n20707) );
  nand_x1_sg U48051 ( .A(n19255), .B(n19256), .X(n19253) );
  nand_x1_sg U48052 ( .A(n5449), .B(n19257), .X(n19256) );
  nand_x1_sg U48053 ( .A(n20236), .B(n20237), .X(n20235) );
  nand_x1_sg U48054 ( .A(n5544), .B(n20238), .X(n20237) );
  nand_x1_sg U48055 ( .A(n46032), .B(n19865), .X(n19864) );
  nand_x1_sg U48056 ( .A(n20059), .B(n20060), .X(n20057) );
  nand_x1_sg U48057 ( .A(n5525), .B(n20061), .X(n20060) );
  nand_x1_sg U48058 ( .A(n46050), .B(n21291), .X(n21290) );
  nand_x1_sg U48059 ( .A(n20879), .B(n20880), .X(n20878) );
  nand_x1_sg U48060 ( .A(n5620), .B(n20881), .X(n20880) );
  nand_x1_sg U48061 ( .A(n46041), .B(n20522), .X(n20521) );
  nand_x1_sg U48062 ( .A(n20699), .B(n20700), .X(n20697) );
  nand_x1_sg U48063 ( .A(n5601), .B(n20701), .X(n20700) );
  nand_x1_sg U48064 ( .A(n19248), .B(n19249), .X(n19246) );
  nand_x1_sg U48065 ( .A(n5450), .B(n19250), .X(n19249) );
  nand_x1_sg U48066 ( .A(n20229), .B(n20230), .X(n20228) );
  nand_x1_sg U48067 ( .A(n5545), .B(n20231), .X(n20230) );
  nand_x1_sg U48068 ( .A(n45987), .B(n19860), .X(n19859) );
  nand_x1_sg U48069 ( .A(n20052), .B(n20053), .X(n20050) );
  nand_x1_sg U48070 ( .A(n5526), .B(n20054), .X(n20053) );
  nor_x1_sg U48071 ( .A(n21617), .B(n21618), .X(n21616) );
  nand_x1_sg U48072 ( .A(n46005), .B(n21286), .X(n21285) );
  nand_x1_sg U48073 ( .A(n20872), .B(n20873), .X(n20871) );
  nand_x1_sg U48074 ( .A(n5621), .B(n20874), .X(n20873) );
  nand_x1_sg U48075 ( .A(n45996), .B(n20517), .X(n20516) );
  nand_x1_sg U48076 ( .A(n20692), .B(n20693), .X(n20690) );
  nand_x1_sg U48077 ( .A(n5602), .B(n20694), .X(n20693) );
  nand_x1_sg U48078 ( .A(n19241), .B(n19242), .X(n19239) );
  nand_x1_sg U48079 ( .A(n5451), .B(n19243), .X(n19242) );
  nand_x1_sg U48080 ( .A(n20222), .B(n20223), .X(n20221) );
  nand_x1_sg U48081 ( .A(n45942), .B(n19855), .X(n19854) );
  nand_x1_sg U48082 ( .A(n20045), .B(n20046), .X(n20043) );
  nand_x1_sg U48083 ( .A(n5527), .B(n20047), .X(n20046) );
  nand_x1_sg U48084 ( .A(n45960), .B(n21281), .X(n21280) );
  nand_x1_sg U48085 ( .A(n20865), .B(n20866), .X(n20864) );
  nand_x1_sg U48086 ( .A(n45951), .B(n20512), .X(n20511) );
  nand_x1_sg U48087 ( .A(n20685), .B(n20686), .X(n20683) );
  nand_x1_sg U48088 ( .A(n5603), .B(n20687), .X(n20686) );
  nor_x1_sg U48089 ( .A(n45884), .B(n19208), .X(n6671) );
  inv_x1_sg U48090 ( .A(n19210), .X(n45884) );
  nand_x1_sg U48091 ( .A(n45892), .B(n19643), .X(n19642) );
  nand_x1_sg U48092 ( .A(n19234), .B(n19235), .X(n19232) );
  nand_x1_sg U48093 ( .A(n45899), .B(n20216), .X(n20215) );
  nand_x1_sg U48094 ( .A(n20038), .B(n20039), .X(n20036) );
  nand_x1_sg U48095 ( .A(n19849), .B(n45895), .X(n19847) );
  nand_x1_sg U48096 ( .A(n45902), .B(n20376), .X(n20375) );
  nand_x1_sg U48097 ( .A(n21448), .B(n21449), .X(n21446) );
  nand_x1_sg U48098 ( .A(n5680), .B(n21450), .X(n21449) );
  nor_x1_sg U48099 ( .A(n21605), .B(n21606), .X(n21604) );
  nand_x4_sg U48100 ( .A(out_L2[2]), .B(n21714), .X(n21713) );
  nand_x2_sg U48101 ( .A(n5700), .B(n45869), .X(n21714) );
  nand_x1_sg U48102 ( .A(n21275), .B(n45915), .X(n21273) );
  nand_x1_sg U48103 ( .A(n45909), .B(n20859), .X(n20858) );
  nand_x1_sg U48104 ( .A(n20506), .B(n45905), .X(n20504) );
  nand_x1_sg U48105 ( .A(n20678), .B(n20679), .X(n20676) );
  nand_x1_sg U48106 ( .A(n45912), .B(n21085), .X(n21084) );
  inv_x1_sg U48107 ( .A(n19228), .X(n45863) );
  nand_x1_sg U48108 ( .A(n20210), .B(n20211), .X(n20209) );
  nand_x1_sg U48109 ( .A(n21441), .B(n21442), .X(n21440) );
  nand_x1_sg U48110 ( .A(n20853), .B(n20854), .X(n20852) );
  nor_x1_sg U48111 ( .A(n19831), .B(n19832), .X(n19626) );
  nor_x1_sg U48112 ( .A(n20488), .B(n20489), .X(n20359) );
  nor_x1_sg U48113 ( .A(n21256), .B(n21257), .X(n21068) );
  inv_x1_sg U48114 ( .A(n7187), .X(n46900) );
  inv_x1_sg U48115 ( .A(n22818), .X(n46867) );
  inv_x1_sg U48116 ( .A(n7140), .X(n46875) );
  inv_x1_sg U48117 ( .A(n7254), .X(n46945) );
  nand_x1_sg U48118 ( .A(n7247), .B(n46934), .X(n7230) );
  nand_x1_sg U48119 ( .A(n7180), .B(n7181), .X(n7178) );
  nand_x1_sg U48120 ( .A(n46927), .B(n7190), .X(n7179) );
  nor_x1_sg U48121 ( .A(n7208), .B(n46917), .X(n7192) );
  inv_x1_sg U48122 ( .A(n7209), .X(n46917) );
  nor_x1_sg U48123 ( .A(n7273), .B(n7274), .X(n7244) );
  nand_x1_sg U48124 ( .A(n7269), .B(n46975), .X(n7245) );
  nand_x1_sg U48125 ( .A(n7306), .B(n46997), .X(n7292) );
  nand_x1_sg U48126 ( .A(n7325), .B(n7326), .X(n7324) );
  nand_x1_sg U48127 ( .A(n7309), .B(n46994), .X(n7326) );
  nand_x1_sg U48128 ( .A(n7355), .B(n7356), .X(n7321) );
  nand_x1_sg U48129 ( .A(n7385), .B(n7362), .X(n7383) );
  nand_x1_sg U48130 ( .A(n7446), .B(n47030), .X(n7413) );
  nand_x2_sg U48131 ( .A(n7418), .B(n7419), .X(n7412) );
  nand_x1_sg U48132 ( .A(n7475), .B(n7476), .X(n7417) );
  nor_x1_sg U48133 ( .A(n47058), .B(n7518), .X(n7512) );
  nand_x1_sg U48134 ( .A(n7567), .B(n47110), .X(n7544) );
  nand_x1_sg U48135 ( .A(n7545), .B(n7521), .X(n7543) );
  nand_x1_sg U48136 ( .A(n47051), .B(n7555), .X(n7545) );
  nand_x1_sg U48137 ( .A(n47087), .B(n7510), .X(n7484) );
  nand_x1_sg U48138 ( .A(n7485), .B(n7486), .X(n7483) );
  nand_x1_sg U48139 ( .A(n47029), .B(n7448), .X(n7486) );
  nand_x1_sg U48140 ( .A(n7045), .B(n7046), .X(n7040) );
  nand_x1_sg U48141 ( .A(n47116), .B(n6924), .X(n7046) );
  nand_x1_sg U48142 ( .A(n7041), .B(n7042), .X(n7039) );
  nand_x1_sg U48143 ( .A(n47112), .B(n7043), .X(n7042) );
  inv_x1_sg U48144 ( .A(n6981), .X(n47122) );
  nor_x1_sg U48145 ( .A(n47048), .B(n7577), .X(n6949) );
  nand_x1_sg U48146 ( .A(n23121), .B(n47139), .X(n23115) );
  inv_x1_sg U48147 ( .A(n8006), .X(n47185) );
  inv_x1_sg U48148 ( .A(n7958), .X(n47168) );
  inv_x1_sg U48149 ( .A(n8073), .X(n47236) );
  nand_x1_sg U48150 ( .A(n8066), .B(n47226), .X(n8049) );
  inv_x1_sg U48151 ( .A(n23095), .X(n47160) );
  nand_x1_sg U48152 ( .A(n7999), .B(n8000), .X(n7997) );
  nand_x1_sg U48153 ( .A(n47219), .B(n8009), .X(n7998) );
  nor_x1_sg U48154 ( .A(n8027), .B(n47209), .X(n8011) );
  inv_x1_sg U48155 ( .A(n8028), .X(n47209) );
  nor_x1_sg U48156 ( .A(n8092), .B(n8093), .X(n8063) );
  nand_x1_sg U48157 ( .A(n8088), .B(n47265), .X(n8064) );
  nand_x1_sg U48158 ( .A(n8124), .B(n47286), .X(n8110) );
  nand_x1_sg U48159 ( .A(n8143), .B(n8144), .X(n8142) );
  nand_x1_sg U48160 ( .A(n8127), .B(n47283), .X(n8144) );
  nand_x1_sg U48161 ( .A(n8173), .B(n8174), .X(n8139) );
  nand_x1_sg U48162 ( .A(n8203), .B(n8180), .X(n8201) );
  nand_x1_sg U48163 ( .A(n8264), .B(n47317), .X(n8231) );
  nand_x2_sg U48164 ( .A(n8236), .B(n8237), .X(n8230) );
  nand_x1_sg U48165 ( .A(n8293), .B(n8294), .X(n8235) );
  nor_x1_sg U48166 ( .A(n47344), .B(n8336), .X(n8330) );
  nand_x1_sg U48167 ( .A(n8385), .B(n47396), .X(n8362) );
  nand_x1_sg U48168 ( .A(n8363), .B(n8339), .X(n8361) );
  nand_x1_sg U48169 ( .A(n47338), .B(n8373), .X(n8363) );
  nand_x1_sg U48170 ( .A(n47373), .B(n8328), .X(n8302) );
  nand_x1_sg U48171 ( .A(n8303), .B(n8304), .X(n8301) );
  nand_x1_sg U48172 ( .A(n47316), .B(n8266), .X(n8304) );
  nand_x1_sg U48173 ( .A(n7863), .B(n7864), .X(n7858) );
  nand_x1_sg U48174 ( .A(n47402), .B(n7741), .X(n7864) );
  nand_x1_sg U48175 ( .A(n7859), .B(n7860), .X(n7857) );
  nand_x1_sg U48176 ( .A(n47398), .B(n7861), .X(n7860) );
  inv_x1_sg U48177 ( .A(n7798), .X(n47408) );
  nor_x1_sg U48178 ( .A(n47335), .B(n8395), .X(n7766) );
  nand_x1_sg U48179 ( .A(n23401), .B(n47424), .X(n23395) );
  inv_x1_sg U48180 ( .A(n8824), .X(n47470) );
  inv_x1_sg U48181 ( .A(n8776), .X(n47453) );
  inv_x1_sg U48182 ( .A(n8891), .X(n47521) );
  nand_x1_sg U48183 ( .A(n8884), .B(n47511), .X(n8867) );
  inv_x1_sg U48184 ( .A(n23375), .X(n47445) );
  nand_x1_sg U48185 ( .A(n8817), .B(n8818), .X(n8815) );
  nand_x1_sg U48186 ( .A(n47504), .B(n8827), .X(n8816) );
  nor_x1_sg U48187 ( .A(n8845), .B(n47494), .X(n8829) );
  inv_x1_sg U48188 ( .A(n8846), .X(n47494) );
  nor_x1_sg U48189 ( .A(n8910), .B(n8911), .X(n8881) );
  nand_x1_sg U48190 ( .A(n8906), .B(n47550), .X(n8882) );
  nand_x1_sg U48191 ( .A(n8942), .B(n47571), .X(n8928) );
  nand_x1_sg U48192 ( .A(n8961), .B(n8962), .X(n8960) );
  nand_x1_sg U48193 ( .A(n8945), .B(n47568), .X(n8962) );
  nand_x1_sg U48194 ( .A(n8991), .B(n8992), .X(n8957) );
  nand_x1_sg U48195 ( .A(n9021), .B(n8998), .X(n9019) );
  nand_x1_sg U48196 ( .A(n9082), .B(n47602), .X(n9049) );
  nand_x2_sg U48197 ( .A(n9054), .B(n9055), .X(n9048) );
  nand_x1_sg U48198 ( .A(n9111), .B(n9112), .X(n9053) );
  nor_x1_sg U48199 ( .A(n47629), .B(n9154), .X(n9148) );
  nand_x1_sg U48200 ( .A(n9203), .B(n47681), .X(n9180) );
  nand_x1_sg U48201 ( .A(n9181), .B(n9157), .X(n9179) );
  nand_x1_sg U48202 ( .A(n47623), .B(n9191), .X(n9181) );
  nand_x1_sg U48203 ( .A(n47658), .B(n9146), .X(n9120) );
  nand_x1_sg U48204 ( .A(n9121), .B(n9122), .X(n9119) );
  nand_x1_sg U48205 ( .A(n47601), .B(n9084), .X(n9122) );
  nand_x1_sg U48206 ( .A(n8681), .B(n8682), .X(n8676) );
  nand_x1_sg U48207 ( .A(n47687), .B(n8559), .X(n8682) );
  nand_x1_sg U48208 ( .A(n8677), .B(n8678), .X(n8675) );
  nand_x1_sg U48209 ( .A(n47683), .B(n8679), .X(n8678) );
  inv_x1_sg U48210 ( .A(n8616), .X(n47693) );
  nor_x1_sg U48211 ( .A(n47620), .B(n9213), .X(n8584) );
  nand_x1_sg U48212 ( .A(n23680), .B(n47709), .X(n23674) );
  inv_x1_sg U48213 ( .A(n9644), .X(n47755) );
  inv_x1_sg U48214 ( .A(n9596), .X(n47738) );
  inv_x1_sg U48215 ( .A(n9711), .X(n47806) );
  nand_x1_sg U48216 ( .A(n9704), .B(n47796), .X(n9687) );
  inv_x1_sg U48217 ( .A(n23654), .X(n47730) );
  nand_x1_sg U48218 ( .A(n9637), .B(n9638), .X(n9635) );
  nand_x1_sg U48219 ( .A(n47789), .B(n9647), .X(n9636) );
  nor_x1_sg U48220 ( .A(n9665), .B(n47779), .X(n9649) );
  inv_x1_sg U48221 ( .A(n9666), .X(n47779) );
  nor_x1_sg U48222 ( .A(n9730), .B(n9731), .X(n9701) );
  nand_x1_sg U48223 ( .A(n9726), .B(n47835), .X(n9702) );
  nand_x1_sg U48224 ( .A(n9762), .B(n47856), .X(n9748) );
  nand_x1_sg U48225 ( .A(n9781), .B(n9782), .X(n9780) );
  nand_x1_sg U48226 ( .A(n9765), .B(n47853), .X(n9782) );
  nand_x1_sg U48227 ( .A(n9811), .B(n9812), .X(n9777) );
  nand_x1_sg U48228 ( .A(n9841), .B(n9818), .X(n9839) );
  nand_x1_sg U48229 ( .A(n9902), .B(n47887), .X(n9869) );
  nand_x2_sg U48230 ( .A(n9874), .B(n9875), .X(n9868) );
  nand_x1_sg U48231 ( .A(n9931), .B(n9932), .X(n9873) );
  nor_x1_sg U48232 ( .A(n47914), .B(n9974), .X(n9968) );
  nand_x1_sg U48233 ( .A(n10023), .B(n47966), .X(n10000) );
  nand_x1_sg U48234 ( .A(n10001), .B(n9977), .X(n9999) );
  nand_x1_sg U48235 ( .A(n47908), .B(n10011), .X(n10001) );
  nand_x1_sg U48236 ( .A(n47943), .B(n9966), .X(n9940) );
  nand_x1_sg U48237 ( .A(n9941), .B(n9942), .X(n9939) );
  nand_x1_sg U48238 ( .A(n47886), .B(n9904), .X(n9942) );
  nand_x1_sg U48239 ( .A(n9501), .B(n9502), .X(n9496) );
  nand_x1_sg U48240 ( .A(n47972), .B(n9379), .X(n9502) );
  nand_x1_sg U48241 ( .A(n9497), .B(n9498), .X(n9495) );
  nand_x1_sg U48242 ( .A(n47968), .B(n9499), .X(n9498) );
  inv_x1_sg U48243 ( .A(n9436), .X(n47978) );
  nor_x1_sg U48244 ( .A(n47905), .B(n10033), .X(n9404) );
  nand_x1_sg U48245 ( .A(n23959), .B(n47994), .X(n23953) );
  inv_x1_sg U48246 ( .A(n10463), .X(n48040) );
  inv_x1_sg U48247 ( .A(n10415), .X(n48023) );
  inv_x1_sg U48248 ( .A(n10530), .X(n48091) );
  nand_x1_sg U48249 ( .A(n10523), .B(n48081), .X(n10506) );
  inv_x1_sg U48250 ( .A(n23933), .X(n48015) );
  nand_x1_sg U48251 ( .A(n10456), .B(n10457), .X(n10454) );
  nand_x1_sg U48252 ( .A(n48074), .B(n10466), .X(n10455) );
  nor_x1_sg U48253 ( .A(n10484), .B(n48064), .X(n10468) );
  inv_x1_sg U48254 ( .A(n10485), .X(n48064) );
  nor_x1_sg U48255 ( .A(n10549), .B(n10550), .X(n10520) );
  nand_x1_sg U48256 ( .A(n10545), .B(n48120), .X(n10521) );
  nand_x1_sg U48257 ( .A(n10581), .B(n48141), .X(n10567) );
  nand_x1_sg U48258 ( .A(n10600), .B(n10601), .X(n10599) );
  nand_x1_sg U48259 ( .A(n10584), .B(n48138), .X(n10601) );
  nand_x1_sg U48260 ( .A(n10630), .B(n10631), .X(n10596) );
  nand_x1_sg U48261 ( .A(n10660), .B(n10637), .X(n10658) );
  nand_x1_sg U48262 ( .A(n10721), .B(n48172), .X(n10688) );
  nand_x2_sg U48263 ( .A(n10693), .B(n10694), .X(n10687) );
  nand_x1_sg U48264 ( .A(n10750), .B(n10751), .X(n10692) );
  nor_x1_sg U48265 ( .A(n48199), .B(n10793), .X(n10787) );
  nand_x1_sg U48266 ( .A(n10842), .B(n48251), .X(n10819) );
  nand_x1_sg U48267 ( .A(n10820), .B(n10796), .X(n10818) );
  nand_x1_sg U48268 ( .A(n48193), .B(n10830), .X(n10820) );
  nand_x1_sg U48269 ( .A(n48228), .B(n10785), .X(n10759) );
  nand_x1_sg U48270 ( .A(n10760), .B(n10761), .X(n10758) );
  nand_x1_sg U48271 ( .A(n48171), .B(n10723), .X(n10761) );
  nand_x1_sg U48272 ( .A(n10320), .B(n10321), .X(n10315) );
  nand_x1_sg U48273 ( .A(n48257), .B(n10198), .X(n10321) );
  nand_x1_sg U48274 ( .A(n10316), .B(n10317), .X(n10314) );
  nand_x1_sg U48275 ( .A(n48253), .B(n10318), .X(n10317) );
  inv_x1_sg U48276 ( .A(n10255), .X(n48263) );
  nor_x1_sg U48277 ( .A(n48190), .B(n10852), .X(n10223) );
  nand_x1_sg U48278 ( .A(n24238), .B(n48279), .X(n24232) );
  inv_x1_sg U48279 ( .A(n11282), .X(n48325) );
  inv_x1_sg U48280 ( .A(n11234), .X(n48308) );
  inv_x1_sg U48281 ( .A(n11349), .X(n48376) );
  nand_x1_sg U48282 ( .A(n11342), .B(n48366), .X(n11325) );
  inv_x1_sg U48283 ( .A(n24212), .X(n48300) );
  nand_x1_sg U48284 ( .A(n11275), .B(n11276), .X(n11273) );
  nand_x1_sg U48285 ( .A(n48359), .B(n11285), .X(n11274) );
  nor_x1_sg U48286 ( .A(n11303), .B(n48349), .X(n11287) );
  inv_x1_sg U48287 ( .A(n11304), .X(n48349) );
  nor_x1_sg U48288 ( .A(n11368), .B(n11369), .X(n11339) );
  nand_x1_sg U48289 ( .A(n11364), .B(n48405), .X(n11340) );
  nand_x1_sg U48290 ( .A(n11400), .B(n48426), .X(n11386) );
  nand_x1_sg U48291 ( .A(n11419), .B(n11420), .X(n11418) );
  nand_x1_sg U48292 ( .A(n11403), .B(n48423), .X(n11420) );
  nand_x1_sg U48293 ( .A(n11449), .B(n11450), .X(n11415) );
  nand_x1_sg U48294 ( .A(n11479), .B(n11456), .X(n11477) );
  nand_x1_sg U48295 ( .A(n11540), .B(n48457), .X(n11507) );
  nand_x2_sg U48296 ( .A(n11512), .B(n11513), .X(n11506) );
  nand_x1_sg U48297 ( .A(n11569), .B(n11570), .X(n11511) );
  nor_x1_sg U48298 ( .A(n48484), .B(n11612), .X(n11606) );
  nand_x1_sg U48299 ( .A(n11661), .B(n48536), .X(n11638) );
  nand_x1_sg U48300 ( .A(n11639), .B(n11615), .X(n11637) );
  nand_x1_sg U48301 ( .A(n48478), .B(n11649), .X(n11639) );
  nand_x1_sg U48302 ( .A(n48513), .B(n11604), .X(n11578) );
  nand_x1_sg U48303 ( .A(n11579), .B(n11580), .X(n11577) );
  nand_x1_sg U48304 ( .A(n48456), .B(n11542), .X(n11580) );
  nand_x1_sg U48305 ( .A(n11139), .B(n11140), .X(n11134) );
  nand_x1_sg U48306 ( .A(n48542), .B(n11017), .X(n11140) );
  nand_x1_sg U48307 ( .A(n11135), .B(n11136), .X(n11133) );
  nand_x1_sg U48308 ( .A(n48538), .B(n11137), .X(n11136) );
  inv_x1_sg U48309 ( .A(n11074), .X(n48548) );
  nor_x1_sg U48310 ( .A(n48475), .B(n11671), .X(n11042) );
  nand_x1_sg U48311 ( .A(n24517), .B(n48564), .X(n24511) );
  inv_x1_sg U48312 ( .A(n12101), .X(n48610) );
  inv_x1_sg U48313 ( .A(n12053), .X(n48593) );
  inv_x1_sg U48314 ( .A(n12168), .X(n48661) );
  nand_x1_sg U48315 ( .A(n12161), .B(n48651), .X(n12144) );
  inv_x1_sg U48316 ( .A(n24491), .X(n48585) );
  nand_x1_sg U48317 ( .A(n12094), .B(n12095), .X(n12092) );
  nand_x1_sg U48318 ( .A(n48644), .B(n12104), .X(n12093) );
  nor_x1_sg U48319 ( .A(n12122), .B(n48634), .X(n12106) );
  inv_x1_sg U48320 ( .A(n12123), .X(n48634) );
  nor_x1_sg U48321 ( .A(n12187), .B(n12188), .X(n12158) );
  nand_x1_sg U48322 ( .A(n12183), .B(n48690), .X(n12159) );
  nand_x1_sg U48323 ( .A(n12219), .B(n48711), .X(n12205) );
  nand_x1_sg U48324 ( .A(n12238), .B(n12239), .X(n12237) );
  nand_x1_sg U48325 ( .A(n12222), .B(n48708), .X(n12239) );
  nand_x1_sg U48326 ( .A(n12268), .B(n12269), .X(n12234) );
  nand_x1_sg U48327 ( .A(n12298), .B(n12275), .X(n12296) );
  nand_x1_sg U48328 ( .A(n12359), .B(n48742), .X(n12326) );
  nand_x2_sg U48329 ( .A(n12331), .B(n12332), .X(n12325) );
  nand_x1_sg U48330 ( .A(n12388), .B(n12389), .X(n12330) );
  nor_x1_sg U48331 ( .A(n48769), .B(n12431), .X(n12425) );
  nand_x1_sg U48332 ( .A(n12480), .B(n48821), .X(n12457) );
  nand_x1_sg U48333 ( .A(n12458), .B(n12434), .X(n12456) );
  nand_x1_sg U48334 ( .A(n48763), .B(n12468), .X(n12458) );
  nand_x1_sg U48335 ( .A(n48798), .B(n12423), .X(n12397) );
  nand_x1_sg U48336 ( .A(n12398), .B(n12399), .X(n12396) );
  nand_x1_sg U48337 ( .A(n48741), .B(n12361), .X(n12399) );
  nand_x1_sg U48338 ( .A(n11958), .B(n11959), .X(n11953) );
  nand_x1_sg U48339 ( .A(n48827), .B(n11836), .X(n11959) );
  nand_x1_sg U48340 ( .A(n11954), .B(n11955), .X(n11952) );
  nand_x1_sg U48341 ( .A(n48823), .B(n11956), .X(n11955) );
  inv_x1_sg U48342 ( .A(n11893), .X(n48833) );
  nor_x1_sg U48343 ( .A(n48760), .B(n12490), .X(n11861) );
  nand_x1_sg U48344 ( .A(n24795), .B(n48849), .X(n24789) );
  inv_x1_sg U48345 ( .A(n12920), .X(n48896) );
  inv_x1_sg U48346 ( .A(n12872), .X(n48879) );
  inv_x1_sg U48347 ( .A(n12987), .X(n48947) );
  nand_x1_sg U48348 ( .A(n12980), .B(n48937), .X(n12963) );
  nand_x1_sg U48349 ( .A(n12913), .B(n12914), .X(n12911) );
  nand_x1_sg U48350 ( .A(n48930), .B(n12923), .X(n12912) );
  nor_x1_sg U48351 ( .A(n12941), .B(n48920), .X(n12925) );
  inv_x1_sg U48352 ( .A(n12942), .X(n48920) );
  nor_x1_sg U48353 ( .A(n13006), .B(n13007), .X(n12977) );
  nand_x1_sg U48354 ( .A(n13002), .B(n48976), .X(n12978) );
  nand_x1_sg U48355 ( .A(n13038), .B(n48997), .X(n13024) );
  nand_x1_sg U48356 ( .A(n13057), .B(n13058), .X(n13056) );
  nand_x1_sg U48357 ( .A(n13041), .B(n48994), .X(n13058) );
  nand_x1_sg U48358 ( .A(n13087), .B(n13088), .X(n13053) );
  nand_x1_sg U48359 ( .A(n13117), .B(n13094), .X(n13115) );
  nand_x1_sg U48360 ( .A(n13178), .B(n49028), .X(n13145) );
  nand_x2_sg U48361 ( .A(n13150), .B(n13151), .X(n13144) );
  nand_x1_sg U48362 ( .A(n13207), .B(n13208), .X(n13149) );
  nor_x1_sg U48363 ( .A(n49056), .B(n13250), .X(n13244) );
  nand_x1_sg U48364 ( .A(n13299), .B(n49108), .X(n13276) );
  nand_x1_sg U48365 ( .A(n13277), .B(n13253), .X(n13275) );
  nand_x1_sg U48366 ( .A(n49049), .B(n13287), .X(n13277) );
  nand_x1_sg U48367 ( .A(n49085), .B(n13242), .X(n13216) );
  nand_x1_sg U48368 ( .A(n13217), .B(n13218), .X(n13215) );
  nand_x1_sg U48369 ( .A(n49027), .B(n13180), .X(n13218) );
  nand_x1_sg U48370 ( .A(n12777), .B(n12778), .X(n12772) );
  nand_x1_sg U48371 ( .A(n49114), .B(n12655), .X(n12778) );
  nand_x1_sg U48372 ( .A(n12773), .B(n12774), .X(n12771) );
  nand_x1_sg U48373 ( .A(n49110), .B(n12775), .X(n12774) );
  inv_x1_sg U48374 ( .A(n12712), .X(n49120) );
  nor_x1_sg U48375 ( .A(n49046), .B(n13309), .X(n12680) );
  nand_x1_sg U48376 ( .A(n25074), .B(n49136), .X(n25068) );
  inv_x1_sg U48377 ( .A(n13739), .X(n49183) );
  inv_x1_sg U48378 ( .A(n13691), .X(n49166) );
  inv_x1_sg U48379 ( .A(n13806), .X(n49234) );
  nand_x1_sg U48380 ( .A(n13799), .B(n49224), .X(n13782) );
  inv_x1_sg U48381 ( .A(n25048), .X(n49158) );
  nand_x1_sg U48382 ( .A(n13732), .B(n13733), .X(n13730) );
  nand_x1_sg U48383 ( .A(n49217), .B(n13742), .X(n13731) );
  nor_x1_sg U48384 ( .A(n13760), .B(n49207), .X(n13744) );
  inv_x1_sg U48385 ( .A(n13761), .X(n49207) );
  nor_x1_sg U48386 ( .A(n13825), .B(n13826), .X(n13796) );
  nand_x1_sg U48387 ( .A(n13821), .B(n49263), .X(n13797) );
  nand_x1_sg U48388 ( .A(n13857), .B(n49284), .X(n13843) );
  nand_x1_sg U48389 ( .A(n13876), .B(n13877), .X(n13875) );
  nand_x1_sg U48390 ( .A(n13860), .B(n49281), .X(n13877) );
  nand_x1_sg U48391 ( .A(n13906), .B(n13907), .X(n13872) );
  nand_x1_sg U48392 ( .A(n13936), .B(n13913), .X(n13934) );
  nand_x1_sg U48393 ( .A(n13997), .B(n49315), .X(n13964) );
  nand_x2_sg U48394 ( .A(n13969), .B(n13970), .X(n13963) );
  nand_x1_sg U48395 ( .A(n14026), .B(n14027), .X(n13968) );
  nor_x1_sg U48396 ( .A(n49342), .B(n14069), .X(n14063) );
  nand_x1_sg U48397 ( .A(n14118), .B(n49394), .X(n14095) );
  nand_x1_sg U48398 ( .A(n14096), .B(n14072), .X(n14094) );
  nand_x1_sg U48399 ( .A(n49336), .B(n14106), .X(n14096) );
  nand_x1_sg U48400 ( .A(n49371), .B(n14061), .X(n14035) );
  nand_x1_sg U48401 ( .A(n14036), .B(n14037), .X(n14034) );
  nand_x1_sg U48402 ( .A(n49314), .B(n13999), .X(n14037) );
  nand_x1_sg U48403 ( .A(n13596), .B(n13597), .X(n13591) );
  nand_x1_sg U48404 ( .A(n49400), .B(n13474), .X(n13597) );
  nand_x1_sg U48405 ( .A(n13592), .B(n13593), .X(n13590) );
  nand_x1_sg U48406 ( .A(n49396), .B(n13594), .X(n13593) );
  inv_x1_sg U48407 ( .A(n13531), .X(n49406) );
  nor_x1_sg U48408 ( .A(n49333), .B(n14128), .X(n13499) );
  nand_x1_sg U48409 ( .A(n25353), .B(n49422), .X(n25347) );
  inv_x1_sg U48410 ( .A(n14558), .X(n49469) );
  inv_x1_sg U48411 ( .A(n14510), .X(n49452) );
  inv_x1_sg U48412 ( .A(n14625), .X(n49520) );
  nand_x1_sg U48413 ( .A(n14618), .B(n49510), .X(n14601) );
  inv_x1_sg U48414 ( .A(n25327), .X(n49444) );
  nand_x1_sg U48415 ( .A(n14551), .B(n14552), .X(n14549) );
  nand_x1_sg U48416 ( .A(n49503), .B(n14561), .X(n14550) );
  nor_x1_sg U48417 ( .A(n14579), .B(n49493), .X(n14563) );
  inv_x1_sg U48418 ( .A(n14580), .X(n49493) );
  nor_x1_sg U48419 ( .A(n14644), .B(n14645), .X(n14615) );
  nand_x1_sg U48420 ( .A(n14640), .B(n49549), .X(n14616) );
  nand_x1_sg U48421 ( .A(n14676), .B(n49570), .X(n14662) );
  nand_x1_sg U48422 ( .A(n14695), .B(n14696), .X(n14694) );
  nand_x1_sg U48423 ( .A(n14679), .B(n49567), .X(n14696) );
  nand_x1_sg U48424 ( .A(n14725), .B(n14726), .X(n14691) );
  nand_x1_sg U48425 ( .A(n14755), .B(n14732), .X(n14753) );
  nand_x1_sg U48426 ( .A(n14816), .B(n49601), .X(n14783) );
  nand_x2_sg U48427 ( .A(n14788), .B(n14789), .X(n14782) );
  nand_x1_sg U48428 ( .A(n14845), .B(n14846), .X(n14787) );
  nor_x1_sg U48429 ( .A(n49628), .B(n14888), .X(n14882) );
  nand_x1_sg U48430 ( .A(n14937), .B(n49680), .X(n14914) );
  nand_x1_sg U48431 ( .A(n14915), .B(n14891), .X(n14913) );
  nand_x1_sg U48432 ( .A(n49622), .B(n14925), .X(n14915) );
  nand_x1_sg U48433 ( .A(n49657), .B(n14880), .X(n14854) );
  nand_x1_sg U48434 ( .A(n14855), .B(n14856), .X(n14853) );
  nand_x1_sg U48435 ( .A(n49600), .B(n14818), .X(n14856) );
  nand_x1_sg U48436 ( .A(n14415), .B(n14416), .X(n14410) );
  nand_x1_sg U48437 ( .A(n49686), .B(n14293), .X(n14416) );
  nand_x1_sg U48438 ( .A(n14411), .B(n14412), .X(n14409) );
  nand_x1_sg U48439 ( .A(n49682), .B(n14413), .X(n14412) );
  inv_x1_sg U48440 ( .A(n14350), .X(n49692) );
  nor_x1_sg U48441 ( .A(n49619), .B(n14947), .X(n14318) );
  nand_x1_sg U48442 ( .A(n25632), .B(n49708), .X(n25626) );
  inv_x1_sg U48443 ( .A(n15377), .X(n49755) );
  inv_x1_sg U48444 ( .A(n15329), .X(n49737) );
  inv_x1_sg U48445 ( .A(n15444), .X(n49806) );
  nand_x1_sg U48446 ( .A(n15437), .B(n49796), .X(n15420) );
  inv_x1_sg U48447 ( .A(n25606), .X(n49729) );
  nand_x1_sg U48448 ( .A(n15370), .B(n15371), .X(n15368) );
  nand_x1_sg U48449 ( .A(n49789), .B(n15380), .X(n15369) );
  nor_x1_sg U48450 ( .A(n15398), .B(n49779), .X(n15382) );
  inv_x1_sg U48451 ( .A(n15399), .X(n49779) );
  nor_x1_sg U48452 ( .A(n15463), .B(n15464), .X(n15434) );
  nand_x1_sg U48453 ( .A(n15459), .B(n49835), .X(n15435) );
  nand_x1_sg U48454 ( .A(n15495), .B(n49856), .X(n15481) );
  nand_x1_sg U48455 ( .A(n15514), .B(n15515), .X(n15513) );
  nand_x1_sg U48456 ( .A(n15498), .B(n49853), .X(n15515) );
  nand_x1_sg U48457 ( .A(n15544), .B(n15545), .X(n15510) );
  nand_x1_sg U48458 ( .A(n15574), .B(n15551), .X(n15572) );
  nand_x1_sg U48459 ( .A(n15635), .B(n49887), .X(n15602) );
  nand_x2_sg U48460 ( .A(n15607), .B(n15608), .X(n15601) );
  nand_x1_sg U48461 ( .A(n15664), .B(n15665), .X(n15606) );
  nor_x1_sg U48462 ( .A(n49914), .B(n15707), .X(n15701) );
  nand_x1_sg U48463 ( .A(n15756), .B(n49966), .X(n15733) );
  nand_x1_sg U48464 ( .A(n15734), .B(n15710), .X(n15732) );
  nand_x1_sg U48465 ( .A(n49908), .B(n15744), .X(n15734) );
  nand_x1_sg U48466 ( .A(n49943), .B(n15699), .X(n15673) );
  nand_x1_sg U48467 ( .A(n15674), .B(n15675), .X(n15672) );
  nand_x1_sg U48468 ( .A(n49886), .B(n15637), .X(n15675) );
  nand_x1_sg U48469 ( .A(n15234), .B(n15235), .X(n15229) );
  nand_x1_sg U48470 ( .A(n49972), .B(n15112), .X(n15235) );
  nand_x1_sg U48471 ( .A(n15230), .B(n15231), .X(n15228) );
  nand_x1_sg U48472 ( .A(n49968), .B(n15232), .X(n15231) );
  inv_x1_sg U48473 ( .A(n15169), .X(n49978) );
  nor_x1_sg U48474 ( .A(n49905), .B(n15766), .X(n15137) );
  nand_x1_sg U48475 ( .A(n25909), .B(n49994), .X(n25903) );
  inv_x1_sg U48476 ( .A(n16196), .X(n50041) );
  inv_x1_sg U48477 ( .A(n16148), .X(n50024) );
  inv_x1_sg U48478 ( .A(n16263), .X(n50092) );
  nand_x1_sg U48479 ( .A(n16256), .B(n50082), .X(n16239) );
  inv_x1_sg U48480 ( .A(n25883), .X(n50016) );
  nand_x1_sg U48481 ( .A(n16189), .B(n16190), .X(n16187) );
  nand_x1_sg U48482 ( .A(n50075), .B(n16199), .X(n16188) );
  nor_x1_sg U48483 ( .A(n16217), .B(n50065), .X(n16201) );
  inv_x1_sg U48484 ( .A(n16218), .X(n50065) );
  nor_x1_sg U48485 ( .A(n16282), .B(n16283), .X(n16253) );
  nand_x1_sg U48486 ( .A(n16278), .B(n50121), .X(n16254) );
  nand_x1_sg U48487 ( .A(n16314), .B(n50142), .X(n16300) );
  nand_x1_sg U48488 ( .A(n16333), .B(n16334), .X(n16332) );
  nand_x1_sg U48489 ( .A(n16317), .B(n50139), .X(n16334) );
  nand_x1_sg U48490 ( .A(n16363), .B(n16364), .X(n16329) );
  nand_x1_sg U48491 ( .A(n16393), .B(n16370), .X(n16391) );
  nand_x1_sg U48492 ( .A(n16454), .B(n50173), .X(n16421) );
  nand_x2_sg U48493 ( .A(n16426), .B(n16427), .X(n16420) );
  nand_x1_sg U48494 ( .A(n16483), .B(n16484), .X(n16425) );
  nor_x1_sg U48495 ( .A(n50200), .B(n16526), .X(n16520) );
  nand_x1_sg U48496 ( .A(n16575), .B(n50252), .X(n16552) );
  nand_x1_sg U48497 ( .A(n16553), .B(n16529), .X(n16551) );
  nand_x1_sg U48498 ( .A(n50194), .B(n16563), .X(n16553) );
  nand_x1_sg U48499 ( .A(n50229), .B(n16518), .X(n16492) );
  nand_x1_sg U48500 ( .A(n16493), .B(n16494), .X(n16491) );
  nand_x1_sg U48501 ( .A(n50172), .B(n16456), .X(n16494) );
  nand_x1_sg U48502 ( .A(n16053), .B(n16054), .X(n16048) );
  nand_x1_sg U48503 ( .A(n50258), .B(n15931), .X(n16054) );
  nand_x1_sg U48504 ( .A(n16049), .B(n16050), .X(n16047) );
  nand_x1_sg U48505 ( .A(n50254), .B(n16051), .X(n16050) );
  inv_x1_sg U48506 ( .A(n15988), .X(n50264) );
  nor_x1_sg U48507 ( .A(n50191), .B(n16585), .X(n15956) );
  inv_x1_sg U48508 ( .A(n17012), .X(n50333) );
  inv_x1_sg U48509 ( .A(n16965), .X(n50309) );
  inv_x1_sg U48510 ( .A(n17079), .X(n50377) );
  nand_x1_sg U48511 ( .A(n17072), .B(n50367), .X(n17055) );
  nand_x1_sg U48512 ( .A(n17005), .B(n17006), .X(n17003) );
  nand_x1_sg U48513 ( .A(n50360), .B(n17015), .X(n17004) );
  nor_x1_sg U48514 ( .A(n17033), .B(n50350), .X(n17017) );
  inv_x1_sg U48515 ( .A(n17034), .X(n50350) );
  nor_x1_sg U48516 ( .A(n17098), .B(n17099), .X(n17069) );
  nand_x1_sg U48517 ( .A(n17094), .B(n50406), .X(n17070) );
  nand_x1_sg U48518 ( .A(n17150), .B(n17151), .X(n17149) );
  nand_x1_sg U48519 ( .A(n17134), .B(n50424), .X(n17151) );
  nand_x1_sg U48520 ( .A(n17180), .B(n17181), .X(n17146) );
  nand_x1_sg U48521 ( .A(n17210), .B(n17187), .X(n17208) );
  nand_x1_sg U48522 ( .A(n17223), .B(n17224), .X(n17209) );
  nand_x1_sg U48523 ( .A(n17271), .B(n50458), .X(n17238) );
  nand_x2_sg U48524 ( .A(n17243), .B(n17244), .X(n17237) );
  nand_x1_sg U48525 ( .A(n17300), .B(n17301), .X(n17242) );
  nor_x1_sg U48526 ( .A(n50485), .B(n17343), .X(n17337) );
  nand_x1_sg U48527 ( .A(n17392), .B(n50537), .X(n17369) );
  nand_x1_sg U48528 ( .A(n17370), .B(n17346), .X(n17368) );
  nand_x1_sg U48529 ( .A(n50479), .B(n17380), .X(n17370) );
  nand_x1_sg U48530 ( .A(n50514), .B(n17335), .X(n17309) );
  nand_x1_sg U48531 ( .A(n17310), .B(n17311), .X(n17308) );
  nand_x1_sg U48532 ( .A(n50457), .B(n17273), .X(n17311) );
  nand_x1_sg U48533 ( .A(n16872), .B(n16873), .X(n16867) );
  nand_x1_sg U48534 ( .A(n50543), .B(n16748), .X(n16873) );
  nand_x1_sg U48535 ( .A(n16868), .B(n16869), .X(n16866) );
  nand_x1_sg U48536 ( .A(n50539), .B(n16870), .X(n16869) );
  inv_x1_sg U48537 ( .A(n16805), .X(n50550) );
  nand_x1_sg U48538 ( .A(n50536), .B(n16841), .X(n16803) );
  nor_x1_sg U48539 ( .A(n50476), .B(n17402), .X(n16773) );
  nand_x1_sg U48540 ( .A(n26469), .B(n50569), .X(n26463) );
  inv_x1_sg U48541 ( .A(n17834), .X(n50615) );
  inv_x1_sg U48542 ( .A(n17786), .X(n50598) );
  inv_x1_sg U48543 ( .A(n17901), .X(n50666) );
  nand_x1_sg U48544 ( .A(n17894), .B(n50656), .X(n17877) );
  inv_x1_sg U48545 ( .A(n26443), .X(n50590) );
  nand_x1_sg U48546 ( .A(n17827), .B(n17828), .X(n17825) );
  nand_x1_sg U48547 ( .A(n50649), .B(n17837), .X(n17826) );
  nor_x1_sg U48548 ( .A(n17855), .B(n50639), .X(n17839) );
  inv_x1_sg U48549 ( .A(n17856), .X(n50639) );
  nor_x1_sg U48550 ( .A(n17920), .B(n17921), .X(n17891) );
  nand_x1_sg U48551 ( .A(n17916), .B(n50695), .X(n17892) );
  nand_x1_sg U48552 ( .A(n17952), .B(n50716), .X(n17938) );
  nand_x1_sg U48553 ( .A(n17971), .B(n17972), .X(n17970) );
  nand_x1_sg U48554 ( .A(n17955), .B(n50713), .X(n17972) );
  nand_x1_sg U48555 ( .A(n18001), .B(n18002), .X(n17967) );
  nand_x1_sg U48556 ( .A(n18031), .B(n18008), .X(n18029) );
  nand_x1_sg U48557 ( .A(n18092), .B(n50747), .X(n18059) );
  nand_x2_sg U48558 ( .A(n18064), .B(n18065), .X(n18058) );
  nand_x1_sg U48559 ( .A(n18121), .B(n18122), .X(n18063) );
  nor_x1_sg U48560 ( .A(n50774), .B(n18164), .X(n18158) );
  nand_x1_sg U48561 ( .A(n18213), .B(n50826), .X(n18190) );
  nand_x1_sg U48562 ( .A(n18191), .B(n18167), .X(n18189) );
  nand_x1_sg U48563 ( .A(n50768), .B(n18201), .X(n18191) );
  nand_x1_sg U48564 ( .A(n50803), .B(n18156), .X(n18130) );
  nand_x1_sg U48565 ( .A(n18131), .B(n18132), .X(n18129) );
  nand_x1_sg U48566 ( .A(n50746), .B(n18094), .X(n18132) );
  nand_x1_sg U48567 ( .A(n17691), .B(n17692), .X(n17686) );
  nand_x1_sg U48568 ( .A(n50832), .B(n17569), .X(n17692) );
  nand_x1_sg U48569 ( .A(n17687), .B(n17688), .X(n17685) );
  nand_x1_sg U48570 ( .A(n50828), .B(n17689), .X(n17688) );
  inv_x1_sg U48571 ( .A(n17626), .X(n50838) );
  nor_x1_sg U48572 ( .A(n50765), .B(n18223), .X(n17594) );
  nand_x1_sg U48573 ( .A(n26747), .B(n50855), .X(n26741) );
  inv_x1_sg U48574 ( .A(n18655), .X(n50902) );
  inv_x1_sg U48575 ( .A(n18607), .X(n50885) );
  inv_x1_sg U48576 ( .A(n18722), .X(n50953) );
  nand_x1_sg U48577 ( .A(n18715), .B(n50943), .X(n18698) );
  inv_x1_sg U48578 ( .A(n26721), .X(n50877) );
  nand_x1_sg U48579 ( .A(n18648), .B(n18649), .X(n18646) );
  nand_x1_sg U48580 ( .A(n50936), .B(n18658), .X(n18647) );
  nor_x1_sg U48581 ( .A(n18676), .B(n50926), .X(n18660) );
  inv_x1_sg U48582 ( .A(n18677), .X(n50926) );
  nor_x1_sg U48583 ( .A(n18741), .B(n18742), .X(n18712) );
  nand_x1_sg U48584 ( .A(n18737), .B(n50982), .X(n18713) );
  nand_x1_sg U48585 ( .A(n18773), .B(n51003), .X(n18759) );
  nand_x1_sg U48586 ( .A(n18792), .B(n18793), .X(n18791) );
  nand_x1_sg U48587 ( .A(n18776), .B(n51000), .X(n18793) );
  nand_x1_sg U48588 ( .A(n18822), .B(n18823), .X(n18788) );
  nand_x1_sg U48589 ( .A(n18852), .B(n18829), .X(n18850) );
  nand_x1_sg U48590 ( .A(n18913), .B(n51034), .X(n18880) );
  nand_x2_sg U48591 ( .A(n18885), .B(n18886), .X(n18879) );
  nand_x1_sg U48592 ( .A(n18942), .B(n18943), .X(n18884) );
  nor_x1_sg U48593 ( .A(n51061), .B(n18985), .X(n18979) );
  nand_x1_sg U48594 ( .A(n19034), .B(n51113), .X(n19011) );
  nand_x1_sg U48595 ( .A(n19012), .B(n18988), .X(n19010) );
  nand_x1_sg U48596 ( .A(n51055), .B(n19022), .X(n19012) );
  nand_x1_sg U48597 ( .A(n51090), .B(n18977), .X(n18951) );
  nand_x1_sg U48598 ( .A(n18952), .B(n18953), .X(n18950) );
  nand_x1_sg U48599 ( .A(n51033), .B(n18915), .X(n18953) );
  nand_x1_sg U48600 ( .A(n18512), .B(n18513), .X(n18507) );
  nand_x1_sg U48601 ( .A(n51119), .B(n18390), .X(n18513) );
  nand_x1_sg U48602 ( .A(n18508), .B(n18509), .X(n18506) );
  nand_x1_sg U48603 ( .A(n51115), .B(n18510), .X(n18509) );
  inv_x1_sg U48604 ( .A(n18447), .X(n51125) );
  nor_x1_sg U48605 ( .A(n51052), .B(n19044), .X(n18415) );
  nand_x1_sg U48606 ( .A(n26883), .B(n26884), .X(n26882) );
  inv_x1_sg U48607 ( .A(n26867), .X(n45773) );
  nand_x1_sg U48608 ( .A(n45754), .B(n26844), .X(n26822) );
  inv_x1_sg U48609 ( .A(n26838), .X(n45776) );
  inv_x1_sg U48610 ( .A(n26860), .X(n45774) );
  inv_x1_sg U48611 ( .A(n26853), .X(n45775) );
  inv_x1_sg U48612 ( .A(n26874), .X(n45772) );
  nand_x1_sg U48613 ( .A(n27100), .B(n27101), .X(n27075) );
  nand_x1_sg U48614 ( .A(n27119), .B(n27120), .X(n27066) );
  nand_x1_sg U48615 ( .A(n5209), .B(n26872), .X(n27120) );
  nand_x1_sg U48616 ( .A(n27113), .B(n27114), .X(n27069) );
  nand_x1_sg U48617 ( .A(n5228), .B(n26865), .X(n27114) );
  nand_x1_sg U48618 ( .A(n27131), .B(n27132), .X(n27060) );
  nand_x1_sg U48619 ( .A(n5171), .B(n26886), .X(n27132) );
  nand_x1_sg U48620 ( .A(n27107), .B(n27108), .X(n27072) );
  nand_x1_sg U48621 ( .A(n5247), .B(n26858), .X(n27108) );
  nand_x1_sg U48622 ( .A(n27125), .B(n27126), .X(n27063) );
  nand_x1_sg U48623 ( .A(n5190), .B(n26879), .X(n27126) );
  nand_x1_sg U48624 ( .A(n45667), .B(n27330), .X(n27305) );
  nand_x1_sg U48625 ( .A(n27349), .B(n27350), .X(n27296) );
  nand_x1_sg U48626 ( .A(n5210), .B(n27124), .X(n27350) );
  nand_x1_sg U48627 ( .A(n27343), .B(n27344), .X(n27299) );
  nand_x1_sg U48628 ( .A(n5229), .B(n27118), .X(n27344) );
  nand_x1_sg U48629 ( .A(n27361), .B(n27362), .X(n27290) );
  nand_x1_sg U48630 ( .A(n5172), .B(n27136), .X(n27362) );
  nand_x1_sg U48631 ( .A(n27337), .B(n27338), .X(n27302) );
  nand_x1_sg U48632 ( .A(n5248), .B(n27112), .X(n27338) );
  nand_x1_sg U48633 ( .A(n27355), .B(n27356), .X(n27293) );
  nand_x1_sg U48634 ( .A(n5191), .B(n27130), .X(n27356) );
  nand_x1_sg U48635 ( .A(n45623), .B(n27543), .X(n27518) );
  nand_x1_sg U48636 ( .A(n27562), .B(n27563), .X(n27509) );
  nand_x1_sg U48637 ( .A(n5211), .B(n27354), .X(n27563) );
  nand_x1_sg U48638 ( .A(n27556), .B(n27557), .X(n27512) );
  nand_x1_sg U48639 ( .A(n5230), .B(n27348), .X(n27557) );
  nand_x1_sg U48640 ( .A(n27285), .B(n27286), .X(n27284) );
  nand_x1_sg U48641 ( .A(n5173), .B(n27287), .X(n27286) );
  nand_x1_sg U48642 ( .A(n27550), .B(n27551), .X(n27515) );
  nand_x1_sg U48643 ( .A(n5249), .B(n27342), .X(n27551) );
  nand_x1_sg U48644 ( .A(n27568), .B(n27569), .X(n27506) );
  nand_x1_sg U48645 ( .A(n5192), .B(n27360), .X(n27569) );
  nand_x1_sg U48646 ( .A(n27756), .B(n27757), .X(n27703) );
  nand_x1_sg U48647 ( .A(n5212), .B(n27567), .X(n27757) );
  nand_x1_sg U48648 ( .A(n45579), .B(n27737), .X(n27712) );
  nand_x1_sg U48649 ( .A(n27750), .B(n27751), .X(n27706) );
  nand_x1_sg U48650 ( .A(n5231), .B(n27561), .X(n27751) );
  nand_x1_sg U48651 ( .A(n27279), .B(n27280), .X(n27278) );
  nand_x1_sg U48652 ( .A(n5174), .B(n27281), .X(n27280) );
  nand_x1_sg U48653 ( .A(n27744), .B(n27745), .X(n27709) );
  nand_x1_sg U48654 ( .A(n5250), .B(n27555), .X(n27745) );
  nand_x1_sg U48655 ( .A(n27501), .B(n27502), .X(n27500) );
  nand_x1_sg U48656 ( .A(n5193), .B(n27503), .X(n27502) );
  nand_x1_sg U48657 ( .A(n27698), .B(n27699), .X(n27697) );
  nand_x1_sg U48658 ( .A(n5213), .B(n27700), .X(n27699) );
  nand_x1_sg U48659 ( .A(n45534), .B(n27914), .X(n27889) );
  nand_x1_sg U48660 ( .A(n27927), .B(n27928), .X(n27883) );
  nand_x1_sg U48661 ( .A(n5232), .B(n27755), .X(n27928) );
  nand_x1_sg U48662 ( .A(n27273), .B(n27274), .X(n27272) );
  nand_x1_sg U48663 ( .A(n5175), .B(n27275), .X(n27274) );
  nand_x1_sg U48664 ( .A(n27921), .B(n27922), .X(n27886) );
  nand_x1_sg U48665 ( .A(n5251), .B(n27749), .X(n27922) );
  nand_x1_sg U48666 ( .A(n27495), .B(n27496), .X(n27494) );
  nand_x1_sg U48667 ( .A(n5194), .B(n27497), .X(n27496) );
  nand_x1_sg U48668 ( .A(n27692), .B(n27693), .X(n27691) );
  nand_x1_sg U48669 ( .A(n5214), .B(n27694), .X(n27693) );
  nand_x1_sg U48670 ( .A(n45490), .B(n28076), .X(n28051) );
  nand_x1_sg U48671 ( .A(n27878), .B(n27879), .X(n27877) );
  nand_x1_sg U48672 ( .A(n5233), .B(n27880), .X(n27879) );
  nand_x1_sg U48673 ( .A(n27267), .B(n27268), .X(n27266) );
  nand_x1_sg U48674 ( .A(n5176), .B(n27269), .X(n27268) );
  nand_x1_sg U48675 ( .A(n28083), .B(n28084), .X(n28048) );
  nand_x1_sg U48676 ( .A(n5252), .B(n27926), .X(n28084) );
  nand_x1_sg U48677 ( .A(n27489), .B(n27490), .X(n27488) );
  nand_x1_sg U48678 ( .A(n5195), .B(n27491), .X(n27490) );
  nand_x1_sg U48679 ( .A(n27686), .B(n27687), .X(n27685) );
  nand_x1_sg U48680 ( .A(n5215), .B(n27688), .X(n27687) );
  nand_x1_sg U48681 ( .A(n45466), .B(n28211), .X(n28186) );
  nand_x1_sg U48682 ( .A(n27872), .B(n27873), .X(n27871) );
  nand_x1_sg U48683 ( .A(n5234), .B(n27874), .X(n27873) );
  nand_x1_sg U48684 ( .A(n27261), .B(n27262), .X(n27260) );
  nand_x1_sg U48685 ( .A(n5177), .B(n27263), .X(n27262) );
  nand_x1_sg U48686 ( .A(n28043), .B(n28044), .X(n28042) );
  nand_x1_sg U48687 ( .A(n5253), .B(n28045), .X(n28044) );
  nand_x1_sg U48688 ( .A(n27483), .B(n27484), .X(n27482) );
  nand_x1_sg U48689 ( .A(n5196), .B(n27485), .X(n27484) );
  nand_x1_sg U48690 ( .A(n27680), .B(n27681), .X(n27679) );
  nand_x1_sg U48691 ( .A(n5216), .B(n27682), .X(n27681) );
  nand_x1_sg U48692 ( .A(n45422), .B(n28182), .X(n28181) );
  nand_x1_sg U48693 ( .A(n27866), .B(n27867), .X(n27865) );
  nand_x1_sg U48694 ( .A(n5235), .B(n27868), .X(n27867) );
  nand_x1_sg U48695 ( .A(n27255), .B(n27256), .X(n27254) );
  nand_x1_sg U48696 ( .A(n5178), .B(n27257), .X(n27256) );
  nand_x1_sg U48697 ( .A(n28037), .B(n28038), .X(n28036) );
  nand_x1_sg U48698 ( .A(n5254), .B(n28039), .X(n28038) );
  nand_x1_sg U48699 ( .A(n27477), .B(n27478), .X(n27476) );
  nand_x1_sg U48700 ( .A(n5197), .B(n27479), .X(n27478) );
  nand_x1_sg U48701 ( .A(n27674), .B(n27675), .X(n27673) );
  nand_x1_sg U48702 ( .A(n5217), .B(n27676), .X(n27675) );
  nand_x1_sg U48703 ( .A(n45376), .B(n28176), .X(n28175) );
  nand_x1_sg U48704 ( .A(n28313), .B(n28314), .X(n28311) );
  nand_x1_sg U48705 ( .A(n5293), .B(n28315), .X(n28314) );
  nand_x1_sg U48706 ( .A(n27860), .B(n27861), .X(n27859) );
  nand_x1_sg U48707 ( .A(n5236), .B(n27862), .X(n27861) );
  nand_x1_sg U48708 ( .A(n27249), .B(n27250), .X(n27248) );
  nand_x1_sg U48709 ( .A(n5179), .B(n27251), .X(n27250) );
  nand_x1_sg U48710 ( .A(n28031), .B(n28032), .X(n28030) );
  nand_x1_sg U48711 ( .A(n5255), .B(n28033), .X(n28032) );
  nand_x1_sg U48712 ( .A(n27471), .B(n27472), .X(n27470) );
  nand_x1_sg U48713 ( .A(n5198), .B(n27473), .X(n27472) );
  nand_x1_sg U48714 ( .A(n27668), .B(n27669), .X(n27667) );
  nand_x1_sg U48715 ( .A(n5218), .B(n27670), .X(n27669) );
  nand_x1_sg U48716 ( .A(n45331), .B(n28171), .X(n28170) );
  nand_x1_sg U48717 ( .A(n28307), .B(n28308), .X(n28305) );
  nand_x1_sg U48718 ( .A(n5294), .B(n28309), .X(n28308) );
  nand_x1_sg U48719 ( .A(n27854), .B(n27855), .X(n27853) );
  nand_x1_sg U48720 ( .A(n5237), .B(n27856), .X(n27855) );
  nand_x1_sg U48721 ( .A(n27243), .B(n27244), .X(n27242) );
  nand_x1_sg U48722 ( .A(n5180), .B(n27245), .X(n27244) );
  nand_x1_sg U48723 ( .A(n28025), .B(n28026), .X(n28024) );
  nand_x1_sg U48724 ( .A(n5256), .B(n28027), .X(n28026) );
  nand_x1_sg U48725 ( .A(n27465), .B(n27466), .X(n27464) );
  nand_x1_sg U48726 ( .A(n5199), .B(n27467), .X(n27466) );
  nand_x1_sg U48727 ( .A(n27662), .B(n27663), .X(n27661) );
  nand_x1_sg U48728 ( .A(n5219), .B(n27664), .X(n27663) );
  nand_x1_sg U48729 ( .A(n45286), .B(n28166), .X(n28165) );
  nand_x1_sg U48730 ( .A(n28301), .B(n28302), .X(n28299) );
  nand_x1_sg U48731 ( .A(n5295), .B(n28303), .X(n28302) );
  nand_x1_sg U48732 ( .A(n27848), .B(n27849), .X(n27847) );
  nand_x1_sg U48733 ( .A(n5238), .B(n27850), .X(n27849) );
  nand_x1_sg U48734 ( .A(n27237), .B(n27238), .X(n27236) );
  nand_x1_sg U48735 ( .A(n5181), .B(n27239), .X(n27238) );
  nand_x1_sg U48736 ( .A(n28019), .B(n28020), .X(n28018) );
  nand_x1_sg U48737 ( .A(n5257), .B(n28021), .X(n28020) );
  nand_x1_sg U48738 ( .A(n27459), .B(n27460), .X(n27458) );
  nand_x1_sg U48739 ( .A(n5200), .B(n27461), .X(n27460) );
  nand_x1_sg U48740 ( .A(n27656), .B(n27657), .X(n27655) );
  nand_x1_sg U48741 ( .A(n5220), .B(n27658), .X(n27657) );
  nand_x1_sg U48742 ( .A(n45241), .B(n28161), .X(n28160) );
  nand_x1_sg U48743 ( .A(n28295), .B(n28296), .X(n28293) );
  nand_x1_sg U48744 ( .A(n5296), .B(n28297), .X(n28296) );
  nand_x1_sg U48745 ( .A(n27842), .B(n27843), .X(n27841) );
  nand_x1_sg U48746 ( .A(n5239), .B(n27844), .X(n27843) );
  nand_x1_sg U48747 ( .A(n27231), .B(n27232), .X(n27230) );
  nand_x1_sg U48748 ( .A(n5182), .B(n27233), .X(n27232) );
  nand_x1_sg U48749 ( .A(n28013), .B(n28014), .X(n28012) );
  nand_x1_sg U48750 ( .A(n5258), .B(n28015), .X(n28014) );
  nand_x1_sg U48751 ( .A(n27453), .B(n27454), .X(n27452) );
  nand_x1_sg U48752 ( .A(n5201), .B(n27455), .X(n27454) );
  nand_x1_sg U48753 ( .A(n27650), .B(n27651), .X(n27649) );
  nand_x1_sg U48754 ( .A(n5221), .B(n27652), .X(n27651) );
  nand_x1_sg U48755 ( .A(n45195), .B(n28156), .X(n28155) );
  nand_x1_sg U48756 ( .A(n28289), .B(n28290), .X(n28287) );
  nand_x1_sg U48757 ( .A(n5297), .B(n28291), .X(n28290) );
  nand_x1_sg U48758 ( .A(n27836), .B(n27837), .X(n27835) );
  nand_x1_sg U48759 ( .A(n5240), .B(n27838), .X(n27837) );
  nand_x1_sg U48760 ( .A(n27225), .B(n27226), .X(n27224) );
  nand_x1_sg U48761 ( .A(n5183), .B(n27227), .X(n27226) );
  nand_x1_sg U48762 ( .A(n28007), .B(n28008), .X(n28006) );
  nand_x1_sg U48763 ( .A(n5259), .B(n28009), .X(n28008) );
  nand_x1_sg U48764 ( .A(n27447), .B(n27448), .X(n27446) );
  nand_x1_sg U48765 ( .A(n5202), .B(n27449), .X(n27448) );
  nand_x1_sg U48766 ( .A(n27644), .B(n27645), .X(n27643) );
  nand_x1_sg U48767 ( .A(n5222), .B(n27646), .X(n27645) );
  nand_x1_sg U48768 ( .A(n45150), .B(n28151), .X(n28150) );
  nand_x1_sg U48769 ( .A(n28283), .B(n28284), .X(n28281) );
  nand_x1_sg U48770 ( .A(n5298), .B(n28285), .X(n28284) );
  nand_x1_sg U48771 ( .A(n27830), .B(n27831), .X(n27829) );
  nand_x1_sg U48772 ( .A(n5241), .B(n27832), .X(n27831) );
  nand_x1_sg U48773 ( .A(n27219), .B(n27220), .X(n27218) );
  nand_x1_sg U48774 ( .A(n5184), .B(n27221), .X(n27220) );
  nand_x1_sg U48775 ( .A(n28001), .B(n28002), .X(n28000) );
  nand_x1_sg U48776 ( .A(n5260), .B(n28003), .X(n28002) );
  nand_x1_sg U48777 ( .A(n27441), .B(n27442), .X(n27440) );
  nand_x1_sg U48778 ( .A(n5203), .B(n27443), .X(n27442) );
  nand_x1_sg U48779 ( .A(n27638), .B(n27639), .X(n27637) );
  nand_x1_sg U48780 ( .A(n5223), .B(n27640), .X(n27639) );
  nand_x1_sg U48781 ( .A(n45104), .B(n28146), .X(n28145) );
  nand_x1_sg U48782 ( .A(n28277), .B(n28278), .X(n28275) );
  nand_x1_sg U48783 ( .A(n5299), .B(n28279), .X(n28278) );
  nand_x1_sg U48784 ( .A(n27824), .B(n27825), .X(n27823) );
  nand_x1_sg U48785 ( .A(n5242), .B(n27826), .X(n27825) );
  nand_x1_sg U48786 ( .A(n27213), .B(n27214), .X(n27212) );
  nand_x1_sg U48787 ( .A(n5185), .B(n27215), .X(n27214) );
  nand_x1_sg U48788 ( .A(n27995), .B(n27996), .X(n27994) );
  nand_x1_sg U48789 ( .A(n5261), .B(n27997), .X(n27996) );
  nand_x1_sg U48790 ( .A(n27435), .B(n27436), .X(n27434) );
  nand_x1_sg U48791 ( .A(n5204), .B(n27437), .X(n27436) );
  nand_x1_sg U48792 ( .A(n27632), .B(n27633), .X(n27631) );
  nand_x1_sg U48793 ( .A(n5224), .B(n27634), .X(n27633) );
  nand_x1_sg U48794 ( .A(n27818), .B(n27819), .X(n27817) );
  nand_x1_sg U48795 ( .A(n5243), .B(n27820), .X(n27819) );
  nand_x1_sg U48796 ( .A(n27207), .B(n27208), .X(n27206) );
  nand_x1_sg U48797 ( .A(n5186), .B(n27209), .X(n27208) );
  nor_x1_sg U48798 ( .A(n45080), .B(n28137), .X(n27987) );
  inv_x1_sg U48799 ( .A(n28139), .X(n45080) );
  nand_x1_sg U48800 ( .A(n27989), .B(n27990), .X(n27988) );
  nand_x1_sg U48801 ( .A(n5262), .B(n27991), .X(n27990) );
  nand_x1_sg U48802 ( .A(n27429), .B(n27430), .X(n27428) );
  nand_x1_sg U48803 ( .A(n5205), .B(n27431), .X(n27430) );
  nand_x1_sg U48804 ( .A(n27626), .B(n27627), .X(n27625) );
  nand_x1_sg U48805 ( .A(n27812), .B(n27813), .X(n27811) );
  nand_x1_sg U48806 ( .A(n27201), .B(n27202), .X(n27200) );
  nor_x1_sg U48807 ( .A(n28130), .B(n28131), .X(n27980) );
  nand_x1_sg U48808 ( .A(n27982), .B(n27983), .X(n27981) );
  nand_x1_sg U48809 ( .A(n27423), .B(n27424), .X(n27422) );
  inv_x1_sg U48810 ( .A(n28125), .X(n44999) );
  inv_x1_sg U48811 ( .A(n27618), .X(n45008) );
  inv_x1_sg U48812 ( .A(n27803), .X(n45005) );
  inv_x1_sg U48813 ( .A(n27972), .X(n45002) );
  inv_x1_sg U48814 ( .A(n27414), .X(n45011) );
  nor_x1_sg U48815 ( .A(n44968), .B(n28254), .X(n28123) );
  nor_x1_sg U48816 ( .A(n28121), .B(n28122), .X(n27970) );
  nand_x1_sg U48817 ( .A(n22844), .B(n46847), .X(n22838) );
  nand_x1_sg U48818 ( .A(n22776), .B(n22777), .X(n22774) );
  nand_x1_sg U48819 ( .A(n23053), .B(n23054), .X(n23051) );
  nand_x1_sg U48820 ( .A(n23039), .B(n23040), .X(n23037) );
  nand_x1_sg U48821 ( .A(n23025), .B(n23026), .X(n23023) );
  inv_x1_sg U48822 ( .A(n22994), .X(n47414) );
  nor_x1_sg U48823 ( .A(n22989), .B(n22990), .X(n22987) );
  inv_x1_sg U48824 ( .A(n22991), .X(n47382) );
  nand_x1_sg U48825 ( .A(n23333), .B(n23334), .X(n23331) );
  nand_x1_sg U48826 ( .A(n23319), .B(n23320), .X(n23317) );
  nand_x1_sg U48827 ( .A(n23305), .B(n23306), .X(n23303) );
  inv_x1_sg U48828 ( .A(n23274), .X(n47699) );
  nor_x1_sg U48829 ( .A(n23269), .B(n23270), .X(n23267) );
  inv_x1_sg U48830 ( .A(n23271), .X(n47667) );
  nand_x1_sg U48831 ( .A(n23612), .B(n23613), .X(n23610) );
  nand_x1_sg U48832 ( .A(n23598), .B(n23599), .X(n23596) );
  nand_x1_sg U48833 ( .A(n23584), .B(n23585), .X(n23582) );
  inv_x1_sg U48834 ( .A(n23553), .X(n47984) );
  nor_x1_sg U48835 ( .A(n23548), .B(n23549), .X(n23546) );
  inv_x1_sg U48836 ( .A(n23550), .X(n47952) );
  nand_x1_sg U48837 ( .A(n23891), .B(n23892), .X(n23889) );
  nand_x1_sg U48838 ( .A(n23877), .B(n23878), .X(n23875) );
  nand_x1_sg U48839 ( .A(n23863), .B(n23864), .X(n23861) );
  inv_x1_sg U48840 ( .A(n23832), .X(n48269) );
  nor_x1_sg U48841 ( .A(n23827), .B(n23828), .X(n23825) );
  inv_x1_sg U48842 ( .A(n23829), .X(n48237) );
  nand_x1_sg U48843 ( .A(n24170), .B(n24171), .X(n24168) );
  nand_x1_sg U48844 ( .A(n24156), .B(n24157), .X(n24154) );
  nand_x1_sg U48845 ( .A(n24142), .B(n24143), .X(n24140) );
  inv_x1_sg U48846 ( .A(n24111), .X(n48554) );
  nor_x1_sg U48847 ( .A(n24106), .B(n24107), .X(n24104) );
  inv_x1_sg U48848 ( .A(n24108), .X(n48522) );
  nand_x1_sg U48849 ( .A(n24449), .B(n24450), .X(n24447) );
  nand_x1_sg U48850 ( .A(n24435), .B(n24436), .X(n24433) );
  nand_x1_sg U48851 ( .A(n24421), .B(n24422), .X(n24419) );
  inv_x1_sg U48852 ( .A(n24390), .X(n48839) );
  nor_x1_sg U48853 ( .A(n24385), .B(n24386), .X(n24383) );
  inv_x1_sg U48854 ( .A(n24387), .X(n48807) );
  inv_x1_sg U48855 ( .A(n24769), .X(n48871) );
  nand_x1_sg U48856 ( .A(n24727), .B(n24728), .X(n24725) );
  nand_x1_sg U48857 ( .A(n24713), .B(n24714), .X(n24711) );
  nand_x1_sg U48858 ( .A(n24699), .B(n24700), .X(n24697) );
  inv_x1_sg U48859 ( .A(n24668), .X(n49126) );
  nor_x1_sg U48860 ( .A(n24663), .B(n24664), .X(n24661) );
  inv_x1_sg U48861 ( .A(n24665), .X(n49094) );
  nand_x1_sg U48862 ( .A(n25006), .B(n25007), .X(n25004) );
  nand_x1_sg U48863 ( .A(n24992), .B(n24993), .X(n24990) );
  nand_x1_sg U48864 ( .A(n24978), .B(n24979), .X(n24976) );
  inv_x1_sg U48865 ( .A(n24947), .X(n49412) );
  nor_x1_sg U48866 ( .A(n24942), .B(n24943), .X(n24940) );
  inv_x1_sg U48867 ( .A(n24944), .X(n49380) );
  nand_x1_sg U48868 ( .A(n25285), .B(n25286), .X(n25283) );
  nand_x1_sg U48869 ( .A(n25271), .B(n25272), .X(n25269) );
  nand_x1_sg U48870 ( .A(n25257), .B(n25258), .X(n25255) );
  inv_x1_sg U48871 ( .A(n25226), .X(n49698) );
  nor_x1_sg U48872 ( .A(n25221), .B(n25222), .X(n25219) );
  inv_x1_sg U48873 ( .A(n25223), .X(n49666) );
  nand_x1_sg U48874 ( .A(n25564), .B(n25565), .X(n25562) );
  nand_x1_sg U48875 ( .A(n25550), .B(n25551), .X(n25548) );
  nand_x1_sg U48876 ( .A(n25536), .B(n25537), .X(n25534) );
  inv_x1_sg U48877 ( .A(n25505), .X(n49984) );
  nor_x1_sg U48878 ( .A(n25500), .B(n25501), .X(n25498) );
  inv_x1_sg U48879 ( .A(n25502), .X(n49952) );
  nand_x1_sg U48880 ( .A(n25841), .B(n25842), .X(n25839) );
  nand_x1_sg U48881 ( .A(n25827), .B(n25828), .X(n25825) );
  nand_x1_sg U48882 ( .A(n25813), .B(n25814), .X(n25811) );
  inv_x1_sg U48883 ( .A(n25782), .X(n50270) );
  nor_x1_sg U48884 ( .A(n25777), .B(n25778), .X(n25775) );
  inv_x1_sg U48885 ( .A(n25779), .X(n50238) );
  nand_x1_sg U48886 ( .A(n26115), .B(n26116), .X(n26112) );
  nand_x1_sg U48887 ( .A(n26080), .B(n26156), .X(n26071) );
  nand_x1_sg U48888 ( .A(n26401), .B(n26402), .X(n26399) );
  nand_x1_sg U48889 ( .A(n26387), .B(n26388), .X(n26385) );
  nand_x1_sg U48890 ( .A(n26373), .B(n26374), .X(n26371) );
  inv_x1_sg U48891 ( .A(n26342), .X(n50845) );
  nor_x1_sg U48892 ( .A(n26337), .B(n26338), .X(n26335) );
  inv_x1_sg U48893 ( .A(n26339), .X(n50812) );
  nand_x1_sg U48894 ( .A(n26679), .B(n26680), .X(n26677) );
  nand_x1_sg U48895 ( .A(n26665), .B(n26666), .X(n26663) );
  nand_x1_sg U48896 ( .A(n26651), .B(n26652), .X(n26649) );
  inv_x1_sg U48897 ( .A(n26620), .X(n51131) );
  nor_x1_sg U48898 ( .A(n26615), .B(n26616), .X(n26613) );
  inv_x1_sg U48899 ( .A(n26617), .X(n51099) );
  nand_x1_sg U48900 ( .A(n46607), .B(n19140), .X(n19138) );
  nor_x1_sg U48901 ( .A(n46629), .B(n19514), .X(n19510) );
  inv_x1_sg U48902 ( .A(n19516), .X(n46629) );
  nor_x1_sg U48903 ( .A(n46630), .B(n19511), .X(n19137) );
  inv_x1_sg U48904 ( .A(n19513), .X(n46630) );
  nand_x1_sg U48905 ( .A(n46610), .B(n19147), .X(n19135) );
  nand_x1_sg U48906 ( .A(n46597), .B(n19537), .X(n19524) );
  nor_x1_sg U48907 ( .A(n46628), .B(n19517), .X(n19119) );
  inv_x1_sg U48908 ( .A(n19519), .X(n46628) );
  nor_x1_sg U48909 ( .A(n46627), .B(n19520), .X(n19117) );
  inv_x1_sg U48910 ( .A(n19522), .X(n46627) );
  nor_x1_sg U48911 ( .A(n46625), .B(n19526), .X(n19123) );
  inv_x1_sg U48912 ( .A(n19529), .X(n46625) );
  inv_x1_sg U48913 ( .A(n20986), .X(n46616) );
  nand_x2_sg U48914 ( .A(out_L2[18]), .B(n20981), .X(n20980) );
  nand_x1_sg U48915 ( .A(n20983), .B(n46617), .X(n20978) );
  nor_x1_sg U48916 ( .A(n46620), .B(n20969), .X(n20568) );
  inv_x1_sg U48917 ( .A(n20971), .X(n46620) );
  nand_x1_sg U48918 ( .A(n46615), .B(n21007), .X(n20964) );
  nor_x1_sg U48919 ( .A(n46624), .B(n20576), .X(n19527) );
  inv_x1_sg U48920 ( .A(n20578), .X(n46624) );
  nor_x1_sg U48921 ( .A(n46623), .B(n20579), .X(n20574) );
  inv_x1_sg U48922 ( .A(n20582), .X(n46623) );
  nor_x1_sg U48923 ( .A(n46621), .B(n20966), .X(n20960) );
  inv_x1_sg U48924 ( .A(n20968), .X(n46621) );
  inv_x1_sg U48925 ( .A(n19331), .X(n46608) );
  nand_x1_sg U48926 ( .A(n5981), .B(n5982), .X(n5980) );
  nor_x1_sg U48927 ( .A(n21187), .B(n21188), .X(n21181) );
  nand_x1_sg U48928 ( .A(n46524), .B(n6033), .X(n6032) );
  nand_x1_sg U48929 ( .A(n19946), .B(n19947), .X(n19929) );
  nand_x1_sg U48930 ( .A(n5533), .B(n46513), .X(n19947) );
  nor_x1_sg U48931 ( .A(n46566), .B(n19922), .X(n6020) );
  inv_x1_sg U48932 ( .A(n19924), .X(n46566) );
  nand_x1_sg U48933 ( .A(n42081), .B(n21357), .X(n21352) );
  inv_x1_sg U48934 ( .A(n19936), .X(n46556) );
  nor_x1_sg U48935 ( .A(n20772), .B(n46551), .X(n6051) );
  inv_x1_sg U48936 ( .A(n20773), .X(n46551) );
  inv_x1_sg U48937 ( .A(n19319), .X(n46521) );
  nand_x1_sg U48938 ( .A(n6082), .B(n6083), .X(n6081) );
  nand_x1_sg U48939 ( .A(n5420), .B(n6084), .X(n6083) );
  nor_x1_sg U48940 ( .A(n46517), .B(n20122), .X(n6068) );
  inv_x1_sg U48941 ( .A(n20124), .X(n46517) );
  inv_x1_sg U48942 ( .A(n20130), .X(n46512) );
  nand_x1_sg U48943 ( .A(n46501), .B(n21539), .X(n21534) );
  nor_x1_sg U48944 ( .A(n20131), .B(n20132), .X(n6102) );
  nor_x1_sg U48945 ( .A(n20765), .B(n20766), .X(n6101) );
  nor_x1_sg U48946 ( .A(n19488), .B(n46478), .X(n6134) );
  inv_x1_sg U48947 ( .A(n19489), .X(n46478) );
  nand_x1_sg U48948 ( .A(n6129), .B(n6130), .X(n6128) );
  nand_x1_sg U48949 ( .A(n20311), .B(n46449), .X(n20294) );
  nand_x1_sg U48950 ( .A(n21526), .B(n21527), .X(n21524) );
  nand_x1_sg U48951 ( .A(n5668), .B(n21528), .X(n21527) );
  nor_x1_sg U48952 ( .A(n21673), .B(n21674), .X(n21523) );
  nor_x1_sg U48953 ( .A(n20758), .B(n20759), .X(n6147) );
  nand_x1_sg U48954 ( .A(n46387), .B(n6174), .X(n6173) );
  inv_x1_sg U48955 ( .A(n19308), .X(n46432) );
  nor_x1_sg U48956 ( .A(n46429), .B(n19904), .X(n6162) );
  inv_x1_sg U48957 ( .A(n19906), .X(n46429) );
  nand_x1_sg U48958 ( .A(n21519), .B(n21520), .X(n21517) );
  nand_x1_sg U48959 ( .A(n5669), .B(n21521), .X(n21520) );
  nand_x1_sg U48960 ( .A(n46416), .B(n21671), .X(n21669) );
  nor_x1_sg U48961 ( .A(n20751), .B(n20752), .X(n6193) );
  nand_x1_sg U48962 ( .A(n19303), .B(n19304), .X(n19301) );
  nand_x1_sg U48963 ( .A(n5442), .B(n19305), .X(n19304) );
  nand_x1_sg U48964 ( .A(n6221), .B(n6222), .X(n6220) );
  nand_x1_sg U48965 ( .A(n20284), .B(n20285), .X(n20282) );
  nand_x1_sg U48966 ( .A(n5537), .B(n20286), .X(n20285) );
  inv_x1_sg U48967 ( .A(n19898), .X(n46382) );
  nand_x1_sg U48968 ( .A(n21513), .B(n21514), .X(n21511) );
  nand_x1_sg U48969 ( .A(n5670), .B(n21515), .X(n21514) );
  nor_x1_sg U48970 ( .A(n21661), .B(n21662), .X(n21510) );
  nor_x1_sg U48971 ( .A(n20554), .B(n20555), .X(n6240) );
  nand_x1_sg U48972 ( .A(n46296), .B(n6267), .X(n6266) );
  nand_x1_sg U48973 ( .A(n21506), .B(n21507), .X(n21504) );
  nand_x1_sg U48974 ( .A(n5671), .B(n21508), .X(n21507) );
  nand_x1_sg U48975 ( .A(n46327), .B(n21659), .X(n21657) );
  nand_x1_sg U48976 ( .A(n46251), .B(n6312), .X(n6311) );
  nand_x1_sg U48977 ( .A(n21500), .B(n21501), .X(n21498) );
  nand_x1_sg U48978 ( .A(n5672), .B(n21502), .X(n21501) );
  nor_x1_sg U48979 ( .A(n21649), .B(n21650), .X(n21497) );
  nand_x1_sg U48980 ( .A(n46205), .B(n6356), .X(n6355) );
  nand_x1_sg U48981 ( .A(n21493), .B(n21494), .X(n21491) );
  nand_x1_sg U48982 ( .A(n5673), .B(n21495), .X(n21494) );
  nand_x1_sg U48983 ( .A(n46236), .B(n21647), .X(n21645) );
  nand_x1_sg U48984 ( .A(n46160), .B(n6401), .X(n6400) );
  nand_x1_sg U48985 ( .A(n21487), .B(n21488), .X(n21485) );
  nand_x1_sg U48986 ( .A(n5674), .B(n21489), .X(n21488) );
  nor_x1_sg U48987 ( .A(n21637), .B(n21638), .X(n21484) );
  nand_x1_sg U48988 ( .A(n19269), .B(n19270), .X(n19267) );
  nand_x1_sg U48989 ( .A(n5447), .B(n19271), .X(n19270) );
  nand_x1_sg U48990 ( .A(n46114), .B(n6445), .X(n6444) );
  nand_x1_sg U48991 ( .A(n21480), .B(n21481), .X(n21478) );
  nand_x1_sg U48992 ( .A(n5675), .B(n21482), .X(n21481) );
  nand_x1_sg U48993 ( .A(n46145), .B(n21635), .X(n21633) );
  nand_x1_sg U48994 ( .A(n46069), .B(n6490), .X(n6489) );
  nand_x1_sg U48995 ( .A(n21474), .B(n21475), .X(n21472) );
  nand_x1_sg U48996 ( .A(n5676), .B(n21476), .X(n21475) );
  nor_x1_sg U48997 ( .A(n21625), .B(n21626), .X(n21471) );
  nand_x1_sg U48998 ( .A(n46023), .B(n6534), .X(n6533) );
  nand_x1_sg U48999 ( .A(n21467), .B(n21468), .X(n21465) );
  nand_x1_sg U49000 ( .A(n5677), .B(n21469), .X(n21468) );
  nand_x1_sg U49001 ( .A(n46054), .B(n21623), .X(n21621) );
  nand_x1_sg U49002 ( .A(n45978), .B(n6579), .X(n6578) );
  nand_x1_sg U49003 ( .A(n21461), .B(n21462), .X(n21459) );
  nand_x1_sg U49004 ( .A(n5678), .B(n21463), .X(n21462) );
  nor_x1_sg U49005 ( .A(n21613), .B(n21614), .X(n21458) );
  nand_x1_sg U49006 ( .A(n45933), .B(n6623), .X(n6622) );
  nand_x1_sg U49007 ( .A(n21454), .B(n21455), .X(n21452) );
  nand_x1_sg U49008 ( .A(n5679), .B(n21456), .X(n21455) );
  nand_x1_sg U49009 ( .A(n42076), .B(n21611), .X(n21609) );
  nand_x1_sg U49010 ( .A(n6669), .B(n45885), .X(n6668) );
  nor_x1_sg U49011 ( .A(n19640), .B(n19641), .X(n6674) );
  inv_x1_sg U49012 ( .A(n19848), .X(n45927) );
  nor_x1_sg U49013 ( .A(n20373), .B(n20374), .X(n6659) );
  nor_x1_sg U49014 ( .A(n21601), .B(n21602), .X(n21445) );
  inv_x1_sg U49015 ( .A(n21274), .X(n45921) );
  inv_x1_sg U49016 ( .A(n20505), .X(n45924) );
  nor_x1_sg U49017 ( .A(n21082), .B(n21083), .X(n6691) );
  nand_x1_sg U49018 ( .A(n45866), .B(n6714), .X(n6713) );
  nand_x1_sg U49019 ( .A(n45871), .B(n21599), .X(n21597) );
  nor_x1_sg U49020 ( .A(n19627), .B(n45856), .X(n6763) );
  inv_x1_sg U49021 ( .A(n19628), .X(n45856) );
  nor_x1_sg U49022 ( .A(n19394), .B(n45860), .X(n6764) );
  inv_x1_sg U49023 ( .A(n19395), .X(n45860) );
  nor_x1_sg U49024 ( .A(n19217), .B(n45864), .X(n6753) );
  inv_x1_sg U49025 ( .A(n19218), .X(n45864) );
  nor_x1_sg U49026 ( .A(n19833), .B(n45852), .X(n6744) );
  inv_x1_sg U49027 ( .A(n19834), .X(n45852) );
  nor_x1_sg U49028 ( .A(n20021), .B(n45848), .X(n6743) );
  inv_x1_sg U49029 ( .A(n20022), .X(n45848) );
  nor_x1_sg U49030 ( .A(n20360), .B(n45840), .X(n6747) );
  inv_x1_sg U49031 ( .A(n20361), .X(n45840) );
  inv_x1_sg U49032 ( .A(n21591), .X(n45813) );
  nor_x1_sg U49033 ( .A(n21259), .B(n45820), .X(n6772) );
  inv_x1_sg U49034 ( .A(n21260), .X(n45820) );
  nor_x1_sg U49035 ( .A(n20490), .B(n45836), .X(n6778) );
  inv_x1_sg U49036 ( .A(n20491), .X(n45836) );
  nor_x1_sg U49037 ( .A(n20661), .B(n45832), .X(n6777) );
  inv_x1_sg U49038 ( .A(n20662), .X(n45832) );
  nor_x1_sg U49039 ( .A(n21069), .B(n45824), .X(n6781) );
  inv_x1_sg U49040 ( .A(n21070), .X(n45824) );
  nor_x1_sg U49041 ( .A(n19392), .B(n19393), .X(n19216) );
  nor_x1_sg U49042 ( .A(n19624), .B(n19625), .X(n6807) );
  nor_x1_sg U49043 ( .A(n20198), .B(n20199), .X(n20020) );
  nor_x1_sg U49044 ( .A(n20018), .B(n20019), .X(n6794) );
  nor_x1_sg U49045 ( .A(n20357), .B(n20358), .X(n6797) );
  nor_x1_sg U49046 ( .A(n20841), .B(n20842), .X(n20660) );
  nor_x1_sg U49047 ( .A(n20658), .B(n20659), .X(n6818) );
  nor_x1_sg U49048 ( .A(n21066), .B(n21067), .X(n6821) );
  nand_x1_sg U49049 ( .A(n22849), .B(n22850), .X(n22848) );
  nand_x1_sg U49050 ( .A(n46859), .B(n7073), .X(n7072) );
  nor_x1_sg U49051 ( .A(n7084), .B(n7085), .X(n7082) );
  nor_x1_sg U49052 ( .A(n7099), .B(n7100), .X(n7095) );
  inv_x1_sg U49053 ( .A(n7116), .X(n46886) );
  nor_x1_sg U49054 ( .A(n7163), .B(n7164), .X(n7160) );
  nand_x1_sg U49055 ( .A(n7123), .B(n7124), .X(n7116) );
  nand_x1_sg U49056 ( .A(n46864), .B(n7107), .X(n7123) );
  nor_x1_sg U49057 ( .A(n7134), .B(n46894), .X(n7114) );
  nand_x1_sg U49058 ( .A(n7139), .B(n7150), .X(n7144) );
  nand_x1_sg U49059 ( .A(n46908), .B(n7159), .X(n7145) );
  nand_x2_sg U49060 ( .A(n7202), .B(n7203), .X(n7196) );
  nand_x1_sg U49061 ( .A(n7218), .B(n46948), .X(n7197) );
  nor_x1_sg U49062 ( .A(n47013), .B(n7319), .X(n7312) );
  nor_x1_sg U49063 ( .A(n47044), .B(n7411), .X(n7404) );
  nand_x1_sg U49064 ( .A(n7459), .B(n7414), .X(n7452) );
  nor_x1_sg U49065 ( .A(n7037), .B(n7038), .X(n6975) );
  nand_x1_sg U49066 ( .A(n6976), .B(n47123), .X(n6974) );
  nand_x1_sg U49067 ( .A(n6947), .B(n6948), .X(n6940) );
  nand_x2_sg U49068 ( .A(n6941), .B(n6942), .X(n6939) );
  nand_x1_sg U49069 ( .A(n6959), .B(n6960), .X(n6952) );
  nand_x1_sg U49070 ( .A(n46961), .B(n6961), .X(n6960) );
  nand_x1_sg U49071 ( .A(n6955), .B(n6956), .X(n6954) );
  nand_x1_sg U49072 ( .A(n47152), .B(n7891), .X(n7890) );
  nor_x1_sg U49073 ( .A(n7902), .B(n7903), .X(n7900) );
  nand_x4_sg U49074 ( .A(n7945), .B(n47174), .X(n7925) );
  nor_x1_sg U49075 ( .A(n7917), .B(n7918), .X(n7913) );
  inv_x1_sg U49076 ( .A(n7934), .X(n47179) );
  nor_x1_sg U49077 ( .A(n7982), .B(n7983), .X(n7979) );
  nand_x1_sg U49078 ( .A(n7941), .B(n7942), .X(n7934) );
  nand_x1_sg U49079 ( .A(n47157), .B(n7925), .X(n7941) );
  nor_x1_sg U49080 ( .A(n7952), .B(n47189), .X(n7932) );
  nand_x1_sg U49081 ( .A(n7957), .B(n7968), .X(n7962) );
  nand_x1_sg U49082 ( .A(n47201), .B(n7978), .X(n7963) );
  nand_x2_sg U49083 ( .A(n8021), .B(n8022), .X(n8015) );
  nand_x1_sg U49084 ( .A(n8037), .B(n47239), .X(n8016) );
  nor_x1_sg U49085 ( .A(n47301), .B(n8137), .X(n8130) );
  nor_x1_sg U49086 ( .A(n47331), .B(n8229), .X(n8222) );
  nand_x1_sg U49087 ( .A(n8277), .B(n8232), .X(n8270) );
  nor_x1_sg U49088 ( .A(n7855), .B(n7856), .X(n7792) );
  nand_x1_sg U49089 ( .A(n7793), .B(n47409), .X(n7791) );
  nand_x1_sg U49090 ( .A(n7764), .B(n7765), .X(n7757) );
  nand_x2_sg U49091 ( .A(n7758), .B(n7759), .X(n7756) );
  nand_x1_sg U49092 ( .A(n7776), .B(n7777), .X(n7769) );
  nand_x1_sg U49093 ( .A(n47252), .B(n7778), .X(n7777) );
  nand_x1_sg U49094 ( .A(n7772), .B(n7773), .X(n7771) );
  nand_x1_sg U49095 ( .A(n47437), .B(n8709), .X(n8708) );
  nor_x1_sg U49096 ( .A(n8720), .B(n8721), .X(n8718) );
  nand_x4_sg U49097 ( .A(n8763), .B(n47459), .X(n8743) );
  nor_x1_sg U49098 ( .A(n8735), .B(n8736), .X(n8731) );
  inv_x1_sg U49099 ( .A(n8752), .X(n47464) );
  nor_x1_sg U49100 ( .A(n8800), .B(n8801), .X(n8797) );
  nand_x1_sg U49101 ( .A(n8759), .B(n8760), .X(n8752) );
  nand_x1_sg U49102 ( .A(n47442), .B(n8743), .X(n8759) );
  nor_x1_sg U49103 ( .A(n8770), .B(n47474), .X(n8750) );
  nand_x1_sg U49104 ( .A(n8775), .B(n8786), .X(n8780) );
  nand_x1_sg U49105 ( .A(n47486), .B(n8796), .X(n8781) );
  nand_x2_sg U49106 ( .A(n8839), .B(n8840), .X(n8833) );
  nand_x1_sg U49107 ( .A(n8855), .B(n47524), .X(n8834) );
  nor_x1_sg U49108 ( .A(n47586), .B(n8955), .X(n8948) );
  nor_x1_sg U49109 ( .A(n47616), .B(n9047), .X(n9040) );
  nand_x1_sg U49110 ( .A(n9095), .B(n9050), .X(n9088) );
  nor_x1_sg U49111 ( .A(n8673), .B(n8674), .X(n8610) );
  nand_x1_sg U49112 ( .A(n8611), .B(n47694), .X(n8609) );
  nand_x1_sg U49113 ( .A(n8582), .B(n8583), .X(n8575) );
  nand_x2_sg U49114 ( .A(n8576), .B(n8577), .X(n8574) );
  nand_x1_sg U49115 ( .A(n8594), .B(n8595), .X(n8587) );
  nand_x1_sg U49116 ( .A(n47537), .B(n8596), .X(n8595) );
  nand_x1_sg U49117 ( .A(n8590), .B(n8591), .X(n8589) );
  nand_x1_sg U49118 ( .A(n47722), .B(n9529), .X(n9528) );
  nor_x1_sg U49119 ( .A(n9540), .B(n9541), .X(n9538) );
  nand_x4_sg U49120 ( .A(n9583), .B(n47744), .X(n9563) );
  nor_x1_sg U49121 ( .A(n9555), .B(n9556), .X(n9551) );
  inv_x1_sg U49122 ( .A(n9572), .X(n47749) );
  nor_x1_sg U49123 ( .A(n9620), .B(n9621), .X(n9617) );
  nand_x1_sg U49124 ( .A(n9579), .B(n9580), .X(n9572) );
  nand_x1_sg U49125 ( .A(n47727), .B(n9563), .X(n9579) );
  nor_x1_sg U49126 ( .A(n9590), .B(n47759), .X(n9570) );
  nand_x1_sg U49127 ( .A(n9595), .B(n9606), .X(n9600) );
  nand_x1_sg U49128 ( .A(n47771), .B(n9616), .X(n9601) );
  nand_x2_sg U49129 ( .A(n9659), .B(n9660), .X(n9653) );
  nand_x1_sg U49130 ( .A(n9675), .B(n47809), .X(n9654) );
  nor_x1_sg U49131 ( .A(n47871), .B(n9775), .X(n9768) );
  nor_x1_sg U49132 ( .A(n47901), .B(n9867), .X(n9860) );
  nand_x1_sg U49133 ( .A(n9915), .B(n9870), .X(n9908) );
  nor_x1_sg U49134 ( .A(n9493), .B(n9494), .X(n9430) );
  nand_x1_sg U49135 ( .A(n9431), .B(n47979), .X(n9429) );
  nand_x1_sg U49136 ( .A(n9402), .B(n9403), .X(n9395) );
  nand_x2_sg U49137 ( .A(n9396), .B(n9397), .X(n9394) );
  nand_x1_sg U49138 ( .A(n9414), .B(n9415), .X(n9407) );
  nand_x1_sg U49139 ( .A(n47822), .B(n9416), .X(n9415) );
  nand_x1_sg U49140 ( .A(n9410), .B(n9411), .X(n9409) );
  nand_x1_sg U49141 ( .A(n48007), .B(n10348), .X(n10347) );
  nor_x1_sg U49142 ( .A(n10359), .B(n10360), .X(n10357) );
  nand_x4_sg U49143 ( .A(n10402), .B(n48029), .X(n10382) );
  nor_x1_sg U49144 ( .A(n10374), .B(n10375), .X(n10370) );
  inv_x1_sg U49145 ( .A(n10391), .X(n48034) );
  nor_x1_sg U49146 ( .A(n10439), .B(n10440), .X(n10436) );
  nand_x1_sg U49147 ( .A(n10398), .B(n10399), .X(n10391) );
  nand_x1_sg U49148 ( .A(n48012), .B(n10382), .X(n10398) );
  nor_x1_sg U49149 ( .A(n10409), .B(n48044), .X(n10389) );
  nand_x1_sg U49150 ( .A(n10414), .B(n10425), .X(n10419) );
  nand_x1_sg U49151 ( .A(n48056), .B(n10435), .X(n10420) );
  nand_x2_sg U49152 ( .A(n10478), .B(n10479), .X(n10472) );
  nand_x1_sg U49153 ( .A(n10494), .B(n48094), .X(n10473) );
  nor_x1_sg U49154 ( .A(n48156), .B(n10594), .X(n10587) );
  nor_x1_sg U49155 ( .A(n48186), .B(n10686), .X(n10679) );
  nand_x1_sg U49156 ( .A(n10734), .B(n10689), .X(n10727) );
  nor_x1_sg U49157 ( .A(n10312), .B(n10313), .X(n10249) );
  nand_x1_sg U49158 ( .A(n10250), .B(n48264), .X(n10248) );
  nand_x1_sg U49159 ( .A(n10221), .B(n10222), .X(n10214) );
  nand_x2_sg U49160 ( .A(n10215), .B(n10216), .X(n10213) );
  nand_x1_sg U49161 ( .A(n10233), .B(n10234), .X(n10226) );
  nand_x1_sg U49162 ( .A(n48107), .B(n10235), .X(n10234) );
  nand_x1_sg U49163 ( .A(n10229), .B(n10230), .X(n10228) );
  nand_x1_sg U49164 ( .A(n48292), .B(n11167), .X(n11166) );
  nor_x1_sg U49165 ( .A(n11178), .B(n11179), .X(n11176) );
  nand_x4_sg U49166 ( .A(n11221), .B(n48314), .X(n11201) );
  nor_x1_sg U49167 ( .A(n11193), .B(n11194), .X(n11189) );
  inv_x1_sg U49168 ( .A(n11210), .X(n48319) );
  nor_x1_sg U49169 ( .A(n11258), .B(n11259), .X(n11255) );
  nand_x1_sg U49170 ( .A(n11217), .B(n11218), .X(n11210) );
  nand_x1_sg U49171 ( .A(n48297), .B(n11201), .X(n11217) );
  nor_x1_sg U49172 ( .A(n11228), .B(n48329), .X(n11208) );
  nand_x1_sg U49173 ( .A(n11233), .B(n11244), .X(n11238) );
  nand_x1_sg U49174 ( .A(n48341), .B(n11254), .X(n11239) );
  nand_x2_sg U49175 ( .A(n11297), .B(n11298), .X(n11291) );
  nand_x1_sg U49176 ( .A(n11313), .B(n48379), .X(n11292) );
  nor_x1_sg U49177 ( .A(n48441), .B(n11413), .X(n11406) );
  nor_x1_sg U49178 ( .A(n48471), .B(n11505), .X(n11498) );
  nand_x1_sg U49179 ( .A(n11553), .B(n11508), .X(n11546) );
  nor_x1_sg U49180 ( .A(n11131), .B(n11132), .X(n11068) );
  nand_x1_sg U49181 ( .A(n11069), .B(n48549), .X(n11067) );
  nand_x1_sg U49182 ( .A(n11040), .B(n11041), .X(n11033) );
  nand_x2_sg U49183 ( .A(n11034), .B(n11035), .X(n11032) );
  nand_x1_sg U49184 ( .A(n11052), .B(n11053), .X(n11045) );
  nand_x1_sg U49185 ( .A(n48392), .B(n11054), .X(n11053) );
  nand_x1_sg U49186 ( .A(n11048), .B(n11049), .X(n11047) );
  nand_x1_sg U49187 ( .A(n48577), .B(n11986), .X(n11985) );
  nor_x1_sg U49188 ( .A(n11997), .B(n11998), .X(n11995) );
  nand_x4_sg U49189 ( .A(n12040), .B(n48599), .X(n12020) );
  nor_x1_sg U49190 ( .A(n12012), .B(n12013), .X(n12008) );
  inv_x1_sg U49191 ( .A(n12029), .X(n48604) );
  nor_x1_sg U49192 ( .A(n12077), .B(n12078), .X(n12074) );
  nand_x1_sg U49193 ( .A(n12036), .B(n12037), .X(n12029) );
  nand_x1_sg U49194 ( .A(n48582), .B(n12020), .X(n12036) );
  nor_x1_sg U49195 ( .A(n12047), .B(n48614), .X(n12027) );
  nand_x1_sg U49196 ( .A(n12052), .B(n12063), .X(n12057) );
  nand_x1_sg U49197 ( .A(n48626), .B(n12073), .X(n12058) );
  nand_x2_sg U49198 ( .A(n12116), .B(n12117), .X(n12110) );
  nand_x1_sg U49199 ( .A(n12132), .B(n48664), .X(n12111) );
  nor_x1_sg U49200 ( .A(n48726), .B(n12232), .X(n12225) );
  nor_x1_sg U49201 ( .A(n48756), .B(n12324), .X(n12317) );
  nand_x1_sg U49202 ( .A(n12372), .B(n12327), .X(n12365) );
  nor_x1_sg U49203 ( .A(n11950), .B(n11951), .X(n11887) );
  nand_x1_sg U49204 ( .A(n11888), .B(n48834), .X(n11886) );
  nand_x1_sg U49205 ( .A(n11859), .B(n11860), .X(n11852) );
  nand_x2_sg U49206 ( .A(n11853), .B(n11854), .X(n11851) );
  nand_x1_sg U49207 ( .A(n11871), .B(n11872), .X(n11864) );
  nand_x1_sg U49208 ( .A(n48677), .B(n11873), .X(n11872) );
  nand_x1_sg U49209 ( .A(n11867), .B(n11868), .X(n11866) );
  nand_x1_sg U49210 ( .A(n48863), .B(n12805), .X(n12804) );
  nor_x1_sg U49211 ( .A(n12816), .B(n12817), .X(n12814) );
  nand_x4_sg U49212 ( .A(n12859), .B(n48885), .X(n12839) );
  nor_x1_sg U49213 ( .A(n12831), .B(n12832), .X(n12827) );
  inv_x1_sg U49214 ( .A(n12848), .X(n48890) );
  nor_x1_sg U49215 ( .A(n12896), .B(n12897), .X(n12893) );
  nand_x1_sg U49216 ( .A(n12855), .B(n12856), .X(n12848) );
  nand_x1_sg U49217 ( .A(n48868), .B(n12839), .X(n12855) );
  nor_x1_sg U49218 ( .A(n12866), .B(n48900), .X(n12846) );
  nand_x1_sg U49219 ( .A(n12871), .B(n12882), .X(n12876) );
  nand_x1_sg U49220 ( .A(n48912), .B(n12892), .X(n12877) );
  nand_x2_sg U49221 ( .A(n12935), .B(n12936), .X(n12929) );
  nand_x1_sg U49222 ( .A(n12951), .B(n48950), .X(n12930) );
  nor_x1_sg U49223 ( .A(n49012), .B(n13051), .X(n13044) );
  nor_x1_sg U49224 ( .A(n49042), .B(n13143), .X(n13136) );
  nand_x1_sg U49225 ( .A(n13191), .B(n13146), .X(n13184) );
  nor_x1_sg U49226 ( .A(n12769), .B(n12770), .X(n12706) );
  nand_x1_sg U49227 ( .A(n12707), .B(n49121), .X(n12705) );
  nand_x1_sg U49228 ( .A(n12678), .B(n12679), .X(n12671) );
  nand_x2_sg U49229 ( .A(n12672), .B(n12673), .X(n12670) );
  nand_x1_sg U49230 ( .A(n12690), .B(n12691), .X(n12683) );
  nand_x1_sg U49231 ( .A(n48963), .B(n12692), .X(n12691) );
  nand_x1_sg U49232 ( .A(n12686), .B(n12687), .X(n12685) );
  nand_x1_sg U49233 ( .A(n49150), .B(n13624), .X(n13623) );
  nor_x1_sg U49234 ( .A(n13635), .B(n13636), .X(n13633) );
  nand_x4_sg U49235 ( .A(n13678), .B(n49172), .X(n13658) );
  nor_x1_sg U49236 ( .A(n13650), .B(n13651), .X(n13646) );
  inv_x1_sg U49237 ( .A(n13667), .X(n49177) );
  nor_x1_sg U49238 ( .A(n13715), .B(n13716), .X(n13712) );
  nand_x1_sg U49239 ( .A(n13674), .B(n13675), .X(n13667) );
  nand_x1_sg U49240 ( .A(n49155), .B(n13658), .X(n13674) );
  nor_x1_sg U49241 ( .A(n13685), .B(n49187), .X(n13665) );
  nand_x1_sg U49242 ( .A(n13690), .B(n13701), .X(n13695) );
  nand_x1_sg U49243 ( .A(n49199), .B(n13711), .X(n13696) );
  nand_x2_sg U49244 ( .A(n13754), .B(n13755), .X(n13748) );
  nand_x1_sg U49245 ( .A(n13770), .B(n49237), .X(n13749) );
  nor_x1_sg U49246 ( .A(n49299), .B(n13870), .X(n13863) );
  nor_x1_sg U49247 ( .A(n49329), .B(n13962), .X(n13955) );
  nand_x1_sg U49248 ( .A(n14010), .B(n13965), .X(n14003) );
  nor_x1_sg U49249 ( .A(n13588), .B(n13589), .X(n13525) );
  nand_x1_sg U49250 ( .A(n13526), .B(n49407), .X(n13524) );
  nand_x1_sg U49251 ( .A(n13497), .B(n13498), .X(n13490) );
  nand_x2_sg U49252 ( .A(n13491), .B(n13492), .X(n13489) );
  nand_x1_sg U49253 ( .A(n13509), .B(n13510), .X(n13502) );
  nand_x1_sg U49254 ( .A(n49250), .B(n13511), .X(n13510) );
  nand_x1_sg U49255 ( .A(n13505), .B(n13506), .X(n13504) );
  nand_x1_sg U49256 ( .A(n49436), .B(n14443), .X(n14442) );
  nor_x1_sg U49257 ( .A(n14454), .B(n14455), .X(n14452) );
  nor_x1_sg U49258 ( .A(n14469), .B(n14470), .X(n14465) );
  inv_x1_sg U49259 ( .A(n14486), .X(n49463) );
  nor_x1_sg U49260 ( .A(n14534), .B(n14535), .X(n14531) );
  nand_x1_sg U49261 ( .A(n14493), .B(n14494), .X(n14486) );
  nand_x1_sg U49262 ( .A(n49441), .B(n14477), .X(n14493) );
  nor_x1_sg U49263 ( .A(n14504), .B(n49473), .X(n14484) );
  nand_x1_sg U49264 ( .A(n14509), .B(n14520), .X(n14514) );
  nand_x1_sg U49265 ( .A(n49485), .B(n14530), .X(n14515) );
  nand_x2_sg U49266 ( .A(n14573), .B(n14574), .X(n14567) );
  nand_x1_sg U49267 ( .A(n14589), .B(n49523), .X(n14568) );
  nor_x1_sg U49268 ( .A(n49585), .B(n14689), .X(n14682) );
  nor_x1_sg U49269 ( .A(n49615), .B(n14781), .X(n14774) );
  nand_x1_sg U49270 ( .A(n14829), .B(n14784), .X(n14822) );
  nor_x1_sg U49271 ( .A(n14407), .B(n14408), .X(n14344) );
  nand_x1_sg U49272 ( .A(n14345), .B(n49693), .X(n14343) );
  nand_x1_sg U49273 ( .A(n14316), .B(n14317), .X(n14309) );
  nand_x2_sg U49274 ( .A(n14310), .B(n14311), .X(n14308) );
  nand_x1_sg U49275 ( .A(n14328), .B(n14329), .X(n14321) );
  nand_x1_sg U49276 ( .A(n49536), .B(n14330), .X(n14329) );
  nand_x1_sg U49277 ( .A(n14324), .B(n14325), .X(n14323) );
  nand_x1_sg U49278 ( .A(n49721), .B(n15262), .X(n15261) );
  nor_x1_sg U49279 ( .A(n15273), .B(n15274), .X(n15271) );
  nor_x1_sg U49280 ( .A(n15288), .B(n15289), .X(n15284) );
  inv_x1_sg U49281 ( .A(n15305), .X(n49748) );
  nor_x1_sg U49282 ( .A(n15353), .B(n15354), .X(n15350) );
  nand_x1_sg U49283 ( .A(n15312), .B(n15313), .X(n15305) );
  nand_x1_sg U49284 ( .A(n49726), .B(n15296), .X(n15312) );
  nor_x1_sg U49285 ( .A(n15323), .B(n49759), .X(n15303) );
  nand_x1_sg U49286 ( .A(n15328), .B(n15339), .X(n15333) );
  nand_x1_sg U49287 ( .A(n49771), .B(n15349), .X(n15334) );
  nand_x2_sg U49288 ( .A(n15392), .B(n15393), .X(n15386) );
  nand_x1_sg U49289 ( .A(n15408), .B(n49809), .X(n15387) );
  nor_x1_sg U49290 ( .A(n49871), .B(n15508), .X(n15501) );
  nor_x1_sg U49291 ( .A(n49901), .B(n15600), .X(n15593) );
  nand_x1_sg U49292 ( .A(n15648), .B(n15603), .X(n15641) );
  nor_x1_sg U49293 ( .A(n15226), .B(n15227), .X(n15163) );
  nand_x1_sg U49294 ( .A(n15164), .B(n49979), .X(n15162) );
  nand_x1_sg U49295 ( .A(n15135), .B(n15136), .X(n15128) );
  nand_x2_sg U49296 ( .A(n15129), .B(n15130), .X(n15127) );
  nand_x1_sg U49297 ( .A(n15147), .B(n15148), .X(n15140) );
  nand_x1_sg U49298 ( .A(n49822), .B(n15149), .X(n15148) );
  nand_x1_sg U49299 ( .A(n15143), .B(n15144), .X(n15142) );
  nand_x1_sg U49300 ( .A(n50008), .B(n16081), .X(n16080) );
  nor_x1_sg U49301 ( .A(n16092), .B(n16093), .X(n16090) );
  nor_x1_sg U49302 ( .A(n16107), .B(n16108), .X(n16103) );
  inv_x1_sg U49303 ( .A(n16124), .X(n50035) );
  nor_x1_sg U49304 ( .A(n16172), .B(n16173), .X(n16169) );
  nand_x1_sg U49305 ( .A(n16131), .B(n16132), .X(n16124) );
  nand_x1_sg U49306 ( .A(n50013), .B(n16115), .X(n16131) );
  nor_x1_sg U49307 ( .A(n16142), .B(n50045), .X(n16122) );
  nand_x1_sg U49308 ( .A(n16147), .B(n16158), .X(n16152) );
  nand_x1_sg U49309 ( .A(n50057), .B(n16168), .X(n16153) );
  nand_x2_sg U49310 ( .A(n16211), .B(n16212), .X(n16205) );
  nand_x1_sg U49311 ( .A(n16227), .B(n50095), .X(n16206) );
  nor_x1_sg U49312 ( .A(n50157), .B(n16327), .X(n16320) );
  nor_x1_sg U49313 ( .A(n50187), .B(n16419), .X(n16412) );
  nand_x1_sg U49314 ( .A(n16467), .B(n16422), .X(n16460) );
  nor_x1_sg U49315 ( .A(n16045), .B(n16046), .X(n15982) );
  nand_x1_sg U49316 ( .A(n15983), .B(n50265), .X(n15981) );
  nand_x1_sg U49317 ( .A(n15954), .B(n15955), .X(n15947) );
  nand_x2_sg U49318 ( .A(n15948), .B(n15949), .X(n15946) );
  nand_x1_sg U49319 ( .A(n15966), .B(n15967), .X(n15959) );
  nand_x1_sg U49320 ( .A(n50108), .B(n15968), .X(n15967) );
  nand_x1_sg U49321 ( .A(n15962), .B(n15963), .X(n15961) );
  nand_x1_sg U49322 ( .A(n50292), .B(n16900), .X(n16899) );
  nor_x1_sg U49323 ( .A(n16910), .B(n16911), .X(n16909) );
  nor_x1_sg U49324 ( .A(n16924), .B(n16925), .X(n16920) );
  inv_x1_sg U49325 ( .A(n16941), .X(n50320) );
  nor_x1_sg U49326 ( .A(n16988), .B(n16989), .X(n16985) );
  nand_x1_sg U49327 ( .A(n16948), .B(n16949), .X(n16941) );
  nand_x1_sg U49328 ( .A(n50297), .B(n16932), .X(n16948) );
  nor_x1_sg U49329 ( .A(n16959), .B(n50327), .X(n16939) );
  nand_x1_sg U49330 ( .A(n16964), .B(n16975), .X(n16969) );
  nand_x1_sg U49331 ( .A(n50342), .B(n16984), .X(n16970) );
  nand_x2_sg U49332 ( .A(n17027), .B(n17028), .X(n17021) );
  nand_x1_sg U49333 ( .A(n17043), .B(n50380), .X(n17022) );
  nor_x1_sg U49334 ( .A(n50442), .B(n17144), .X(n17137) );
  nor_x1_sg U49335 ( .A(n50472), .B(n17236), .X(n17229) );
  nand_x1_sg U49336 ( .A(n17284), .B(n17239), .X(n17277) );
  nor_x1_sg U49337 ( .A(n16864), .B(n16865), .X(n16799) );
  nand_x1_sg U49338 ( .A(n16800), .B(n50551), .X(n16798) );
  nand_x1_sg U49339 ( .A(n16771), .B(n16772), .X(n16764) );
  nand_x2_sg U49340 ( .A(n16765), .B(n16766), .X(n16763) );
  nand_x1_sg U49341 ( .A(n16783), .B(n16784), .X(n16776) );
  nand_x1_sg U49342 ( .A(n50393), .B(n16785), .X(n16784) );
  nand_x1_sg U49343 ( .A(n16779), .B(n16780), .X(n16778) );
  nand_x1_sg U49344 ( .A(n50582), .B(n17719), .X(n17718) );
  nor_x1_sg U49345 ( .A(n17730), .B(n17731), .X(n17728) );
  nor_x1_sg U49346 ( .A(n17745), .B(n17746), .X(n17741) );
  inv_x1_sg U49347 ( .A(n17762), .X(n50609) );
  nor_x1_sg U49348 ( .A(n17810), .B(n17811), .X(n17807) );
  nand_x1_sg U49349 ( .A(n17769), .B(n17770), .X(n17762) );
  nand_x1_sg U49350 ( .A(n50587), .B(n17753), .X(n17769) );
  nor_x1_sg U49351 ( .A(n17780), .B(n50619), .X(n17760) );
  nand_x1_sg U49352 ( .A(n17785), .B(n17796), .X(n17790) );
  nand_x1_sg U49353 ( .A(n50631), .B(n17806), .X(n17791) );
  nand_x2_sg U49354 ( .A(n17849), .B(n17850), .X(n17843) );
  nand_x1_sg U49355 ( .A(n17865), .B(n50669), .X(n17844) );
  nor_x1_sg U49356 ( .A(n50731), .B(n17965), .X(n17958) );
  nor_x1_sg U49357 ( .A(n50761), .B(n18057), .X(n18050) );
  nand_x1_sg U49358 ( .A(n18105), .B(n18060), .X(n18098) );
  nor_x1_sg U49359 ( .A(n17683), .B(n17684), .X(n17620) );
  nand_x1_sg U49360 ( .A(n17621), .B(n50839), .X(n17619) );
  nand_x1_sg U49361 ( .A(n17592), .B(n17593), .X(n17585) );
  nand_x2_sg U49362 ( .A(n17586), .B(n17587), .X(n17584) );
  nand_x1_sg U49363 ( .A(n17604), .B(n17605), .X(n17597) );
  nand_x1_sg U49364 ( .A(n50682), .B(n17606), .X(n17605) );
  nand_x1_sg U49365 ( .A(n17600), .B(n17601), .X(n17599) );
  nand_x1_sg U49366 ( .A(n50869), .B(n18540), .X(n18539) );
  nor_x1_sg U49367 ( .A(n18551), .B(n18552), .X(n18549) );
  nor_x1_sg U49368 ( .A(n18566), .B(n18567), .X(n18562) );
  inv_x1_sg U49369 ( .A(n18583), .X(n50896) );
  nor_x1_sg U49370 ( .A(n18631), .B(n18632), .X(n18628) );
  nand_x1_sg U49371 ( .A(n18590), .B(n18591), .X(n18583) );
  nand_x1_sg U49372 ( .A(n50874), .B(n18574), .X(n18590) );
  nor_x1_sg U49373 ( .A(n18601), .B(n50906), .X(n18581) );
  nand_x1_sg U49374 ( .A(n18606), .B(n18617), .X(n18611) );
  nand_x1_sg U49375 ( .A(n50918), .B(n18627), .X(n18612) );
  nand_x2_sg U49376 ( .A(n18670), .B(n18671), .X(n18664) );
  nand_x1_sg U49377 ( .A(n18686), .B(n50956), .X(n18665) );
  nor_x1_sg U49378 ( .A(n51018), .B(n18786), .X(n18779) );
  nor_x1_sg U49379 ( .A(n51048), .B(n18878), .X(n18871) );
  nand_x1_sg U49380 ( .A(n18926), .B(n18881), .X(n18919) );
  nor_x1_sg U49381 ( .A(n18504), .B(n18505), .X(n18441) );
  nand_x1_sg U49382 ( .A(n18442), .B(n51126), .X(n18440) );
  nand_x1_sg U49383 ( .A(n18413), .B(n18414), .X(n18406) );
  nand_x2_sg U49384 ( .A(n18407), .B(n18408), .X(n18405) );
  nand_x1_sg U49385 ( .A(n18425), .B(n18426), .X(n18418) );
  nand_x1_sg U49386 ( .A(n50969), .B(n18427), .X(n18426) );
  nand_x1_sg U49387 ( .A(n18421), .B(n18422), .X(n18420) );
  nand_x1_sg U49388 ( .A(n28553), .B(n28554), .X(n28552) );
  nand_x1_sg U49389 ( .A(n26833), .B(n26834), .X(n26832) );
  nand_x1_sg U49390 ( .A(n26897), .B(n26898), .X(n26896) );
  nand_x1_sg U49391 ( .A(n26890), .B(n26891), .X(n26889) );
  inv_x1_sg U49392 ( .A(n26881), .X(n45771) );
  nand_x1_sg U49393 ( .A(n28560), .B(n28561), .X(n28559) );
  nor_x1_sg U49394 ( .A(n26823), .B(n45789), .X(n26781) );
  inv_x1_sg U49395 ( .A(n26824), .X(n45789) );
  nand_x1_sg U49396 ( .A(n28546), .B(n28547), .X(n28545) );
  nand_x1_sg U49397 ( .A(n28567), .B(n28568), .X(n28566) );
  nor_x1_sg U49398 ( .A(n29268), .B(n29269), .X(n29226) );
  nor_x1_sg U49399 ( .A(n29216), .B(n29217), .X(n29215) );
  nor_x1_sg U49400 ( .A(n29204), .B(n29205), .X(n29203) );
  nor_x1_sg U49401 ( .A(n45398), .B(n28310), .X(n22116) );
  inv_x1_sg U49402 ( .A(n28312), .X(n45398) );
  nor_x1_sg U49403 ( .A(n45352), .B(n28304), .X(n22164) );
  inv_x1_sg U49404 ( .A(n28306), .X(n45352) );
  nor_x1_sg U49405 ( .A(n29192), .B(n29193), .X(n29191) );
  nor_x1_sg U49406 ( .A(n45307), .B(n28298), .X(n22211) );
  inv_x1_sg U49407 ( .A(n28300), .X(n45307) );
  nor_x1_sg U49408 ( .A(n45262), .B(n28292), .X(n22259) );
  inv_x1_sg U49409 ( .A(n28294), .X(n45262) );
  nor_x1_sg U49410 ( .A(n29180), .B(n29181), .X(n29179) );
  nor_x1_sg U49411 ( .A(n45217), .B(n28286), .X(n22306) );
  inv_x1_sg U49412 ( .A(n28288), .X(n45217) );
  nor_x1_sg U49413 ( .A(n45171), .B(n28280), .X(n22354) );
  inv_x1_sg U49414 ( .A(n28282), .X(n45171) );
  nor_x1_sg U49415 ( .A(n29168), .B(n29169), .X(n29167) );
  nor_x1_sg U49416 ( .A(n45126), .B(n28274), .X(n22401) );
  inv_x1_sg U49417 ( .A(n28276), .X(n45126) );
  nor_x1_sg U49418 ( .A(n29156), .B(n29157), .X(n29155) );
  nand_x1_sg U49419 ( .A(n28458), .B(n28459), .X(n28380) );
  nand_x1_sg U49420 ( .A(n28976), .B(n28977), .X(n28823) );
  nand_x1_sg U49421 ( .A(n27187), .B(n27188), .X(n26964) );
  nand_x1_sg U49422 ( .A(n22550), .B(n26948), .X(n22513) );
  nand_x1_sg U49423 ( .A(n26949), .B(n22589), .X(n26948) );
  nand_x1_sg U49424 ( .A(n28806), .B(n28807), .X(n28635) );
  nand_x1_sg U49425 ( .A(n28618), .B(n28619), .X(n28474) );
  nand_x1_sg U49426 ( .A(n29136), .B(n29137), .X(n28994) );
  inv_x1_sg U49427 ( .A(n27193), .X(n45014) );
  nor_x1_sg U49428 ( .A(n28256), .B(n44995), .X(n22535) );
  inv_x1_sg U49429 ( .A(n28257), .X(n44995) );
  nor_x1_sg U49430 ( .A(n22804), .B(n22805), .X(n22800) );
  nor_x1_sg U49431 ( .A(n22808), .B(n22809), .X(n22803) );
  nor_x1_sg U49432 ( .A(n22797), .B(n22798), .X(n22792) );
  inv_x1_sg U49433 ( .A(n22781), .X(n46903) );
  nand_x1_sg U49434 ( .A(n22783), .B(n22784), .X(n22781) );
  nand_x1_sg U49435 ( .A(n22769), .B(n22770), .X(n22767) );
  nand_x1_sg U49436 ( .A(n22762), .B(n22763), .X(n22760) );
  inv_x1_sg U49437 ( .A(n22753), .X(n46984) );
  nand_x1_sg U49438 ( .A(n22755), .B(n22756), .X(n22753) );
  inv_x1_sg U49439 ( .A(n22746), .X(n47007) );
  nand_x1_sg U49440 ( .A(n22748), .B(n22749), .X(n22746) );
  nand_x1_sg U49441 ( .A(n22741), .B(n22742), .X(n22739) );
  inv_x1_sg U49442 ( .A(n22718), .X(n47120) );
  inv_x1_sg U49443 ( .A(n23104), .X(n47150) );
  nor_x1_sg U49444 ( .A(n23081), .B(n23082), .X(n23077) );
  nor_x1_sg U49445 ( .A(n23085), .B(n23086), .X(n23080) );
  nor_x1_sg U49446 ( .A(n23074), .B(n23075), .X(n23069) );
  inv_x1_sg U49447 ( .A(n23058), .X(n47196) );
  nand_x1_sg U49448 ( .A(n23060), .B(n23061), .X(n23058) );
  inv_x1_sg U49449 ( .A(n23044), .X(n47233) );
  nand_x1_sg U49450 ( .A(n23046), .B(n23047), .X(n23044) );
  inv_x1_sg U49451 ( .A(n23030), .X(n47273) );
  nand_x1_sg U49452 ( .A(n23032), .B(n23033), .X(n23030) );
  nand_x1_sg U49453 ( .A(n23018), .B(n23019), .X(n23016) );
  inv_x1_sg U49454 ( .A(n23384), .X(n47435) );
  nor_x1_sg U49455 ( .A(n23361), .B(n23362), .X(n23357) );
  nor_x1_sg U49456 ( .A(n23365), .B(n23366), .X(n23360) );
  nor_x1_sg U49457 ( .A(n23354), .B(n23355), .X(n23349) );
  inv_x1_sg U49458 ( .A(n23338), .X(n47481) );
  nand_x1_sg U49459 ( .A(n23340), .B(n23341), .X(n23338) );
  inv_x1_sg U49460 ( .A(n23324), .X(n47518) );
  nand_x1_sg U49461 ( .A(n23326), .B(n23327), .X(n23324) );
  inv_x1_sg U49462 ( .A(n23310), .X(n47558) );
  nand_x1_sg U49463 ( .A(n23312), .B(n23313), .X(n23310) );
  nand_x1_sg U49464 ( .A(n23298), .B(n23299), .X(n23296) );
  inv_x1_sg U49465 ( .A(n23663), .X(n47720) );
  nor_x1_sg U49466 ( .A(n23640), .B(n23641), .X(n23636) );
  nor_x1_sg U49467 ( .A(n23644), .B(n23645), .X(n23639) );
  nor_x1_sg U49468 ( .A(n23633), .B(n23634), .X(n23628) );
  inv_x1_sg U49469 ( .A(n23617), .X(n47766) );
  nand_x1_sg U49470 ( .A(n23619), .B(n23620), .X(n23617) );
  inv_x1_sg U49471 ( .A(n23603), .X(n47803) );
  nand_x1_sg U49472 ( .A(n23605), .B(n23606), .X(n23603) );
  inv_x1_sg U49473 ( .A(n23589), .X(n47843) );
  nand_x1_sg U49474 ( .A(n23591), .B(n23592), .X(n23589) );
  nand_x1_sg U49475 ( .A(n23577), .B(n23578), .X(n23575) );
  inv_x1_sg U49476 ( .A(n23942), .X(n48005) );
  nor_x1_sg U49477 ( .A(n23919), .B(n23920), .X(n23915) );
  nor_x1_sg U49478 ( .A(n23923), .B(n23924), .X(n23918) );
  nor_x1_sg U49479 ( .A(n23912), .B(n23913), .X(n23907) );
  inv_x1_sg U49480 ( .A(n23896), .X(n48051) );
  nand_x1_sg U49481 ( .A(n23898), .B(n23899), .X(n23896) );
  inv_x1_sg U49482 ( .A(n23882), .X(n48088) );
  nand_x1_sg U49483 ( .A(n23884), .B(n23885), .X(n23882) );
  inv_x1_sg U49484 ( .A(n23868), .X(n48128) );
  nand_x1_sg U49485 ( .A(n23870), .B(n23871), .X(n23868) );
  nand_x1_sg U49486 ( .A(n23856), .B(n23857), .X(n23854) );
  inv_x1_sg U49487 ( .A(n24221), .X(n48290) );
  nor_x1_sg U49488 ( .A(n24198), .B(n24199), .X(n24194) );
  nor_x1_sg U49489 ( .A(n24202), .B(n24203), .X(n24197) );
  nor_x1_sg U49490 ( .A(n24191), .B(n24192), .X(n24186) );
  inv_x1_sg U49491 ( .A(n24175), .X(n48336) );
  nand_x1_sg U49492 ( .A(n24177), .B(n24178), .X(n24175) );
  inv_x1_sg U49493 ( .A(n24147), .X(n48413) );
  nand_x1_sg U49494 ( .A(n24149), .B(n24150), .X(n24147) );
  nand_x1_sg U49495 ( .A(n24135), .B(n24136), .X(n24133) );
  inv_x1_sg U49496 ( .A(n24500), .X(n48575) );
  nor_x1_sg U49497 ( .A(n24477), .B(n24478), .X(n24473) );
  nor_x1_sg U49498 ( .A(n24481), .B(n24482), .X(n24476) );
  nor_x1_sg U49499 ( .A(n24470), .B(n24471), .X(n24465) );
  inv_x1_sg U49500 ( .A(n24454), .X(n48621) );
  nand_x1_sg U49501 ( .A(n24456), .B(n24457), .X(n24454) );
  inv_x1_sg U49502 ( .A(n24440), .X(n48658) );
  nand_x1_sg U49503 ( .A(n24442), .B(n24443), .X(n24440) );
  inv_x1_sg U49504 ( .A(n24426), .X(n48698) );
  nand_x1_sg U49505 ( .A(n24428), .B(n24429), .X(n24426) );
  nand_x1_sg U49506 ( .A(n24414), .B(n24415), .X(n24412) );
  inv_x1_sg U49507 ( .A(n24778), .X(n48861) );
  nor_x1_sg U49508 ( .A(n24755), .B(n24756), .X(n24751) );
  nor_x1_sg U49509 ( .A(n24759), .B(n24760), .X(n24754) );
  nor_x1_sg U49510 ( .A(n24748), .B(n24749), .X(n24743) );
  inv_x1_sg U49511 ( .A(n24732), .X(n48907) );
  nand_x1_sg U49512 ( .A(n24734), .B(n24735), .X(n24732) );
  inv_x1_sg U49513 ( .A(n24718), .X(n48944) );
  nand_x1_sg U49514 ( .A(n24720), .B(n24721), .X(n24718) );
  inv_x1_sg U49515 ( .A(n24704), .X(n48984) );
  nand_x1_sg U49516 ( .A(n24706), .B(n24707), .X(n24704) );
  nand_x1_sg U49517 ( .A(n24692), .B(n24693), .X(n24690) );
  inv_x1_sg U49518 ( .A(n25057), .X(n49148) );
  nor_x1_sg U49519 ( .A(n25034), .B(n25035), .X(n25030) );
  nor_x1_sg U49520 ( .A(n25038), .B(n25039), .X(n25033) );
  nor_x1_sg U49521 ( .A(n25027), .B(n25028), .X(n25022) );
  inv_x1_sg U49522 ( .A(n25011), .X(n49194) );
  nand_x1_sg U49523 ( .A(n25013), .B(n25014), .X(n25011) );
  inv_x1_sg U49524 ( .A(n24997), .X(n49231) );
  nand_x1_sg U49525 ( .A(n24999), .B(n25000), .X(n24997) );
  inv_x1_sg U49526 ( .A(n24983), .X(n49271) );
  nand_x1_sg U49527 ( .A(n24985), .B(n24986), .X(n24983) );
  nand_x1_sg U49528 ( .A(n24971), .B(n24972), .X(n24969) );
  inv_x1_sg U49529 ( .A(n25336), .X(n49434) );
  nor_x1_sg U49530 ( .A(n25313), .B(n25314), .X(n25309) );
  nor_x1_sg U49531 ( .A(n25317), .B(n25318), .X(n25312) );
  nor_x1_sg U49532 ( .A(n25306), .B(n25307), .X(n25301) );
  inv_x1_sg U49533 ( .A(n25290), .X(n49480) );
  nand_x1_sg U49534 ( .A(n25292), .B(n25293), .X(n25290) );
  inv_x1_sg U49535 ( .A(n25276), .X(n49517) );
  nand_x1_sg U49536 ( .A(n25278), .B(n25279), .X(n25276) );
  inv_x1_sg U49537 ( .A(n25262), .X(n49557) );
  nand_x1_sg U49538 ( .A(n25264), .B(n25265), .X(n25262) );
  nand_x1_sg U49539 ( .A(n25250), .B(n25251), .X(n25248) );
  inv_x1_sg U49540 ( .A(n25615), .X(n49719) );
  nor_x1_sg U49541 ( .A(n25592), .B(n25593), .X(n25588) );
  nor_x1_sg U49542 ( .A(n25596), .B(n25597), .X(n25591) );
  nor_x1_sg U49543 ( .A(n25585), .B(n25586), .X(n25580) );
  inv_x1_sg U49544 ( .A(n25569), .X(n49766) );
  nand_x1_sg U49545 ( .A(n25571), .B(n25572), .X(n25569) );
  inv_x1_sg U49546 ( .A(n25555), .X(n49803) );
  nand_x1_sg U49547 ( .A(n25557), .B(n25558), .X(n25555) );
  inv_x1_sg U49548 ( .A(n25541), .X(n49843) );
  nand_x1_sg U49549 ( .A(n25543), .B(n25544), .X(n25541) );
  nand_x1_sg U49550 ( .A(n25529), .B(n25530), .X(n25527) );
  inv_x1_sg U49551 ( .A(n25892), .X(n50006) );
  nor_x1_sg U49552 ( .A(n25869), .B(n25870), .X(n25865) );
  nor_x1_sg U49553 ( .A(n25873), .B(n25874), .X(n25868) );
  nor_x1_sg U49554 ( .A(n25862), .B(n25863), .X(n25857) );
  inv_x1_sg U49555 ( .A(n25846), .X(n50052) );
  nand_x1_sg U49556 ( .A(n25848), .B(n25849), .X(n25846) );
  inv_x1_sg U49557 ( .A(n25832), .X(n50089) );
  nand_x1_sg U49558 ( .A(n25834), .B(n25835), .X(n25832) );
  inv_x1_sg U49559 ( .A(n25818), .X(n50129) );
  nand_x1_sg U49560 ( .A(n25820), .B(n25821), .X(n25818) );
  nand_x1_sg U49561 ( .A(n25806), .B(n25807), .X(n25804) );
  inv_x1_sg U49562 ( .A(n26110), .X(n50290) );
  nor_x1_sg U49563 ( .A(n26168), .B(n26169), .X(n26107) );
  nor_x1_sg U49564 ( .A(n26162), .B(n50310), .X(n26096) );
  inv_x1_sg U49565 ( .A(n26163), .X(n50310) );
  nor_x1_sg U49566 ( .A(n26097), .B(n26098), .X(n26095) );
  inv_x1_sg U49567 ( .A(n26179), .X(n50558) );
  nor_x1_sg U49568 ( .A(n26145), .B(n26146), .X(n26143) );
  nor_x1_sg U49569 ( .A(n26159), .B(n26160), .X(n26089) );
  inv_x1_sg U49570 ( .A(n26078), .X(n50356) );
  nand_x1_sg U49571 ( .A(n26086), .B(n26157), .X(n26078) );
  inv_x1_sg U49572 ( .A(n26066), .X(n50395) );
  nand_x1_sg U49573 ( .A(n26074), .B(n26155), .X(n26066) );
  inv_x1_sg U49574 ( .A(n26059), .X(n50413) );
  nand_x1_sg U49575 ( .A(n26068), .B(n26154), .X(n26059) );
  inv_x1_sg U49576 ( .A(n26054), .X(n50435) );
  nand_x1_sg U49577 ( .A(n26062), .B(n26153), .X(n26054) );
  inv_x1_sg U49578 ( .A(n26047), .X(n50453) );
  nand_x1_sg U49579 ( .A(n26056), .B(n26152), .X(n26047) );
  inv_x1_sg U49580 ( .A(n26042), .X(n50482) );
  nand_x1_sg U49581 ( .A(n26050), .B(n26151), .X(n26042) );
  nand_x1_sg U49582 ( .A(n26044), .B(n26150), .X(n26136) );
  inv_x1_sg U49583 ( .A(n26452), .X(n50580) );
  nor_x1_sg U49584 ( .A(n26429), .B(n26430), .X(n26425) );
  nor_x1_sg U49585 ( .A(n26433), .B(n26434), .X(n26428) );
  nor_x1_sg U49586 ( .A(n26422), .B(n26423), .X(n26417) );
  inv_x1_sg U49587 ( .A(n26406), .X(n50626) );
  nand_x1_sg U49588 ( .A(n26408), .B(n26409), .X(n26406) );
  inv_x1_sg U49589 ( .A(n26392), .X(n50663) );
  nand_x1_sg U49590 ( .A(n26394), .B(n26395), .X(n26392) );
  inv_x1_sg U49591 ( .A(n26378), .X(n50703) );
  nand_x1_sg U49592 ( .A(n26380), .B(n26381), .X(n26378) );
  nand_x1_sg U49593 ( .A(n26366), .B(n26367), .X(n26364) );
  inv_x1_sg U49594 ( .A(n26730), .X(n50867) );
  nor_x1_sg U49595 ( .A(n26707), .B(n26708), .X(n26703) );
  nor_x1_sg U49596 ( .A(n26711), .B(n26712), .X(n26706) );
  nor_x1_sg U49597 ( .A(n26700), .B(n26701), .X(n26695) );
  inv_x1_sg U49598 ( .A(n26684), .X(n50913) );
  nand_x1_sg U49599 ( .A(n26686), .B(n26687), .X(n26684) );
  inv_x1_sg U49600 ( .A(n26670), .X(n50950) );
  nand_x1_sg U49601 ( .A(n26672), .B(n26673), .X(n26670) );
  inv_x1_sg U49602 ( .A(n26656), .X(n50990) );
  nand_x1_sg U49603 ( .A(n26658), .B(n26659), .X(n26656) );
  nand_x1_sg U49604 ( .A(n26644), .B(n26645), .X(n26642) );
  nor_x1_sg U49605 ( .A(n46631), .B(n19136), .X(n19131) );
  inv_x1_sg U49606 ( .A(n19139), .X(n46631) );
  inv_x1_sg U49607 ( .A(n19134), .X(n46632) );
  nor_x1_sg U49608 ( .A(n46626), .B(n19523), .X(n19125) );
  inv_x1_sg U49609 ( .A(n19525), .X(n46626) );
  nor_x1_sg U49610 ( .A(n20972), .B(n46619), .X(n20566) );
  inv_x1_sg U49611 ( .A(n20973), .X(n46619) );
  nor_x1_sg U49612 ( .A(n46622), .B(n20963), .X(n20580) );
  inv_x1_sg U49613 ( .A(n20965), .X(n46622) );
  inv_x1_sg U49614 ( .A(n5979), .X(n46609) );
  inv_x1_sg U49615 ( .A(n6031), .X(n46571) );
  inv_x1_sg U49616 ( .A(n19930), .X(n46561) );
  inv_x1_sg U49617 ( .A(n6080), .X(n46522) );
  nor_x1_sg U49618 ( .A(n46475), .B(n20293), .X(n6119) );
  inv_x1_sg U49619 ( .A(n20295), .X(n46475) );
  inv_x1_sg U49620 ( .A(n21525), .X(n46466) );
  inv_x1_sg U49621 ( .A(n6172), .X(n46433) );
  inv_x1_sg U49622 ( .A(n21518), .X(n46419) );
  nor_x1_sg U49623 ( .A(n46384), .B(n19300), .X(n6216) );
  inv_x1_sg U49624 ( .A(n19302), .X(n46384) );
  inv_x1_sg U49625 ( .A(n20283), .X(n46380) );
  inv_x1_sg U49626 ( .A(n21512), .X(n46371) );
  inv_x1_sg U49627 ( .A(n21505), .X(n46330) );
  inv_x1_sg U49628 ( .A(n21499), .X(n46284) );
  inv_x1_sg U49629 ( .A(n21492), .X(n46239) );
  inv_x1_sg U49630 ( .A(n21486), .X(n46193) );
  inv_x1_sg U49631 ( .A(n21479), .X(n46148) );
  inv_x1_sg U49632 ( .A(n21473), .X(n46102) );
  inv_x1_sg U49633 ( .A(n21466), .X(n46057) );
  inv_x1_sg U49634 ( .A(n21460), .X(n46011) );
  inv_x1_sg U49635 ( .A(n21453), .X(n45966) );
  inv_x1_sg U49636 ( .A(n6667), .X(n45930) );
  inv_x1_sg U49637 ( .A(n6758), .X(n45868) );
  nor_x1_sg U49638 ( .A(n20200), .B(n45844), .X(n6748) );
  inv_x1_sg U49639 ( .A(n20201), .X(n45844) );
  nor_x1_sg U49640 ( .A(n21431), .B(n45816), .X(n6771) );
  inv_x1_sg U49641 ( .A(n21432), .X(n45816) );
  nor_x1_sg U49642 ( .A(n20843), .B(n45828), .X(n6782) );
  inv_x1_sg U49643 ( .A(n20844), .X(n45828) );
  nor_x1_sg U49644 ( .A(n19214), .B(n19215), .X(n6802) );
  nand_x1_sg U49645 ( .A(n7070), .B(n46860), .X(n6848) );
  nor_x1_sg U49646 ( .A(n7080), .B(n7081), .X(n6854) );
  nand_x1_sg U49647 ( .A(n7105), .B(n46882), .X(n7090) );
  nand_x1_sg U49648 ( .A(n7091), .B(n7092), .X(n7089) );
  nand_x1_sg U49649 ( .A(n7168), .B(n7169), .X(n7148) );
  nand_x1_sg U49650 ( .A(n7231), .B(n7232), .X(n7200) );
  nand_x1_sg U49651 ( .A(n7201), .B(n7194), .X(n7199) );
  nand_x1_sg U49652 ( .A(n46947), .B(n7220), .X(n7201) );
  nand_x1_sg U49653 ( .A(n7238), .B(n7239), .X(n7236) );
  nand_x1_sg U49654 ( .A(n47014), .B(n7310), .X(n7265) );
  nand_x1_sg U49655 ( .A(n7266), .B(n7267), .X(n7264) );
  nand_x1_sg U49656 ( .A(n46999), .B(n42255), .X(n7267) );
  nand_x1_sg U49657 ( .A(n7317), .B(n7318), .X(n7315) );
  nand_x1_sg U49658 ( .A(n47068), .B(n7402), .X(n7351) );
  nand_x1_sg U49659 ( .A(n7352), .B(n7353), .X(n7350) );
  nand_x1_sg U49660 ( .A(n47039), .B(n42254), .X(n7353) );
  nand_x1_sg U49661 ( .A(n7450), .B(n47090), .X(n7408) );
  nand_x1_sg U49662 ( .A(n7409), .B(n7410), .X(n7407) );
  nand_x1_sg U49663 ( .A(n7514), .B(n47114), .X(n7456) );
  nand_x1_sg U49664 ( .A(n7457), .B(n7458), .X(n7455) );
  nand_x1_sg U49665 ( .A(n47089), .B(n7452), .X(n7458) );
  inv_x1_sg U49666 ( .A(n6973), .X(n47124) );
  nand_x1_sg U49667 ( .A(n47098), .B(n6967), .X(n6965) );
  nor_x1_sg U49668 ( .A(n6937), .B(n6938), .X(n6935) );
  nand_x1_sg U49669 ( .A(n47046), .B(n6951), .X(n6936) );
  nand_x1_sg U49670 ( .A(n7888), .B(n47153), .X(n7665) );
  nor_x1_sg U49671 ( .A(n7898), .B(n7899), .X(n7671) );
  nand_x1_sg U49672 ( .A(n7923), .B(n47175), .X(n7908) );
  nand_x1_sg U49673 ( .A(n7909), .B(n7910), .X(n7907) );
  nand_x1_sg U49674 ( .A(n7987), .B(n7988), .X(n7966) );
  nand_x1_sg U49675 ( .A(n8050), .B(n8051), .X(n8019) );
  nand_x1_sg U49676 ( .A(n8020), .B(n8013), .X(n8018) );
  nand_x1_sg U49677 ( .A(n47238), .B(n8039), .X(n8020) );
  nand_x1_sg U49678 ( .A(n8057), .B(n8058), .X(n8055) );
  nand_x1_sg U49679 ( .A(n47302), .B(n8128), .X(n8084) );
  nand_x1_sg U49680 ( .A(n8135), .B(n8136), .X(n8133) );
  nand_x1_sg U49681 ( .A(n47354), .B(n8220), .X(n8169) );
  nand_x1_sg U49682 ( .A(n8170), .B(n8171), .X(n8168) );
  nand_x1_sg U49683 ( .A(n47326), .B(n42253), .X(n8171) );
  nand_x1_sg U49684 ( .A(n8268), .B(n47376), .X(n8226) );
  nand_x1_sg U49685 ( .A(n8227), .B(n8228), .X(n8225) );
  nand_x1_sg U49686 ( .A(n8332), .B(n47400), .X(n8274) );
  nand_x1_sg U49687 ( .A(n8275), .B(n8276), .X(n8273) );
  nand_x1_sg U49688 ( .A(n47375), .B(n8270), .X(n8276) );
  inv_x1_sg U49689 ( .A(n7790), .X(n47410) );
  nand_x1_sg U49690 ( .A(n47384), .B(n7784), .X(n7782) );
  nor_x1_sg U49691 ( .A(n7754), .B(n7755), .X(n7752) );
  nand_x1_sg U49692 ( .A(n47333), .B(n7768), .X(n7753) );
  nand_x1_sg U49693 ( .A(n8706), .B(n47438), .X(n8483) );
  nor_x1_sg U49694 ( .A(n8716), .B(n8717), .X(n8489) );
  nand_x1_sg U49695 ( .A(n8741), .B(n47460), .X(n8726) );
  nand_x1_sg U49696 ( .A(n8727), .B(n8728), .X(n8725) );
  nand_x1_sg U49697 ( .A(n8805), .B(n8806), .X(n8784) );
  nand_x1_sg U49698 ( .A(n8868), .B(n8869), .X(n8837) );
  nand_x1_sg U49699 ( .A(n8838), .B(n8831), .X(n8836) );
  nand_x1_sg U49700 ( .A(n47523), .B(n8857), .X(n8838) );
  nand_x1_sg U49701 ( .A(n8875), .B(n8876), .X(n8873) );
  nand_x1_sg U49702 ( .A(n47587), .B(n8946), .X(n8902) );
  nand_x1_sg U49703 ( .A(n8953), .B(n8954), .X(n8951) );
  nand_x1_sg U49704 ( .A(n47639), .B(n9038), .X(n8987) );
  nand_x1_sg U49705 ( .A(n8988), .B(n8989), .X(n8986) );
  nand_x1_sg U49706 ( .A(n47611), .B(n42252), .X(n8989) );
  nand_x1_sg U49707 ( .A(n9086), .B(n47661), .X(n9044) );
  nand_x1_sg U49708 ( .A(n9045), .B(n9046), .X(n9043) );
  nand_x1_sg U49709 ( .A(n9150), .B(n47685), .X(n9092) );
  nand_x1_sg U49710 ( .A(n9093), .B(n9094), .X(n9091) );
  nand_x1_sg U49711 ( .A(n47660), .B(n9088), .X(n9094) );
  inv_x1_sg U49712 ( .A(n8608), .X(n47695) );
  nand_x1_sg U49713 ( .A(n47669), .B(n8602), .X(n8600) );
  nor_x1_sg U49714 ( .A(n8572), .B(n8573), .X(n8570) );
  nand_x1_sg U49715 ( .A(n47618), .B(n8586), .X(n8571) );
  nand_x1_sg U49716 ( .A(n9526), .B(n47723), .X(n9303) );
  nor_x1_sg U49717 ( .A(n9536), .B(n9537), .X(n9309) );
  nand_x1_sg U49718 ( .A(n9561), .B(n47745), .X(n9546) );
  nand_x1_sg U49719 ( .A(n9547), .B(n9548), .X(n9545) );
  nand_x1_sg U49720 ( .A(n9625), .B(n9626), .X(n9604) );
  nand_x1_sg U49721 ( .A(n9688), .B(n9689), .X(n9657) );
  nand_x1_sg U49722 ( .A(n9658), .B(n9651), .X(n9656) );
  nand_x1_sg U49723 ( .A(n47808), .B(n9677), .X(n9658) );
  nand_x1_sg U49724 ( .A(n9695), .B(n9696), .X(n9693) );
  nand_x1_sg U49725 ( .A(n47872), .B(n9766), .X(n9722) );
  nand_x1_sg U49726 ( .A(n9773), .B(n9774), .X(n9771) );
  nand_x1_sg U49727 ( .A(n47924), .B(n9858), .X(n9807) );
  nand_x1_sg U49728 ( .A(n9808), .B(n9809), .X(n9806) );
  nand_x1_sg U49729 ( .A(n47896), .B(n42251), .X(n9809) );
  nand_x1_sg U49730 ( .A(n9906), .B(n47946), .X(n9864) );
  nand_x1_sg U49731 ( .A(n9865), .B(n9866), .X(n9863) );
  nand_x1_sg U49732 ( .A(n9970), .B(n47970), .X(n9912) );
  nand_x1_sg U49733 ( .A(n9913), .B(n9914), .X(n9911) );
  nand_x1_sg U49734 ( .A(n47945), .B(n9908), .X(n9914) );
  inv_x1_sg U49735 ( .A(n9428), .X(n47980) );
  nand_x1_sg U49736 ( .A(n47954), .B(n9422), .X(n9420) );
  nor_x1_sg U49737 ( .A(n9392), .B(n9393), .X(n9390) );
  nand_x1_sg U49738 ( .A(n47903), .B(n9406), .X(n9391) );
  nand_x1_sg U49739 ( .A(n10345), .B(n48008), .X(n10122) );
  nor_x1_sg U49740 ( .A(n10355), .B(n10356), .X(n10128) );
  nand_x1_sg U49741 ( .A(n10380), .B(n48030), .X(n10365) );
  nand_x1_sg U49742 ( .A(n10366), .B(n10367), .X(n10364) );
  nand_x1_sg U49743 ( .A(n10444), .B(n10445), .X(n10423) );
  nand_x1_sg U49744 ( .A(n10507), .B(n10508), .X(n10476) );
  nand_x1_sg U49745 ( .A(n10477), .B(n10470), .X(n10475) );
  nand_x1_sg U49746 ( .A(n48093), .B(n10496), .X(n10477) );
  nand_x1_sg U49747 ( .A(n10514), .B(n10515), .X(n10512) );
  nand_x1_sg U49748 ( .A(n48157), .B(n10585), .X(n10541) );
  nand_x1_sg U49749 ( .A(n10592), .B(n10593), .X(n10590) );
  nand_x1_sg U49750 ( .A(n48209), .B(n10677), .X(n10626) );
  nand_x1_sg U49751 ( .A(n10627), .B(n10628), .X(n10625) );
  nand_x1_sg U49752 ( .A(n48181), .B(n42250), .X(n10628) );
  nand_x1_sg U49753 ( .A(n10725), .B(n48231), .X(n10683) );
  nand_x1_sg U49754 ( .A(n10684), .B(n10685), .X(n10682) );
  nand_x1_sg U49755 ( .A(n10789), .B(n48255), .X(n10731) );
  nand_x1_sg U49756 ( .A(n10732), .B(n10733), .X(n10730) );
  nand_x1_sg U49757 ( .A(n48230), .B(n10727), .X(n10733) );
  inv_x1_sg U49758 ( .A(n10247), .X(n48265) );
  nand_x1_sg U49759 ( .A(n48239), .B(n10241), .X(n10239) );
  nor_x1_sg U49760 ( .A(n10211), .B(n10212), .X(n10209) );
  nand_x1_sg U49761 ( .A(n48188), .B(n10225), .X(n10210) );
  nand_x1_sg U49762 ( .A(n11164), .B(n48293), .X(n10941) );
  nor_x1_sg U49763 ( .A(n11174), .B(n11175), .X(n10947) );
  nand_x1_sg U49764 ( .A(n11199), .B(n48315), .X(n11184) );
  nand_x1_sg U49765 ( .A(n11185), .B(n11186), .X(n11183) );
  nand_x1_sg U49766 ( .A(n11263), .B(n11264), .X(n11242) );
  nand_x1_sg U49767 ( .A(n11326), .B(n11327), .X(n11295) );
  nand_x1_sg U49768 ( .A(n11296), .B(n11289), .X(n11294) );
  nand_x1_sg U49769 ( .A(n48378), .B(n11315), .X(n11296) );
  nand_x1_sg U49770 ( .A(n11333), .B(n11334), .X(n11331) );
  nand_x1_sg U49771 ( .A(n48442), .B(n11404), .X(n11360) );
  nand_x1_sg U49772 ( .A(n11411), .B(n11412), .X(n11409) );
  nand_x1_sg U49773 ( .A(n48494), .B(n11496), .X(n11445) );
  nand_x1_sg U49774 ( .A(n11446), .B(n11447), .X(n11444) );
  nand_x1_sg U49775 ( .A(n48466), .B(n42249), .X(n11447) );
  nand_x1_sg U49776 ( .A(n11544), .B(n48516), .X(n11502) );
  nand_x1_sg U49777 ( .A(n11503), .B(n11504), .X(n11501) );
  nand_x1_sg U49778 ( .A(n11608), .B(n48540), .X(n11550) );
  nand_x1_sg U49779 ( .A(n11551), .B(n11552), .X(n11549) );
  nand_x1_sg U49780 ( .A(n48515), .B(n11546), .X(n11552) );
  inv_x1_sg U49781 ( .A(n11066), .X(n48550) );
  nand_x1_sg U49782 ( .A(n48524), .B(n11060), .X(n11058) );
  nor_x1_sg U49783 ( .A(n11030), .B(n11031), .X(n11028) );
  nand_x1_sg U49784 ( .A(n48473), .B(n11044), .X(n11029) );
  nand_x1_sg U49785 ( .A(n11983), .B(n48578), .X(n11760) );
  nor_x1_sg U49786 ( .A(n11993), .B(n11994), .X(n11766) );
  nand_x1_sg U49787 ( .A(n12018), .B(n48600), .X(n12003) );
  nand_x1_sg U49788 ( .A(n12004), .B(n12005), .X(n12002) );
  nand_x1_sg U49789 ( .A(n12082), .B(n12083), .X(n12061) );
  nand_x1_sg U49790 ( .A(n12145), .B(n12146), .X(n12114) );
  nand_x1_sg U49791 ( .A(n12115), .B(n12108), .X(n12113) );
  nand_x1_sg U49792 ( .A(n48663), .B(n12134), .X(n12115) );
  nand_x1_sg U49793 ( .A(n12152), .B(n12153), .X(n12150) );
  nand_x1_sg U49794 ( .A(n48727), .B(n12223), .X(n12179) );
  nand_x1_sg U49795 ( .A(n12230), .B(n12231), .X(n12228) );
  nand_x1_sg U49796 ( .A(n48779), .B(n12315), .X(n12264) );
  nand_x1_sg U49797 ( .A(n12265), .B(n12266), .X(n12263) );
  nand_x1_sg U49798 ( .A(n48751), .B(n42248), .X(n12266) );
  nand_x1_sg U49799 ( .A(n12363), .B(n48801), .X(n12321) );
  nand_x1_sg U49800 ( .A(n12322), .B(n12323), .X(n12320) );
  nand_x1_sg U49801 ( .A(n12427), .B(n48825), .X(n12369) );
  nand_x1_sg U49802 ( .A(n12370), .B(n12371), .X(n12368) );
  nand_x1_sg U49803 ( .A(n48800), .B(n12365), .X(n12371) );
  inv_x1_sg U49804 ( .A(n11885), .X(n48835) );
  nand_x1_sg U49805 ( .A(n48809), .B(n11879), .X(n11877) );
  nor_x1_sg U49806 ( .A(n11849), .B(n11850), .X(n11847) );
  nand_x1_sg U49807 ( .A(n48758), .B(n11863), .X(n11848) );
  nand_x1_sg U49808 ( .A(n12802), .B(n48864), .X(n12579) );
  nor_x1_sg U49809 ( .A(n12812), .B(n12813), .X(n12585) );
  nand_x1_sg U49810 ( .A(n12837), .B(n48886), .X(n12822) );
  nand_x1_sg U49811 ( .A(n12823), .B(n12824), .X(n12821) );
  nand_x1_sg U49812 ( .A(n12901), .B(n12902), .X(n12880) );
  nand_x1_sg U49813 ( .A(n12964), .B(n12965), .X(n12933) );
  nand_x1_sg U49814 ( .A(n12934), .B(n12927), .X(n12932) );
  nand_x1_sg U49815 ( .A(n48949), .B(n12953), .X(n12934) );
  nand_x1_sg U49816 ( .A(n12971), .B(n12972), .X(n12969) );
  nand_x1_sg U49817 ( .A(n49013), .B(n13042), .X(n12998) );
  nand_x1_sg U49818 ( .A(n13049), .B(n13050), .X(n13047) );
  nand_x1_sg U49819 ( .A(n49066), .B(n13134), .X(n13083) );
  nand_x1_sg U49820 ( .A(n13084), .B(n13085), .X(n13082) );
  nand_x1_sg U49821 ( .A(n49037), .B(n42247), .X(n13085) );
  nand_x1_sg U49822 ( .A(n13182), .B(n49088), .X(n13140) );
  nand_x1_sg U49823 ( .A(n13141), .B(n13142), .X(n13139) );
  nand_x1_sg U49824 ( .A(n13246), .B(n49112), .X(n13188) );
  nand_x1_sg U49825 ( .A(n13189), .B(n13190), .X(n13187) );
  nand_x1_sg U49826 ( .A(n49087), .B(n13184), .X(n13190) );
  inv_x1_sg U49827 ( .A(n12704), .X(n49122) );
  nand_x1_sg U49828 ( .A(n49096), .B(n12698), .X(n12696) );
  nor_x1_sg U49829 ( .A(n12668), .B(n12669), .X(n12666) );
  nand_x1_sg U49830 ( .A(n49044), .B(n12682), .X(n12667) );
  nand_x1_sg U49831 ( .A(n13621), .B(n49151), .X(n13398) );
  nor_x1_sg U49832 ( .A(n13631), .B(n13632), .X(n13404) );
  nand_x1_sg U49833 ( .A(n13656), .B(n49173), .X(n13641) );
  nand_x1_sg U49834 ( .A(n13642), .B(n13643), .X(n13640) );
  nand_x1_sg U49835 ( .A(n13720), .B(n13721), .X(n13699) );
  nand_x1_sg U49836 ( .A(n13783), .B(n13784), .X(n13752) );
  nand_x1_sg U49837 ( .A(n13753), .B(n13746), .X(n13751) );
  nand_x1_sg U49838 ( .A(n49236), .B(n13772), .X(n13753) );
  nand_x1_sg U49839 ( .A(n13790), .B(n13791), .X(n13788) );
  nand_x1_sg U49840 ( .A(n49300), .B(n13861), .X(n13817) );
  nand_x1_sg U49841 ( .A(n13868), .B(n13869), .X(n13866) );
  nand_x1_sg U49842 ( .A(n49352), .B(n13953), .X(n13902) );
  nand_x1_sg U49843 ( .A(n13903), .B(n13904), .X(n13901) );
  nand_x1_sg U49844 ( .A(n49324), .B(n42246), .X(n13904) );
  nand_x1_sg U49845 ( .A(n14001), .B(n49374), .X(n13959) );
  nand_x1_sg U49846 ( .A(n13960), .B(n13961), .X(n13958) );
  nand_x1_sg U49847 ( .A(n14065), .B(n49398), .X(n14007) );
  nand_x1_sg U49848 ( .A(n14008), .B(n14009), .X(n14006) );
  nand_x1_sg U49849 ( .A(n49373), .B(n14003), .X(n14009) );
  inv_x1_sg U49850 ( .A(n13523), .X(n49408) );
  nand_x1_sg U49851 ( .A(n49382), .B(n13517), .X(n13515) );
  nor_x1_sg U49852 ( .A(n13487), .B(n13488), .X(n13485) );
  nand_x1_sg U49853 ( .A(n49331), .B(n13501), .X(n13486) );
  nand_x1_sg U49854 ( .A(n14440), .B(n49437), .X(n14217) );
  nor_x1_sg U49855 ( .A(n14450), .B(n14451), .X(n14223) );
  nand_x1_sg U49856 ( .A(n14475), .B(n49459), .X(n14460) );
  nand_x1_sg U49857 ( .A(n14461), .B(n14462), .X(n14459) );
  nand_x1_sg U49858 ( .A(n14539), .B(n14540), .X(n14518) );
  nand_x1_sg U49859 ( .A(n14602), .B(n14603), .X(n14571) );
  nand_x1_sg U49860 ( .A(n14572), .B(n14565), .X(n14570) );
  nand_x1_sg U49861 ( .A(n49522), .B(n14591), .X(n14572) );
  nand_x1_sg U49862 ( .A(n14609), .B(n14610), .X(n14607) );
  nand_x1_sg U49863 ( .A(n49586), .B(n14680), .X(n14636) );
  nand_x1_sg U49864 ( .A(n14687), .B(n14688), .X(n14685) );
  nand_x1_sg U49865 ( .A(n49638), .B(n14772), .X(n14721) );
  nand_x1_sg U49866 ( .A(n14722), .B(n14723), .X(n14720) );
  nand_x1_sg U49867 ( .A(n49610), .B(n42245), .X(n14723) );
  nand_x1_sg U49868 ( .A(n14820), .B(n49660), .X(n14778) );
  nand_x1_sg U49869 ( .A(n14779), .B(n14780), .X(n14777) );
  nand_x1_sg U49870 ( .A(n14884), .B(n49684), .X(n14826) );
  nand_x1_sg U49871 ( .A(n14827), .B(n14828), .X(n14825) );
  nand_x1_sg U49872 ( .A(n49659), .B(n14822), .X(n14828) );
  inv_x1_sg U49873 ( .A(n14342), .X(n49694) );
  nand_x1_sg U49874 ( .A(n49668), .B(n14336), .X(n14334) );
  nor_x1_sg U49875 ( .A(n14306), .B(n14307), .X(n14304) );
  nand_x1_sg U49876 ( .A(n49617), .B(n14320), .X(n14305) );
  nand_x1_sg U49877 ( .A(n15259), .B(n49722), .X(n15036) );
  nor_x1_sg U49878 ( .A(n15269), .B(n15270), .X(n15042) );
  nand_x1_sg U49879 ( .A(n15294), .B(n49744), .X(n15279) );
  nand_x1_sg U49880 ( .A(n15280), .B(n15281), .X(n15278) );
  nand_x1_sg U49881 ( .A(n15358), .B(n15359), .X(n15337) );
  nand_x1_sg U49882 ( .A(n15421), .B(n15422), .X(n15390) );
  nand_x1_sg U49883 ( .A(n15391), .B(n15384), .X(n15389) );
  nand_x1_sg U49884 ( .A(n49808), .B(n15410), .X(n15391) );
  nand_x1_sg U49885 ( .A(n15428), .B(n15429), .X(n15426) );
  nand_x1_sg U49886 ( .A(n49872), .B(n15499), .X(n15455) );
  nand_x1_sg U49887 ( .A(n15506), .B(n15507), .X(n15504) );
  nand_x1_sg U49888 ( .A(n49924), .B(n15591), .X(n15540) );
  nand_x1_sg U49889 ( .A(n15541), .B(n15542), .X(n15539) );
  nand_x1_sg U49890 ( .A(n49896), .B(n42244), .X(n15542) );
  nand_x1_sg U49891 ( .A(n15639), .B(n49946), .X(n15597) );
  nand_x1_sg U49892 ( .A(n15598), .B(n15599), .X(n15596) );
  nand_x1_sg U49893 ( .A(n15703), .B(n49970), .X(n15645) );
  nand_x1_sg U49894 ( .A(n15646), .B(n15647), .X(n15644) );
  nand_x1_sg U49895 ( .A(n49945), .B(n15641), .X(n15647) );
  inv_x1_sg U49896 ( .A(n15161), .X(n49980) );
  nand_x1_sg U49897 ( .A(n49954), .B(n15155), .X(n15153) );
  nor_x1_sg U49898 ( .A(n15125), .B(n15126), .X(n15123) );
  nand_x1_sg U49899 ( .A(n49903), .B(n15139), .X(n15124) );
  nand_x1_sg U49900 ( .A(n16078), .B(n50009), .X(n15855) );
  nor_x1_sg U49901 ( .A(n16088), .B(n16089), .X(n15861) );
  nand_x1_sg U49902 ( .A(n16113), .B(n50031), .X(n16098) );
  nand_x1_sg U49903 ( .A(n16099), .B(n16100), .X(n16097) );
  nand_x1_sg U49904 ( .A(n16177), .B(n16178), .X(n16156) );
  nand_x1_sg U49905 ( .A(n16240), .B(n16241), .X(n16209) );
  nand_x1_sg U49906 ( .A(n16210), .B(n16203), .X(n16208) );
  nand_x1_sg U49907 ( .A(n50094), .B(n16229), .X(n16210) );
  nand_x1_sg U49908 ( .A(n16247), .B(n16248), .X(n16245) );
  nand_x1_sg U49909 ( .A(n50158), .B(n16318), .X(n16274) );
  nand_x1_sg U49910 ( .A(n16325), .B(n16326), .X(n16323) );
  nand_x1_sg U49911 ( .A(n50210), .B(n16410), .X(n16359) );
  nand_x1_sg U49912 ( .A(n16360), .B(n16361), .X(n16358) );
  nand_x1_sg U49913 ( .A(n50182), .B(n42243), .X(n16361) );
  nand_x1_sg U49914 ( .A(n16458), .B(n50232), .X(n16416) );
  nand_x1_sg U49915 ( .A(n16417), .B(n16418), .X(n16415) );
  nand_x1_sg U49916 ( .A(n16522), .B(n50256), .X(n16464) );
  nand_x1_sg U49917 ( .A(n16465), .B(n16466), .X(n16463) );
  nand_x1_sg U49918 ( .A(n50231), .B(n16460), .X(n16466) );
  inv_x1_sg U49919 ( .A(n15980), .X(n50266) );
  nand_x1_sg U49920 ( .A(n50240), .B(n15974), .X(n15972) );
  nor_x1_sg U49921 ( .A(n15944), .B(n15945), .X(n15942) );
  nand_x1_sg U49922 ( .A(n50189), .B(n15958), .X(n15943) );
  nand_x1_sg U49923 ( .A(n26126), .B(n26127), .X(n26125) );
  nand_x1_sg U49924 ( .A(n16897), .B(n50293), .X(n16672) );
  nor_x1_sg U49925 ( .A(n16907), .B(n16908), .X(n16678) );
  nand_x1_sg U49926 ( .A(n16930), .B(n50316), .X(n16916) );
  nand_x1_sg U49927 ( .A(n16917), .B(n16918), .X(n16915) );
  nand_x1_sg U49928 ( .A(n16993), .B(n16994), .X(n16973) );
  nand_x1_sg U49929 ( .A(n17056), .B(n17057), .X(n17025) );
  nand_x1_sg U49930 ( .A(n17026), .B(n17019), .X(n17024) );
  nand_x1_sg U49931 ( .A(n50379), .B(n17045), .X(n17026) );
  nand_x1_sg U49932 ( .A(n17063), .B(n17064), .X(n17061) );
  nand_x1_sg U49933 ( .A(n50443), .B(n17135), .X(n17090) );
  nand_x1_sg U49934 ( .A(n17091), .B(n17092), .X(n17089) );
  nand_x1_sg U49935 ( .A(n50429), .B(n42242), .X(n17092) );
  nand_x1_sg U49936 ( .A(n17142), .B(n17143), .X(n17140) );
  nand_x1_sg U49937 ( .A(n50495), .B(n17227), .X(n17176) );
  nand_x1_sg U49938 ( .A(n17177), .B(n17178), .X(n17175) );
  nand_x1_sg U49939 ( .A(n50467), .B(n42241), .X(n17178) );
  nand_x1_sg U49940 ( .A(n17275), .B(n50517), .X(n17233) );
  nand_x1_sg U49941 ( .A(n17234), .B(n17235), .X(n17232) );
  nand_x1_sg U49942 ( .A(n17339), .B(n50541), .X(n17281) );
  nand_x1_sg U49943 ( .A(n17282), .B(n17283), .X(n17280) );
  nand_x1_sg U49944 ( .A(n50516), .B(n17277), .X(n17283) );
  inv_x1_sg U49945 ( .A(n16797), .X(n50552) );
  nand_x1_sg U49946 ( .A(n50526), .B(n16791), .X(n16789) );
  nor_x1_sg U49947 ( .A(n16761), .B(n16762), .X(n16759) );
  nand_x1_sg U49948 ( .A(n50474), .B(n16775), .X(n16760) );
  nand_x1_sg U49949 ( .A(n17716), .B(n50583), .X(n17493) );
  nor_x1_sg U49950 ( .A(n17726), .B(n17727), .X(n17499) );
  nand_x1_sg U49951 ( .A(n17751), .B(n50605), .X(n17736) );
  nand_x1_sg U49952 ( .A(n17737), .B(n17738), .X(n17735) );
  nand_x1_sg U49953 ( .A(n17815), .B(n17816), .X(n17794) );
  nand_x1_sg U49954 ( .A(n17878), .B(n17879), .X(n17847) );
  nand_x1_sg U49955 ( .A(n17848), .B(n17841), .X(n17846) );
  nand_x1_sg U49956 ( .A(n50668), .B(n17867), .X(n17848) );
  nand_x1_sg U49957 ( .A(n17885), .B(n17886), .X(n17883) );
  nand_x1_sg U49958 ( .A(n50732), .B(n17956), .X(n17912) );
  nand_x1_sg U49959 ( .A(n17963), .B(n17964), .X(n17961) );
  nand_x1_sg U49960 ( .A(n50784), .B(n18048), .X(n17997) );
  nand_x1_sg U49961 ( .A(n17998), .B(n17999), .X(n17996) );
  nand_x1_sg U49962 ( .A(n50756), .B(n42240), .X(n17999) );
  nand_x1_sg U49963 ( .A(n18096), .B(n50806), .X(n18054) );
  nand_x1_sg U49964 ( .A(n18055), .B(n18056), .X(n18053) );
  nand_x1_sg U49965 ( .A(n18160), .B(n50830), .X(n18102) );
  nand_x1_sg U49966 ( .A(n18103), .B(n18104), .X(n18101) );
  nand_x1_sg U49967 ( .A(n50805), .B(n18098), .X(n18104) );
  inv_x1_sg U49968 ( .A(n17618), .X(n50840) );
  nand_x1_sg U49969 ( .A(n50814), .B(n17612), .X(n17610) );
  nor_x1_sg U49970 ( .A(n17582), .B(n17583), .X(n17580) );
  nand_x1_sg U49971 ( .A(n50763), .B(n17596), .X(n17581) );
  nand_x1_sg U49972 ( .A(n18537), .B(n50870), .X(n18314) );
  nor_x1_sg U49973 ( .A(n18547), .B(n18548), .X(n18320) );
  nand_x1_sg U49974 ( .A(n18572), .B(n50892), .X(n18557) );
  nand_x1_sg U49975 ( .A(n18558), .B(n18559), .X(n18556) );
  nand_x1_sg U49976 ( .A(n18636), .B(n18637), .X(n18615) );
  nand_x1_sg U49977 ( .A(n18699), .B(n18700), .X(n18668) );
  nand_x1_sg U49978 ( .A(n18669), .B(n18662), .X(n18667) );
  nand_x1_sg U49979 ( .A(n50955), .B(n18688), .X(n18669) );
  nand_x1_sg U49980 ( .A(n18706), .B(n18707), .X(n18704) );
  nand_x1_sg U49981 ( .A(n51019), .B(n18777), .X(n18733) );
  nand_x1_sg U49982 ( .A(n18784), .B(n18785), .X(n18782) );
  nand_x1_sg U49983 ( .A(n51071), .B(n18869), .X(n18818) );
  nand_x1_sg U49984 ( .A(n18819), .B(n18820), .X(n18817) );
  nand_x1_sg U49985 ( .A(n51043), .B(n42239), .X(n18820) );
  nand_x1_sg U49986 ( .A(n18917), .B(n51093), .X(n18875) );
  nand_x1_sg U49987 ( .A(n18876), .B(n18877), .X(n18874) );
  nand_x1_sg U49988 ( .A(n18981), .B(n51117), .X(n18923) );
  nand_x1_sg U49989 ( .A(n18924), .B(n18925), .X(n18922) );
  nand_x1_sg U49990 ( .A(n51092), .B(n18919), .X(n18925) );
  inv_x1_sg U49991 ( .A(n18439), .X(n51127) );
  nand_x1_sg U49992 ( .A(n51101), .B(n18433), .X(n18431) );
  nor_x1_sg U49993 ( .A(n18403), .B(n18404), .X(n18401) );
  nand_x1_sg U49994 ( .A(n51050), .B(n18417), .X(n18402) );
  inv_x1_sg U49995 ( .A(n28551), .X(n45780) );
  inv_x1_sg U49996 ( .A(n26831), .X(n45777) );
  inv_x1_sg U49997 ( .A(n26895), .X(n45769) );
  inv_x1_sg U49998 ( .A(n26888), .X(n45770) );
  nand_x2_sg U49999 ( .A(out_L1[18]), .B(n28539), .X(n28538) );
  nand_x1_sg U50000 ( .A(n28541), .B(n45782), .X(n28536) );
  inv_x1_sg U50001 ( .A(n28558), .X(n45779) );
  nand_x1_sg U50002 ( .A(n26775), .B(n26776), .X(n26774) );
  nand_x1_sg U50003 ( .A(n39260), .B(n26777), .X(n26776) );
  nand_x1_sg U50004 ( .A(n38932), .B(n26765), .X(n26764) );
  inv_x1_sg U50005 ( .A(n28544), .X(n45781) );
  inv_x1_sg U50006 ( .A(n28565), .X(n45778) );
  nand_x1_sg U50007 ( .A(n28750), .B(n28751), .X(n28731) );
  nand_x1_sg U50008 ( .A(n5361), .B(n28556), .X(n28751) );
  nand_x1_sg U50009 ( .A(n27088), .B(n27089), .X(n27081) );
  nand_x1_sg U50010 ( .A(n5304), .B(n26836), .X(n27089) );
  nand_x1_sg U50011 ( .A(n27137), .B(n27138), .X(n27057) );
  nand_x1_sg U50012 ( .A(n5152), .B(n26893), .X(n27138) );
  nand_x1_sg U50013 ( .A(n21760), .B(n21761), .X(n21759) );
  nand_x1_sg U50014 ( .A(n5133), .B(n21762), .X(n21761) );
  nor_x1_sg U50015 ( .A(n28742), .B(n28743), .X(n28736) );
  nand_x1_sg U50016 ( .A(n28756), .B(n28757), .X(n28728) );
  nand_x1_sg U50017 ( .A(n5342), .B(n28563), .X(n28757) );
  nand_x1_sg U50018 ( .A(n21739), .B(n21740), .X(n21738) );
  nand_x1_sg U50019 ( .A(n28744), .B(n28745), .X(n28734) );
  nand_x1_sg U50020 ( .A(n5380), .B(n28549), .X(n28745) );
  nand_x1_sg U50021 ( .A(n27085), .B(n27086), .X(n27084) );
  nand_x1_sg U50022 ( .A(n5323), .B(n27087), .X(n27086) );
  nand_x1_sg U50023 ( .A(n28929), .B(n28930), .X(n28910) );
  nand_x1_sg U50024 ( .A(n5362), .B(n28755), .X(n28930) );
  nand_x1_sg U50025 ( .A(n27318), .B(n27319), .X(n27311) );
  nand_x1_sg U50026 ( .A(n5305), .B(n27093), .X(n27319) );
  nand_x1_sg U50027 ( .A(n27052), .B(n27053), .X(n27051) );
  nand_x1_sg U50028 ( .A(n5153), .B(n27054), .X(n27053) );
  nand_x1_sg U50029 ( .A(n21807), .B(n21808), .X(n21806) );
  nand_x1_sg U50030 ( .A(n5134), .B(n21809), .X(n21808) );
  nand_x1_sg U50031 ( .A(n42086), .B(n28921), .X(n28916) );
  nand_x1_sg U50032 ( .A(n28723), .B(n28724), .X(n28722) );
  nand_x1_sg U50033 ( .A(n5343), .B(n28725), .X(n28724) );
  nand_x1_sg U50034 ( .A(n21786), .B(n21787), .X(n21785) );
  nand_x1_sg U50035 ( .A(n28923), .B(n28924), .X(n28913) );
  nand_x1_sg U50036 ( .A(n5381), .B(n28749), .X(n28924) );
  nand_x1_sg U50037 ( .A(n27315), .B(n27316), .X(n27314) );
  nand_x1_sg U50038 ( .A(n5324), .B(n27317), .X(n27316) );
  nand_x1_sg U50039 ( .A(n28905), .B(n28906), .X(n28904) );
  nand_x1_sg U50040 ( .A(n5363), .B(n28907), .X(n28906) );
  nand_x1_sg U50041 ( .A(n27531), .B(n27532), .X(n27524) );
  nand_x1_sg U50042 ( .A(n5306), .B(n27323), .X(n27532) );
  nand_x1_sg U50043 ( .A(n27046), .B(n27047), .X(n27045) );
  nand_x1_sg U50044 ( .A(n5154), .B(n27048), .X(n27047) );
  nand_x1_sg U50045 ( .A(n21854), .B(n21855), .X(n21853) );
  nand_x1_sg U50046 ( .A(n5135), .B(n21856), .X(n21855) );
  nand_x1_sg U50047 ( .A(n45652), .B(n29090), .X(n29085) );
  nand_x1_sg U50048 ( .A(n28717), .B(n28718), .X(n28716) );
  nand_x1_sg U50049 ( .A(n5344), .B(n28719), .X(n28718) );
  nand_x1_sg U50050 ( .A(n21833), .B(n21834), .X(n21832) );
  nand_x1_sg U50051 ( .A(n29092), .B(n29093), .X(n29082) );
  nand_x1_sg U50052 ( .A(n5382), .B(n28928), .X(n29093) );
  nand_x1_sg U50053 ( .A(n27528), .B(n27529), .X(n27527) );
  nand_x1_sg U50054 ( .A(n5325), .B(n27530), .X(n27529) );
  nand_x1_sg U50055 ( .A(n28899), .B(n28900), .X(n28898) );
  nand_x1_sg U50056 ( .A(n5364), .B(n28901), .X(n28900) );
  nand_x1_sg U50057 ( .A(n27725), .B(n27726), .X(n27718) );
  nand_x1_sg U50058 ( .A(n5307), .B(n27536), .X(n27726) );
  nand_x1_sg U50059 ( .A(n27040), .B(n27041), .X(n27039) );
  nand_x1_sg U50060 ( .A(n5155), .B(n27042), .X(n27041) );
  nand_x1_sg U50061 ( .A(n21900), .B(n21901), .X(n21899) );
  nand_x1_sg U50062 ( .A(n5136), .B(n21902), .X(n21901) );
  nand_x1_sg U50063 ( .A(n28711), .B(n28712), .X(n28710) );
  nand_x1_sg U50064 ( .A(n5345), .B(n28713), .X(n28712) );
  nand_x1_sg U50065 ( .A(n41102), .B(n21877), .X(n21874) );
  nand_x1_sg U50066 ( .A(n21880), .B(n21881), .X(n21879) );
  nor_x1_sg U50067 ( .A(n29224), .B(n29225), .X(n29075) );
  nand_x1_sg U50068 ( .A(n29077), .B(n29078), .X(n29076) );
  nand_x1_sg U50069 ( .A(n5383), .B(n29079), .X(n29078) );
  nand_x1_sg U50070 ( .A(n27722), .B(n27723), .X(n27721) );
  nand_x1_sg U50071 ( .A(n5326), .B(n27724), .X(n27723) );
  nand_x1_sg U50072 ( .A(n28893), .B(n28894), .X(n28892) );
  nand_x1_sg U50073 ( .A(n5365), .B(n28895), .X(n28894) );
  nand_x1_sg U50074 ( .A(n27902), .B(n27903), .X(n27895) );
  nand_x1_sg U50075 ( .A(n5308), .B(n27730), .X(n27903) );
  nand_x1_sg U50076 ( .A(n21947), .B(n21948), .X(n21946) );
  nand_x1_sg U50077 ( .A(n5137), .B(n21949), .X(n21948) );
  nand_x1_sg U50078 ( .A(n27034), .B(n27035), .X(n27033) );
  nand_x1_sg U50079 ( .A(n5156), .B(n27036), .X(n27035) );
  nand_x1_sg U50080 ( .A(n45564), .B(n29222), .X(n29220) );
  nand_x1_sg U50081 ( .A(n28705), .B(n28706), .X(n28704) );
  nand_x1_sg U50082 ( .A(n5346), .B(n28707), .X(n28706) );
  nand_x1_sg U50083 ( .A(n19124), .B(n21923), .X(n21920) );
  nand_x1_sg U50084 ( .A(n21926), .B(n21927), .X(n21925) );
  nand_x1_sg U50085 ( .A(n29070), .B(n29071), .X(n29069) );
  nand_x1_sg U50086 ( .A(n5384), .B(n29072), .X(n29071) );
  nand_x1_sg U50087 ( .A(n27899), .B(n27900), .X(n27898) );
  nand_x1_sg U50088 ( .A(n5327), .B(n27901), .X(n27900) );
  nand_x1_sg U50089 ( .A(n28887), .B(n28888), .X(n28886) );
  nand_x1_sg U50090 ( .A(n5366), .B(n28889), .X(n28888) );
  nand_x1_sg U50091 ( .A(n28064), .B(n28065), .X(n28057) );
  nand_x1_sg U50092 ( .A(n5309), .B(n27907), .X(n28065) );
  nand_x1_sg U50093 ( .A(n27028), .B(n27029), .X(n27027) );
  nand_x1_sg U50094 ( .A(n5157), .B(n27030), .X(n27029) );
  nand_x1_sg U50095 ( .A(n21993), .B(n21994), .X(n21992) );
  nand_x1_sg U50096 ( .A(n5138), .B(n21995), .X(n21994) );
  nand_x1_sg U50097 ( .A(n28699), .B(n28700), .X(n28698) );
  nand_x1_sg U50098 ( .A(n5347), .B(n28701), .X(n28700) );
  nand_x1_sg U50099 ( .A(n41101), .B(n21970), .X(n21967) );
  nand_x1_sg U50100 ( .A(n21973), .B(n21974), .X(n21972) );
  nand_x1_sg U50101 ( .A(n41090), .B(n21975), .X(n21974) );
  nor_x1_sg U50102 ( .A(n29212), .B(n29213), .X(n29062) );
  nand_x1_sg U50103 ( .A(n29064), .B(n29065), .X(n29063) );
  nand_x1_sg U50104 ( .A(n5385), .B(n29066), .X(n29065) );
  nand_x1_sg U50105 ( .A(n28061), .B(n28062), .X(n28060) );
  nand_x1_sg U50106 ( .A(n5328), .B(n28063), .X(n28062) );
  nand_x1_sg U50107 ( .A(n28881), .B(n28882), .X(n28880) );
  nand_x1_sg U50108 ( .A(n5367), .B(n28883), .X(n28882) );
  nand_x1_sg U50109 ( .A(n28199), .B(n28200), .X(n28192) );
  nand_x1_sg U50110 ( .A(n5310), .B(n28069), .X(n28200) );
  nand_x1_sg U50111 ( .A(n27022), .B(n27023), .X(n27021) );
  nand_x1_sg U50112 ( .A(n5158), .B(n27024), .X(n27023) );
  nand_x1_sg U50113 ( .A(n22040), .B(n22041), .X(n22039) );
  nand_x1_sg U50114 ( .A(n5139), .B(n22042), .X(n22041) );
  nand_x1_sg U50115 ( .A(n45475), .B(n29210), .X(n29208) );
  nand_x1_sg U50116 ( .A(n28693), .B(n28694), .X(n28692) );
  nand_x1_sg U50117 ( .A(n5348), .B(n28695), .X(n28694) );
  nand_x1_sg U50118 ( .A(n41102), .B(n22016), .X(n22013) );
  nand_x1_sg U50119 ( .A(n22019), .B(n22020), .X(n22018) );
  nand_x1_sg U50120 ( .A(n29057), .B(n29058), .X(n29056) );
  nand_x1_sg U50121 ( .A(n5386), .B(n29059), .X(n29058) );
  nand_x1_sg U50122 ( .A(n28196), .B(n28197), .X(n28195) );
  nand_x1_sg U50123 ( .A(n5329), .B(n28198), .X(n28197) );
  nand_x1_sg U50124 ( .A(n28875), .B(n28876), .X(n28874) );
  nand_x1_sg U50125 ( .A(n5368), .B(n28877), .X(n28876) );
  nand_x1_sg U50126 ( .A(n28328), .B(n28329), .X(n28321) );
  nand_x1_sg U50127 ( .A(n5311), .B(n28204), .X(n28329) );
  nand_x1_sg U50128 ( .A(n27016), .B(n27017), .X(n27015) );
  nand_x1_sg U50129 ( .A(n5159), .B(n27018), .X(n27017) );
  nand_x1_sg U50130 ( .A(n22086), .B(n22087), .X(n22085) );
  nand_x1_sg U50131 ( .A(n5140), .B(n22088), .X(n22087) );
  nand_x1_sg U50132 ( .A(n28687), .B(n28688), .X(n28686) );
  nand_x1_sg U50133 ( .A(n5349), .B(n28689), .X(n28688) );
  nand_x1_sg U50134 ( .A(n41103), .B(n22063), .X(n22060) );
  nand_x1_sg U50135 ( .A(n22066), .B(n22067), .X(n22065) );
  nand_x1_sg U50136 ( .A(n39260), .B(n22068), .X(n22067) );
  nor_x1_sg U50137 ( .A(n29200), .B(n29201), .X(n29049) );
  nand_x1_sg U50138 ( .A(n29051), .B(n29052), .X(n29050) );
  nand_x1_sg U50139 ( .A(n5387), .B(n29053), .X(n29052) );
  nand_x1_sg U50140 ( .A(n28325), .B(n28326), .X(n28324) );
  nand_x1_sg U50141 ( .A(n5330), .B(n28327), .X(n28326) );
  nand_x1_sg U50142 ( .A(n28869), .B(n28870), .X(n28868) );
  nand_x1_sg U50143 ( .A(n5369), .B(n28871), .X(n28870) );
  nand_x1_sg U50144 ( .A(n28432), .B(n28433), .X(n28425) );
  nand_x1_sg U50145 ( .A(n5312), .B(n28333), .X(n28433) );
  nand_x1_sg U50146 ( .A(n27010), .B(n27011), .X(n27009) );
  nand_x1_sg U50147 ( .A(n5160), .B(n27012), .X(n27011) );
  nand_x1_sg U50148 ( .A(n22134), .B(n22135), .X(n22133) );
  nand_x1_sg U50149 ( .A(n5141), .B(n22136), .X(n22135) );
  nand_x1_sg U50150 ( .A(n45385), .B(n29198), .X(n29196) );
  nand_x1_sg U50151 ( .A(n28681), .B(n28682), .X(n28680) );
  nand_x1_sg U50152 ( .A(n5350), .B(n28683), .X(n28682) );
  nand_x1_sg U50153 ( .A(n39257), .B(n22109), .X(n22106) );
  nand_x1_sg U50154 ( .A(n22112), .B(n22113), .X(n22111) );
  nand_x1_sg U50155 ( .A(n29044), .B(n29045), .X(n29043) );
  nand_x1_sg U50156 ( .A(n5388), .B(n29046), .X(n29045) );
  nand_x1_sg U50157 ( .A(n28429), .B(n28430), .X(n28428) );
  nand_x1_sg U50158 ( .A(n5331), .B(n28431), .X(n28430) );
  nand_x1_sg U50159 ( .A(n28863), .B(n28864), .X(n28862) );
  nand_x1_sg U50160 ( .A(n5370), .B(n28865), .X(n28864) );
  nand_x1_sg U50161 ( .A(n28420), .B(n28421), .X(n28419) );
  nand_x1_sg U50162 ( .A(n5313), .B(n28422), .X(n28421) );
  nand_x1_sg U50163 ( .A(n27004), .B(n27005), .X(n27003) );
  nand_x1_sg U50164 ( .A(n5161), .B(n27006), .X(n27005) );
  nand_x1_sg U50165 ( .A(n22181), .B(n22182), .X(n22180) );
  nand_x1_sg U50166 ( .A(n5142), .B(n22183), .X(n22182) );
  nand_x1_sg U50167 ( .A(n28675), .B(n28676), .X(n28674) );
  nand_x1_sg U50168 ( .A(n5351), .B(n28677), .X(n28676) );
  nand_x1_sg U50169 ( .A(n39257), .B(n22157), .X(n22154) );
  nand_x1_sg U50170 ( .A(n22160), .B(n22161), .X(n22159) );
  nor_x1_sg U50171 ( .A(n29188), .B(n29189), .X(n29036) );
  nand_x1_sg U50172 ( .A(n29038), .B(n29039), .X(n29037) );
  nand_x1_sg U50173 ( .A(n5389), .B(n29040), .X(n29039) );
  nand_x1_sg U50174 ( .A(n28514), .B(n28515), .X(n28513) );
  nand_x1_sg U50175 ( .A(n5332), .B(n28516), .X(n28515) );
  nand_x1_sg U50176 ( .A(n28857), .B(n28858), .X(n28856) );
  nand_x1_sg U50177 ( .A(n5371), .B(n28859), .X(n28858) );
  nand_x1_sg U50178 ( .A(n28414), .B(n28415), .X(n28413) );
  nand_x1_sg U50179 ( .A(n5314), .B(n28416), .X(n28415) );
  nand_x1_sg U50180 ( .A(n26998), .B(n26999), .X(n26997) );
  nand_x1_sg U50181 ( .A(n5162), .B(n27000), .X(n26999) );
  nand_x1_sg U50182 ( .A(n22229), .B(n22230), .X(n22228) );
  nand_x1_sg U50183 ( .A(n5143), .B(n22231), .X(n22230) );
  nand_x1_sg U50184 ( .A(n42085), .B(n29186), .X(n29184) );
  nand_x1_sg U50185 ( .A(n28669), .B(n28670), .X(n28668) );
  nand_x1_sg U50186 ( .A(n5352), .B(n28671), .X(n28670) );
  nand_x1_sg U50187 ( .A(n41101), .B(n22204), .X(n22201) );
  nand_x1_sg U50188 ( .A(n22207), .B(n22208), .X(n22206) );
  nand_x1_sg U50189 ( .A(n41090), .B(n22209), .X(n22208) );
  nand_x1_sg U50190 ( .A(n29031), .B(n29032), .X(n29030) );
  nand_x1_sg U50191 ( .A(n5390), .B(n29033), .X(n29032) );
  nand_x1_sg U50192 ( .A(n28508), .B(n28509), .X(n28507) );
  nand_x1_sg U50193 ( .A(n5333), .B(n28510), .X(n28509) );
  nand_x1_sg U50194 ( .A(n28851), .B(n28852), .X(n28850) );
  nand_x1_sg U50195 ( .A(n5372), .B(n28853), .X(n28852) );
  nand_x1_sg U50196 ( .A(n28408), .B(n28409), .X(n28407) );
  nand_x1_sg U50197 ( .A(n5315), .B(n28410), .X(n28409) );
  nand_x1_sg U50198 ( .A(n26992), .B(n26993), .X(n26991) );
  nand_x1_sg U50199 ( .A(n5163), .B(n26994), .X(n26993) );
  nand_x1_sg U50200 ( .A(n22276), .B(n22277), .X(n22275) );
  nand_x1_sg U50201 ( .A(n5144), .B(n22278), .X(n22277) );
  nand_x1_sg U50202 ( .A(n28663), .B(n28664), .X(n28662) );
  nand_x1_sg U50203 ( .A(n5353), .B(n28665), .X(n28664) );
  nand_x1_sg U50204 ( .A(n38934), .B(n22252), .X(n22249) );
  nand_x1_sg U50205 ( .A(n22255), .B(n22256), .X(n22254) );
  nand_x1_sg U50206 ( .A(n38928), .B(n22257), .X(n22256) );
  nor_x1_sg U50207 ( .A(n29176), .B(n29177), .X(n29023) );
  nand_x1_sg U50208 ( .A(n29025), .B(n29026), .X(n29024) );
  nand_x1_sg U50209 ( .A(n5391), .B(n29027), .X(n29026) );
  nand_x1_sg U50210 ( .A(n28502), .B(n28503), .X(n28501) );
  nand_x1_sg U50211 ( .A(n5334), .B(n28504), .X(n28503) );
  nand_x1_sg U50212 ( .A(n28845), .B(n28846), .X(n28844) );
  nand_x1_sg U50213 ( .A(n5373), .B(n28847), .X(n28846) );
  nand_x1_sg U50214 ( .A(n28402), .B(n28403), .X(n28401) );
  nand_x1_sg U50215 ( .A(n5316), .B(n28404), .X(n28403) );
  nand_x1_sg U50216 ( .A(n26986), .B(n26987), .X(n26985) );
  nand_x1_sg U50217 ( .A(n5164), .B(n26988), .X(n26987) );
  nand_x1_sg U50218 ( .A(n22324), .B(n22325), .X(n22323) );
  nand_x1_sg U50219 ( .A(n5145), .B(n22326), .X(n22325) );
  nand_x1_sg U50220 ( .A(n45204), .B(n29174), .X(n29172) );
  nand_x1_sg U50221 ( .A(n28657), .B(n28658), .X(n28656) );
  nand_x1_sg U50222 ( .A(n5354), .B(n28659), .X(n28658) );
  nand_x1_sg U50223 ( .A(n19124), .B(n22299), .X(n22296) );
  nand_x1_sg U50224 ( .A(n22302), .B(n22303), .X(n22301) );
  nand_x1_sg U50225 ( .A(n29018), .B(n29019), .X(n29017) );
  nand_x1_sg U50226 ( .A(n5392), .B(n29020), .X(n29019) );
  nand_x1_sg U50227 ( .A(n28496), .B(n28497), .X(n28495) );
  nand_x1_sg U50228 ( .A(n5335), .B(n28498), .X(n28497) );
  nand_x1_sg U50229 ( .A(n28839), .B(n28840), .X(n28838) );
  nand_x1_sg U50230 ( .A(n5374), .B(n28841), .X(n28840) );
  nand_x1_sg U50231 ( .A(n28396), .B(n28397), .X(n28395) );
  nand_x1_sg U50232 ( .A(n5317), .B(n28398), .X(n28397) );
  nand_x1_sg U50233 ( .A(n26980), .B(n26981), .X(n26979) );
  nand_x1_sg U50234 ( .A(n5165), .B(n26982), .X(n26981) );
  nand_x1_sg U50235 ( .A(n22371), .B(n22372), .X(n22370) );
  nand_x1_sg U50236 ( .A(n5146), .B(n22373), .X(n22372) );
  nand_x1_sg U50237 ( .A(n28651), .B(n28652), .X(n28650) );
  nand_x1_sg U50238 ( .A(n5355), .B(n28653), .X(n28652) );
  nand_x1_sg U50239 ( .A(n41102), .B(n22347), .X(n22344) );
  nand_x1_sg U50240 ( .A(n22350), .B(n22351), .X(n22349) );
  nand_x1_sg U50241 ( .A(n41091), .B(n22352), .X(n22351) );
  nor_x1_sg U50242 ( .A(n29164), .B(n29165), .X(n29010) );
  nand_x1_sg U50243 ( .A(n29012), .B(n29013), .X(n29011) );
  nand_x1_sg U50244 ( .A(n5393), .B(n29014), .X(n29013) );
  nand_x1_sg U50245 ( .A(n28490), .B(n28491), .X(n28489) );
  nand_x1_sg U50246 ( .A(n5336), .B(n28492), .X(n28491) );
  nand_x1_sg U50247 ( .A(n28833), .B(n28834), .X(n28832) );
  nand_x1_sg U50248 ( .A(n5375), .B(n28835), .X(n28834) );
  nand_x1_sg U50249 ( .A(n28390), .B(n28391), .X(n28389) );
  nand_x1_sg U50250 ( .A(n5318), .B(n28392), .X(n28391) );
  nand_x1_sg U50251 ( .A(n26974), .B(n26975), .X(n26973) );
  nand_x1_sg U50252 ( .A(n5166), .B(n26976), .X(n26975) );
  nand_x1_sg U50253 ( .A(n22419), .B(n22420), .X(n22418) );
  nand_x1_sg U50254 ( .A(n5147), .B(n22421), .X(n22420) );
  nand_x1_sg U50255 ( .A(n45113), .B(n29162), .X(n29160) );
  nand_x1_sg U50256 ( .A(n28645), .B(n28646), .X(n28644) );
  nand_x1_sg U50257 ( .A(n5356), .B(n28647), .X(n28646) );
  nand_x1_sg U50258 ( .A(n41103), .B(n22394), .X(n22391) );
  nand_x1_sg U50259 ( .A(n22397), .B(n22398), .X(n22396) );
  nand_x1_sg U50260 ( .A(n41091), .B(n22399), .X(n22398) );
  nand_x1_sg U50261 ( .A(n29005), .B(n29006), .X(n29004) );
  nand_x1_sg U50262 ( .A(n5394), .B(n29007), .X(n29006) );
  nand_x1_sg U50263 ( .A(n28484), .B(n28485), .X(n28483) );
  nand_x1_sg U50264 ( .A(n5337), .B(n28486), .X(n28485) );
  nand_x1_sg U50265 ( .A(n28384), .B(n28385), .X(n28383) );
  nand_x1_sg U50266 ( .A(n5319), .B(n28386), .X(n28385) );
  nand_x1_sg U50267 ( .A(n28827), .B(n28828), .X(n28826) );
  nand_x1_sg U50268 ( .A(n5376), .B(n28829), .X(n28828) );
  nand_x1_sg U50269 ( .A(n26968), .B(n26969), .X(n26967) );
  nand_x1_sg U50270 ( .A(n5167), .B(n26970), .X(n26969) );
  nand_x1_sg U50271 ( .A(n22465), .B(n22466), .X(n22464) );
  nand_x1_sg U50272 ( .A(n5148), .B(n22467), .X(n22466) );
  nand_x1_sg U50273 ( .A(n28639), .B(n28640), .X(n28638) );
  nand_x1_sg U50274 ( .A(n5357), .B(n28641), .X(n28640) );
  nand_x1_sg U50275 ( .A(n22444), .B(n22445), .X(n22443) );
  nand_x1_sg U50276 ( .A(n38928), .B(n22446), .X(n22445) );
  nand_x1_sg U50277 ( .A(n28478), .B(n28479), .X(n28477) );
  nand_x1_sg U50278 ( .A(n5338), .B(n28480), .X(n28479) );
  nor_x1_sg U50279 ( .A(n29152), .B(n29153), .X(n28997) );
  nand_x1_sg U50280 ( .A(n28999), .B(n29000), .X(n28998) );
  nand_x1_sg U50281 ( .A(n5395), .B(n29001), .X(n29000) );
  nand_x1_sg U50282 ( .A(n28378), .B(n28379), .X(n28377) );
  nand_x1_sg U50283 ( .A(n28821), .B(n28822), .X(n28820) );
  nand_x1_sg U50284 ( .A(n26962), .B(n26963), .X(n26961) );
  nand_x1_sg U50285 ( .A(n22511), .B(n22512), .X(n22510) );
  nand_x1_sg U50286 ( .A(n28633), .B(n28634), .X(n28632) );
  nand_x1_sg U50287 ( .A(n45023), .B(n29150), .X(n29148) );
  nand_x1_sg U50288 ( .A(n22490), .B(n22491), .X(n22489) );
  nand_x1_sg U50289 ( .A(n28472), .B(n28473), .X(n28471) );
  nand_x1_sg U50290 ( .A(n28992), .B(n28993), .X(n28991) );
  inv_x1_sg U50291 ( .A(n28812), .X(n44983) );
  inv_x1_sg U50292 ( .A(n28369), .X(n44992) );
  nand_x1_sg U50293 ( .A(n45018), .B(n22550), .X(n22548) );
  inv_x1_sg U50294 ( .A(n29142), .X(n44977) );
  inv_x1_sg U50295 ( .A(n28624), .X(n44986) );
  nand_x1_sg U50296 ( .A(n22533), .B(n22534), .X(n22532) );
  inv_x1_sg U50297 ( .A(n28983), .X(n44980) );
  inv_x1_sg U50298 ( .A(n28464), .X(n44989) );
  nand_x1_sg U50299 ( .A(n22572), .B(n22573), .X(n22571) );
  nor_x1_sg U50300 ( .A(n22831), .B(n22832), .X(n22824) );
  inv_x1_sg U50301 ( .A(n22836), .X(n46852) );
  inv_x1_sg U50302 ( .A(n22827), .X(n46857) );
  nor_x1_sg U50303 ( .A(n46846), .B(n22822), .X(n22816) );
  inv_x1_sg U50304 ( .A(n22825), .X(n46846) );
  inv_x1_sg U50305 ( .A(n22786), .X(n46891) );
  nand_x1_sg U50306 ( .A(n22790), .B(n22791), .X(n22786) );
  inv_x1_sg U50307 ( .A(n22732), .X(n47056) );
  nand_x1_sg U50308 ( .A(n22734), .B(n22735), .X(n22732) );
  inv_x1_sg U50309 ( .A(n22716), .X(n47129) );
  nor_x1_sg U50310 ( .A(n22711), .B(n22712), .X(n22709) );
  nor_x1_sg U50311 ( .A(n22722), .B(n22723), .X(n22718) );
  nor_x1_sg U50312 ( .A(n23108), .B(n47137), .X(n23102) );
  inv_x1_sg U50313 ( .A(n23109), .X(n47137) );
  inv_x1_sg U50314 ( .A(n23113), .X(n47145) );
  inv_x1_sg U50315 ( .A(n23063), .X(n47184) );
  nand_x1_sg U50316 ( .A(n23067), .B(n23068), .X(n23063) );
  inv_x1_sg U50317 ( .A(n23009), .X(n47342) );
  nand_x1_sg U50318 ( .A(n23011), .B(n23012), .X(n23009) );
  nor_x1_sg U50319 ( .A(n23388), .B(n47422), .X(n23382) );
  inv_x1_sg U50320 ( .A(n23389), .X(n47422) );
  inv_x1_sg U50321 ( .A(n23393), .X(n47430) );
  inv_x1_sg U50322 ( .A(n23343), .X(n47469) );
  nand_x1_sg U50323 ( .A(n23347), .B(n23348), .X(n23343) );
  inv_x1_sg U50324 ( .A(n23289), .X(n47627) );
  nand_x1_sg U50325 ( .A(n23291), .B(n23292), .X(n23289) );
  nor_x1_sg U50326 ( .A(n23667), .B(n47707), .X(n23661) );
  inv_x1_sg U50327 ( .A(n23668), .X(n47707) );
  inv_x1_sg U50328 ( .A(n23672), .X(n47715) );
  inv_x1_sg U50329 ( .A(n23622), .X(n47754) );
  nand_x1_sg U50330 ( .A(n23626), .B(n23627), .X(n23622) );
  inv_x1_sg U50331 ( .A(n23568), .X(n47912) );
  nand_x1_sg U50332 ( .A(n23570), .B(n23571), .X(n23568) );
  nor_x1_sg U50333 ( .A(n23946), .B(n47992), .X(n23940) );
  inv_x1_sg U50334 ( .A(n23947), .X(n47992) );
  inv_x1_sg U50335 ( .A(n23951), .X(n48000) );
  inv_x1_sg U50336 ( .A(n23901), .X(n48039) );
  nand_x1_sg U50337 ( .A(n23905), .B(n23906), .X(n23901) );
  inv_x1_sg U50338 ( .A(n23847), .X(n48197) );
  nand_x1_sg U50339 ( .A(n23849), .B(n23850), .X(n23847) );
  nor_x1_sg U50340 ( .A(n24225), .B(n48277), .X(n24219) );
  inv_x1_sg U50341 ( .A(n24226), .X(n48277) );
  inv_x1_sg U50342 ( .A(n24230), .X(n48285) );
  inv_x1_sg U50343 ( .A(n24180), .X(n48324) );
  nand_x1_sg U50344 ( .A(n24184), .B(n24185), .X(n24180) );
  inv_x1_sg U50345 ( .A(n24161), .X(n48373) );
  nand_x1_sg U50346 ( .A(n24163), .B(n24164), .X(n24161) );
  inv_x1_sg U50347 ( .A(n24126), .X(n48482) );
  nand_x1_sg U50348 ( .A(n24128), .B(n24129), .X(n24126) );
  nand_x1_sg U50349 ( .A(n39081), .B(n29270), .X(n24101) );
  nor_x1_sg U50350 ( .A(n24504), .B(n48562), .X(n24498) );
  inv_x1_sg U50351 ( .A(n24505), .X(n48562) );
  inv_x1_sg U50352 ( .A(n24509), .X(n48570) );
  inv_x1_sg U50353 ( .A(n24459), .X(n48609) );
  nand_x1_sg U50354 ( .A(n24463), .B(n24464), .X(n24459) );
  inv_x1_sg U50355 ( .A(n24405), .X(n48767) );
  nand_x1_sg U50356 ( .A(n24407), .B(n24408), .X(n24405) );
  nor_x1_sg U50357 ( .A(n24782), .B(n48847), .X(n24776) );
  inv_x1_sg U50358 ( .A(n24783), .X(n48847) );
  inv_x1_sg U50359 ( .A(n24787), .X(n48855) );
  inv_x1_sg U50360 ( .A(n24737), .X(n48895) );
  nand_x1_sg U50361 ( .A(n24741), .B(n24742), .X(n24737) );
  inv_x1_sg U50362 ( .A(n24683), .X(n49053) );
  nand_x1_sg U50363 ( .A(n24685), .B(n24686), .X(n24683) );
  nor_x1_sg U50364 ( .A(n25061), .B(n49134), .X(n25055) );
  inv_x1_sg U50365 ( .A(n25062), .X(n49134) );
  inv_x1_sg U50366 ( .A(n25066), .X(n49142) );
  inv_x1_sg U50367 ( .A(n25016), .X(n49182) );
  nand_x1_sg U50368 ( .A(n25020), .B(n25021), .X(n25016) );
  inv_x1_sg U50369 ( .A(n24962), .X(n49340) );
  nand_x1_sg U50370 ( .A(n24964), .B(n24965), .X(n24962) );
  nor_x1_sg U50371 ( .A(n25340), .B(n49420), .X(n25334) );
  inv_x1_sg U50372 ( .A(n25341), .X(n49420) );
  inv_x1_sg U50373 ( .A(n25345), .X(n49428) );
  inv_x1_sg U50374 ( .A(n25295), .X(n49468) );
  nand_x1_sg U50375 ( .A(n25299), .B(n25300), .X(n25295) );
  inv_x1_sg U50376 ( .A(n25241), .X(n49626) );
  nand_x1_sg U50377 ( .A(n25243), .B(n25244), .X(n25241) );
  nor_x1_sg U50378 ( .A(n25619), .B(n49706), .X(n25613) );
  inv_x1_sg U50379 ( .A(n25620), .X(n49706) );
  inv_x1_sg U50380 ( .A(n25624), .X(n49714) );
  inv_x1_sg U50381 ( .A(n25574), .X(n49753) );
  nand_x1_sg U50382 ( .A(n25578), .B(n25579), .X(n25574) );
  inv_x1_sg U50383 ( .A(n25520), .X(n49912) );
  nand_x1_sg U50384 ( .A(n25522), .B(n25523), .X(n25520) );
  nand_x1_sg U50385 ( .A(n51138), .B(n26778), .X(n25495) );
  nor_x1_sg U50386 ( .A(n25896), .B(n49992), .X(n25890) );
  inv_x1_sg U50387 ( .A(n25897), .X(n49992) );
  inv_x1_sg U50388 ( .A(n25901), .X(n50000) );
  inv_x1_sg U50389 ( .A(n25851), .X(n50040) );
  nand_x1_sg U50390 ( .A(n25855), .B(n25856), .X(n25851) );
  inv_x1_sg U50391 ( .A(n25797), .X(n50198) );
  nand_x1_sg U50392 ( .A(n25799), .B(n25800), .X(n25797) );
  nand_x1_sg U50393 ( .A(n50280), .B(n26121), .X(n26119) );
  nand_x1_sg U50394 ( .A(n26103), .B(n26104), .X(n26101) );
  inv_x1_sg U50395 ( .A(n26084), .X(n50336) );
  nand_x1_sg U50396 ( .A(n26092), .B(n26158), .X(n26084) );
  nor_x1_sg U50397 ( .A(n26036), .B(n26037), .X(n26035) );
  nor_x1_sg U50398 ( .A(n26456), .B(n50567), .X(n26450) );
  inv_x1_sg U50399 ( .A(n26457), .X(n50567) );
  inv_x1_sg U50400 ( .A(n26461), .X(n50575) );
  inv_x1_sg U50401 ( .A(n26411), .X(n50614) );
  nand_x1_sg U50402 ( .A(n26415), .B(n26416), .X(n26411) );
  inv_x1_sg U50403 ( .A(n26357), .X(n50772) );
  nand_x1_sg U50404 ( .A(n26359), .B(n26360), .X(n26357) );
  nor_x1_sg U50405 ( .A(n26734), .B(n50853), .X(n26728) );
  inv_x1_sg U50406 ( .A(n26735), .X(n50853) );
  inv_x1_sg U50407 ( .A(n26739), .X(n50861) );
  inv_x1_sg U50408 ( .A(n26689), .X(n50901) );
  nand_x1_sg U50409 ( .A(n26693), .B(n26694), .X(n26689) );
  inv_x1_sg U50410 ( .A(n26635), .X(n51059) );
  nand_x1_sg U50411 ( .A(n26637), .B(n26638), .X(n26635) );
  nand_x1_sg U50412 ( .A(n19127), .B(n19128), .X(n19111) );
  nand_x1_sg U50413 ( .A(n19113), .B(n19114), .X(n19112) );
  nand_x1_sg U50414 ( .A(n20561), .B(n20562), .X(n20560) );
  nand_x1_sg U50415 ( .A(n20570), .B(n20571), .X(n20559) );
  nand_x1_sg U50416 ( .A(n5970), .B(n5971), .X(n5958) );
  nand_x1_sg U50417 ( .A(n5960), .B(n5961), .X(n5959) );
  nand_x1_sg U50418 ( .A(n5992), .B(n5993), .X(n5991) );
  nand_x1_sg U50419 ( .A(n5999), .B(n6000), .X(n5990) );
  nand_x1_sg U50420 ( .A(n6025), .B(n6026), .X(n6013) );
  nand_x1_sg U50421 ( .A(n6015), .B(n6016), .X(n6014) );
  nand_x1_sg U50422 ( .A(n6041), .B(n6042), .X(n6040) );
  nand_x1_sg U50423 ( .A(n6047), .B(n6048), .X(n6039) );
  nand_x1_sg U50424 ( .A(n6073), .B(n6074), .X(n6062) );
  nand_x1_sg U50425 ( .A(n6064), .B(n6065), .X(n6063) );
  nand_x1_sg U50426 ( .A(n6091), .B(n6092), .X(n6090) );
  nand_x1_sg U50427 ( .A(n6097), .B(n6098), .X(n6089) );
  nand_x1_sg U50428 ( .A(n6120), .B(n6121), .X(n6110) );
  nand_x1_sg U50429 ( .A(n6112), .B(n6113), .X(n6111) );
  nand_x1_sg U50430 ( .A(n6137), .B(n6138), .X(n6136) );
  nand_x1_sg U50431 ( .A(n6143), .B(n6144), .X(n6135) );
  nand_x1_sg U50432 ( .A(n6165), .B(n6166), .X(n6155) );
  nand_x1_sg U50433 ( .A(n6157), .B(n6158), .X(n6156) );
  nand_x1_sg U50434 ( .A(n6182), .B(n6183), .X(n6181) );
  nand_x1_sg U50435 ( .A(n6189), .B(n6190), .X(n6180) );
  nand_x1_sg U50436 ( .A(n6212), .B(n6213), .X(n6201) );
  nand_x1_sg U50437 ( .A(n6203), .B(n6204), .X(n6202) );
  nand_x1_sg U50438 ( .A(n6229), .B(n6230), .X(n6228) );
  nand_x1_sg U50439 ( .A(n6235), .B(n6236), .X(n6227) );
  nand_x1_sg U50440 ( .A(n6258), .B(n6259), .X(n6248) );
  nand_x1_sg U50441 ( .A(n6250), .B(n6251), .X(n6249) );
  nand_x1_sg U50442 ( .A(n6273), .B(n6274), .X(n6272) );
  nand_x1_sg U50443 ( .A(n6280), .B(n6281), .X(n6271) );
  nand_x1_sg U50444 ( .A(n6303), .B(n6304), .X(n6293) );
  nand_x1_sg U50445 ( .A(n6295), .B(n6296), .X(n6294) );
  nand_x1_sg U50446 ( .A(n6318), .B(n6319), .X(n6317) );
  nand_x1_sg U50447 ( .A(n6324), .B(n6325), .X(n6316) );
  nand_x1_sg U50448 ( .A(n6347), .B(n6348), .X(n6337) );
  nand_x1_sg U50449 ( .A(n6339), .B(n6340), .X(n6338) );
  nand_x1_sg U50450 ( .A(n6362), .B(n6363), .X(n6361) );
  nand_x1_sg U50451 ( .A(n6369), .B(n6370), .X(n6360) );
  nand_x1_sg U50452 ( .A(n6392), .B(n6393), .X(n6382) );
  nand_x1_sg U50453 ( .A(n6384), .B(n6385), .X(n6383) );
  nand_x1_sg U50454 ( .A(n6407), .B(n6408), .X(n6406) );
  nand_x1_sg U50455 ( .A(n6413), .B(n6414), .X(n6405) );
  nand_x1_sg U50456 ( .A(n6436), .B(n6437), .X(n6426) );
  nand_x1_sg U50457 ( .A(n6428), .B(n6429), .X(n6427) );
  nand_x1_sg U50458 ( .A(n6451), .B(n6452), .X(n6450) );
  nand_x1_sg U50459 ( .A(n6458), .B(n6459), .X(n6449) );
  nand_x1_sg U50460 ( .A(n6481), .B(n6482), .X(n6471) );
  nand_x1_sg U50461 ( .A(n6473), .B(n6474), .X(n6472) );
  nand_x1_sg U50462 ( .A(n6496), .B(n6497), .X(n6495) );
  nand_x1_sg U50463 ( .A(n6502), .B(n6503), .X(n6494) );
  nand_x1_sg U50464 ( .A(n6525), .B(n6526), .X(n6515) );
  nand_x1_sg U50465 ( .A(n6517), .B(n6518), .X(n6516) );
  nand_x1_sg U50466 ( .A(n6540), .B(n6541), .X(n6539) );
  nand_x1_sg U50467 ( .A(n6547), .B(n6548), .X(n6538) );
  nand_x1_sg U50468 ( .A(n6570), .B(n6571), .X(n6560) );
  nand_x1_sg U50469 ( .A(n6562), .B(n6563), .X(n6561) );
  nand_x1_sg U50470 ( .A(n6585), .B(n6586), .X(n6584) );
  nand_x1_sg U50471 ( .A(n6591), .B(n6592), .X(n6583) );
  nand_x1_sg U50472 ( .A(n6614), .B(n6615), .X(n6604) );
  nand_x1_sg U50473 ( .A(n6606), .B(n6607), .X(n6605) );
  nand_x1_sg U50474 ( .A(n6629), .B(n6630), .X(n6628) );
  nand_x1_sg U50475 ( .A(n6636), .B(n6637), .X(n6627) );
  nand_x1_sg U50476 ( .A(n6660), .B(n6661), .X(n6649) );
  nand_x1_sg U50477 ( .A(n6651), .B(n6652), .X(n6650) );
  nand_x1_sg U50478 ( .A(n6677), .B(n6678), .X(n6676) );
  nand_x1_sg U50479 ( .A(n6683), .B(n6684), .X(n6675) );
  nand_x1_sg U50480 ( .A(n6705), .B(n6706), .X(n6697) );
  nand_x1_sg U50481 ( .A(n6699), .B(n6700), .X(n6698) );
  nand_x1_sg U50482 ( .A(n6721), .B(n6722), .X(n6720) );
  nand_x1_sg U50483 ( .A(n6726), .B(n6727), .X(n6719) );
  nand_x1_sg U50484 ( .A(n6749), .B(n6750), .X(n6737) );
  nand_x1_sg U50485 ( .A(n6739), .B(n6740), .X(n6738) );
  nand_x1_sg U50486 ( .A(n6767), .B(n6768), .X(n6766) );
  nand_x1_sg U50487 ( .A(n6773), .B(n6774), .X(n6765) );
  nand_x1_sg U50488 ( .A(n6798), .B(n6799), .X(n6788) );
  nand_x1_sg U50489 ( .A(n6790), .B(n6791), .X(n6789) );
  nand_x1_sg U50490 ( .A(n6810), .B(n6811), .X(n6809) );
  nand_x1_sg U50491 ( .A(n6814), .B(n6815), .X(n6808) );
  nor_x1_sg U50492 ( .A(n7077), .B(n7078), .X(n6840) );
  nand_x1_sg U50493 ( .A(n7068), .B(n7069), .X(n6852) );
  nand_x1_sg U50494 ( .A(n7109), .B(n7110), .X(n6866) );
  nand_x1_sg U50495 ( .A(n6866), .B(n6865), .X(n6863) );
  nand_x1_sg U50496 ( .A(n7063), .B(n6863), .X(n6871) );
  nand_x1_sg U50497 ( .A(n7171), .B(n46951), .X(n6884) );
  nand_x1_sg U50498 ( .A(n7060), .B(n7061), .X(n6883) );
  nand_x1_sg U50499 ( .A(n46931), .B(n6876), .X(n7061) );
  inv_x1_sg U50500 ( .A(n6964), .X(n47125) );
  nand_x1_sg U50501 ( .A(n6933), .B(n47102), .X(n6931) );
  nand_x1_sg U50502 ( .A(n6936), .B(n6935), .X(n6933) );
  nor_x1_sg U50503 ( .A(n7895), .B(n7896), .X(n7657) );
  nand_x1_sg U50504 ( .A(n7886), .B(n7887), .X(n7669) );
  nand_x1_sg U50505 ( .A(n7927), .B(n7928), .X(n7683) );
  nand_x1_sg U50506 ( .A(n7683), .B(n7682), .X(n7680) );
  nand_x1_sg U50507 ( .A(n7881), .B(n7680), .X(n7688) );
  nand_x1_sg U50508 ( .A(n7990), .B(n47242), .X(n7701) );
  nand_x1_sg U50509 ( .A(n7878), .B(n7879), .X(n7700) );
  nand_x1_sg U50510 ( .A(n47223), .B(n7693), .X(n7879) );
  inv_x1_sg U50511 ( .A(n7781), .X(n47411) );
  nand_x1_sg U50512 ( .A(n7750), .B(n47388), .X(n7748) );
  nand_x1_sg U50513 ( .A(n7753), .B(n7752), .X(n7750) );
  nand_x1_sg U50514 ( .A(n23407), .B(n23408), .X(n23406) );
  nor_x1_sg U50515 ( .A(n8713), .B(n8714), .X(n8475) );
  nand_x1_sg U50516 ( .A(n8704), .B(n8705), .X(n8487) );
  nand_x1_sg U50517 ( .A(n8745), .B(n8746), .X(n8501) );
  nand_x1_sg U50518 ( .A(n8501), .B(n8500), .X(n8498) );
  nand_x1_sg U50519 ( .A(n8699), .B(n8498), .X(n8506) );
  nand_x1_sg U50520 ( .A(n8808), .B(n47527), .X(n8519) );
  nand_x1_sg U50521 ( .A(n8696), .B(n8697), .X(n8518) );
  nand_x1_sg U50522 ( .A(n47508), .B(n8511), .X(n8697) );
  inv_x1_sg U50523 ( .A(n8599), .X(n47696) );
  nand_x1_sg U50524 ( .A(n8568), .B(n47673), .X(n8566) );
  nand_x1_sg U50525 ( .A(n8571), .B(n8570), .X(n8568) );
  nand_x1_sg U50526 ( .A(n23686), .B(n23687), .X(n23685) );
  nor_x1_sg U50527 ( .A(n9533), .B(n9534), .X(n9295) );
  nand_x1_sg U50528 ( .A(n9524), .B(n9525), .X(n9307) );
  nand_x1_sg U50529 ( .A(n9565), .B(n9566), .X(n9321) );
  nand_x1_sg U50530 ( .A(n9321), .B(n9320), .X(n9318) );
  nand_x1_sg U50531 ( .A(n9519), .B(n9318), .X(n9326) );
  nand_x1_sg U50532 ( .A(n9628), .B(n47812), .X(n9339) );
  nand_x1_sg U50533 ( .A(n9516), .B(n9517), .X(n9338) );
  nand_x1_sg U50534 ( .A(n47793), .B(n9331), .X(n9517) );
  inv_x1_sg U50535 ( .A(n9419), .X(n47981) );
  nand_x1_sg U50536 ( .A(n9388), .B(n47958), .X(n9386) );
  nand_x1_sg U50537 ( .A(n9391), .B(n9390), .X(n9388) );
  nand_x1_sg U50538 ( .A(n23965), .B(n23966), .X(n23964) );
  nor_x1_sg U50539 ( .A(n10352), .B(n10353), .X(n10114) );
  nand_x1_sg U50540 ( .A(n10343), .B(n10344), .X(n10126) );
  nand_x1_sg U50541 ( .A(n10384), .B(n10385), .X(n10140) );
  nand_x1_sg U50542 ( .A(n10140), .B(n10139), .X(n10137) );
  nand_x1_sg U50543 ( .A(n10338), .B(n10137), .X(n10145) );
  nand_x1_sg U50544 ( .A(n10447), .B(n48097), .X(n10158) );
  nand_x1_sg U50545 ( .A(n10335), .B(n10336), .X(n10157) );
  nand_x1_sg U50546 ( .A(n48078), .B(n10150), .X(n10336) );
  inv_x1_sg U50547 ( .A(n10238), .X(n48266) );
  nand_x1_sg U50548 ( .A(n10207), .B(n48243), .X(n10205) );
  nand_x1_sg U50549 ( .A(n10210), .B(n10209), .X(n10207) );
  nand_x1_sg U50550 ( .A(n24244), .B(n24245), .X(n24243) );
  nor_x1_sg U50551 ( .A(n11171), .B(n11172), .X(n10933) );
  nand_x1_sg U50552 ( .A(n11162), .B(n11163), .X(n10945) );
  nand_x1_sg U50553 ( .A(n11203), .B(n11204), .X(n10959) );
  nand_x1_sg U50554 ( .A(n10959), .B(n10958), .X(n10956) );
  nand_x1_sg U50555 ( .A(n11157), .B(n10956), .X(n10964) );
  nand_x1_sg U50556 ( .A(n11266), .B(n48382), .X(n10977) );
  nand_x1_sg U50557 ( .A(n11154), .B(n11155), .X(n10976) );
  nand_x1_sg U50558 ( .A(n48363), .B(n10969), .X(n11155) );
  inv_x1_sg U50559 ( .A(n11057), .X(n48551) );
  nand_x1_sg U50560 ( .A(n11026), .B(n48528), .X(n11024) );
  nand_x1_sg U50561 ( .A(n11029), .B(n11028), .X(n11026) );
  nand_x1_sg U50562 ( .A(n24523), .B(n24524), .X(n24522) );
  nor_x1_sg U50563 ( .A(n11990), .B(n11991), .X(n11752) );
  nand_x1_sg U50564 ( .A(n11981), .B(n11982), .X(n11764) );
  nand_x1_sg U50565 ( .A(n12022), .B(n12023), .X(n11778) );
  nand_x1_sg U50566 ( .A(n11778), .B(n11777), .X(n11775) );
  nand_x1_sg U50567 ( .A(n11976), .B(n11775), .X(n11783) );
  nand_x1_sg U50568 ( .A(n12085), .B(n48667), .X(n11796) );
  nand_x1_sg U50569 ( .A(n11973), .B(n11974), .X(n11795) );
  nand_x1_sg U50570 ( .A(n48648), .B(n11788), .X(n11974) );
  inv_x1_sg U50571 ( .A(n11876), .X(n48836) );
  nand_x1_sg U50572 ( .A(n11845), .B(n48813), .X(n11843) );
  nand_x1_sg U50573 ( .A(n11848), .B(n11847), .X(n11845) );
  nand_x1_sg U50574 ( .A(n24801), .B(n24802), .X(n24800) );
  nor_x1_sg U50575 ( .A(n12809), .B(n12810), .X(n12571) );
  nand_x1_sg U50576 ( .A(n12800), .B(n12801), .X(n12583) );
  nand_x1_sg U50577 ( .A(n12841), .B(n12842), .X(n12597) );
  nand_x1_sg U50578 ( .A(n12597), .B(n12596), .X(n12594) );
  nand_x1_sg U50579 ( .A(n12795), .B(n12594), .X(n12602) );
  nand_x1_sg U50580 ( .A(n12904), .B(n48953), .X(n12615) );
  nand_x1_sg U50581 ( .A(n12792), .B(n12793), .X(n12614) );
  nand_x1_sg U50582 ( .A(n48934), .B(n12607), .X(n12793) );
  inv_x1_sg U50583 ( .A(n12695), .X(n49123) );
  nand_x1_sg U50584 ( .A(n12664), .B(n49100), .X(n12662) );
  nand_x1_sg U50585 ( .A(n12667), .B(n12666), .X(n12664) );
  nand_x1_sg U50586 ( .A(n25080), .B(n25081), .X(n25079) );
  nor_x1_sg U50587 ( .A(n13628), .B(n13629), .X(n13390) );
  nand_x1_sg U50588 ( .A(n13619), .B(n13620), .X(n13402) );
  nand_x1_sg U50589 ( .A(n13660), .B(n13661), .X(n13416) );
  nand_x1_sg U50590 ( .A(n13416), .B(n13415), .X(n13413) );
  nand_x1_sg U50591 ( .A(n13614), .B(n13413), .X(n13421) );
  nand_x1_sg U50592 ( .A(n13723), .B(n49240), .X(n13434) );
  nand_x1_sg U50593 ( .A(n13611), .B(n13612), .X(n13433) );
  nand_x1_sg U50594 ( .A(n49221), .B(n13426), .X(n13612) );
  inv_x1_sg U50595 ( .A(n13514), .X(n49409) );
  nand_x1_sg U50596 ( .A(n13483), .B(n49386), .X(n13481) );
  nand_x1_sg U50597 ( .A(n13486), .B(n13485), .X(n13483) );
  nand_x1_sg U50598 ( .A(n25359), .B(n25360), .X(n25358) );
  nor_x1_sg U50599 ( .A(n14447), .B(n14448), .X(n14209) );
  nand_x1_sg U50600 ( .A(n14438), .B(n14439), .X(n14221) );
  nand_x1_sg U50601 ( .A(n14479), .B(n14480), .X(n14235) );
  nand_x1_sg U50602 ( .A(n14235), .B(n14234), .X(n14232) );
  nand_x1_sg U50603 ( .A(n14433), .B(n14232), .X(n14240) );
  nand_x1_sg U50604 ( .A(n14542), .B(n49526), .X(n14253) );
  nand_x1_sg U50605 ( .A(n14430), .B(n14431), .X(n14252) );
  nand_x1_sg U50606 ( .A(n49507), .B(n14245), .X(n14431) );
  inv_x1_sg U50607 ( .A(n14333), .X(n49695) );
  nand_x1_sg U50608 ( .A(n14302), .B(n49672), .X(n14300) );
  nand_x1_sg U50609 ( .A(n14305), .B(n14304), .X(n14302) );
  nand_x1_sg U50610 ( .A(n25638), .B(n25639), .X(n25637) );
  nor_x1_sg U50611 ( .A(n15266), .B(n15267), .X(n15028) );
  nand_x1_sg U50612 ( .A(n15257), .B(n15258), .X(n15040) );
  nand_x1_sg U50613 ( .A(n15298), .B(n15299), .X(n15054) );
  nand_x1_sg U50614 ( .A(n15054), .B(n15053), .X(n15051) );
  nand_x1_sg U50615 ( .A(n15252), .B(n15051), .X(n15059) );
  nand_x1_sg U50616 ( .A(n15361), .B(n49812), .X(n15072) );
  nand_x1_sg U50617 ( .A(n15249), .B(n15250), .X(n15071) );
  nand_x1_sg U50618 ( .A(n49793), .B(n15064), .X(n15250) );
  inv_x1_sg U50619 ( .A(n15152), .X(n49981) );
  nand_x1_sg U50620 ( .A(n15121), .B(n49958), .X(n15119) );
  nand_x1_sg U50621 ( .A(n15124), .B(n15123), .X(n15121) );
  nand_x1_sg U50622 ( .A(n25915), .B(n25916), .X(n25914) );
  nor_x1_sg U50623 ( .A(n16085), .B(n16086), .X(n15847) );
  nand_x1_sg U50624 ( .A(n16076), .B(n16077), .X(n15859) );
  nand_x1_sg U50625 ( .A(n16117), .B(n16118), .X(n15873) );
  nand_x1_sg U50626 ( .A(n15873), .B(n15872), .X(n15870) );
  nand_x1_sg U50627 ( .A(n16071), .B(n15870), .X(n15878) );
  nand_x1_sg U50628 ( .A(n16180), .B(n50098), .X(n15891) );
  nand_x1_sg U50629 ( .A(n16068), .B(n16069), .X(n15890) );
  nand_x1_sg U50630 ( .A(n50079), .B(n15883), .X(n16069) );
  inv_x1_sg U50631 ( .A(n15971), .X(n50267) );
  nand_x1_sg U50632 ( .A(n15940), .B(n50244), .X(n15938) );
  nand_x1_sg U50633 ( .A(n15943), .B(n15942), .X(n15940) );
  nor_x1_sg U50634 ( .A(n16904), .B(n16905), .X(n16664) );
  nand_x1_sg U50635 ( .A(n16895), .B(n16896), .X(n16676) );
  nand_x1_sg U50636 ( .A(n16934), .B(n16935), .X(n16690) );
  nand_x1_sg U50637 ( .A(n16690), .B(n16689), .X(n16687) );
  nand_x1_sg U50638 ( .A(n16890), .B(n16687), .X(n16695) );
  nand_x1_sg U50639 ( .A(n16996), .B(n50383), .X(n16708) );
  nand_x1_sg U50640 ( .A(n16887), .B(n16888), .X(n16707) );
  nand_x1_sg U50641 ( .A(n50364), .B(n16700), .X(n16888) );
  inv_x1_sg U50642 ( .A(n16788), .X(n50553) );
  nand_x1_sg U50643 ( .A(n16757), .B(n50529), .X(n16755) );
  nand_x1_sg U50644 ( .A(n16760), .B(n16759), .X(n16757) );
  nand_x1_sg U50645 ( .A(n26475), .B(n26476), .X(n26474) );
  nor_x1_sg U50646 ( .A(n17723), .B(n17724), .X(n17485) );
  nand_x1_sg U50647 ( .A(n17714), .B(n17715), .X(n17497) );
  nand_x1_sg U50648 ( .A(n17755), .B(n17756), .X(n17511) );
  nand_x1_sg U50649 ( .A(n17511), .B(n17510), .X(n17508) );
  nand_x1_sg U50650 ( .A(n17709), .B(n17508), .X(n17516) );
  nand_x1_sg U50651 ( .A(n17818), .B(n50672), .X(n17529) );
  nand_x1_sg U50652 ( .A(n17706), .B(n17707), .X(n17528) );
  nand_x1_sg U50653 ( .A(n50653), .B(n17521), .X(n17707) );
  inv_x1_sg U50654 ( .A(n17609), .X(n50841) );
  nand_x1_sg U50655 ( .A(n17578), .B(n50818), .X(n17576) );
  nand_x1_sg U50656 ( .A(n17581), .B(n17580), .X(n17578) );
  nand_x1_sg U50657 ( .A(n26753), .B(n26754), .X(n26752) );
  nor_x1_sg U50658 ( .A(n18544), .B(n18545), .X(n18306) );
  nand_x1_sg U50659 ( .A(n18535), .B(n18536), .X(n18318) );
  nand_x1_sg U50660 ( .A(n18576), .B(n18577), .X(n18332) );
  nand_x1_sg U50661 ( .A(n18332), .B(n18331), .X(n18329) );
  nand_x1_sg U50662 ( .A(n18530), .B(n18329), .X(n18337) );
  nand_x1_sg U50663 ( .A(n18639), .B(n50959), .X(n18350) );
  nand_x1_sg U50664 ( .A(n18527), .B(n18528), .X(n18349) );
  nand_x1_sg U50665 ( .A(n50940), .B(n18342), .X(n18528) );
  inv_x1_sg U50666 ( .A(n18430), .X(n51128) );
  nand_x1_sg U50667 ( .A(n18399), .B(n51105), .X(n18397) );
  nand_x1_sg U50668 ( .A(n18402), .B(n18401), .X(n18399) );
  nor_x1_sg U50669 ( .A(n26761), .B(n26762), .X(n26760) );
  nand_x1_sg U50670 ( .A(n26768), .B(n26769), .X(n26761) );
  nand_x1_sg U50671 ( .A(n21757), .B(n45768), .X(n21756) );
  inv_x1_sg U50672 ( .A(n21758), .X(n45768) );
  nor_x1_sg U50673 ( .A(n21727), .B(n21728), .X(n21726) );
  nand_x1_sg U50674 ( .A(n21733), .B(n21734), .X(n21727) );
  nand_x1_sg U50675 ( .A(n21804), .B(n45725), .X(n21803) );
  inv_x1_sg U50676 ( .A(n21805), .X(n45725) );
  nor_x1_sg U50677 ( .A(n21774), .B(n21775), .X(n21773) );
  nand_x1_sg U50678 ( .A(n21780), .B(n21781), .X(n21774) );
  nand_x1_sg U50679 ( .A(n21851), .B(n45682), .X(n21850) );
  inv_x1_sg U50680 ( .A(n21852), .X(n45682) );
  nor_x1_sg U50681 ( .A(n21821), .B(n21822), .X(n21820) );
  nand_x1_sg U50682 ( .A(n21827), .B(n21828), .X(n21821) );
  nand_x1_sg U50683 ( .A(n21897), .B(n45638), .X(n21896) );
  inv_x1_sg U50684 ( .A(n21898), .X(n45638) );
  nor_x1_sg U50685 ( .A(n21868), .B(n21869), .X(n21867) );
  nand_x1_sg U50686 ( .A(n21874), .B(n21875), .X(n21868) );
  nand_x1_sg U50687 ( .A(n21944), .B(n45594), .X(n21943) );
  inv_x1_sg U50688 ( .A(n21945), .X(n45594) );
  nor_x1_sg U50689 ( .A(n21914), .B(n21915), .X(n21913) );
  nand_x1_sg U50690 ( .A(n21920), .B(n21921), .X(n21914) );
  nand_x1_sg U50691 ( .A(n21990), .B(n45549), .X(n21989) );
  inv_x1_sg U50692 ( .A(n21991), .X(n45549) );
  nor_x1_sg U50693 ( .A(n21961), .B(n21962), .X(n21960) );
  nand_x1_sg U50694 ( .A(n21967), .B(n21968), .X(n21961) );
  nand_x1_sg U50695 ( .A(n22037), .B(n45505), .X(n22036) );
  inv_x1_sg U50696 ( .A(n22038), .X(n45505) );
  nor_x1_sg U50697 ( .A(n22007), .B(n22008), .X(n22006) );
  nand_x1_sg U50698 ( .A(n22013), .B(n22014), .X(n22007) );
  nand_x1_sg U50699 ( .A(n22083), .B(n45457), .X(n22082) );
  inv_x1_sg U50700 ( .A(n22084), .X(n45457) );
  nor_x1_sg U50701 ( .A(n22054), .B(n22055), .X(n22053) );
  nand_x1_sg U50702 ( .A(n22060), .B(n22061), .X(n22054) );
  nand_x1_sg U50703 ( .A(n22131), .B(n45413), .X(n22130) );
  inv_x1_sg U50704 ( .A(n22132), .X(n45413) );
  nor_x1_sg U50705 ( .A(n22100), .B(n22101), .X(n22099) );
  nand_x1_sg U50706 ( .A(n22106), .B(n22107), .X(n22100) );
  nand_x1_sg U50707 ( .A(n22178), .B(n45367), .X(n22177) );
  inv_x1_sg U50708 ( .A(n22179), .X(n45367) );
  nor_x1_sg U50709 ( .A(n22148), .B(n22149), .X(n22147) );
  nand_x1_sg U50710 ( .A(n22154), .B(n22155), .X(n22148) );
  nand_x1_sg U50711 ( .A(n22226), .B(n45322), .X(n22225) );
  inv_x1_sg U50712 ( .A(n22227), .X(n45322) );
  nor_x1_sg U50713 ( .A(n22195), .B(n22196), .X(n22194) );
  nand_x1_sg U50714 ( .A(n22201), .B(n22202), .X(n22195) );
  nand_x1_sg U50715 ( .A(n22273), .B(n45277), .X(n22272) );
  inv_x1_sg U50716 ( .A(n22274), .X(n45277) );
  nor_x1_sg U50717 ( .A(n22243), .B(n22244), .X(n22242) );
  nand_x1_sg U50718 ( .A(n22249), .B(n22250), .X(n22243) );
  nand_x1_sg U50719 ( .A(n22321), .B(n45232), .X(n22320) );
  inv_x1_sg U50720 ( .A(n22322), .X(n45232) );
  nor_x1_sg U50721 ( .A(n22290), .B(n22291), .X(n22289) );
  nand_x1_sg U50722 ( .A(n22296), .B(n22297), .X(n22290) );
  nand_x1_sg U50723 ( .A(n22368), .B(n45186), .X(n22367) );
  inv_x1_sg U50724 ( .A(n22369), .X(n45186) );
  nor_x1_sg U50725 ( .A(n22338), .B(n22339), .X(n22337) );
  nand_x1_sg U50726 ( .A(n22344), .B(n22345), .X(n22338) );
  nand_x1_sg U50727 ( .A(n22416), .B(n45141), .X(n22415) );
  inv_x1_sg U50728 ( .A(n22417), .X(n45141) );
  nor_x1_sg U50729 ( .A(n22385), .B(n22386), .X(n22384) );
  nand_x1_sg U50730 ( .A(n22391), .B(n22392), .X(n22385) );
  nand_x1_sg U50731 ( .A(n22462), .B(n45094), .X(n22461) );
  inv_x1_sg U50732 ( .A(n22463), .X(n45094) );
  nor_x1_sg U50733 ( .A(n22433), .B(n22434), .X(n22432) );
  nand_x1_sg U50734 ( .A(n22439), .B(n22440), .X(n22433) );
  nand_x1_sg U50735 ( .A(n22508), .B(n45050), .X(n22507) );
  inv_x1_sg U50736 ( .A(n22509), .X(n45050) );
  nor_x1_sg U50737 ( .A(n22479), .B(n22480), .X(n22478) );
  nand_x1_sg U50738 ( .A(n22485), .B(n22486), .X(n22479) );
  nor_x1_sg U50739 ( .A(n22525), .B(n22526), .X(n22524) );
  nand_x1_sg U50740 ( .A(n22529), .B(n22530), .X(n22525) );
  nor_x1_sg U50741 ( .A(n22561), .B(n22562), .X(n22560) );
  nand_x1_sg U50742 ( .A(n22567), .B(n22568), .X(n22561) );
  nand_x1_sg U50743 ( .A(n7009), .B(n22717), .X(n22702) );
  nor_x1_sg U50744 ( .A(n26033), .B(n26034), .X(n26029) );
  nand_x1_sg U50745 ( .A(n40221), .B(n19108), .X(n19106) );
  nor_x1_sg U50746 ( .A(n20559), .B(n20560), .X(n19109) );
  nor_x1_sg U50747 ( .A(n19111), .B(n19112), .X(n19110) );
  nand_x1_sg U50748 ( .A(n40222), .B(n5955), .X(n5952) );
  nor_x1_sg U50749 ( .A(n5990), .B(n5991), .X(n5956) );
  nor_x1_sg U50750 ( .A(n5958), .B(n5959), .X(n5957) );
  nand_x1_sg U50751 ( .A(n40090), .B(n6010), .X(n6008) );
  nor_x1_sg U50752 ( .A(n6039), .B(n6040), .X(n6011) );
  nor_x1_sg U50753 ( .A(n6013), .B(n6014), .X(n6012) );
  nand_x1_sg U50754 ( .A(n41417), .B(n6059), .X(n6057) );
  nor_x1_sg U50755 ( .A(n6089), .B(n6090), .X(n6060) );
  nor_x1_sg U50756 ( .A(n6062), .B(n6063), .X(n6061) );
  nand_x1_sg U50757 ( .A(n41419), .B(n6107), .X(n6105) );
  nor_x1_sg U50758 ( .A(n6135), .B(n6136), .X(n6108) );
  nor_x1_sg U50759 ( .A(n6110), .B(n6111), .X(n6109) );
  nand_x1_sg U50760 ( .A(n40221), .B(n6152), .X(n6150) );
  nor_x1_sg U50761 ( .A(n6180), .B(n6181), .X(n6153) );
  nor_x1_sg U50762 ( .A(n6155), .B(n6156), .X(n6154) );
  nand_x1_sg U50763 ( .A(n40222), .B(n6198), .X(n6196) );
  nor_x1_sg U50764 ( .A(n6227), .B(n6228), .X(n6199) );
  nor_x1_sg U50765 ( .A(n6201), .B(n6202), .X(n6200) );
  nand_x1_sg U50766 ( .A(n41419), .B(n6245), .X(n6243) );
  nor_x1_sg U50767 ( .A(n6271), .B(n6272), .X(n6246) );
  nor_x1_sg U50768 ( .A(n6248), .B(n6249), .X(n6247) );
  nand_x1_sg U50769 ( .A(n41418), .B(n6290), .X(n6288) );
  nor_x1_sg U50770 ( .A(n6316), .B(n6317), .X(n6291) );
  nor_x1_sg U50771 ( .A(n6293), .B(n6294), .X(n6292) );
  nand_x1_sg U50772 ( .A(n40222), .B(n6334), .X(n6332) );
  nor_x1_sg U50773 ( .A(n6360), .B(n6361), .X(n6335) );
  nor_x1_sg U50774 ( .A(n6337), .B(n6338), .X(n6336) );
  nand_x1_sg U50775 ( .A(n40090), .B(n6379), .X(n6377) );
  nor_x1_sg U50776 ( .A(n6405), .B(n6406), .X(n6380) );
  nor_x1_sg U50777 ( .A(n6382), .B(n6383), .X(n6381) );
  nand_x1_sg U50778 ( .A(n40222), .B(n6423), .X(n6421) );
  nor_x1_sg U50779 ( .A(n6449), .B(n6450), .X(n6424) );
  nor_x1_sg U50780 ( .A(n6426), .B(n6427), .X(n6425) );
  nand_x1_sg U50781 ( .A(n39434), .B(n6468), .X(n6466) );
  nor_x1_sg U50782 ( .A(n6494), .B(n6495), .X(n6469) );
  nor_x1_sg U50783 ( .A(n6471), .B(n6472), .X(n6470) );
  nand_x1_sg U50784 ( .A(n39435), .B(n6512), .X(n6510) );
  nor_x1_sg U50785 ( .A(n6538), .B(n6539), .X(n6513) );
  nor_x1_sg U50786 ( .A(n6515), .B(n6516), .X(n6514) );
  nand_x1_sg U50787 ( .A(n40089), .B(n6557), .X(n6555) );
  nor_x1_sg U50788 ( .A(n6583), .B(n6584), .X(n6558) );
  nor_x1_sg U50789 ( .A(n6560), .B(n6561), .X(n6559) );
  nand_x1_sg U50790 ( .A(n41420), .B(n6601), .X(n6599) );
  nor_x1_sg U50791 ( .A(n6627), .B(n6628), .X(n6602) );
  nor_x1_sg U50792 ( .A(n6604), .B(n6605), .X(n6603) );
  nand_x1_sg U50793 ( .A(n38983), .B(n6646), .X(n6644) );
  nor_x1_sg U50794 ( .A(n6675), .B(n6676), .X(n6647) );
  nor_x1_sg U50795 ( .A(n6649), .B(n6650), .X(n6648) );
  nand_x1_sg U50796 ( .A(n38983), .B(n6694), .X(n6692) );
  nor_x1_sg U50797 ( .A(n6719), .B(n6720), .X(n6695) );
  nor_x1_sg U50798 ( .A(n6697), .B(n6698), .X(n6696) );
  nand_x1_sg U50799 ( .A(n41420), .B(n6734), .X(n6732) );
  nor_x1_sg U50800 ( .A(n6765), .B(n6766), .X(n6735) );
  nor_x1_sg U50801 ( .A(n6737), .B(n6738), .X(n6736) );
  nand_x1_sg U50802 ( .A(n40090), .B(n6785), .X(n6783) );
  nor_x1_sg U50803 ( .A(n6808), .B(n6809), .X(n6786) );
  nor_x1_sg U50804 ( .A(n6788), .B(n6789), .X(n6787) );
  inv_x1_sg U50805 ( .A(n6838), .X(n46855) );
  nand_x1_sg U50806 ( .A(n46862), .B(n6844), .X(n6842) );
  inv_x1_sg U50807 ( .A(n6853), .X(n46873) );
  inv_x1_sg U50808 ( .A(n6860), .X(n46885) );
  inv_x1_sg U50809 ( .A(n6878), .X(n46932) );
  inv_x1_sg U50810 ( .A(n6890), .X(n46980) );
  inv_x1_sg U50811 ( .A(n6896), .X(n47003) );
  inv_x1_sg U50812 ( .A(n6902), .X(n47017) );
  inv_x1_sg U50813 ( .A(n6908), .X(n47043) );
  inv_x1_sg U50814 ( .A(n6914), .X(n47071) );
  inv_x1_sg U50815 ( .A(n6920), .X(n47093) );
  inv_x1_sg U50816 ( .A(n6926), .X(n47118) );
  inv_x1_sg U50817 ( .A(n6930), .X(n47126) );
  inv_x1_sg U50818 ( .A(n7655), .X(n47148) );
  inv_x1_sg U50819 ( .A(n7670), .X(n47166) );
  inv_x1_sg U50820 ( .A(n7677), .X(n47178) );
  inv_x1_sg U50821 ( .A(n7695), .X(n47224) );
  inv_x1_sg U50822 ( .A(n7707), .X(n47270) );
  inv_x1_sg U50823 ( .A(n7713), .X(n47292) );
  inv_x1_sg U50824 ( .A(n7719), .X(n47305) );
  inv_x1_sg U50825 ( .A(n7725), .X(n47330) );
  inv_x1_sg U50826 ( .A(n7731), .X(n47357) );
  inv_x1_sg U50827 ( .A(n7737), .X(n47379) );
  inv_x1_sg U50828 ( .A(n7743), .X(n47404) );
  inv_x1_sg U50829 ( .A(n7747), .X(n47412) );
  inv_x1_sg U50830 ( .A(n8473), .X(n47433) );
  inv_x1_sg U50831 ( .A(n8488), .X(n47451) );
  inv_x1_sg U50832 ( .A(n8495), .X(n47463) );
  inv_x1_sg U50833 ( .A(n8513), .X(n47509) );
  inv_x1_sg U50834 ( .A(n8525), .X(n47555) );
  inv_x1_sg U50835 ( .A(n8531), .X(n47577) );
  inv_x1_sg U50836 ( .A(n8537), .X(n47590) );
  inv_x1_sg U50837 ( .A(n8543), .X(n47615) );
  inv_x1_sg U50838 ( .A(n8549), .X(n47642) );
  inv_x1_sg U50839 ( .A(n8555), .X(n47664) );
  inv_x1_sg U50840 ( .A(n8561), .X(n47689) );
  inv_x1_sg U50841 ( .A(n8565), .X(n47697) );
  inv_x1_sg U50842 ( .A(n9293), .X(n47718) );
  inv_x1_sg U50843 ( .A(n9308), .X(n47736) );
  inv_x1_sg U50844 ( .A(n9315), .X(n47748) );
  inv_x1_sg U50845 ( .A(n9333), .X(n47794) );
  inv_x1_sg U50846 ( .A(n9345), .X(n47840) );
  inv_x1_sg U50847 ( .A(n9351), .X(n47862) );
  inv_x1_sg U50848 ( .A(n9357), .X(n47875) );
  inv_x1_sg U50849 ( .A(n9363), .X(n47900) );
  inv_x1_sg U50850 ( .A(n9369), .X(n47927) );
  inv_x1_sg U50851 ( .A(n9375), .X(n47949) );
  inv_x1_sg U50852 ( .A(n9381), .X(n47974) );
  inv_x1_sg U50853 ( .A(n9385), .X(n47982) );
  inv_x1_sg U50854 ( .A(n10112), .X(n48003) );
  inv_x1_sg U50855 ( .A(n10127), .X(n48021) );
  inv_x1_sg U50856 ( .A(n10134), .X(n48033) );
  inv_x1_sg U50857 ( .A(n10152), .X(n48079) );
  inv_x1_sg U50858 ( .A(n10164), .X(n48125) );
  inv_x1_sg U50859 ( .A(n10170), .X(n48147) );
  inv_x1_sg U50860 ( .A(n10176), .X(n48160) );
  inv_x1_sg U50861 ( .A(n10182), .X(n48185) );
  inv_x1_sg U50862 ( .A(n10188), .X(n48212) );
  inv_x1_sg U50863 ( .A(n10194), .X(n48234) );
  inv_x1_sg U50864 ( .A(n10200), .X(n48259) );
  inv_x1_sg U50865 ( .A(n10204), .X(n48267) );
  inv_x1_sg U50866 ( .A(n10931), .X(n48288) );
  inv_x1_sg U50867 ( .A(n10946), .X(n48306) );
  inv_x1_sg U50868 ( .A(n10953), .X(n48318) );
  inv_x1_sg U50869 ( .A(n10971), .X(n48364) );
  inv_x1_sg U50870 ( .A(n10983), .X(n48410) );
  inv_x1_sg U50871 ( .A(n10989), .X(n48432) );
  inv_x1_sg U50872 ( .A(n10995), .X(n48445) );
  inv_x1_sg U50873 ( .A(n11001), .X(n48470) );
  inv_x1_sg U50874 ( .A(n11007), .X(n48497) );
  inv_x1_sg U50875 ( .A(n11013), .X(n48519) );
  inv_x1_sg U50876 ( .A(n11019), .X(n48544) );
  inv_x1_sg U50877 ( .A(n11023), .X(n48552) );
  inv_x1_sg U50878 ( .A(n11750), .X(n48573) );
  inv_x1_sg U50879 ( .A(n11765), .X(n48591) );
  inv_x1_sg U50880 ( .A(n11772), .X(n48603) );
  inv_x1_sg U50881 ( .A(n11790), .X(n48649) );
  inv_x1_sg U50882 ( .A(n11802), .X(n48695) );
  inv_x1_sg U50883 ( .A(n11808), .X(n48717) );
  inv_x1_sg U50884 ( .A(n11814), .X(n48730) );
  inv_x1_sg U50885 ( .A(n11820), .X(n48755) );
  inv_x1_sg U50886 ( .A(n11826), .X(n48782) );
  inv_x1_sg U50887 ( .A(n11832), .X(n48804) );
  inv_x1_sg U50888 ( .A(n11838), .X(n48829) );
  inv_x1_sg U50889 ( .A(n11842), .X(n48837) );
  inv_x1_sg U50890 ( .A(n12569), .X(n48859) );
  inv_x1_sg U50891 ( .A(n12584), .X(n48877) );
  inv_x1_sg U50892 ( .A(n12591), .X(n48889) );
  inv_x1_sg U50893 ( .A(n12609), .X(n48935) );
  inv_x1_sg U50894 ( .A(n12621), .X(n48981) );
  inv_x1_sg U50895 ( .A(n12627), .X(n49003) );
  inv_x1_sg U50896 ( .A(n12633), .X(n49016) );
  inv_x1_sg U50897 ( .A(n12639), .X(n49041) );
  inv_x1_sg U50898 ( .A(n12645), .X(n49069) );
  inv_x1_sg U50899 ( .A(n12651), .X(n49091) );
  inv_x1_sg U50900 ( .A(n12657), .X(n49116) );
  inv_x1_sg U50901 ( .A(n12661), .X(n49124) );
  inv_x1_sg U50902 ( .A(n13388), .X(n49146) );
  inv_x1_sg U50903 ( .A(n13403), .X(n49164) );
  inv_x1_sg U50904 ( .A(n13410), .X(n49176) );
  inv_x1_sg U50905 ( .A(n13428), .X(n49222) );
  inv_x1_sg U50906 ( .A(n13440), .X(n49268) );
  inv_x1_sg U50907 ( .A(n13446), .X(n49290) );
  inv_x1_sg U50908 ( .A(n13452), .X(n49303) );
  inv_x1_sg U50909 ( .A(n13458), .X(n49328) );
  inv_x1_sg U50910 ( .A(n13464), .X(n49355) );
  inv_x1_sg U50911 ( .A(n13470), .X(n49377) );
  inv_x1_sg U50912 ( .A(n13476), .X(n49402) );
  inv_x1_sg U50913 ( .A(n13480), .X(n49410) );
  inv_x1_sg U50914 ( .A(n14207), .X(n49432) );
  inv_x1_sg U50915 ( .A(n14222), .X(n49450) );
  inv_x1_sg U50916 ( .A(n14229), .X(n49462) );
  inv_x1_sg U50917 ( .A(n14247), .X(n49508) );
  inv_x1_sg U50918 ( .A(n14259), .X(n49554) );
  inv_x1_sg U50919 ( .A(n14265), .X(n49576) );
  inv_x1_sg U50920 ( .A(n14271), .X(n49589) );
  inv_x1_sg U50921 ( .A(n14277), .X(n49614) );
  inv_x1_sg U50922 ( .A(n14283), .X(n49641) );
  inv_x1_sg U50923 ( .A(n14289), .X(n49663) );
  inv_x1_sg U50924 ( .A(n14295), .X(n49688) );
  inv_x1_sg U50925 ( .A(n14299), .X(n49696) );
  inv_x1_sg U50926 ( .A(n15026), .X(n49717) );
  inv_x1_sg U50927 ( .A(n15041), .X(n49735) );
  inv_x1_sg U50928 ( .A(n15048), .X(n49747) );
  inv_x1_sg U50929 ( .A(n15066), .X(n49794) );
  inv_x1_sg U50930 ( .A(n15078), .X(n49840) );
  inv_x1_sg U50931 ( .A(n15084), .X(n49862) );
  inv_x1_sg U50932 ( .A(n15090), .X(n49875) );
  inv_x1_sg U50933 ( .A(n15096), .X(n49900) );
  inv_x1_sg U50934 ( .A(n15102), .X(n49927) );
  inv_x1_sg U50935 ( .A(n15108), .X(n49949) );
  inv_x1_sg U50936 ( .A(n15114), .X(n49974) );
  inv_x1_sg U50937 ( .A(n15118), .X(n49982) );
  inv_x1_sg U50938 ( .A(n15845), .X(n50004) );
  inv_x1_sg U50939 ( .A(n15860), .X(n50022) );
  inv_x1_sg U50940 ( .A(n15867), .X(n50034) );
  inv_x1_sg U50941 ( .A(n15885), .X(n50080) );
  inv_x1_sg U50942 ( .A(n15897), .X(n50126) );
  inv_x1_sg U50943 ( .A(n15903), .X(n50148) );
  inv_x1_sg U50944 ( .A(n15909), .X(n50161) );
  inv_x1_sg U50945 ( .A(n15915), .X(n50186) );
  inv_x1_sg U50946 ( .A(n15921), .X(n50213) );
  inv_x1_sg U50947 ( .A(n15927), .X(n50235) );
  inv_x1_sg U50948 ( .A(n15933), .X(n50260) );
  inv_x1_sg U50949 ( .A(n15937), .X(n50268) );
  inv_x1_sg U50950 ( .A(n16662), .X(n50287) );
  inv_x1_sg U50951 ( .A(n16677), .X(n50307) );
  inv_x1_sg U50952 ( .A(n16684), .X(n50319) );
  inv_x1_sg U50953 ( .A(n16702), .X(n50365) );
  inv_x1_sg U50954 ( .A(n16714), .X(n50411) );
  inv_x1_sg U50955 ( .A(n16720), .X(n50433) );
  inv_x1_sg U50956 ( .A(n16726), .X(n50446) );
  inv_x1_sg U50957 ( .A(n16732), .X(n50471) );
  inv_x1_sg U50958 ( .A(n16738), .X(n50498) );
  inv_x1_sg U50959 ( .A(n16744), .X(n50520) );
  inv_x1_sg U50960 ( .A(n16750), .X(n50545) );
  inv_x1_sg U50961 ( .A(n16754), .X(n50554) );
  inv_x1_sg U50962 ( .A(n17483), .X(n50578) );
  inv_x1_sg U50963 ( .A(n17498), .X(n50596) );
  inv_x1_sg U50964 ( .A(n17505), .X(n50608) );
  inv_x1_sg U50965 ( .A(n17523), .X(n50654) );
  inv_x1_sg U50966 ( .A(n17535), .X(n50700) );
  inv_x1_sg U50967 ( .A(n17541), .X(n50722) );
  inv_x1_sg U50968 ( .A(n17547), .X(n50735) );
  inv_x1_sg U50969 ( .A(n17553), .X(n50760) );
  inv_x1_sg U50970 ( .A(n17559), .X(n50787) );
  inv_x1_sg U50971 ( .A(n17565), .X(n50809) );
  inv_x1_sg U50972 ( .A(n17571), .X(n50834) );
  nand_x1_sg U50973 ( .A(n41117), .B(n41418), .X(n17466) );
  inv_x1_sg U50974 ( .A(n17575), .X(n50842) );
  inv_x1_sg U50975 ( .A(n18304), .X(n50865) );
  inv_x1_sg U50976 ( .A(n18319), .X(n50883) );
  inv_x1_sg U50977 ( .A(n18326), .X(n50895) );
  inv_x1_sg U50978 ( .A(n18344), .X(n50941) );
  inv_x1_sg U50979 ( .A(n18356), .X(n50987) );
  inv_x1_sg U50980 ( .A(n18362), .X(n51009) );
  inv_x1_sg U50981 ( .A(n18368), .X(n51022) );
  inv_x1_sg U50982 ( .A(n18374), .X(n51047) );
  inv_x1_sg U50983 ( .A(n18380), .X(n51074) );
  inv_x1_sg U50984 ( .A(n18386), .X(n51096) );
  inv_x1_sg U50985 ( .A(n18392), .X(n51121) );
  inv_x1_sg U50986 ( .A(n18396), .X(n51129) );
  nand_x1_sg U50987 ( .A(n26788), .B(n26789), .X(n26787) );
  nand_x1_sg U50988 ( .A(n26794), .B(n26795), .X(n26793) );
  nand_x1_sg U50989 ( .A(n26782), .B(n26783), .X(n5941) );
  nand_x1_sg U50990 ( .A(n28517), .B(n28518), .X(n5938) );
  nand_x1_sg U50991 ( .A(n20962), .B(n26827), .X(n28517) );
  nand_x1_sg U50992 ( .A(n21749), .B(n21750), .X(n21748) );
  nand_x1_sg U50993 ( .A(n21754), .B(n21755), .X(n21753) );
  nand_x1_sg U50994 ( .A(n21743), .B(n21744), .X(n5897) );
  nand_x1_sg U50995 ( .A(n21764), .B(n21765), .X(n5894) );
  nand_x1_sg U50996 ( .A(n21796), .B(n21797), .X(n21795) );
  nand_x1_sg U50997 ( .A(n21801), .B(n21802), .X(n21800) );
  nand_x1_sg U50998 ( .A(n21790), .B(n21791), .X(n5920) );
  nand_x1_sg U50999 ( .A(n21811), .B(n21812), .X(n5917) );
  nand_x1_sg U51000 ( .A(n21843), .B(n21844), .X(n21842) );
  nand_x1_sg U51001 ( .A(n21848), .B(n21849), .X(n21847) );
  nand_x1_sg U51002 ( .A(n21837), .B(n21838), .X(n5785) );
  nand_x1_sg U51003 ( .A(n21858), .B(n21859), .X(n5782) );
  nand_x1_sg U51004 ( .A(n21889), .B(n21890), .X(n21888) );
  nand_x1_sg U51005 ( .A(n21894), .B(n21895), .X(n21893) );
  nand_x1_sg U51006 ( .A(n21884), .B(n21885), .X(n5856) );
  nand_x1_sg U51007 ( .A(n21904), .B(n21905), .X(n5853) );
  nand_x1_sg U51008 ( .A(n21936), .B(n21937), .X(n21935) );
  nand_x1_sg U51009 ( .A(n21941), .B(n21942), .X(n21940) );
  nand_x1_sg U51010 ( .A(n21930), .B(n21931), .X(n5849) );
  nand_x1_sg U51011 ( .A(n21951), .B(n21952), .X(n5846) );
  nand_x1_sg U51012 ( .A(n21982), .B(n21983), .X(n21981) );
  nand_x1_sg U51013 ( .A(n21987), .B(n21988), .X(n21986) );
  nand_x1_sg U51014 ( .A(n21977), .B(n21978), .X(n5911) );
  nand_x1_sg U51015 ( .A(n21997), .B(n21998), .X(n5908) );
  nand_x1_sg U51016 ( .A(n38930), .B(n21999), .X(n21998) );
  nand_x1_sg U51017 ( .A(n22029), .B(n22030), .X(n22028) );
  nand_x1_sg U51018 ( .A(n22034), .B(n22035), .X(n22033) );
  nand_x1_sg U51019 ( .A(n22023), .B(n22024), .X(n5872) );
  nand_x1_sg U51020 ( .A(n22044), .B(n22045), .X(n5869) );
  nand_x1_sg U51021 ( .A(n22075), .B(n22076), .X(n22074) );
  nand_x1_sg U51022 ( .A(n22080), .B(n22081), .X(n22079) );
  nand_x1_sg U51023 ( .A(n22070), .B(n22071), .X(n5890) );
  nand_x1_sg U51024 ( .A(n22090), .B(n22091), .X(n5887) );
  nand_x1_sg U51025 ( .A(n41095), .B(n22092), .X(n22091) );
  nand_x1_sg U51026 ( .A(n22123), .B(n22124), .X(n22122) );
  nand_x1_sg U51027 ( .A(n22128), .B(n22129), .X(n22127) );
  nand_x1_sg U51028 ( .A(n22117), .B(n22118), .X(n5795) );
  nand_x1_sg U51029 ( .A(n22138), .B(n22139), .X(n5792) );
  nand_x1_sg U51030 ( .A(n22170), .B(n22171), .X(n22169) );
  nand_x1_sg U51031 ( .A(n22175), .B(n22176), .X(n22174) );
  nand_x1_sg U51032 ( .A(n22165), .B(n22166), .X(n5818) );
  nand_x1_sg U51033 ( .A(n22185), .B(n22186), .X(n5815) );
  nand_x1_sg U51034 ( .A(n22218), .B(n22219), .X(n22217) );
  nand_x1_sg U51035 ( .A(n22223), .B(n22224), .X(n22222) );
  nand_x1_sg U51036 ( .A(n22212), .B(n22213), .X(n5927) );
  nand_x1_sg U51037 ( .A(n22233), .B(n22234), .X(n5924) );
  nand_x1_sg U51038 ( .A(n41095), .B(n22235), .X(n22234) );
  nand_x1_sg U51039 ( .A(n22265), .B(n22266), .X(n22264) );
  nand_x1_sg U51040 ( .A(n22270), .B(n22271), .X(n22269) );
  nand_x1_sg U51041 ( .A(n22260), .B(n22261), .X(n5811) );
  nand_x1_sg U51042 ( .A(n22280), .B(n22281), .X(n5808) );
  nand_x1_sg U51043 ( .A(n38930), .B(n22282), .X(n22281) );
  nand_x1_sg U51044 ( .A(n22313), .B(n22314), .X(n22312) );
  nand_x1_sg U51045 ( .A(n22318), .B(n22319), .X(n22317) );
  nand_x1_sg U51046 ( .A(n22307), .B(n22308), .X(n5881) );
  nand_x1_sg U51047 ( .A(n22328), .B(n22329), .X(n5878) );
  nand_x1_sg U51048 ( .A(n22360), .B(n22361), .X(n22359) );
  nand_x1_sg U51049 ( .A(n22365), .B(n22366), .X(n22364) );
  nand_x1_sg U51050 ( .A(n22355), .B(n22356), .X(n5840) );
  nand_x1_sg U51051 ( .A(n22375), .B(n22376), .X(n5837) );
  nand_x1_sg U51052 ( .A(n41094), .B(n22377), .X(n22376) );
  nand_x1_sg U51053 ( .A(n22408), .B(n22409), .X(n22407) );
  nand_x1_sg U51054 ( .A(n22413), .B(n22414), .X(n22412) );
  nand_x1_sg U51055 ( .A(n22402), .B(n22403), .X(n5804) );
  nand_x1_sg U51056 ( .A(n22423), .B(n22424), .X(n5801) );
  nand_x1_sg U51057 ( .A(n38930), .B(n22425), .X(n22424) );
  nand_x1_sg U51058 ( .A(n22454), .B(n22455), .X(n22453) );
  nand_x1_sg U51059 ( .A(n38938), .B(n22456), .X(n22455) );
  nand_x1_sg U51060 ( .A(n22459), .B(n22460), .X(n22458) );
  nand_x1_sg U51061 ( .A(n22449), .B(n22450), .X(n5825) );
  nand_x1_sg U51062 ( .A(n22469), .B(n22470), .X(n5822) );
  nand_x1_sg U51063 ( .A(n39259), .B(n22471), .X(n22470) );
  nand_x1_sg U51064 ( .A(n22500), .B(n22501), .X(n22499) );
  nand_x1_sg U51065 ( .A(n41110), .B(n22502), .X(n22501) );
  nand_x1_sg U51066 ( .A(n22505), .B(n22506), .X(n22504) );
  nand_x1_sg U51067 ( .A(n22494), .B(n22495), .X(n5904) );
  nand_x1_sg U51068 ( .A(n22515), .B(n22516), .X(n5901) );
  nand_x1_sg U51069 ( .A(n22540), .B(n22541), .X(n22539) );
  nand_x1_sg U51070 ( .A(n22543), .B(n22544), .X(n22542) );
  nand_x1_sg U51071 ( .A(n22536), .B(n22537), .X(n5948) );
  nand_x1_sg U51072 ( .A(n22553), .B(n22554), .X(n5945) );
  nand_x1_sg U51073 ( .A(n22581), .B(n22582), .X(n22580) );
  nand_x1_sg U51074 ( .A(n22586), .B(n22587), .X(n22585) );
  nand_x1_sg U51075 ( .A(n22576), .B(n22577), .X(n5934) );
  nand_x1_sg U51076 ( .A(n22592), .B(n22593), .X(n5931) );
  nand_x2_sg U51077 ( .A(n22596), .B(n22597), .X(n5771) );
  nand_x2_sg U51078 ( .A(n22602), .B(n22603), .X(n5788) );
  nand_x2_sg U51079 ( .A(n22608), .B(n22609), .X(n5913) );
  nand_x2_sg U51080 ( .A(n22614), .B(n22615), .X(n5865) );
  nand_x2_sg U51081 ( .A(n22620), .B(n22621), .X(n5842) );
  nand_x2_sg U51082 ( .A(n22626), .B(n22627), .X(n5773) );
  nor_x1_sg U51083 ( .A(n22633), .B(n22634), .X(n5786) );
  nand_x2_sg U51084 ( .A(n22640), .B(n22641), .X(n5874) );
  nand_x2_sg U51085 ( .A(n22646), .B(n22647), .X(n5829) );
  nand_x2_sg U51086 ( .A(n22651), .B(n22652), .X(n5777) );
  nand_x2_sg U51087 ( .A(n22658), .B(n22659), .X(n5863) );
  nand_x2_sg U51088 ( .A(n22664), .B(n22665), .X(n5827) );
  nand_x2_sg U51089 ( .A(n22670), .B(n22671), .X(n5775) );
  nand_x2_sg U51090 ( .A(n22676), .B(n22677), .X(n5833) );
  nand_x2_sg U51091 ( .A(n22682), .B(n22683), .X(n5883) );
  nand_x1_sg U51092 ( .A(n39478), .B(n22688), .X(n5950) );
  nand_x1_sg U51093 ( .A(n22692), .B(n40217), .X(n5797) );
  nand_x2_sg U51094 ( .A(n22699), .B(n22700), .X(n5831) );
  nand_x4_sg U51095 ( .A(n22856), .B(n22857), .X(n22855) );
  nand_x4_sg U51096 ( .A(n22864), .B(n22865), .X(n22863) );
  nand_x4_sg U51097 ( .A(n22871), .B(n22872), .X(n22870) );
  nand_x4_sg U51098 ( .A(n22878), .B(n22879), .X(n22877) );
  nand_x4_sg U51099 ( .A(n22885), .B(n22886), .X(n22884) );
  nand_x4_sg U51100 ( .A(n22892), .B(n22893), .X(n22891) );
  nor_x1_sg U51101 ( .A(n22899), .B(n22900), .X(n22898) );
  nor_x1_sg U51102 ( .A(n22906), .B(n22907), .X(n22905) );
  nand_x4_sg U51103 ( .A(n22913), .B(n22914), .X(n22912) );
  nor_x1_sg U51104 ( .A(n22920), .B(n22921), .X(n22919) );
  nand_x4_sg U51105 ( .A(n22927), .B(n22928), .X(n22926) );
  nor_x1_sg U51106 ( .A(n22934), .B(n22935), .X(n22933) );
  nand_x4_sg U51107 ( .A(n22941), .B(n22942), .X(n22940) );
  nor_x1_sg U51108 ( .A(n22948), .B(n22949), .X(n22947) );
  nand_x4_sg U51109 ( .A(n22955), .B(n22956), .X(n22954) );
  nand_x1_sg U51110 ( .A(n40217), .B(n22962), .X(n22961) );
  nand_x1_sg U51111 ( .A(n22967), .B(n39928), .X(n22966) );
  nor_x1_sg U51112 ( .A(n22974), .B(n22975), .X(n22973) );
  nand_x4_sg U51113 ( .A(n23133), .B(n23134), .X(n23132) );
  nand_x4_sg U51114 ( .A(n23141), .B(n23142), .X(n23140) );
  nand_x4_sg U51115 ( .A(n23148), .B(n23149), .X(n23147) );
  nand_x4_sg U51116 ( .A(n23155), .B(n23156), .X(n23154) );
  nand_x4_sg U51117 ( .A(n23162), .B(n23163), .X(n23161) );
  nand_x4_sg U51118 ( .A(n23169), .B(n23170), .X(n23168) );
  nor_x1_sg U51119 ( .A(n23176), .B(n23177), .X(n23175) );
  nor_x1_sg U51120 ( .A(n23183), .B(n23184), .X(n23182) );
  nand_x4_sg U51121 ( .A(n23190), .B(n23191), .X(n23189) );
  nor_x1_sg U51122 ( .A(n23197), .B(n23198), .X(n23196) );
  nand_x4_sg U51123 ( .A(n23204), .B(n23205), .X(n23203) );
  nor_x1_sg U51124 ( .A(n23211), .B(n23212), .X(n23210) );
  nand_x4_sg U51125 ( .A(n23218), .B(n23219), .X(n23217) );
  nor_x1_sg U51126 ( .A(n23225), .B(n23226), .X(n23224) );
  nand_x4_sg U51127 ( .A(n23232), .B(n23233), .X(n23231) );
  nand_x1_sg U51128 ( .A(n40217), .B(n23239), .X(n23238) );
  nand_x1_sg U51129 ( .A(n23244), .B(n39279), .X(n23243) );
  nor_x1_sg U51130 ( .A(n23251), .B(n23252), .X(n23250) );
  nand_x4_sg U51131 ( .A(n23413), .B(n23414), .X(n23412) );
  nand_x4_sg U51132 ( .A(n23421), .B(n23422), .X(n23420) );
  nand_x4_sg U51133 ( .A(n23428), .B(n23429), .X(n23427) );
  nand_x4_sg U51134 ( .A(n23435), .B(n23436), .X(n23434) );
  nand_x4_sg U51135 ( .A(n23442), .B(n23443), .X(n23441) );
  nand_x4_sg U51136 ( .A(n23449), .B(n23450), .X(n23448) );
  nor_x1_sg U51137 ( .A(n23456), .B(n23457), .X(n23455) );
  nor_x1_sg U51138 ( .A(n23463), .B(n23464), .X(n23462) );
  nand_x4_sg U51139 ( .A(n23470), .B(n23471), .X(n23469) );
  nor_x1_sg U51140 ( .A(n23477), .B(n23478), .X(n23476) );
  nand_x4_sg U51141 ( .A(n23484), .B(n23485), .X(n23483) );
  nor_x1_sg U51142 ( .A(n23491), .B(n23492), .X(n23490) );
  nand_x4_sg U51143 ( .A(n23498), .B(n23499), .X(n23497) );
  nor_x1_sg U51144 ( .A(n23505), .B(n23506), .X(n23504) );
  nand_x4_sg U51145 ( .A(n23512), .B(n23513), .X(n23511) );
  nand_x1_sg U51146 ( .A(n41318), .B(n23519), .X(n23518) );
  nor_x1_sg U51147 ( .A(n23531), .B(n23532), .X(n23530) );
  nand_x4_sg U51148 ( .A(n23692), .B(n23693), .X(n23691) );
  nand_x4_sg U51149 ( .A(n23700), .B(n23701), .X(n23699) );
  nand_x4_sg U51150 ( .A(n23707), .B(n23708), .X(n23706) );
  nand_x4_sg U51151 ( .A(n23714), .B(n23715), .X(n23713) );
  nand_x4_sg U51152 ( .A(n23721), .B(n23722), .X(n23720) );
  nand_x4_sg U51153 ( .A(n23728), .B(n23729), .X(n23727) );
  nor_x1_sg U51154 ( .A(n23735), .B(n23736), .X(n23734) );
  nor_x1_sg U51155 ( .A(n23742), .B(n23743), .X(n23741) );
  nand_x4_sg U51156 ( .A(n23749), .B(n23750), .X(n23748) );
  nor_x1_sg U51157 ( .A(n23756), .B(n23757), .X(n23755) );
  nand_x4_sg U51158 ( .A(n23763), .B(n23764), .X(n23762) );
  nor_x1_sg U51159 ( .A(n23770), .B(n23771), .X(n23769) );
  nand_x4_sg U51160 ( .A(n23777), .B(n23778), .X(n23776) );
  nor_x1_sg U51161 ( .A(n23784), .B(n23785), .X(n23783) );
  nand_x4_sg U51162 ( .A(n23791), .B(n23792), .X(n23790) );
  nand_x1_sg U51163 ( .A(n41311), .B(n23798), .X(n23797) );
  nor_x1_sg U51164 ( .A(n23810), .B(n23811), .X(n23809) );
  nand_x4_sg U51165 ( .A(n23971), .B(n23972), .X(n23970) );
  nand_x4_sg U51166 ( .A(n23979), .B(n23980), .X(n23978) );
  nand_x4_sg U51167 ( .A(n23986), .B(n23987), .X(n23985) );
  nand_x4_sg U51168 ( .A(n23993), .B(n23994), .X(n23992) );
  nand_x4_sg U51169 ( .A(n24000), .B(n24001), .X(n23999) );
  nand_x4_sg U51170 ( .A(n24007), .B(n24008), .X(n24006) );
  nor_x1_sg U51171 ( .A(n24014), .B(n24015), .X(n24013) );
  nor_x1_sg U51172 ( .A(n24021), .B(n24022), .X(n24020) );
  nand_x4_sg U51173 ( .A(n24028), .B(n24029), .X(n24027) );
  nor_x1_sg U51174 ( .A(n24035), .B(n24036), .X(n24034) );
  nand_x4_sg U51175 ( .A(n24042), .B(n24043), .X(n24041) );
  nor_x1_sg U51176 ( .A(n24049), .B(n24050), .X(n24048) );
  nand_x4_sg U51177 ( .A(n24056), .B(n24057), .X(n24055) );
  nor_x1_sg U51178 ( .A(n24063), .B(n24064), .X(n24062) );
  nand_x4_sg U51179 ( .A(n24070), .B(n24071), .X(n24069) );
  nand_x1_sg U51180 ( .A(n41464), .B(n24077), .X(n24076) );
  nor_x1_sg U51181 ( .A(n24089), .B(n24090), .X(n24088) );
  nand_x4_sg U51182 ( .A(n24250), .B(n24251), .X(n24249) );
  nand_x4_sg U51183 ( .A(n24258), .B(n24259), .X(n24257) );
  nand_x4_sg U51184 ( .A(n24265), .B(n24266), .X(n24264) );
  nand_x4_sg U51185 ( .A(n24272), .B(n24273), .X(n24271) );
  nand_x4_sg U51186 ( .A(n24279), .B(n24280), .X(n24278) );
  nand_x4_sg U51187 ( .A(n24286), .B(n24287), .X(n24285) );
  nor_x1_sg U51188 ( .A(n24293), .B(n24294), .X(n24292) );
  nor_x1_sg U51189 ( .A(n24300), .B(n24301), .X(n24299) );
  nand_x4_sg U51190 ( .A(n24307), .B(n24308), .X(n24306) );
  nor_x1_sg U51191 ( .A(n24314), .B(n24315), .X(n24313) );
  nand_x4_sg U51192 ( .A(n24321), .B(n24322), .X(n24320) );
  nor_x1_sg U51193 ( .A(n24328), .B(n24329), .X(n24327) );
  nand_x4_sg U51194 ( .A(n24335), .B(n24336), .X(n24334) );
  nor_x1_sg U51195 ( .A(n24342), .B(n24343), .X(n24341) );
  nand_x4_sg U51196 ( .A(n24349), .B(n24350), .X(n24348) );
  nand_x1_sg U51197 ( .A(n39658), .B(n24356), .X(n24355) );
  nor_x1_sg U51198 ( .A(n24368), .B(n24369), .X(n24367) );
  nand_x4_sg U51199 ( .A(n24529), .B(n24530), .X(n24528) );
  nand_x4_sg U51200 ( .A(n24537), .B(n24538), .X(n24536) );
  nand_x4_sg U51201 ( .A(n24544), .B(n24545), .X(n24543) );
  nand_x4_sg U51202 ( .A(n24551), .B(n24552), .X(n24550) );
  nand_x4_sg U51203 ( .A(n24558), .B(n24559), .X(n24557) );
  nand_x4_sg U51204 ( .A(n24565), .B(n24566), .X(n24564) );
  nor_x1_sg U51205 ( .A(n24572), .B(n24573), .X(n24571) );
  nor_x1_sg U51206 ( .A(n24579), .B(n24580), .X(n24578) );
  nand_x4_sg U51207 ( .A(n24586), .B(n24587), .X(n24585) );
  nor_x1_sg U51208 ( .A(n24593), .B(n24594), .X(n24592) );
  nand_x4_sg U51209 ( .A(n24600), .B(n24601), .X(n24599) );
  nor_x1_sg U51210 ( .A(n24607), .B(n24608), .X(n24606) );
  nand_x4_sg U51211 ( .A(n24614), .B(n24615), .X(n24613) );
  nor_x1_sg U51212 ( .A(n24621), .B(n24622), .X(n24620) );
  nand_x4_sg U51213 ( .A(n24628), .B(n24629), .X(n24627) );
  nand_x1_sg U51214 ( .A(n41308), .B(n24635), .X(n24634) );
  nand_x1_sg U51215 ( .A(n24640), .B(n41308), .X(n24639) );
  nor_x1_sg U51216 ( .A(n24647), .B(n24648), .X(n24646) );
  nand_x4_sg U51217 ( .A(n24807), .B(n24808), .X(n24806) );
  nand_x4_sg U51218 ( .A(n24815), .B(n24816), .X(n24814) );
  nand_x4_sg U51219 ( .A(n24822), .B(n24823), .X(n24821) );
  nand_x4_sg U51220 ( .A(n24829), .B(n24830), .X(n24828) );
  nand_x4_sg U51221 ( .A(n24836), .B(n24837), .X(n24835) );
  nand_x4_sg U51222 ( .A(n24843), .B(n24844), .X(n24842) );
  nor_x1_sg U51223 ( .A(n24850), .B(n24851), .X(n24849) );
  nor_x1_sg U51224 ( .A(n24857), .B(n24858), .X(n24856) );
  nand_x4_sg U51225 ( .A(n24864), .B(n24865), .X(n24863) );
  nor_x1_sg U51226 ( .A(n24871), .B(n24872), .X(n24870) );
  nand_x4_sg U51227 ( .A(n24878), .B(n24879), .X(n24877) );
  nor_x1_sg U51228 ( .A(n24885), .B(n24886), .X(n24884) );
  nand_x4_sg U51229 ( .A(n24892), .B(n24893), .X(n24891) );
  nor_x1_sg U51230 ( .A(n24899), .B(n24900), .X(n24898) );
  nand_x4_sg U51231 ( .A(n24906), .B(n24907), .X(n24905) );
  nand_x1_sg U51232 ( .A(n39658), .B(n24913), .X(n24912) );
  nor_x1_sg U51233 ( .A(n24925), .B(n24926), .X(n24924) );
  nand_x4_sg U51234 ( .A(n25086), .B(n25087), .X(n25085) );
  nand_x4_sg U51235 ( .A(n25094), .B(n25095), .X(n25093) );
  nand_x4_sg U51236 ( .A(n25101), .B(n25102), .X(n25100) );
  nand_x4_sg U51237 ( .A(n25108), .B(n25109), .X(n25107) );
  nand_x4_sg U51238 ( .A(n25115), .B(n25116), .X(n25114) );
  nand_x4_sg U51239 ( .A(n25122), .B(n25123), .X(n25121) );
  nor_x1_sg U51240 ( .A(n25129), .B(n25130), .X(n25128) );
  nor_x1_sg U51241 ( .A(n25136), .B(n25137), .X(n25135) );
  nand_x4_sg U51242 ( .A(n25143), .B(n25144), .X(n25142) );
  nor_x1_sg U51243 ( .A(n25150), .B(n25151), .X(n25149) );
  nand_x4_sg U51244 ( .A(n25157), .B(n25158), .X(n25156) );
  nor_x1_sg U51245 ( .A(n25164), .B(n25165), .X(n25163) );
  nand_x4_sg U51246 ( .A(n25171), .B(n25172), .X(n25170) );
  nor_x1_sg U51247 ( .A(n25178), .B(n25179), .X(n25177) );
  nand_x4_sg U51248 ( .A(n25185), .B(n25186), .X(n25184) );
  nand_x1_sg U51249 ( .A(n39929), .B(n25192), .X(n25191) );
  nand_x1_sg U51250 ( .A(n25197), .B(n41309), .X(n25196) );
  nor_x1_sg U51251 ( .A(n25204), .B(n25205), .X(n25203) );
  nand_x4_sg U51252 ( .A(n25365), .B(n25366), .X(n25364) );
  nand_x4_sg U51253 ( .A(n25373), .B(n25374), .X(n25372) );
  nand_x4_sg U51254 ( .A(n25380), .B(n25381), .X(n25379) );
  nand_x4_sg U51255 ( .A(n25387), .B(n25388), .X(n25386) );
  nand_x4_sg U51256 ( .A(n25394), .B(n25395), .X(n25393) );
  nand_x4_sg U51257 ( .A(n25401), .B(n25402), .X(n25400) );
  nor_x1_sg U51258 ( .A(n25408), .B(n25409), .X(n25407) );
  nor_x1_sg U51259 ( .A(n25415), .B(n25416), .X(n25414) );
  nand_x4_sg U51260 ( .A(n25422), .B(n25423), .X(n25421) );
  nor_x1_sg U51261 ( .A(n25429), .B(n25430), .X(n25428) );
  nand_x4_sg U51262 ( .A(n25436), .B(n25437), .X(n25435) );
  nor_x1_sg U51263 ( .A(n25443), .B(n25444), .X(n25442) );
  nand_x4_sg U51264 ( .A(n25450), .B(n25451), .X(n25449) );
  nor_x1_sg U51265 ( .A(n25457), .B(n25458), .X(n25456) );
  nand_x4_sg U51266 ( .A(n25464), .B(n25465), .X(n25463) );
  nand_x1_sg U51267 ( .A(n38943), .B(n25471), .X(n25470) );
  nor_x1_sg U51268 ( .A(n25483), .B(n25484), .X(n25482) );
  nand_x4_sg U51269 ( .A(n25644), .B(n25645), .X(n25643) );
  nand_x4_sg U51270 ( .A(n25652), .B(n25653), .X(n25651) );
  nand_x4_sg U51271 ( .A(n25659), .B(n25660), .X(n25658) );
  nand_x4_sg U51272 ( .A(n25666), .B(n25667), .X(n25665) );
  nand_x4_sg U51273 ( .A(n25673), .B(n25674), .X(n25672) );
  nand_x4_sg U51274 ( .A(n25680), .B(n25681), .X(n25679) );
  nor_x1_sg U51275 ( .A(n25687), .B(n25688), .X(n25686) );
  nor_x1_sg U51276 ( .A(n25694), .B(n25695), .X(n25693) );
  nand_x4_sg U51277 ( .A(n25701), .B(n25702), .X(n25700) );
  nor_x1_sg U51278 ( .A(n25708), .B(n25709), .X(n25707) );
  nand_x4_sg U51279 ( .A(n25715), .B(n25716), .X(n25714) );
  nor_x1_sg U51280 ( .A(n25722), .B(n25723), .X(n25721) );
  nand_x4_sg U51281 ( .A(n25729), .B(n25730), .X(n25728) );
  nor_x1_sg U51282 ( .A(n25736), .B(n25737), .X(n25735) );
  nand_x4_sg U51283 ( .A(n25743), .B(n25744), .X(n25742) );
  nand_x1_sg U51284 ( .A(n40218), .B(n25750), .X(n25749) );
  nand_x1_sg U51285 ( .A(n25755), .B(n39658), .X(n25754) );
  nor_x1_sg U51286 ( .A(n25762), .B(n25763), .X(n25761) );
  nand_x2_sg U51287 ( .A(n25918), .B(n25919), .X(n5753) );
  nand_x2_sg U51288 ( .A(n25925), .B(n25926), .X(n5760) );
  nand_x2_sg U51289 ( .A(n25931), .B(n25932), .X(n5734) );
  nand_x2_sg U51290 ( .A(n25937), .B(n25938), .X(n5738) );
  nand_x2_sg U51291 ( .A(n25943), .B(n25944), .X(n5749) );
  nand_x2_sg U51292 ( .A(n25949), .B(n25950), .X(n5736) );
  nor_x1_sg U51293 ( .A(n25956), .B(n25957), .X(n5755) );
  nor_x1_sg U51294 ( .A(n25963), .B(n25964), .X(n5739) );
  nand_x2_sg U51295 ( .A(n25969), .B(n25970), .X(n5741) );
  nand_x1_sg U51296 ( .A(n25981), .B(n38943), .X(n25976) );
  nand_x2_sg U51297 ( .A(n25982), .B(n25983), .X(n5768) );
  nor_x1_sg U51298 ( .A(n51312), .B(n25989), .X(n5754) );
  nand_x2_sg U51299 ( .A(n25995), .B(n25996), .X(n5757) );
  nor_x1_sg U51300 ( .A(n51313), .B(n26002), .X(n5742) );
  nand_x2_sg U51301 ( .A(n26008), .B(n26009), .X(n5751) );
  nand_x1_sg U51302 ( .A(n41312), .B(n26014), .X(n5764) );
  nand_x1_sg U51303 ( .A(n26018), .B(n41318), .X(n5762) );
  nand_x2_sg U51304 ( .A(n26025), .B(n26026), .X(n5766) );
  nand_x2_sg U51305 ( .A(n26185), .B(n26186), .X(n26182) );
  nand_x2_sg U51306 ( .A(n26194), .B(n26195), .X(n26192) );
  nand_x2_sg U51307 ( .A(n26202), .B(n26203), .X(n26200) );
  nand_x2_sg U51308 ( .A(n26210), .B(n26211), .X(n26208) );
  nand_x2_sg U51309 ( .A(n26218), .B(n26219), .X(n26216) );
  nand_x2_sg U51310 ( .A(n26226), .B(n26227), .X(n26224) );
  nor_x1_sg U51311 ( .A(n26234), .B(n26235), .X(n26233) );
  nor_x1_sg U51312 ( .A(n26242), .B(n26243), .X(n26241) );
  nand_x2_sg U51313 ( .A(n26250), .B(n26251), .X(n26248) );
  nor_x1_sg U51314 ( .A(n26258), .B(n26259), .X(n26257) );
  nand_x2_sg U51315 ( .A(n26266), .B(n26267), .X(n26264) );
  nor_x1_sg U51316 ( .A(n26274), .B(n26275), .X(n26273) );
  nand_x2_sg U51317 ( .A(n26282), .B(n26283), .X(n26280) );
  nor_x1_sg U51318 ( .A(n26290), .B(n26291), .X(n26289) );
  nand_x2_sg U51319 ( .A(n26298), .B(n26299), .X(n26296) );
  nand_x1_sg U51320 ( .A(n39276), .B(n26306), .X(n26304) );
  inv_x1_sg U51321 ( .A(n26325), .X(n51412) );
  nand_x4_sg U51322 ( .A(n26481), .B(n26482), .X(n26480) );
  nand_x4_sg U51323 ( .A(n26489), .B(n26490), .X(n26488) );
  nand_x4_sg U51324 ( .A(n26496), .B(n26497), .X(n26495) );
  nand_x4_sg U51325 ( .A(n26503), .B(n26504), .X(n26502) );
  nand_x4_sg U51326 ( .A(n26510), .B(n26511), .X(n26509) );
  nand_x4_sg U51327 ( .A(n26517), .B(n26518), .X(n26516) );
  nor_x1_sg U51328 ( .A(n26524), .B(n26525), .X(n26523) );
  nor_x1_sg U51329 ( .A(n26531), .B(n26532), .X(n26530) );
  nand_x4_sg U51330 ( .A(n26538), .B(n26539), .X(n26537) );
  nor_x1_sg U51331 ( .A(n26545), .B(n26546), .X(n26544) );
  nand_x4_sg U51332 ( .A(n26552), .B(n26553), .X(n26551) );
  nor_x1_sg U51333 ( .A(n26559), .B(n26560), .X(n26558) );
  nand_x4_sg U51334 ( .A(n26566), .B(n26567), .X(n26565) );
  nor_x1_sg U51335 ( .A(n26573), .B(n26574), .X(n26572) );
  nand_x4_sg U51336 ( .A(n26580), .B(n26581), .X(n26579) );
  nand_x1_sg U51337 ( .A(n41312), .B(n26587), .X(n26586) );
  nand_x1_sg U51338 ( .A(n26592), .B(n41309), .X(n26591) );
  nor_x1_sg U51339 ( .A(n26599), .B(n26600), .X(n26598) );
  nand_x1_sg U51340 ( .A(out_L1[1]), .B(n41268), .X(n36879) );
  nand_x1_sg U51341 ( .A(out_L1[16]), .B(n41268), .X(n36887) );
  inv_x1_sg U51342 ( .A(n17470), .X(n51421) );
  nor_x1_sg U51343 ( .A(n5936), .B(n5937), .X(n5935) );
  nor_x1_sg U51344 ( .A(n5892), .B(n5893), .X(n5891) );
  nor_x1_sg U51345 ( .A(n5915), .B(n5916), .X(n5914) );
  nor_x1_sg U51346 ( .A(n5780), .B(n5781), .X(n5778) );
  nor_x1_sg U51347 ( .A(n5851), .B(n5852), .X(n5850) );
  nor_x1_sg U51348 ( .A(n5844), .B(n5845), .X(n5843) );
  nor_x1_sg U51349 ( .A(n5906), .B(n5907), .X(n5905) );
  nor_x1_sg U51350 ( .A(n5867), .B(n5868), .X(n5866) );
  nor_x1_sg U51351 ( .A(n5885), .B(n5886), .X(n5884) );
  nor_x1_sg U51352 ( .A(n5790), .B(n5791), .X(n5789) );
  nor_x1_sg U51353 ( .A(n5813), .B(n5814), .X(n5812) );
  nor_x1_sg U51354 ( .A(n5922), .B(n5923), .X(n5921) );
  nor_x1_sg U51355 ( .A(n5806), .B(n5807), .X(n5805) );
  nor_x1_sg U51356 ( .A(n5876), .B(n5877), .X(n5875) );
  nor_x1_sg U51357 ( .A(n5835), .B(n5836), .X(n5834) );
  nor_x1_sg U51358 ( .A(n5799), .B(n5800), .X(n5798) );
  nor_x1_sg U51359 ( .A(n5820), .B(n5821), .X(n5819) );
  nor_x1_sg U51360 ( .A(n5899), .B(n5900), .X(n5898) );
  nor_x1_sg U51361 ( .A(n5943), .B(n5944), .X(n5942) );
  nor_x1_sg U51362 ( .A(n5929), .B(n5930), .X(n5928) );
  nand_x1_sg U51363 ( .A(n39126), .B(n5865), .X(n5864) );
  nand_x1_sg U51364 ( .A(n41280), .B(n5797), .X(n5796) );
  inv_x1_sg U51365 ( .A(n22983), .X(n51489) );
  inv_x1_sg U51366 ( .A(n23260), .X(n51442) );
  inv_x1_sg U51367 ( .A(n23540), .X(n51443) );
  inv_x1_sg U51368 ( .A(n23819), .X(n51444) );
  inv_x1_sg U51369 ( .A(n24098), .X(n51445) );
  inv_x1_sg U51370 ( .A(n24377), .X(n51446) );
  inv_x1_sg U51371 ( .A(n24656), .X(n51447) );
  inv_x1_sg U51372 ( .A(n24934), .X(n51448) );
  inv_x1_sg U51373 ( .A(n25213), .X(n51449) );
  inv_x1_sg U51374 ( .A(n25492), .X(n51450) );
  inv_x1_sg U51375 ( .A(n25771), .X(n51451) );
  inv_x1_sg U51376 ( .A(n26608), .X(n51488) );
  nand_x1_sg U51377 ( .A(n39259), .B(n22187), .X(n22186) );
  nand_x1_sg U51378 ( .A(n41093), .B(n22046), .X(n22045) );
  nand_x1_sg U51379 ( .A(n39260), .B(n22162), .X(n22161) );
  nand_x1_sg U51380 ( .A(n38928), .B(n22021), .X(n22020) );
  nand_x1_sg U51381 ( .A(n36878), .B(n36879), .X(out[1]) );
  nor_x1_sg U51382 ( .A(n46602), .B(n19731), .X(n5965) );
  nand_x1_sg U51383 ( .A(n36886), .B(n36887), .X(out[16]) );
  inv_x1_sg U51384 ( .A(n25975), .X(n51467) );
  nor_x1_sg U51385 ( .A(n44973), .B(n27190), .X(n22575) );
  nor_x1_sg U51386 ( .A(n44966), .B(n28461), .X(n22594) );
  nor_x1_sg U51387 ( .A(n27968), .B(n27969), .X(n22565) );
  nor_x1_sg U51388 ( .A(n46598), .B(n19737), .X(n5969) );
  nor_x1_sg U51389 ( .A(n19931), .B(n19932), .X(n6023) );
  nand_x1_sg U51390 ( .A(n40026), .B(n6057), .X(n6058) );
  nor_x1_sg U51391 ( .A(n44971), .B(n27615), .X(n22569) );
  nor_x1_sg U51392 ( .A(n46600), .B(n19734), .X(n5964) );
  nor_x1_sg U51393 ( .A(n19743), .B(n19744), .X(n6003) );
  nor_x1_sg U51394 ( .A(n20432), .B(n20433), .X(n6210) );
  nor_x1_sg U51395 ( .A(n21174), .B(n21175), .X(n5998) );
  nor_x1_sg U51396 ( .A(n46563), .B(n19925), .X(n42330) );
  inv_x1_sg U51397 ( .A(n19927), .X(n46563) );
  nor_x1_sg U51398 ( .A(n19897), .B(n46382), .X(n6207) );
  nor_x1_sg U51399 ( .A(n46514), .B(n20125), .X(n42331) );
  inv_x1_sg U51400 ( .A(n20127), .X(n46514) );
  nor_x1_sg U51401 ( .A(n21278), .B(n21279), .X(n6635) );
  nor_x1_sg U51402 ( .A(n21283), .B(n21284), .X(n6590) );
  nor_x1_sg U51403 ( .A(n21288), .B(n21289), .X(n6546) );
  nor_x1_sg U51404 ( .A(n21293), .B(n21294), .X(n6501) );
  nor_x1_sg U51405 ( .A(n21298), .B(n21299), .X(n6457) );
  nor_x1_sg U51406 ( .A(n21303), .B(n21304), .X(n6412) );
  nor_x1_sg U51407 ( .A(n21308), .B(n21309), .X(n6368) );
  nor_x1_sg U51408 ( .A(n21313), .B(n21314), .X(n6323) );
  nor_x1_sg U51409 ( .A(n21318), .B(n21319), .X(n6279) );
  nor_x1_sg U51410 ( .A(n21323), .B(n21324), .X(n6234) );
  nor_x1_sg U51411 ( .A(n21328), .B(n21329), .X(n6188) );
  nor_x1_sg U51412 ( .A(n21333), .B(n21334), .X(n6142) );
  nor_x1_sg U51413 ( .A(n21338), .B(n21339), .X(n6096) );
  nor_x1_sg U51414 ( .A(n24937), .B(n51138), .X(n19126) );
  nand_x1_sg U51415 ( .A(n39259), .B(n22517), .X(n22516) );
  nand_x1_sg U51416 ( .A(n20962), .B(n22330), .X(n22329) );
  nand_x1_sg U51417 ( .A(n38930), .B(n22140), .X(n22139) );
  nor_x1_sg U51418 ( .A(n42058), .B(n42020), .X(n20962) );
  nand_x1_sg U51419 ( .A(n41090), .B(n22492), .X(n22491) );
  nand_x1_sg U51420 ( .A(n38928), .B(n22304), .X(n22303) );
  nand_x1_sg U51421 ( .A(n39260), .B(n22114), .X(n22113) );
  nor_x1_sg U51422 ( .A(n25216), .B(n51139), .X(n19118) );
  nor_x1_sg U51423 ( .A(n22707), .B(n47130), .X(n22638) );
  inv_x1_sg U51424 ( .A(n22708), .X(n47130) );
  inv_x1_sg U51425 ( .A(n41085), .X(n42332) );
  inv_x1_sg U51426 ( .A(n26305), .X(n51485) );
  inv_x1_sg U51427 ( .A(n5949), .X(n51526) );
  nor_x1_sg U51428 ( .A(n46521), .B(n19317), .X(n6077) );
  nor_x1_sg U51429 ( .A(n19716), .B(n19717), .X(n6087) );
  nor_x1_sg U51430 ( .A(n46608), .B(n19329), .X(n5974) );
  nor_x1_sg U51431 ( .A(n20110), .B(n20111), .X(n6161) );
  nor_x1_sg U51432 ( .A(n46596), .B(n19740), .X(n5968) );
  nor_x1_sg U51433 ( .A(n20034), .B(n20035), .X(n6655) );
  nor_x1_sg U51434 ( .A(n46431), .B(n19482), .X(n42333) );
  inv_x1_sg U51435 ( .A(n19484), .X(n46431) );
  nor_x1_sg U51436 ( .A(n19857), .B(n19858), .X(n6567) );
  nor_x1_sg U51437 ( .A(n19862), .B(n19863), .X(n6522) );
  nor_x1_sg U51438 ( .A(n19867), .B(n19868), .X(n6478) );
  nor_x1_sg U51439 ( .A(n19872), .B(n19873), .X(n6433) );
  nor_x1_sg U51440 ( .A(n19877), .B(n19878), .X(n6389) );
  nor_x1_sg U51441 ( .A(n19882), .B(n19883), .X(n6344) );
  nor_x1_sg U51442 ( .A(n19852), .B(n19853), .X(n6611) );
  nor_x1_sg U51443 ( .A(n19887), .B(n19888), .X(n6300) );
  nor_x1_sg U51444 ( .A(n21165), .B(n21166), .X(n6055) );
  nor_x1_sg U51445 ( .A(n46604), .B(n19728), .X(n42334) );
  inv_x1_sg U51446 ( .A(n19730), .X(n46604) );
  nor_x1_sg U51447 ( .A(n19892), .B(n19893), .X(n6255) );
  nor_x1_sg U51448 ( .A(n20296), .B(n20297), .X(n6118) );
  nor_x1_sg U51449 ( .A(n20674), .B(n20675), .X(n6687) );
  nor_x1_sg U51450 ( .A(n46591), .B(n20781), .X(n42335) );
  inv_x1_sg U51451 ( .A(n20783), .X(n46591) );
  nor_x1_sg U51452 ( .A(n20519), .B(n20520), .X(n6552) );
  nor_x1_sg U51453 ( .A(n20534), .B(n20535), .X(n6418) );
  nor_x1_sg U51454 ( .A(n20549), .B(n20550), .X(n6285) );
  nor_x1_sg U51455 ( .A(n46561), .B(n19928), .X(n6024) );
  nor_x1_sg U51456 ( .A(n46380), .B(n20281), .X(n6211) );
  nor_x1_sg U51457 ( .A(n46512), .B(n20128), .X(n6071) );
  nor_x1_sg U51458 ( .A(n26087), .B(n50325), .X(n42337) );
  inv_x1_sg U51459 ( .A(n26088), .X(n50325) );
  nand_x1_sg U51460 ( .A(n42059), .B(n17464), .X(n42338) );
  nand_x1_sg U51461 ( .A(n39434), .B(n41197), .X(n10095) );
  inv_x1_sg U51462 ( .A(n6784), .X(n51440) );
  inv_x1_sg U51463 ( .A(n6733), .X(n51439) );
  inv_x1_sg U51464 ( .A(n6693), .X(n51438) );
  inv_x1_sg U51465 ( .A(n6645), .X(n51437) );
  inv_x1_sg U51466 ( .A(n6600), .X(n51436) );
  inv_x1_sg U51467 ( .A(n6556), .X(n51435) );
  inv_x1_sg U51468 ( .A(n6511), .X(n51434) );
  inv_x1_sg U51469 ( .A(n6467), .X(n51433) );
  inv_x1_sg U51470 ( .A(n6422), .X(n51432) );
  inv_x1_sg U51471 ( .A(n6378), .X(n51431) );
  inv_x1_sg U51472 ( .A(n6333), .X(n51430) );
  inv_x1_sg U51473 ( .A(n6289), .X(n51429) );
  inv_x1_sg U51474 ( .A(n6244), .X(n51428) );
  inv_x1_sg U51475 ( .A(n6197), .X(n51427) );
  inv_x1_sg U51476 ( .A(n6151), .X(n51426) );
  inv_x1_sg U51477 ( .A(n6106), .X(n51425) );
  inv_x1_sg U51478 ( .A(n6058), .X(n51424) );
  inv_x1_sg U51479 ( .A(n6009), .X(n51423) );
  inv_x1_sg U51480 ( .A(n5953), .X(n51422) );
  inv_x1_sg U51481 ( .A(n19107), .X(n51441) );
  nor_x1_sg U51482 ( .A(n45079), .B(n28268), .X(n42340) );
  inv_x1_sg U51483 ( .A(n28270), .X(n45079) );
  nor_x1_sg U51484 ( .A(n46520), .B(n19495), .X(n42341) );
  inv_x1_sg U51485 ( .A(n19497), .X(n46520) );
  nor_x1_sg U51486 ( .A(n46605), .B(n19332), .X(n42342) );
  inv_x1_sg U51487 ( .A(n19334), .X(n46605) );
  nor_x1_sg U51488 ( .A(n45920), .B(n21444), .X(n42343) );
  inv_x1_sg U51489 ( .A(n21447), .X(n45920) );
  nor_x1_sg U51490 ( .A(n20509), .B(n20510), .X(n6641) );
  nor_x1_sg U51491 ( .A(n20544), .B(n20545), .X(n6329) );
  nor_x1_sg U51492 ( .A(n46432), .B(n19306), .X(n6169) );
  nor_x1_sg U51493 ( .A(n22794), .B(n46892), .X(n42369) );
  inv_x1_sg U51494 ( .A(n22795), .X(n46892) );
  nor_x1_sg U51495 ( .A(n26141), .B(n50559), .X(n42370) );
  inv_x1_sg U51496 ( .A(n26142), .X(n50559) );
  nand_x1_sg U51497 ( .A(n42119), .B(n39391), .X(n42386) );
  nand_x1_sg U51498 ( .A(n39434), .B(n41261), .X(n18287) );
  nand_x1_sg U51499 ( .A(n41418), .B(n41291), .X(n15828) );
  nand_x1_sg U51500 ( .A(n41417), .B(n41232), .X(n15009) );
  nand_x1_sg U51501 ( .A(n38983), .B(n41228), .X(n14190) );
  nand_x1_sg U51502 ( .A(n40220), .B(n41241), .X(n13371) );
  nand_x1_sg U51503 ( .A(n40090), .B(n41257), .X(n12552) );
  nand_x1_sg U51504 ( .A(n40089), .B(n41203), .X(n11733) );
  nand_x1_sg U51505 ( .A(n39435), .B(n41222), .X(n10914) );
  nand_x1_sg U51506 ( .A(n41417), .B(n39095), .X(n16646) );
  nand_x1_sg U51507 ( .A(n41417), .B(n40023), .X(n6822) );
  nand_x1_sg U51508 ( .A(n7345), .B(n47040), .X(n7316) );
  nand_x1_sg U51509 ( .A(n8163), .B(n47327), .X(n8134) );
  nand_x1_sg U51510 ( .A(n8981), .B(n47612), .X(n8952) );
  nand_x1_sg U51511 ( .A(n9801), .B(n47897), .X(n9772) );
  nand_x1_sg U51512 ( .A(n10620), .B(n48182), .X(n10591) );
  nand_x1_sg U51513 ( .A(n11439), .B(n48467), .X(n11410) );
  nand_x1_sg U51514 ( .A(n12258), .B(n48752), .X(n12229) );
  nand_x1_sg U51515 ( .A(n13077), .B(n49038), .X(n13048) );
  nand_x1_sg U51516 ( .A(n13896), .B(n49325), .X(n13867) );
  nand_x1_sg U51517 ( .A(n14715), .B(n49611), .X(n14686) );
  nand_x1_sg U51518 ( .A(n15534), .B(n49897), .X(n15505) );
  nand_x1_sg U51519 ( .A(n16353), .B(n50183), .X(n16324) );
  nand_x1_sg U51520 ( .A(n17170), .B(n50468), .X(n17141) );
  nand_x1_sg U51521 ( .A(n17991), .B(n50757), .X(n17962) );
  nand_x1_sg U51522 ( .A(n18812), .B(n51044), .X(n18783) );
  nand_x1_sg U51523 ( .A(n16705), .B(n50384), .X(n16703) );
  nand_x1_sg U51524 ( .A(n47109), .B(n7016), .X(n6979) );
  nand_x1_sg U51525 ( .A(n47395), .B(n7834), .X(n7796) );
  nand_x1_sg U51526 ( .A(n47680), .B(n8652), .X(n8614) );
  nand_x1_sg U51527 ( .A(n47965), .B(n9472), .X(n9434) );
  nand_x1_sg U51528 ( .A(n48250), .B(n10291), .X(n10253) );
  nand_x1_sg U51529 ( .A(n48535), .B(n11110), .X(n11072) );
  nand_x1_sg U51530 ( .A(n48820), .B(n11929), .X(n11891) );
  nand_x1_sg U51531 ( .A(n49107), .B(n12748), .X(n12710) );
  nand_x1_sg U51532 ( .A(n49393), .B(n13567), .X(n13529) );
  nand_x1_sg U51533 ( .A(n49679), .B(n14386), .X(n14348) );
  nand_x1_sg U51534 ( .A(n49965), .B(n15205), .X(n15167) );
  nand_x1_sg U51535 ( .A(n50251), .B(n16024), .X(n15986) );
  nand_x1_sg U51536 ( .A(n50825), .B(n17662), .X(n17624) );
  nand_x1_sg U51537 ( .A(n51112), .B(n18483), .X(n18445) );
  nand_x1_sg U51538 ( .A(n17131), .B(n50427), .X(n17117) );
  nand_x1_sg U51539 ( .A(n17084), .B(n50430), .X(n17062) );
  nand_x1_sg U51540 ( .A(n7259), .B(n47000), .X(n7237) );
  nand_x1_sg U51541 ( .A(n8078), .B(n47289), .X(n8056) );
  nand_x1_sg U51542 ( .A(n8896), .B(n47574), .X(n8874) );
  nand_x1_sg U51543 ( .A(n9716), .B(n47859), .X(n9694) );
  nand_x1_sg U51544 ( .A(n10535), .B(n48144), .X(n10513) );
  nand_x1_sg U51545 ( .A(n11354), .B(n48429), .X(n11332) );
  nand_x1_sg U51546 ( .A(n12173), .B(n48714), .X(n12151) );
  nand_x1_sg U51547 ( .A(n12992), .B(n49000), .X(n12970) );
  nand_x1_sg U51548 ( .A(n13811), .B(n49287), .X(n13789) );
  nand_x1_sg U51549 ( .A(n14630), .B(n49573), .X(n14608) );
  nand_x1_sg U51550 ( .A(n15449), .B(n49859), .X(n15427) );
  nand_x1_sg U51551 ( .A(n16268), .B(n50145), .X(n16246) );
  nand_x1_sg U51552 ( .A(n17906), .B(n50719), .X(n17884) );
  nand_x1_sg U51553 ( .A(n18727), .B(n51006), .X(n18705) );
  nand_x1_sg U51554 ( .A(n7117), .B(n46911), .X(n6872) );
  nand_x1_sg U51555 ( .A(n7935), .B(n47204), .X(n7689) );
  nand_x1_sg U51556 ( .A(n8753), .B(n47489), .X(n8507) );
  nand_x1_sg U51557 ( .A(n9573), .B(n47774), .X(n9327) );
  nand_x1_sg U51558 ( .A(n10392), .B(n48059), .X(n10146) );
  nand_x1_sg U51559 ( .A(n11211), .B(n48344), .X(n10965) );
  nand_x1_sg U51560 ( .A(n12030), .B(n48629), .X(n11784) );
  nand_x1_sg U51561 ( .A(n12849), .B(n48915), .X(n12603) );
  nand_x1_sg U51562 ( .A(n13668), .B(n49202), .X(n13422) );
  nand_x1_sg U51563 ( .A(n14487), .B(n49488), .X(n14241) );
  nand_x1_sg U51564 ( .A(n15306), .B(n49774), .X(n15060) );
  nand_x1_sg U51565 ( .A(n16125), .B(n50060), .X(n15879) );
  nand_x1_sg U51566 ( .A(n16942), .B(n50345), .X(n16696) );
  nand_x1_sg U51567 ( .A(n17763), .B(n50634), .X(n17517) );
  nand_x1_sg U51568 ( .A(n18584), .B(n50921), .X(n18338) );
  nand_x1_sg U51569 ( .A(n7588), .B(n47047), .X(n7579) );
  nand_x1_sg U51570 ( .A(n17413), .B(n50475), .X(n17404) );
  nand_x1_sg U51571 ( .A(n50295), .B(n16668), .X(n16666) );
  nand_x1_sg U51572 ( .A(n47155), .B(n7661), .X(n7659) );
  nand_x1_sg U51573 ( .A(n47440), .B(n8479), .X(n8477) );
  nand_x1_sg U51574 ( .A(n47725), .B(n9299), .X(n9297) );
  nand_x1_sg U51575 ( .A(n48010), .B(n10118), .X(n10116) );
  nand_x1_sg U51576 ( .A(n48295), .B(n10937), .X(n10935) );
  nand_x1_sg U51577 ( .A(n48580), .B(n11756), .X(n11754) );
  nand_x1_sg U51578 ( .A(n48866), .B(n12575), .X(n12573) );
  nand_x1_sg U51579 ( .A(n49153), .B(n13394), .X(n13392) );
  nand_x1_sg U51580 ( .A(n49439), .B(n14213), .X(n14211) );
  nand_x1_sg U51581 ( .A(n49724), .B(n15032), .X(n15030) );
  nand_x1_sg U51582 ( .A(n50011), .B(n15851), .X(n15849) );
  nand_x1_sg U51583 ( .A(n50585), .B(n17489), .X(n17487) );
  nand_x1_sg U51584 ( .A(n50872), .B(n18310), .X(n18308) );
  nand_x1_sg U51585 ( .A(n7175), .B(n46928), .X(n7170) );
  nand_x1_sg U51586 ( .A(n7994), .B(n47220), .X(n7989) );
  nand_x1_sg U51587 ( .A(n8812), .B(n47505), .X(n8807) );
  nand_x1_sg U51588 ( .A(n9632), .B(n47790), .X(n9627) );
  nand_x1_sg U51589 ( .A(n10451), .B(n48075), .X(n10446) );
  nand_x1_sg U51590 ( .A(n11270), .B(n48360), .X(n11265) );
  nand_x1_sg U51591 ( .A(n12089), .B(n48645), .X(n12084) );
  nand_x1_sg U51592 ( .A(n12908), .B(n48931), .X(n12903) );
  nand_x1_sg U51593 ( .A(n13727), .B(n49218), .X(n13722) );
  nand_x1_sg U51594 ( .A(n14546), .B(n49504), .X(n14541) );
  nand_x1_sg U51595 ( .A(n15365), .B(n49790), .X(n15360) );
  nand_x1_sg U51596 ( .A(n16184), .B(n50076), .X(n16179) );
  nand_x1_sg U51597 ( .A(n17822), .B(n50650), .X(n17817) );
  nand_x1_sg U51598 ( .A(n18643), .B(n50937), .X(n18638) );
  nand_x1_sg U51599 ( .A(n17000), .B(n50361), .X(n16995) );
  nand_x1_sg U51600 ( .A(n6881), .B(n46952), .X(n6879) );
  nand_x1_sg U51601 ( .A(n7698), .B(n47243), .X(n7696) );
  nand_x1_sg U51602 ( .A(n8516), .B(n47528), .X(n8514) );
  nand_x1_sg U51603 ( .A(n9336), .B(n47813), .X(n9334) );
  nand_x1_sg U51604 ( .A(n10155), .B(n48098), .X(n10153) );
  nand_x1_sg U51605 ( .A(n10974), .B(n48383), .X(n10972) );
  nand_x1_sg U51606 ( .A(n11793), .B(n48668), .X(n11791) );
  nand_x1_sg U51607 ( .A(n12612), .B(n48954), .X(n12610) );
  nand_x1_sg U51608 ( .A(n13431), .B(n49241), .X(n13429) );
  nand_x1_sg U51609 ( .A(n14250), .B(n49527), .X(n14248) );
  nand_x1_sg U51610 ( .A(n15069), .B(n49813), .X(n15067) );
  nand_x1_sg U51611 ( .A(n15888), .B(n50099), .X(n15886) );
  nand_x1_sg U51612 ( .A(n17526), .B(n50673), .X(n17524) );
  nand_x1_sg U51613 ( .A(n18347), .B(n50960), .X(n18345) );
  nand_x1_sg U51614 ( .A(n7553), .B(n47052), .X(n7520) );
  nand_x1_sg U51615 ( .A(n8371), .B(n47339), .X(n8338) );
  nand_x1_sg U51616 ( .A(n9189), .B(n47624), .X(n9156) );
  nand_x1_sg U51617 ( .A(n10009), .B(n47909), .X(n9976) );
  nand_x1_sg U51618 ( .A(n10828), .B(n48194), .X(n10795) );
  nand_x1_sg U51619 ( .A(n11647), .B(n48479), .X(n11614) );
  nand_x1_sg U51620 ( .A(n12466), .B(n48764), .X(n12433) );
  nand_x1_sg U51621 ( .A(n13285), .B(n49050), .X(n13252) );
  nand_x1_sg U51622 ( .A(n14104), .B(n49337), .X(n14071) );
  nand_x1_sg U51623 ( .A(n14923), .B(n49623), .X(n14890) );
  nand_x1_sg U51624 ( .A(n15742), .B(n49909), .X(n15709) );
  nand_x1_sg U51625 ( .A(n16561), .B(n50195), .X(n16528) );
  nand_x1_sg U51626 ( .A(n17378), .B(n50480), .X(n17345) );
  nand_x1_sg U51627 ( .A(n18199), .B(n50769), .X(n18166) );
  nand_x1_sg U51628 ( .A(n19020), .B(n51056), .X(n18987) );
  nand_x1_sg U51629 ( .A(n47077), .B(n6984), .X(n6982) );
  nand_x1_sg U51630 ( .A(n47363), .B(n7801), .X(n7799) );
  nand_x1_sg U51631 ( .A(n47648), .B(n8619), .X(n8617) );
  nand_x1_sg U51632 ( .A(n47933), .B(n9439), .X(n9437) );
  nand_x1_sg U51633 ( .A(n48218), .B(n10258), .X(n10256) );
  nand_x1_sg U51634 ( .A(n48503), .B(n11077), .X(n11075) );
  nand_x1_sg U51635 ( .A(n48788), .B(n11896), .X(n11894) );
  nand_x1_sg U51636 ( .A(n49075), .B(n12715), .X(n12713) );
  nand_x1_sg U51637 ( .A(n49361), .B(n13534), .X(n13532) );
  nand_x1_sg U51638 ( .A(n49647), .B(n14353), .X(n14351) );
  nand_x1_sg U51639 ( .A(n49933), .B(n15172), .X(n15170) );
  nand_x1_sg U51640 ( .A(n50219), .B(n15991), .X(n15989) );
  nand_x1_sg U51641 ( .A(n50504), .B(n16808), .X(n16806) );
  nand_x1_sg U51642 ( .A(n50793), .B(n17629), .X(n17627) );
  nand_x1_sg U51643 ( .A(n51080), .B(n18450), .X(n18448) );
  nand_x1_sg U51644 ( .A(n6863), .B(n46897), .X(n6861) );
  nand_x1_sg U51645 ( .A(n7680), .B(n47192), .X(n7678) );
  nand_x1_sg U51646 ( .A(n8498), .B(n47477), .X(n8496) );
  nand_x1_sg U51647 ( .A(n9318), .B(n47762), .X(n9316) );
  nand_x1_sg U51648 ( .A(n10137), .B(n48047), .X(n10135) );
  nand_x1_sg U51649 ( .A(n10956), .B(n48332), .X(n10954) );
  nand_x1_sg U51650 ( .A(n11775), .B(n48617), .X(n11773) );
  nand_x1_sg U51651 ( .A(n12594), .B(n48903), .X(n12592) );
  nand_x1_sg U51652 ( .A(n13413), .B(n49190), .X(n13411) );
  nand_x1_sg U51653 ( .A(n14232), .B(n49476), .X(n14230) );
  nand_x1_sg U51654 ( .A(n15051), .B(n49762), .X(n15049) );
  nand_x1_sg U51655 ( .A(n15870), .B(n50048), .X(n15868) );
  nand_x1_sg U51656 ( .A(n16687), .B(n50330), .X(n16685) );
  nand_x1_sg U51657 ( .A(n17508), .B(n50622), .X(n17506) );
  nand_x1_sg U51658 ( .A(n18329), .B(n50909), .X(n18327) );
  nand_x1_sg U51659 ( .A(n6869), .B(n46912), .X(n6867) );
  nand_x1_sg U51660 ( .A(n7686), .B(n47205), .X(n7684) );
  nand_x1_sg U51661 ( .A(n8504), .B(n47490), .X(n8502) );
  nand_x1_sg U51662 ( .A(n9324), .B(n47775), .X(n9322) );
  nand_x1_sg U51663 ( .A(n10143), .B(n48060), .X(n10141) );
  nand_x1_sg U51664 ( .A(n10962), .B(n48345), .X(n10960) );
  nand_x1_sg U51665 ( .A(n11781), .B(n48630), .X(n11779) );
  nand_x1_sg U51666 ( .A(n12600), .B(n48916), .X(n12598) );
  nand_x1_sg U51667 ( .A(n13419), .B(n49203), .X(n13417) );
  nand_x1_sg U51668 ( .A(n14238), .B(n49489), .X(n14236) );
  nand_x1_sg U51669 ( .A(n15057), .B(n49775), .X(n15055) );
  nand_x1_sg U51670 ( .A(n15876), .B(n50061), .X(n15874) );
  nand_x1_sg U51671 ( .A(n16693), .B(n50346), .X(n16691) );
  nand_x1_sg U51672 ( .A(n17514), .B(n50635), .X(n17512) );
  nand_x1_sg U51673 ( .A(n18335), .B(n50922), .X(n18333) );
  nand_x1_sg U51674 ( .A(n7238), .B(n46953), .X(n7234) );
  nand_x1_sg U51675 ( .A(n8057), .B(n47244), .X(n8053) );
  nand_x1_sg U51676 ( .A(n8875), .B(n47529), .X(n8871) );
  nand_x1_sg U51677 ( .A(n9695), .B(n47814), .X(n9691) );
  nand_x1_sg U51678 ( .A(n10514), .B(n48099), .X(n10510) );
  nand_x1_sg U51679 ( .A(n11333), .B(n48384), .X(n11329) );
  nand_x1_sg U51680 ( .A(n12152), .B(n48669), .X(n12148) );
  nand_x1_sg U51681 ( .A(n12971), .B(n48955), .X(n12967) );
  nand_x1_sg U51682 ( .A(n13790), .B(n49242), .X(n13786) );
  nand_x1_sg U51683 ( .A(n14609), .B(n49528), .X(n14605) );
  nand_x1_sg U51684 ( .A(n15428), .B(n49814), .X(n15424) );
  nand_x1_sg U51685 ( .A(n16247), .B(n50100), .X(n16243) );
  nand_x1_sg U51686 ( .A(n17063), .B(n50385), .X(n17059) );
  nand_x1_sg U51687 ( .A(n17885), .B(n50674), .X(n17881) );
  nand_x1_sg U51688 ( .A(n18706), .B(n50961), .X(n18702) );
  nand_x1_sg U51689 ( .A(n20592), .B(n46613), .X(n20590) );
  inv_x1_sg U51690 ( .A(n7406), .X(n47091) );
  inv_x1_sg U51691 ( .A(n7454), .X(n47115) );
  inv_x1_sg U51692 ( .A(n8224), .X(n47377) );
  inv_x1_sg U51693 ( .A(n8272), .X(n47401) );
  inv_x1_sg U51694 ( .A(n9042), .X(n47662) );
  inv_x1_sg U51695 ( .A(n9090), .X(n47686) );
  inv_x1_sg U51696 ( .A(n9862), .X(n47947) );
  inv_x1_sg U51697 ( .A(n9910), .X(n47971) );
  inv_x1_sg U51698 ( .A(n10681), .X(n48232) );
  inv_x1_sg U51699 ( .A(n10729), .X(n48256) );
  inv_x1_sg U51700 ( .A(n11500), .X(n48517) );
  inv_x1_sg U51701 ( .A(n11548), .X(n48541) );
  inv_x1_sg U51702 ( .A(n12319), .X(n48802) );
  inv_x1_sg U51703 ( .A(n12367), .X(n48826) );
  inv_x1_sg U51704 ( .A(n13138), .X(n49089) );
  inv_x1_sg U51705 ( .A(n13186), .X(n49113) );
  inv_x1_sg U51706 ( .A(n13957), .X(n49375) );
  inv_x1_sg U51707 ( .A(n14005), .X(n49399) );
  inv_x1_sg U51708 ( .A(n14776), .X(n49661) );
  inv_x1_sg U51709 ( .A(n14824), .X(n49685) );
  inv_x1_sg U51710 ( .A(n15595), .X(n49947) );
  inv_x1_sg U51711 ( .A(n15643), .X(n49971) );
  inv_x1_sg U51712 ( .A(n16414), .X(n50233) );
  inv_x1_sg U51713 ( .A(n16462), .X(n50257) );
  inv_x1_sg U51714 ( .A(n17231), .X(n50518) );
  inv_x1_sg U51715 ( .A(n17279), .X(n50542) );
  inv_x1_sg U51716 ( .A(n18052), .X(n50807) );
  inv_x1_sg U51717 ( .A(n18100), .X(n50831) );
  inv_x1_sg U51718 ( .A(n18873), .X(n51094) );
  inv_x1_sg U51719 ( .A(n18921), .X(n51118) );
  inv_x1_sg U51720 ( .A(n17207), .X(n50466) );
  inv_x1_sg U51721 ( .A(n7349), .X(n47069) );
  inv_x1_sg U51722 ( .A(n8167), .X(n47355) );
  inv_x1_sg U51723 ( .A(n8985), .X(n47640) );
  inv_x1_sg U51724 ( .A(n9805), .X(n47925) );
  inv_x1_sg U51725 ( .A(n10624), .X(n48210) );
  inv_x1_sg U51726 ( .A(n11443), .X(n48495) );
  inv_x1_sg U51727 ( .A(n12262), .X(n48780) );
  inv_x1_sg U51728 ( .A(n13081), .X(n49067) );
  inv_x1_sg U51729 ( .A(n13900), .X(n49353) );
  inv_x1_sg U51730 ( .A(n14719), .X(n49639) );
  inv_x1_sg U51731 ( .A(n15538), .X(n49925) );
  inv_x1_sg U51732 ( .A(n16357), .X(n50211) );
  inv_x1_sg U51733 ( .A(n17174), .X(n50496) );
  inv_x1_sg U51734 ( .A(n17995), .X(n50785) );
  inv_x1_sg U51735 ( .A(n18816), .X(n51072) );
  inv_x1_sg U51736 ( .A(n7382), .X(n47038) );
  inv_x1_sg U51737 ( .A(n8200), .X(n47325) );
  inv_x1_sg U51738 ( .A(n9018), .X(n47610) );
  inv_x1_sg U51739 ( .A(n9838), .X(n47895) );
  inv_x1_sg U51740 ( .A(n10657), .X(n48180) );
  inv_x1_sg U51741 ( .A(n11476), .X(n48465) );
  inv_x1_sg U51742 ( .A(n12295), .X(n48750) );
  inv_x1_sg U51743 ( .A(n13114), .X(n49036) );
  inv_x1_sg U51744 ( .A(n13933), .X(n49323) );
  inv_x1_sg U51745 ( .A(n14752), .X(n49609) );
  inv_x1_sg U51746 ( .A(n15571), .X(n49895) );
  inv_x1_sg U51747 ( .A(n16390), .X(n50181) );
  inv_x1_sg U51748 ( .A(n18028), .X(n50755) );
  inv_x1_sg U51749 ( .A(n18849), .X(n51042) );
  inv_x1_sg U51750 ( .A(n7346), .X(n47040) );
  inv_x1_sg U51751 ( .A(n8164), .X(n47327) );
  inv_x1_sg U51752 ( .A(n8982), .X(n47612) );
  inv_x1_sg U51753 ( .A(n9802), .X(n47897) );
  inv_x1_sg U51754 ( .A(n10621), .X(n48182) );
  inv_x1_sg U51755 ( .A(n11440), .X(n48467) );
  inv_x1_sg U51756 ( .A(n12259), .X(n48752) );
  inv_x1_sg U51757 ( .A(n13078), .X(n49038) );
  inv_x1_sg U51758 ( .A(n13897), .X(n49325) );
  inv_x1_sg U51759 ( .A(n14716), .X(n49611) );
  inv_x1_sg U51760 ( .A(n15535), .X(n49897) );
  inv_x1_sg U51761 ( .A(n16354), .X(n50183) );
  inv_x1_sg U51762 ( .A(n17171), .X(n50468) );
  inv_x1_sg U51763 ( .A(n17992), .X(n50757) );
  inv_x1_sg U51764 ( .A(n18813), .X(n51044) );
  inv_x1_sg U51765 ( .A(n7522), .X(n47085) );
  inv_x1_sg U51766 ( .A(n8340), .X(n47371) );
  inv_x1_sg U51767 ( .A(n9158), .X(n47656) );
  inv_x1_sg U51768 ( .A(n9978), .X(n47941) );
  inv_x1_sg U51769 ( .A(n10797), .X(n48226) );
  inv_x1_sg U51770 ( .A(n11616), .X(n48511) );
  inv_x1_sg U51771 ( .A(n12435), .X(n48796) );
  inv_x1_sg U51772 ( .A(n13254), .X(n49083) );
  inv_x1_sg U51773 ( .A(n14073), .X(n49369) );
  inv_x1_sg U51774 ( .A(n14892), .X(n49655) );
  inv_x1_sg U51775 ( .A(n15711), .X(n49941) );
  inv_x1_sg U51776 ( .A(n16530), .X(n50227) );
  inv_x1_sg U51777 ( .A(n17347), .X(n50512) );
  inv_x1_sg U51778 ( .A(n18168), .X(n50801) );
  inv_x1_sg U51779 ( .A(n18989), .X(n51088) );
  inv_x1_sg U51780 ( .A(n7314), .X(n47041) );
  inv_x1_sg U51781 ( .A(n17139), .X(n50469) );
  inv_x1_sg U51782 ( .A(n7542), .X(n47111) );
  inv_x1_sg U51783 ( .A(n8360), .X(n47397) );
  inv_x1_sg U51784 ( .A(n9178), .X(n47682) );
  inv_x1_sg U51785 ( .A(n9998), .X(n47967) );
  inv_x1_sg U51786 ( .A(n10817), .X(n48252) );
  inv_x1_sg U51787 ( .A(n11636), .X(n48537) );
  inv_x1_sg U51788 ( .A(n12455), .X(n48822) );
  inv_x1_sg U51789 ( .A(n13274), .X(n49109) );
  inv_x1_sg U51790 ( .A(n14093), .X(n49395) );
  inv_x1_sg U51791 ( .A(n14912), .X(n49681) );
  inv_x1_sg U51792 ( .A(n15731), .X(n49967) );
  inv_x1_sg U51793 ( .A(n16550), .X(n50253) );
  inv_x1_sg U51794 ( .A(n17367), .X(n50538) );
  inv_x1_sg U51795 ( .A(n18188), .X(n50827) );
  inv_x1_sg U51796 ( .A(n19009), .X(n51114) );
  inv_x1_sg U51797 ( .A(n7195), .X(n46949) );
  inv_x1_sg U51798 ( .A(n8014), .X(n47240) );
  inv_x1_sg U51799 ( .A(n8832), .X(n47525) );
  inv_x1_sg U51800 ( .A(n9652), .X(n47810) );
  inv_x1_sg U51801 ( .A(n10471), .X(n48095) );
  inv_x1_sg U51802 ( .A(n11290), .X(n48380) );
  inv_x1_sg U51803 ( .A(n12109), .X(n48665) );
  inv_x1_sg U51804 ( .A(n12928), .X(n48951) );
  inv_x1_sg U51805 ( .A(n13747), .X(n49238) );
  inv_x1_sg U51806 ( .A(n14566), .X(n49524) );
  inv_x1_sg U51807 ( .A(n15385), .X(n49810) );
  inv_x1_sg U51808 ( .A(n16204), .X(n50096) );
  inv_x1_sg U51809 ( .A(n17020), .X(n50381) );
  inv_x1_sg U51810 ( .A(n17842), .X(n50670) );
  inv_x1_sg U51811 ( .A(n18663), .X(n50957) );
  inv_x1_sg U51812 ( .A(n7482), .X(n47088) );
  inv_x1_sg U51813 ( .A(n8300), .X(n47374) );
  inv_x1_sg U51814 ( .A(n9118), .X(n47659) );
  inv_x1_sg U51815 ( .A(n9938), .X(n47944) );
  inv_x1_sg U51816 ( .A(n10757), .X(n48229) );
  inv_x1_sg U51817 ( .A(n11576), .X(n48514) );
  inv_x1_sg U51818 ( .A(n12395), .X(n48799) );
  inv_x1_sg U51819 ( .A(n13214), .X(n49086) );
  inv_x1_sg U51820 ( .A(n14033), .X(n49372) );
  inv_x1_sg U51821 ( .A(n14852), .X(n49658) );
  inv_x1_sg U51822 ( .A(n15671), .X(n49944) );
  inv_x1_sg U51823 ( .A(n16490), .X(n50230) );
  inv_x1_sg U51824 ( .A(n17307), .X(n50515) );
  inv_x1_sg U51825 ( .A(n18128), .X(n50804) );
  inv_x1_sg U51826 ( .A(n18949), .X(n51091) );
  inv_x1_sg U51827 ( .A(n7263), .X(n47015) );
  inv_x1_sg U51828 ( .A(n17088), .X(n50444) );
  inv_x1_sg U51829 ( .A(n16706), .X(n50384) );
  inv_x1_sg U51830 ( .A(n8047), .X(n47237) );
  inv_x1_sg U51831 ( .A(n8865), .X(n47522) );
  inv_x1_sg U51832 ( .A(n9685), .X(n47807) );
  inv_x1_sg U51833 ( .A(n10504), .X(n48092) );
  inv_x1_sg U51834 ( .A(n11323), .X(n48377) );
  inv_x1_sg U51835 ( .A(n12142), .X(n48662) );
  inv_x1_sg U51836 ( .A(n12961), .X(n48948) );
  inv_x1_sg U51837 ( .A(n13780), .X(n49235) );
  inv_x1_sg U51838 ( .A(n14599), .X(n49521) );
  inv_x1_sg U51839 ( .A(n15418), .X(n49807) );
  inv_x1_sg U51840 ( .A(n16237), .X(n50093) );
  inv_x1_sg U51841 ( .A(n17875), .X(n50667) );
  inv_x1_sg U51842 ( .A(n18696), .X(n50954) );
  inv_x1_sg U51843 ( .A(n7421), .X(n47019) );
  inv_x1_sg U51844 ( .A(n8239), .X(n47307) );
  inv_x1_sg U51845 ( .A(n9057), .X(n47592) );
  inv_x1_sg U51846 ( .A(n9877), .X(n47877) );
  inv_x1_sg U51847 ( .A(n10696), .X(n48162) );
  inv_x1_sg U51848 ( .A(n11515), .X(n48447) );
  inv_x1_sg U51849 ( .A(n12334), .X(n48732) );
  inv_x1_sg U51850 ( .A(n13153), .X(n49018) );
  inv_x1_sg U51851 ( .A(n13972), .X(n49305) );
  inv_x1_sg U51852 ( .A(n14791), .X(n49591) );
  inv_x1_sg U51853 ( .A(n15610), .X(n49877) );
  inv_x1_sg U51854 ( .A(n16429), .X(n50163) );
  inv_x1_sg U51855 ( .A(n18067), .X(n50737) );
  inv_x1_sg U51856 ( .A(n18888), .X(n51024) );
  inv_x1_sg U51857 ( .A(n17132), .X(n50427) );
  inv_x1_sg U51858 ( .A(n7260), .X(n47000) );
  inv_x1_sg U51859 ( .A(n17085), .X(n50430) );
  inv_x1_sg U51860 ( .A(n8079), .X(n47289) );
  inv_x1_sg U51861 ( .A(n8897), .X(n47574) );
  inv_x1_sg U51862 ( .A(n9717), .X(n47859) );
  inv_x1_sg U51863 ( .A(n10536), .X(n48144) );
  inv_x1_sg U51864 ( .A(n11355), .X(n48429) );
  inv_x1_sg U51865 ( .A(n12174), .X(n48714) );
  inv_x1_sg U51866 ( .A(n12993), .X(n49000) );
  inv_x1_sg U51867 ( .A(n13812), .X(n49287) );
  inv_x1_sg U51868 ( .A(n14631), .X(n49573) );
  inv_x1_sg U51869 ( .A(n15450), .X(n49859) );
  inv_x1_sg U51870 ( .A(n16269), .X(n50145) );
  inv_x1_sg U51871 ( .A(n17907), .X(n50719) );
  inv_x1_sg U51872 ( .A(n18728), .X(n51006) );
  inv_x1_sg U51873 ( .A(n7118), .X(n46911) );
  inv_x1_sg U51874 ( .A(n7936), .X(n47204) );
  inv_x1_sg U51875 ( .A(n8754), .X(n47489) );
  inv_x1_sg U51876 ( .A(n9574), .X(n47774) );
  inv_x1_sg U51877 ( .A(n10393), .X(n48059) );
  inv_x1_sg U51878 ( .A(n11212), .X(n48344) );
  inv_x1_sg U51879 ( .A(n12031), .X(n48629) );
  inv_x1_sg U51880 ( .A(n12850), .X(n48915) );
  inv_x1_sg U51881 ( .A(n13669), .X(n49202) );
  inv_x1_sg U51882 ( .A(n14488), .X(n49488) );
  inv_x1_sg U51883 ( .A(n15307), .X(n49774) );
  inv_x1_sg U51884 ( .A(n16126), .X(n50060) );
  inv_x1_sg U51885 ( .A(n16943), .X(n50345) );
  inv_x1_sg U51886 ( .A(n17764), .X(n50634) );
  inv_x1_sg U51887 ( .A(n18585), .X(n50921) );
  inv_x1_sg U51888 ( .A(n7515), .X(n47114) );
  inv_x1_sg U51889 ( .A(n8333), .X(n47400) );
  inv_x1_sg U51890 ( .A(n9151), .X(n47685) );
  inv_x1_sg U51891 ( .A(n9971), .X(n47970) );
  inv_x1_sg U51892 ( .A(n10790), .X(n48255) );
  inv_x1_sg U51893 ( .A(n11609), .X(n48540) );
  inv_x1_sg U51894 ( .A(n12428), .X(n48825) );
  inv_x1_sg U51895 ( .A(n13247), .X(n49112) );
  inv_x1_sg U51896 ( .A(n14066), .X(n49398) );
  inv_x1_sg U51897 ( .A(n14885), .X(n49684) );
  inv_x1_sg U51898 ( .A(n15704), .X(n49970) );
  inv_x1_sg U51899 ( .A(n16523), .X(n50256) );
  inv_x1_sg U51900 ( .A(n17340), .X(n50541) );
  inv_x1_sg U51901 ( .A(n18161), .X(n50830) );
  inv_x1_sg U51902 ( .A(n18982), .X(n51117) );
  inv_x1_sg U51903 ( .A(n7451), .X(n47090) );
  inv_x1_sg U51904 ( .A(n8269), .X(n47376) );
  inv_x1_sg U51905 ( .A(n9087), .X(n47661) );
  inv_x1_sg U51906 ( .A(n9907), .X(n47946) );
  inv_x1_sg U51907 ( .A(n10726), .X(n48231) );
  inv_x1_sg U51908 ( .A(n11545), .X(n48516) );
  inv_x1_sg U51909 ( .A(n12364), .X(n48801) );
  inv_x1_sg U51910 ( .A(n13183), .X(n49088) );
  inv_x1_sg U51911 ( .A(n14002), .X(n49374) );
  inv_x1_sg U51912 ( .A(n14821), .X(n49660) );
  inv_x1_sg U51913 ( .A(n15640), .X(n49946) );
  inv_x1_sg U51914 ( .A(n16459), .X(n50232) );
  inv_x1_sg U51915 ( .A(n17276), .X(n50517) );
  inv_x1_sg U51916 ( .A(n18097), .X(n50806) );
  inv_x1_sg U51917 ( .A(n18918), .X(n51093) );
  inv_x1_sg U51918 ( .A(n6934), .X(n47102) );
  inv_x1_sg U51919 ( .A(n7751), .X(n47388) );
  inv_x1_sg U51920 ( .A(n8569), .X(n47673) );
  inv_x1_sg U51921 ( .A(n9389), .X(n47958) );
  inv_x1_sg U51922 ( .A(n10208), .X(n48243) );
  inv_x1_sg U51923 ( .A(n11027), .X(n48528) );
  inv_x1_sg U51924 ( .A(n11846), .X(n48813) );
  inv_x1_sg U51925 ( .A(n12665), .X(n49100) );
  inv_x1_sg U51926 ( .A(n13484), .X(n49386) );
  inv_x1_sg U51927 ( .A(n14303), .X(n49672) );
  inv_x1_sg U51928 ( .A(n15122), .X(n49958) );
  inv_x1_sg U51929 ( .A(n15941), .X(n50244) );
  inv_x1_sg U51930 ( .A(n16758), .X(n50529) );
  inv_x1_sg U51931 ( .A(n17579), .X(n50818) );
  inv_x1_sg U51932 ( .A(n18400), .X(n51105) );
  inv_x1_sg U51933 ( .A(n7568), .X(n47110) );
  inv_x1_sg U51934 ( .A(n8386), .X(n47396) );
  inv_x1_sg U51935 ( .A(n9204), .X(n47681) );
  inv_x1_sg U51936 ( .A(n10024), .X(n47966) );
  inv_x1_sg U51937 ( .A(n10843), .X(n48251) );
  inv_x1_sg U51938 ( .A(n11662), .X(n48536) );
  inv_x1_sg U51939 ( .A(n12481), .X(n48821) );
  inv_x1_sg U51940 ( .A(n13300), .X(n49108) );
  inv_x1_sg U51941 ( .A(n14119), .X(n49394) );
  inv_x1_sg U51942 ( .A(n14938), .X(n49680) );
  inv_x1_sg U51943 ( .A(n15757), .X(n49966) );
  inv_x1_sg U51944 ( .A(n16576), .X(n50252) );
  inv_x1_sg U51945 ( .A(n17393), .X(n50537) );
  inv_x1_sg U51946 ( .A(n18214), .X(n50826) );
  inv_x1_sg U51947 ( .A(n19035), .X(n51113) );
  inv_x1_sg U51948 ( .A(n7019), .X(n47109) );
  inv_x1_sg U51949 ( .A(n7837), .X(n47395) );
  inv_x1_sg U51950 ( .A(n8655), .X(n47680) );
  inv_x1_sg U51951 ( .A(n9475), .X(n47965) );
  inv_x1_sg U51952 ( .A(n10294), .X(n48250) );
  inv_x1_sg U51953 ( .A(n11113), .X(n48535) );
  inv_x1_sg U51954 ( .A(n11932), .X(n48820) );
  inv_x1_sg U51955 ( .A(n12751), .X(n49107) );
  inv_x1_sg U51956 ( .A(n13570), .X(n49393) );
  inv_x1_sg U51957 ( .A(n14389), .X(n49679) );
  inv_x1_sg U51958 ( .A(n15208), .X(n49965) );
  inv_x1_sg U51959 ( .A(n16027), .X(n50251) );
  inv_x1_sg U51960 ( .A(n17665), .X(n50825) );
  inv_x1_sg U51961 ( .A(n18486), .X(n51112) );
  inv_x1_sg U51962 ( .A(n7426), .X(n47036) );
  inv_x1_sg U51963 ( .A(n8244), .X(n47323) );
  inv_x1_sg U51964 ( .A(n9062), .X(n47608) );
  inv_x1_sg U51965 ( .A(n9882), .X(n47893) );
  inv_x1_sg U51966 ( .A(n10701), .X(n48178) );
  inv_x1_sg U51967 ( .A(n11520), .X(n48463) );
  inv_x1_sg U51968 ( .A(n12339), .X(n48748) );
  inv_x1_sg U51969 ( .A(n13158), .X(n49034) );
  inv_x1_sg U51970 ( .A(n13977), .X(n49321) );
  inv_x1_sg U51971 ( .A(n14796), .X(n49607) );
  inv_x1_sg U51972 ( .A(n15615), .X(n49893) );
  inv_x1_sg U51973 ( .A(n16434), .X(n50179) );
  inv_x1_sg U51974 ( .A(n18072), .X(n50753) );
  inv_x1_sg U51975 ( .A(n18893), .X(n51040) );
  inv_x1_sg U51976 ( .A(n17251), .X(n50464) );
  inv_x1_sg U51977 ( .A(n7115), .X(n46895) );
  inv_x1_sg U51978 ( .A(n7933), .X(n47190) );
  inv_x1_sg U51979 ( .A(n8751), .X(n47475) );
  inv_x1_sg U51980 ( .A(n9571), .X(n47760) );
  inv_x1_sg U51981 ( .A(n10390), .X(n48045) );
  inv_x1_sg U51982 ( .A(n11209), .X(n48330) );
  inv_x1_sg U51983 ( .A(n12028), .X(n48615) );
  inv_x1_sg U51984 ( .A(n12847), .X(n48901) );
  inv_x1_sg U51985 ( .A(n13666), .X(n49188) );
  inv_x1_sg U51986 ( .A(n14485), .X(n49474) );
  inv_x1_sg U51987 ( .A(n15304), .X(n49760) );
  inv_x1_sg U51988 ( .A(n16123), .X(n50046) );
  inv_x1_sg U51989 ( .A(n16940), .X(n50328) );
  inv_x1_sg U51990 ( .A(n17761), .X(n50620) );
  inv_x1_sg U51991 ( .A(n18582), .X(n50907) );
  inv_x1_sg U51992 ( .A(n7405), .X(n47068) );
  inv_x1_sg U51993 ( .A(n8223), .X(n47354) );
  inv_x1_sg U51994 ( .A(n9041), .X(n47639) );
  inv_x1_sg U51995 ( .A(n9861), .X(n47924) );
  inv_x1_sg U51996 ( .A(n10680), .X(n48209) );
  inv_x1_sg U51997 ( .A(n11499), .X(n48494) );
  inv_x1_sg U51998 ( .A(n12318), .X(n48779) );
  inv_x1_sg U51999 ( .A(n13137), .X(n49066) );
  inv_x1_sg U52000 ( .A(n13956), .X(n49352) );
  inv_x1_sg U52001 ( .A(n14775), .X(n49638) );
  inv_x1_sg U52002 ( .A(n15594), .X(n49924) );
  inv_x1_sg U52003 ( .A(n16413), .X(n50210) );
  inv_x1_sg U52004 ( .A(n17230), .X(n50495) );
  inv_x1_sg U52005 ( .A(n18051), .X(n50784) );
  inv_x1_sg U52006 ( .A(n18872), .X(n51071) );
  inv_x1_sg U52007 ( .A(n6953), .X(n47046) );
  inv_x1_sg U52008 ( .A(n16777), .X(n50474) );
  inv_x1_sg U52009 ( .A(n8082), .X(n47303) );
  inv_x1_sg U52010 ( .A(n8900), .X(n47588) );
  inv_x1_sg U52011 ( .A(n9720), .X(n47873) );
  inv_x1_sg U52012 ( .A(n10539), .X(n48158) );
  inv_x1_sg U52013 ( .A(n11358), .X(n48443) );
  inv_x1_sg U52014 ( .A(n12177), .X(n48728) );
  inv_x1_sg U52015 ( .A(n12996), .X(n49014) );
  inv_x1_sg U52016 ( .A(n13815), .X(n49301) );
  inv_x1_sg U52017 ( .A(n14634), .X(n49587) );
  inv_x1_sg U52018 ( .A(n15453), .X(n49873) );
  inv_x1_sg U52019 ( .A(n16272), .X(n50159) );
  inv_x1_sg U52020 ( .A(n17910), .X(n50733) );
  inv_x1_sg U52021 ( .A(n18731), .X(n51020) );
  inv_x1_sg U52022 ( .A(n7235), .X(n47001) );
  inv_x1_sg U52023 ( .A(n8054), .X(n47290) );
  inv_x1_sg U52024 ( .A(n8132), .X(n47328) );
  inv_x1_sg U52025 ( .A(n8872), .X(n47575) );
  inv_x1_sg U52026 ( .A(n8950), .X(n47613) );
  inv_x1_sg U52027 ( .A(n9692), .X(n47860) );
  inv_x1_sg U52028 ( .A(n9770), .X(n47898) );
  inv_x1_sg U52029 ( .A(n10511), .X(n48145) );
  inv_x1_sg U52030 ( .A(n10589), .X(n48183) );
  inv_x1_sg U52031 ( .A(n11330), .X(n48430) );
  inv_x1_sg U52032 ( .A(n11408), .X(n48468) );
  inv_x1_sg U52033 ( .A(n12149), .X(n48715) );
  inv_x1_sg U52034 ( .A(n12227), .X(n48753) );
  inv_x1_sg U52035 ( .A(n12968), .X(n49001) );
  inv_x1_sg U52036 ( .A(n13046), .X(n49039) );
  inv_x1_sg U52037 ( .A(n13787), .X(n49288) );
  inv_x1_sg U52038 ( .A(n13865), .X(n49326) );
  inv_x1_sg U52039 ( .A(n14606), .X(n49574) );
  inv_x1_sg U52040 ( .A(n14684), .X(n49612) );
  inv_x1_sg U52041 ( .A(n15425), .X(n49860) );
  inv_x1_sg U52042 ( .A(n15503), .X(n49898) );
  inv_x1_sg U52043 ( .A(n16244), .X(n50146) );
  inv_x1_sg U52044 ( .A(n16322), .X(n50184) );
  inv_x1_sg U52045 ( .A(n17060), .X(n50431) );
  inv_x1_sg U52046 ( .A(n17882), .X(n50720) );
  inv_x1_sg U52047 ( .A(n17960), .X(n50758) );
  inv_x1_sg U52048 ( .A(n18703), .X(n51007) );
  inv_x1_sg U52049 ( .A(n18781), .X(n51045) );
  inv_x1_sg U52050 ( .A(n17115), .X(n50428) );
  inv_x1_sg U52051 ( .A(n7415), .X(n47066) );
  inv_x1_sg U52052 ( .A(n8233), .X(n47352) );
  inv_x1_sg U52053 ( .A(n9051), .X(n47637) );
  inv_x1_sg U52054 ( .A(n9871), .X(n47922) );
  inv_x1_sg U52055 ( .A(n10690), .X(n48207) );
  inv_x1_sg U52056 ( .A(n11509), .X(n48492) );
  inv_x1_sg U52057 ( .A(n12328), .X(n48777) );
  inv_x1_sg U52058 ( .A(n13147), .X(n49064) );
  inv_x1_sg U52059 ( .A(n13966), .X(n49350) );
  inv_x1_sg U52060 ( .A(n14785), .X(n49636) );
  inv_x1_sg U52061 ( .A(n15604), .X(n49922) );
  inv_x1_sg U52062 ( .A(n16423), .X(n50208) );
  inv_x1_sg U52063 ( .A(n17240), .X(n50493) );
  inv_x1_sg U52064 ( .A(n18061), .X(n50782) );
  inv_x1_sg U52065 ( .A(n18882), .X(n51069) );
  inv_x1_sg U52066 ( .A(n7615), .X(n47104) );
  inv_x1_sg U52067 ( .A(n8433), .X(n47390) );
  inv_x1_sg U52068 ( .A(n9251), .X(n47675) );
  inv_x1_sg U52069 ( .A(n10071), .X(n47960) );
  inv_x1_sg U52070 ( .A(n10890), .X(n48245) );
  inv_x1_sg U52071 ( .A(n11709), .X(n48530) );
  inv_x1_sg U52072 ( .A(n12528), .X(n48815) );
  inv_x1_sg U52073 ( .A(n13347), .X(n49102) );
  inv_x1_sg U52074 ( .A(n14166), .X(n49388) );
  inv_x1_sg U52075 ( .A(n14985), .X(n49674) );
  inv_x1_sg U52076 ( .A(n15804), .X(n49960) );
  inv_x1_sg U52077 ( .A(n16623), .X(n50246) );
  inv_x1_sg U52078 ( .A(n17440), .X(n50531) );
  inv_x1_sg U52079 ( .A(n18261), .X(n50820) );
  inv_x1_sg U52080 ( .A(n19082), .X(n51107) );
  inv_x1_sg U52081 ( .A(n7198), .X(n46978) );
  inv_x1_sg U52082 ( .A(n8017), .X(n47268) );
  inv_x1_sg U52083 ( .A(n8835), .X(n47553) );
  inv_x1_sg U52084 ( .A(n9655), .X(n47838) );
  inv_x1_sg U52085 ( .A(n10474), .X(n48123) );
  inv_x1_sg U52086 ( .A(n11293), .X(n48408) );
  inv_x1_sg U52087 ( .A(n12112), .X(n48693) );
  inv_x1_sg U52088 ( .A(n12931), .X(n48979) );
  inv_x1_sg U52089 ( .A(n13750), .X(n49266) );
  inv_x1_sg U52090 ( .A(n14569), .X(n49552) );
  inv_x1_sg U52091 ( .A(n15388), .X(n49838) );
  inv_x1_sg U52092 ( .A(n16207), .X(n50124) );
  inv_x1_sg U52093 ( .A(n17023), .X(n50409) );
  inv_x1_sg U52094 ( .A(n17845), .X(n50698) );
  inv_x1_sg U52095 ( .A(n18666), .X(n50985) );
  inv_x1_sg U52096 ( .A(n7290), .X(n46998) );
  nand_x1_sg U52097 ( .A(n7064), .B(n7065), .X(n6865) );
  nand_x1_sg U52098 ( .A(n7882), .B(n7883), .X(n7682) );
  nand_x1_sg U52099 ( .A(n8700), .B(n8701), .X(n8500) );
  nand_x1_sg U52100 ( .A(n9520), .B(n9521), .X(n9320) );
  nand_x1_sg U52101 ( .A(n10339), .B(n10340), .X(n10139) );
  nand_x1_sg U52102 ( .A(n11158), .B(n11159), .X(n10958) );
  nand_x1_sg U52103 ( .A(n11977), .B(n11978), .X(n11777) );
  nand_x1_sg U52104 ( .A(n12796), .B(n12797), .X(n12596) );
  nand_x1_sg U52105 ( .A(n13615), .B(n13616), .X(n13415) );
  nand_x1_sg U52106 ( .A(n14434), .B(n14435), .X(n14234) );
  nand_x1_sg U52107 ( .A(n15253), .B(n15254), .X(n15053) );
  nand_x1_sg U52108 ( .A(n16072), .B(n16073), .X(n15872) );
  nand_x1_sg U52109 ( .A(n16891), .B(n16892), .X(n16689) );
  nand_x1_sg U52110 ( .A(n17710), .B(n17711), .X(n17510) );
  nand_x1_sg U52111 ( .A(n18531), .B(n18532), .X(n18331) );
  inv_x1_sg U52112 ( .A(n6882), .X(n46952) );
  inv_x1_sg U52113 ( .A(n7699), .X(n47243) );
  inv_x1_sg U52114 ( .A(n8517), .X(n47528) );
  inv_x1_sg U52115 ( .A(n9337), .X(n47813) );
  inv_x1_sg U52116 ( .A(n10156), .X(n48098) );
  inv_x1_sg U52117 ( .A(n10975), .X(n48383) );
  inv_x1_sg U52118 ( .A(n11794), .X(n48668) );
  inv_x1_sg U52119 ( .A(n12613), .X(n48954) );
  inv_x1_sg U52120 ( .A(n13432), .X(n49241) );
  inv_x1_sg U52121 ( .A(n14251), .X(n49527) );
  inv_x1_sg U52122 ( .A(n15070), .X(n49813) );
  inv_x1_sg U52123 ( .A(n15889), .X(n50099) );
  inv_x1_sg U52124 ( .A(n17527), .X(n50673) );
  inv_x1_sg U52125 ( .A(n18348), .X(n50960) );
  nand_x1_sg U52126 ( .A(n7246), .B(n7227), .X(n7241) );
  nand_x1_sg U52127 ( .A(n8065), .B(n8046), .X(n8060) );
  nand_x1_sg U52128 ( .A(n8883), .B(n8864), .X(n8878) );
  nand_x1_sg U52129 ( .A(n9703), .B(n9684), .X(n9698) );
  nand_x1_sg U52130 ( .A(n10522), .B(n10503), .X(n10517) );
  nand_x1_sg U52131 ( .A(n11341), .B(n11322), .X(n11336) );
  nand_x1_sg U52132 ( .A(n12160), .B(n12141), .X(n12155) );
  nand_x1_sg U52133 ( .A(n12979), .B(n12960), .X(n12974) );
  nand_x1_sg U52134 ( .A(n13798), .B(n13779), .X(n13793) );
  nand_x1_sg U52135 ( .A(n14617), .B(n14598), .X(n14612) );
  nand_x1_sg U52136 ( .A(n15436), .B(n15417), .X(n15431) );
  nand_x1_sg U52137 ( .A(n16255), .B(n16236), .X(n16250) );
  nand_x1_sg U52138 ( .A(n17071), .B(n17052), .X(n17066) );
  nand_x1_sg U52139 ( .A(n17893), .B(n17874), .X(n17888) );
  nand_x1_sg U52140 ( .A(n18714), .B(n18695), .X(n18709) );
  nand_x1_sg U52141 ( .A(n7149), .B(n7142), .X(n7147) );
  nand_x1_sg U52142 ( .A(n7967), .B(n7960), .X(n7965) );
  nand_x1_sg U52143 ( .A(n8785), .B(n8778), .X(n8783) );
  nand_x1_sg U52144 ( .A(n9605), .B(n9598), .X(n9603) );
  nand_x1_sg U52145 ( .A(n10424), .B(n10417), .X(n10422) );
  nand_x1_sg U52146 ( .A(n11243), .B(n11236), .X(n11241) );
  nand_x1_sg U52147 ( .A(n12062), .B(n12055), .X(n12060) );
  nand_x1_sg U52148 ( .A(n12881), .B(n12874), .X(n12879) );
  nand_x1_sg U52149 ( .A(n13700), .B(n13693), .X(n13698) );
  nand_x1_sg U52150 ( .A(n14519), .B(n14512), .X(n14517) );
  nand_x1_sg U52151 ( .A(n15338), .B(n15331), .X(n15336) );
  nand_x1_sg U52152 ( .A(n16157), .B(n16150), .X(n16155) );
  nand_x1_sg U52153 ( .A(n16974), .B(n16967), .X(n16972) );
  nand_x1_sg U52154 ( .A(n17795), .B(n17788), .X(n17793) );
  nand_x1_sg U52155 ( .A(n18616), .B(n18609), .X(n18614) );
  inv_x1_sg U52156 ( .A(n7228), .X(n46946) );
  inv_x1_sg U52157 ( .A(n17053), .X(n50378) );
  inv_x1_sg U52158 ( .A(n8108), .X(n47287) );
  inv_x1_sg U52159 ( .A(n8926), .X(n47572) );
  inv_x1_sg U52160 ( .A(n9746), .X(n47857) );
  inv_x1_sg U52161 ( .A(n10565), .X(n48142) );
  inv_x1_sg U52162 ( .A(n11384), .X(n48427) );
  inv_x1_sg U52163 ( .A(n12203), .X(n48712) );
  inv_x1_sg U52164 ( .A(n13022), .X(n48998) );
  inv_x1_sg U52165 ( .A(n13841), .X(n49285) );
  inv_x1_sg U52166 ( .A(n14660), .X(n49571) );
  inv_x1_sg U52167 ( .A(n15479), .X(n49857) );
  inv_x1_sg U52168 ( .A(n16298), .X(n50143) );
  inv_x1_sg U52169 ( .A(n17936), .X(n50717) );
  inv_x1_sg U52170 ( .A(n18757), .X(n51004) );
  inv_x1_sg U52171 ( .A(n7143), .X(n46909) );
  inv_x1_sg U52172 ( .A(n7961), .X(n47202) );
  inv_x1_sg U52173 ( .A(n8779), .X(n47487) );
  inv_x1_sg U52174 ( .A(n9599), .X(n47772) );
  inv_x1_sg U52175 ( .A(n10418), .X(n48057) );
  inv_x1_sg U52176 ( .A(n11237), .X(n48342) );
  inv_x1_sg U52177 ( .A(n12056), .X(n48627) );
  inv_x1_sg U52178 ( .A(n12875), .X(n48913) );
  inv_x1_sg U52179 ( .A(n13694), .X(n49200) );
  inv_x1_sg U52180 ( .A(n14513), .X(n49486) );
  inv_x1_sg U52181 ( .A(n15332), .X(n49772) );
  inv_x1_sg U52182 ( .A(n16151), .X(n50058) );
  inv_x1_sg U52183 ( .A(n16968), .X(n50343) );
  inv_x1_sg U52184 ( .A(n17789), .X(n50632) );
  inv_x1_sg U52185 ( .A(n18610), .X(n50919) );
  inv_x1_sg U52186 ( .A(n7177), .X(n46928) );
  inv_x1_sg U52187 ( .A(n7996), .X(n47220) );
  inv_x1_sg U52188 ( .A(n8814), .X(n47505) );
  inv_x1_sg U52189 ( .A(n9634), .X(n47790) );
  inv_x1_sg U52190 ( .A(n10453), .X(n48075) );
  inv_x1_sg U52191 ( .A(n11272), .X(n48360) );
  inv_x1_sg U52192 ( .A(n12091), .X(n48645) );
  inv_x1_sg U52193 ( .A(n12910), .X(n48931) );
  inv_x1_sg U52194 ( .A(n13729), .X(n49218) );
  inv_x1_sg U52195 ( .A(n14548), .X(n49504) );
  inv_x1_sg U52196 ( .A(n15367), .X(n49790) );
  inv_x1_sg U52197 ( .A(n16186), .X(n50076) );
  inv_x1_sg U52198 ( .A(n17002), .X(n50361) );
  inv_x1_sg U52199 ( .A(n17824), .X(n50650) );
  inv_x1_sg U52200 ( .A(n18645), .X(n50937) );
  inv_x1_sg U52201 ( .A(n7589), .X(n47047) );
  inv_x1_sg U52202 ( .A(n17414), .X(n50475) );
  inv_x1_sg U52203 ( .A(n7564), .X(n47050) );
  inv_x1_sg U52204 ( .A(n17389), .X(n50478) );
  inv_x1_sg U52205 ( .A(n8382), .X(n47337) );
  inv_x1_sg U52206 ( .A(n9200), .X(n47622) );
  inv_x1_sg U52207 ( .A(n10020), .X(n47907) );
  inv_x1_sg U52208 ( .A(n10839), .X(n48192) );
  inv_x1_sg U52209 ( .A(n11658), .X(n48477) );
  inv_x1_sg U52210 ( .A(n12477), .X(n48762) );
  inv_x1_sg U52211 ( .A(n13296), .X(n49048) );
  inv_x1_sg U52212 ( .A(n14115), .X(n49335) );
  inv_x1_sg U52213 ( .A(n14934), .X(n49621) );
  inv_x1_sg U52214 ( .A(n15753), .X(n49907) );
  inv_x1_sg U52215 ( .A(n16572), .X(n50193) );
  inv_x1_sg U52216 ( .A(n18210), .X(n50767) );
  inv_x1_sg U52217 ( .A(n19031), .X(n51054) );
  inv_x1_sg U52218 ( .A(n7071), .X(n46860) );
  inv_x1_sg U52219 ( .A(n7889), .X(n47153) );
  inv_x1_sg U52220 ( .A(n8707), .X(n47438) );
  inv_x1_sg U52221 ( .A(n9527), .X(n47723) );
  inv_x1_sg U52222 ( .A(n10346), .X(n48008) );
  inv_x1_sg U52223 ( .A(n11165), .X(n48293) );
  inv_x1_sg U52224 ( .A(n11984), .X(n48578) );
  inv_x1_sg U52225 ( .A(n12803), .X(n48864) );
  inv_x1_sg U52226 ( .A(n13622), .X(n49151) );
  inv_x1_sg U52227 ( .A(n14441), .X(n49437) );
  inv_x1_sg U52228 ( .A(n15260), .X(n49722) );
  inv_x1_sg U52229 ( .A(n16079), .X(n50009) );
  inv_x1_sg U52230 ( .A(n16898), .X(n50293) );
  inv_x1_sg U52231 ( .A(n17717), .X(n50583) );
  inv_x1_sg U52232 ( .A(n18538), .X(n50870) );
  inv_x1_sg U52233 ( .A(n17246), .X(n50448) );
  inv_x1_sg U52234 ( .A(n7595), .X(n47106) );
  inv_x1_sg U52235 ( .A(n8413), .X(n47392) );
  inv_x1_sg U52236 ( .A(n9231), .X(n47677) );
  inv_x1_sg U52237 ( .A(n10051), .X(n47962) );
  inv_x1_sg U52238 ( .A(n10870), .X(n48247) );
  inv_x1_sg U52239 ( .A(n11689), .X(n48532) );
  inv_x1_sg U52240 ( .A(n12508), .X(n48817) );
  inv_x1_sg U52241 ( .A(n13327), .X(n49104) );
  inv_x1_sg U52242 ( .A(n14146), .X(n49390) );
  inv_x1_sg U52243 ( .A(n14965), .X(n49676) );
  inv_x1_sg U52244 ( .A(n15784), .X(n49962) );
  inv_x1_sg U52245 ( .A(n16603), .X(n50248) );
  inv_x1_sg U52246 ( .A(n17420), .X(n50533) );
  inv_x1_sg U52247 ( .A(n18241), .X(n50822) );
  inv_x1_sg U52248 ( .A(n19062), .X(n51109) );
  inv_x1_sg U52249 ( .A(n7463), .X(n47023) );
  inv_x1_sg U52250 ( .A(n8281), .X(n47311) );
  inv_x1_sg U52251 ( .A(n9099), .X(n47596) );
  inv_x1_sg U52252 ( .A(n9919), .X(n47881) );
  inv_x1_sg U52253 ( .A(n10738), .X(n48166) );
  inv_x1_sg U52254 ( .A(n11557), .X(n48451) );
  inv_x1_sg U52255 ( .A(n12376), .X(n48736) );
  inv_x1_sg U52256 ( .A(n13195), .X(n49022) );
  inv_x1_sg U52257 ( .A(n14014), .X(n49309) );
  inv_x1_sg U52258 ( .A(n14833), .X(n49595) );
  inv_x1_sg U52259 ( .A(n15652), .X(n49881) );
  inv_x1_sg U52260 ( .A(n16471), .X(n50167) );
  inv_x1_sg U52261 ( .A(n18109), .X(n50741) );
  inv_x1_sg U52262 ( .A(n18930), .X(n51028) );
  inv_x1_sg U52263 ( .A(n17288), .X(n50452) );
  inv_x1_sg U52264 ( .A(n7554), .X(n47052) );
  inv_x1_sg U52265 ( .A(n8372), .X(n47339) );
  inv_x1_sg U52266 ( .A(n9190), .X(n47624) );
  inv_x1_sg U52267 ( .A(n10010), .X(n47909) );
  inv_x1_sg U52268 ( .A(n10829), .X(n48194) );
  inv_x1_sg U52269 ( .A(n11648), .X(n48479) );
  inv_x1_sg U52270 ( .A(n12467), .X(n48764) );
  inv_x1_sg U52271 ( .A(n13286), .X(n49050) );
  inv_x1_sg U52272 ( .A(n14105), .X(n49337) );
  inv_x1_sg U52273 ( .A(n14924), .X(n49623) );
  inv_x1_sg U52274 ( .A(n15743), .X(n49909) );
  inv_x1_sg U52275 ( .A(n16562), .X(n50195) );
  inv_x1_sg U52276 ( .A(n17379), .X(n50480) );
  inv_x1_sg U52277 ( .A(n18200), .X(n50769) );
  inv_x1_sg U52278 ( .A(n19021), .X(n51056) );
  inv_x1_sg U52279 ( .A(n17204), .X(n50398) );
  inv_x1_sg U52280 ( .A(n17114), .X(n50352) );
  inv_x1_sg U52281 ( .A(n6977), .X(n47123) );
  inv_x1_sg U52282 ( .A(n7794), .X(n47409) );
  inv_x1_sg U52283 ( .A(n8612), .X(n47694) );
  inv_x1_sg U52284 ( .A(n9432), .X(n47979) );
  inv_x1_sg U52285 ( .A(n10251), .X(n48264) );
  inv_x1_sg U52286 ( .A(n11070), .X(n48549) );
  inv_x1_sg U52287 ( .A(n11889), .X(n48834) );
  inv_x1_sg U52288 ( .A(n12708), .X(n49121) );
  inv_x1_sg U52289 ( .A(n13527), .X(n49407) );
  inv_x1_sg U52290 ( .A(n14346), .X(n49693) );
  inv_x1_sg U52291 ( .A(n15165), .X(n49979) );
  inv_x1_sg U52292 ( .A(n15984), .X(n50265) );
  inv_x1_sg U52293 ( .A(n16801), .X(n50551) );
  inv_x1_sg U52294 ( .A(n17622), .X(n50839) );
  inv_x1_sg U52295 ( .A(n18443), .X(n51126) );
  inv_x1_sg U52296 ( .A(n7663), .X(n47155) );
  inv_x1_sg U52297 ( .A(n8481), .X(n47440) );
  inv_x1_sg U52298 ( .A(n9301), .X(n47725) );
  inv_x1_sg U52299 ( .A(n10120), .X(n48010) );
  inv_x1_sg U52300 ( .A(n10939), .X(n48295) );
  inv_x1_sg U52301 ( .A(n11758), .X(n48580) );
  inv_x1_sg U52302 ( .A(n12577), .X(n48866) );
  inv_x1_sg U52303 ( .A(n13396), .X(n49153) );
  inv_x1_sg U52304 ( .A(n14215), .X(n49439) );
  inv_x1_sg U52305 ( .A(n15034), .X(n49724) );
  inv_x1_sg U52306 ( .A(n15853), .X(n50011) );
  inv_x1_sg U52307 ( .A(n16670), .X(n50295) );
  inv_x1_sg U52308 ( .A(n17491), .X(n50585) );
  inv_x1_sg U52309 ( .A(n18312), .X(n50872) );
  inv_x1_sg U52310 ( .A(n7307), .X(n46997) );
  inv_x1_sg U52311 ( .A(n8125), .X(n47286) );
  inv_x1_sg U52312 ( .A(n8943), .X(n47571) );
  inv_x1_sg U52313 ( .A(n9763), .X(n47856) );
  inv_x1_sg U52314 ( .A(n10582), .X(n48141) );
  inv_x1_sg U52315 ( .A(n11401), .X(n48426) );
  inv_x1_sg U52316 ( .A(n12220), .X(n48711) );
  inv_x1_sg U52317 ( .A(n13039), .X(n48997) );
  inv_x1_sg U52318 ( .A(n13858), .X(n49284) );
  inv_x1_sg U52319 ( .A(n14677), .X(n49570) );
  inv_x1_sg U52320 ( .A(n15496), .X(n49856) );
  inv_x1_sg U52321 ( .A(n16315), .X(n50142) );
  inv_x1_sg U52322 ( .A(n17953), .X(n50716) );
  inv_x1_sg U52323 ( .A(n18774), .X(n51003) );
  inv_x1_sg U52324 ( .A(n7447), .X(n47030) );
  inv_x1_sg U52325 ( .A(n8265), .X(n47317) );
  inv_x1_sg U52326 ( .A(n9083), .X(n47602) );
  inv_x1_sg U52327 ( .A(n9903), .X(n47887) );
  inv_x1_sg U52328 ( .A(n10722), .X(n48172) );
  inv_x1_sg U52329 ( .A(n11541), .X(n48457) );
  inv_x1_sg U52330 ( .A(n12360), .X(n48742) );
  inv_x1_sg U52331 ( .A(n13179), .X(n49028) );
  inv_x1_sg U52332 ( .A(n13998), .X(n49315) );
  inv_x1_sg U52333 ( .A(n14817), .X(n49601) );
  inv_x1_sg U52334 ( .A(n15636), .X(n49887) );
  inv_x1_sg U52335 ( .A(n16455), .X(n50173) );
  inv_x1_sg U52336 ( .A(n17272), .X(n50458) );
  inv_x1_sg U52337 ( .A(n18093), .X(n50747) );
  inv_x1_sg U52338 ( .A(n18914), .X(n51034) );
  inv_x1_sg U52339 ( .A(n16997), .X(n50383) );
  inv_x1_sg U52340 ( .A(n7248), .X(n46934) );
  inv_x1_sg U52341 ( .A(n8067), .X(n47226) );
  inv_x1_sg U52342 ( .A(n8885), .X(n47511) );
  inv_x1_sg U52343 ( .A(n9705), .X(n47796) );
  inv_x1_sg U52344 ( .A(n10524), .X(n48081) );
  inv_x1_sg U52345 ( .A(n11343), .X(n48366) );
  inv_x1_sg U52346 ( .A(n12162), .X(n48651) );
  inv_x1_sg U52347 ( .A(n12981), .X(n48937) );
  inv_x1_sg U52348 ( .A(n13800), .X(n49224) );
  inv_x1_sg U52349 ( .A(n14619), .X(n49510) );
  inv_x1_sg U52350 ( .A(n15438), .X(n49796) );
  inv_x1_sg U52351 ( .A(n16257), .X(n50082) );
  inv_x1_sg U52352 ( .A(n17895), .X(n50656) );
  inv_x1_sg U52353 ( .A(n18716), .X(n50943) );
  inv_x1_sg U52354 ( .A(n17073), .X(n50367) );
  inv_x1_sg U52355 ( .A(n7219), .X(n46948) );
  inv_x1_sg U52356 ( .A(n8038), .X(n47239) );
  inv_x1_sg U52357 ( .A(n8856), .X(n47524) );
  inv_x1_sg U52358 ( .A(n9676), .X(n47809) );
  inv_x1_sg U52359 ( .A(n10495), .X(n48094) );
  inv_x1_sg U52360 ( .A(n11314), .X(n48379) );
  inv_x1_sg U52361 ( .A(n12133), .X(n48664) );
  inv_x1_sg U52362 ( .A(n12952), .X(n48950) );
  inv_x1_sg U52363 ( .A(n13771), .X(n49237) );
  inv_x1_sg U52364 ( .A(n14590), .X(n49523) );
  inv_x1_sg U52365 ( .A(n15409), .X(n49809) );
  inv_x1_sg U52366 ( .A(n16228), .X(n50095) );
  inv_x1_sg U52367 ( .A(n17044), .X(n50380) );
  inv_x1_sg U52368 ( .A(n17866), .X(n50669) );
  inv_x1_sg U52369 ( .A(n18687), .X(n50956) );
  inv_x1_sg U52370 ( .A(n7539), .X(n47084) );
  inv_x1_sg U52371 ( .A(n8357), .X(n47370) );
  inv_x1_sg U52372 ( .A(n9175), .X(n47655) );
  inv_x1_sg U52373 ( .A(n9995), .X(n47940) );
  inv_x1_sg U52374 ( .A(n10814), .X(n48225) );
  inv_x1_sg U52375 ( .A(n11633), .X(n48510) );
  inv_x1_sg U52376 ( .A(n12452), .X(n48795) );
  inv_x1_sg U52377 ( .A(n13271), .X(n49082) );
  inv_x1_sg U52378 ( .A(n14090), .X(n49368) );
  inv_x1_sg U52379 ( .A(n14909), .X(n49654) );
  inv_x1_sg U52380 ( .A(n15728), .X(n49940) );
  inv_x1_sg U52381 ( .A(n16547), .X(n50226) );
  inv_x1_sg U52382 ( .A(n17364), .X(n50511) );
  inv_x1_sg U52383 ( .A(n18185), .X(n50800) );
  inv_x1_sg U52384 ( .A(n19006), .X(n51087) );
  inv_x1_sg U52385 ( .A(n17387), .X(n50392) );
  inv_x1_sg U52386 ( .A(n7304), .X(n46944) );
  inv_x1_sg U52387 ( .A(n17950), .X(n50665) );
  inv_x1_sg U52388 ( .A(n8122), .X(n47235) );
  inv_x1_sg U52389 ( .A(n8940), .X(n47520) );
  inv_x1_sg U52390 ( .A(n9760), .X(n47805) );
  inv_x1_sg U52391 ( .A(n10579), .X(n48090) );
  inv_x1_sg U52392 ( .A(n11398), .X(n48375) );
  inv_x1_sg U52393 ( .A(n12217), .X(n48660) );
  inv_x1_sg U52394 ( .A(n13036), .X(n48946) );
  inv_x1_sg U52395 ( .A(n13855), .X(n49233) );
  inv_x1_sg U52396 ( .A(n14674), .X(n49519) );
  inv_x1_sg U52397 ( .A(n15493), .X(n49805) );
  inv_x1_sg U52398 ( .A(n16312), .X(n50091) );
  inv_x1_sg U52399 ( .A(n18771), .X(n50952) );
  inv_x1_sg U52400 ( .A(n6986), .X(n47077) );
  inv_x1_sg U52401 ( .A(n7803), .X(n47363) );
  inv_x1_sg U52402 ( .A(n8621), .X(n47648) );
  inv_x1_sg U52403 ( .A(n9441), .X(n47933) );
  inv_x1_sg U52404 ( .A(n10260), .X(n48218) );
  inv_x1_sg U52405 ( .A(n11079), .X(n48503) );
  inv_x1_sg U52406 ( .A(n11898), .X(n48788) );
  inv_x1_sg U52407 ( .A(n12717), .X(n49075) );
  inv_x1_sg U52408 ( .A(n13536), .X(n49361) );
  inv_x1_sg U52409 ( .A(n14355), .X(n49647) );
  inv_x1_sg U52410 ( .A(n15174), .X(n49933) );
  inv_x1_sg U52411 ( .A(n15993), .X(n50219) );
  inv_x1_sg U52412 ( .A(n16810), .X(n50504) );
  inv_x1_sg U52413 ( .A(n17631), .X(n50793) );
  inv_x1_sg U52414 ( .A(n18452), .X(n51080) );
  inv_x1_sg U52415 ( .A(n7613), .X(n47059) );
  inv_x1_sg U52416 ( .A(n17438), .X(n50486) );
  inv_x1_sg U52417 ( .A(n17258), .X(n50368) );
  inv_x1_sg U52418 ( .A(n17330), .X(n50417) );
  inv_x1_sg U52419 ( .A(n7505), .X(n46987) );
  inv_x1_sg U52420 ( .A(n8323), .X(n47276) );
  inv_x1_sg U52421 ( .A(n9141), .X(n47561) );
  inv_x1_sg U52422 ( .A(n9961), .X(n47846) );
  inv_x1_sg U52423 ( .A(n10780), .X(n48131) );
  inv_x1_sg U52424 ( .A(n11599), .X(n48416) );
  inv_x1_sg U52425 ( .A(n12418), .X(n48701) );
  inv_x1_sg U52426 ( .A(n13237), .X(n48987) );
  inv_x1_sg U52427 ( .A(n14056), .X(n49274) );
  inv_x1_sg U52428 ( .A(n14875), .X(n49560) );
  inv_x1_sg U52429 ( .A(n15694), .X(n49846) );
  inv_x1_sg U52430 ( .A(n16513), .X(n50132) );
  inv_x1_sg U52431 ( .A(n18151), .X(n50706) );
  inv_x1_sg U52432 ( .A(n18972), .X(n50993) );
  inv_x1_sg U52433 ( .A(n17317), .X(n50387) );
  inv_x1_sg U52434 ( .A(n6970), .X(n47098) );
  inv_x1_sg U52435 ( .A(n17615), .X(n50814) );
  inv_x1_sg U52436 ( .A(n7787), .X(n47384) );
  inv_x1_sg U52437 ( .A(n8605), .X(n47669) );
  inv_x1_sg U52438 ( .A(n9425), .X(n47954) );
  inv_x1_sg U52439 ( .A(n10244), .X(n48239) );
  inv_x1_sg U52440 ( .A(n11063), .X(n48524) );
  inv_x1_sg U52441 ( .A(n11882), .X(n48809) );
  inv_x1_sg U52442 ( .A(n12701), .X(n49096) );
  inv_x1_sg U52443 ( .A(n13520), .X(n49382) );
  inv_x1_sg U52444 ( .A(n14339), .X(n49668) );
  inv_x1_sg U52445 ( .A(n15158), .X(n49954) );
  inv_x1_sg U52446 ( .A(n15977), .X(n50240) );
  inv_x1_sg U52447 ( .A(n16794), .X(n50526) );
  inv_x1_sg U52448 ( .A(n18436), .X(n51101) );
  inv_x1_sg U52449 ( .A(n7023), .X(n47062) );
  inv_x1_sg U52450 ( .A(n7841), .X(n47348) );
  inv_x1_sg U52451 ( .A(n8659), .X(n47633) );
  inv_x1_sg U52452 ( .A(n9479), .X(n47918) );
  inv_x1_sg U52453 ( .A(n10298), .X(n48203) );
  inv_x1_sg U52454 ( .A(n11117), .X(n48488) );
  inv_x1_sg U52455 ( .A(n11936), .X(n48773) );
  inv_x1_sg U52456 ( .A(n12755), .X(n49060) );
  inv_x1_sg U52457 ( .A(n13574), .X(n49346) );
  inv_x1_sg U52458 ( .A(n14393), .X(n49632) );
  inv_x1_sg U52459 ( .A(n15212), .X(n49918) );
  inv_x1_sg U52460 ( .A(n16031), .X(n50204) );
  inv_x1_sg U52461 ( .A(n17669), .X(n50778) );
  inv_x1_sg U52462 ( .A(n18490), .X(n51065) );
  inv_x1_sg U52463 ( .A(n6846), .X(n46862) );
  inv_x1_sg U52464 ( .A(n7162), .X(n46908) );
  inv_x1_sg U52465 ( .A(n7981), .X(n47201) );
  inv_x1_sg U52466 ( .A(n8799), .X(n47486) );
  inv_x1_sg U52467 ( .A(n9619), .X(n47771) );
  inv_x1_sg U52468 ( .A(n10438), .X(n48056) );
  inv_x1_sg U52469 ( .A(n11257), .X(n48341) );
  inv_x1_sg U52470 ( .A(n12076), .X(n48626) );
  inv_x1_sg U52471 ( .A(n12895), .X(n48912) );
  inv_x1_sg U52472 ( .A(n13714), .X(n49199) );
  inv_x1_sg U52473 ( .A(n14533), .X(n49485) );
  inv_x1_sg U52474 ( .A(n15352), .X(n49771) );
  inv_x1_sg U52475 ( .A(n16171), .X(n50057) );
  inv_x1_sg U52476 ( .A(n16987), .X(n50342) );
  inv_x1_sg U52477 ( .A(n17809), .X(n50631) );
  inv_x1_sg U52478 ( .A(n18630), .X(n50918) );
  inv_x1_sg U52479 ( .A(n7313), .X(n47014) );
  inv_x1_sg U52480 ( .A(n17138), .X(n50443) );
  inv_x1_sg U52481 ( .A(n7513), .X(n47087) );
  inv_x1_sg U52482 ( .A(n8331), .X(n47373) );
  inv_x1_sg U52483 ( .A(n9149), .X(n47658) );
  inv_x1_sg U52484 ( .A(n9969), .X(n47943) );
  inv_x1_sg U52485 ( .A(n10788), .X(n48228) );
  inv_x1_sg U52486 ( .A(n11607), .X(n48513) );
  inv_x1_sg U52487 ( .A(n12426), .X(n48798) );
  inv_x1_sg U52488 ( .A(n13245), .X(n49085) );
  inv_x1_sg U52489 ( .A(n14064), .X(n49371) );
  inv_x1_sg U52490 ( .A(n14883), .X(n49657) );
  inv_x1_sg U52491 ( .A(n15702), .X(n49943) );
  inv_x1_sg U52492 ( .A(n16521), .X(n50229) );
  inv_x1_sg U52493 ( .A(n17338), .X(n50514) );
  inv_x1_sg U52494 ( .A(n18159), .X(n50803) );
  inv_x1_sg U52495 ( .A(n18980), .X(n51090) );
  inv_x1_sg U52496 ( .A(n7193), .X(n46927) );
  inv_x1_sg U52497 ( .A(n8012), .X(n47219) );
  inv_x1_sg U52498 ( .A(n8830), .X(n47504) );
  inv_x1_sg U52499 ( .A(n9650), .X(n47789) );
  inv_x1_sg U52500 ( .A(n10469), .X(n48074) );
  inv_x1_sg U52501 ( .A(n11288), .X(n48359) );
  inv_x1_sg U52502 ( .A(n12107), .X(n48644) );
  inv_x1_sg U52503 ( .A(n12926), .X(n48930) );
  inv_x1_sg U52504 ( .A(n13745), .X(n49217) );
  inv_x1_sg U52505 ( .A(n14564), .X(n49503) );
  inv_x1_sg U52506 ( .A(n15383), .X(n49789) );
  inv_x1_sg U52507 ( .A(n16202), .X(n50075) );
  inv_x1_sg U52508 ( .A(n17018), .X(n50360) );
  inv_x1_sg U52509 ( .A(n17840), .X(n50649) );
  inv_x1_sg U52510 ( .A(n18661), .X(n50936) );
  inv_x1_sg U52511 ( .A(n16844), .X(n50536) );
  inv_x1_sg U52512 ( .A(n7770), .X(n47333) );
  inv_x1_sg U52513 ( .A(n8588), .X(n47618) );
  inv_x1_sg U52514 ( .A(n9408), .X(n47903) );
  inv_x1_sg U52515 ( .A(n10227), .X(n48188) );
  inv_x1_sg U52516 ( .A(n11046), .X(n48473) );
  inv_x1_sg U52517 ( .A(n11865), .X(n48758) );
  inv_x1_sg U52518 ( .A(n12684), .X(n49044) );
  inv_x1_sg U52519 ( .A(n13503), .X(n49331) );
  inv_x1_sg U52520 ( .A(n14322), .X(n49617) );
  inv_x1_sg U52521 ( .A(n15141), .X(n49903) );
  inv_x1_sg U52522 ( .A(n15960), .X(n50189) );
  inv_x1_sg U52523 ( .A(n17598), .X(n50763) );
  inv_x1_sg U52524 ( .A(n18419), .X(n51050) );
  nand_x1_sg U52525 ( .A(n6957), .B(n46991), .X(n6956) );
  nand_x1_sg U52526 ( .A(n7774), .B(n47280), .X(n7773) );
  nand_x1_sg U52527 ( .A(n8592), .B(n47565), .X(n8591) );
  nand_x1_sg U52528 ( .A(n9412), .B(n47850), .X(n9411) );
  nand_x1_sg U52529 ( .A(n10231), .B(n48135), .X(n10230) );
  nand_x1_sg U52530 ( .A(n11050), .B(n48420), .X(n11049) );
  nand_x1_sg U52531 ( .A(n11869), .B(n48705), .X(n11868) );
  nand_x1_sg U52532 ( .A(n12688), .B(n48991), .X(n12687) );
  nand_x1_sg U52533 ( .A(n13507), .B(n49278), .X(n13506) );
  nand_x1_sg U52534 ( .A(n14326), .B(n49564), .X(n14325) );
  nand_x1_sg U52535 ( .A(n15145), .B(n49850), .X(n15144) );
  nand_x1_sg U52536 ( .A(n15964), .B(n50136), .X(n15963) );
  nand_x1_sg U52537 ( .A(n17602), .B(n50710), .X(n17601) );
  nand_x1_sg U52538 ( .A(n18423), .B(n50997), .X(n18422) );
  nand_x1_sg U52539 ( .A(n16781), .B(n50421), .X(n16780) );
  inv_x1_sg U52540 ( .A(n7323), .X(n46995) );
  inv_x1_sg U52541 ( .A(n17148), .X(n50425) );
  inv_x1_sg U52542 ( .A(n16971), .X(n50363) );
  inv_x1_sg U52543 ( .A(n7497), .X(n47028) );
  inv_x1_sg U52544 ( .A(n8315), .X(n47315) );
  inv_x1_sg U52545 ( .A(n9133), .X(n47600) );
  inv_x1_sg U52546 ( .A(n9953), .X(n47885) );
  inv_x1_sg U52547 ( .A(n10772), .X(n48170) );
  inv_x1_sg U52548 ( .A(n11591), .X(n48455) );
  inv_x1_sg U52549 ( .A(n12410), .X(n48740) );
  inv_x1_sg U52550 ( .A(n13229), .X(n49026) );
  inv_x1_sg U52551 ( .A(n14048), .X(n49313) );
  inv_x1_sg U52552 ( .A(n14867), .X(n49599) );
  inv_x1_sg U52553 ( .A(n15686), .X(n49885) );
  inv_x1_sg U52554 ( .A(n16505), .X(n50171) );
  inv_x1_sg U52555 ( .A(n17322), .X(n50456) );
  inv_x1_sg U52556 ( .A(n18143), .X(n50745) );
  inv_x1_sg U52557 ( .A(n18964), .X(n51032) );
  inv_x1_sg U52558 ( .A(n7146), .X(n46930) );
  inv_x1_sg U52559 ( .A(n7964), .X(n47222) );
  inv_x1_sg U52560 ( .A(n8782), .X(n47507) );
  inv_x1_sg U52561 ( .A(n9602), .X(n47792) );
  inv_x1_sg U52562 ( .A(n10421), .X(n48077) );
  inv_x1_sg U52563 ( .A(n11240), .X(n48362) );
  inv_x1_sg U52564 ( .A(n12059), .X(n48647) );
  inv_x1_sg U52565 ( .A(n12878), .X(n48933) );
  inv_x1_sg U52566 ( .A(n13697), .X(n49220) );
  inv_x1_sg U52567 ( .A(n14516), .X(n49506) );
  inv_x1_sg U52568 ( .A(n15335), .X(n49792) );
  inv_x1_sg U52569 ( .A(n16154), .X(n50078) );
  inv_x1_sg U52570 ( .A(n17792), .X(n50652) );
  inv_x1_sg U52571 ( .A(n18613), .X(n50939) );
  inv_x1_sg U52572 ( .A(n6864), .X(n46897) );
  inv_x1_sg U52573 ( .A(n7681), .X(n47192) );
  inv_x1_sg U52574 ( .A(n8499), .X(n47477) );
  inv_x1_sg U52575 ( .A(n9319), .X(n47762) );
  inv_x1_sg U52576 ( .A(n10138), .X(n48047) );
  inv_x1_sg U52577 ( .A(n10957), .X(n48332) );
  inv_x1_sg U52578 ( .A(n11776), .X(n48617) );
  inv_x1_sg U52579 ( .A(n12595), .X(n48903) );
  inv_x1_sg U52580 ( .A(n13414), .X(n49190) );
  inv_x1_sg U52581 ( .A(n14233), .X(n49476) );
  inv_x1_sg U52582 ( .A(n15052), .X(n49762) );
  inv_x1_sg U52583 ( .A(n15871), .X(n50048) );
  inv_x1_sg U52584 ( .A(n16688), .X(n50330) );
  inv_x1_sg U52585 ( .A(n17509), .X(n50622) );
  inv_x1_sg U52586 ( .A(n18330), .X(n50909) );
  inv_x1_sg U52587 ( .A(n6870), .X(n46912) );
  inv_x1_sg U52588 ( .A(n7687), .X(n47205) );
  inv_x1_sg U52589 ( .A(n8505), .X(n47490) );
  inv_x1_sg U52590 ( .A(n9325), .X(n47775) );
  inv_x1_sg U52591 ( .A(n10144), .X(n48060) );
  inv_x1_sg U52592 ( .A(n10963), .X(n48345) );
  inv_x1_sg U52593 ( .A(n11782), .X(n48630) );
  inv_x1_sg U52594 ( .A(n12601), .X(n48916) );
  inv_x1_sg U52595 ( .A(n13420), .X(n49203) );
  inv_x1_sg U52596 ( .A(n14239), .X(n49489) );
  inv_x1_sg U52597 ( .A(n15058), .X(n49775) );
  inv_x1_sg U52598 ( .A(n15877), .X(n50061) );
  inv_x1_sg U52599 ( .A(n16694), .X(n50346) );
  inv_x1_sg U52600 ( .A(n17515), .X(n50635) );
  inv_x1_sg U52601 ( .A(n18336), .X(n50922) );
  inv_x1_sg U52602 ( .A(n25993), .X(n51312) );
  inv_x1_sg U52603 ( .A(n26006), .X(n51313) );
  inv_x1_sg U52604 ( .A(n7088), .X(n46883) );
  inv_x1_sg U52605 ( .A(n7906), .X(n47176) );
  inv_x1_sg U52606 ( .A(n8724), .X(n47461) );
  inv_x1_sg U52607 ( .A(n9544), .X(n47746) );
  inv_x1_sg U52608 ( .A(n10363), .X(n48031) );
  inv_x1_sg U52609 ( .A(n11182), .X(n48316) );
  inv_x1_sg U52610 ( .A(n12001), .X(n48601) );
  inv_x1_sg U52611 ( .A(n12820), .X(n48887) );
  inv_x1_sg U52612 ( .A(n13639), .X(n49174) );
  inv_x1_sg U52613 ( .A(n14458), .X(n49460) );
  inv_x1_sg U52614 ( .A(n15277), .X(n49745) );
  inv_x1_sg U52615 ( .A(n16096), .X(n50032) );
  inv_x1_sg U52616 ( .A(n16914), .X(n50317) );
  inv_x1_sg U52617 ( .A(n17734), .X(n50606) );
  inv_x1_sg U52618 ( .A(n18555), .X(n50893) );
  inv_x1_sg U52619 ( .A(n17460), .X(n50521) );
  inv_x1_sg U52620 ( .A(n7635), .X(n47094) );
  inv_x1_sg U52621 ( .A(n8453), .X(n47380) );
  inv_x1_sg U52622 ( .A(n9271), .X(n47665) );
  inv_x1_sg U52623 ( .A(n10091), .X(n47950) );
  inv_x1_sg U52624 ( .A(n10910), .X(n48235) );
  inv_x1_sg U52625 ( .A(n11729), .X(n48520) );
  inv_x1_sg U52626 ( .A(n12548), .X(n48805) );
  inv_x1_sg U52627 ( .A(n13367), .X(n49092) );
  inv_x1_sg U52628 ( .A(n14186), .X(n49378) );
  inv_x1_sg U52629 ( .A(n15005), .X(n49664) );
  inv_x1_sg U52630 ( .A(n15824), .X(n49950) );
  inv_x1_sg U52631 ( .A(n16643), .X(n50236) );
  inv_x1_sg U52632 ( .A(n18281), .X(n50810) );
  inv_x1_sg U52633 ( .A(n19102), .X(n51097) );
  nand_x1_sg U52634 ( .A(n26307), .B(n50848), .X(n26306) );
  inv_x1_sg U52635 ( .A(n26308), .X(n50848) );
  inv_x1_sg U52636 ( .A(n7342), .X(n46992) );
  inv_x1_sg U52637 ( .A(n17167), .X(n50422) );
  inv_x1_sg U52638 ( .A(n8160), .X(n47281) );
  inv_x1_sg U52639 ( .A(n8978), .X(n47566) );
  inv_x1_sg U52640 ( .A(n9798), .X(n47851) );
  inv_x1_sg U52641 ( .A(n10617), .X(n48136) );
  inv_x1_sg U52642 ( .A(n11436), .X(n48421) );
  inv_x1_sg U52643 ( .A(n12255), .X(n48706) );
  inv_x1_sg U52644 ( .A(n13074), .X(n48992) );
  inv_x1_sg U52645 ( .A(n13893), .X(n49279) );
  inv_x1_sg U52646 ( .A(n14712), .X(n49565) );
  inv_x1_sg U52647 ( .A(n15531), .X(n49851) );
  inv_x1_sg U52648 ( .A(n16350), .X(n50137) );
  inv_x1_sg U52649 ( .A(n17988), .X(n50711) );
  inv_x1_sg U52650 ( .A(n18809), .X(n50998) );
  inv_x1_sg U52651 ( .A(n8407), .X(n47334) );
  inv_x1_sg U52652 ( .A(n9225), .X(n47619) );
  inv_x1_sg U52653 ( .A(n10045), .X(n47904) );
  inv_x1_sg U52654 ( .A(n10864), .X(n48189) );
  inv_x1_sg U52655 ( .A(n11683), .X(n48474) );
  inv_x1_sg U52656 ( .A(n12502), .X(n48759) );
  inv_x1_sg U52657 ( .A(n13321), .X(n49045) );
  inv_x1_sg U52658 ( .A(n14140), .X(n49332) );
  inv_x1_sg U52659 ( .A(n14959), .X(n49618) );
  inv_x1_sg U52660 ( .A(n15778), .X(n49904) );
  inv_x1_sg U52661 ( .A(n16597), .X(n50190) );
  inv_x1_sg U52662 ( .A(n18235), .X(n50764) );
  inv_x1_sg U52663 ( .A(n19056), .X(n51051) );
  inv_x1_sg U52664 ( .A(n7467), .X(n47034) );
  inv_x1_sg U52665 ( .A(n8285), .X(n47321) );
  inv_x1_sg U52666 ( .A(n9103), .X(n47606) );
  inv_x1_sg U52667 ( .A(n9923), .X(n47891) );
  inv_x1_sg U52668 ( .A(n10742), .X(n48176) );
  inv_x1_sg U52669 ( .A(n11561), .X(n48461) );
  inv_x1_sg U52670 ( .A(n12380), .X(n48746) );
  inv_x1_sg U52671 ( .A(n13199), .X(n49032) );
  inv_x1_sg U52672 ( .A(n14018), .X(n49319) );
  inv_x1_sg U52673 ( .A(n14837), .X(n49605) );
  inv_x1_sg U52674 ( .A(n15656), .X(n49891) );
  inv_x1_sg U52675 ( .A(n16475), .X(n50177) );
  inv_x1_sg U52676 ( .A(n18113), .X(n50751) );
  inv_x1_sg U52677 ( .A(n18934), .X(n51038) );
  inv_x1_sg U52678 ( .A(n17292), .X(n50462) );
  inv_x1_sg U52679 ( .A(n7098), .X(n46869) );
  inv_x1_sg U52680 ( .A(n7916), .X(n47162) );
  inv_x1_sg U52681 ( .A(n8734), .X(n47447) );
  inv_x1_sg U52682 ( .A(n9554), .X(n47732) );
  inv_x1_sg U52683 ( .A(n10373), .X(n48017) );
  inv_x1_sg U52684 ( .A(n11192), .X(n48302) );
  inv_x1_sg U52685 ( .A(n12011), .X(n48587) );
  inv_x1_sg U52686 ( .A(n12830), .X(n48873) );
  inv_x1_sg U52687 ( .A(n13649), .X(n49160) );
  inv_x1_sg U52688 ( .A(n14468), .X(n49446) );
  inv_x1_sg U52689 ( .A(n15287), .X(n49731) );
  inv_x1_sg U52690 ( .A(n16106), .X(n50018) );
  inv_x1_sg U52691 ( .A(n16923), .X(n50303) );
  inv_x1_sg U52692 ( .A(n17744), .X(n50592) );
  inv_x1_sg U52693 ( .A(n18565), .X(n50879) );
  inv_x1_sg U52694 ( .A(n16931), .X(n50316) );
  inv_x1_sg U52695 ( .A(n7289), .X(n46919) );
  inv_x1_sg U52696 ( .A(n8107), .X(n47211) );
  inv_x1_sg U52697 ( .A(n8925), .X(n47496) );
  inv_x1_sg U52698 ( .A(n9745), .X(n47781) );
  inv_x1_sg U52699 ( .A(n10564), .X(n48066) );
  inv_x1_sg U52700 ( .A(n11383), .X(n48351) );
  inv_x1_sg U52701 ( .A(n12202), .X(n48636) );
  inv_x1_sg U52702 ( .A(n13021), .X(n48922) );
  inv_x1_sg U52703 ( .A(n13840), .X(n49209) );
  inv_x1_sg U52704 ( .A(n14659), .X(n49495) );
  inv_x1_sg U52705 ( .A(n15478), .X(n49781) );
  inv_x1_sg U52706 ( .A(n16297), .X(n50067) );
  inv_x1_sg U52707 ( .A(n17935), .X(n50641) );
  inv_x1_sg U52708 ( .A(n18756), .X(n50928) );
  inv_x1_sg U52709 ( .A(n7106), .X(n46882) );
  inv_x1_sg U52710 ( .A(n7924), .X(n47175) );
  inv_x1_sg U52711 ( .A(n8742), .X(n47460) );
  inv_x1_sg U52712 ( .A(n9562), .X(n47745) );
  inv_x1_sg U52713 ( .A(n10381), .X(n48030) );
  inv_x1_sg U52714 ( .A(n11200), .X(n48315) );
  inv_x1_sg U52715 ( .A(n12019), .X(n48600) );
  inv_x1_sg U52716 ( .A(n12838), .X(n48886) );
  inv_x1_sg U52717 ( .A(n13657), .X(n49173) );
  inv_x1_sg U52718 ( .A(n14476), .X(n49459) );
  inv_x1_sg U52719 ( .A(n15295), .X(n49744) );
  inv_x1_sg U52720 ( .A(n16114), .X(n50031) );
  inv_x1_sg U52721 ( .A(n17752), .X(n50605) );
  inv_x1_sg U52722 ( .A(n18573), .X(n50892) );
  inv_x1_sg U52723 ( .A(n7270), .X(n46975) );
  inv_x1_sg U52724 ( .A(n17095), .X(n50406) );
  inv_x1_sg U52725 ( .A(n8089), .X(n47265) );
  inv_x1_sg U52726 ( .A(n8907), .X(n47550) );
  inv_x1_sg U52727 ( .A(n9727), .X(n47835) );
  inv_x1_sg U52728 ( .A(n10546), .X(n48120) );
  inv_x1_sg U52729 ( .A(n11365), .X(n48405) );
  inv_x1_sg U52730 ( .A(n12184), .X(n48690) );
  inv_x1_sg U52731 ( .A(n13003), .X(n48976) );
  inv_x1_sg U52732 ( .A(n13822), .X(n49263) );
  inv_x1_sg U52733 ( .A(n14641), .X(n49549) );
  inv_x1_sg U52734 ( .A(n15460), .X(n49835) );
  inv_x1_sg U52735 ( .A(n16279), .X(n50121) );
  inv_x1_sg U52736 ( .A(n17917), .X(n50695) );
  inv_x1_sg U52737 ( .A(n18738), .X(n50982) );
  inv_x1_sg U52738 ( .A(n7379), .X(n46967) );
  inv_x1_sg U52739 ( .A(n8197), .X(n47257) );
  inv_x1_sg U52740 ( .A(n9015), .X(n47542) );
  inv_x1_sg U52741 ( .A(n9835), .X(n47827) );
  inv_x1_sg U52742 ( .A(n10654), .X(n48112) );
  inv_x1_sg U52743 ( .A(n11473), .X(n48397) );
  inv_x1_sg U52744 ( .A(n12292), .X(n48682) );
  inv_x1_sg U52745 ( .A(n13111), .X(n48968) );
  inv_x1_sg U52746 ( .A(n13930), .X(n49255) );
  inv_x1_sg U52747 ( .A(n14749), .X(n49541) );
  inv_x1_sg U52748 ( .A(n15568), .X(n49827) );
  inv_x1_sg U52749 ( .A(n16387), .X(n50113) );
  inv_x1_sg U52750 ( .A(n18025), .X(n50687) );
  inv_x1_sg U52751 ( .A(n18846), .X(n50974) );
  inv_x1_sg U52752 ( .A(n7507), .X(n46981) );
  inv_x1_sg U52753 ( .A(n8325), .X(n47271) );
  inv_x1_sg U52754 ( .A(n9143), .X(n47556) );
  inv_x1_sg U52755 ( .A(n9963), .X(n47841) );
  inv_x1_sg U52756 ( .A(n10782), .X(n48126) );
  inv_x1_sg U52757 ( .A(n11601), .X(n48411) );
  inv_x1_sg U52758 ( .A(n12420), .X(n48696) );
  inv_x1_sg U52759 ( .A(n13239), .X(n48982) );
  inv_x1_sg U52760 ( .A(n14058), .X(n49269) );
  inv_x1_sg U52761 ( .A(n14877), .X(n49555) );
  inv_x1_sg U52762 ( .A(n15696), .X(n49841) );
  inv_x1_sg U52763 ( .A(n16515), .X(n50127) );
  inv_x1_sg U52764 ( .A(n17332), .X(n50412) );
  inv_x1_sg U52765 ( .A(n18153), .X(n50701) );
  inv_x1_sg U52766 ( .A(n18974), .X(n50988) );
  nand_x1_sg U52767 ( .A(n26588), .B(n51134), .X(n26587) );
  inv_x1_sg U52768 ( .A(n26589), .X(n51134) );
  nand_x1_sg U52769 ( .A(n22689), .B(n47131), .X(n22688) );
  inv_x1_sg U52770 ( .A(n22690), .X(n47131) );
  inv_x1_sg U52771 ( .A(n7495), .X(n47022) );
  inv_x1_sg U52772 ( .A(n7172), .X(n46951) );
  inv_x1_sg U52773 ( .A(n7991), .X(n47242) );
  inv_x1_sg U52774 ( .A(n8809), .X(n47527) );
  inv_x1_sg U52775 ( .A(n9629), .X(n47812) );
  inv_x1_sg U52776 ( .A(n10448), .X(n48097) );
  inv_x1_sg U52777 ( .A(n11267), .X(n48382) );
  inv_x1_sg U52778 ( .A(n12086), .X(n48667) );
  inv_x1_sg U52779 ( .A(n12905), .X(n48953) );
  inv_x1_sg U52780 ( .A(n13724), .X(n49240) );
  inv_x1_sg U52781 ( .A(n14543), .X(n49526) );
  inv_x1_sg U52782 ( .A(n15362), .X(n49812) );
  inv_x1_sg U52783 ( .A(n16181), .X(n50098) );
  inv_x1_sg U52784 ( .A(n17819), .X(n50672) );
  inv_x1_sg U52785 ( .A(n18640), .X(n50959) );
  inv_x1_sg U52786 ( .A(n7133), .X(n46874) );
  inv_x1_sg U52787 ( .A(n17779), .X(n50597) );
  inv_x1_sg U52788 ( .A(n8313), .X(n47310) );
  inv_x1_sg U52789 ( .A(n9131), .X(n47595) );
  inv_x1_sg U52790 ( .A(n9951), .X(n47880) );
  inv_x1_sg U52791 ( .A(n10770), .X(n48165) );
  inv_x1_sg U52792 ( .A(n11589), .X(n48450) );
  inv_x1_sg U52793 ( .A(n12408), .X(n48735) );
  inv_x1_sg U52794 ( .A(n13227), .X(n49021) );
  inv_x1_sg U52795 ( .A(n14046), .X(n49308) );
  inv_x1_sg U52796 ( .A(n14865), .X(n49594) );
  inv_x1_sg U52797 ( .A(n15684), .X(n49880) );
  inv_x1_sg U52798 ( .A(n16503), .X(n50166) );
  inv_x1_sg U52799 ( .A(n18141), .X(n50740) );
  inv_x1_sg U52800 ( .A(n18962), .X(n51027) );
  inv_x1_sg U52801 ( .A(n7226), .X(n46888) );
  inv_x1_sg U52802 ( .A(n17051), .X(n50322) );
  inv_x1_sg U52803 ( .A(n7951), .X(n47167) );
  inv_x1_sg U52804 ( .A(n8769), .X(n47452) );
  inv_x1_sg U52805 ( .A(n9589), .X(n47737) );
  inv_x1_sg U52806 ( .A(n10408), .X(n48022) );
  inv_x1_sg U52807 ( .A(n11227), .X(n48307) );
  inv_x1_sg U52808 ( .A(n12046), .X(n48592) );
  inv_x1_sg U52809 ( .A(n12865), .X(n48878) );
  inv_x1_sg U52810 ( .A(n13684), .X(n49165) );
  inv_x1_sg U52811 ( .A(n14503), .X(n49451) );
  inv_x1_sg U52812 ( .A(n15322), .X(n49736) );
  inv_x1_sg U52813 ( .A(n16141), .X(n50023) );
  inv_x1_sg U52814 ( .A(n16958), .X(n50308) );
  inv_x1_sg U52815 ( .A(n18600), .X(n50884) );
  inv_x1_sg U52816 ( .A(n8045), .X(n47181) );
  inv_x1_sg U52817 ( .A(n8863), .X(n47466) );
  inv_x1_sg U52818 ( .A(n9683), .X(n47751) );
  inv_x1_sg U52819 ( .A(n10502), .X(n48036) );
  inv_x1_sg U52820 ( .A(n11321), .X(n48321) );
  inv_x1_sg U52821 ( .A(n12140), .X(n48606) );
  inv_x1_sg U52822 ( .A(n12959), .X(n48892) );
  inv_x1_sg U52823 ( .A(n13778), .X(n49179) );
  inv_x1_sg U52824 ( .A(n14597), .X(n49465) );
  inv_x1_sg U52825 ( .A(n15416), .X(n49750) );
  inv_x1_sg U52826 ( .A(n16235), .X(n50037) );
  inv_x1_sg U52827 ( .A(n17873), .X(n50611) );
  inv_x1_sg U52828 ( .A(n18694), .X(n50898) );
  inv_x1_sg U52829 ( .A(n7628), .X(n47103) );
  inv_x1_sg U52830 ( .A(n8446), .X(n47389) );
  inv_x1_sg U52831 ( .A(n9264), .X(n47674) );
  inv_x1_sg U52832 ( .A(n10084), .X(n47959) );
  inv_x1_sg U52833 ( .A(n10903), .X(n48244) );
  inv_x1_sg U52834 ( .A(n11722), .X(n48529) );
  inv_x1_sg U52835 ( .A(n12541), .X(n48814) );
  inv_x1_sg U52836 ( .A(n13360), .X(n49101) );
  inv_x1_sg U52837 ( .A(n14179), .X(n49387) );
  inv_x1_sg U52838 ( .A(n14998), .X(n49673) );
  inv_x1_sg U52839 ( .A(n15817), .X(n49959) );
  inv_x1_sg U52840 ( .A(n16636), .X(n50245) );
  inv_x1_sg U52841 ( .A(n17453), .X(n50530) );
  inv_x1_sg U52842 ( .A(n18274), .X(n50819) );
  inv_x1_sg U52843 ( .A(n19095), .X(n51106) );
  inv_x1_sg U52844 ( .A(n7562), .X(n46960) );
  inv_x1_sg U52845 ( .A(n8380), .X(n47251) );
  inv_x1_sg U52846 ( .A(n9198), .X(n47536) );
  inv_x1_sg U52847 ( .A(n10018), .X(n47821) );
  inv_x1_sg U52848 ( .A(n10837), .X(n48106) );
  inv_x1_sg U52849 ( .A(n11656), .X(n48391) );
  inv_x1_sg U52850 ( .A(n12475), .X(n48676) );
  inv_x1_sg U52851 ( .A(n13294), .X(n48962) );
  inv_x1_sg U52852 ( .A(n14113), .X(n49249) );
  inv_x1_sg U52853 ( .A(n14932), .X(n49535) );
  inv_x1_sg U52854 ( .A(n15751), .X(n49821) );
  inv_x1_sg U52855 ( .A(n16570), .X(n50107) );
  inv_x1_sg U52856 ( .A(n18208), .X(n50681) );
  inv_x1_sg U52857 ( .A(n19029), .X(n50968) );
  inv_x1_sg U52858 ( .A(n17129), .X(n50376) );
  nand_x2_sg U52859 ( .A(n26756), .B(n26757), .X(n26755) );
  nand_x2_sg U52860 ( .A(n21769), .B(n21770), .X(n21768) );
  nand_x2_sg U52861 ( .A(n21909), .B(n21910), .X(n21908) );
  nand_x2_sg U52862 ( .A(n22049), .B(n22050), .X(n22048) );
  nand_x2_sg U52863 ( .A(n22190), .B(n22191), .X(n22189) );
  nand_x2_sg U52864 ( .A(n22333), .B(n22334), .X(n22332) );
  nand_x2_sg U52865 ( .A(n22474), .B(n22475), .X(n22473) );
  inv_x1_sg U52866 ( .A(n18259), .X(n50775) );
  inv_x1_sg U52867 ( .A(n8431), .X(n47345) );
  inv_x1_sg U52868 ( .A(n9249), .X(n47630) );
  inv_x1_sg U52869 ( .A(n10069), .X(n47915) );
  inv_x1_sg U52870 ( .A(n10888), .X(n48200) );
  inv_x1_sg U52871 ( .A(n11707), .X(n48485) );
  inv_x1_sg U52872 ( .A(n12526), .X(n48770) );
  inv_x1_sg U52873 ( .A(n13345), .X(n49057) );
  inv_x1_sg U52874 ( .A(n14164), .X(n49343) );
  inv_x1_sg U52875 ( .A(n14983), .X(n49629) );
  inv_x1_sg U52876 ( .A(n15802), .X(n49915) );
  inv_x1_sg U52877 ( .A(n16621), .X(n50201) );
  inv_x1_sg U52878 ( .A(n19080), .X(n51062) );
  inv_x1_sg U52879 ( .A(n7433), .X(n46935) );
  inv_x1_sg U52880 ( .A(n8251), .X(n47227) );
  inv_x1_sg U52881 ( .A(n9069), .X(n47512) );
  inv_x1_sg U52882 ( .A(n9889), .X(n47797) );
  inv_x1_sg U52883 ( .A(n10708), .X(n48082) );
  inv_x1_sg U52884 ( .A(n11527), .X(n48367) );
  inv_x1_sg U52885 ( .A(n12346), .X(n48652) );
  inv_x1_sg U52886 ( .A(n13165), .X(n48938) );
  inv_x1_sg U52887 ( .A(n13984), .X(n49225) );
  inv_x1_sg U52888 ( .A(n14803), .X(n49511) );
  inv_x1_sg U52889 ( .A(n15622), .X(n49797) );
  inv_x1_sg U52890 ( .A(n16441), .X(n50083) );
  inv_x1_sg U52891 ( .A(n18079), .X(n50657) );
  inv_x1_sg U52892 ( .A(n18900), .X(n50944) );
  nand_x2_sg U52893 ( .A(n21722), .B(n21723), .X(n21721) );
  nand_x2_sg U52894 ( .A(n21863), .B(n21864), .X(n21862) );
  nand_x2_sg U52895 ( .A(n22002), .B(n22003), .X(n22001) );
  nand_x2_sg U52896 ( .A(n22143), .B(n22144), .X(n22142) );
  nand_x2_sg U52897 ( .A(n22285), .B(n22286), .X(n22284) );
  nand_x2_sg U52898 ( .A(n22428), .B(n22429), .X(n22427) );
  nand_x2_sg U52899 ( .A(n21816), .B(n21817), .X(n21815) );
  nand_x2_sg U52900 ( .A(n21956), .B(n21957), .X(n21955) );
  nand_x2_sg U52901 ( .A(n22095), .B(n22096), .X(n22094) );
  nand_x2_sg U52902 ( .A(n22238), .B(n22239), .X(n22237) );
  nand_x2_sg U52903 ( .A(n22380), .B(n22381), .X(n22379) );
  nand_x2_sg U52904 ( .A(n22520), .B(n22521), .X(n22519) );
  inv_x1_sg U52905 ( .A(n17320), .X(n50451) );
  inv_x1_sg U52906 ( .A(n7258), .X(n46933) );
  inv_x1_sg U52907 ( .A(n17905), .X(n50655) );
  inv_x1_sg U52908 ( .A(n8077), .X(n47225) );
  inv_x1_sg U52909 ( .A(n8895), .X(n47510) );
  inv_x1_sg U52910 ( .A(n9715), .X(n47795) );
  inv_x1_sg U52911 ( .A(n10534), .X(n48080) );
  inv_x1_sg U52912 ( .A(n11353), .X(n48365) );
  inv_x1_sg U52913 ( .A(n12172), .X(n48650) );
  inv_x1_sg U52914 ( .A(n12991), .X(n48936) );
  inv_x1_sg U52915 ( .A(n13810), .X(n49223) );
  inv_x1_sg U52916 ( .A(n14629), .X(n49509) );
  inv_x1_sg U52917 ( .A(n15448), .X(n49795) );
  inv_x1_sg U52918 ( .A(n16267), .X(n50081) );
  inv_x1_sg U52919 ( .A(n17083), .X(n50366) );
  inv_x1_sg U52920 ( .A(n18726), .X(n50942) );
  nand_x1_sg U52921 ( .A(n23520), .B(n47987), .X(n23519) );
  inv_x1_sg U52922 ( .A(n23521), .X(n47987) );
  nand_x1_sg U52923 ( .A(n23799), .B(n48272), .X(n23798) );
  inv_x1_sg U52924 ( .A(n23800), .X(n48272) );
  nand_x1_sg U52925 ( .A(n22963), .B(n47417), .X(n22962) );
  inv_x1_sg U52926 ( .A(n22964), .X(n47417) );
  nand_x1_sg U52927 ( .A(n23240), .B(n47702), .X(n23239) );
  inv_x1_sg U52928 ( .A(n23241), .X(n47702) );
  nand_x1_sg U52929 ( .A(n24078), .B(n48557), .X(n24077) );
  inv_x1_sg U52930 ( .A(n24079), .X(n48557) );
  nand_x1_sg U52931 ( .A(n24357), .B(n48842), .X(n24356) );
  inv_x1_sg U52932 ( .A(n24358), .X(n48842) );
  nand_x1_sg U52933 ( .A(n24914), .B(n49415), .X(n24913) );
  inv_x1_sg U52934 ( .A(n24915), .X(n49415) );
  nand_x1_sg U52935 ( .A(n25193), .B(n49701), .X(n25192) );
  inv_x1_sg U52936 ( .A(n25194), .X(n49701) );
  nand_x1_sg U52937 ( .A(n25472), .B(n49987), .X(n25471) );
  inv_x1_sg U52938 ( .A(n25473), .X(n49987) );
  nand_x1_sg U52939 ( .A(n25751), .B(n50273), .X(n25750) );
  inv_x1_sg U52940 ( .A(n25752), .X(n50273) );
  nand_x1_sg U52941 ( .A(n24636), .B(n49129), .X(n24635) );
  inv_x1_sg U52942 ( .A(n24637), .X(n49129) );
  inv_x1_sg U52943 ( .A(n7076), .X(n46859) );
  inv_x1_sg U52944 ( .A(n7894), .X(n47152) );
  inv_x1_sg U52945 ( .A(n8712), .X(n47437) );
  inv_x1_sg U52946 ( .A(n9532), .X(n47722) );
  inv_x1_sg U52947 ( .A(n10351), .X(n48007) );
  inv_x1_sg U52948 ( .A(n11170), .X(n48292) );
  inv_x1_sg U52949 ( .A(n11989), .X(n48577) );
  inv_x1_sg U52950 ( .A(n12808), .X(n48863) );
  inv_x1_sg U52951 ( .A(n13627), .X(n49150) );
  inv_x1_sg U52952 ( .A(n14446), .X(n49436) );
  inv_x1_sg U52953 ( .A(n15265), .X(n49721) );
  inv_x1_sg U52954 ( .A(n16084), .X(n50008) );
  inv_x1_sg U52955 ( .A(n17722), .X(n50582) );
  inv_x1_sg U52956 ( .A(n18543), .X(n50869) );
  inv_x1_sg U52957 ( .A(n16903), .X(n50292) );
  inv_x1_sg U52958 ( .A(n7158), .X(n46880) );
  inv_x1_sg U52959 ( .A(n17805), .X(n50603) );
  inv_x1_sg U52960 ( .A(n7977), .X(n47173) );
  inv_x1_sg U52961 ( .A(n8795), .X(n47458) );
  inv_x1_sg U52962 ( .A(n9615), .X(n47743) );
  inv_x1_sg U52963 ( .A(n10434), .X(n48028) );
  inv_x1_sg U52964 ( .A(n11253), .X(n48313) );
  inv_x1_sg U52965 ( .A(n12072), .X(n48598) );
  inv_x1_sg U52966 ( .A(n12891), .X(n48884) );
  inv_x1_sg U52967 ( .A(n13710), .X(n49171) );
  inv_x1_sg U52968 ( .A(n14529), .X(n49457) );
  inv_x1_sg U52969 ( .A(n15348), .X(n49742) );
  inv_x1_sg U52970 ( .A(n16167), .X(n50029) );
  inv_x1_sg U52971 ( .A(n16983), .X(n50314) );
  inv_x1_sg U52972 ( .A(n18626), .X(n50890) );
  inv_x1_sg U52973 ( .A(n7617), .X(n47053) );
  inv_x1_sg U52974 ( .A(n8435), .X(n47340) );
  inv_x1_sg U52975 ( .A(n9253), .X(n47625) );
  inv_x1_sg U52976 ( .A(n10073), .X(n47910) );
  inv_x1_sg U52977 ( .A(n10892), .X(n48195) );
  inv_x1_sg U52978 ( .A(n11711), .X(n48480) );
  inv_x1_sg U52979 ( .A(n12530), .X(n48765) );
  inv_x1_sg U52980 ( .A(n13349), .X(n49051) );
  inv_x1_sg U52981 ( .A(n14168), .X(n49338) );
  inv_x1_sg U52982 ( .A(n14987), .X(n49624) );
  inv_x1_sg U52983 ( .A(n15806), .X(n49910) );
  inv_x1_sg U52984 ( .A(n16625), .X(n50196) );
  inv_x1_sg U52985 ( .A(n18263), .X(n50770) );
  inv_x1_sg U52986 ( .A(n19084), .X(n51057) );
  inv_x1_sg U52987 ( .A(n16848), .X(n50489) );
  inv_x1_sg U52988 ( .A(n17442), .X(n50481) );
  nand_x1_sg U52989 ( .A(n26015), .B(n50561), .X(n26014) );
  inv_x1_sg U52990 ( .A(n26016), .X(n50561) );
  inv_x1_sg U52991 ( .A(n8131), .X(n47302) );
  inv_x1_sg U52992 ( .A(n8949), .X(n47587) );
  inv_x1_sg U52993 ( .A(n9769), .X(n47872) );
  inv_x1_sg U52994 ( .A(n10588), .X(n48157) );
  inv_x1_sg U52995 ( .A(n11407), .X(n48442) );
  inv_x1_sg U52996 ( .A(n12226), .X(n48727) );
  inv_x1_sg U52997 ( .A(n13045), .X(n49013) );
  inv_x1_sg U52998 ( .A(n13864), .X(n49300) );
  inv_x1_sg U52999 ( .A(n14683), .X(n49586) );
  inv_x1_sg U53000 ( .A(n15502), .X(n49872) );
  inv_x1_sg U53001 ( .A(n16321), .X(n50158) );
  inv_x1_sg U53002 ( .A(n17959), .X(n50732) );
  inv_x1_sg U53003 ( .A(n18780), .X(n51019) );
  inv_x1_sg U53004 ( .A(n7479), .X(n47064) );
  inv_x1_sg U53005 ( .A(n8297), .X(n47350) );
  inv_x1_sg U53006 ( .A(n9115), .X(n47635) );
  inv_x1_sg U53007 ( .A(n9935), .X(n47920) );
  inv_x1_sg U53008 ( .A(n10754), .X(n48205) );
  inv_x1_sg U53009 ( .A(n11573), .X(n48490) );
  inv_x1_sg U53010 ( .A(n12392), .X(n48775) );
  inv_x1_sg U53011 ( .A(n13211), .X(n49062) );
  inv_x1_sg U53012 ( .A(n14030), .X(n49348) );
  inv_x1_sg U53013 ( .A(n14849), .X(n49634) );
  inv_x1_sg U53014 ( .A(n15668), .X(n49920) );
  inv_x1_sg U53015 ( .A(n16487), .X(n50206) );
  inv_x1_sg U53016 ( .A(n17304), .X(n50491) );
  inv_x1_sg U53017 ( .A(n18125), .X(n50780) );
  inv_x1_sg U53018 ( .A(n18946), .X(n51067) );
  inv_x1_sg U53019 ( .A(n7492), .X(n46955) );
  inv_x1_sg U53020 ( .A(n8310), .X(n47246) );
  inv_x1_sg U53021 ( .A(n9128), .X(n47531) );
  inv_x1_sg U53022 ( .A(n9948), .X(n47816) );
  inv_x1_sg U53023 ( .A(n10767), .X(n48101) );
  inv_x1_sg U53024 ( .A(n11586), .X(n48386) );
  inv_x1_sg U53025 ( .A(n12405), .X(n48671) );
  inv_x1_sg U53026 ( .A(n13224), .X(n48957) );
  inv_x1_sg U53027 ( .A(n14043), .X(n49244) );
  inv_x1_sg U53028 ( .A(n14862), .X(n49530) );
  inv_x1_sg U53029 ( .A(n15681), .X(n49816) );
  inv_x1_sg U53030 ( .A(n16500), .X(n50102) );
  inv_x1_sg U53031 ( .A(n18138), .X(n50676) );
  inv_x1_sg U53032 ( .A(n18959), .X(n50963) );
  inv_x1_sg U53033 ( .A(n26758), .X(n51509) );
  inv_x1_sg U53034 ( .A(n21724), .X(n51490) );
  inv_x1_sg U53035 ( .A(n21771), .X(n51491) );
  inv_x1_sg U53036 ( .A(n21818), .X(n51492) );
  inv_x1_sg U53037 ( .A(n21865), .X(n51493) );
  inv_x1_sg U53038 ( .A(n21911), .X(n51494) );
  inv_x1_sg U53039 ( .A(n21958), .X(n51495) );
  inv_x1_sg U53040 ( .A(n22004), .X(n51496) );
  inv_x1_sg U53041 ( .A(n22051), .X(n51497) );
  inv_x1_sg U53042 ( .A(n22097), .X(n51498) );
  inv_x1_sg U53043 ( .A(n22145), .X(n51499) );
  inv_x1_sg U53044 ( .A(n22192), .X(n51500) );
  inv_x1_sg U53045 ( .A(n22240), .X(n51501) );
  inv_x1_sg U53046 ( .A(n22287), .X(n51502) );
  inv_x1_sg U53047 ( .A(n22335), .X(n51503) );
  inv_x1_sg U53048 ( .A(n22382), .X(n51504) );
  inv_x1_sg U53049 ( .A(n22430), .X(n51505) );
  inv_x1_sg U53050 ( .A(n22476), .X(n51506) );
  inv_x1_sg U53051 ( .A(n22522), .X(n51507) );
  inv_x1_sg U53052 ( .A(n22558), .X(n51508) );
  nand_x1_sg U53053 ( .A(n17078), .B(n17077), .X(n17079) );
  inv_x1_sg U53054 ( .A(n5752), .X(n51458) );
  inv_x1_sg U53055 ( .A(n5759), .X(n51460) );
  inv_x1_sg U53056 ( .A(n5732), .X(n51452) );
  inv_x1_sg U53057 ( .A(n5737), .X(n51454) );
  inv_x1_sg U53058 ( .A(n5748), .X(n51456) );
  inv_x1_sg U53059 ( .A(n25955), .X(n51465) );
  inv_x1_sg U53060 ( .A(n25962), .X(n51466) );
  inv_x1_sg U53061 ( .A(n5767), .X(n51464) );
  inv_x1_sg U53062 ( .A(n25988), .X(n51468) );
  inv_x1_sg U53063 ( .A(n26001), .X(n51469) );
  inv_x1_sg U53064 ( .A(n5763), .X(n51462) );
  inv_x1_sg U53065 ( .A(n5735), .X(n51453) );
  inv_x1_sg U53066 ( .A(n5740), .X(n51455) );
  inv_x1_sg U53067 ( .A(n5756), .X(n51459) );
  inv_x1_sg U53068 ( .A(n5750), .X(n51457) );
  inv_x1_sg U53069 ( .A(n5761), .X(n51461) );
  inv_x1_sg U53070 ( .A(n5765), .X(n51463) );
  nand_x1_sg U53071 ( .A(n40586), .B(n39129), .X(n7639) );
  inv_x1_sg U53072 ( .A(n8141), .X(n47284) );
  inv_x1_sg U53073 ( .A(n8959), .X(n47569) );
  inv_x1_sg U53074 ( .A(n9779), .X(n47854) );
  inv_x1_sg U53075 ( .A(n10598), .X(n48139) );
  inv_x1_sg U53076 ( .A(n11417), .X(n48424) );
  inv_x1_sg U53077 ( .A(n12236), .X(n48709) );
  inv_x1_sg U53078 ( .A(n13055), .X(n48995) );
  inv_x1_sg U53079 ( .A(n13874), .X(n49282) );
  inv_x1_sg U53080 ( .A(n14693), .X(n49568) );
  inv_x1_sg U53081 ( .A(n15512), .X(n49854) );
  inv_x1_sg U53082 ( .A(n16331), .X(n50140) );
  inv_x1_sg U53083 ( .A(n17969), .X(n50714) );
  inv_x1_sg U53084 ( .A(n18790), .X(n51001) );
  inv_x1_sg U53085 ( .A(n8059), .X(n47244) );
  inv_x1_sg U53086 ( .A(n8877), .X(n47529) );
  inv_x1_sg U53087 ( .A(n9697), .X(n47814) );
  inv_x1_sg U53088 ( .A(n10516), .X(n48099) );
  inv_x1_sg U53089 ( .A(n11335), .X(n48384) );
  inv_x1_sg U53090 ( .A(n12154), .X(n48669) );
  inv_x1_sg U53091 ( .A(n12973), .X(n48955) );
  inv_x1_sg U53092 ( .A(n13792), .X(n49242) );
  inv_x1_sg U53093 ( .A(n14611), .X(n49528) );
  inv_x1_sg U53094 ( .A(n15430), .X(n49814) );
  inv_x1_sg U53095 ( .A(n16249), .X(n50100) );
  inv_x1_sg U53096 ( .A(n17887), .X(n50674) );
  inv_x1_sg U53097 ( .A(n18708), .X(n50961) );
  inv_x1_sg U53098 ( .A(n7240), .X(n46953) );
  inv_x1_sg U53099 ( .A(n17065), .X(n50385) );
  inv_x1_sg U53100 ( .A(n7527), .X(n47063) );
  inv_x1_sg U53101 ( .A(n8345), .X(n47349) );
  inv_x1_sg U53102 ( .A(n9163), .X(n47634) );
  inv_x1_sg U53103 ( .A(n9983), .X(n47919) );
  inv_x1_sg U53104 ( .A(n10802), .X(n48204) );
  inv_x1_sg U53105 ( .A(n11621), .X(n48489) );
  inv_x1_sg U53106 ( .A(n12440), .X(n48774) );
  inv_x1_sg U53107 ( .A(n13259), .X(n49061) );
  inv_x1_sg U53108 ( .A(n14078), .X(n49347) );
  inv_x1_sg U53109 ( .A(n14897), .X(n49633) );
  inv_x1_sg U53110 ( .A(n15716), .X(n49919) );
  inv_x1_sg U53111 ( .A(n16535), .X(n50205) );
  inv_x1_sg U53112 ( .A(n17352), .X(n50490) );
  inv_x1_sg U53113 ( .A(n18173), .X(n50779) );
  inv_x1_sg U53114 ( .A(n18994), .X(n51066) );
  inv_x1_sg U53115 ( .A(n7128), .X(n46881) );
  inv_x1_sg U53116 ( .A(n7946), .X(n47174) );
  inv_x1_sg U53117 ( .A(n8764), .X(n47459) );
  inv_x1_sg U53118 ( .A(n9584), .X(n47744) );
  inv_x1_sg U53119 ( .A(n10403), .X(n48029) );
  inv_x1_sg U53120 ( .A(n11222), .X(n48314) );
  inv_x1_sg U53121 ( .A(n12041), .X(n48599) );
  inv_x1_sg U53122 ( .A(n12860), .X(n48885) );
  inv_x1_sg U53123 ( .A(n13679), .X(n49172) );
  inv_x1_sg U53124 ( .A(n14498), .X(n49458) );
  inv_x1_sg U53125 ( .A(n15317), .X(n49743) );
  inv_x1_sg U53126 ( .A(n16136), .X(n50030) );
  inv_x1_sg U53127 ( .A(n16953), .X(n50315) );
  inv_x1_sg U53128 ( .A(n17774), .X(n50604) );
  inv_x1_sg U53129 ( .A(n18595), .X(n50891) );
  inv_x1_sg U53130 ( .A(n17456), .X(n50527) );
  inv_x1_sg U53131 ( .A(n7631), .X(n47100) );
  inv_x1_sg U53132 ( .A(n8449), .X(n47386) );
  inv_x1_sg U53133 ( .A(n9267), .X(n47671) );
  inv_x1_sg U53134 ( .A(n10087), .X(n47956) );
  inv_x1_sg U53135 ( .A(n10906), .X(n48241) );
  inv_x1_sg U53136 ( .A(n11725), .X(n48526) );
  inv_x1_sg U53137 ( .A(n12544), .X(n48811) );
  inv_x1_sg U53138 ( .A(n13363), .X(n49098) );
  inv_x1_sg U53139 ( .A(n14182), .X(n49384) );
  inv_x1_sg U53140 ( .A(n15001), .X(n49670) );
  inv_x1_sg U53141 ( .A(n15820), .X(n49956) );
  inv_x1_sg U53142 ( .A(n16639), .X(n50242) );
  inv_x1_sg U53143 ( .A(n18277), .X(n50816) );
  inv_x1_sg U53144 ( .A(n19098), .X(n51103) );
  inv_x1_sg U53145 ( .A(n21160), .X(n46505) );
  inv_x1_sg U53146 ( .A(n21154), .X(n46468) );
  inv_x1_sg U53147 ( .A(n21148), .X(n46421) );
  inv_x1_sg U53148 ( .A(n21136), .X(n46332) );
  inv_x1_sg U53149 ( .A(n21142), .X(n46373) );
  inv_x1_sg U53150 ( .A(n21130), .X(n46286) );
  inv_x1_sg U53151 ( .A(n21124), .X(n46241) );
  inv_x1_sg U53152 ( .A(n21118), .X(n46195) );
  inv_x1_sg U53153 ( .A(n21112), .X(n46150) );
  inv_x1_sg U53154 ( .A(n21106), .X(n46104) );
  inv_x1_sg U53155 ( .A(n21100), .X(n46059) );
  inv_x1_sg U53156 ( .A(n21094), .X(n46013) );
  inv_x1_sg U53157 ( .A(n21088), .X(n45968) );
  inv_x1_sg U53158 ( .A(n20427), .X(n46335) );
  inv_x1_sg U53159 ( .A(n20379), .X(n45971) );
  inv_x1_sg U53160 ( .A(n20421), .X(n46289) );
  inv_x1_sg U53161 ( .A(n20415), .X(n46244) );
  inv_x1_sg U53162 ( .A(n20409), .X(n46198) );
  inv_x1_sg U53163 ( .A(n20403), .X(n46153) );
  inv_x1_sg U53164 ( .A(n20397), .X(n46107) );
  inv_x1_sg U53165 ( .A(n20391), .X(n46062) );
  inv_x1_sg U53166 ( .A(n20385), .X(n46016) );
  inv_x1_sg U53167 ( .A(n19694), .X(n46338) );
  inv_x1_sg U53168 ( .A(n19688), .X(n46292) );
  inv_x1_sg U53169 ( .A(n19682), .X(n46247) );
  inv_x1_sg U53170 ( .A(n19676), .X(n46201) );
  inv_x1_sg U53171 ( .A(n19670), .X(n46156) );
  inv_x1_sg U53172 ( .A(n19664), .X(n46110) );
  inv_x1_sg U53173 ( .A(n19658), .X(n46065) );
  inv_x1_sg U53174 ( .A(n19652), .X(n46019) );
  inv_x1_sg U53175 ( .A(n19646), .X(n45974) );
  inv_x1_sg U53176 ( .A(n7298), .X(n46974) );
  inv_x1_sg U53177 ( .A(n8116), .X(n47264) );
  inv_x1_sg U53178 ( .A(n8934), .X(n47549) );
  inv_x1_sg U53179 ( .A(n9754), .X(n47834) );
  inv_x1_sg U53180 ( .A(n10573), .X(n48119) );
  inv_x1_sg U53181 ( .A(n11392), .X(n48404) );
  inv_x1_sg U53182 ( .A(n12211), .X(n48689) );
  inv_x1_sg U53183 ( .A(n13030), .X(n48975) );
  inv_x1_sg U53184 ( .A(n13849), .X(n49262) );
  inv_x1_sg U53185 ( .A(n14668), .X(n49548) );
  inv_x1_sg U53186 ( .A(n15487), .X(n49834) );
  inv_x1_sg U53187 ( .A(n16306), .X(n50120) );
  inv_x1_sg U53188 ( .A(n17123), .X(n50405) );
  inv_x1_sg U53189 ( .A(n17944), .X(n50694) );
  inv_x1_sg U53190 ( .A(n18765), .X(n50981) );
  inv_x1_sg U53191 ( .A(n7471), .X(n47033) );
  inv_x1_sg U53192 ( .A(n17296), .X(n50461) );
  inv_x1_sg U53193 ( .A(n8289), .X(n47320) );
  inv_x1_sg U53194 ( .A(n9107), .X(n47605) );
  inv_x1_sg U53195 ( .A(n9927), .X(n47890) );
  inv_x1_sg U53196 ( .A(n10746), .X(n48175) );
  inv_x1_sg U53197 ( .A(n11565), .X(n48460) );
  inv_x1_sg U53198 ( .A(n12384), .X(n48745) );
  inv_x1_sg U53199 ( .A(n13203), .X(n49031) );
  inv_x1_sg U53200 ( .A(n14022), .X(n49318) );
  inv_x1_sg U53201 ( .A(n14841), .X(n49604) );
  inv_x1_sg U53202 ( .A(n15660), .X(n49890) );
  inv_x1_sg U53203 ( .A(n16479), .X(n50176) );
  inv_x1_sg U53204 ( .A(n18117), .X(n50750) );
  inv_x1_sg U53205 ( .A(n18938), .X(n51037) );
  nand_x2_sg U53206 ( .A(n17327), .B(n17298), .X(n17326) );
  nand_x2_sg U53207 ( .A(n7502), .B(n7473), .X(n7501) );
  nand_x2_sg U53208 ( .A(n8320), .B(n8291), .X(n8319) );
  nand_x2_sg U53209 ( .A(n9138), .B(n9109), .X(n9137) );
  nand_x2_sg U53210 ( .A(n9958), .B(n9929), .X(n9957) );
  nand_x2_sg U53211 ( .A(n10777), .B(n10748), .X(n10776) );
  nand_x2_sg U53212 ( .A(n11596), .B(n11567), .X(n11595) );
  nand_x2_sg U53213 ( .A(n12415), .B(n12386), .X(n12414) );
  nand_x2_sg U53214 ( .A(n13234), .B(n13205), .X(n13233) );
  nand_x2_sg U53215 ( .A(n14053), .B(n14024), .X(n14052) );
  nand_x2_sg U53216 ( .A(n14872), .B(n14843), .X(n14871) );
  nand_x2_sg U53217 ( .A(n15691), .B(n15662), .X(n15690) );
  nand_x2_sg U53218 ( .A(n16510), .B(n16481), .X(n16509) );
  nand_x2_sg U53219 ( .A(n18148), .B(n18119), .X(n18147) );
  nand_x2_sg U53220 ( .A(n18969), .B(n18940), .X(n18968) );
  nand_x2_sg U53221 ( .A(n22556), .B(n22557), .X(n22555) );
  nand_x1_sg U53222 ( .A(n39256), .B(n28519), .X(n28518) );
  inv_x1_sg U53223 ( .A(n23254), .X(n47703) );
  inv_x1_sg U53224 ( .A(n5769), .X(n51510) );
  inv_x1_sg U53225 ( .A(n5787), .X(n51514) );
  inv_x1_sg U53226 ( .A(n5864), .X(n51522) );
  inv_x1_sg U53227 ( .A(n5841), .X(n51520) );
  inv_x1_sg U53228 ( .A(n5826), .X(n51516) );
  inv_x1_sg U53229 ( .A(n5774), .X(n51512) );
  inv_x1_sg U53230 ( .A(n5882), .X(n51524) );
  inv_x1_sg U53231 ( .A(n5830), .X(n51518) );
  inv_x1_sg U53232 ( .A(n22705), .X(n51528) );
  inv_x1_sg U53233 ( .A(n5912), .X(n51525) );
  inv_x1_sg U53234 ( .A(n5772), .X(n51511) );
  inv_x1_sg U53235 ( .A(n22632), .X(n51527) );
  inv_x1_sg U53236 ( .A(n5873), .X(n51523) );
  inv_x1_sg U53237 ( .A(n5828), .X(n51517) );
  inv_x1_sg U53238 ( .A(n5776), .X(n51513) );
  inv_x1_sg U53239 ( .A(n5862), .X(n51521) );
  inv_x1_sg U53240 ( .A(n5832), .X(n51519) );
  inv_x1_sg U53241 ( .A(n5796), .X(n51515) );
  nand_x1_sg U53242 ( .A(n6832), .B(n6833), .X(n6830) );
  nand_x1_sg U53243 ( .A(n17477), .B(n17478), .X(n17476) );
  nand_x1_sg U53244 ( .A(n7649), .B(n7650), .X(n7648) );
  nand_x1_sg U53245 ( .A(n8467), .B(n8468), .X(n8466) );
  nand_x1_sg U53246 ( .A(n9287), .B(n9288), .X(n9286) );
  nand_x1_sg U53247 ( .A(n10106), .B(n10107), .X(n10105) );
  nand_x1_sg U53248 ( .A(n10925), .B(n10926), .X(n10924) );
  nand_x1_sg U53249 ( .A(n11744), .B(n11745), .X(n11743) );
  nand_x1_sg U53250 ( .A(n12563), .B(n12564), .X(n12562) );
  nand_x1_sg U53251 ( .A(n13382), .B(n13383), .X(n13381) );
  nand_x1_sg U53252 ( .A(n14201), .B(n14202), .X(n14200) );
  nand_x1_sg U53253 ( .A(n15020), .B(n15021), .X(n15019) );
  nand_x1_sg U53254 ( .A(n15839), .B(n15840), .X(n15838) );
  nand_x1_sg U53255 ( .A(n16656), .B(n16657), .X(n16654) );
  nand_x1_sg U53256 ( .A(n18298), .B(n18299), .X(n18297) );
  inv_x1_sg U53257 ( .A(n24781), .X(n48856) );
  inv_x1_sg U53258 ( .A(n25060), .X(n49143) );
  inv_x1_sg U53259 ( .A(n25339), .X(n49429) );
  inv_x1_sg U53260 ( .A(n25895), .X(n50001) );
  inv_x1_sg U53261 ( .A(n26733), .X(n50862) );
  inv_x1_sg U53262 ( .A(n26118), .X(n50281) );
  inv_x1_sg U53263 ( .A(n26473), .X(n50564) );
  inv_x1_sg U53264 ( .A(n22847), .X(n46844) );
  inv_x1_sg U53265 ( .A(n20953), .X(n46550) );
  inv_x1_sg U53266 ( .A(n26108), .X(n50291) );
  inv_x1_sg U53267 ( .A(n23275), .X(n47691) );
  inv_x1_sg U53268 ( .A(n22995), .X(n47406) );
  inv_x1_sg U53269 ( .A(n23554), .X(n47976) );
  inv_x1_sg U53270 ( .A(n23833), .X(n48261) );
  inv_x1_sg U53271 ( .A(n24112), .X(n48546) );
  inv_x1_sg U53272 ( .A(n24391), .X(n48831) );
  inv_x1_sg U53273 ( .A(n24669), .X(n49118) );
  inv_x1_sg U53274 ( .A(n24948), .X(n49404) );
  inv_x1_sg U53275 ( .A(n25227), .X(n49690) );
  inv_x1_sg U53276 ( .A(n25506), .X(n49976) );
  inv_x1_sg U53277 ( .A(n25783), .X(n50262) );
  inv_x1_sg U53278 ( .A(n26343), .X(n50836) );
  inv_x1_sg U53279 ( .A(n26621), .X(n51123) );
  inv_x1_sg U53280 ( .A(n20105), .X(n46381) );
  inv_x1_sg U53281 ( .A(n20779), .X(n46594) );
  inv_x1_sg U53282 ( .A(n19700), .X(n46383) );
  nand_x1_sg U53283 ( .A(n19168), .B(n38200), .X(n19167) );
  nand_x1_sg U53284 ( .A(n20164), .B(n38218), .X(n20163) );
  nand_x1_sg U53285 ( .A(n19582), .B(n38438), .X(n19581) );
  inv_x1_sg U53286 ( .A(n28263), .X(n45036) );
  nand_x1_sg U53287 ( .A(n19159), .B(n38440), .X(n19158) );
  inv_x1_sg U53288 ( .A(n25584), .X(n49754) );
  inv_x1_sg U53289 ( .A(n19226), .X(n45883) );
  inv_x1_sg U53290 ( .A(n21530), .X(n46504) );
  inv_x1_sg U53291 ( .A(n21348), .X(n46546) );
  nand_x1_sg U53292 ( .A(n20600), .B(n38199), .X(n20599) );
  nand_x1_sg U53293 ( .A(n20795), .B(n38217), .X(n20794) );
  nand_x1_sg U53294 ( .A(n19589), .B(n38260), .X(n19588) );
  inv_x1_sg U53295 ( .A(n19919), .X(n46519) );
  inv_x1_sg U53296 ( .A(n19725), .X(n46568) );
  inv_x1_sg U53297 ( .A(n20290), .X(n46428) );
  inv_x1_sg U53298 ( .A(n20453), .X(n46352) );
  inv_x1_sg U53299 ( .A(n21439), .X(n45874) );
  inv_x1_sg U53300 ( .A(n20670), .X(n45877) );
  inv_x1_sg U53301 ( .A(n20030), .X(n45880) );
  inv_x1_sg U53302 ( .A(n21178), .X(n46586) );
  inv_x1_sg U53303 ( .A(n28317), .X(n45443) );
  inv_x1_sg U53304 ( .A(n28188), .X(n45488) );
  inv_x1_sg U53305 ( .A(n28053), .X(n45532) );
  inv_x1_sg U53306 ( .A(n27891), .X(n45577) );
  inv_x1_sg U53307 ( .A(n27714), .X(n45621) );
  inv_x1_sg U53308 ( .A(n27520), .X(n45665) );
  inv_x1_sg U53309 ( .A(n27307), .X(n45709) );
  nand_x1_sg U53310 ( .A(n26842), .B(n38396), .X(n26841) );
  nand_x1_sg U53311 ( .A(n26857), .B(n38412), .X(n26856) );
  nand_x1_sg U53312 ( .A(n26864), .B(n38420), .X(n26863) );
  nand_x1_sg U53313 ( .A(n26871), .B(n38427), .X(n26870) );
  nand_x1_sg U53314 ( .A(n28562), .B(n38430), .X(n28561) );
  nand_x1_sg U53315 ( .A(n26878), .B(n38433), .X(n26877) );
  nand_x1_sg U53316 ( .A(n28569), .B(n38435), .X(n28568) );
  nand_x1_sg U53317 ( .A(n26885), .B(n38437), .X(n26884) );
  nand_x1_sg U53318 ( .A(n26835), .B(n38453), .X(n26834) );
  nand_x1_sg U53319 ( .A(n28555), .B(n38454), .X(n28554) );
  nand_x1_sg U53320 ( .A(n26899), .B(n38455), .X(n26898) );
  nand_x1_sg U53321 ( .A(n26892), .B(n38456), .X(n26891) );
  nand_x1_sg U53322 ( .A(n20990), .B(n38434), .X(n20989) );
  nand_x1_sg U53323 ( .A(n28548), .B(n38436), .X(n28547) );
  inv_x1_sg U53324 ( .A(n26821), .X(n45790) );
  inv_x1_sg U53325 ( .A(n27986), .X(n45082) );
  inv_x1_sg U53326 ( .A(n27979), .X(n45038) );
  inv_x1_sg U53327 ( .A(n28996), .X(n45069) );
  inv_x1_sg U53328 ( .A(n29009), .X(n45161) );
  inv_x1_sg U53329 ( .A(n29022), .X(n45252) );
  inv_x1_sg U53330 ( .A(n29035), .X(n45342) );
  inv_x1_sg U53331 ( .A(n29048), .X(n45433) );
  inv_x1_sg U53332 ( .A(n29061), .X(n45522) );
  inv_x1_sg U53333 ( .A(n29074), .X(n45611) );
  nand_x1_sg U53334 ( .A(n20834), .B(n38202), .X(n20833) );
  nand_x1_sg U53335 ( .A(n20191), .B(n38203), .X(n20190) );
  nand_x1_sg U53336 ( .A(n19385), .B(n38204), .X(n19384) );
  nand_x1_sg U53337 ( .A(n19162), .B(n38198), .X(n19161) );
  nand_x1_sg U53338 ( .A(n20798), .B(n38216), .X(n20797) );
  nand_x1_sg U53339 ( .A(n20801), .B(n38215), .X(n20800) );
  nand_x1_sg U53340 ( .A(n20804), .B(n38205), .X(n20803) );
  nand_x1_sg U53341 ( .A(n20807), .B(n38206), .X(n20806) );
  nand_x1_sg U53342 ( .A(n20810), .B(n38207), .X(n20809) );
  nand_x1_sg U53343 ( .A(n20813), .B(n38208), .X(n20812) );
  nand_x1_sg U53344 ( .A(n20816), .B(n38209), .X(n20815) );
  nand_x1_sg U53345 ( .A(n20819), .B(n38210), .X(n20818) );
  nand_x1_sg U53346 ( .A(n20822), .B(n38211), .X(n20821) );
  nand_x1_sg U53347 ( .A(n20825), .B(n38212), .X(n20824) );
  nand_x1_sg U53348 ( .A(n20828), .B(n38213), .X(n20827) );
  nand_x1_sg U53349 ( .A(n20831), .B(n38214), .X(n20830) );
  nand_x1_sg U53350 ( .A(n20188), .B(n38226), .X(n20187) );
  nand_x1_sg U53351 ( .A(n20185), .B(n38225), .X(n20184) );
  nand_x1_sg U53352 ( .A(n20182), .B(n38224), .X(n20181) );
  nand_x1_sg U53353 ( .A(n20179), .B(n38223), .X(n20178) );
  nand_x1_sg U53354 ( .A(n19382), .B(n38235), .X(n19381) );
  nand_x1_sg U53355 ( .A(n20176), .B(n38222), .X(n20175) );
  nand_x1_sg U53356 ( .A(n19379), .B(n38234), .X(n19378) );
  nand_x1_sg U53357 ( .A(n20173), .B(n38221), .X(n20172) );
  nand_x1_sg U53358 ( .A(n19376), .B(n38233), .X(n19375) );
  nand_x1_sg U53359 ( .A(n20170), .B(n38220), .X(n20169) );
  nand_x1_sg U53360 ( .A(n19373), .B(n38232), .X(n19372) );
  nand_x1_sg U53361 ( .A(n20167), .B(n38219), .X(n20166) );
  nand_x1_sg U53362 ( .A(n19370), .B(n38231), .X(n19369) );
  nand_x1_sg U53363 ( .A(n19367), .B(n38230), .X(n19366) );
  nand_x1_sg U53364 ( .A(n19364), .B(n38229), .X(n19363) );
  nand_x1_sg U53365 ( .A(n19361), .B(n38228), .X(n19360) );
  nand_x1_sg U53366 ( .A(n21022), .B(n38250), .X(n21021) );
  nand_x1_sg U53367 ( .A(n21025), .B(n38249), .X(n21024) );
  nand_x1_sg U53368 ( .A(n21028), .B(n38240), .X(n21027) );
  nand_x1_sg U53369 ( .A(n21031), .B(n38241), .X(n21030) );
  nand_x1_sg U53370 ( .A(n21034), .B(n38242), .X(n21033) );
  nand_x1_sg U53371 ( .A(n21037), .B(n38243), .X(n21036) );
  nand_x1_sg U53372 ( .A(n21040), .B(n38244), .X(n21039) );
  nand_x1_sg U53373 ( .A(n21043), .B(n38245), .X(n21042) );
  nand_x1_sg U53374 ( .A(n21046), .B(n38246), .X(n21045) );
  nand_x1_sg U53375 ( .A(n21049), .B(n38247), .X(n21048) );
  nand_x1_sg U53376 ( .A(n21052), .B(n38248), .X(n21051) );
  nand_x1_sg U53377 ( .A(n21055), .B(n38236), .X(n21054) );
  nand_x1_sg U53378 ( .A(n19592), .B(n38261), .X(n19591) );
  nand_x1_sg U53379 ( .A(n28090), .B(n38350), .X(n28089) );
  nand_x1_sg U53380 ( .A(n28087), .B(n38359), .X(n28086) );
  nand_x1_sg U53381 ( .A(n27925), .B(n38368), .X(n27924) );
  nand_x1_sg U53382 ( .A(n27748), .B(n38377), .X(n27747) );
  nand_x1_sg U53383 ( .A(n27554), .B(n38386), .X(n27553) );
  nand_x1_sg U53384 ( .A(n27341), .B(n38395), .X(n27340) );
  nand_x1_sg U53385 ( .A(n27111), .B(n38404), .X(n27110) );
  nand_x1_sg U53386 ( .A(n20343), .B(n38259), .X(n20342) );
  nand_x1_sg U53387 ( .A(n20337), .B(n38257), .X(n20336) );
  nand_x1_sg U53388 ( .A(n20334), .B(n38256), .X(n20333) );
  nand_x1_sg U53389 ( .A(n19613), .B(n38238), .X(n19612) );
  nand_x1_sg U53390 ( .A(n20331), .B(n38255), .X(n20330) );
  nand_x1_sg U53391 ( .A(n19610), .B(n38267), .X(n19609) );
  nand_x1_sg U53392 ( .A(n20328), .B(n38254), .X(n20327) );
  nand_x1_sg U53393 ( .A(n19607), .B(n38266), .X(n19606) );
  nand_x1_sg U53394 ( .A(n20325), .B(n38253), .X(n20324) );
  nand_x1_sg U53395 ( .A(n19604), .B(n38265), .X(n19603) );
  nand_x1_sg U53396 ( .A(n19601), .B(n38264), .X(n19600) );
  nand_x1_sg U53397 ( .A(n19598), .B(n38263), .X(n19597) );
  nand_x1_sg U53398 ( .A(n19595), .B(n38262), .X(n19594) );
  nand_x1_sg U53399 ( .A(n28972), .B(n38514), .X(n28971) );
  nand_x1_sg U53400 ( .A(n28966), .B(n38506), .X(n28965) );
  nand_x1_sg U53401 ( .A(n28960), .B(n38498), .X(n28959) );
  nand_x1_sg U53402 ( .A(n28954), .B(n38490), .X(n28953) );
  nand_x1_sg U53403 ( .A(n28948), .B(n38482), .X(n28947) );
  nand_x1_sg U53404 ( .A(n28942), .B(n38474), .X(n28941) );
  nand_x1_sg U53405 ( .A(n28936), .B(n38466), .X(n28935) );
  nand_x1_sg U53406 ( .A(n27964), .B(n38285), .X(n27963) );
  nand_x1_sg U53407 ( .A(n27961), .B(n38288), .X(n27960) );
  nand_x1_sg U53408 ( .A(n28111), .B(n38292), .X(n28110) );
  nand_x1_sg U53409 ( .A(n28108), .B(n38296), .X(n28107) );
  nand_x1_sg U53410 ( .A(n28105), .B(n38305), .X(n28104) );
  nand_x1_sg U53411 ( .A(n28102), .B(n38314), .X(n28101) );
  nand_x1_sg U53412 ( .A(n28099), .B(n38323), .X(n28098) );
  nand_x1_sg U53413 ( .A(n28096), .B(n38332), .X(n28095) );
  nand_x1_sg U53414 ( .A(n28093), .B(n38341), .X(n28092) );
  nand_x1_sg U53415 ( .A(n20346), .B(n38237), .X(n20345) );
  nand_x1_sg U53416 ( .A(n20340), .B(n38258), .X(n20339) );
  inv_x1_sg U53417 ( .A(n21668), .X(n46417) );
  nand_x1_sg U53418 ( .A(n21548), .B(n38442), .X(n21547) );
  nand_x1_sg U53419 ( .A(n21554), .B(n38444), .X(n21553) );
  nand_x1_sg U53420 ( .A(n21560), .B(n38446), .X(n21559) );
  nand_x1_sg U53421 ( .A(n21566), .B(n38448), .X(n21565) );
  nand_x1_sg U53422 ( .A(n21572), .B(n38450), .X(n21571) );
  nand_x1_sg U53423 ( .A(n21578), .B(n38452), .X(n21577) );
  nand_x1_sg U53424 ( .A(n21584), .B(n38428), .X(n21583) );
  nand_x1_sg U53425 ( .A(n21193), .B(n38421), .X(n21192) );
  nand_x1_sg U53426 ( .A(n28457), .B(n38517), .X(n28456) );
  nand_x1_sg U53427 ( .A(n21363), .B(n38413), .X(n21362) );
  nand_x1_sg U53428 ( .A(n28454), .B(n38513), .X(n28453) );
  nand_x1_sg U53429 ( .A(n28451), .B(n38509), .X(n28450) );
  nand_x1_sg U53430 ( .A(n28448), .B(n38505), .X(n28447) );
  nand_x1_sg U53431 ( .A(n28445), .B(n38501), .X(n28444) );
  nand_x1_sg U53432 ( .A(n28442), .B(n38497), .X(n28441) );
  nand_x1_sg U53433 ( .A(n28439), .B(n38493), .X(n28438) );
  nand_x1_sg U53434 ( .A(n28436), .B(n38489), .X(n28435) );
  nand_x1_sg U53435 ( .A(n28338), .B(n38324), .X(n28337) );
  nand_x1_sg U53436 ( .A(n28209), .B(n38333), .X(n28208) );
  nand_x1_sg U53437 ( .A(n28074), .B(n38342), .X(n28073) );
  nand_x1_sg U53438 ( .A(n27912), .B(n38351), .X(n27911) );
  nand_x1_sg U53439 ( .A(n27735), .B(n38360), .X(n27734) );
  nand_x1_sg U53440 ( .A(n27541), .B(n38369), .X(n27540) );
  nand_x1_sg U53441 ( .A(n27328), .B(n38378), .X(n27327) );
  nand_x1_sg U53442 ( .A(n27098), .B(n38387), .X(n27097) );
  nand_x1_sg U53443 ( .A(n27186), .B(n38519), .X(n27185) );
  nand_x1_sg U53444 ( .A(n27183), .B(n38516), .X(n27182) );
  nand_x1_sg U53445 ( .A(n27180), .B(n38512), .X(n27179) );
  nand_x1_sg U53446 ( .A(n27177), .B(n38508), .X(n27176) );
  nand_x1_sg U53447 ( .A(n27174), .B(n38504), .X(n27173) );
  nand_x1_sg U53448 ( .A(n27171), .B(n38500), .X(n27170) );
  nand_x1_sg U53449 ( .A(n27168), .B(n38496), .X(n27167) );
  nand_x1_sg U53450 ( .A(n27165), .B(n38492), .X(n27164) );
  nand_x1_sg U53451 ( .A(n27162), .B(n38488), .X(n27161) );
  nand_x1_sg U53452 ( .A(n27159), .B(n38484), .X(n27158) );
  nand_x1_sg U53453 ( .A(n27156), .B(n38480), .X(n27155) );
  nand_x1_sg U53454 ( .A(n27153), .B(n38476), .X(n27152) );
  nand_x1_sg U53455 ( .A(n27150), .B(n38472), .X(n27149) );
  nand_x1_sg U53456 ( .A(n27147), .B(n38468), .X(n27146) );
  nand_x1_sg U53457 ( .A(n27144), .B(n38464), .X(n27143) );
  nand_x1_sg U53458 ( .A(n27141), .B(n38460), .X(n27140) );
  inv_x1_sg U53459 ( .A(n21533), .X(n46502) );
  nand_x1_sg U53460 ( .A(n28975), .B(n38518), .X(n28974) );
  nand_x1_sg U53461 ( .A(n28969), .B(n38510), .X(n28968) );
  nand_x1_sg U53462 ( .A(n28963), .B(n38502), .X(n28962) );
  nand_x1_sg U53463 ( .A(n28957), .B(n38494), .X(n28956) );
  nand_x1_sg U53464 ( .A(n28332), .B(n38485), .X(n28331) );
  nand_x1_sg U53465 ( .A(n28951), .B(n38486), .X(n28950) );
  nand_x1_sg U53466 ( .A(n28203), .B(n38481), .X(n28202) );
  nand_x1_sg U53467 ( .A(n28068), .B(n38477), .X(n28067) );
  nand_x1_sg U53468 ( .A(n28945), .B(n38478), .X(n28944) );
  nand_x1_sg U53469 ( .A(n27906), .B(n38473), .X(n27905) );
  nand_x1_sg U53470 ( .A(n27729), .B(n38469), .X(n27728) );
  nand_x1_sg U53471 ( .A(n28939), .B(n38470), .X(n28938) );
  nand_x1_sg U53472 ( .A(n27535), .B(n38465), .X(n27534) );
  nand_x1_sg U53473 ( .A(n27322), .B(n38461), .X(n27321) );
  nand_x1_sg U53474 ( .A(n28933), .B(n38462), .X(n28932) );
  nand_x1_sg U53475 ( .A(n27092), .B(n38457), .X(n27091) );
  nand_x1_sg U53476 ( .A(n28754), .B(n38458), .X(n28753) );
  nand_x1_sg U53477 ( .A(n28617), .B(n38298), .X(n28616) );
  nand_x1_sg U53478 ( .A(n28614), .B(n38307), .X(n28613) );
  nand_x1_sg U53479 ( .A(n28611), .B(n38316), .X(n28610) );
  nand_x1_sg U53480 ( .A(n28608), .B(n38325), .X(n28607) );
  nand_x1_sg U53481 ( .A(n28605), .B(n38334), .X(n28604) );
  nand_x1_sg U53482 ( .A(n28602), .B(n38343), .X(n28601) );
  nand_x1_sg U53483 ( .A(n28599), .B(n38352), .X(n28598) );
  nand_x1_sg U53484 ( .A(n28362), .B(n38281), .X(n28361) );
  nand_x1_sg U53485 ( .A(n27793), .B(n38294), .X(n27792) );
  nand_x1_sg U53486 ( .A(n28802), .B(n38299), .X(n28801) );
  nand_x1_sg U53487 ( .A(n27790), .B(n38303), .X(n27789) );
  nand_x1_sg U53488 ( .A(n27787), .B(n38312), .X(n27786) );
  nand_x1_sg U53489 ( .A(n28796), .B(n38317), .X(n28795) );
  nand_x1_sg U53490 ( .A(n27784), .B(n38321), .X(n27783) );
  nand_x1_sg U53491 ( .A(n27781), .B(n38330), .X(n27780) );
  nand_x1_sg U53492 ( .A(n28790), .B(n38335), .X(n28789) );
  nand_x1_sg U53493 ( .A(n27778), .B(n38339), .X(n27777) );
  nand_x1_sg U53494 ( .A(n27775), .B(n38348), .X(n27774) );
  nand_x1_sg U53495 ( .A(n28784), .B(n38353), .X(n28783) );
  nand_x1_sg U53496 ( .A(n27772), .B(n38357), .X(n27771) );
  nand_x1_sg U53497 ( .A(n27769), .B(n38366), .X(n27768) );
  nand_x1_sg U53498 ( .A(n28778), .B(n38371), .X(n28777) );
  nand_x1_sg U53499 ( .A(n27766), .B(n38375), .X(n27765) );
  nand_x1_sg U53500 ( .A(n27763), .B(n38384), .X(n27762) );
  nand_x1_sg U53501 ( .A(n28772), .B(n38389), .X(n28771) );
  nand_x1_sg U53502 ( .A(n27760), .B(n38393), .X(n27759) );
  nand_x1_sg U53503 ( .A(n27566), .B(n38402), .X(n27565) );
  nand_x1_sg U53504 ( .A(n28766), .B(n38406), .X(n28765) );
  nand_x1_sg U53505 ( .A(n27353), .B(n38410), .X(n27352) );
  nand_x1_sg U53506 ( .A(n28763), .B(n38415), .X(n28762) );
  nand_x1_sg U53507 ( .A(n27123), .B(n38419), .X(n27122) );
  nand_x1_sg U53508 ( .A(n28760), .B(n38423), .X(n28759) );
  nand_x1_sg U53509 ( .A(n28596), .B(n38361), .X(n28595) );
  nand_x1_sg U53510 ( .A(n28593), .B(n38370), .X(n28592) );
  nand_x1_sg U53511 ( .A(n28590), .B(n38379), .X(n28589) );
  nand_x1_sg U53512 ( .A(n28587), .B(n38388), .X(n28586) );
  nand_x1_sg U53513 ( .A(n28584), .B(n38397), .X(n28583) );
  nand_x1_sg U53514 ( .A(n28581), .B(n38405), .X(n28580) );
  nand_x1_sg U53515 ( .A(n28578), .B(n38414), .X(n28577) );
  nand_x1_sg U53516 ( .A(n28575), .B(n38422), .X(n28574) );
  nand_x1_sg U53517 ( .A(n28927), .B(n38424), .X(n28926) );
  nand_x1_sg U53518 ( .A(n28572), .B(n38429), .X(n28571) );
  nand_x1_sg U53519 ( .A(n28748), .B(n38431), .X(n28747) );
  nand_x1_sg U53520 ( .A(n28359), .B(n38282), .X(n28358) );
  nand_x1_sg U53521 ( .A(n28356), .B(n38284), .X(n28355) );
  nand_x1_sg U53522 ( .A(n28353), .B(n38286), .X(n28352) );
  nand_x1_sg U53523 ( .A(n28350), .B(n38293), .X(n28349) );
  nand_x1_sg U53524 ( .A(n28347), .B(n38297), .X(n28346) );
  nand_x1_sg U53525 ( .A(n28344), .B(n38306), .X(n28343) );
  nand_x1_sg U53526 ( .A(n28341), .B(n38315), .X(n28340) );
  inv_x1_sg U53527 ( .A(n29195), .X(n45386) );
  inv_x1_sg U53528 ( .A(n29207), .X(n45476) );
  inv_x1_sg U53529 ( .A(n29219), .X(n45565) );
  inv_x1_sg U53530 ( .A(n29084), .X(n45653) );
  nand_x1_sg U53531 ( .A(n27796), .B(n38287), .X(n27795) );
  nand_x1_sg U53532 ( .A(n28805), .B(n38289), .X(n28804) );
  nand_x1_sg U53533 ( .A(n27958), .B(n38295), .X(n27957) );
  nand_x1_sg U53534 ( .A(n27407), .B(n38301), .X(n27406) );
  nand_x1_sg U53535 ( .A(n27955), .B(n38304), .X(n27954) );
  nand_x1_sg U53536 ( .A(n28799), .B(n38308), .X(n28798) );
  nand_x1_sg U53537 ( .A(n27404), .B(n38310), .X(n27403) );
  nand_x1_sg U53538 ( .A(n27952), .B(n38313), .X(n27951) );
  nand_x1_sg U53539 ( .A(n27401), .B(n38319), .X(n27400) );
  nand_x1_sg U53540 ( .A(n27949), .B(n38322), .X(n27948) );
  nand_x1_sg U53541 ( .A(n28793), .B(n38326), .X(n28792) );
  nand_x1_sg U53542 ( .A(n27398), .B(n38328), .X(n27397) );
  nand_x1_sg U53543 ( .A(n27946), .B(n38331), .X(n27945) );
  nand_x1_sg U53544 ( .A(n27395), .B(n38337), .X(n27394) );
  nand_x1_sg U53545 ( .A(n27943), .B(n38340), .X(n27942) );
  nand_x1_sg U53546 ( .A(n28787), .B(n38344), .X(n28786) );
  nand_x1_sg U53547 ( .A(n27392), .B(n38346), .X(n27391) );
  nand_x1_sg U53548 ( .A(n27940), .B(n38349), .X(n27939) );
  nand_x1_sg U53549 ( .A(n27389), .B(n38355), .X(n27388) );
  nand_x1_sg U53550 ( .A(n27937), .B(n38358), .X(n27936) );
  nand_x1_sg U53551 ( .A(n28781), .B(n38362), .X(n28780) );
  nand_x1_sg U53552 ( .A(n27386), .B(n38364), .X(n27385) );
  nand_x1_sg U53553 ( .A(n27934), .B(n38367), .X(n27933) );
  nand_x1_sg U53554 ( .A(n27383), .B(n38373), .X(n27382) );
  nand_x1_sg U53555 ( .A(n27931), .B(n38376), .X(n27930) );
  nand_x1_sg U53556 ( .A(n28775), .B(n38380), .X(n28774) );
  nand_x1_sg U53557 ( .A(n27380), .B(n38382), .X(n27379) );
  nand_x1_sg U53558 ( .A(n27754), .B(n38385), .X(n27753) );
  nand_x1_sg U53559 ( .A(n27377), .B(n38391), .X(n27376) );
  nand_x1_sg U53560 ( .A(n27560), .B(n38394), .X(n27559) );
  nand_x1_sg U53561 ( .A(n28769), .B(n38398), .X(n28768) );
  nand_x1_sg U53562 ( .A(n27374), .B(n38400), .X(n27373) );
  nand_x1_sg U53563 ( .A(n27347), .B(n38403), .X(n27346) );
  nand_x1_sg U53564 ( .A(n27371), .B(n38408), .X(n27370) );
  nand_x1_sg U53565 ( .A(n27117), .B(n38411), .X(n27116) );
  nand_x1_sg U53566 ( .A(n27368), .B(n38417), .X(n27367) );
  nand_x1_sg U53567 ( .A(n27365), .B(n38425), .X(n27364) );
  nand_x1_sg U53568 ( .A(n27135), .B(n38432), .X(n27134) );
  nand_x1_sg U53569 ( .A(n27611), .B(n38290), .X(n27610) );
  nand_x1_sg U53570 ( .A(n27608), .B(n38302), .X(n27607) );
  nand_x1_sg U53571 ( .A(n27605), .B(n38311), .X(n27604) );
  nand_x1_sg U53572 ( .A(n27602), .B(n38320), .X(n27601) );
  nand_x1_sg U53573 ( .A(n27599), .B(n38329), .X(n27598) );
  nand_x1_sg U53574 ( .A(n27596), .B(n38338), .X(n27595) );
  nand_x1_sg U53575 ( .A(n27593), .B(n38347), .X(n27592) );
  nand_x1_sg U53576 ( .A(n27590), .B(n38356), .X(n27589) );
  nand_x1_sg U53577 ( .A(n27587), .B(n38365), .X(n27586) );
  nand_x1_sg U53578 ( .A(n27584), .B(n38374), .X(n27583) );
  nand_x1_sg U53579 ( .A(n27581), .B(n38383), .X(n27580) );
  nand_x1_sg U53580 ( .A(n27578), .B(n38392), .X(n27577) );
  nand_x1_sg U53581 ( .A(n27575), .B(n38401), .X(n27574) );
  nand_x1_sg U53582 ( .A(n27572), .B(n38409), .X(n27571) );
  nand_x1_sg U53583 ( .A(n27359), .B(n38418), .X(n27358) );
  nand_x1_sg U53584 ( .A(n27129), .B(n38426), .X(n27128) );
  nand_x1_sg U53585 ( .A(n29135), .B(n38300), .X(n29134) );
  nand_x1_sg U53586 ( .A(n26947), .B(n38280), .X(n26946) );
  nand_x1_sg U53587 ( .A(n29129), .B(n38318), .X(n29128) );
  nand_x1_sg U53588 ( .A(n26944), .B(n38515), .X(n26943) );
  nand_x1_sg U53589 ( .A(n26941), .B(n38511), .X(n26940) );
  nand_x1_sg U53590 ( .A(n29123), .B(n38336), .X(n29122) );
  nand_x1_sg U53591 ( .A(n26938), .B(n38507), .X(n26937) );
  nand_x1_sg U53592 ( .A(n26935), .B(n38503), .X(n26934) );
  nand_x1_sg U53593 ( .A(n29117), .B(n38354), .X(n29116) );
  nand_x1_sg U53594 ( .A(n26932), .B(n38499), .X(n26931) );
  nand_x1_sg U53595 ( .A(n26929), .B(n38495), .X(n26928) );
  nand_x1_sg U53596 ( .A(n29111), .B(n38372), .X(n29110) );
  nand_x1_sg U53597 ( .A(n26926), .B(n38491), .X(n26925) );
  nand_x1_sg U53598 ( .A(n26923), .B(n38487), .X(n26922) );
  nand_x1_sg U53599 ( .A(n29105), .B(n38390), .X(n29104) );
  nand_x1_sg U53600 ( .A(n26920), .B(n38483), .X(n26919) );
  nand_x1_sg U53601 ( .A(n26917), .B(n38479), .X(n26916) );
  nand_x1_sg U53602 ( .A(n29099), .B(n38407), .X(n29098) );
  nand_x1_sg U53603 ( .A(n26914), .B(n38475), .X(n26913) );
  nand_x1_sg U53604 ( .A(n26911), .B(n38471), .X(n26910) );
  nand_x1_sg U53605 ( .A(n26908), .B(n38467), .X(n26907) );
  nand_x1_sg U53606 ( .A(n26905), .B(n38463), .X(n26904) );
  nand_x1_sg U53607 ( .A(n26902), .B(n38459), .X(n26901) );
  inv_x1_sg U53608 ( .A(n21656), .X(n46328) );
  inv_x1_sg U53609 ( .A(n21644), .X(n46237) );
  inv_x1_sg U53610 ( .A(n21632), .X(n46146) );
  inv_x1_sg U53611 ( .A(n21620), .X(n46055) );
  inv_x1_sg U53612 ( .A(n21608), .X(n45964) );
  inv_x1_sg U53613 ( .A(n28382), .X(n45077) );
  inv_x1_sg U53614 ( .A(n28424), .X(n45396) );
  inv_x1_sg U53615 ( .A(n28418), .X(n45350) );
  inv_x1_sg U53616 ( .A(n28412), .X(n45305) );
  inv_x1_sg U53617 ( .A(n28406), .X(n45260) );
  inv_x1_sg U53618 ( .A(n28400), .X(n45215) );
  inv_x1_sg U53619 ( .A(n28394), .X(n45169) );
  inv_x1_sg U53620 ( .A(n28388), .X(n45124) );
  inv_x1_sg U53621 ( .A(n27077), .X(n45752) );
  inv_x1_sg U53622 ( .A(n27056), .X(n45766) );
  inv_x1_sg U53623 ( .A(n27050), .X(n45723) );
  inv_x1_sg U53624 ( .A(n27044), .X(n45680) );
  inv_x1_sg U53625 ( .A(n27038), .X(n45636) );
  inv_x1_sg U53626 ( .A(n27032), .X(n45592) );
  inv_x1_sg U53627 ( .A(n27026), .X(n45547) );
  inv_x1_sg U53628 ( .A(n27020), .X(n45503) );
  inv_x1_sg U53629 ( .A(n27014), .X(n45455) );
  inv_x1_sg U53630 ( .A(n27008), .X(n45411) );
  inv_x1_sg U53631 ( .A(n27002), .X(n45365) );
  inv_x1_sg U53632 ( .A(n26996), .X(n45320) );
  inv_x1_sg U53633 ( .A(n26990), .X(n45275) );
  inv_x1_sg U53634 ( .A(n26984), .X(n45230) );
  inv_x1_sg U53635 ( .A(n26978), .X(n45184) );
  inv_x1_sg U53636 ( .A(n26972), .X(n45139) );
  inv_x1_sg U53637 ( .A(n26966), .X(n45092) );
  inv_x1_sg U53638 ( .A(n26960), .X(n45048) );
  inv_x1_sg U53639 ( .A(n21351), .X(n46544) );
  inv_x1_sg U53640 ( .A(n27080), .X(n45750) );
  inv_x1_sg U53641 ( .A(n28730), .X(n45744) );
  inv_x1_sg U53642 ( .A(n27310), .X(n45707) );
  inv_x1_sg U53643 ( .A(n28909), .X(n45701) );
  inv_x1_sg U53644 ( .A(n27523), .X(n45663) );
  inv_x1_sg U53645 ( .A(n28903), .X(n45657) );
  inv_x1_sg U53646 ( .A(n27717), .X(n45619) );
  inv_x1_sg U53647 ( .A(n28897), .X(n45613) );
  inv_x1_sg U53648 ( .A(n27894), .X(n45575) );
  inv_x1_sg U53649 ( .A(n28891), .X(n45569) );
  inv_x1_sg U53650 ( .A(n28056), .X(n45530) );
  inv_x1_sg U53651 ( .A(n28885), .X(n45524) );
  inv_x1_sg U53652 ( .A(n28191), .X(n45486) );
  inv_x1_sg U53653 ( .A(n28879), .X(n45480) );
  inv_x1_sg U53654 ( .A(n28320), .X(n45441) );
  inv_x1_sg U53655 ( .A(n28873), .X(n45435) );
  inv_x1_sg U53656 ( .A(n28867), .X(n45390) );
  inv_x1_sg U53657 ( .A(n28861), .X(n45344) );
  inv_x1_sg U53658 ( .A(n28855), .X(n45299) );
  inv_x1_sg U53659 ( .A(n28849), .X(n45254) );
  inv_x1_sg U53660 ( .A(n28843), .X(n45209) );
  inv_x1_sg U53661 ( .A(n28837), .X(n45163) );
  inv_x1_sg U53662 ( .A(n28831), .X(n45118) );
  inv_x1_sg U53663 ( .A(n28825), .X(n45071) );
  inv_x1_sg U53664 ( .A(n28376), .X(n45034) );
  inv_x1_sg U53665 ( .A(n28819), .X(n45028) );
  inv_x1_sg U53666 ( .A(n28470), .X(n45032) );
  inv_x1_sg U53667 ( .A(n28476), .X(n45075) );
  inv_x1_sg U53668 ( .A(n28482), .X(n45122) );
  inv_x1_sg U53669 ( .A(n28488), .X(n45167) );
  inv_x1_sg U53670 ( .A(n28494), .X(n45213) );
  inv_x1_sg U53671 ( .A(n28500), .X(n45258) );
  inv_x1_sg U53672 ( .A(n28506), .X(n45303) );
  inv_x1_sg U53673 ( .A(n28512), .X(n45348) );
  inv_x1_sg U53674 ( .A(n28631), .X(n45030) );
  inv_x1_sg U53675 ( .A(n27636), .X(n45133) );
  inv_x1_sg U53676 ( .A(n28643), .X(n45120) );
  inv_x1_sg U53677 ( .A(n29159), .X(n45114) );
  inv_x1_sg U53678 ( .A(n27642), .X(n45178) );
  inv_x1_sg U53679 ( .A(n27648), .X(n45224) );
  inv_x1_sg U53680 ( .A(n28655), .X(n45211) );
  inv_x1_sg U53681 ( .A(n29171), .X(n45205) );
  inv_x1_sg U53682 ( .A(n27654), .X(n45269) );
  inv_x1_sg U53683 ( .A(n27660), .X(n45314) );
  inv_x1_sg U53684 ( .A(n28667), .X(n45301) );
  inv_x1_sg U53685 ( .A(n29183), .X(n45295) );
  inv_x1_sg U53686 ( .A(n27666), .X(n45359) );
  inv_x1_sg U53687 ( .A(n27672), .X(n45405) );
  inv_x1_sg U53688 ( .A(n28679), .X(n45392) );
  inv_x1_sg U53689 ( .A(n27678), .X(n45449) );
  inv_x1_sg U53690 ( .A(n27684), .X(n45497) );
  inv_x1_sg U53691 ( .A(n28691), .X(n45482) );
  inv_x1_sg U53692 ( .A(n27690), .X(n45541) );
  inv_x1_sg U53693 ( .A(n27696), .X(n45586) );
  inv_x1_sg U53694 ( .A(n28703), .X(n45571) );
  inv_x1_sg U53695 ( .A(n27702), .X(n45630) );
  inv_x1_sg U53696 ( .A(n27508), .X(n45674) );
  inv_x1_sg U53697 ( .A(n28715), .X(n45659) );
  inv_x1_sg U53698 ( .A(n27295), .X(n45717) );
  inv_x1_sg U53699 ( .A(n28721), .X(n45703) );
  inv_x1_sg U53700 ( .A(n28915), .X(n45697) );
  inv_x1_sg U53701 ( .A(n27065), .X(n45760) );
  inv_x1_sg U53702 ( .A(n28727), .X(n45746) );
  inv_x1_sg U53703 ( .A(n28990), .X(n45026) );
  inv_x1_sg U53704 ( .A(n29003), .X(n45116) );
  inv_x1_sg U53705 ( .A(n29016), .X(n45207) );
  inv_x1_sg U53706 ( .A(n29029), .X(n45297) );
  inv_x1_sg U53707 ( .A(n28427), .X(n45394) );
  inv_x1_sg U53708 ( .A(n29042), .X(n45388) );
  inv_x1_sg U53709 ( .A(n28323), .X(n45439) );
  inv_x1_sg U53710 ( .A(n28194), .X(n45484) );
  inv_x1_sg U53711 ( .A(n29055), .X(n45478) );
  inv_x1_sg U53712 ( .A(n28059), .X(n45528) );
  inv_x1_sg U53713 ( .A(n27897), .X(n45573) );
  inv_x1_sg U53714 ( .A(n29068), .X(n45567) );
  inv_x1_sg U53715 ( .A(n27720), .X(n45617) );
  inv_x1_sg U53716 ( .A(n27526), .X(n45661) );
  inv_x1_sg U53717 ( .A(n29081), .X(n45655) );
  inv_x1_sg U53718 ( .A(n27313), .X(n45705) );
  inv_x1_sg U53719 ( .A(n28912), .X(n45699) );
  inv_x1_sg U53720 ( .A(n27083), .X(n45748) );
  inv_x1_sg U53721 ( .A(n28733), .X(n45742) );
  inv_x1_sg U53722 ( .A(n27810), .X(n45040) );
  inv_x1_sg U53723 ( .A(n27624), .X(n45042) );
  inv_x1_sg U53724 ( .A(n27816), .X(n45084) );
  inv_x1_sg U53725 ( .A(n27630), .X(n45086) );
  inv_x1_sg U53726 ( .A(n27822), .X(n45131) );
  inv_x1_sg U53727 ( .A(n28637), .X(n45073) );
  inv_x1_sg U53728 ( .A(n27199), .X(n45046) );
  inv_x1_sg U53729 ( .A(n27828), .X(n45176) );
  inv_x1_sg U53730 ( .A(n27205), .X(n45090) );
  inv_x1_sg U53731 ( .A(n27834), .X(n45222) );
  inv_x1_sg U53732 ( .A(n28649), .X(n45165) );
  inv_x1_sg U53733 ( .A(n27211), .X(n45137) );
  inv_x1_sg U53734 ( .A(n27840), .X(n45267) );
  inv_x1_sg U53735 ( .A(n27217), .X(n45182) );
  inv_x1_sg U53736 ( .A(n27846), .X(n45312) );
  inv_x1_sg U53737 ( .A(n28661), .X(n45256) );
  inv_x1_sg U53738 ( .A(n27223), .X(n45228) );
  inv_x1_sg U53739 ( .A(n27852), .X(n45357) );
  inv_x1_sg U53740 ( .A(n27229), .X(n45273) );
  inv_x1_sg U53741 ( .A(n27858), .X(n45403) );
  inv_x1_sg U53742 ( .A(n28673), .X(n45346) );
  inv_x1_sg U53743 ( .A(n27235), .X(n45318) );
  inv_x1_sg U53744 ( .A(n27864), .X(n45447) );
  inv_x1_sg U53745 ( .A(n27241), .X(n45363) );
  inv_x1_sg U53746 ( .A(n27870), .X(n45495) );
  inv_x1_sg U53747 ( .A(n28685), .X(n45437) );
  inv_x1_sg U53748 ( .A(n27247), .X(n45409) );
  inv_x1_sg U53749 ( .A(n27876), .X(n45539) );
  inv_x1_sg U53750 ( .A(n27253), .X(n45453) );
  inv_x1_sg U53751 ( .A(n27882), .X(n45584) );
  inv_x1_sg U53752 ( .A(n28697), .X(n45526) );
  inv_x1_sg U53753 ( .A(n27259), .X(n45501) );
  inv_x1_sg U53754 ( .A(n27705), .X(n45628) );
  inv_x1_sg U53755 ( .A(n27265), .X(n45545) );
  inv_x1_sg U53756 ( .A(n27511), .X(n45672) );
  inv_x1_sg U53757 ( .A(n28709), .X(n45615) );
  inv_x1_sg U53758 ( .A(n27271), .X(n45590) );
  inv_x1_sg U53759 ( .A(n27298), .X(n45715) );
  inv_x1_sg U53760 ( .A(n27277), .X(n45634) );
  inv_x1_sg U53761 ( .A(n27068), .X(n45758) );
  inv_x1_sg U53762 ( .A(n27283), .X(n45678) );
  inv_x1_sg U53763 ( .A(n27289), .X(n45721) );
  inv_x1_sg U53764 ( .A(n27059), .X(n45764) );
  inv_x1_sg U53765 ( .A(n27993), .X(n45129) );
  inv_x1_sg U53766 ( .A(n27421), .X(n45044) );
  inv_x1_sg U53767 ( .A(n27999), .X(n45174) );
  inv_x1_sg U53768 ( .A(n27427), .X(n45088) );
  inv_x1_sg U53769 ( .A(n28005), .X(n45220) );
  inv_x1_sg U53770 ( .A(n27433), .X(n45135) );
  inv_x1_sg U53771 ( .A(n28011), .X(n45265) );
  inv_x1_sg U53772 ( .A(n27439), .X(n45180) );
  inv_x1_sg U53773 ( .A(n28017), .X(n45310) );
  inv_x1_sg U53774 ( .A(n27445), .X(n45226) );
  inv_x1_sg U53775 ( .A(n28023), .X(n45355) );
  inv_x1_sg U53776 ( .A(n27451), .X(n45271) );
  inv_x1_sg U53777 ( .A(n28029), .X(n45401) );
  inv_x1_sg U53778 ( .A(n27457), .X(n45316) );
  inv_x1_sg U53779 ( .A(n28035), .X(n45445) );
  inv_x1_sg U53780 ( .A(n27463), .X(n45361) );
  inv_x1_sg U53781 ( .A(n28041), .X(n45493) );
  inv_x1_sg U53782 ( .A(n27469), .X(n45407) );
  inv_x1_sg U53783 ( .A(n28047), .X(n45537) );
  inv_x1_sg U53784 ( .A(n27475), .X(n45451) );
  inv_x1_sg U53785 ( .A(n27885), .X(n45582) );
  inv_x1_sg U53786 ( .A(n27481), .X(n45499) );
  inv_x1_sg U53787 ( .A(n27708), .X(n45626) );
  inv_x1_sg U53788 ( .A(n27487), .X(n45543) );
  inv_x1_sg U53789 ( .A(n27514), .X(n45670) );
  inv_x1_sg U53790 ( .A(n27493), .X(n45588) );
  inv_x1_sg U53791 ( .A(n27301), .X(n45713) );
  inv_x1_sg U53792 ( .A(n27499), .X(n45632) );
  inv_x1_sg U53793 ( .A(n27071), .X(n45756) );
  inv_x1_sg U53794 ( .A(n27505), .X(n45676) );
  inv_x1_sg U53795 ( .A(n27292), .X(n45719) );
  inv_x1_sg U53796 ( .A(n27062), .X(n45762) );
  nand_x1_sg U53797 ( .A(n21545), .B(n38441), .X(n21544) );
  nand_x1_sg U53798 ( .A(n21551), .B(n38443), .X(n21550) );
  nand_x1_sg U53799 ( .A(n21557), .B(n38445), .X(n21556) );
  nand_x1_sg U53800 ( .A(n21563), .B(n38447), .X(n21562) );
  nand_x1_sg U53801 ( .A(n21569), .B(n38449), .X(n21568) );
  nand_x1_sg U53802 ( .A(n21575), .B(n38451), .X(n21574) );
  nand_x1_sg U53803 ( .A(n21581), .B(n38439), .X(n21580) );
  nand_x1_sg U53804 ( .A(n29132), .B(n38309), .X(n29131) );
  nand_x1_sg U53805 ( .A(n29126), .B(n38327), .X(n29125) );
  nand_x1_sg U53806 ( .A(n29120), .B(n38345), .X(n29119) );
  nand_x1_sg U53807 ( .A(n29114), .B(n38363), .X(n29113) );
  nand_x1_sg U53808 ( .A(n29108), .B(n38381), .X(n29107) );
  nand_x1_sg U53809 ( .A(n29102), .B(n38399), .X(n29101) );
  nand_x1_sg U53810 ( .A(n29096), .B(n38416), .X(n29095) );
  nand_x1_sg U53811 ( .A(n28114), .B(n38291), .X(n28113) );
  nand_x1_sg U53812 ( .A(n28117), .B(n38283), .X(n28116) );
  inv_x1_sg U53813 ( .A(n21596), .X(n45872) );
  inv_x1_sg U53814 ( .A(n29147), .X(n45024) );
  inv_x1_sg U53815 ( .A(n19324), .X(n46569) );
  inv_x1_sg U53816 ( .A(n28534), .X(n45783) );
  inv_x1_sg U53817 ( .A(n20976), .X(n46618) );
  inv_x1_sg U53818 ( .A(n20119), .X(n46477) );
  inv_x1_sg U53819 ( .A(n21078), .X(n45876) );
  inv_x1_sg U53820 ( .A(n20369), .X(n45879) );
  inv_x1_sg U53821 ( .A(n19636), .X(n45882) );
  inv_x1_sg U53822 ( .A(n21172), .X(n46590) );
  inv_x1_sg U53823 ( .A(n20149), .X(n46473) );
  inv_x1_sg U53824 ( .A(n19957), .X(n46515) );
  nand_x1_sg U53825 ( .A(n19358), .B(n38227), .X(n19357) );
  nand_x1_sg U53826 ( .A(n21019), .B(n38251), .X(n21018) );
  nand_x1_sg U53827 ( .A(n20322), .B(n38252), .X(n20321) );
  inv_x1_sg U53828 ( .A(n21276), .X(n45915) );
  inv_x1_sg U53829 ( .A(n20507), .X(n45905) );
  inv_x1_sg U53830 ( .A(n19850), .X(n45895) );
  inv_x1_sg U53831 ( .A(n28141), .X(n45059) );
  inv_x1_sg U53832 ( .A(n6670), .X(n45885) );
  inv_x1_sg U53833 ( .A(n21163), .X(n46496) );
  inv_x1_sg U53834 ( .A(n21157), .X(n46458) );
  inv_x1_sg U53835 ( .A(n21151), .X(n46410) );
  inv_x1_sg U53836 ( .A(n21139), .X(n46321) );
  inv_x1_sg U53837 ( .A(n21145), .X(n46363) );
  inv_x1_sg U53838 ( .A(n21133), .X(n46276) );
  inv_x1_sg U53839 ( .A(n21127), .X(n46230) );
  inv_x1_sg U53840 ( .A(n21121), .X(n46185) );
  inv_x1_sg U53841 ( .A(n21115), .X(n46139) );
  inv_x1_sg U53842 ( .A(n21109), .X(n46094) );
  inv_x1_sg U53843 ( .A(n21103), .X(n46048) );
  inv_x1_sg U53844 ( .A(n21097), .X(n46003) );
  inv_x1_sg U53845 ( .A(n21091), .X(n45957) );
  inv_x1_sg U53846 ( .A(n20430), .X(n46312) );
  inv_x1_sg U53847 ( .A(n20382), .X(n45948) );
  inv_x1_sg U53848 ( .A(n20424), .X(n46267) );
  inv_x1_sg U53849 ( .A(n20418), .X(n46221) );
  inv_x1_sg U53850 ( .A(n20412), .X(n46176) );
  inv_x1_sg U53851 ( .A(n20406), .X(n46130) );
  inv_x1_sg U53852 ( .A(n20400), .X(n46085) );
  inv_x1_sg U53853 ( .A(n20394), .X(n46039) );
  inv_x1_sg U53854 ( .A(n20388), .X(n45994) );
  inv_x1_sg U53855 ( .A(n20312), .X(n46449) );
  inv_x1_sg U53856 ( .A(n19697), .X(n46303) );
  inv_x1_sg U53857 ( .A(n19691), .X(n46258) );
  inv_x1_sg U53858 ( .A(n19685), .X(n46212) );
  inv_x1_sg U53859 ( .A(n19679), .X(n46167) );
  inv_x1_sg U53860 ( .A(n19673), .X(n46121) );
  inv_x1_sg U53861 ( .A(n19667), .X(n46076) );
  inv_x1_sg U53862 ( .A(n19661), .X(n46030) );
  inv_x1_sg U53863 ( .A(n19655), .X(n45985) );
  inv_x1_sg U53864 ( .A(n19649), .X(n45939) );
  inv_x1_sg U53865 ( .A(n20151), .X(n46488) );
  inv_x1_sg U53866 ( .A(n19959), .X(n46532) );
  nand_x1_sg U53867 ( .A(n20997), .B(n38201), .X(n20996) );
  nand_x1_sg U53868 ( .A(n26849), .B(n38239), .X(n26848) );
  nand_x1_sg U53869 ( .A(n21012), .B(n38274), .X(n21011) );
  inv_x1_sg U53870 ( .A(n26816), .X(n45792) );
  inv_x1_sg U53871 ( .A(n26819), .X(n45791) );
  inv_x1_sg U53872 ( .A(n28523), .X(n45787) );
  inv_x1_sg U53873 ( .A(n28532), .X(n45784) );
  inv_x1_sg U53874 ( .A(n21182), .X(n46584) );
  inv_x1_sg U53875 ( .A(n28737), .X(n45740) );
  inv_x1_sg U53876 ( .A(n26955), .X(n45017) );
  inv_x1_sg U53877 ( .A(n28529), .X(n45785) );
  inv_x1_sg U53878 ( .A(n26813), .X(n45793) );
  inv_x1_sg U53879 ( .A(n26829), .X(n45788) );
  inv_x1_sg U53880 ( .A(n28526), .X(n45786) );
  inv_x1_sg U53881 ( .A(n26810), .X(n45794) );
  inv_x1_sg U53882 ( .A(n26807), .X(n45795) );
  inv_x1_sg U53883 ( .A(n26804), .X(n45796) );
  inv_x1_sg U53884 ( .A(n21006), .X(n46588) );
  nand_x1_sg U53885 ( .A(n21004), .B(n38270), .X(n21003) );
  inv_x1_sg U53886 ( .A(n19146), .X(n46606) );
  nand_x1_sg U53887 ( .A(n19144), .B(n38269), .X(n19143) );
  inv_x1_sg U53888 ( .A(n19570), .X(n46611) );
  nand_x1_sg U53889 ( .A(n19569), .B(n38271), .X(n19568) );
  inv_x1_sg U53890 ( .A(n20588), .X(n46592) );
  nand_x1_sg U53891 ( .A(n20587), .B(n38279), .X(n20586) );
  inv_x1_sg U53892 ( .A(n19796), .X(n46346) );
  nand_x1_sg U53893 ( .A(n41544), .B(n46558), .X(n19533) );
  nand_x1_sg U53894 ( .A(n19535), .B(n38276), .X(n19534) );
  nand_x1_sg U53895 ( .A(n41542), .B(n46562), .X(n19547) );
  nand_x1_sg U53896 ( .A(n19549), .B(n38272), .X(n19548) );
  nand_x1_sg U53897 ( .A(n41543), .B(n46565), .X(n19554) );
  nand_x1_sg U53898 ( .A(n19556), .B(n38273), .X(n19555) );
  nand_x1_sg U53899 ( .A(n41541), .B(n46576), .X(n19561) );
  nand_x1_sg U53900 ( .A(n19563), .B(n38277), .X(n19562) );
  nand_x1_sg U53901 ( .A(n41547), .B(n46572), .X(n19150) );
  nand_x1_sg U53902 ( .A(n19152), .B(n38278), .X(n19151) );
  nand_x1_sg U53903 ( .A(n41549), .B(n46560), .X(n19540) );
  nand_x1_sg U53904 ( .A(n19542), .B(n38275), .X(n19541) );
  nand_x1_sg U53905 ( .A(n22546), .B(n45019), .X(n22545) );
  inv_x1_sg U53906 ( .A(n22547), .X(n45019) );
  nand_x1_sg U53907 ( .A(n45797), .B(n26799), .X(n26798) );
  inv_x1_sg U53908 ( .A(n26801), .X(n45797) );
  inv_x1_sg U53909 ( .A(n26183), .X(n51470) );
  inv_x1_sg U53910 ( .A(n26193), .X(n51471) );
  inv_x1_sg U53911 ( .A(n26201), .X(n51472) );
  inv_x1_sg U53912 ( .A(n26209), .X(n51473) );
  inv_x1_sg U53913 ( .A(n26217), .X(n51474) );
  inv_x1_sg U53914 ( .A(n26225), .X(n51475) );
  inv_x1_sg U53915 ( .A(n26249), .X(n51478) );
  inv_x1_sg U53916 ( .A(n26265), .X(n51480) );
  inv_x1_sg U53917 ( .A(n26281), .X(n51482) );
  inv_x1_sg U53918 ( .A(n26297), .X(n51484) );
  inv_x1_sg U53919 ( .A(n26311), .X(n51486) );
  inv_x1_sg U53920 ( .A(n26319), .X(n51487) );
  inv_x1_sg U53921 ( .A(n26232), .X(n51476) );
  inv_x1_sg U53922 ( .A(n26240), .X(n51477) );
  inv_x1_sg U53923 ( .A(n26256), .X(n51479) );
  inv_x1_sg U53924 ( .A(n26272), .X(n51481) );
  inv_x1_sg U53925 ( .A(n26288), .X(n51483) );
  nand_x1_sg U53926 ( .A(n36925), .B(n36924), .X(n1990) );
  nand_x1_sg U53927 ( .A(n36949), .B(n36948), .X(n1978) );
  nand_x1_sg U53928 ( .A(n37405), .B(n37404), .X(n1750) );
  nand_x1_sg U53929 ( .A(n37429), .B(n37428), .X(n1738) );
  nand_x1_sg U53930 ( .A(n37549), .B(n37548), .X(n1658) );
  nand_x1_sg U53931 ( .A(n38029), .B(n38028), .X(n1418) );
  nand_x1_sg U53932 ( .A(n36916), .B(n36917), .X(n1994) );
  nand_x1_sg U53933 ( .A(n36918), .B(n36919), .X(n1993) );
  nand_x1_sg U53934 ( .A(n38118), .B(n38119), .X(n1353) );
  nand_x1_sg U53935 ( .A(n37522), .B(n37523), .X(n1671) );
  nand_x1_sg U53936 ( .A(n36946), .B(n36947), .X(n1979) );
  nand_x1_sg U53937 ( .A(n37396), .B(n37397), .X(n1754) );
  nand_x1_sg U53938 ( .A(n37398), .B(n37399), .X(n1753) );
  nand_x1_sg U53939 ( .A(n37426), .B(n37427), .X(n1739) );
  nand_x1_sg U53940 ( .A(n37546), .B(n37547), .X(n1659) );
  nand_x1_sg U53941 ( .A(n37998), .B(n37999), .X(n1433) );
  nand_x1_sg U53942 ( .A(n38026), .B(n38027), .X(n1419) );
  nand_x1_sg U53943 ( .A(n38112), .B(n38113), .X(n1356) );
  nand_x1_sg U53944 ( .A(n36922), .B(n36923), .X(n1991) );
  nand_x1_sg U53945 ( .A(n37518), .B(n37519), .X(n1673) );
  nand_x1_sg U53946 ( .A(n37524), .B(n37525), .X(n1670) );
  nand_x1_sg U53947 ( .A(n38004), .B(n38005), .X(n1430) );
  nand_x1_sg U53948 ( .A(n38116), .B(n38117), .X(n1354) );
  nand_x1_sg U53949 ( .A(n37520), .B(n37521), .X(n1672) );
  nand_x1_sg U53950 ( .A(n37996), .B(n37997), .X(n1434) );
  nand_x1_sg U53951 ( .A(n38000), .B(n38001), .X(n1432) );
  nand_x1_sg U53952 ( .A(n36912), .B(n36913), .X(n1996) );
  nand_x1_sg U53953 ( .A(n36950), .B(n36951), .X(n1977) );
  nand_x1_sg U53954 ( .A(n37392), .B(n37393), .X(n1756) );
  nand_x1_sg U53955 ( .A(n37430), .B(n37431), .X(n1737) );
  nand_x1_sg U53956 ( .A(n36909), .B(n36910), .X(n1997) );
  nand_x1_sg U53957 ( .A(n36914), .B(n36915), .X(n1995) );
  nand_x1_sg U53958 ( .A(n36920), .B(n36921), .X(n1992) );
  nand_x1_sg U53959 ( .A(n36926), .B(n36927), .X(n1989) );
  nand_x1_sg U53960 ( .A(n36928), .B(n36929), .X(n1988) );
  nand_x1_sg U53961 ( .A(n36930), .B(n36931), .X(n1987) );
  nand_x1_sg U53962 ( .A(n36932), .B(n36933), .X(n1986) );
  nand_x1_sg U53963 ( .A(n36934), .B(n36935), .X(n1985) );
  nand_x1_sg U53964 ( .A(n36936), .B(n36937), .X(n1984) );
  nand_x1_sg U53965 ( .A(n36938), .B(n36939), .X(n1983) );
  nand_x1_sg U53966 ( .A(n36940), .B(n36941), .X(n1982) );
  nand_x1_sg U53967 ( .A(n36942), .B(n36943), .X(n1981) );
  nand_x1_sg U53968 ( .A(n36944), .B(n36945), .X(n1980) );
  nand_x1_sg U53969 ( .A(n37394), .B(n37395), .X(n1755) );
  nand_x1_sg U53970 ( .A(n37400), .B(n37401), .X(n1752) );
  nand_x1_sg U53971 ( .A(n37402), .B(n37403), .X(n1751) );
  nand_x1_sg U53972 ( .A(n37406), .B(n37407), .X(n1749) );
  nand_x1_sg U53973 ( .A(n37408), .B(n37409), .X(n1748) );
  nand_x1_sg U53974 ( .A(n37410), .B(n37411), .X(n1747) );
  nand_x1_sg U53975 ( .A(n37412), .B(n37413), .X(n1746) );
  nand_x1_sg U53976 ( .A(n37414), .B(n37415), .X(n1745) );
  nand_x1_sg U53977 ( .A(n37416), .B(n37417), .X(n1744) );
  nand_x1_sg U53978 ( .A(n37418), .B(n37419), .X(n1743) );
  nand_x1_sg U53979 ( .A(n37420), .B(n37421), .X(n1742) );
  nand_x1_sg U53980 ( .A(n37422), .B(n37423), .X(n1741) );
  nand_x1_sg U53981 ( .A(n37424), .B(n37425), .X(n1740) );
  nand_x1_sg U53982 ( .A(n37512), .B(n37513), .X(n1676) );
  nand_x1_sg U53983 ( .A(n37514), .B(n37515), .X(n1675) );
  nand_x1_sg U53984 ( .A(n37516), .B(n37517), .X(n1674) );
  nand_x1_sg U53985 ( .A(n37526), .B(n37527), .X(n1669) );
  nand_x1_sg U53986 ( .A(n37528), .B(n37529), .X(n1668) );
  nand_x1_sg U53987 ( .A(n37530), .B(n37531), .X(n1667) );
  nand_x1_sg U53988 ( .A(n37532), .B(n37533), .X(n1666) );
  nand_x1_sg U53989 ( .A(n37534), .B(n37535), .X(n1665) );
  nand_x1_sg U53990 ( .A(n37536), .B(n37537), .X(n1664) );
  nand_x1_sg U53991 ( .A(n37538), .B(n37539), .X(n1663) );
  nand_x1_sg U53992 ( .A(n37540), .B(n37541), .X(n1662) );
  nand_x1_sg U53993 ( .A(n37542), .B(n37543), .X(n1661) );
  nand_x1_sg U53994 ( .A(n37544), .B(n37545), .X(n1660) );
  nand_x1_sg U53995 ( .A(n37550), .B(n37551), .X(n1657) );
  nand_x1_sg U53996 ( .A(n37992), .B(n37993), .X(n1436) );
  nand_x1_sg U53997 ( .A(n37994), .B(n37995), .X(n1435) );
  nand_x1_sg U53998 ( .A(n38002), .B(n38003), .X(n1431) );
  nand_x1_sg U53999 ( .A(n38006), .B(n38007), .X(n1429) );
  nand_x1_sg U54000 ( .A(n38008), .B(n38009), .X(n1428) );
  nand_x1_sg U54001 ( .A(n38010), .B(n38011), .X(n1427) );
  nand_x1_sg U54002 ( .A(n38012), .B(n38013), .X(n1426) );
  nand_x1_sg U54003 ( .A(n38014), .B(n38015), .X(n1425) );
  nand_x1_sg U54004 ( .A(n38016), .B(n38017), .X(n1424) );
  nand_x1_sg U54005 ( .A(n38018), .B(n38019), .X(n1423) );
  nand_x1_sg U54006 ( .A(n38020), .B(n38021), .X(n1422) );
  nand_x1_sg U54007 ( .A(n38022), .B(n38023), .X(n1421) );
  nand_x1_sg U54008 ( .A(n38024), .B(n38025), .X(n1420) );
  nand_x1_sg U54009 ( .A(n38030), .B(n38031), .X(n1417) );
  nand_x1_sg U54010 ( .A(n38114), .B(n38115), .X(n1355) );
  nand_x1_sg U54011 ( .A(n36964), .B(n36965), .X(n1970) );
  nand_x1_sg U54012 ( .A(n37004), .B(n37005), .X(n1950) );
  nand_x1_sg U54013 ( .A(n37084), .B(n37085), .X(n1910) );
  nand_x1_sg U54014 ( .A(n37164), .B(n37165), .X(n1870) );
  nand_x1_sg U54015 ( .A(n37204), .B(n37205), .X(n1850) );
  nand_x1_sg U54016 ( .A(n37244), .B(n37245), .X(n1830) );
  nand_x1_sg U54017 ( .A(n37284), .B(n37285), .X(n1810) );
  nand_x1_sg U54018 ( .A(n37324), .B(n37325), .X(n1790) );
  nand_x1_sg U54019 ( .A(n37444), .B(n37445), .X(n1730) );
  nand_x1_sg U54020 ( .A(n37484), .B(n37485), .X(n1710) );
  nand_x1_sg U54021 ( .A(n36956), .B(n36957), .X(n1974) );
  nand_x1_sg U54022 ( .A(n36958), .B(n36959), .X(n1973) );
  nand_x1_sg U54023 ( .A(n36996), .B(n36997), .X(n1954) );
  nand_x1_sg U54024 ( .A(n36998), .B(n36999), .X(n1953) );
  nand_x1_sg U54025 ( .A(n37076), .B(n37077), .X(n1914) );
  nand_x1_sg U54026 ( .A(n37078), .B(n37079), .X(n1913) );
  nand_x1_sg U54027 ( .A(n37116), .B(n37117), .X(n1894) );
  nand_x1_sg U54028 ( .A(n37118), .B(n37119), .X(n1893) );
  nand_x1_sg U54029 ( .A(n37156), .B(n37157), .X(n1874) );
  nand_x1_sg U54030 ( .A(n37158), .B(n37159), .X(n1873) );
  nand_x1_sg U54031 ( .A(n37196), .B(n37197), .X(n1854) );
  nand_x1_sg U54032 ( .A(n37198), .B(n37199), .X(n1853) );
  nand_x1_sg U54033 ( .A(n37236), .B(n37237), .X(n1834) );
  nand_x1_sg U54034 ( .A(n37238), .B(n37239), .X(n1833) );
  nand_x1_sg U54035 ( .A(n37276), .B(n37277), .X(n1814) );
  nand_x1_sg U54036 ( .A(n37278), .B(n37279), .X(n1813) );
  nand_x1_sg U54037 ( .A(n37316), .B(n37317), .X(n1794) );
  nand_x1_sg U54038 ( .A(n37318), .B(n37319), .X(n1793) );
  nand_x1_sg U54039 ( .A(n37436), .B(n37437), .X(n1734) );
  nand_x1_sg U54040 ( .A(n37438), .B(n37439), .X(n1733) );
  nand_x1_sg U54041 ( .A(n37476), .B(n37477), .X(n1714) );
  nand_x1_sg U54042 ( .A(n37478), .B(n37479), .X(n1713) );
  nand_x1_sg U54043 ( .A(n36952), .B(n36953), .X(n1976) );
  nand_x1_sg U54044 ( .A(n36990), .B(n36991), .X(n1957) );
  nand_x1_sg U54045 ( .A(n36992), .B(n36993), .X(n1956) );
  nand_x1_sg U54046 ( .A(n37070), .B(n37071), .X(n1917) );
  nand_x1_sg U54047 ( .A(n37072), .B(n37073), .X(n1916) );
  nand_x1_sg U54048 ( .A(n37110), .B(n37111), .X(n1897) );
  nand_x1_sg U54049 ( .A(n37112), .B(n37113), .X(n1896) );
  nand_x1_sg U54050 ( .A(n37150), .B(n37151), .X(n1877) );
  nand_x1_sg U54051 ( .A(n37152), .B(n37153), .X(n1876) );
  nand_x1_sg U54052 ( .A(n37190), .B(n37191), .X(n1857) );
  nand_x1_sg U54053 ( .A(n37192), .B(n37193), .X(n1856) );
  nand_x1_sg U54054 ( .A(n37230), .B(n37231), .X(n1837) );
  nand_x1_sg U54055 ( .A(n37232), .B(n37233), .X(n1836) );
  nand_x1_sg U54056 ( .A(n37270), .B(n37271), .X(n1817) );
  nand_x1_sg U54057 ( .A(n37272), .B(n37273), .X(n1816) );
  nand_x1_sg U54058 ( .A(n37310), .B(n37311), .X(n1797) );
  nand_x1_sg U54059 ( .A(n37312), .B(n37313), .X(n1796) );
  nand_x1_sg U54060 ( .A(n37390), .B(n37391), .X(n1757) );
  nand_x1_sg U54061 ( .A(n37432), .B(n37433), .X(n1736) );
  nand_x1_sg U54062 ( .A(n37470), .B(n37471), .X(n1717) );
  nand_x1_sg U54063 ( .A(n37472), .B(n37473), .X(n1716) );
  nand_x1_sg U54064 ( .A(n37510), .B(n37511), .X(n1697) );
  nand_x1_sg U54065 ( .A(n36954), .B(n36955), .X(n1975) );
  nand_x1_sg U54066 ( .A(n36994), .B(n36995), .X(n1955) );
  nand_x1_sg U54067 ( .A(n37074), .B(n37075), .X(n1915) );
  nand_x1_sg U54068 ( .A(n37114), .B(n37115), .X(n1895) );
  nand_x1_sg U54069 ( .A(n37154), .B(n37155), .X(n1875) );
  nand_x1_sg U54070 ( .A(n37194), .B(n37195), .X(n1855) );
  nand_x1_sg U54071 ( .A(n37234), .B(n37235), .X(n1835) );
  nand_x1_sg U54072 ( .A(n37274), .B(n37275), .X(n1815) );
  nand_x1_sg U54073 ( .A(n37314), .B(n37315), .X(n1795) );
  nand_x1_sg U54074 ( .A(n37434), .B(n37435), .X(n1735) );
  nand_x1_sg U54075 ( .A(n37474), .B(n37475), .X(n1715) );
  nand_x1_sg U54076 ( .A(n36960), .B(n36961), .X(n1972) );
  nand_x1_sg U54077 ( .A(n36966), .B(n36967), .X(n1969) );
  nand_x1_sg U54078 ( .A(n36968), .B(n36969), .X(n1968) );
  nand_x1_sg U54079 ( .A(n36970), .B(n36971), .X(n1967) );
  nand_x1_sg U54080 ( .A(n36972), .B(n36973), .X(n1966) );
  nand_x1_sg U54081 ( .A(n36974), .B(n36975), .X(n1965) );
  nand_x1_sg U54082 ( .A(n36976), .B(n36977), .X(n1964) );
  nand_x1_sg U54083 ( .A(n36978), .B(n36979), .X(n1963) );
  nand_x1_sg U54084 ( .A(n36980), .B(n36981), .X(n1962) );
  nand_x1_sg U54085 ( .A(n36982), .B(n36983), .X(n1961) );
  nand_x1_sg U54086 ( .A(n36984), .B(n36985), .X(n1960) );
  nand_x1_sg U54087 ( .A(n37000), .B(n37001), .X(n1952) );
  nand_x1_sg U54088 ( .A(n37006), .B(n37007), .X(n1949) );
  nand_x1_sg U54089 ( .A(n37008), .B(n37009), .X(n1948) );
  nand_x1_sg U54090 ( .A(n37010), .B(n37011), .X(n1947) );
  nand_x1_sg U54091 ( .A(n37012), .B(n37013), .X(n1946) );
  nand_x1_sg U54092 ( .A(n37014), .B(n37015), .X(n1945) );
  nand_x1_sg U54093 ( .A(n37016), .B(n37017), .X(n1944) );
  nand_x1_sg U54094 ( .A(n37018), .B(n37019), .X(n1943) );
  nand_x1_sg U54095 ( .A(n37020), .B(n37021), .X(n1942) );
  nand_x1_sg U54096 ( .A(n37022), .B(n37023), .X(n1941) );
  nand_x1_sg U54097 ( .A(n37024), .B(n37025), .X(n1940) );
  nand_x1_sg U54098 ( .A(n37080), .B(n37081), .X(n1912) );
  nand_x1_sg U54099 ( .A(n37086), .B(n37087), .X(n1909) );
  nand_x1_sg U54100 ( .A(n37088), .B(n37089), .X(n1908) );
  nand_x1_sg U54101 ( .A(n37090), .B(n37091), .X(n1907) );
  nand_x1_sg U54102 ( .A(n37092), .B(n37093), .X(n1906) );
  nand_x1_sg U54103 ( .A(n37094), .B(n37095), .X(n1905) );
  nand_x1_sg U54104 ( .A(n37096), .B(n37097), .X(n1904) );
  nand_x1_sg U54105 ( .A(n37098), .B(n37099), .X(n1903) );
  nand_x1_sg U54106 ( .A(n37100), .B(n37101), .X(n1902) );
  nand_x1_sg U54107 ( .A(n37102), .B(n37103), .X(n1901) );
  nand_x1_sg U54108 ( .A(n37104), .B(n37105), .X(n1900) );
  nand_x1_sg U54109 ( .A(n37130), .B(n37131), .X(n1887) );
  nand_x1_sg U54110 ( .A(n37132), .B(n37133), .X(n1886) );
  nand_x1_sg U54111 ( .A(n37134), .B(n37135), .X(n1885) );
  nand_x1_sg U54112 ( .A(n37136), .B(n37137), .X(n1884) );
  nand_x1_sg U54113 ( .A(n37138), .B(n37139), .X(n1883) );
  nand_x1_sg U54114 ( .A(n37140), .B(n37141), .X(n1882) );
  nand_x1_sg U54115 ( .A(n37142), .B(n37143), .X(n1881) );
  nand_x1_sg U54116 ( .A(n37144), .B(n37145), .X(n1880) );
  nand_x1_sg U54117 ( .A(n37160), .B(n37161), .X(n1872) );
  nand_x1_sg U54118 ( .A(n37166), .B(n37167), .X(n1869) );
  nand_x1_sg U54119 ( .A(n37168), .B(n37169), .X(n1868) );
  nand_x1_sg U54120 ( .A(n37170), .B(n37171), .X(n1867) );
  nand_x1_sg U54121 ( .A(n37172), .B(n37173), .X(n1866) );
  nand_x1_sg U54122 ( .A(n37174), .B(n37175), .X(n1865) );
  nand_x1_sg U54123 ( .A(n37176), .B(n37177), .X(n1864) );
  nand_x1_sg U54124 ( .A(n37178), .B(n37179), .X(n1863) );
  nand_x1_sg U54125 ( .A(n37180), .B(n37181), .X(n1862) );
  nand_x1_sg U54126 ( .A(n37182), .B(n37183), .X(n1861) );
  nand_x1_sg U54127 ( .A(n37184), .B(n37185), .X(n1860) );
  nand_x1_sg U54128 ( .A(n37200), .B(n37201), .X(n1852) );
  nand_x1_sg U54129 ( .A(n37206), .B(n37207), .X(n1849) );
  nand_x1_sg U54130 ( .A(n37208), .B(n37209), .X(n1848) );
  nand_x1_sg U54131 ( .A(n37210), .B(n37211), .X(n1847) );
  nand_x1_sg U54132 ( .A(n37212), .B(n37213), .X(n1846) );
  nand_x1_sg U54133 ( .A(n37214), .B(n37215), .X(n1845) );
  nand_x1_sg U54134 ( .A(n37216), .B(n37217), .X(n1844) );
  nand_x1_sg U54135 ( .A(n37218), .B(n37219), .X(n1843) );
  nand_x1_sg U54136 ( .A(n37220), .B(n37221), .X(n1842) );
  nand_x1_sg U54137 ( .A(n37222), .B(n37223), .X(n1841) );
  nand_x1_sg U54138 ( .A(n37224), .B(n37225), .X(n1840) );
  nand_x1_sg U54139 ( .A(n37240), .B(n37241), .X(n1832) );
  nand_x1_sg U54140 ( .A(n37246), .B(n37247), .X(n1829) );
  nand_x1_sg U54141 ( .A(n37248), .B(n37249), .X(n1828) );
  nand_x1_sg U54142 ( .A(n37250), .B(n37251), .X(n1827) );
  nand_x1_sg U54143 ( .A(n37252), .B(n37253), .X(n1826) );
  nand_x1_sg U54144 ( .A(n37254), .B(n37255), .X(n1825) );
  nand_x1_sg U54145 ( .A(n37256), .B(n37257), .X(n1824) );
  nand_x1_sg U54146 ( .A(n37258), .B(n37259), .X(n1823) );
  nand_x1_sg U54147 ( .A(n37260), .B(n37261), .X(n1822) );
  nand_x1_sg U54148 ( .A(n37262), .B(n37263), .X(n1821) );
  nand_x1_sg U54149 ( .A(n37264), .B(n37265), .X(n1820) );
  nand_x1_sg U54150 ( .A(n37280), .B(n37281), .X(n1812) );
  nand_x1_sg U54151 ( .A(n37286), .B(n37287), .X(n1809) );
  nand_x1_sg U54152 ( .A(n37288), .B(n37289), .X(n1808) );
  nand_x1_sg U54153 ( .A(n37290), .B(n37291), .X(n1807) );
  nand_x1_sg U54154 ( .A(n37292), .B(n37293), .X(n1806) );
  nand_x1_sg U54155 ( .A(n37294), .B(n37295), .X(n1805) );
  nand_x1_sg U54156 ( .A(n37296), .B(n37297), .X(n1804) );
  nand_x1_sg U54157 ( .A(n37298), .B(n37299), .X(n1803) );
  nand_x1_sg U54158 ( .A(n37300), .B(n37301), .X(n1802) );
  nand_x1_sg U54159 ( .A(n37302), .B(n37303), .X(n1801) );
  nand_x1_sg U54160 ( .A(n37304), .B(n37305), .X(n1800) );
  nand_x1_sg U54161 ( .A(n37320), .B(n37321), .X(n1792) );
  nand_x1_sg U54162 ( .A(n37326), .B(n37327), .X(n1789) );
  nand_x1_sg U54163 ( .A(n37328), .B(n37329), .X(n1788) );
  nand_x1_sg U54164 ( .A(n37330), .B(n37331), .X(n1787) );
  nand_x1_sg U54165 ( .A(n37332), .B(n37333), .X(n1786) );
  nand_x1_sg U54166 ( .A(n37334), .B(n37335), .X(n1785) );
  nand_x1_sg U54167 ( .A(n37336), .B(n37337), .X(n1784) );
  nand_x1_sg U54168 ( .A(n37338), .B(n37339), .X(n1783) );
  nand_x1_sg U54169 ( .A(n37440), .B(n37441), .X(n1732) );
  nand_x1_sg U54170 ( .A(n37446), .B(n37447), .X(n1729) );
  nand_x1_sg U54171 ( .A(n37448), .B(n37449), .X(n1728) );
  nand_x1_sg U54172 ( .A(n37450), .B(n37451), .X(n1727) );
  nand_x1_sg U54173 ( .A(n37452), .B(n37453), .X(n1726) );
  nand_x1_sg U54174 ( .A(n37454), .B(n37455), .X(n1725) );
  nand_x1_sg U54175 ( .A(n37456), .B(n37457), .X(n1724) );
  nand_x1_sg U54176 ( .A(n37458), .B(n37459), .X(n1723) );
  nand_x1_sg U54177 ( .A(n37460), .B(n37461), .X(n1722) );
  nand_x1_sg U54178 ( .A(n37462), .B(n37463), .X(n1721) );
  nand_x1_sg U54179 ( .A(n37464), .B(n37465), .X(n1720) );
  nand_x1_sg U54180 ( .A(n37480), .B(n37481), .X(n1712) );
  nand_x1_sg U54181 ( .A(n37486), .B(n37487), .X(n1709) );
  nand_x1_sg U54182 ( .A(n37488), .B(n37489), .X(n1708) );
  nand_x1_sg U54183 ( .A(n37490), .B(n37491), .X(n1707) );
  nand_x1_sg U54184 ( .A(n37492), .B(n37493), .X(n1706) );
  nand_x1_sg U54185 ( .A(n37494), .B(n37495), .X(n1705) );
  nand_x1_sg U54186 ( .A(n37496), .B(n37497), .X(n1704) );
  nand_x1_sg U54187 ( .A(n37498), .B(n37499), .X(n1703) );
  nand_x1_sg U54188 ( .A(n37500), .B(n37501), .X(n1702) );
  nand_x1_sg U54189 ( .A(n37502), .B(n37503), .X(n1701) );
  nand_x1_sg U54190 ( .A(n37504), .B(n37505), .X(n1700) );
  nand_x1_sg U54191 ( .A(n37554), .B(n37555), .X(n1655) );
  nand_x1_sg U54192 ( .A(n37556), .B(n37557), .X(n1654) );
  nand_x1_sg U54193 ( .A(n37566), .B(n37567), .X(n1649) );
  nand_x1_sg U54194 ( .A(n37568), .B(n37569), .X(n1648) );
  nand_x1_sg U54195 ( .A(n37570), .B(n37571), .X(n1647) );
  nand_x1_sg U54196 ( .A(n37572), .B(n37573), .X(n1646) );
  nand_x1_sg U54197 ( .A(n37574), .B(n37575), .X(n1645) );
  nand_x1_sg U54198 ( .A(n37576), .B(n37577), .X(n1644) );
  nand_x1_sg U54199 ( .A(n37578), .B(n37579), .X(n1643) );
  nand_x1_sg U54200 ( .A(n37580), .B(n37581), .X(n1642) );
  nand_x1_sg U54201 ( .A(n37582), .B(n37583), .X(n1641) );
  nand_x1_sg U54202 ( .A(n37584), .B(n37585), .X(n1640) );
  nand_x1_sg U54203 ( .A(n37594), .B(n37595), .X(n1635) );
  nand_x1_sg U54204 ( .A(n37596), .B(n37597), .X(n1634) );
  nand_x1_sg U54205 ( .A(n37650), .B(n37651), .X(n1607) );
  nand_x1_sg U54206 ( .A(n37652), .B(n37653), .X(n1606) );
  nand_x1_sg U54207 ( .A(n37654), .B(n37655), .X(n1605) );
  nand_x1_sg U54208 ( .A(n37656), .B(n37657), .X(n1604) );
  nand_x1_sg U54209 ( .A(n37658), .B(n37659), .X(n1603) );
  nand_x1_sg U54210 ( .A(n37660), .B(n37661), .X(n1602) );
  nand_x1_sg U54211 ( .A(n37662), .B(n37663), .X(n1601) );
  nand_x1_sg U54212 ( .A(n37664), .B(n37665), .X(n1600) );
  nand_x1_sg U54213 ( .A(n37674), .B(n37675), .X(n1595) );
  nand_x1_sg U54214 ( .A(n37676), .B(n37677), .X(n1594) );
  nand_x1_sg U54215 ( .A(n37686), .B(n37687), .X(n1589) );
  nand_x1_sg U54216 ( .A(n37688), .B(n37689), .X(n1588) );
  nand_x1_sg U54217 ( .A(n37690), .B(n37691), .X(n1587) );
  nand_x1_sg U54218 ( .A(n37692), .B(n37693), .X(n1586) );
  nand_x1_sg U54219 ( .A(n37694), .B(n37695), .X(n1585) );
  nand_x1_sg U54220 ( .A(n37696), .B(n37697), .X(n1584) );
  nand_x1_sg U54221 ( .A(n37698), .B(n37699), .X(n1583) );
  nand_x1_sg U54222 ( .A(n37700), .B(n37701), .X(n1582) );
  nand_x1_sg U54223 ( .A(n37702), .B(n37703), .X(n1581) );
  nand_x1_sg U54224 ( .A(n37704), .B(n37705), .X(n1580) );
  nand_x1_sg U54225 ( .A(n37754), .B(n37755), .X(n1555) );
  nand_x1_sg U54226 ( .A(n37756), .B(n37757), .X(n1554) );
  nand_x1_sg U54227 ( .A(n37766), .B(n37767), .X(n1549) );
  nand_x1_sg U54228 ( .A(n37768), .B(n37769), .X(n1548) );
  nand_x1_sg U54229 ( .A(n37770), .B(n37771), .X(n1547) );
  nand_x1_sg U54230 ( .A(n37772), .B(n37773), .X(n1546) );
  nand_x1_sg U54231 ( .A(n37774), .B(n37775), .X(n1545) );
  nand_x1_sg U54232 ( .A(n37776), .B(n37777), .X(n1544) );
  nand_x1_sg U54233 ( .A(n37778), .B(n37779), .X(n1543) );
  nand_x1_sg U54234 ( .A(n37780), .B(n37781), .X(n1542) );
  nand_x1_sg U54235 ( .A(n37782), .B(n37783), .X(n1541) );
  nand_x1_sg U54236 ( .A(n37784), .B(n37785), .X(n1540) );
  nand_x1_sg U54237 ( .A(n37794), .B(n37795), .X(n1535) );
  nand_x1_sg U54238 ( .A(n37796), .B(n37797), .X(n1534) );
  nand_x1_sg U54239 ( .A(n37806), .B(n37807), .X(n1529) );
  nand_x1_sg U54240 ( .A(n37808), .B(n37809), .X(n1528) );
  nand_x1_sg U54241 ( .A(n37810), .B(n37811), .X(n1527) );
  nand_x1_sg U54242 ( .A(n37812), .B(n37813), .X(n1526) );
  nand_x1_sg U54243 ( .A(n37814), .B(n37815), .X(n1525) );
  nand_x1_sg U54244 ( .A(n37816), .B(n37817), .X(n1524) );
  nand_x1_sg U54245 ( .A(n37818), .B(n37819), .X(n1523) );
  nand_x1_sg U54246 ( .A(n37820), .B(n37821), .X(n1522) );
  nand_x1_sg U54247 ( .A(n37822), .B(n37823), .X(n1521) );
  nand_x1_sg U54248 ( .A(n37824), .B(n37825), .X(n1520) );
  nand_x1_sg U54249 ( .A(n37834), .B(n37835), .X(n1515) );
  nand_x1_sg U54250 ( .A(n37836), .B(n37837), .X(n1514) );
  nand_x1_sg U54251 ( .A(n37846), .B(n37847), .X(n1509) );
  nand_x1_sg U54252 ( .A(n37848), .B(n37849), .X(n1508) );
  nand_x1_sg U54253 ( .A(n37850), .B(n37851), .X(n1507) );
  nand_x1_sg U54254 ( .A(n37852), .B(n37853), .X(n1506) );
  nand_x1_sg U54255 ( .A(n37854), .B(n37855), .X(n1505) );
  nand_x1_sg U54256 ( .A(n37856), .B(n37857), .X(n1504) );
  nand_x1_sg U54257 ( .A(n37858), .B(n37859), .X(n1503) );
  nand_x1_sg U54258 ( .A(n37926), .B(n37927), .X(n1469) );
  nand_x1_sg U54259 ( .A(n37928), .B(n37929), .X(n1468) );
  nand_x1_sg U54260 ( .A(n37930), .B(n37931), .X(n1467) );
  nand_x1_sg U54261 ( .A(n37932), .B(n37933), .X(n1466) );
  nand_x1_sg U54262 ( .A(n37934), .B(n37935), .X(n1465) );
  nand_x1_sg U54263 ( .A(n37936), .B(n37937), .X(n1464) );
  nand_x1_sg U54264 ( .A(n37938), .B(n37939), .X(n1463) );
  nand_x1_sg U54265 ( .A(n37940), .B(n37941), .X(n1462) );
  nand_x1_sg U54266 ( .A(n37942), .B(n37943), .X(n1461) );
  nand_x1_sg U54267 ( .A(n37944), .B(n37945), .X(n1460) );
  nand_x1_sg U54268 ( .A(n37954), .B(n37955), .X(n1455) );
  nand_x1_sg U54269 ( .A(n37956), .B(n37957), .X(n1454) );
  nand_x1_sg U54270 ( .A(n37966), .B(n37967), .X(n1449) );
  nand_x1_sg U54271 ( .A(n37968), .B(n37969), .X(n1448) );
  nand_x1_sg U54272 ( .A(n37970), .B(n37971), .X(n1447) );
  nand_x1_sg U54273 ( .A(n37972), .B(n37973), .X(n1446) );
  nand_x1_sg U54274 ( .A(n37974), .B(n37975), .X(n1445) );
  nand_x1_sg U54275 ( .A(n37976), .B(n37977), .X(n1444) );
  nand_x1_sg U54276 ( .A(n37978), .B(n37979), .X(n1443) );
  nand_x1_sg U54277 ( .A(n37980), .B(n37981), .X(n1442) );
  nand_x1_sg U54278 ( .A(n37982), .B(n37983), .X(n1441) );
  nand_x1_sg U54279 ( .A(n37984), .B(n37985), .X(n1440) );
  nand_x1_sg U54280 ( .A(n38034), .B(n38035), .X(n1415) );
  nand_x1_sg U54281 ( .A(n38036), .B(n38037), .X(n1414) );
  nand_x1_sg U54282 ( .A(n38046), .B(n38047), .X(n1409) );
  nand_x1_sg U54283 ( .A(n38048), .B(n38049), .X(n1408) );
  nand_x1_sg U54284 ( .A(n38050), .B(n38051), .X(n1407) );
  nand_x1_sg U54285 ( .A(n38052), .B(n38053), .X(n1406) );
  nand_x1_sg U54286 ( .A(n38054), .B(n38055), .X(n1405) );
  nand_x1_sg U54287 ( .A(n38056), .B(n38057), .X(n1404) );
  nand_x1_sg U54288 ( .A(n38058), .B(n38059), .X(n1403) );
  nand_x1_sg U54289 ( .A(n38060), .B(n38061), .X(n1402) );
  nand_x1_sg U54290 ( .A(n38062), .B(n38063), .X(n1401) );
  nand_x1_sg U54291 ( .A(n38064), .B(n38065), .X(n1400) );
  nand_x1_sg U54292 ( .A(n38074), .B(n38075), .X(n1395) );
  nand_x1_sg U54293 ( .A(n38076), .B(n38077), .X(n1394) );
  nand_x1_sg U54294 ( .A(n38086), .B(n38087), .X(n1389) );
  nand_x1_sg U54295 ( .A(n38088), .B(n38089), .X(n1388) );
  nand_x1_sg U54296 ( .A(n38090), .B(n38091), .X(n1387) );
  nand_x1_sg U54297 ( .A(n38092), .B(n38093), .X(n1386) );
  nand_x1_sg U54298 ( .A(n38094), .B(n38095), .X(n1385) );
  nand_x1_sg U54299 ( .A(n38096), .B(n38097), .X(n1384) );
  nand_x1_sg U54300 ( .A(n38098), .B(n38099), .X(n1383) );
  nand_x1_sg U54301 ( .A(n38100), .B(n38101), .X(n1382) );
  nand_x1_sg U54302 ( .A(n38102), .B(n38103), .X(n1381) );
  nand_x1_sg U54303 ( .A(n38104), .B(n38105), .X(n1380) );
  nand_x1_sg U54304 ( .A(n36988), .B(n36989), .X(n1958) );
  nand_x1_sg U54305 ( .A(n37028), .B(n37029), .X(n1938) );
  nand_x1_sg U54306 ( .A(n37108), .B(n37109), .X(n1898) );
  nand_x1_sg U54307 ( .A(n37148), .B(n37149), .X(n1878) );
  nand_x1_sg U54308 ( .A(n37188), .B(n37189), .X(n1858) );
  nand_x1_sg U54309 ( .A(n37228), .B(n37229), .X(n1838) );
  nand_x1_sg U54310 ( .A(n37268), .B(n37269), .X(n1818) );
  nand_x1_sg U54311 ( .A(n37308), .B(n37309), .X(n1798) );
  nand_x1_sg U54312 ( .A(n37468), .B(n37469), .X(n1718) );
  nand_x1_sg U54313 ( .A(n37508), .B(n37509), .X(n1698) );
  nand_x1_sg U54314 ( .A(n37552), .B(n37553), .X(n1656) );
  nand_x1_sg U54315 ( .A(n37590), .B(n37591), .X(n1637) );
  nand_x1_sg U54316 ( .A(n37592), .B(n37593), .X(n1636) );
  nand_x1_sg U54317 ( .A(n37670), .B(n37671), .X(n1597) );
  nand_x1_sg U54318 ( .A(n37672), .B(n37673), .X(n1596) );
  nand_x1_sg U54319 ( .A(n37750), .B(n37751), .X(n1557) );
  nand_x1_sg U54320 ( .A(n37752), .B(n37753), .X(n1556) );
  nand_x1_sg U54321 ( .A(n37790), .B(n37791), .X(n1537) );
  nand_x1_sg U54322 ( .A(n37792), .B(n37793), .X(n1536) );
  nand_x1_sg U54323 ( .A(n37830), .B(n37831), .X(n1517) );
  nand_x1_sg U54324 ( .A(n37832), .B(n37833), .X(n1516) );
  nand_x1_sg U54325 ( .A(n37950), .B(n37951), .X(n1457) );
  nand_x1_sg U54326 ( .A(n37952), .B(n37953), .X(n1456) );
  nand_x1_sg U54327 ( .A(n37990), .B(n37991), .X(n1437) );
  nand_x1_sg U54328 ( .A(n38032), .B(n38033), .X(n1416) );
  nand_x1_sg U54329 ( .A(n38070), .B(n38071), .X(n1397) );
  nand_x1_sg U54330 ( .A(n38072), .B(n38073), .X(n1396) );
  nand_x1_sg U54331 ( .A(n38110), .B(n38111), .X(n1377) );
  nand_x1_sg U54332 ( .A(n36962), .B(n36963), .X(n1971) );
  nand_x1_sg U54333 ( .A(n36986), .B(n36987), .X(n1959) );
  nand_x1_sg U54334 ( .A(n37002), .B(n37003), .X(n1951) );
  nand_x1_sg U54335 ( .A(n37026), .B(n37027), .X(n1939) );
  nand_x1_sg U54336 ( .A(n37082), .B(n37083), .X(n1911) );
  nand_x1_sg U54337 ( .A(n37106), .B(n37107), .X(n1899) );
  nand_x1_sg U54338 ( .A(n37186), .B(n37187), .X(n1859) );
  nand_x1_sg U54339 ( .A(n37202), .B(n37203), .X(n1851) );
  nand_x1_sg U54340 ( .A(n37226), .B(n37227), .X(n1839) );
  nand_x1_sg U54341 ( .A(n37242), .B(n37243), .X(n1831) );
  nand_x1_sg U54342 ( .A(n37266), .B(n37267), .X(n1819) );
  nand_x1_sg U54343 ( .A(n37282), .B(n37283), .X(n1811) );
  nand_x1_sg U54344 ( .A(n37306), .B(n37307), .X(n1799) );
  nand_x1_sg U54345 ( .A(n37322), .B(n37323), .X(n1791) );
  nand_x1_sg U54346 ( .A(n37442), .B(n37443), .X(n1731) );
  nand_x1_sg U54347 ( .A(n37466), .B(n37467), .X(n1719) );
  nand_x1_sg U54348 ( .A(n37482), .B(n37483), .X(n1711) );
  nand_x1_sg U54349 ( .A(n37506), .B(n37507), .X(n1699) );
  nand_x1_sg U54350 ( .A(n37558), .B(n37559), .X(n1653) );
  nand_x1_sg U54351 ( .A(n37560), .B(n37561), .X(n1652) );
  nand_x1_sg U54352 ( .A(n37562), .B(n37563), .X(n1651) );
  nand_x1_sg U54353 ( .A(n37564), .B(n37565), .X(n1650) );
  nand_x1_sg U54354 ( .A(n37586), .B(n37587), .X(n1639) );
  nand_x1_sg U54355 ( .A(n37588), .B(n37589), .X(n1638) );
  nand_x1_sg U54356 ( .A(n37598), .B(n37599), .X(n1633) );
  nand_x1_sg U54357 ( .A(n37706), .B(n37707), .X(n1579) );
  nand_x1_sg U54358 ( .A(n37708), .B(n37709), .X(n1578) );
  nand_x1_sg U54359 ( .A(n37758), .B(n37759), .X(n1553) );
  nand_x1_sg U54360 ( .A(n37760), .B(n37761), .X(n1552) );
  nand_x1_sg U54361 ( .A(n37762), .B(n37763), .X(n1551) );
  nand_x1_sg U54362 ( .A(n37764), .B(n37765), .X(n1550) );
  nand_x1_sg U54363 ( .A(n37786), .B(n37787), .X(n1539) );
  nand_x1_sg U54364 ( .A(n37788), .B(n37789), .X(n1538) );
  nand_x1_sg U54365 ( .A(n37798), .B(n37799), .X(n1533) );
  nand_x1_sg U54366 ( .A(n37800), .B(n37801), .X(n1532) );
  nand_x1_sg U54367 ( .A(n37802), .B(n37803), .X(n1531) );
  nand_x1_sg U54368 ( .A(n37804), .B(n37805), .X(n1530) );
  nand_x1_sg U54369 ( .A(n37826), .B(n37827), .X(n1519) );
  nand_x1_sg U54370 ( .A(n37828), .B(n37829), .X(n1518) );
  nand_x1_sg U54371 ( .A(n37838), .B(n37839), .X(n1513) );
  nand_x1_sg U54372 ( .A(n37840), .B(n37841), .X(n1512) );
  nand_x1_sg U54373 ( .A(n37842), .B(n37843), .X(n1511) );
  nand_x1_sg U54374 ( .A(n37844), .B(n37845), .X(n1510) );
  nand_x1_sg U54375 ( .A(n37958), .B(n37959), .X(n1453) );
  nand_x1_sg U54376 ( .A(n38038), .B(n38039), .X(n1413) );
  nand_x1_sg U54377 ( .A(n38040), .B(n38041), .X(n1412) );
  nand_x1_sg U54378 ( .A(n38042), .B(n38043), .X(n1411) );
  nand_x1_sg U54379 ( .A(n38044), .B(n38045), .X(n1410) );
  nand_x1_sg U54380 ( .A(n38066), .B(n38067), .X(n1399) );
  nand_x1_sg U54381 ( .A(n38068), .B(n38069), .X(n1398) );
  nand_x1_sg U54382 ( .A(n38078), .B(n38079), .X(n1393) );
  nand_x1_sg U54383 ( .A(n38080), .B(n38081), .X(n1392) );
  nand_x1_sg U54384 ( .A(n38082), .B(n38083), .X(n1391) );
  nand_x1_sg U54385 ( .A(n38084), .B(n38085), .X(n1390) );
  nand_x1_sg U54386 ( .A(n38106), .B(n38107), .X(n1379) );
  nand_x1_sg U54387 ( .A(n38108), .B(n38109), .X(n1378) );
  nand_x1_sg U54388 ( .A(n37146), .B(n37147), .X(n1879) );
  nand_x1_sg U54389 ( .A(n37162), .B(n37163), .X(n1871) );
  nand_x1_sg U54390 ( .A(n37666), .B(n37667), .X(n1599) );
  nand_x1_sg U54391 ( .A(n37668), .B(n37669), .X(n1598) );
  nand_x1_sg U54392 ( .A(n37678), .B(n37679), .X(n1593) );
  nand_x1_sg U54393 ( .A(n37680), .B(n37681), .X(n1592) );
  nand_x1_sg U54394 ( .A(n37682), .B(n37683), .X(n1591) );
  nand_x1_sg U54395 ( .A(n37684), .B(n37685), .X(n1590) );
  nand_x1_sg U54396 ( .A(n37920), .B(n37921), .X(n1472) );
  nand_x1_sg U54397 ( .A(n37922), .B(n37923), .X(n1471) );
  nand_x1_sg U54398 ( .A(n37924), .B(n37925), .X(n1470) );
  nand_x1_sg U54399 ( .A(n37946), .B(n37947), .X(n1459) );
  nand_x1_sg U54400 ( .A(n37948), .B(n37949), .X(n1458) );
  nand_x1_sg U54401 ( .A(n37960), .B(n37961), .X(n1452) );
  nand_x1_sg U54402 ( .A(n37962), .B(n37963), .X(n1451) );
  nand_x1_sg U54403 ( .A(n37964), .B(n37965), .X(n1450) );
  nand_x1_sg U54404 ( .A(n37986), .B(n37987), .X(n1439) );
  nand_x1_sg U54405 ( .A(n37988), .B(n37989), .X(n1438) );
  nand_x1_sg U54406 ( .A(n37044), .B(n37045), .X(n1930) );
  nand_x1_sg U54407 ( .A(n37124), .B(n37125), .X(n1890) );
  nand_x1_sg U54408 ( .A(n37364), .B(n37365), .X(n1770) );
  nand_x1_sg U54409 ( .A(n37036), .B(n37037), .X(n1934) );
  nand_x1_sg U54410 ( .A(n37038), .B(n37039), .X(n1933) );
  nand_x1_sg U54411 ( .A(n37356), .B(n37357), .X(n1774) );
  nand_x1_sg U54412 ( .A(n37358), .B(n37359), .X(n1773) );
  nand_x1_sg U54413 ( .A(n37030), .B(n37031), .X(n1937) );
  nand_x1_sg U54414 ( .A(n37032), .B(n37033), .X(n1936) );
  nand_x1_sg U54415 ( .A(n37350), .B(n37351), .X(n1777) );
  nand_x1_sg U54416 ( .A(n37352), .B(n37353), .X(n1776) );
  nand_x1_sg U54417 ( .A(n37034), .B(n37035), .X(n1935) );
  nand_x1_sg U54418 ( .A(n37354), .B(n37355), .X(n1775) );
  nand_x1_sg U54419 ( .A(n37040), .B(n37041), .X(n1932) );
  nand_x1_sg U54420 ( .A(n37046), .B(n37047), .X(n1929) );
  nand_x1_sg U54421 ( .A(n37048), .B(n37049), .X(n1928) );
  nand_x1_sg U54422 ( .A(n37050), .B(n37051), .X(n1927) );
  nand_x1_sg U54423 ( .A(n37052), .B(n37053), .X(n1926) );
  nand_x1_sg U54424 ( .A(n37054), .B(n37055), .X(n1925) );
  nand_x1_sg U54425 ( .A(n37056), .B(n37057), .X(n1924) );
  nand_x1_sg U54426 ( .A(n37058), .B(n37059), .X(n1923) );
  nand_x1_sg U54427 ( .A(n37060), .B(n37061), .X(n1922) );
  nand_x1_sg U54428 ( .A(n37062), .B(n37063), .X(n1921) );
  nand_x1_sg U54429 ( .A(n37064), .B(n37065), .X(n1920) );
  nand_x1_sg U54430 ( .A(n37120), .B(n37121), .X(n1892) );
  nand_x1_sg U54431 ( .A(n37126), .B(n37127), .X(n1889) );
  nand_x1_sg U54432 ( .A(n37128), .B(n37129), .X(n1888) );
  nand_x1_sg U54433 ( .A(n37340), .B(n37341), .X(n1782) );
  nand_x1_sg U54434 ( .A(n37342), .B(n37343), .X(n1781) );
  nand_x1_sg U54435 ( .A(n37344), .B(n37345), .X(n1780) );
  nand_x1_sg U54436 ( .A(n37360), .B(n37361), .X(n1772) );
  nand_x1_sg U54437 ( .A(n37366), .B(n37367), .X(n1769) );
  nand_x1_sg U54438 ( .A(n37368), .B(n37369), .X(n1768) );
  nand_x1_sg U54439 ( .A(n37370), .B(n37371), .X(n1767) );
  nand_x1_sg U54440 ( .A(n37372), .B(n37373), .X(n1766) );
  nand_x1_sg U54441 ( .A(n37374), .B(n37375), .X(n1765) );
  nand_x1_sg U54442 ( .A(n37376), .B(n37377), .X(n1764) );
  nand_x1_sg U54443 ( .A(n37378), .B(n37379), .X(n1763) );
  nand_x1_sg U54444 ( .A(n37380), .B(n37381), .X(n1762) );
  nand_x1_sg U54445 ( .A(n37382), .B(n37383), .X(n1761) );
  nand_x1_sg U54446 ( .A(n37384), .B(n37385), .X(n1760) );
  nand_x1_sg U54447 ( .A(n37606), .B(n37607), .X(n1629) );
  nand_x1_sg U54448 ( .A(n37608), .B(n37609), .X(n1628) );
  nand_x1_sg U54449 ( .A(n37610), .B(n37611), .X(n1627) );
  nand_x1_sg U54450 ( .A(n37612), .B(n37613), .X(n1626) );
  nand_x1_sg U54451 ( .A(n37614), .B(n37615), .X(n1625) );
  nand_x1_sg U54452 ( .A(n37616), .B(n37617), .X(n1624) );
  nand_x1_sg U54453 ( .A(n37618), .B(n37619), .X(n1623) );
  nand_x1_sg U54454 ( .A(n37620), .B(n37621), .X(n1622) );
  nand_x1_sg U54455 ( .A(n37622), .B(n37623), .X(n1621) );
  nand_x1_sg U54456 ( .A(n37624), .B(n37625), .X(n1620) );
  nand_x1_sg U54457 ( .A(n37634), .B(n37635), .X(n1615) );
  nand_x1_sg U54458 ( .A(n37636), .B(n37637), .X(n1614) );
  nand_x1_sg U54459 ( .A(n37646), .B(n37647), .X(n1609) );
  nand_x1_sg U54460 ( .A(n37648), .B(n37649), .X(n1608) );
  nand_x1_sg U54461 ( .A(n37714), .B(n37715), .X(n1575) );
  nand_x1_sg U54462 ( .A(n37716), .B(n37717), .X(n1574) );
  nand_x1_sg U54463 ( .A(n37726), .B(n37727), .X(n1569) );
  nand_x1_sg U54464 ( .A(n37728), .B(n37729), .X(n1568) );
  nand_x1_sg U54465 ( .A(n37730), .B(n37731), .X(n1567) );
  nand_x1_sg U54466 ( .A(n37732), .B(n37733), .X(n1566) );
  nand_x1_sg U54467 ( .A(n37734), .B(n37735), .X(n1565) );
  nand_x1_sg U54468 ( .A(n37736), .B(n37737), .X(n1564) );
  nand_x1_sg U54469 ( .A(n37738), .B(n37739), .X(n1563) );
  nand_x1_sg U54470 ( .A(n37740), .B(n37741), .X(n1562) );
  nand_x1_sg U54471 ( .A(n37742), .B(n37743), .X(n1561) );
  nand_x1_sg U54472 ( .A(n37744), .B(n37745), .X(n1560) );
  nand_x1_sg U54473 ( .A(n37860), .B(n37861), .X(n1502) );
  nand_x1_sg U54474 ( .A(n37862), .B(n37863), .X(n1501) );
  nand_x1_sg U54475 ( .A(n37864), .B(n37865), .X(n1500) );
  nand_x1_sg U54476 ( .A(n37874), .B(n37875), .X(n1495) );
  nand_x1_sg U54477 ( .A(n37876), .B(n37877), .X(n1494) );
  nand_x1_sg U54478 ( .A(n37886), .B(n37887), .X(n1489) );
  nand_x1_sg U54479 ( .A(n37888), .B(n37889), .X(n1488) );
  nand_x1_sg U54480 ( .A(n37890), .B(n37891), .X(n1487) );
  nand_x1_sg U54481 ( .A(n37892), .B(n37893), .X(n1486) );
  nand_x1_sg U54482 ( .A(n37894), .B(n37895), .X(n1485) );
  nand_x1_sg U54483 ( .A(n37896), .B(n37897), .X(n1484) );
  nand_x1_sg U54484 ( .A(n37898), .B(n37899), .X(n1483) );
  nand_x1_sg U54485 ( .A(n37900), .B(n37901), .X(n1482) );
  nand_x1_sg U54486 ( .A(n37902), .B(n37903), .X(n1481) );
  nand_x1_sg U54487 ( .A(n37904), .B(n37905), .X(n1480) );
  nand_x1_sg U54488 ( .A(n37914), .B(n37915), .X(n1475) );
  nand_x1_sg U54489 ( .A(n37916), .B(n37917), .X(n1474) );
  nand_x1_sg U54490 ( .A(n37068), .B(n37069), .X(n1918) );
  nand_x1_sg U54491 ( .A(n37348), .B(n37349), .X(n1778) );
  nand_x1_sg U54492 ( .A(n37388), .B(n37389), .X(n1758) );
  nand_x1_sg U54493 ( .A(n37630), .B(n37631), .X(n1617) );
  nand_x1_sg U54494 ( .A(n37632), .B(n37633), .X(n1616) );
  nand_x1_sg U54495 ( .A(n37710), .B(n37711), .X(n1577) );
  nand_x1_sg U54496 ( .A(n37712), .B(n37713), .X(n1576) );
  nand_x1_sg U54497 ( .A(n37870), .B(n37871), .X(n1497) );
  nand_x1_sg U54498 ( .A(n37872), .B(n37873), .X(n1496) );
  nand_x1_sg U54499 ( .A(n37910), .B(n37911), .X(n1477) );
  nand_x1_sg U54500 ( .A(n37912), .B(n37913), .X(n1476) );
  nand_x1_sg U54501 ( .A(n37122), .B(n37123), .X(n1891) );
  nand_x1_sg U54502 ( .A(n37386), .B(n37387), .X(n1759) );
  nand_x1_sg U54503 ( .A(n37640), .B(n37641), .X(n1612) );
  nand_x1_sg U54504 ( .A(n37642), .B(n37643), .X(n1611) );
  nand_x1_sg U54505 ( .A(n37644), .B(n37645), .X(n1610) );
  nand_x1_sg U54506 ( .A(n37906), .B(n37907), .X(n1479) );
  nand_x1_sg U54507 ( .A(n37042), .B(n37043), .X(n1931) );
  nand_x1_sg U54508 ( .A(n37066), .B(n37067), .X(n1919) );
  nand_x1_sg U54509 ( .A(n37346), .B(n37347), .X(n1779) );
  nand_x1_sg U54510 ( .A(n37362), .B(n37363), .X(n1771) );
  nand_x1_sg U54511 ( .A(n37600), .B(n37601), .X(n1632) );
  nand_x1_sg U54512 ( .A(n37602), .B(n37603), .X(n1631) );
  nand_x1_sg U54513 ( .A(n37604), .B(n37605), .X(n1630) );
  nand_x1_sg U54514 ( .A(n37626), .B(n37627), .X(n1619) );
  nand_x1_sg U54515 ( .A(n37628), .B(n37629), .X(n1618) );
  nand_x1_sg U54516 ( .A(n37638), .B(n37639), .X(n1613) );
  nand_x1_sg U54517 ( .A(n37718), .B(n37719), .X(n1573) );
  nand_x1_sg U54518 ( .A(n37720), .B(n37721), .X(n1572) );
  nand_x1_sg U54519 ( .A(n37722), .B(n37723), .X(n1571) );
  nand_x1_sg U54520 ( .A(n37724), .B(n37725), .X(n1570) );
  nand_x1_sg U54521 ( .A(n37746), .B(n37747), .X(n1559) );
  nand_x1_sg U54522 ( .A(n37748), .B(n37749), .X(n1558) );
  nand_x1_sg U54523 ( .A(n37866), .B(n37867), .X(n1499) );
  nand_x1_sg U54524 ( .A(n37868), .B(n37869), .X(n1498) );
  nand_x1_sg U54525 ( .A(n37878), .B(n37879), .X(n1493) );
  nand_x1_sg U54526 ( .A(n37880), .B(n37881), .X(n1492) );
  nand_x1_sg U54527 ( .A(n37882), .B(n37883), .X(n1491) );
  nand_x1_sg U54528 ( .A(n37884), .B(n37885), .X(n1490) );
  nand_x1_sg U54529 ( .A(n37908), .B(n37909), .X(n1478) );
  nand_x1_sg U54530 ( .A(n37918), .B(n37919), .X(n1473) );
  nand_x1_sg U54531 ( .A(n36874), .B(n36875), .X(out[3]) );
  nand_x1_sg U54532 ( .A(n36872), .B(n36873), .X(out[4]) );
  nand_x1_sg U54533 ( .A(n36870), .B(n36871), .X(out[5]) );
  nand_x1_sg U54534 ( .A(n36868), .B(n36869), .X(out[6]) );
  nand_x1_sg U54535 ( .A(n36866), .B(n36867), .X(out[7]) );
  nand_x1_sg U54536 ( .A(n36864), .B(n36865), .X(out[8]) );
  nand_x1_sg U54537 ( .A(n36862), .B(n36863), .X(out[9]) );
  nand_x1_sg U54538 ( .A(n36900), .B(n36901), .X(out[0]) );
  nand_x1_sg U54539 ( .A(n36876), .B(n36877), .X(out[2]) );
  nand_x1_sg U54540 ( .A(n36898), .B(n36899), .X(out[10]) );
  nand_x1_sg U54541 ( .A(n36896), .B(n36897), .X(out[11]) );
  nand_x1_sg U54542 ( .A(n36894), .B(n36895), .X(out[12]) );
  nand_x1_sg U54543 ( .A(n36892), .B(n36893), .X(out[13]) );
  nand_x1_sg U54544 ( .A(n36890), .B(n36891), .X(out[14]) );
  nand_x1_sg U54545 ( .A(n36888), .B(n36889), .X(out[15]) );
  nand_x1_sg U54546 ( .A(n36884), .B(n36885), .X(out[17]) );
  nand_x1_sg U54547 ( .A(n36882), .B(n36883), .X(out[18]) );
  nand_x1_sg U54548 ( .A(n36880), .B(n36881), .X(out[19]) );
  nand_x2_sg U54549 ( .A(n6757), .B(n6804), .X(n6803) );
  inv_x1_sg U54550 ( .A(n26173), .X(n50278) );
  inv_x1_sg U54551 ( .A(n20449), .X(n46377) );
  inv_x1_sg U54552 ( .A(n20596), .X(n46553) );
  inv_x1_sg U54553 ( .A(n20140), .X(n46471) );
  inv_x1_sg U54554 ( .A(n20307), .X(n46425) );
  inv_x1_sg U54555 ( .A(n21355), .X(n46463) );
  inv_x1_sg U54556 ( .A(n28919), .X(n45608) );
  inv_x1_sg U54557 ( .A(n23000), .X(n47405) );
  inv_x1_sg U54558 ( .A(n23280), .X(n47690) );
  inv_x1_sg U54559 ( .A(n23559), .X(n47975) );
  inv_x1_sg U54560 ( .A(n23838), .X(n48260) );
  inv_x1_sg U54561 ( .A(n24117), .X(n48545) );
  inv_x1_sg U54562 ( .A(n24396), .X(n48830) );
  inv_x1_sg U54563 ( .A(n24674), .X(n49117) );
  inv_x1_sg U54564 ( .A(n24953), .X(n49403) );
  inv_x1_sg U54565 ( .A(n25232), .X(n49689) );
  inv_x1_sg U54566 ( .A(n25511), .X(n49975) );
  inv_x1_sg U54567 ( .A(n25788), .X(n50261) );
  inv_x1_sg U54568 ( .A(n26348), .X(n50835) );
  inv_x1_sg U54569 ( .A(n26626), .X(n51122) );
  inv_x1_sg U54570 ( .A(n21678), .X(n46368) );
  inv_x1_sg U54571 ( .A(n29241), .X(n45339) );
  inv_x1_sg U54572 ( .A(n29235), .X(n45430) );
  inv_x1_sg U54573 ( .A(n29229), .X(n45519) );
  inv_x1_sg U54574 ( .A(n23100), .X(n47142) );
  inv_x1_sg U54575 ( .A(n23380), .X(n47427) );
  inv_x1_sg U54576 ( .A(n23659), .X(n47712) );
  inv_x1_sg U54577 ( .A(n23938), .X(n47997) );
  inv_x1_sg U54578 ( .A(n24217), .X(n48282) );
  inv_x1_sg U54579 ( .A(n24496), .X(n48567) );
  inv_x1_sg U54580 ( .A(n24774), .X(n48852) );
  inv_x1_sg U54581 ( .A(n25053), .X(n49139) );
  inv_x1_sg U54582 ( .A(n25332), .X(n49425) );
  inv_x1_sg U54583 ( .A(n25611), .X(n49711) );
  inv_x1_sg U54584 ( .A(n25888), .X(n49997) );
  inv_x1_sg U54585 ( .A(n26448), .X(n50572) );
  inv_x1_sg U54586 ( .A(n26726), .X(n50858) );
  inv_x1_sg U54587 ( .A(n20593), .X(n46613) );
  inv_x1_sg U54588 ( .A(n20791), .X(n46577) );
  inv_x1_sg U54589 ( .A(n28367), .X(n44967) );
  inv_x1_sg U54590 ( .A(n27412), .X(n44972) );
  inv_x1_sg U54591 ( .A(n28622), .X(n44965) );
  inv_x1_sg U54592 ( .A(n27801), .X(n44970) );
  inv_x1_sg U54593 ( .A(n23122), .X(n47139) );
  inv_x1_sg U54594 ( .A(n23402), .X(n47424) );
  inv_x1_sg U54595 ( .A(n23681), .X(n47709) );
  inv_x1_sg U54596 ( .A(n23960), .X(n47994) );
  inv_x1_sg U54597 ( .A(n24239), .X(n48279) );
  inv_x1_sg U54598 ( .A(n24518), .X(n48564) );
  inv_x1_sg U54599 ( .A(n24796), .X(n48849) );
  inv_x1_sg U54600 ( .A(n25075), .X(n49136) );
  inv_x1_sg U54601 ( .A(n25354), .X(n49422) );
  inv_x1_sg U54602 ( .A(n25633), .X(n49708) );
  inv_x1_sg U54603 ( .A(n25910), .X(n49994) );
  inv_x1_sg U54604 ( .A(n26470), .X(n50569) );
  inv_x1_sg U54605 ( .A(n26748), .X(n50855) );
  inv_x1_sg U54606 ( .A(n22845), .X(n46847) );
  inv_x1_sg U54607 ( .A(n28542), .X(n45782) );
  inv_x1_sg U54608 ( .A(n20984), .X(n46617) );
  inv_x1_sg U54609 ( .A(n19585), .X(n46390) );
  inv_x1_sg U54610 ( .A(n26951), .X(n44974) );
  inv_x1_sg U54611 ( .A(n21343), .X(n46498) );
  inv_x1_sg U54612 ( .A(n21337), .X(n46460) );
  inv_x1_sg U54613 ( .A(n21332), .X(n46412) );
  inv_x1_sg U54614 ( .A(n21327), .X(n46365) );
  inv_x1_sg U54615 ( .A(n20553), .X(n46314) );
  inv_x1_sg U54616 ( .A(n21322), .X(n46323) );
  inv_x1_sg U54617 ( .A(n21317), .X(n46278) );
  inv_x1_sg U54618 ( .A(n20548), .X(n46269) );
  inv_x1_sg U54619 ( .A(n21312), .X(n46232) );
  inv_x1_sg U54620 ( .A(n21307), .X(n46187) );
  inv_x1_sg U54621 ( .A(n20543), .X(n46223) );
  inv_x1_sg U54622 ( .A(n21302), .X(n46141) );
  inv_x1_sg U54623 ( .A(n20538), .X(n46178) );
  inv_x1_sg U54624 ( .A(n21297), .X(n46096) );
  inv_x1_sg U54625 ( .A(n20533), .X(n46132) );
  inv_x1_sg U54626 ( .A(n21292), .X(n46050) );
  inv_x1_sg U54627 ( .A(n20528), .X(n46087) );
  inv_x1_sg U54628 ( .A(n21287), .X(n46005) );
  inv_x1_sg U54629 ( .A(n20523), .X(n46041) );
  inv_x1_sg U54630 ( .A(n21282), .X(n45960) );
  inv_x1_sg U54631 ( .A(n20518), .X(n45996) );
  inv_x1_sg U54632 ( .A(n20513), .X(n45951) );
  inv_x1_sg U54633 ( .A(n21086), .X(n45912) );
  inv_x1_sg U54634 ( .A(n19749), .X(n46554) );
  inv_x1_sg U54635 ( .A(n20305), .X(n46426) );
  inv_x1_sg U54636 ( .A(n21366), .X(n46540) );
  inv_x1_sg U54637 ( .A(n20558), .X(n46356) );
  inv_x1_sg U54638 ( .A(n20377), .X(n45902) );
  inv_x1_sg U54639 ( .A(n19896), .X(n46305) );
  inv_x1_sg U54640 ( .A(n19644), .X(n45892) );
  inv_x1_sg U54641 ( .A(n19856), .X(n45942) );
  inv_x1_sg U54642 ( .A(n19891), .X(n46260) );
  inv_x1_sg U54643 ( .A(n19886), .X(n46214) );
  inv_x1_sg U54644 ( .A(n19881), .X(n46169) );
  inv_x1_sg U54645 ( .A(n19876), .X(n46123) );
  inv_x1_sg U54646 ( .A(n19871), .X(n46078) );
  inv_x1_sg U54647 ( .A(n19866), .X(n46032) );
  inv_x1_sg U54648 ( .A(n19861), .X(n45987) );
  inv_x1_sg U54649 ( .A(n19481), .X(n46344) );
  inv_x1_sg U54650 ( .A(n28136), .X(n44997) );
  inv_x1_sg U54651 ( .A(n6716), .X(n45866) );
  inv_x1_sg U54652 ( .A(n6268), .X(n46296) );
  inv_x1_sg U54653 ( .A(n6313), .X(n46251) );
  inv_x1_sg U54654 ( .A(n6357), .X(n46205) );
  inv_x1_sg U54655 ( .A(n6402), .X(n46160) );
  inv_x1_sg U54656 ( .A(n6446), .X(n46114) );
  inv_x1_sg U54657 ( .A(n6491), .X(n46069) );
  inv_x1_sg U54658 ( .A(n6535), .X(n46023) );
  inv_x1_sg U54659 ( .A(n6580), .X(n45978) );
  inv_x1_sg U54660 ( .A(n6624), .X(n45933) );
  inv_x1_sg U54661 ( .A(n21271), .X(n45818) );
  inv_x1_sg U54662 ( .A(n20502), .X(n45834) );
  inv_x1_sg U54663 ( .A(n20303), .X(n46451) );
  inv_x1_sg U54664 ( .A(n19845), .X(n45850) );
  inv_x1_sg U54665 ( .A(n20445), .X(n46403) );
  inv_x1_sg U54666 ( .A(n20860), .X(n45909) );
  inv_x1_sg U54667 ( .A(n20447), .X(n46378) );
  inv_x1_sg U54668 ( .A(n19709), .X(n46394) );
  inv_x1_sg U54669 ( .A(n20217), .X(n45899) );
  inv_x1_sg U54670 ( .A(n19411), .X(n45889) );
  inv_x1_sg U54671 ( .A(n28147), .X(n45104) );
  inv_x1_sg U54672 ( .A(n28152), .X(n45150) );
  inv_x1_sg U54673 ( .A(n28157), .X(n45195) );
  inv_x1_sg U54674 ( .A(n28162), .X(n45241) );
  inv_x1_sg U54675 ( .A(n28167), .X(n45286) );
  inv_x1_sg U54676 ( .A(n28172), .X(n45331) );
  inv_x1_sg U54677 ( .A(n28177), .X(n45376) );
  inv_x1_sg U54678 ( .A(n28183), .X(n45422) );
  inv_x1_sg U54679 ( .A(n28212), .X(n45466) );
  inv_x1_sg U54680 ( .A(n28077), .X(n45490) );
  inv_x1_sg U54681 ( .A(n27915), .X(n45534) );
  inv_x1_sg U54682 ( .A(n27738), .X(n45579) );
  inv_x1_sg U54683 ( .A(n27544), .X(n45623) );
  inv_x1_sg U54684 ( .A(n27331), .X(n45667) );
  inv_x1_sg U54685 ( .A(n19715), .X(n46443) );
  inv_x1_sg U54686 ( .A(n26122), .X(n50280) );
  inv_x1_sg U54687 ( .A(n21672), .X(n46416) );
  inv_x1_sg U54688 ( .A(n20109), .X(n46350) );
  inv_x1_sg U54689 ( .A(n19939), .X(n46533) );
  inv_x1_sg U54690 ( .A(n26846), .X(n45754) );
  inv_x1_sg U54691 ( .A(n21540), .X(n46501) );
  inv_x1_sg U54692 ( .A(n19321), .X(n46482) );
  inv_x1_sg U54693 ( .A(n20138), .X(n46472) );
  inv_x1_sg U54694 ( .A(n29199), .X(n45385) );
  inv_x1_sg U54695 ( .A(n29211), .X(n45475) );
  inv_x1_sg U54696 ( .A(n29223), .X(n45564) );
  inv_x1_sg U54697 ( .A(n29091), .X(n45652) );
  inv_x1_sg U54698 ( .A(n19327), .X(n46527) );
  inv_x1_sg U54699 ( .A(n19142), .X(n46607) );
  inv_x1_sg U54700 ( .A(n19567), .X(n46612) );
  inv_x1_sg U54701 ( .A(n19560), .X(n46603) );
  inv_x1_sg U54702 ( .A(n19553), .X(n46601) );
  inv_x1_sg U54703 ( .A(n19546), .X(n46599) );
  inv_x1_sg U54704 ( .A(n20585), .X(n46593) );
  inv_x1_sg U54705 ( .A(n20591), .X(n46614) );
  inv_x1_sg U54706 ( .A(n19532), .X(n46595) );
  inv_x1_sg U54707 ( .A(n21002), .X(n46589) );
  inv_x1_sg U54708 ( .A(n19539), .X(n46597) );
  inv_x1_sg U54709 ( .A(n20994), .X(n46587) );
  inv_x1_sg U54710 ( .A(n21009), .X(n46615) );
  inv_x1_sg U54711 ( .A(n19149), .X(n46610) );
  inv_x1_sg U54712 ( .A(n6035), .X(n46524) );
  inv_x1_sg U54713 ( .A(n6176), .X(n46387) );
  nand_x2_sg U54714 ( .A(n21588), .B(n21589), .X(n21430) );
  nand_x2_sg U54715 ( .A(n29139), .B(n29140), .X(n28981) );
  nor_x1_sg U54716 ( .A(n22570), .B(n22571), .X(n22559) );
  nor_x1_sg U54717 ( .A(n19943), .B(n5553), .X(n19942) );
  nor_x1_sg U54718 ( .A(n28249), .B(n5282), .X(n28248) );
  nor_x1_sg U54719 ( .A(n20653), .B(n5586), .X(n20652) );
  nor_x1_sg U54720 ( .A(n20013), .B(n5510), .X(n20012) );
  nor_x1_sg U54721 ( .A(n19209), .B(n5434), .X(n19208) );
  nor_x1_sg U54722 ( .A(n21423), .B(n5662), .X(n21422) );
  nand_x4_sg U54723 ( .A(n29267), .B(out_L1[0]), .X(n29266) );
  nand_x4_sg U54724 ( .A(n21716), .B(out_L2[0]), .X(n21715) );
  inv_x1_sg U54725 ( .A(n7040), .X(n47117) );
  inv_x1_sg U54726 ( .A(n7858), .X(n47403) );
  inv_x1_sg U54727 ( .A(n8676), .X(n47688) );
  inv_x1_sg U54728 ( .A(n9496), .X(n47973) );
  inv_x1_sg U54729 ( .A(n10315), .X(n48258) );
  inv_x1_sg U54730 ( .A(n11134), .X(n48543) );
  inv_x1_sg U54731 ( .A(n11953), .X(n48828) );
  inv_x1_sg U54732 ( .A(n12772), .X(n49115) );
  inv_x1_sg U54733 ( .A(n13591), .X(n49401) );
  inv_x1_sg U54734 ( .A(n14410), .X(n49687) );
  inv_x1_sg U54735 ( .A(n15229), .X(n49973) );
  inv_x1_sg U54736 ( .A(n16048), .X(n50259) );
  inv_x1_sg U54737 ( .A(n16867), .X(n50544) );
  inv_x1_sg U54738 ( .A(n17686), .X(n50833) );
  inv_x1_sg U54739 ( .A(n18507), .X(n51120) );
  nor_x1_sg U54740 ( .A(n47071), .B(n6911), .X(n6909) );
  nor_x1_sg U54741 ( .A(n6912), .B(n6913), .X(n6911) );
  nand_x1_sg U54742 ( .A(n6913), .B(n6912), .X(n6914) );
  nor_x1_sg U54743 ( .A(n47093), .B(n6917), .X(n6915) );
  nor_x1_sg U54744 ( .A(n6918), .B(n6919), .X(n6917) );
  nand_x1_sg U54745 ( .A(n6919), .B(n6918), .X(n6920) );
  nor_x1_sg U54746 ( .A(n47118), .B(n6923), .X(n6921) );
  nor_x1_sg U54747 ( .A(n6924), .B(n6925), .X(n6923) );
  nand_x1_sg U54748 ( .A(n6925), .B(n6924), .X(n6926) );
  nor_x1_sg U54749 ( .A(n47379), .B(n7734), .X(n7732) );
  nor_x1_sg U54750 ( .A(n7735), .B(n7736), .X(n7734) );
  nand_x1_sg U54751 ( .A(n7736), .B(n7735), .X(n7737) );
  nor_x1_sg U54752 ( .A(n47404), .B(n7740), .X(n7738) );
  nor_x1_sg U54753 ( .A(n7741), .B(n7742), .X(n7740) );
  nand_x1_sg U54754 ( .A(n7742), .B(n7741), .X(n7743) );
  nor_x1_sg U54755 ( .A(n47664), .B(n8552), .X(n8550) );
  nor_x1_sg U54756 ( .A(n8553), .B(n8554), .X(n8552) );
  nand_x1_sg U54757 ( .A(n8554), .B(n8553), .X(n8555) );
  nor_x1_sg U54758 ( .A(n47689), .B(n8558), .X(n8556) );
  nor_x1_sg U54759 ( .A(n8559), .B(n8560), .X(n8558) );
  nand_x1_sg U54760 ( .A(n8560), .B(n8559), .X(n8561) );
  nor_x1_sg U54761 ( .A(n47949), .B(n9372), .X(n9370) );
  nor_x1_sg U54762 ( .A(n9373), .B(n9374), .X(n9372) );
  nand_x1_sg U54763 ( .A(n9374), .B(n9373), .X(n9375) );
  nor_x1_sg U54764 ( .A(n47974), .B(n9378), .X(n9376) );
  nor_x1_sg U54765 ( .A(n9379), .B(n9380), .X(n9378) );
  nand_x1_sg U54766 ( .A(n9380), .B(n9379), .X(n9381) );
  nor_x1_sg U54767 ( .A(n48234), .B(n10191), .X(n10189) );
  nor_x1_sg U54768 ( .A(n10192), .B(n10193), .X(n10191) );
  nand_x1_sg U54769 ( .A(n10193), .B(n10192), .X(n10194) );
  nor_x1_sg U54770 ( .A(n48259), .B(n10197), .X(n10195) );
  nor_x1_sg U54771 ( .A(n10198), .B(n10199), .X(n10197) );
  nand_x1_sg U54772 ( .A(n10199), .B(n10198), .X(n10200) );
  nor_x1_sg U54773 ( .A(n48519), .B(n11010), .X(n11008) );
  nor_x1_sg U54774 ( .A(n11011), .B(n11012), .X(n11010) );
  nand_x1_sg U54775 ( .A(n11012), .B(n11011), .X(n11013) );
  nor_x1_sg U54776 ( .A(n48544), .B(n11016), .X(n11014) );
  nor_x1_sg U54777 ( .A(n11017), .B(n11018), .X(n11016) );
  nand_x1_sg U54778 ( .A(n11018), .B(n11017), .X(n11019) );
  nor_x1_sg U54779 ( .A(n48804), .B(n11829), .X(n11827) );
  nor_x1_sg U54780 ( .A(n11830), .B(n11831), .X(n11829) );
  nand_x1_sg U54781 ( .A(n11831), .B(n11830), .X(n11832) );
  nor_x1_sg U54782 ( .A(n48829), .B(n11835), .X(n11833) );
  nor_x1_sg U54783 ( .A(n11836), .B(n11837), .X(n11835) );
  nand_x1_sg U54784 ( .A(n11837), .B(n11836), .X(n11838) );
  nor_x1_sg U54785 ( .A(n49091), .B(n12648), .X(n12646) );
  nor_x1_sg U54786 ( .A(n12649), .B(n12650), .X(n12648) );
  nand_x1_sg U54787 ( .A(n12650), .B(n12649), .X(n12651) );
  nor_x1_sg U54788 ( .A(n49116), .B(n12654), .X(n12652) );
  nor_x1_sg U54789 ( .A(n12655), .B(n12656), .X(n12654) );
  nand_x1_sg U54790 ( .A(n12656), .B(n12655), .X(n12657) );
  nor_x1_sg U54791 ( .A(n49377), .B(n13467), .X(n13465) );
  nor_x1_sg U54792 ( .A(n13468), .B(n13469), .X(n13467) );
  nand_x1_sg U54793 ( .A(n13469), .B(n13468), .X(n13470) );
  nor_x1_sg U54794 ( .A(n49402), .B(n13473), .X(n13471) );
  nor_x1_sg U54795 ( .A(n13474), .B(n13475), .X(n13473) );
  nand_x1_sg U54796 ( .A(n13475), .B(n13474), .X(n13476) );
  nor_x1_sg U54797 ( .A(n49663), .B(n14286), .X(n14284) );
  nor_x1_sg U54798 ( .A(n14287), .B(n14288), .X(n14286) );
  nand_x1_sg U54799 ( .A(n14288), .B(n14287), .X(n14289) );
  nor_x1_sg U54800 ( .A(n49688), .B(n14292), .X(n14290) );
  nor_x1_sg U54801 ( .A(n14293), .B(n14294), .X(n14292) );
  nand_x1_sg U54802 ( .A(n14294), .B(n14293), .X(n14295) );
  nor_x1_sg U54803 ( .A(n49949), .B(n15105), .X(n15103) );
  nor_x1_sg U54804 ( .A(n15106), .B(n15107), .X(n15105) );
  nand_x1_sg U54805 ( .A(n15107), .B(n15106), .X(n15108) );
  nor_x1_sg U54806 ( .A(n49974), .B(n15111), .X(n15109) );
  nor_x1_sg U54807 ( .A(n15112), .B(n15113), .X(n15111) );
  nand_x1_sg U54808 ( .A(n15113), .B(n15112), .X(n15114) );
  nor_x1_sg U54809 ( .A(n50235), .B(n15924), .X(n15922) );
  nor_x1_sg U54810 ( .A(n15925), .B(n15926), .X(n15924) );
  nand_x1_sg U54811 ( .A(n15926), .B(n15925), .X(n15927) );
  nor_x1_sg U54812 ( .A(n50260), .B(n15930), .X(n15928) );
  nor_x1_sg U54813 ( .A(n15931), .B(n15932), .X(n15930) );
  nand_x1_sg U54814 ( .A(n15932), .B(n15931), .X(n15933) );
  nor_x1_sg U54815 ( .A(n50498), .B(n16735), .X(n16733) );
  nor_x1_sg U54816 ( .A(n16736), .B(n16737), .X(n16735) );
  nand_x1_sg U54817 ( .A(n16737), .B(n16736), .X(n16738) );
  nor_x1_sg U54818 ( .A(n50520), .B(n16741), .X(n16739) );
  nor_x1_sg U54819 ( .A(n16742), .B(n16743), .X(n16741) );
  nand_x1_sg U54820 ( .A(n16743), .B(n16742), .X(n16744) );
  nor_x1_sg U54821 ( .A(n50545), .B(n16747), .X(n16745) );
  nor_x1_sg U54822 ( .A(n16748), .B(n16749), .X(n16747) );
  nand_x1_sg U54823 ( .A(n16749), .B(n16748), .X(n16750) );
  nor_x1_sg U54824 ( .A(n50809), .B(n17562), .X(n17560) );
  nor_x1_sg U54825 ( .A(n17563), .B(n17564), .X(n17562) );
  nand_x1_sg U54826 ( .A(n17564), .B(n17563), .X(n17565) );
  nor_x1_sg U54827 ( .A(n50834), .B(n17568), .X(n17566) );
  nor_x1_sg U54828 ( .A(n17569), .B(n17570), .X(n17568) );
  nand_x1_sg U54829 ( .A(n17570), .B(n17569), .X(n17571) );
  nor_x1_sg U54830 ( .A(n51096), .B(n18383), .X(n18381) );
  nor_x1_sg U54831 ( .A(n18384), .B(n18385), .X(n18383) );
  nand_x1_sg U54832 ( .A(n18385), .B(n18384), .X(n18386) );
  nor_x1_sg U54833 ( .A(n51121), .B(n18389), .X(n18387) );
  nor_x1_sg U54834 ( .A(n18390), .B(n18391), .X(n18389) );
  nand_x1_sg U54835 ( .A(n18391), .B(n18390), .X(n18392) );
  inv_x1_sg U54836 ( .A(n6919), .X(n47092) );
  inv_x1_sg U54837 ( .A(n7736), .X(n47378) );
  inv_x1_sg U54838 ( .A(n8554), .X(n47663) );
  inv_x1_sg U54839 ( .A(n9374), .X(n47948) );
  inv_x1_sg U54840 ( .A(n10193), .X(n48233) );
  inv_x1_sg U54841 ( .A(n11012), .X(n48518) );
  inv_x1_sg U54842 ( .A(n11831), .X(n48803) );
  inv_x1_sg U54843 ( .A(n12650), .X(n49090) );
  inv_x1_sg U54844 ( .A(n13469), .X(n49376) );
  inv_x1_sg U54845 ( .A(n14288), .X(n49662) );
  inv_x1_sg U54846 ( .A(n15107), .X(n49948) );
  inv_x1_sg U54847 ( .A(n15926), .X(n50234) );
  inv_x1_sg U54848 ( .A(n16743), .X(n50519) );
  inv_x1_sg U54849 ( .A(n17564), .X(n50808) );
  inv_x1_sg U54850 ( .A(n18385), .X(n51095) );
  inv_x1_sg U54851 ( .A(n6913), .X(n47070) );
  inv_x1_sg U54852 ( .A(n16737), .X(n50497) );
  inv_x1_sg U54853 ( .A(n6925), .X(n47116) );
  inv_x1_sg U54854 ( .A(n7742), .X(n47402) );
  inv_x1_sg U54855 ( .A(n8560), .X(n47687) );
  inv_x1_sg U54856 ( .A(n9380), .X(n47972) );
  inv_x1_sg U54857 ( .A(n10199), .X(n48257) );
  inv_x1_sg U54858 ( .A(n11018), .X(n48542) );
  inv_x1_sg U54859 ( .A(n11837), .X(n48827) );
  inv_x1_sg U54860 ( .A(n12656), .X(n49114) );
  inv_x1_sg U54861 ( .A(n13475), .X(n49400) );
  inv_x1_sg U54862 ( .A(n14294), .X(n49686) );
  inv_x1_sg U54863 ( .A(n15113), .X(n49972) );
  inv_x1_sg U54864 ( .A(n15932), .X(n50258) );
  inv_x1_sg U54865 ( .A(n16749), .X(n50543) );
  inv_x1_sg U54866 ( .A(n17570), .X(n50832) );
  inv_x1_sg U54867 ( .A(n18391), .X(n51119) );
  nor_x1_sg U54868 ( .A(n6929), .B(n47126), .X(n6927) );
  nor_x1_sg U54869 ( .A(n6932), .B(n6931), .X(n6929) );
  nand_x1_sg U54870 ( .A(n6931), .B(n6932), .X(n6930) );
  nor_x1_sg U54871 ( .A(n7746), .B(n47412), .X(n7744) );
  nor_x1_sg U54872 ( .A(n7749), .B(n7748), .X(n7746) );
  nand_x1_sg U54873 ( .A(n7748), .B(n7749), .X(n7747) );
  nor_x1_sg U54874 ( .A(n8564), .B(n47697), .X(n8562) );
  nor_x1_sg U54875 ( .A(n8567), .B(n8566), .X(n8564) );
  nand_x1_sg U54876 ( .A(n8566), .B(n8567), .X(n8565) );
  nor_x1_sg U54877 ( .A(n9384), .B(n47982), .X(n9382) );
  nor_x1_sg U54878 ( .A(n9387), .B(n9386), .X(n9384) );
  nand_x1_sg U54879 ( .A(n9386), .B(n9387), .X(n9385) );
  nor_x1_sg U54880 ( .A(n10203), .B(n48267), .X(n10201) );
  nor_x1_sg U54881 ( .A(n10206), .B(n10205), .X(n10203) );
  nand_x1_sg U54882 ( .A(n10205), .B(n10206), .X(n10204) );
  nor_x1_sg U54883 ( .A(n11022), .B(n48552), .X(n11020) );
  nor_x1_sg U54884 ( .A(n11025), .B(n11024), .X(n11022) );
  nand_x1_sg U54885 ( .A(n11024), .B(n11025), .X(n11023) );
  nor_x1_sg U54886 ( .A(n11841), .B(n48837), .X(n11839) );
  nor_x1_sg U54887 ( .A(n11844), .B(n11843), .X(n11841) );
  nand_x1_sg U54888 ( .A(n11843), .B(n11844), .X(n11842) );
  nor_x1_sg U54889 ( .A(n12660), .B(n49124), .X(n12658) );
  nor_x1_sg U54890 ( .A(n12663), .B(n12662), .X(n12660) );
  nand_x1_sg U54891 ( .A(n12662), .B(n12663), .X(n12661) );
  nor_x1_sg U54892 ( .A(n13479), .B(n49410), .X(n13477) );
  nor_x1_sg U54893 ( .A(n13482), .B(n13481), .X(n13479) );
  nand_x1_sg U54894 ( .A(n13481), .B(n13482), .X(n13480) );
  nor_x1_sg U54895 ( .A(n14298), .B(n49696), .X(n14296) );
  nor_x1_sg U54896 ( .A(n14301), .B(n14300), .X(n14298) );
  nand_x1_sg U54897 ( .A(n14300), .B(n14301), .X(n14299) );
  nor_x1_sg U54898 ( .A(n15117), .B(n49982), .X(n15115) );
  nor_x1_sg U54899 ( .A(n15120), .B(n15119), .X(n15117) );
  nand_x1_sg U54900 ( .A(n15119), .B(n15120), .X(n15118) );
  nor_x1_sg U54901 ( .A(n15936), .B(n50268), .X(n15934) );
  nor_x1_sg U54902 ( .A(n15939), .B(n15938), .X(n15936) );
  nand_x1_sg U54903 ( .A(n15938), .B(n15939), .X(n15937) );
  nor_x1_sg U54904 ( .A(n16753), .B(n50554), .X(n16751) );
  nor_x1_sg U54905 ( .A(n16756), .B(n16755), .X(n16753) );
  nand_x1_sg U54906 ( .A(n16755), .B(n16756), .X(n16754) );
  nor_x1_sg U54907 ( .A(n17574), .B(n50842), .X(n17572) );
  nor_x1_sg U54908 ( .A(n17577), .B(n17576), .X(n17574) );
  nand_x1_sg U54909 ( .A(n17576), .B(n17577), .X(n17575) );
  nor_x1_sg U54910 ( .A(n18395), .B(n51129), .X(n18393) );
  nor_x1_sg U54911 ( .A(n18398), .B(n18397), .X(n18395) );
  nand_x1_sg U54912 ( .A(n18397), .B(n18398), .X(n18396) );
  nor_x1_sg U54913 ( .A(n7040), .B(n47113), .X(n7037) );
  nor_x1_sg U54914 ( .A(n7039), .B(n47117), .X(n7038) );
  inv_x1_sg U54915 ( .A(n7039), .X(n47113) );
  nor_x1_sg U54916 ( .A(n7858), .B(n47399), .X(n7855) );
  nor_x1_sg U54917 ( .A(n7857), .B(n47403), .X(n7856) );
  inv_x1_sg U54918 ( .A(n7857), .X(n47399) );
  nor_x1_sg U54919 ( .A(n8676), .B(n47684), .X(n8673) );
  nor_x1_sg U54920 ( .A(n8675), .B(n47688), .X(n8674) );
  inv_x1_sg U54921 ( .A(n8675), .X(n47684) );
  nor_x1_sg U54922 ( .A(n9496), .B(n47969), .X(n9493) );
  nor_x1_sg U54923 ( .A(n9495), .B(n47973), .X(n9494) );
  inv_x1_sg U54924 ( .A(n9495), .X(n47969) );
  nor_x1_sg U54925 ( .A(n10315), .B(n48254), .X(n10312) );
  nor_x1_sg U54926 ( .A(n10314), .B(n48258), .X(n10313) );
  inv_x1_sg U54927 ( .A(n10314), .X(n48254) );
  nor_x1_sg U54928 ( .A(n11134), .B(n48539), .X(n11131) );
  nor_x1_sg U54929 ( .A(n11133), .B(n48543), .X(n11132) );
  inv_x1_sg U54930 ( .A(n11133), .X(n48539) );
  nor_x1_sg U54931 ( .A(n11953), .B(n48824), .X(n11950) );
  nor_x1_sg U54932 ( .A(n11952), .B(n48828), .X(n11951) );
  inv_x1_sg U54933 ( .A(n11952), .X(n48824) );
  nor_x1_sg U54934 ( .A(n12772), .B(n49111), .X(n12769) );
  nor_x1_sg U54935 ( .A(n12771), .B(n49115), .X(n12770) );
  inv_x1_sg U54936 ( .A(n12771), .X(n49111) );
  nor_x1_sg U54937 ( .A(n13591), .B(n49397), .X(n13588) );
  nor_x1_sg U54938 ( .A(n13590), .B(n49401), .X(n13589) );
  inv_x1_sg U54939 ( .A(n13590), .X(n49397) );
  nor_x1_sg U54940 ( .A(n14410), .B(n49683), .X(n14407) );
  nor_x1_sg U54941 ( .A(n14409), .B(n49687), .X(n14408) );
  inv_x1_sg U54942 ( .A(n14409), .X(n49683) );
  nor_x1_sg U54943 ( .A(n15229), .B(n49969), .X(n15226) );
  nor_x1_sg U54944 ( .A(n15228), .B(n49973), .X(n15227) );
  inv_x1_sg U54945 ( .A(n15228), .X(n49969) );
  nor_x1_sg U54946 ( .A(n16048), .B(n50255), .X(n16045) );
  nor_x1_sg U54947 ( .A(n16047), .B(n50259), .X(n16046) );
  inv_x1_sg U54948 ( .A(n16047), .X(n50255) );
  nor_x1_sg U54949 ( .A(n16867), .B(n50540), .X(n16864) );
  nor_x1_sg U54950 ( .A(n16866), .B(n50544), .X(n16865) );
  inv_x1_sg U54951 ( .A(n16866), .X(n50540) );
  nor_x1_sg U54952 ( .A(n17686), .B(n50829), .X(n17683) );
  nor_x1_sg U54953 ( .A(n17685), .B(n50833), .X(n17684) );
  inv_x1_sg U54954 ( .A(n17685), .X(n50829) );
  nor_x1_sg U54955 ( .A(n18507), .B(n51116), .X(n18504) );
  nor_x1_sg U54956 ( .A(n18506), .B(n51120), .X(n18505) );
  inv_x1_sg U54957 ( .A(n18506), .X(n51116) );
  nor_x1_sg U54958 ( .A(n47017), .B(n6899), .X(n6897) );
  nor_x1_sg U54959 ( .A(n6900), .B(n6901), .X(n6899) );
  nand_x1_sg U54960 ( .A(n6901), .B(n6900), .X(n6902) );
  nor_x1_sg U54961 ( .A(n47043), .B(n6905), .X(n6903) );
  nor_x1_sg U54962 ( .A(n6906), .B(n6907), .X(n6905) );
  nand_x1_sg U54963 ( .A(n6907), .B(n6906), .X(n6908) );
  nor_x1_sg U54964 ( .A(n47357), .B(n7728), .X(n7726) );
  nor_x1_sg U54965 ( .A(n7729), .B(n7730), .X(n7728) );
  nand_x1_sg U54966 ( .A(n7730), .B(n7729), .X(n7731) );
  nor_x1_sg U54967 ( .A(n47642), .B(n8546), .X(n8544) );
  nor_x1_sg U54968 ( .A(n8547), .B(n8548), .X(n8546) );
  nand_x1_sg U54969 ( .A(n8548), .B(n8547), .X(n8549) );
  nor_x1_sg U54970 ( .A(n47927), .B(n9366), .X(n9364) );
  nor_x1_sg U54971 ( .A(n9367), .B(n9368), .X(n9366) );
  nand_x1_sg U54972 ( .A(n9368), .B(n9367), .X(n9369) );
  nor_x1_sg U54973 ( .A(n48212), .B(n10185), .X(n10183) );
  nor_x1_sg U54974 ( .A(n10186), .B(n10187), .X(n10185) );
  nand_x1_sg U54975 ( .A(n10187), .B(n10186), .X(n10188) );
  nor_x1_sg U54976 ( .A(n48497), .B(n11004), .X(n11002) );
  nor_x1_sg U54977 ( .A(n11005), .B(n11006), .X(n11004) );
  nand_x1_sg U54978 ( .A(n11006), .B(n11005), .X(n11007) );
  nor_x1_sg U54979 ( .A(n48782), .B(n11823), .X(n11821) );
  nor_x1_sg U54980 ( .A(n11824), .B(n11825), .X(n11823) );
  nand_x1_sg U54981 ( .A(n11825), .B(n11824), .X(n11826) );
  nor_x1_sg U54982 ( .A(n49069), .B(n12642), .X(n12640) );
  nor_x1_sg U54983 ( .A(n12643), .B(n12644), .X(n12642) );
  nand_x1_sg U54984 ( .A(n12644), .B(n12643), .X(n12645) );
  nor_x1_sg U54985 ( .A(n49355), .B(n13461), .X(n13459) );
  nor_x1_sg U54986 ( .A(n13462), .B(n13463), .X(n13461) );
  nand_x1_sg U54987 ( .A(n13463), .B(n13462), .X(n13464) );
  nor_x1_sg U54988 ( .A(n49641), .B(n14280), .X(n14278) );
  nor_x1_sg U54989 ( .A(n14281), .B(n14282), .X(n14280) );
  nand_x1_sg U54990 ( .A(n14282), .B(n14281), .X(n14283) );
  nor_x1_sg U54991 ( .A(n49927), .B(n15099), .X(n15097) );
  nor_x1_sg U54992 ( .A(n15100), .B(n15101), .X(n15099) );
  nand_x1_sg U54993 ( .A(n15101), .B(n15100), .X(n15102) );
  nor_x1_sg U54994 ( .A(n50213), .B(n15918), .X(n15916) );
  nor_x1_sg U54995 ( .A(n15919), .B(n15920), .X(n15918) );
  nand_x1_sg U54996 ( .A(n15920), .B(n15919), .X(n15921) );
  nor_x1_sg U54997 ( .A(n50446), .B(n16723), .X(n16721) );
  nor_x1_sg U54998 ( .A(n16724), .B(n16725), .X(n16723) );
  nand_x1_sg U54999 ( .A(n16725), .B(n16724), .X(n16726) );
  nor_x1_sg U55000 ( .A(n50471), .B(n16729), .X(n16727) );
  nor_x1_sg U55001 ( .A(n16730), .B(n16731), .X(n16729) );
  nand_x1_sg U55002 ( .A(n16731), .B(n16730), .X(n16732) );
  nor_x1_sg U55003 ( .A(n50787), .B(n17556), .X(n17554) );
  nor_x1_sg U55004 ( .A(n17557), .B(n17558), .X(n17556) );
  nand_x1_sg U55005 ( .A(n17558), .B(n17557), .X(n17559) );
  nor_x1_sg U55006 ( .A(n51074), .B(n18377), .X(n18375) );
  nor_x1_sg U55007 ( .A(n18378), .B(n18379), .X(n18377) );
  nand_x1_sg U55008 ( .A(n18379), .B(n18378), .X(n18380) );
  nor_x1_sg U55009 ( .A(n7407), .B(n7408), .X(n7406) );
  nor_x1_sg U55010 ( .A(n8225), .B(n8226), .X(n8224) );
  nor_x1_sg U55011 ( .A(n9043), .B(n9044), .X(n9042) );
  nor_x1_sg U55012 ( .A(n9863), .B(n9864), .X(n9862) );
  nor_x1_sg U55013 ( .A(n10682), .B(n10683), .X(n10681) );
  nor_x1_sg U55014 ( .A(n11501), .B(n11502), .X(n11500) );
  nor_x1_sg U55015 ( .A(n12320), .B(n12321), .X(n12319) );
  nor_x1_sg U55016 ( .A(n13139), .B(n13140), .X(n13138) );
  nor_x1_sg U55017 ( .A(n13958), .B(n13959), .X(n13957) );
  nor_x1_sg U55018 ( .A(n14777), .B(n14778), .X(n14776) );
  nor_x1_sg U55019 ( .A(n15596), .B(n15597), .X(n15595) );
  nor_x1_sg U55020 ( .A(n16415), .B(n16416), .X(n16414) );
  nor_x1_sg U55021 ( .A(n17232), .B(n17233), .X(n17231) );
  nor_x1_sg U55022 ( .A(n18053), .B(n18054), .X(n18052) );
  nor_x1_sg U55023 ( .A(n18874), .B(n18875), .X(n18873) );
  nor_x1_sg U55024 ( .A(n7350), .B(n7351), .X(n7349) );
  nor_x1_sg U55025 ( .A(n7455), .B(n7456), .X(n7454) );
  nor_x1_sg U55026 ( .A(n8168), .B(n8169), .X(n8167) );
  nor_x1_sg U55027 ( .A(n8273), .B(n8274), .X(n8272) );
  nor_x1_sg U55028 ( .A(n8986), .B(n8987), .X(n8985) );
  nor_x1_sg U55029 ( .A(n9091), .B(n9092), .X(n9090) );
  nor_x1_sg U55030 ( .A(n9806), .B(n9807), .X(n9805) );
  nor_x1_sg U55031 ( .A(n9911), .B(n9912), .X(n9910) );
  nor_x1_sg U55032 ( .A(n10625), .B(n10626), .X(n10624) );
  nor_x1_sg U55033 ( .A(n10730), .B(n10731), .X(n10729) );
  nor_x1_sg U55034 ( .A(n11444), .B(n11445), .X(n11443) );
  nor_x1_sg U55035 ( .A(n11549), .B(n11550), .X(n11548) );
  nor_x1_sg U55036 ( .A(n12263), .B(n12264), .X(n12262) );
  nor_x1_sg U55037 ( .A(n12368), .B(n12369), .X(n12367) );
  nor_x1_sg U55038 ( .A(n13082), .B(n13083), .X(n13081) );
  nor_x1_sg U55039 ( .A(n13187), .B(n13188), .X(n13186) );
  nor_x1_sg U55040 ( .A(n13901), .B(n13902), .X(n13900) );
  nor_x1_sg U55041 ( .A(n14006), .B(n14007), .X(n14005) );
  nor_x1_sg U55042 ( .A(n14720), .B(n14721), .X(n14719) );
  nor_x1_sg U55043 ( .A(n14825), .B(n14826), .X(n14824) );
  nor_x1_sg U55044 ( .A(n15539), .B(n15540), .X(n15538) );
  nor_x1_sg U55045 ( .A(n15644), .B(n15645), .X(n15643) );
  nor_x1_sg U55046 ( .A(n16358), .B(n16359), .X(n16357) );
  nor_x1_sg U55047 ( .A(n16463), .B(n16464), .X(n16462) );
  nor_x1_sg U55048 ( .A(n17175), .B(n17176), .X(n17174) );
  nor_x1_sg U55049 ( .A(n17280), .B(n17281), .X(n17279) );
  nor_x1_sg U55050 ( .A(n17996), .B(n17997), .X(n17995) );
  nor_x1_sg U55051 ( .A(n18101), .B(n18102), .X(n18100) );
  nor_x1_sg U55052 ( .A(n18817), .B(n18818), .X(n18816) );
  nor_x1_sg U55053 ( .A(n18922), .B(n18923), .X(n18921) );
  nor_x1_sg U55054 ( .A(n7383), .B(n7384), .X(n7382) );
  nor_x1_sg U55055 ( .A(n8201), .B(n8202), .X(n8200) );
  nor_x1_sg U55056 ( .A(n9019), .B(n9020), .X(n9018) );
  nor_x1_sg U55057 ( .A(n9839), .B(n9840), .X(n9838) );
  nor_x1_sg U55058 ( .A(n10658), .B(n10659), .X(n10657) );
  nor_x1_sg U55059 ( .A(n11477), .B(n11478), .X(n11476) );
  nor_x1_sg U55060 ( .A(n12296), .B(n12297), .X(n12295) );
  nor_x1_sg U55061 ( .A(n13115), .B(n13116), .X(n13114) );
  nor_x1_sg U55062 ( .A(n13934), .B(n13935), .X(n13933) );
  nor_x1_sg U55063 ( .A(n14753), .B(n14754), .X(n14752) );
  nor_x1_sg U55064 ( .A(n15572), .B(n15573), .X(n15571) );
  nor_x1_sg U55065 ( .A(n16391), .B(n16392), .X(n16390) );
  nor_x1_sg U55066 ( .A(n17208), .B(n17209), .X(n17207) );
  nor_x1_sg U55067 ( .A(n18029), .B(n18030), .X(n18028) );
  nor_x1_sg U55068 ( .A(n18850), .B(n18851), .X(n18849) );
  inv_x1_sg U55069 ( .A(n6907), .X(n47042) );
  inv_x1_sg U55070 ( .A(n16731), .X(n50470) );
  inv_x1_sg U55071 ( .A(n6901), .X(n47016) );
  inv_x1_sg U55072 ( .A(n7730), .X(n47356) );
  inv_x1_sg U55073 ( .A(n8548), .X(n47641) );
  inv_x1_sg U55074 ( .A(n9368), .X(n47926) );
  inv_x1_sg U55075 ( .A(n10187), .X(n48211) );
  inv_x1_sg U55076 ( .A(n11006), .X(n48496) );
  inv_x1_sg U55077 ( .A(n11825), .X(n48781) );
  inv_x1_sg U55078 ( .A(n12644), .X(n49068) );
  inv_x1_sg U55079 ( .A(n13463), .X(n49354) );
  inv_x1_sg U55080 ( .A(n14282), .X(n49640) );
  inv_x1_sg U55081 ( .A(n15101), .X(n49926) );
  inv_x1_sg U55082 ( .A(n15920), .X(n50212) );
  inv_x1_sg U55083 ( .A(n16725), .X(n50445) );
  inv_x1_sg U55084 ( .A(n17558), .X(n50786) );
  inv_x1_sg U55085 ( .A(n18379), .X(n51073) );
  inv_x1_sg U55086 ( .A(n7348), .X(n47039) );
  inv_x1_sg U55087 ( .A(n8166), .X(n47326) );
  inv_x1_sg U55088 ( .A(n8984), .X(n47611) );
  inv_x1_sg U55089 ( .A(n9804), .X(n47896) );
  inv_x1_sg U55090 ( .A(n10623), .X(n48181) );
  inv_x1_sg U55091 ( .A(n11442), .X(n48466) );
  inv_x1_sg U55092 ( .A(n12261), .X(n48751) );
  inv_x1_sg U55093 ( .A(n13080), .X(n49037) );
  inv_x1_sg U55094 ( .A(n13899), .X(n49324) );
  inv_x1_sg U55095 ( .A(n14718), .X(n49610) );
  inv_x1_sg U55096 ( .A(n15537), .X(n49896) );
  inv_x1_sg U55097 ( .A(n16356), .X(n50182) );
  inv_x1_sg U55098 ( .A(n17173), .X(n50467) );
  inv_x1_sg U55099 ( .A(n17994), .X(n50756) );
  inv_x1_sg U55100 ( .A(n18815), .X(n51043) );
  nand_x1_sg U55101 ( .A(n7348), .B(n42254), .X(n7345) );
  nor_x1_sg U55102 ( .A(n42254), .B(n7348), .X(n7346) );
  nand_x1_sg U55103 ( .A(n8166), .B(n42253), .X(n8163) );
  nor_x1_sg U55104 ( .A(n42253), .B(n8166), .X(n8164) );
  nand_x1_sg U55105 ( .A(n8984), .B(n42252), .X(n8981) );
  nor_x1_sg U55106 ( .A(n42252), .B(n8984), .X(n8982) );
  nand_x1_sg U55107 ( .A(n9804), .B(n42251), .X(n9801) );
  nor_x1_sg U55108 ( .A(n42251), .B(n9804), .X(n9802) );
  nand_x1_sg U55109 ( .A(n10623), .B(n42250), .X(n10620) );
  nor_x1_sg U55110 ( .A(n42250), .B(n10623), .X(n10621) );
  nand_x1_sg U55111 ( .A(n11442), .B(n42249), .X(n11439) );
  nor_x1_sg U55112 ( .A(n42249), .B(n11442), .X(n11440) );
  nand_x1_sg U55113 ( .A(n12261), .B(n42248), .X(n12258) );
  nor_x1_sg U55114 ( .A(n42248), .B(n12261), .X(n12259) );
  nand_x1_sg U55115 ( .A(n13080), .B(n42247), .X(n13077) );
  nor_x1_sg U55116 ( .A(n42247), .B(n13080), .X(n13078) );
  nand_x1_sg U55117 ( .A(n13899), .B(n42246), .X(n13896) );
  nor_x1_sg U55118 ( .A(n42246), .B(n13899), .X(n13897) );
  nand_x1_sg U55119 ( .A(n14718), .B(n42245), .X(n14715) );
  nor_x1_sg U55120 ( .A(n42245), .B(n14718), .X(n14716) );
  nand_x1_sg U55121 ( .A(n15537), .B(n42244), .X(n15534) );
  nor_x1_sg U55122 ( .A(n42244), .B(n15537), .X(n15535) );
  nand_x1_sg U55123 ( .A(n16356), .B(n42243), .X(n16353) );
  nor_x1_sg U55124 ( .A(n42243), .B(n16356), .X(n16354) );
  nand_x1_sg U55125 ( .A(n17173), .B(n42241), .X(n17170) );
  nor_x1_sg U55126 ( .A(n42241), .B(n17173), .X(n17171) );
  nand_x1_sg U55127 ( .A(n17994), .B(n42240), .X(n17991) );
  nor_x1_sg U55128 ( .A(n42240), .B(n17994), .X(n17992) );
  nand_x1_sg U55129 ( .A(n18815), .B(n42239), .X(n18812) );
  nor_x1_sg U55130 ( .A(n42239), .B(n18815), .X(n18813) );
  nand_x1_sg U55131 ( .A(n7400), .B(n47037), .X(n7399) );
  nand_x1_sg U55132 ( .A(n8218), .B(n47324), .X(n8217) );
  nand_x1_sg U55133 ( .A(n9036), .B(n47609), .X(n9035) );
  nand_x1_sg U55134 ( .A(n9856), .B(n47894), .X(n9855) );
  nand_x1_sg U55135 ( .A(n10675), .B(n48179), .X(n10674) );
  nand_x1_sg U55136 ( .A(n11494), .B(n48464), .X(n11493) );
  nand_x1_sg U55137 ( .A(n12313), .B(n48749), .X(n12312) );
  nand_x1_sg U55138 ( .A(n13132), .B(n49035), .X(n13131) );
  nand_x1_sg U55139 ( .A(n13951), .B(n49322), .X(n13950) );
  nand_x1_sg U55140 ( .A(n14770), .B(n49608), .X(n14769) );
  nand_x1_sg U55141 ( .A(n15589), .B(n49894), .X(n15588) );
  nand_x1_sg U55142 ( .A(n16408), .B(n50180), .X(n16407) );
  nand_x1_sg U55143 ( .A(n18046), .B(n50754), .X(n18045) );
  nand_x1_sg U55144 ( .A(n18867), .B(n51041), .X(n18866) );
  inv_x1_sg U55145 ( .A(n7401), .X(n47037) );
  inv_x1_sg U55146 ( .A(n8219), .X(n47324) );
  inv_x1_sg U55147 ( .A(n9037), .X(n47609) );
  inv_x1_sg U55148 ( .A(n9857), .X(n47894) );
  inv_x1_sg U55149 ( .A(n10676), .X(n48179) );
  inv_x1_sg U55150 ( .A(n11495), .X(n48464) );
  inv_x1_sg U55151 ( .A(n12314), .X(n48749) );
  inv_x1_sg U55152 ( .A(n13133), .X(n49035) );
  inv_x1_sg U55153 ( .A(n13952), .X(n49322) );
  inv_x1_sg U55154 ( .A(n14771), .X(n49608) );
  inv_x1_sg U55155 ( .A(n15590), .X(n49894) );
  inv_x1_sg U55156 ( .A(n16409), .X(n50180) );
  inv_x1_sg U55157 ( .A(n18047), .X(n50754) );
  inv_x1_sg U55158 ( .A(n18868), .X(n51041) );
  inv_x1_sg U55159 ( .A(n7322), .X(n47013) );
  nor_x1_sg U55160 ( .A(n7320), .B(n7321), .X(n7319) );
  inv_x1_sg U55161 ( .A(n8140), .X(n47301) );
  nor_x1_sg U55162 ( .A(n8138), .B(n8139), .X(n8137) );
  inv_x1_sg U55163 ( .A(n8958), .X(n47586) );
  nor_x1_sg U55164 ( .A(n8956), .B(n8957), .X(n8955) );
  inv_x1_sg U55165 ( .A(n9778), .X(n47871) );
  nor_x1_sg U55166 ( .A(n9776), .B(n9777), .X(n9775) );
  inv_x1_sg U55167 ( .A(n10597), .X(n48156) );
  nor_x1_sg U55168 ( .A(n10595), .B(n10596), .X(n10594) );
  inv_x1_sg U55169 ( .A(n11416), .X(n48441) );
  nor_x1_sg U55170 ( .A(n11414), .B(n11415), .X(n11413) );
  inv_x1_sg U55171 ( .A(n12235), .X(n48726) );
  nor_x1_sg U55172 ( .A(n12233), .B(n12234), .X(n12232) );
  inv_x1_sg U55173 ( .A(n13054), .X(n49012) );
  nor_x1_sg U55174 ( .A(n13052), .B(n13053), .X(n13051) );
  inv_x1_sg U55175 ( .A(n13873), .X(n49299) );
  nor_x1_sg U55176 ( .A(n13871), .B(n13872), .X(n13870) );
  inv_x1_sg U55177 ( .A(n14692), .X(n49585) );
  nor_x1_sg U55178 ( .A(n14690), .B(n14691), .X(n14689) );
  inv_x1_sg U55179 ( .A(n15511), .X(n49871) );
  nor_x1_sg U55180 ( .A(n15509), .B(n15510), .X(n15508) );
  inv_x1_sg U55181 ( .A(n16330), .X(n50157) );
  nor_x1_sg U55182 ( .A(n16328), .B(n16329), .X(n16327) );
  inv_x1_sg U55183 ( .A(n17147), .X(n50442) );
  nor_x1_sg U55184 ( .A(n17145), .B(n17146), .X(n17144) );
  inv_x1_sg U55185 ( .A(n17968), .X(n50731) );
  nor_x1_sg U55186 ( .A(n17966), .B(n17967), .X(n17965) );
  inv_x1_sg U55187 ( .A(n18789), .X(n51018) );
  nor_x1_sg U55188 ( .A(n18787), .B(n18788), .X(n18786) );
  inv_x1_sg U55189 ( .A(n7409), .X(n47044) );
  nor_x1_sg U55190 ( .A(n7412), .B(n7413), .X(n7411) );
  inv_x1_sg U55191 ( .A(n8227), .X(n47331) );
  nor_x1_sg U55192 ( .A(n8230), .B(n8231), .X(n8229) );
  inv_x1_sg U55193 ( .A(n9045), .X(n47616) );
  nor_x1_sg U55194 ( .A(n9048), .B(n9049), .X(n9047) );
  inv_x1_sg U55195 ( .A(n9865), .X(n47901) );
  nor_x1_sg U55196 ( .A(n9868), .B(n9869), .X(n9867) );
  inv_x1_sg U55197 ( .A(n10684), .X(n48186) );
  nor_x1_sg U55198 ( .A(n10687), .B(n10688), .X(n10686) );
  inv_x1_sg U55199 ( .A(n11503), .X(n48471) );
  nor_x1_sg U55200 ( .A(n11506), .B(n11507), .X(n11505) );
  inv_x1_sg U55201 ( .A(n12322), .X(n48756) );
  nor_x1_sg U55202 ( .A(n12325), .B(n12326), .X(n12324) );
  inv_x1_sg U55203 ( .A(n13141), .X(n49042) );
  nor_x1_sg U55204 ( .A(n13144), .B(n13145), .X(n13143) );
  inv_x1_sg U55205 ( .A(n13960), .X(n49329) );
  nor_x1_sg U55206 ( .A(n13963), .B(n13964), .X(n13962) );
  inv_x1_sg U55207 ( .A(n14779), .X(n49615) );
  nor_x1_sg U55208 ( .A(n14782), .B(n14783), .X(n14781) );
  inv_x1_sg U55209 ( .A(n15598), .X(n49901) );
  nor_x1_sg U55210 ( .A(n15601), .B(n15602), .X(n15600) );
  inv_x1_sg U55211 ( .A(n16417), .X(n50187) );
  nor_x1_sg U55212 ( .A(n16420), .B(n16421), .X(n16419) );
  inv_x1_sg U55213 ( .A(n17234), .X(n50472) );
  nor_x1_sg U55214 ( .A(n17237), .B(n17238), .X(n17236) );
  inv_x1_sg U55215 ( .A(n18055), .X(n50761) );
  nor_x1_sg U55216 ( .A(n18058), .B(n18059), .X(n18057) );
  inv_x1_sg U55217 ( .A(n18876), .X(n51048) );
  nor_x1_sg U55218 ( .A(n18879), .B(n18880), .X(n18878) );
  nor_x1_sg U55219 ( .A(n6963), .B(n47125), .X(n6932) );
  nor_x1_sg U55220 ( .A(n6966), .B(n6965), .X(n6963) );
  nand_x1_sg U55221 ( .A(n6965), .B(n6966), .X(n6964) );
  nor_x1_sg U55222 ( .A(n7780), .B(n47411), .X(n7749) );
  nor_x1_sg U55223 ( .A(n7783), .B(n7782), .X(n7780) );
  nand_x1_sg U55224 ( .A(n7782), .B(n7783), .X(n7781) );
  nor_x1_sg U55225 ( .A(n8598), .B(n47696), .X(n8567) );
  nor_x1_sg U55226 ( .A(n8601), .B(n8600), .X(n8598) );
  nand_x1_sg U55227 ( .A(n8600), .B(n8601), .X(n8599) );
  nor_x1_sg U55228 ( .A(n9418), .B(n47981), .X(n9387) );
  nor_x1_sg U55229 ( .A(n9421), .B(n9420), .X(n9418) );
  nand_x1_sg U55230 ( .A(n9420), .B(n9421), .X(n9419) );
  nor_x1_sg U55231 ( .A(n10237), .B(n48266), .X(n10206) );
  nor_x1_sg U55232 ( .A(n10240), .B(n10239), .X(n10237) );
  nand_x1_sg U55233 ( .A(n10239), .B(n10240), .X(n10238) );
  nor_x1_sg U55234 ( .A(n11056), .B(n48551), .X(n11025) );
  nor_x1_sg U55235 ( .A(n11059), .B(n11058), .X(n11056) );
  nand_x1_sg U55236 ( .A(n11058), .B(n11059), .X(n11057) );
  nor_x1_sg U55237 ( .A(n11875), .B(n48836), .X(n11844) );
  nor_x1_sg U55238 ( .A(n11878), .B(n11877), .X(n11875) );
  nand_x1_sg U55239 ( .A(n11877), .B(n11878), .X(n11876) );
  nor_x1_sg U55240 ( .A(n12694), .B(n49123), .X(n12663) );
  nor_x1_sg U55241 ( .A(n12697), .B(n12696), .X(n12694) );
  nand_x1_sg U55242 ( .A(n12696), .B(n12697), .X(n12695) );
  nor_x1_sg U55243 ( .A(n13513), .B(n49409), .X(n13482) );
  nor_x1_sg U55244 ( .A(n13516), .B(n13515), .X(n13513) );
  nand_x1_sg U55245 ( .A(n13515), .B(n13516), .X(n13514) );
  nor_x1_sg U55246 ( .A(n14332), .B(n49695), .X(n14301) );
  nor_x1_sg U55247 ( .A(n14335), .B(n14334), .X(n14332) );
  nand_x1_sg U55248 ( .A(n14334), .B(n14335), .X(n14333) );
  nor_x1_sg U55249 ( .A(n15151), .B(n49981), .X(n15120) );
  nor_x1_sg U55250 ( .A(n15154), .B(n15153), .X(n15151) );
  nand_x1_sg U55251 ( .A(n15153), .B(n15154), .X(n15152) );
  nor_x1_sg U55252 ( .A(n15970), .B(n50267), .X(n15939) );
  nor_x1_sg U55253 ( .A(n15973), .B(n15972), .X(n15970) );
  nand_x1_sg U55254 ( .A(n15972), .B(n15973), .X(n15971) );
  nor_x1_sg U55255 ( .A(n16787), .B(n50553), .X(n16756) );
  nor_x1_sg U55256 ( .A(n16790), .B(n16789), .X(n16787) );
  nand_x1_sg U55257 ( .A(n16789), .B(n16790), .X(n16788) );
  nor_x1_sg U55258 ( .A(n17608), .B(n50841), .X(n17577) );
  nor_x1_sg U55259 ( .A(n17611), .B(n17610), .X(n17608) );
  nand_x1_sg U55260 ( .A(n17610), .B(n17611), .X(n17609) );
  nor_x1_sg U55261 ( .A(n18429), .B(n51128), .X(n18398) );
  nor_x1_sg U55262 ( .A(n18432), .B(n18431), .X(n18429) );
  nand_x1_sg U55263 ( .A(n18431), .B(n18432), .X(n18430) );
  nor_x1_sg U55264 ( .A(n6972), .B(n47124), .X(n6966) );
  nor_x1_sg U55265 ( .A(n6975), .B(n6974), .X(n6972) );
  nor_x1_sg U55266 ( .A(n7789), .B(n47410), .X(n7783) );
  nor_x1_sg U55267 ( .A(n7792), .B(n7791), .X(n7789) );
  nor_x1_sg U55268 ( .A(n8607), .B(n47695), .X(n8601) );
  nor_x1_sg U55269 ( .A(n8610), .B(n8609), .X(n8607) );
  nor_x1_sg U55270 ( .A(n9427), .B(n47980), .X(n9421) );
  nor_x1_sg U55271 ( .A(n9430), .B(n9429), .X(n9427) );
  nor_x1_sg U55272 ( .A(n10246), .B(n48265), .X(n10240) );
  nor_x1_sg U55273 ( .A(n10249), .B(n10248), .X(n10246) );
  nor_x1_sg U55274 ( .A(n11065), .B(n48550), .X(n11059) );
  nor_x1_sg U55275 ( .A(n11068), .B(n11067), .X(n11065) );
  nor_x1_sg U55276 ( .A(n11884), .B(n48835), .X(n11878) );
  nor_x1_sg U55277 ( .A(n11887), .B(n11886), .X(n11884) );
  nor_x1_sg U55278 ( .A(n12703), .B(n49122), .X(n12697) );
  nor_x1_sg U55279 ( .A(n12706), .B(n12705), .X(n12703) );
  nor_x1_sg U55280 ( .A(n13522), .B(n49408), .X(n13516) );
  nor_x1_sg U55281 ( .A(n13525), .B(n13524), .X(n13522) );
  nor_x1_sg U55282 ( .A(n14341), .B(n49694), .X(n14335) );
  nor_x1_sg U55283 ( .A(n14344), .B(n14343), .X(n14341) );
  nor_x1_sg U55284 ( .A(n15160), .B(n49980), .X(n15154) );
  nor_x1_sg U55285 ( .A(n15163), .B(n15162), .X(n15160) );
  nor_x1_sg U55286 ( .A(n15979), .B(n50266), .X(n15973) );
  nor_x1_sg U55287 ( .A(n15982), .B(n15981), .X(n15979) );
  nor_x1_sg U55288 ( .A(n16796), .B(n50552), .X(n16790) );
  nor_x1_sg U55289 ( .A(n16799), .B(n16798), .X(n16796) );
  nor_x1_sg U55290 ( .A(n17617), .B(n50840), .X(n17611) );
  nor_x1_sg U55291 ( .A(n17620), .B(n17619), .X(n17617) );
  nor_x1_sg U55292 ( .A(n18438), .B(n51127), .X(n18432) );
  nor_x1_sg U55293 ( .A(n18441), .B(n18440), .X(n18438) );
  nor_x1_sg U55294 ( .A(n47003), .B(n6893), .X(n6891) );
  nor_x1_sg U55295 ( .A(n6894), .B(n6895), .X(n6893) );
  nand_x1_sg U55296 ( .A(n6895), .B(n6894), .X(n6896) );
  nor_x1_sg U55297 ( .A(n47292), .B(n7710), .X(n7708) );
  nor_x1_sg U55298 ( .A(n7711), .B(n7712), .X(n7710) );
  nand_x1_sg U55299 ( .A(n7712), .B(n7711), .X(n7713) );
  nor_x1_sg U55300 ( .A(n47305), .B(n7716), .X(n7714) );
  nor_x1_sg U55301 ( .A(n7717), .B(n7718), .X(n7716) );
  nand_x1_sg U55302 ( .A(n7718), .B(n7717), .X(n7719) );
  nor_x1_sg U55303 ( .A(n47330), .B(n7722), .X(n7720) );
  nor_x1_sg U55304 ( .A(n7723), .B(n7724), .X(n7722) );
  nand_x1_sg U55305 ( .A(n7724), .B(n7723), .X(n7725) );
  nor_x1_sg U55306 ( .A(n47577), .B(n8528), .X(n8526) );
  nor_x1_sg U55307 ( .A(n8529), .B(n8530), .X(n8528) );
  nand_x1_sg U55308 ( .A(n8530), .B(n8529), .X(n8531) );
  nor_x1_sg U55309 ( .A(n47590), .B(n8534), .X(n8532) );
  nor_x1_sg U55310 ( .A(n8535), .B(n8536), .X(n8534) );
  nand_x1_sg U55311 ( .A(n8536), .B(n8535), .X(n8537) );
  nor_x1_sg U55312 ( .A(n47615), .B(n8540), .X(n8538) );
  nor_x1_sg U55313 ( .A(n8541), .B(n8542), .X(n8540) );
  nand_x1_sg U55314 ( .A(n8542), .B(n8541), .X(n8543) );
  nor_x1_sg U55315 ( .A(n47862), .B(n9348), .X(n9346) );
  nor_x1_sg U55316 ( .A(n9349), .B(n9350), .X(n9348) );
  nand_x1_sg U55317 ( .A(n9350), .B(n9349), .X(n9351) );
  nor_x1_sg U55318 ( .A(n47875), .B(n9354), .X(n9352) );
  nor_x1_sg U55319 ( .A(n9355), .B(n9356), .X(n9354) );
  nand_x1_sg U55320 ( .A(n9356), .B(n9355), .X(n9357) );
  nor_x1_sg U55321 ( .A(n47900), .B(n9360), .X(n9358) );
  nor_x1_sg U55322 ( .A(n9361), .B(n9362), .X(n9360) );
  nand_x1_sg U55323 ( .A(n9362), .B(n9361), .X(n9363) );
  nor_x1_sg U55324 ( .A(n48147), .B(n10167), .X(n10165) );
  nor_x1_sg U55325 ( .A(n10168), .B(n10169), .X(n10167) );
  nand_x1_sg U55326 ( .A(n10169), .B(n10168), .X(n10170) );
  nor_x1_sg U55327 ( .A(n48160), .B(n10173), .X(n10171) );
  nor_x1_sg U55328 ( .A(n10174), .B(n10175), .X(n10173) );
  nand_x1_sg U55329 ( .A(n10175), .B(n10174), .X(n10176) );
  nor_x1_sg U55330 ( .A(n48185), .B(n10179), .X(n10177) );
  nor_x1_sg U55331 ( .A(n10180), .B(n10181), .X(n10179) );
  nand_x1_sg U55332 ( .A(n10181), .B(n10180), .X(n10182) );
  nor_x1_sg U55333 ( .A(n48432), .B(n10986), .X(n10984) );
  nor_x1_sg U55334 ( .A(n10987), .B(n10988), .X(n10986) );
  nand_x1_sg U55335 ( .A(n10988), .B(n10987), .X(n10989) );
  nor_x1_sg U55336 ( .A(n48445), .B(n10992), .X(n10990) );
  nor_x1_sg U55337 ( .A(n10993), .B(n10994), .X(n10992) );
  nand_x1_sg U55338 ( .A(n10994), .B(n10993), .X(n10995) );
  nor_x1_sg U55339 ( .A(n48470), .B(n10998), .X(n10996) );
  nor_x1_sg U55340 ( .A(n10999), .B(n11000), .X(n10998) );
  nand_x1_sg U55341 ( .A(n11000), .B(n10999), .X(n11001) );
  nor_x1_sg U55342 ( .A(n48717), .B(n11805), .X(n11803) );
  nor_x1_sg U55343 ( .A(n11806), .B(n11807), .X(n11805) );
  nand_x1_sg U55344 ( .A(n11807), .B(n11806), .X(n11808) );
  nor_x1_sg U55345 ( .A(n48730), .B(n11811), .X(n11809) );
  nor_x1_sg U55346 ( .A(n11812), .B(n11813), .X(n11811) );
  nand_x1_sg U55347 ( .A(n11813), .B(n11812), .X(n11814) );
  nor_x1_sg U55348 ( .A(n48755), .B(n11817), .X(n11815) );
  nor_x1_sg U55349 ( .A(n11818), .B(n11819), .X(n11817) );
  nand_x1_sg U55350 ( .A(n11819), .B(n11818), .X(n11820) );
  nor_x1_sg U55351 ( .A(n49003), .B(n12624), .X(n12622) );
  nor_x1_sg U55352 ( .A(n12625), .B(n12626), .X(n12624) );
  nand_x1_sg U55353 ( .A(n12626), .B(n12625), .X(n12627) );
  nor_x1_sg U55354 ( .A(n49016), .B(n12630), .X(n12628) );
  nor_x1_sg U55355 ( .A(n12631), .B(n12632), .X(n12630) );
  nand_x1_sg U55356 ( .A(n12632), .B(n12631), .X(n12633) );
  nor_x1_sg U55357 ( .A(n49041), .B(n12636), .X(n12634) );
  nor_x1_sg U55358 ( .A(n12637), .B(n12638), .X(n12636) );
  nand_x1_sg U55359 ( .A(n12638), .B(n12637), .X(n12639) );
  nor_x1_sg U55360 ( .A(n49290), .B(n13443), .X(n13441) );
  nor_x1_sg U55361 ( .A(n13444), .B(n13445), .X(n13443) );
  nand_x1_sg U55362 ( .A(n13445), .B(n13444), .X(n13446) );
  nor_x1_sg U55363 ( .A(n49303), .B(n13449), .X(n13447) );
  nor_x1_sg U55364 ( .A(n13450), .B(n13451), .X(n13449) );
  nand_x1_sg U55365 ( .A(n13451), .B(n13450), .X(n13452) );
  nor_x1_sg U55366 ( .A(n49328), .B(n13455), .X(n13453) );
  nor_x1_sg U55367 ( .A(n13456), .B(n13457), .X(n13455) );
  nand_x1_sg U55368 ( .A(n13457), .B(n13456), .X(n13458) );
  nor_x1_sg U55369 ( .A(n49576), .B(n14262), .X(n14260) );
  nor_x1_sg U55370 ( .A(n14263), .B(n14264), .X(n14262) );
  nand_x1_sg U55371 ( .A(n14264), .B(n14263), .X(n14265) );
  nor_x1_sg U55372 ( .A(n49589), .B(n14268), .X(n14266) );
  nor_x1_sg U55373 ( .A(n14269), .B(n14270), .X(n14268) );
  nand_x1_sg U55374 ( .A(n14270), .B(n14269), .X(n14271) );
  nor_x1_sg U55375 ( .A(n49614), .B(n14274), .X(n14272) );
  nor_x1_sg U55376 ( .A(n14275), .B(n14276), .X(n14274) );
  nand_x1_sg U55377 ( .A(n14276), .B(n14275), .X(n14277) );
  nor_x1_sg U55378 ( .A(n49862), .B(n15081), .X(n15079) );
  nor_x1_sg U55379 ( .A(n15082), .B(n15083), .X(n15081) );
  nand_x1_sg U55380 ( .A(n15083), .B(n15082), .X(n15084) );
  nor_x1_sg U55381 ( .A(n49875), .B(n15087), .X(n15085) );
  nor_x1_sg U55382 ( .A(n15088), .B(n15089), .X(n15087) );
  nand_x1_sg U55383 ( .A(n15089), .B(n15088), .X(n15090) );
  nor_x1_sg U55384 ( .A(n49900), .B(n15093), .X(n15091) );
  nor_x1_sg U55385 ( .A(n15094), .B(n15095), .X(n15093) );
  nand_x1_sg U55386 ( .A(n15095), .B(n15094), .X(n15096) );
  nor_x1_sg U55387 ( .A(n50148), .B(n15900), .X(n15898) );
  nor_x1_sg U55388 ( .A(n15901), .B(n15902), .X(n15900) );
  nand_x1_sg U55389 ( .A(n15902), .B(n15901), .X(n15903) );
  nor_x1_sg U55390 ( .A(n50161), .B(n15906), .X(n15904) );
  nor_x1_sg U55391 ( .A(n15907), .B(n15908), .X(n15906) );
  nand_x1_sg U55392 ( .A(n15908), .B(n15907), .X(n15909) );
  nor_x1_sg U55393 ( .A(n50186), .B(n15912), .X(n15910) );
  nor_x1_sg U55394 ( .A(n15913), .B(n15914), .X(n15912) );
  nand_x1_sg U55395 ( .A(n15914), .B(n15913), .X(n15915) );
  nor_x1_sg U55396 ( .A(n50307), .B(n16675), .X(n16673) );
  nor_x1_sg U55397 ( .A(n16676), .B(n50306), .X(n16675) );
  nand_x1_sg U55398 ( .A(n50306), .B(n16676), .X(n16677) );
  nor_x1_sg U55399 ( .A(n50411), .B(n16711), .X(n16709) );
  nor_x1_sg U55400 ( .A(n16712), .B(n16713), .X(n16711) );
  nand_x1_sg U55401 ( .A(n16713), .B(n16712), .X(n16714) );
  nor_x1_sg U55402 ( .A(n50433), .B(n16717), .X(n16715) );
  nor_x1_sg U55403 ( .A(n16718), .B(n16719), .X(n16717) );
  nand_x1_sg U55404 ( .A(n16719), .B(n16718), .X(n16720) );
  nor_x1_sg U55405 ( .A(n50722), .B(n17538), .X(n17536) );
  nor_x1_sg U55406 ( .A(n17539), .B(n17540), .X(n17538) );
  nand_x1_sg U55407 ( .A(n17540), .B(n17539), .X(n17541) );
  nor_x1_sg U55408 ( .A(n50735), .B(n17544), .X(n17542) );
  nor_x1_sg U55409 ( .A(n17545), .B(n17546), .X(n17544) );
  nand_x1_sg U55410 ( .A(n17546), .B(n17545), .X(n17547) );
  nor_x1_sg U55411 ( .A(n50760), .B(n17550), .X(n17548) );
  nor_x1_sg U55412 ( .A(n17551), .B(n17552), .X(n17550) );
  nand_x1_sg U55413 ( .A(n17552), .B(n17551), .X(n17553) );
  nor_x1_sg U55414 ( .A(n51009), .B(n18359), .X(n18357) );
  nor_x1_sg U55415 ( .A(n18360), .B(n18361), .X(n18359) );
  nand_x1_sg U55416 ( .A(n18361), .B(n18360), .X(n18362) );
  nor_x1_sg U55417 ( .A(n51022), .B(n18365), .X(n18363) );
  nor_x1_sg U55418 ( .A(n18366), .B(n18367), .X(n18365) );
  nand_x1_sg U55419 ( .A(n18367), .B(n18366), .X(n18368) );
  nor_x1_sg U55420 ( .A(n51047), .B(n18371), .X(n18369) );
  nor_x1_sg U55421 ( .A(n18372), .B(n18373), .X(n18371) );
  nand_x1_sg U55422 ( .A(n18373), .B(n18372), .X(n18374) );
  nor_x1_sg U55423 ( .A(n8048), .B(n8049), .X(n8047) );
  nor_x1_sg U55424 ( .A(n8866), .B(n8867), .X(n8865) );
  nor_x1_sg U55425 ( .A(n9686), .B(n9687), .X(n9685) );
  nor_x1_sg U55426 ( .A(n10505), .B(n10506), .X(n10504) );
  nor_x1_sg U55427 ( .A(n11324), .B(n11325), .X(n11323) );
  nor_x1_sg U55428 ( .A(n12143), .B(n12144), .X(n12142) );
  nor_x1_sg U55429 ( .A(n12962), .B(n12963), .X(n12961) );
  nor_x1_sg U55430 ( .A(n13781), .B(n13782), .X(n13780) );
  nor_x1_sg U55431 ( .A(n14600), .B(n14601), .X(n14599) );
  nor_x1_sg U55432 ( .A(n15419), .B(n15420), .X(n15418) );
  nor_x1_sg U55433 ( .A(n16238), .B(n16239), .X(n16237) );
  nor_x1_sg U55434 ( .A(n17876), .B(n17877), .X(n17875) );
  nor_x1_sg U55435 ( .A(n18697), .B(n18698), .X(n18696) );
  nor_x1_sg U55436 ( .A(n7315), .B(n7316), .X(n7314) );
  nor_x1_sg U55437 ( .A(n7523), .B(n7524), .X(n7522) );
  nor_x1_sg U55438 ( .A(n8341), .B(n8342), .X(n8340) );
  nor_x1_sg U55439 ( .A(n9159), .B(n9160), .X(n9158) );
  nor_x1_sg U55440 ( .A(n9979), .B(n9980), .X(n9978) );
  nor_x1_sg U55441 ( .A(n10798), .B(n10799), .X(n10797) );
  nor_x1_sg U55442 ( .A(n11617), .B(n11618), .X(n11616) );
  nor_x1_sg U55443 ( .A(n12436), .B(n12437), .X(n12435) );
  nor_x1_sg U55444 ( .A(n13255), .B(n13256), .X(n13254) );
  nor_x1_sg U55445 ( .A(n14074), .B(n14075), .X(n14073) );
  nor_x1_sg U55446 ( .A(n14893), .B(n14894), .X(n14892) );
  nor_x1_sg U55447 ( .A(n15712), .B(n15713), .X(n15711) );
  nor_x1_sg U55448 ( .A(n16531), .B(n16532), .X(n16530) );
  nor_x1_sg U55449 ( .A(n17348), .B(n17349), .X(n17347) );
  nor_x1_sg U55450 ( .A(n18169), .B(n18170), .X(n18168) );
  nor_x1_sg U55451 ( .A(n18990), .B(n18991), .X(n18989) );
  nor_x1_sg U55452 ( .A(n17140), .B(n17141), .X(n17139) );
  nor_x1_sg U55453 ( .A(n7483), .B(n7484), .X(n7482) );
  nor_x1_sg U55454 ( .A(n8301), .B(n8302), .X(n8300) );
  nor_x1_sg U55455 ( .A(n9119), .B(n9120), .X(n9118) );
  nor_x1_sg U55456 ( .A(n9939), .B(n9940), .X(n9938) );
  nor_x1_sg U55457 ( .A(n10758), .B(n10759), .X(n10757) );
  nor_x1_sg U55458 ( .A(n11577), .B(n11578), .X(n11576) );
  nor_x1_sg U55459 ( .A(n12396), .B(n12397), .X(n12395) );
  nor_x1_sg U55460 ( .A(n13215), .B(n13216), .X(n13214) );
  nor_x1_sg U55461 ( .A(n14034), .B(n14035), .X(n14033) );
  nor_x1_sg U55462 ( .A(n14853), .B(n14854), .X(n14852) );
  nor_x1_sg U55463 ( .A(n15672), .B(n15673), .X(n15671) );
  nor_x1_sg U55464 ( .A(n16491), .B(n16492), .X(n16490) );
  nor_x1_sg U55465 ( .A(n17308), .B(n17309), .X(n17307) );
  nor_x1_sg U55466 ( .A(n18129), .B(n18130), .X(n18128) );
  nor_x1_sg U55467 ( .A(n18950), .B(n18951), .X(n18949) );
  nor_x1_sg U55468 ( .A(n7264), .B(n7265), .X(n7263) );
  nor_x1_sg U55469 ( .A(n17089), .B(n17090), .X(n17088) );
  nor_x1_sg U55470 ( .A(n7196), .B(n7197), .X(n7195) );
  nor_x1_sg U55471 ( .A(n8015), .B(n8016), .X(n8014) );
  nor_x1_sg U55472 ( .A(n8833), .B(n8834), .X(n8832) );
  nor_x1_sg U55473 ( .A(n9653), .B(n9654), .X(n9652) );
  nor_x1_sg U55474 ( .A(n10472), .B(n10473), .X(n10471) );
  nor_x1_sg U55475 ( .A(n11291), .B(n11292), .X(n11290) );
  nor_x1_sg U55476 ( .A(n12110), .B(n12111), .X(n12109) );
  nor_x1_sg U55477 ( .A(n12929), .B(n12930), .X(n12928) );
  nor_x1_sg U55478 ( .A(n13748), .B(n13749), .X(n13747) );
  nor_x1_sg U55479 ( .A(n14567), .B(n14568), .X(n14566) );
  nor_x1_sg U55480 ( .A(n15386), .B(n15387), .X(n15385) );
  nor_x1_sg U55481 ( .A(n16205), .B(n16206), .X(n16204) );
  nor_x1_sg U55482 ( .A(n17021), .B(n17022), .X(n17020) );
  nor_x1_sg U55483 ( .A(n17843), .B(n17844), .X(n17842) );
  nor_x1_sg U55484 ( .A(n18664), .B(n18665), .X(n18663) );
  nor_x1_sg U55485 ( .A(n7543), .B(n7544), .X(n7542) );
  nor_x1_sg U55486 ( .A(n8361), .B(n8362), .X(n8360) );
  nor_x1_sg U55487 ( .A(n9179), .B(n9180), .X(n9178) );
  nor_x1_sg U55488 ( .A(n9999), .B(n10000), .X(n9998) );
  nor_x1_sg U55489 ( .A(n10818), .B(n10819), .X(n10817) );
  nor_x1_sg U55490 ( .A(n11637), .B(n11638), .X(n11636) );
  nor_x1_sg U55491 ( .A(n12456), .B(n12457), .X(n12455) );
  nor_x1_sg U55492 ( .A(n13275), .B(n13276), .X(n13274) );
  nor_x1_sg U55493 ( .A(n14094), .B(n14095), .X(n14093) );
  nor_x1_sg U55494 ( .A(n14913), .B(n14914), .X(n14912) );
  nor_x1_sg U55495 ( .A(n15732), .B(n15733), .X(n15731) );
  nor_x1_sg U55496 ( .A(n16551), .B(n16552), .X(n16550) );
  nor_x1_sg U55497 ( .A(n17368), .B(n17369), .X(n17367) );
  nor_x1_sg U55498 ( .A(n18189), .B(n18190), .X(n18188) );
  nor_x1_sg U55499 ( .A(n19010), .B(n19011), .X(n19009) );
  nand_x1_sg U55500 ( .A(n50389), .B(n17158), .X(n17197) );
  nand_x1_sg U55501 ( .A(n50371), .B(n17199), .X(n17198) );
  nand_x1_sg U55502 ( .A(n47018), .B(n7422), .X(n7420) );
  nor_x1_sg U55503 ( .A(n7422), .B(n47018), .X(n7421) );
  nand_x1_sg U55504 ( .A(n47306), .B(n8240), .X(n8238) );
  nor_x1_sg U55505 ( .A(n8240), .B(n47306), .X(n8239) );
  nand_x1_sg U55506 ( .A(n47591), .B(n9058), .X(n9056) );
  nor_x1_sg U55507 ( .A(n9058), .B(n47591), .X(n9057) );
  nand_x1_sg U55508 ( .A(n47876), .B(n9878), .X(n9876) );
  nor_x1_sg U55509 ( .A(n9878), .B(n47876), .X(n9877) );
  nand_x1_sg U55510 ( .A(n48161), .B(n10697), .X(n10695) );
  nor_x1_sg U55511 ( .A(n10697), .B(n48161), .X(n10696) );
  nand_x1_sg U55512 ( .A(n48446), .B(n11516), .X(n11514) );
  nor_x1_sg U55513 ( .A(n11516), .B(n48446), .X(n11515) );
  nand_x1_sg U55514 ( .A(n48731), .B(n12335), .X(n12333) );
  nor_x1_sg U55515 ( .A(n12335), .B(n48731), .X(n12334) );
  nand_x1_sg U55516 ( .A(n49017), .B(n13154), .X(n13152) );
  nor_x1_sg U55517 ( .A(n13154), .B(n49017), .X(n13153) );
  nand_x1_sg U55518 ( .A(n49304), .B(n13973), .X(n13971) );
  nor_x1_sg U55519 ( .A(n13973), .B(n49304), .X(n13972) );
  nand_x1_sg U55520 ( .A(n49590), .B(n14792), .X(n14790) );
  nor_x1_sg U55521 ( .A(n14792), .B(n49590), .X(n14791) );
  nand_x1_sg U55522 ( .A(n49876), .B(n15611), .X(n15609) );
  nor_x1_sg U55523 ( .A(n15611), .B(n49876), .X(n15610) );
  nand_x1_sg U55524 ( .A(n50162), .B(n16430), .X(n16428) );
  nor_x1_sg U55525 ( .A(n16430), .B(n50162), .X(n16429) );
  nand_x1_sg U55526 ( .A(n50736), .B(n18068), .X(n18066) );
  nor_x1_sg U55527 ( .A(n18068), .B(n50736), .X(n18067) );
  nand_x1_sg U55528 ( .A(n51023), .B(n18889), .X(n18887) );
  nor_x1_sg U55529 ( .A(n18889), .B(n51023), .X(n18888) );
  nand_x1_sg U55530 ( .A(n49463), .B(n14484), .X(n14483) );
  nor_x1_sg U55531 ( .A(n14484), .B(n49463), .X(n14485) );
  nand_x1_sg U55532 ( .A(n49748), .B(n15303), .X(n15302) );
  nor_x1_sg U55533 ( .A(n15303), .B(n49748), .X(n15304) );
  nand_x1_sg U55534 ( .A(n50035), .B(n16122), .X(n16121) );
  nor_x1_sg U55535 ( .A(n16122), .B(n50035), .X(n16123) );
  nand_x1_sg U55536 ( .A(n50320), .B(n16939), .X(n16938) );
  nor_x1_sg U55537 ( .A(n16939), .B(n50320), .X(n16940) );
  nand_x1_sg U55538 ( .A(n50609), .B(n17760), .X(n17759) );
  nor_x1_sg U55539 ( .A(n17760), .B(n50609), .X(n17761) );
  nand_x1_sg U55540 ( .A(n50896), .B(n18581), .X(n18580) );
  nor_x1_sg U55541 ( .A(n18581), .B(n50896), .X(n18582) );
  nand_x1_sg U55542 ( .A(n7425), .B(n47035), .X(n7424) );
  nor_x1_sg U55543 ( .A(n47035), .B(n7425), .X(n7426) );
  nand_x1_sg U55544 ( .A(n8243), .B(n47322), .X(n8242) );
  nor_x1_sg U55545 ( .A(n47322), .B(n8243), .X(n8244) );
  nand_x1_sg U55546 ( .A(n9061), .B(n47607), .X(n9060) );
  nor_x1_sg U55547 ( .A(n47607), .B(n9061), .X(n9062) );
  nand_x1_sg U55548 ( .A(n9881), .B(n47892), .X(n9880) );
  nor_x1_sg U55549 ( .A(n47892), .B(n9881), .X(n9882) );
  nand_x1_sg U55550 ( .A(n10700), .B(n48177), .X(n10699) );
  nor_x1_sg U55551 ( .A(n48177), .B(n10700), .X(n10701) );
  nand_x1_sg U55552 ( .A(n11519), .B(n48462), .X(n11518) );
  nor_x1_sg U55553 ( .A(n48462), .B(n11519), .X(n11520) );
  nand_x1_sg U55554 ( .A(n12338), .B(n48747), .X(n12337) );
  nor_x1_sg U55555 ( .A(n48747), .B(n12338), .X(n12339) );
  nand_x1_sg U55556 ( .A(n13157), .B(n49033), .X(n13156) );
  nor_x1_sg U55557 ( .A(n49033), .B(n13157), .X(n13158) );
  nand_x1_sg U55558 ( .A(n13976), .B(n49320), .X(n13975) );
  nor_x1_sg U55559 ( .A(n49320), .B(n13976), .X(n13977) );
  nand_x1_sg U55560 ( .A(n14795), .B(n49606), .X(n14794) );
  nor_x1_sg U55561 ( .A(n49606), .B(n14795), .X(n14796) );
  nand_x1_sg U55562 ( .A(n15614), .B(n49892), .X(n15613) );
  nor_x1_sg U55563 ( .A(n49892), .B(n15614), .X(n15615) );
  nand_x1_sg U55564 ( .A(n16433), .B(n50178), .X(n16432) );
  nor_x1_sg U55565 ( .A(n50178), .B(n16433), .X(n16434) );
  nand_x1_sg U55566 ( .A(n17250), .B(n50463), .X(n17249) );
  nor_x1_sg U55567 ( .A(n50463), .B(n17250), .X(n17251) );
  nand_x1_sg U55568 ( .A(n18071), .B(n50752), .X(n18070) );
  nor_x1_sg U55569 ( .A(n50752), .B(n18071), .X(n18072) );
  nand_x1_sg U55570 ( .A(n18892), .B(n51039), .X(n18891) );
  nor_x1_sg U55571 ( .A(n51039), .B(n18892), .X(n18893) );
  nand_x1_sg U55572 ( .A(n46886), .B(n7114), .X(n7113) );
  nor_x1_sg U55573 ( .A(n7114), .B(n46886), .X(n7115) );
  nand_x1_sg U55574 ( .A(n47179), .B(n7932), .X(n7931) );
  nor_x1_sg U55575 ( .A(n7932), .B(n47179), .X(n7933) );
  nand_x1_sg U55576 ( .A(n47464), .B(n8750), .X(n8749) );
  nor_x1_sg U55577 ( .A(n8750), .B(n47464), .X(n8751) );
  nand_x1_sg U55578 ( .A(n47749), .B(n9570), .X(n9569) );
  nor_x1_sg U55579 ( .A(n9570), .B(n47749), .X(n9571) );
  nand_x1_sg U55580 ( .A(n48034), .B(n10389), .X(n10388) );
  nor_x1_sg U55581 ( .A(n10389), .B(n48034), .X(n10390) );
  nand_x1_sg U55582 ( .A(n48319), .B(n11208), .X(n11207) );
  nor_x1_sg U55583 ( .A(n11208), .B(n48319), .X(n11209) );
  nand_x1_sg U55584 ( .A(n48604), .B(n12027), .X(n12026) );
  nor_x1_sg U55585 ( .A(n12027), .B(n48604), .X(n12028) );
  nand_x1_sg U55586 ( .A(n48890), .B(n12846), .X(n12845) );
  nor_x1_sg U55587 ( .A(n12846), .B(n48890), .X(n12847) );
  nand_x1_sg U55588 ( .A(n49177), .B(n13665), .X(n13664) );
  nor_x1_sg U55589 ( .A(n13665), .B(n49177), .X(n13666) );
  inv_x1_sg U55590 ( .A(n6895), .X(n47002) );
  inv_x1_sg U55591 ( .A(n7712), .X(n47291) );
  inv_x1_sg U55592 ( .A(n8530), .X(n47576) );
  inv_x1_sg U55593 ( .A(n9350), .X(n47861) );
  inv_x1_sg U55594 ( .A(n10169), .X(n48146) );
  inv_x1_sg U55595 ( .A(n10988), .X(n48431) );
  inv_x1_sg U55596 ( .A(n11807), .X(n48716) );
  inv_x1_sg U55597 ( .A(n12626), .X(n49002) );
  inv_x1_sg U55598 ( .A(n13445), .X(n49289) );
  inv_x1_sg U55599 ( .A(n14264), .X(n49575) );
  inv_x1_sg U55600 ( .A(n15083), .X(n49861) );
  inv_x1_sg U55601 ( .A(n15902), .X(n50147) );
  inv_x1_sg U55602 ( .A(n16719), .X(n50432) );
  inv_x1_sg U55603 ( .A(n17540), .X(n50721) );
  inv_x1_sg U55604 ( .A(n18361), .X(n51008) );
  inv_x1_sg U55605 ( .A(n7724), .X(n47329) );
  inv_x1_sg U55606 ( .A(n8542), .X(n47614) );
  inv_x1_sg U55607 ( .A(n9362), .X(n47899) );
  inv_x1_sg U55608 ( .A(n10181), .X(n48184) );
  inv_x1_sg U55609 ( .A(n11000), .X(n48469) );
  inv_x1_sg U55610 ( .A(n11819), .X(n48754) );
  inv_x1_sg U55611 ( .A(n12638), .X(n49040) );
  inv_x1_sg U55612 ( .A(n13457), .X(n49327) );
  inv_x1_sg U55613 ( .A(n14276), .X(n49613) );
  inv_x1_sg U55614 ( .A(n15095), .X(n49899) );
  inv_x1_sg U55615 ( .A(n15914), .X(n50185) );
  inv_x1_sg U55616 ( .A(n17552), .X(n50759) );
  inv_x1_sg U55617 ( .A(n18373), .X(n51046) );
  inv_x1_sg U55618 ( .A(n7718), .X(n47304) );
  inv_x1_sg U55619 ( .A(n8536), .X(n47589) );
  inv_x1_sg U55620 ( .A(n9356), .X(n47874) );
  inv_x1_sg U55621 ( .A(n10175), .X(n48159) );
  inv_x1_sg U55622 ( .A(n10994), .X(n48444) );
  inv_x1_sg U55623 ( .A(n11813), .X(n48729) );
  inv_x1_sg U55624 ( .A(n12632), .X(n49015) );
  inv_x1_sg U55625 ( .A(n13451), .X(n49302) );
  inv_x1_sg U55626 ( .A(n14270), .X(n49588) );
  inv_x1_sg U55627 ( .A(n15089), .X(n49874) );
  inv_x1_sg U55628 ( .A(n15908), .X(n50160) );
  inv_x1_sg U55629 ( .A(n17546), .X(n50734) );
  inv_x1_sg U55630 ( .A(n18367), .X(n51021) );
  inv_x1_sg U55631 ( .A(n16713), .X(n50410) );
  nand_x1_sg U55632 ( .A(n47259), .B(n47248), .X(n8150) );
  nand_x1_sg U55633 ( .A(n8151), .B(n8152), .X(n8149) );
  nand_x1_sg U55634 ( .A(n47544), .B(n47533), .X(n8968) );
  nand_x1_sg U55635 ( .A(n8969), .B(n8970), .X(n8967) );
  nand_x1_sg U55636 ( .A(n47829), .B(n47818), .X(n9788) );
  nand_x1_sg U55637 ( .A(n9789), .B(n9790), .X(n9787) );
  nand_x1_sg U55638 ( .A(n48114), .B(n48103), .X(n10607) );
  nand_x1_sg U55639 ( .A(n10608), .B(n10609), .X(n10606) );
  nand_x1_sg U55640 ( .A(n48399), .B(n48388), .X(n11426) );
  nand_x1_sg U55641 ( .A(n11427), .B(n11428), .X(n11425) );
  nand_x1_sg U55642 ( .A(n48684), .B(n48673), .X(n12245) );
  nand_x1_sg U55643 ( .A(n12246), .B(n12247), .X(n12244) );
  nand_x1_sg U55644 ( .A(n48970), .B(n48959), .X(n13064) );
  nand_x1_sg U55645 ( .A(n13065), .B(n13066), .X(n13063) );
  nand_x1_sg U55646 ( .A(n49257), .B(n49246), .X(n13883) );
  nand_x1_sg U55647 ( .A(n13884), .B(n13885), .X(n13882) );
  nand_x1_sg U55648 ( .A(n49543), .B(n49532), .X(n14702) );
  nand_x1_sg U55649 ( .A(n14703), .B(n14704), .X(n14701) );
  nand_x1_sg U55650 ( .A(n49829), .B(n49818), .X(n15521) );
  nand_x1_sg U55651 ( .A(n15522), .B(n15523), .X(n15520) );
  nand_x1_sg U55652 ( .A(n50115), .B(n50104), .X(n16340) );
  nand_x1_sg U55653 ( .A(n16341), .B(n16342), .X(n16339) );
  nand_x1_sg U55654 ( .A(n50400), .B(n50389), .X(n17157) );
  nand_x1_sg U55655 ( .A(n17158), .B(n17159), .X(n17156) );
  nand_x1_sg U55656 ( .A(n50689), .B(n50678), .X(n17978) );
  nand_x1_sg U55657 ( .A(n17979), .B(n17980), .X(n17977) );
  nand_x1_sg U55658 ( .A(n50976), .B(n50965), .X(n18799) );
  nand_x1_sg U55659 ( .A(n18800), .B(n18801), .X(n18798) );
  nand_x1_sg U55660 ( .A(n46969), .B(n46957), .X(n7332) );
  nand_x1_sg U55661 ( .A(n7333), .B(n7334), .X(n7331) );
  nand_x1_sg U55662 ( .A(n7358), .B(n47004), .X(n7354) );
  nand_x1_sg U55663 ( .A(n8176), .B(n47293), .X(n8172) );
  nand_x1_sg U55664 ( .A(n8994), .B(n47578), .X(n8990) );
  nand_x1_sg U55665 ( .A(n9814), .B(n47863), .X(n9810) );
  nand_x1_sg U55666 ( .A(n10633), .B(n48148), .X(n10629) );
  nand_x1_sg U55667 ( .A(n11452), .B(n48433), .X(n11448) );
  nand_x1_sg U55668 ( .A(n12271), .B(n48718), .X(n12267) );
  nand_x1_sg U55669 ( .A(n13090), .B(n49004), .X(n13086) );
  nand_x1_sg U55670 ( .A(n13909), .B(n49291), .X(n13905) );
  nand_x1_sg U55671 ( .A(n14728), .B(n49577), .X(n14724) );
  nand_x1_sg U55672 ( .A(n15547), .B(n49863), .X(n15543) );
  nand_x1_sg U55673 ( .A(n16366), .B(n50149), .X(n16362) );
  nand_x1_sg U55674 ( .A(n17183), .B(n50434), .X(n17179) );
  nand_x1_sg U55675 ( .A(n18004), .B(n50723), .X(n18000) );
  nand_x1_sg U55676 ( .A(n18825), .B(n51010), .X(n18821) );
  inv_x1_sg U55677 ( .A(n7044), .X(n47112) );
  inv_x1_sg U55678 ( .A(n7862), .X(n47398) );
  inv_x1_sg U55679 ( .A(n8680), .X(n47683) );
  inv_x1_sg U55680 ( .A(n9500), .X(n47968) );
  inv_x1_sg U55681 ( .A(n10319), .X(n48253) );
  inv_x1_sg U55682 ( .A(n11138), .X(n48538) );
  inv_x1_sg U55683 ( .A(n11957), .X(n48823) );
  inv_x1_sg U55684 ( .A(n12776), .X(n49110) );
  inv_x1_sg U55685 ( .A(n13595), .X(n49396) );
  inv_x1_sg U55686 ( .A(n14414), .X(n49682) );
  inv_x1_sg U55687 ( .A(n15233), .X(n49968) );
  inv_x1_sg U55688 ( .A(n16052), .X(n50254) );
  inv_x1_sg U55689 ( .A(n16871), .X(n50539) );
  inv_x1_sg U55690 ( .A(n17690), .X(n50828) );
  inv_x1_sg U55691 ( .A(n18511), .X(n51115) );
  nand_x1_sg U55692 ( .A(n47067), .B(n7404), .X(n7410) );
  inv_x1_sg U55693 ( .A(n7403), .X(n47067) );
  nand_x1_sg U55694 ( .A(n47353), .B(n8222), .X(n8228) );
  inv_x1_sg U55695 ( .A(n8221), .X(n47353) );
  nand_x1_sg U55696 ( .A(n47638), .B(n9040), .X(n9046) );
  inv_x1_sg U55697 ( .A(n9039), .X(n47638) );
  nand_x1_sg U55698 ( .A(n47923), .B(n9860), .X(n9866) );
  inv_x1_sg U55699 ( .A(n9859), .X(n47923) );
  nand_x1_sg U55700 ( .A(n48208), .B(n10679), .X(n10685) );
  inv_x1_sg U55701 ( .A(n10678), .X(n48208) );
  nand_x1_sg U55702 ( .A(n48493), .B(n11498), .X(n11504) );
  inv_x1_sg U55703 ( .A(n11497), .X(n48493) );
  nand_x1_sg U55704 ( .A(n48778), .B(n12317), .X(n12323) );
  inv_x1_sg U55705 ( .A(n12316), .X(n48778) );
  nand_x1_sg U55706 ( .A(n49065), .B(n13136), .X(n13142) );
  inv_x1_sg U55707 ( .A(n13135), .X(n49065) );
  nand_x1_sg U55708 ( .A(n49351), .B(n13955), .X(n13961) );
  inv_x1_sg U55709 ( .A(n13954), .X(n49351) );
  nand_x1_sg U55710 ( .A(n49637), .B(n14774), .X(n14780) );
  inv_x1_sg U55711 ( .A(n14773), .X(n49637) );
  nand_x1_sg U55712 ( .A(n49923), .B(n15593), .X(n15599) );
  inv_x1_sg U55713 ( .A(n15592), .X(n49923) );
  nand_x1_sg U55714 ( .A(n50209), .B(n16412), .X(n16418) );
  inv_x1_sg U55715 ( .A(n16411), .X(n50209) );
  nand_x1_sg U55716 ( .A(n50494), .B(n17229), .X(n17235) );
  inv_x1_sg U55717 ( .A(n17228), .X(n50494) );
  nand_x1_sg U55718 ( .A(n50783), .B(n18050), .X(n18056) );
  inv_x1_sg U55719 ( .A(n18049), .X(n50783) );
  nand_x1_sg U55720 ( .A(n51070), .B(n18871), .X(n18877) );
  inv_x1_sg U55721 ( .A(n18870), .X(n51070) );
  inv_x1_sg U55722 ( .A(n7453), .X(n47089) );
  inv_x1_sg U55723 ( .A(n8271), .X(n47375) );
  inv_x1_sg U55724 ( .A(n9089), .X(n47660) );
  inv_x1_sg U55725 ( .A(n9909), .X(n47945) );
  inv_x1_sg U55726 ( .A(n10728), .X(n48230) );
  inv_x1_sg U55727 ( .A(n11547), .X(n48515) );
  inv_x1_sg U55728 ( .A(n12366), .X(n48800) );
  inv_x1_sg U55729 ( .A(n13185), .X(n49087) );
  inv_x1_sg U55730 ( .A(n14004), .X(n49373) );
  inv_x1_sg U55731 ( .A(n14823), .X(n49659) );
  inv_x1_sg U55732 ( .A(n15642), .X(n49945) );
  inv_x1_sg U55733 ( .A(n16461), .X(n50231) );
  inv_x1_sg U55734 ( .A(n17278), .X(n50516) );
  inv_x1_sg U55735 ( .A(n18099), .X(n50805) );
  inv_x1_sg U55736 ( .A(n18920), .X(n51092) );
  nor_x1_sg U55737 ( .A(n16707), .B(n16708), .X(n16706) );
  inv_x1_sg U55738 ( .A(n7262), .X(n46999) );
  inv_x1_sg U55739 ( .A(n8081), .X(n47288) );
  inv_x1_sg U55740 ( .A(n8899), .X(n47573) );
  inv_x1_sg U55741 ( .A(n9719), .X(n47858) );
  inv_x1_sg U55742 ( .A(n10538), .X(n48143) );
  inv_x1_sg U55743 ( .A(n11357), .X(n48428) );
  inv_x1_sg U55744 ( .A(n12176), .X(n48713) );
  inv_x1_sg U55745 ( .A(n12995), .X(n48999) );
  inv_x1_sg U55746 ( .A(n13814), .X(n49286) );
  inv_x1_sg U55747 ( .A(n14633), .X(n49572) );
  inv_x1_sg U55748 ( .A(n15452), .X(n49858) );
  inv_x1_sg U55749 ( .A(n16271), .X(n50144) );
  inv_x1_sg U55750 ( .A(n17087), .X(n50429) );
  inv_x1_sg U55751 ( .A(n17909), .X(n50718) );
  inv_x1_sg U55752 ( .A(n18730), .X(n51005) );
  nand_x1_sg U55753 ( .A(n17134), .B(n17133), .X(n17131) );
  nor_x1_sg U55754 ( .A(n17133), .B(n17134), .X(n17132) );
  nor_x1_sg U55755 ( .A(n6935), .B(n6936), .X(n6934) );
  nor_x1_sg U55756 ( .A(n7752), .B(n7753), .X(n7751) );
  nor_x1_sg U55757 ( .A(n8570), .B(n8571), .X(n8569) );
  nor_x1_sg U55758 ( .A(n9390), .B(n9391), .X(n9389) );
  nor_x1_sg U55759 ( .A(n10209), .B(n10210), .X(n10208) );
  nor_x1_sg U55760 ( .A(n11028), .B(n11029), .X(n11027) );
  nor_x1_sg U55761 ( .A(n11847), .B(n11848), .X(n11846) );
  nor_x1_sg U55762 ( .A(n12666), .B(n12667), .X(n12665) );
  nor_x1_sg U55763 ( .A(n13485), .B(n13486), .X(n13484) );
  nor_x1_sg U55764 ( .A(n14304), .B(n14305), .X(n14303) );
  nor_x1_sg U55765 ( .A(n15123), .B(n15124), .X(n15122) );
  nor_x1_sg U55766 ( .A(n15942), .B(n15943), .X(n15941) );
  nor_x1_sg U55767 ( .A(n16759), .B(n16760), .X(n16758) );
  nor_x1_sg U55768 ( .A(n17580), .B(n17581), .X(n17579) );
  nor_x1_sg U55769 ( .A(n18401), .B(n18402), .X(n18400) );
  nand_x1_sg U55770 ( .A(n47250), .B(n47261), .X(n8205) );
  nand_x1_sg U55771 ( .A(n8206), .B(n8207), .X(n8204) );
  nand_x1_sg U55772 ( .A(n47535), .B(n47546), .X(n9023) );
  nand_x1_sg U55773 ( .A(n9024), .B(n9025), .X(n9022) );
  nand_x1_sg U55774 ( .A(n47820), .B(n47831), .X(n9843) );
  nand_x1_sg U55775 ( .A(n9844), .B(n9845), .X(n9842) );
  nand_x1_sg U55776 ( .A(n48105), .B(n48116), .X(n10662) );
  nand_x1_sg U55777 ( .A(n10663), .B(n10664), .X(n10661) );
  nand_x1_sg U55778 ( .A(n48390), .B(n48401), .X(n11481) );
  nand_x1_sg U55779 ( .A(n11482), .B(n11483), .X(n11480) );
  nand_x1_sg U55780 ( .A(n48675), .B(n48686), .X(n12300) );
  nand_x1_sg U55781 ( .A(n12301), .B(n12302), .X(n12299) );
  nand_x1_sg U55782 ( .A(n48961), .B(n48972), .X(n13119) );
  nand_x1_sg U55783 ( .A(n13120), .B(n13121), .X(n13118) );
  nand_x1_sg U55784 ( .A(n49248), .B(n49259), .X(n13938) );
  nand_x1_sg U55785 ( .A(n13939), .B(n13940), .X(n13937) );
  nand_x1_sg U55786 ( .A(n49534), .B(n49545), .X(n14757) );
  nand_x1_sg U55787 ( .A(n14758), .B(n14759), .X(n14756) );
  nand_x1_sg U55788 ( .A(n49820), .B(n49831), .X(n15576) );
  nand_x1_sg U55789 ( .A(n15577), .B(n15578), .X(n15575) );
  nand_x1_sg U55790 ( .A(n50106), .B(n50117), .X(n16395) );
  nand_x1_sg U55791 ( .A(n16396), .B(n16397), .X(n16394) );
  nand_x1_sg U55792 ( .A(n50680), .B(n50691), .X(n18033) );
  nand_x1_sg U55793 ( .A(n18034), .B(n18035), .X(n18032) );
  nand_x1_sg U55794 ( .A(n50967), .B(n50978), .X(n18854) );
  nand_x1_sg U55795 ( .A(n18855), .B(n18856), .X(n18853) );
  nand_x1_sg U55796 ( .A(n46971), .B(n7388), .X(n7385) );
  nand_x1_sg U55797 ( .A(n47261), .B(n8206), .X(n8203) );
  nand_x1_sg U55798 ( .A(n47546), .B(n9024), .X(n9021) );
  nand_x1_sg U55799 ( .A(n47831), .B(n9844), .X(n9841) );
  nand_x1_sg U55800 ( .A(n48116), .B(n10663), .X(n10660) );
  nand_x1_sg U55801 ( .A(n48401), .B(n11482), .X(n11479) );
  nand_x1_sg U55802 ( .A(n48686), .B(n12301), .X(n12298) );
  nand_x1_sg U55803 ( .A(n48972), .B(n13120), .X(n13117) );
  nand_x1_sg U55804 ( .A(n49259), .B(n13939), .X(n13936) );
  nand_x1_sg U55805 ( .A(n49545), .B(n14758), .X(n14755) );
  nand_x1_sg U55806 ( .A(n49831), .B(n15577), .X(n15574) );
  nand_x1_sg U55807 ( .A(n50117), .B(n16396), .X(n16393) );
  nand_x1_sg U55808 ( .A(n50402), .B(n17213), .X(n17210) );
  nand_x1_sg U55809 ( .A(n50691), .B(n18034), .X(n18031) );
  nand_x1_sg U55810 ( .A(n50978), .B(n18855), .X(n18852) );
  nand_x1_sg U55811 ( .A(n7120), .B(n7119), .X(n7117) );
  nor_x1_sg U55812 ( .A(n7119), .B(n7120), .X(n7118) );
  nand_x1_sg U55813 ( .A(n7938), .B(n7937), .X(n7935) );
  nor_x1_sg U55814 ( .A(n7937), .B(n7938), .X(n7936) );
  nand_x1_sg U55815 ( .A(n8756), .B(n8755), .X(n8753) );
  nor_x1_sg U55816 ( .A(n8755), .B(n8756), .X(n8754) );
  nand_x1_sg U55817 ( .A(n9576), .B(n9575), .X(n9573) );
  nor_x1_sg U55818 ( .A(n9575), .B(n9576), .X(n9574) );
  nand_x1_sg U55819 ( .A(n10395), .B(n10394), .X(n10392) );
  nor_x1_sg U55820 ( .A(n10394), .B(n10395), .X(n10393) );
  nand_x1_sg U55821 ( .A(n11214), .B(n11213), .X(n11211) );
  nor_x1_sg U55822 ( .A(n11213), .B(n11214), .X(n11212) );
  nand_x1_sg U55823 ( .A(n12033), .B(n12032), .X(n12030) );
  nor_x1_sg U55824 ( .A(n12032), .B(n12033), .X(n12031) );
  nand_x1_sg U55825 ( .A(n12852), .B(n12851), .X(n12849) );
  nor_x1_sg U55826 ( .A(n12851), .B(n12852), .X(n12850) );
  nand_x1_sg U55827 ( .A(n13671), .B(n13670), .X(n13668) );
  nor_x1_sg U55828 ( .A(n13670), .B(n13671), .X(n13669) );
  nand_x1_sg U55829 ( .A(n14490), .B(n14489), .X(n14487) );
  nor_x1_sg U55830 ( .A(n14489), .B(n14490), .X(n14488) );
  nand_x1_sg U55831 ( .A(n15309), .B(n15308), .X(n15306) );
  nor_x1_sg U55832 ( .A(n15308), .B(n15309), .X(n15307) );
  nand_x1_sg U55833 ( .A(n16128), .B(n16127), .X(n16125) );
  nor_x1_sg U55834 ( .A(n16127), .B(n16128), .X(n16126) );
  nand_x1_sg U55835 ( .A(n16945), .B(n16944), .X(n16942) );
  nor_x1_sg U55836 ( .A(n16944), .B(n16945), .X(n16943) );
  nand_x1_sg U55837 ( .A(n17766), .B(n17765), .X(n17763) );
  nor_x1_sg U55838 ( .A(n17765), .B(n17766), .X(n17764) );
  nand_x1_sg U55839 ( .A(n18587), .B(n18586), .X(n18584) );
  nor_x1_sg U55840 ( .A(n18586), .B(n18587), .X(n18585) );
  nand_x1_sg U55841 ( .A(n7044), .B(n7043), .X(n7514) );
  nor_x1_sg U55842 ( .A(n7043), .B(n7044), .X(n7515) );
  nand_x1_sg U55843 ( .A(n7862), .B(n7861), .X(n8332) );
  nor_x1_sg U55844 ( .A(n7861), .B(n7862), .X(n8333) );
  nand_x1_sg U55845 ( .A(n8680), .B(n8679), .X(n9150) );
  nor_x1_sg U55846 ( .A(n8679), .B(n8680), .X(n9151) );
  nand_x1_sg U55847 ( .A(n9500), .B(n9499), .X(n9970) );
  nor_x1_sg U55848 ( .A(n9499), .B(n9500), .X(n9971) );
  nand_x1_sg U55849 ( .A(n10319), .B(n10318), .X(n10789) );
  nor_x1_sg U55850 ( .A(n10318), .B(n10319), .X(n10790) );
  nand_x1_sg U55851 ( .A(n11138), .B(n11137), .X(n11608) );
  nor_x1_sg U55852 ( .A(n11137), .B(n11138), .X(n11609) );
  nand_x1_sg U55853 ( .A(n11957), .B(n11956), .X(n12427) );
  nor_x1_sg U55854 ( .A(n11956), .B(n11957), .X(n12428) );
  nand_x1_sg U55855 ( .A(n12776), .B(n12775), .X(n13246) );
  nor_x1_sg U55856 ( .A(n12775), .B(n12776), .X(n13247) );
  nand_x1_sg U55857 ( .A(n13595), .B(n13594), .X(n14065) );
  nor_x1_sg U55858 ( .A(n13594), .B(n13595), .X(n14066) );
  nand_x1_sg U55859 ( .A(n14414), .B(n14413), .X(n14884) );
  nor_x1_sg U55860 ( .A(n14413), .B(n14414), .X(n14885) );
  nand_x1_sg U55861 ( .A(n15233), .B(n15232), .X(n15703) );
  nor_x1_sg U55862 ( .A(n15232), .B(n15233), .X(n15704) );
  nand_x1_sg U55863 ( .A(n16052), .B(n16051), .X(n16522) );
  nor_x1_sg U55864 ( .A(n16051), .B(n16052), .X(n16523) );
  nand_x1_sg U55865 ( .A(n16871), .B(n16870), .X(n17339) );
  nor_x1_sg U55866 ( .A(n16870), .B(n16871), .X(n17340) );
  nand_x1_sg U55867 ( .A(n17690), .B(n17689), .X(n18160) );
  nor_x1_sg U55868 ( .A(n17689), .B(n17690), .X(n18161) );
  nand_x1_sg U55869 ( .A(n18511), .B(n18510), .X(n18981) );
  nor_x1_sg U55870 ( .A(n18510), .B(n18511), .X(n18982) );
  nand_x1_sg U55871 ( .A(n8271), .B(n8270), .X(n8268) );
  nor_x1_sg U55872 ( .A(n8270), .B(n8271), .X(n8269) );
  nand_x1_sg U55873 ( .A(n9089), .B(n9088), .X(n9086) );
  nor_x1_sg U55874 ( .A(n9088), .B(n9089), .X(n9087) );
  nand_x1_sg U55875 ( .A(n9909), .B(n9908), .X(n9906) );
  nor_x1_sg U55876 ( .A(n9908), .B(n9909), .X(n9907) );
  nand_x1_sg U55877 ( .A(n10728), .B(n10727), .X(n10725) );
  nor_x1_sg U55878 ( .A(n10727), .B(n10728), .X(n10726) );
  nand_x1_sg U55879 ( .A(n11547), .B(n11546), .X(n11544) );
  nor_x1_sg U55880 ( .A(n11546), .B(n11547), .X(n11545) );
  nand_x1_sg U55881 ( .A(n12366), .B(n12365), .X(n12363) );
  nor_x1_sg U55882 ( .A(n12365), .B(n12366), .X(n12364) );
  nand_x1_sg U55883 ( .A(n13185), .B(n13184), .X(n13182) );
  nor_x1_sg U55884 ( .A(n13184), .B(n13185), .X(n13183) );
  nand_x1_sg U55885 ( .A(n14004), .B(n14003), .X(n14001) );
  nor_x1_sg U55886 ( .A(n14003), .B(n14004), .X(n14002) );
  nand_x1_sg U55887 ( .A(n14823), .B(n14822), .X(n14820) );
  nor_x1_sg U55888 ( .A(n14822), .B(n14823), .X(n14821) );
  nand_x1_sg U55889 ( .A(n15642), .B(n15641), .X(n15639) );
  nor_x1_sg U55890 ( .A(n15641), .B(n15642), .X(n15640) );
  nand_x1_sg U55891 ( .A(n16461), .B(n16460), .X(n16458) );
  nor_x1_sg U55892 ( .A(n16460), .B(n16461), .X(n16459) );
  nand_x1_sg U55893 ( .A(n17278), .B(n17277), .X(n17275) );
  nor_x1_sg U55894 ( .A(n17277), .B(n17278), .X(n17276) );
  nand_x1_sg U55895 ( .A(n18099), .B(n18098), .X(n18096) );
  nor_x1_sg U55896 ( .A(n18098), .B(n18099), .X(n18097) );
  nand_x1_sg U55897 ( .A(n18920), .B(n18919), .X(n18917) );
  nor_x1_sg U55898 ( .A(n18919), .B(n18920), .X(n18918) );
  nand_x1_sg U55899 ( .A(n7453), .B(n7452), .X(n7450) );
  nor_x1_sg U55900 ( .A(n7452), .B(n7453), .X(n7451) );
  nand_x1_sg U55901 ( .A(n7262), .B(n42255), .X(n7259) );
  nor_x1_sg U55902 ( .A(n42255), .B(n7262), .X(n7260) );
  nand_x1_sg U55903 ( .A(n8081), .B(n8080), .X(n8078) );
  nor_x1_sg U55904 ( .A(n8080), .B(n8081), .X(n8079) );
  nand_x1_sg U55905 ( .A(n8899), .B(n8898), .X(n8896) );
  nor_x1_sg U55906 ( .A(n8898), .B(n8899), .X(n8897) );
  nand_x1_sg U55907 ( .A(n9719), .B(n9718), .X(n9716) );
  nor_x1_sg U55908 ( .A(n9718), .B(n9719), .X(n9717) );
  nand_x1_sg U55909 ( .A(n10538), .B(n10537), .X(n10535) );
  nor_x1_sg U55910 ( .A(n10537), .B(n10538), .X(n10536) );
  nand_x1_sg U55911 ( .A(n11357), .B(n11356), .X(n11354) );
  nor_x1_sg U55912 ( .A(n11356), .B(n11357), .X(n11355) );
  nand_x1_sg U55913 ( .A(n12176), .B(n12175), .X(n12173) );
  nor_x1_sg U55914 ( .A(n12175), .B(n12176), .X(n12174) );
  nand_x1_sg U55915 ( .A(n12995), .B(n12994), .X(n12992) );
  nor_x1_sg U55916 ( .A(n12994), .B(n12995), .X(n12993) );
  nand_x1_sg U55917 ( .A(n13814), .B(n13813), .X(n13811) );
  nor_x1_sg U55918 ( .A(n13813), .B(n13814), .X(n13812) );
  nand_x1_sg U55919 ( .A(n14633), .B(n14632), .X(n14630) );
  nor_x1_sg U55920 ( .A(n14632), .B(n14633), .X(n14631) );
  nand_x1_sg U55921 ( .A(n15452), .B(n15451), .X(n15449) );
  nor_x1_sg U55922 ( .A(n15451), .B(n15452), .X(n15450) );
  nand_x1_sg U55923 ( .A(n16271), .B(n16270), .X(n16268) );
  nor_x1_sg U55924 ( .A(n16270), .B(n16271), .X(n16269) );
  nand_x1_sg U55925 ( .A(n17087), .B(n42242), .X(n17084) );
  nor_x1_sg U55926 ( .A(n42242), .B(n17087), .X(n17085) );
  nand_x1_sg U55927 ( .A(n17909), .B(n17908), .X(n17906) );
  nor_x1_sg U55928 ( .A(n17908), .B(n17909), .X(n17907) );
  nand_x1_sg U55929 ( .A(n18730), .B(n18729), .X(n18727) );
  nor_x1_sg U55930 ( .A(n18729), .B(n18730), .X(n18728) );
  nand_x1_sg U55931 ( .A(n17226), .B(n50449), .X(n17223) );
  nand_x1_sg U55932 ( .A(n17225), .B(n50465), .X(n17224) );
  nand_x1_sg U55933 ( .A(n7034), .B(n47082), .X(n7567) );
  nor_x1_sg U55934 ( .A(n47082), .B(n7034), .X(n7568) );
  nand_x1_sg U55935 ( .A(n7852), .B(n47368), .X(n8385) );
  nor_x1_sg U55936 ( .A(n47368), .B(n7852), .X(n8386) );
  nand_x1_sg U55937 ( .A(n8670), .B(n47653), .X(n9203) );
  nor_x1_sg U55938 ( .A(n47653), .B(n8670), .X(n9204) );
  nand_x1_sg U55939 ( .A(n9490), .B(n47938), .X(n10023) );
  nor_x1_sg U55940 ( .A(n47938), .B(n9490), .X(n10024) );
  nand_x1_sg U55941 ( .A(n10309), .B(n48223), .X(n10842) );
  nor_x1_sg U55942 ( .A(n48223), .B(n10309), .X(n10843) );
  nand_x1_sg U55943 ( .A(n11128), .B(n48508), .X(n11661) );
  nor_x1_sg U55944 ( .A(n48508), .B(n11128), .X(n11662) );
  nand_x1_sg U55945 ( .A(n11947), .B(n48793), .X(n12480) );
  nor_x1_sg U55946 ( .A(n48793), .B(n11947), .X(n12481) );
  nand_x1_sg U55947 ( .A(n12766), .B(n49080), .X(n13299) );
  nor_x1_sg U55948 ( .A(n49080), .B(n12766), .X(n13300) );
  nand_x1_sg U55949 ( .A(n13585), .B(n49366), .X(n14118) );
  nor_x1_sg U55950 ( .A(n49366), .B(n13585), .X(n14119) );
  nand_x1_sg U55951 ( .A(n14404), .B(n49652), .X(n14937) );
  nor_x1_sg U55952 ( .A(n49652), .B(n14404), .X(n14938) );
  nand_x1_sg U55953 ( .A(n15223), .B(n49938), .X(n15756) );
  nor_x1_sg U55954 ( .A(n49938), .B(n15223), .X(n15757) );
  nand_x1_sg U55955 ( .A(n16042), .B(n50224), .X(n16575) );
  nor_x1_sg U55956 ( .A(n50224), .B(n16042), .X(n16576) );
  nand_x1_sg U55957 ( .A(n16861), .B(n50509), .X(n17392) );
  nor_x1_sg U55958 ( .A(n50509), .B(n16861), .X(n17393) );
  nand_x1_sg U55959 ( .A(n17680), .B(n50798), .X(n18213) );
  nor_x1_sg U55960 ( .A(n50798), .B(n17680), .X(n18214) );
  nand_x1_sg U55961 ( .A(n18501), .B(n51085), .X(n19034) );
  nor_x1_sg U55962 ( .A(n51085), .B(n18501), .X(n19035) );
  inv_x1_sg U55963 ( .A(n22656), .X(n46938) );
  nand_x1_sg U55964 ( .A(n7403), .B(n7404), .X(n7402) );
  nor_x1_sg U55965 ( .A(n7404), .B(n7403), .X(n7405) );
  nand_x1_sg U55966 ( .A(n8221), .B(n8222), .X(n8220) );
  nor_x1_sg U55967 ( .A(n8222), .B(n8221), .X(n8223) );
  nand_x1_sg U55968 ( .A(n9039), .B(n9040), .X(n9038) );
  nor_x1_sg U55969 ( .A(n9040), .B(n9039), .X(n9041) );
  nand_x1_sg U55970 ( .A(n9859), .B(n9860), .X(n9858) );
  nor_x1_sg U55971 ( .A(n9860), .B(n9859), .X(n9861) );
  nand_x1_sg U55972 ( .A(n10678), .B(n10679), .X(n10677) );
  nor_x1_sg U55973 ( .A(n10679), .B(n10678), .X(n10680) );
  nand_x1_sg U55974 ( .A(n11497), .B(n11498), .X(n11496) );
  nor_x1_sg U55975 ( .A(n11498), .B(n11497), .X(n11499) );
  nand_x1_sg U55976 ( .A(n12316), .B(n12317), .X(n12315) );
  nor_x1_sg U55977 ( .A(n12317), .B(n12316), .X(n12318) );
  nand_x1_sg U55978 ( .A(n13135), .B(n13136), .X(n13134) );
  nor_x1_sg U55979 ( .A(n13136), .B(n13135), .X(n13137) );
  nand_x1_sg U55980 ( .A(n13954), .B(n13955), .X(n13953) );
  nor_x1_sg U55981 ( .A(n13955), .B(n13954), .X(n13956) );
  nand_x1_sg U55982 ( .A(n14773), .B(n14774), .X(n14772) );
  nor_x1_sg U55983 ( .A(n14774), .B(n14773), .X(n14775) );
  nand_x1_sg U55984 ( .A(n15592), .B(n15593), .X(n15591) );
  nor_x1_sg U55985 ( .A(n15593), .B(n15592), .X(n15594) );
  nand_x1_sg U55986 ( .A(n16411), .B(n16412), .X(n16410) );
  nor_x1_sg U55987 ( .A(n16412), .B(n16411), .X(n16413) );
  nand_x1_sg U55988 ( .A(n17228), .B(n17229), .X(n17227) );
  nor_x1_sg U55989 ( .A(n17229), .B(n17228), .X(n17230) );
  nand_x1_sg U55990 ( .A(n18049), .B(n18050), .X(n18048) );
  nor_x1_sg U55991 ( .A(n18050), .B(n18049), .X(n18051) );
  nand_x1_sg U55992 ( .A(n18870), .B(n18871), .X(n18869) );
  nor_x1_sg U55993 ( .A(n18871), .B(n18870), .X(n18872) );
  nand_x1_sg U55994 ( .A(n7017), .B(n7018), .X(n7016) );
  nor_x1_sg U55995 ( .A(n7018), .B(n7017), .X(n7019) );
  nand_x1_sg U55996 ( .A(n7835), .B(n7836), .X(n7834) );
  nor_x1_sg U55997 ( .A(n7836), .B(n7835), .X(n7837) );
  nand_x1_sg U55998 ( .A(n8653), .B(n8654), .X(n8652) );
  nor_x1_sg U55999 ( .A(n8654), .B(n8653), .X(n8655) );
  nand_x1_sg U56000 ( .A(n9473), .B(n9474), .X(n9472) );
  nor_x1_sg U56001 ( .A(n9474), .B(n9473), .X(n9475) );
  nand_x1_sg U56002 ( .A(n10292), .B(n10293), .X(n10291) );
  nor_x1_sg U56003 ( .A(n10293), .B(n10292), .X(n10294) );
  nand_x1_sg U56004 ( .A(n11111), .B(n11112), .X(n11110) );
  nor_x1_sg U56005 ( .A(n11112), .B(n11111), .X(n11113) );
  nand_x1_sg U56006 ( .A(n11930), .B(n11931), .X(n11929) );
  nor_x1_sg U56007 ( .A(n11931), .B(n11930), .X(n11932) );
  nand_x1_sg U56008 ( .A(n12749), .B(n12750), .X(n12748) );
  nor_x1_sg U56009 ( .A(n12750), .B(n12749), .X(n12751) );
  nand_x1_sg U56010 ( .A(n13568), .B(n13569), .X(n13567) );
  nor_x1_sg U56011 ( .A(n13569), .B(n13568), .X(n13570) );
  nand_x1_sg U56012 ( .A(n14387), .B(n14388), .X(n14386) );
  nor_x1_sg U56013 ( .A(n14388), .B(n14387), .X(n14389) );
  nand_x1_sg U56014 ( .A(n15206), .B(n15207), .X(n15205) );
  nor_x1_sg U56015 ( .A(n15207), .B(n15206), .X(n15208) );
  nand_x1_sg U56016 ( .A(n16025), .B(n16026), .X(n16024) );
  nor_x1_sg U56017 ( .A(n16026), .B(n16025), .X(n16027) );
  nand_x1_sg U56018 ( .A(n17663), .B(n17664), .X(n17662) );
  nor_x1_sg U56019 ( .A(n17664), .B(n17663), .X(n17665) );
  nand_x1_sg U56020 ( .A(n18484), .B(n18485), .X(n18483) );
  nor_x1_sg U56021 ( .A(n18485), .B(n18484), .X(n18486) );
  nand_x1_sg U56022 ( .A(n47009), .B(n6952), .X(n6951) );
  nor_x1_sg U56023 ( .A(n6952), .B(n47009), .X(n6953) );
  nand_x1_sg U56024 ( .A(n50438), .B(n16776), .X(n16775) );
  nor_x1_sg U56025 ( .A(n16776), .B(n50438), .X(n16777) );
  nor_x1_sg U56026 ( .A(n38892), .B(n6842), .X(\L2_0/n3512 ) );
  nor_x1_sg U56027 ( .A(n6822), .B(n6879), .X(\L2_0/n3488 ) );
  inv_x1_sg U56028 ( .A(n22980), .X(n47385) );
  inv_x1_sg U56029 ( .A(n23257), .X(n47670) );
  inv_x1_sg U56030 ( .A(n23537), .X(n47955) );
  inv_x1_sg U56031 ( .A(n23816), .X(n48240) );
  inv_x1_sg U56032 ( .A(n24095), .X(n48525) );
  inv_x1_sg U56033 ( .A(n24374), .X(n48810) );
  inv_x1_sg U56034 ( .A(n24653), .X(n49097) );
  inv_x1_sg U56035 ( .A(n24931), .X(n49383) );
  inv_x1_sg U56036 ( .A(n25210), .X(n49669) );
  inv_x1_sg U56037 ( .A(n25489), .X(n49955) );
  inv_x1_sg U56038 ( .A(n25768), .X(n50241) );
  inv_x1_sg U56039 ( .A(n26324), .X(n50815) );
  inv_x1_sg U56040 ( .A(n26605), .X(n51102) );
  inv_x1_sg U56041 ( .A(n8207), .X(n47261) );
  inv_x1_sg U56042 ( .A(n9025), .X(n47546) );
  inv_x1_sg U56043 ( .A(n9845), .X(n47831) );
  inv_x1_sg U56044 ( .A(n10664), .X(n48116) );
  inv_x1_sg U56045 ( .A(n11483), .X(n48401) );
  inv_x1_sg U56046 ( .A(n12302), .X(n48686) );
  inv_x1_sg U56047 ( .A(n13121), .X(n48972) );
  inv_x1_sg U56048 ( .A(n13940), .X(n49259) );
  inv_x1_sg U56049 ( .A(n14759), .X(n49545) );
  inv_x1_sg U56050 ( .A(n15578), .X(n49831) );
  inv_x1_sg U56051 ( .A(n16397), .X(n50117) );
  inv_x1_sg U56052 ( .A(n18035), .X(n50691) );
  inv_x1_sg U56053 ( .A(n18856), .X(n50978) );
  inv_x1_sg U56054 ( .A(n8152), .X(n47248) );
  inv_x1_sg U56055 ( .A(n8970), .X(n47533) );
  inv_x1_sg U56056 ( .A(n9790), .X(n47818) );
  inv_x1_sg U56057 ( .A(n10609), .X(n48103) );
  inv_x1_sg U56058 ( .A(n11428), .X(n48388) );
  inv_x1_sg U56059 ( .A(n12247), .X(n48673) );
  inv_x1_sg U56060 ( .A(n13066), .X(n48959) );
  inv_x1_sg U56061 ( .A(n13885), .X(n49246) );
  inv_x1_sg U56062 ( .A(n14704), .X(n49532) );
  inv_x1_sg U56063 ( .A(n15523), .X(n49818) );
  inv_x1_sg U56064 ( .A(n16342), .X(n50104) );
  inv_x1_sg U56065 ( .A(n17159), .X(n50389) );
  inv_x1_sg U56066 ( .A(n17980), .X(n50678) );
  inv_x1_sg U56067 ( .A(n18801), .X(n50965) );
  inv_x1_sg U56068 ( .A(n7334), .X(n46957) );
  inv_x1_sg U56069 ( .A(n7170), .X(n46929) );
  inv_x1_sg U56070 ( .A(n7989), .X(n47221) );
  inv_x1_sg U56071 ( .A(n8807), .X(n47506) );
  inv_x1_sg U56072 ( .A(n9627), .X(n47791) );
  inv_x1_sg U56073 ( .A(n10446), .X(n48076) );
  inv_x1_sg U56074 ( .A(n11265), .X(n48361) );
  inv_x1_sg U56075 ( .A(n12084), .X(n48646) );
  inv_x1_sg U56076 ( .A(n12903), .X(n48932) );
  inv_x1_sg U56077 ( .A(n13722), .X(n49219) );
  inv_x1_sg U56078 ( .A(n14541), .X(n49505) );
  inv_x1_sg U56079 ( .A(n15360), .X(n49791) );
  inv_x1_sg U56080 ( .A(n16179), .X(n50077) );
  inv_x1_sg U56081 ( .A(n16995), .X(n50362) );
  inv_x1_sg U56082 ( .A(n17817), .X(n50651) );
  inv_x1_sg U56083 ( .A(n18638), .X(n50938) );
  nor_x1_sg U56084 ( .A(n22905), .B(n39900), .X(\L1_0/n4323 ) );
  nor_x1_sg U56085 ( .A(n6835), .B(n40923), .X(\L2_0/n3516 ) );
  nor_x1_sg U56086 ( .A(n6927), .B(n40922), .X(\L2_0/n3456 ) );
  inv_x1_sg U56087 ( .A(n7210), .X(n46916) );
  nor_x1_sg U56088 ( .A(n6849), .B(n6822), .X(\L2_0/n3508 ) );
  nor_x1_sg U56089 ( .A(n6855), .B(n40923), .X(\L2_0/n3504 ) );
  nor_x1_sg U56090 ( .A(n6873), .B(n40921), .X(\L2_0/n3492 ) );
  nor_x1_sg U56091 ( .A(n6885), .B(n40921), .X(\L2_0/n3484 ) );
  nor_x1_sg U56092 ( .A(n6891), .B(n40921), .X(\L2_0/n3480 ) );
  nor_x1_sg U56093 ( .A(n6897), .B(n40922), .X(\L2_0/n3476 ) );
  nor_x1_sg U56094 ( .A(n6903), .B(n40923), .X(\L2_0/n3472 ) );
  nor_x1_sg U56095 ( .A(n6909), .B(n40923), .X(\L2_0/n3468 ) );
  nor_x1_sg U56096 ( .A(n6915), .B(n40921), .X(\L2_0/n3464 ) );
  nor_x1_sg U56097 ( .A(n6921), .B(n40922), .X(\L2_0/n3460 ) );
  nor_x1_sg U56098 ( .A(n40029), .B(n51325), .X(\L1_0/n4324 ) );
  inv_x1_sg U56099 ( .A(n22905), .X(n51325) );
  nor_x1_sg U56100 ( .A(n39142), .B(n22912), .X(\L1_0/n4320 ) );
  nor_x1_sg U56101 ( .A(n41386), .B(n22940), .X(\L1_0/n4304 ) );
  nor_x1_sg U56102 ( .A(n42000), .B(n22954), .X(\L1_0/n4296 ) );
  nor_x1_sg U56103 ( .A(n39143), .B(n22926), .X(\L1_0/n4312 ) );
  nor_x1_sg U56104 ( .A(n51209), .B(n42000), .X(\L1_0/n4311 ) );
  inv_x1_sg U56105 ( .A(n22926), .X(n51209) );
  nor_x1_sg U56106 ( .A(n51208), .B(n40029), .X(\L1_0/n4319 ) );
  inv_x1_sg U56107 ( .A(n22912), .X(n51208) );
  nor_x1_sg U56108 ( .A(n51210), .B(n41388), .X(\L1_0/n4303 ) );
  inv_x1_sg U56109 ( .A(n22940), .X(n51210) );
  nor_x1_sg U56110 ( .A(n51211), .B(n41387), .X(\L1_0/n4295 ) );
  inv_x1_sg U56111 ( .A(n22954), .X(n51211) );
  nand_x1_sg U56112 ( .A(n40585), .B(n40023), .X(n6823) );
  nor_x1_sg U56113 ( .A(n7210), .B(n7211), .X(n7208) );
  nand_x1_sg U56114 ( .A(n7210), .B(n7211), .X(n7209) );
  nor_x1_sg U56115 ( .A(n8029), .B(n8030), .X(n8027) );
  nand_x1_sg U56116 ( .A(n8029), .B(n8030), .X(n8028) );
  nor_x1_sg U56117 ( .A(n8847), .B(n8848), .X(n8845) );
  nand_x1_sg U56118 ( .A(n8847), .B(n8848), .X(n8846) );
  nor_x1_sg U56119 ( .A(n9667), .B(n9668), .X(n9665) );
  nand_x1_sg U56120 ( .A(n9667), .B(n9668), .X(n9666) );
  nor_x1_sg U56121 ( .A(n10486), .B(n10487), .X(n10484) );
  nand_x1_sg U56122 ( .A(n10486), .B(n10487), .X(n10485) );
  nor_x1_sg U56123 ( .A(n11305), .B(n11306), .X(n11303) );
  nand_x1_sg U56124 ( .A(n11305), .B(n11306), .X(n11304) );
  nor_x1_sg U56125 ( .A(n12124), .B(n12125), .X(n12122) );
  nand_x1_sg U56126 ( .A(n12124), .B(n12125), .X(n12123) );
  nor_x1_sg U56127 ( .A(n12943), .B(n12944), .X(n12941) );
  nand_x1_sg U56128 ( .A(n12943), .B(n12944), .X(n12942) );
  nor_x1_sg U56129 ( .A(n13762), .B(n13763), .X(n13760) );
  nand_x1_sg U56130 ( .A(n13762), .B(n13763), .X(n13761) );
  nor_x1_sg U56131 ( .A(n14581), .B(n14582), .X(n14579) );
  nand_x1_sg U56132 ( .A(n14581), .B(n14582), .X(n14580) );
  nor_x1_sg U56133 ( .A(n15400), .B(n15401), .X(n15398) );
  nand_x1_sg U56134 ( .A(n15400), .B(n15401), .X(n15399) );
  nor_x1_sg U56135 ( .A(n16219), .B(n16220), .X(n16217) );
  nand_x1_sg U56136 ( .A(n16219), .B(n16220), .X(n16218) );
  nor_x1_sg U56137 ( .A(n17035), .B(n17036), .X(n17033) );
  nand_x1_sg U56138 ( .A(n17035), .B(n17036), .X(n17034) );
  nor_x1_sg U56139 ( .A(n17857), .B(n17858), .X(n17855) );
  nand_x1_sg U56140 ( .A(n17857), .B(n17858), .X(n17856) );
  nor_x1_sg U56141 ( .A(n18678), .B(n18679), .X(n18676) );
  nand_x1_sg U56142 ( .A(n18678), .B(n18679), .X(n18677) );
  nor_x1_sg U56143 ( .A(n7215), .B(n7214), .X(n7212) );
  nand_x1_sg U56144 ( .A(n7214), .B(n7215), .X(n7213) );
  nor_x1_sg U56145 ( .A(n50423), .B(n50347), .X(n17152) );
  nor_x1_sg U56146 ( .A(n17154), .B(n17155), .X(n17153) );
  inv_x1_sg U56147 ( .A(n17154), .X(n50347) );
  nor_x1_sg U56148 ( .A(n39680), .B(n39603), .X(n17377) );
  nor_x1_sg U56149 ( .A(n7242), .B(n46976), .X(n7233) );
  inv_x1_sg U56150 ( .A(n7243), .X(n46976) );
  nor_x1_sg U56151 ( .A(n7244), .B(n7245), .X(n7242) );
  nor_x1_sg U56152 ( .A(n8061), .B(n47266), .X(n8052) );
  inv_x1_sg U56153 ( .A(n8062), .X(n47266) );
  nor_x1_sg U56154 ( .A(n8063), .B(n8064), .X(n8061) );
  nor_x1_sg U56155 ( .A(n8879), .B(n47551), .X(n8870) );
  inv_x1_sg U56156 ( .A(n8880), .X(n47551) );
  nor_x1_sg U56157 ( .A(n8881), .B(n8882), .X(n8879) );
  nor_x1_sg U56158 ( .A(n9699), .B(n47836), .X(n9690) );
  inv_x1_sg U56159 ( .A(n9700), .X(n47836) );
  nor_x1_sg U56160 ( .A(n9701), .B(n9702), .X(n9699) );
  nor_x1_sg U56161 ( .A(n10518), .B(n48121), .X(n10509) );
  inv_x1_sg U56162 ( .A(n10519), .X(n48121) );
  nor_x1_sg U56163 ( .A(n10520), .B(n10521), .X(n10518) );
  nor_x1_sg U56164 ( .A(n11337), .B(n48406), .X(n11328) );
  inv_x1_sg U56165 ( .A(n11338), .X(n48406) );
  nor_x1_sg U56166 ( .A(n11339), .B(n11340), .X(n11337) );
  nor_x1_sg U56167 ( .A(n12156), .B(n48691), .X(n12147) );
  inv_x1_sg U56168 ( .A(n12157), .X(n48691) );
  nor_x1_sg U56169 ( .A(n12158), .B(n12159), .X(n12156) );
  nor_x1_sg U56170 ( .A(n12975), .B(n48977), .X(n12966) );
  inv_x1_sg U56171 ( .A(n12976), .X(n48977) );
  nor_x1_sg U56172 ( .A(n12977), .B(n12978), .X(n12975) );
  nor_x1_sg U56173 ( .A(n13794), .B(n49264), .X(n13785) );
  inv_x1_sg U56174 ( .A(n13795), .X(n49264) );
  nor_x1_sg U56175 ( .A(n13796), .B(n13797), .X(n13794) );
  nor_x1_sg U56176 ( .A(n14613), .B(n49550), .X(n14604) );
  inv_x1_sg U56177 ( .A(n14614), .X(n49550) );
  nor_x1_sg U56178 ( .A(n14615), .B(n14616), .X(n14613) );
  nor_x1_sg U56179 ( .A(n15432), .B(n49836), .X(n15423) );
  inv_x1_sg U56180 ( .A(n15433), .X(n49836) );
  nor_x1_sg U56181 ( .A(n15434), .B(n15435), .X(n15432) );
  nor_x1_sg U56182 ( .A(n16251), .B(n50122), .X(n16242) );
  inv_x1_sg U56183 ( .A(n16252), .X(n50122) );
  nor_x1_sg U56184 ( .A(n16253), .B(n16254), .X(n16251) );
  nor_x1_sg U56185 ( .A(n17067), .B(n50407), .X(n17058) );
  inv_x1_sg U56186 ( .A(n17068), .X(n50407) );
  nor_x1_sg U56187 ( .A(n17069), .B(n17070), .X(n17067) );
  nor_x1_sg U56188 ( .A(n17889), .B(n50696), .X(n17880) );
  inv_x1_sg U56189 ( .A(n17890), .X(n50696) );
  nor_x1_sg U56190 ( .A(n17891), .B(n17892), .X(n17889) );
  nor_x1_sg U56191 ( .A(n18710), .B(n50983), .X(n18701) );
  inv_x1_sg U56192 ( .A(n18711), .X(n50983) );
  nor_x1_sg U56193 ( .A(n18712), .B(n18713), .X(n18710) );
  nor_x1_sg U56194 ( .A(n39606), .B(n39855), .X(n6958) );
  nor_x1_sg U56195 ( .A(n39602), .B(n39884), .X(n16782) );
  nor_x1_sg U56196 ( .A(n39611), .B(n41736), .X(n8199) );
  nor_x1_sg U56197 ( .A(n39609), .B(n41735), .X(n9017) );
  nor_x1_sg U56198 ( .A(n39627), .B(n41734), .X(n9837) );
  nor_x1_sg U56199 ( .A(n39624), .B(n41727), .X(n10656) );
  nor_x1_sg U56200 ( .A(n39621), .B(n41726), .X(n11475) );
  nor_x1_sg U56201 ( .A(n39618), .B(n41730), .X(n12294) );
  nor_x1_sg U56202 ( .A(n39639), .B(n41729), .X(n13113) );
  nor_x1_sg U56203 ( .A(n39635), .B(n41728), .X(n13932) );
  nor_x1_sg U56204 ( .A(n39633), .B(n41731), .X(n14751) );
  nor_x1_sg U56205 ( .A(n39629), .B(n41733), .X(n15570) );
  nor_x1_sg U56206 ( .A(n39648), .B(n41732), .X(n16389) );
  nor_x1_sg U56207 ( .A(n39615), .B(n41739), .X(n17206) );
  nor_x1_sg U56208 ( .A(n39644), .B(n41738), .X(n18027) );
  nor_x1_sg U56209 ( .A(n39641), .B(n41737), .X(n18848) );
  inv_x1_sg U56210 ( .A(n7121), .X(n46894) );
  nor_x1_sg U56211 ( .A(n7135), .B(n46875), .X(n7134) );
  inv_x1_sg U56212 ( .A(n7939), .X(n47189) );
  nor_x1_sg U56213 ( .A(n7953), .B(n47168), .X(n7952) );
  inv_x1_sg U56214 ( .A(n8757), .X(n47474) );
  nor_x1_sg U56215 ( .A(n8771), .B(n47453), .X(n8770) );
  inv_x1_sg U56216 ( .A(n9577), .X(n47759) );
  nor_x1_sg U56217 ( .A(n9591), .B(n47738), .X(n9590) );
  inv_x1_sg U56218 ( .A(n10396), .X(n48044) );
  nor_x1_sg U56219 ( .A(n10410), .B(n48023), .X(n10409) );
  inv_x1_sg U56220 ( .A(n11215), .X(n48329) );
  nor_x1_sg U56221 ( .A(n11229), .B(n48308), .X(n11228) );
  inv_x1_sg U56222 ( .A(n12034), .X(n48614) );
  nor_x1_sg U56223 ( .A(n12048), .B(n48593), .X(n12047) );
  inv_x1_sg U56224 ( .A(n12853), .X(n48900) );
  nor_x1_sg U56225 ( .A(n12867), .B(n48879), .X(n12866) );
  inv_x1_sg U56226 ( .A(n13672), .X(n49187) );
  nor_x1_sg U56227 ( .A(n13686), .B(n49166), .X(n13685) );
  inv_x1_sg U56228 ( .A(n14491), .X(n49473) );
  nor_x1_sg U56229 ( .A(n14505), .B(n49452), .X(n14504) );
  inv_x1_sg U56230 ( .A(n15310), .X(n49759) );
  nor_x1_sg U56231 ( .A(n15324), .B(n49737), .X(n15323) );
  inv_x1_sg U56232 ( .A(n16129), .X(n50045) );
  nor_x1_sg U56233 ( .A(n16143), .B(n50024), .X(n16142) );
  inv_x1_sg U56234 ( .A(n16946), .X(n50327) );
  nor_x1_sg U56235 ( .A(n16960), .B(n50309), .X(n16959) );
  inv_x1_sg U56236 ( .A(n17767), .X(n50619) );
  nor_x1_sg U56237 ( .A(n17781), .B(n50598), .X(n17780) );
  inv_x1_sg U56238 ( .A(n18588), .X(n50906) );
  nor_x1_sg U56239 ( .A(n18602), .B(n50885), .X(n18601) );
  nor_x1_sg U56240 ( .A(n41725), .B(n41709), .X(n7381) );
  nor_x1_sg U56241 ( .A(n39731), .B(n41664), .X(n7775) );
  nor_x1_sg U56242 ( .A(n39734), .B(n41687), .X(n8593) );
  nor_x1_sg U56243 ( .A(n39737), .B(n39858), .X(n9413) );
  nor_x1_sg U56244 ( .A(n39740), .B(n39864), .X(n10232) );
  nor_x1_sg U56245 ( .A(n39743), .B(n39867), .X(n11051) );
  nor_x1_sg U56246 ( .A(n39746), .B(n39870), .X(n11870) );
  nor_x1_sg U56247 ( .A(n39749), .B(n39873), .X(n12689) );
  nor_x1_sg U56248 ( .A(n39752), .B(n39876), .X(n13508) );
  nor_x1_sg U56249 ( .A(n39755), .B(n39879), .X(n14327) );
  nor_x1_sg U56250 ( .A(n39758), .B(n39897), .X(n15146) );
  nor_x1_sg U56251 ( .A(n39761), .B(n39882), .X(n15965) );
  nor_x1_sg U56252 ( .A(n39764), .B(n39888), .X(n17603) );
  nor_x1_sg U56253 ( .A(n39767), .B(n39891), .X(n18424) );
  nand_x1_sg U56254 ( .A(n22901), .B(n22902), .X(n22900) );
  nand_x1_sg U56255 ( .A(n22904), .B(n39477), .X(n22899) );
  nand_x1_sg U56256 ( .A(n41194), .B(n22903), .X(n22902) );
  nand_x1_sg U56257 ( .A(n22908), .B(n47416), .X(n22907) );
  nand_x1_sg U56258 ( .A(n22911), .B(n41464), .X(n22906) );
  inv_x1_sg U56259 ( .A(n22909), .X(n47416) );
  nand_x1_sg U56260 ( .A(n23178), .B(n23179), .X(n23177) );
  nand_x1_sg U56261 ( .A(n23181), .B(n38815), .X(n23176) );
  nand_x1_sg U56262 ( .A(n39224), .B(n23180), .X(n23179) );
  nand_x1_sg U56263 ( .A(n23185), .B(n47701), .X(n23184) );
  nand_x1_sg U56264 ( .A(n23188), .B(n41318), .X(n23183) );
  inv_x1_sg U56265 ( .A(n23186), .X(n47701) );
  nand_x1_sg U56266 ( .A(n23458), .B(n23459), .X(n23457) );
  nand_x1_sg U56267 ( .A(n23461), .B(n41313), .X(n23456) );
  nand_x1_sg U56268 ( .A(n41183), .B(n23460), .X(n23459) );
  nand_x1_sg U56269 ( .A(n23465), .B(n47986), .X(n23464) );
  nand_x1_sg U56270 ( .A(n23468), .B(n40227), .X(n23463) );
  inv_x1_sg U56271 ( .A(n23466), .X(n47986) );
  nand_x1_sg U56272 ( .A(n23737), .B(n23738), .X(n23736) );
  nand_x1_sg U56273 ( .A(n23740), .B(n41463), .X(n23735) );
  nand_x1_sg U56274 ( .A(n41179), .B(n23739), .X(n23738) );
  nand_x1_sg U56275 ( .A(n23744), .B(n48271), .X(n23743) );
  nand_x1_sg U56276 ( .A(n23747), .B(n41308), .X(n23742) );
  inv_x1_sg U56277 ( .A(n23745), .X(n48271) );
  nand_x1_sg U56278 ( .A(n24016), .B(n24017), .X(n24015) );
  nand_x1_sg U56279 ( .A(n24019), .B(n39280), .X(n24014) );
  nand_x1_sg U56280 ( .A(n39230), .B(n24018), .X(n24017) );
  nand_x1_sg U56281 ( .A(n24023), .B(n48556), .X(n24022) );
  nand_x1_sg U56282 ( .A(n24026), .B(n41316), .X(n24021) );
  inv_x1_sg U56283 ( .A(n24024), .X(n48556) );
  nand_x1_sg U56284 ( .A(n24295), .B(n24296), .X(n24294) );
  nand_x1_sg U56285 ( .A(n24298), .B(n38815), .X(n24293) );
  nand_x1_sg U56286 ( .A(n39232), .B(n24297), .X(n24296) );
  nand_x1_sg U56287 ( .A(n24302), .B(n48841), .X(n24301) );
  nand_x1_sg U56288 ( .A(n24305), .B(n41461), .X(n24300) );
  inv_x1_sg U56289 ( .A(n24303), .X(n48841) );
  nand_x1_sg U56290 ( .A(n24574), .B(n24575), .X(n24573) );
  nand_x1_sg U56291 ( .A(n24577), .B(n40226), .X(n24572) );
  nand_x1_sg U56292 ( .A(n39234), .B(n24576), .X(n24575) );
  nand_x1_sg U56293 ( .A(n24581), .B(n49128), .X(n24580) );
  nand_x1_sg U56294 ( .A(n24584), .B(n39277), .X(n24579) );
  inv_x1_sg U56295 ( .A(n24582), .X(n49128) );
  nand_x1_sg U56296 ( .A(n24852), .B(n24853), .X(n24851) );
  nand_x1_sg U56297 ( .A(n24855), .B(n39280), .X(n24850) );
  nand_x1_sg U56298 ( .A(n41160), .B(n24854), .X(n24853) );
  nand_x1_sg U56299 ( .A(n24859), .B(n49414), .X(n24858) );
  nand_x1_sg U56300 ( .A(n24862), .B(n41315), .X(n24857) );
  inv_x1_sg U56301 ( .A(n24860), .X(n49414) );
  nand_x1_sg U56302 ( .A(n25131), .B(n25132), .X(n25130) );
  nand_x1_sg U56303 ( .A(n25134), .B(n40227), .X(n25129) );
  nand_x1_sg U56304 ( .A(n39238), .B(n25133), .X(n25132) );
  nand_x1_sg U56305 ( .A(n25138), .B(n49700), .X(n25137) );
  nand_x1_sg U56306 ( .A(n25141), .B(n41317), .X(n25136) );
  inv_x1_sg U56307 ( .A(n25139), .X(n49700) );
  nand_x1_sg U56308 ( .A(n25410), .B(n25411), .X(n25409) );
  nand_x1_sg U56309 ( .A(n25413), .B(n39926), .X(n25408) );
  nand_x1_sg U56310 ( .A(n41150), .B(n25412), .X(n25411) );
  nand_x1_sg U56311 ( .A(n25417), .B(n49986), .X(n25416) );
  nand_x1_sg U56312 ( .A(n25420), .B(n38944), .X(n25415) );
  inv_x1_sg U56313 ( .A(n25418), .X(n49986) );
  nand_x1_sg U56314 ( .A(n25689), .B(n25690), .X(n25688) );
  nand_x1_sg U56315 ( .A(n25692), .B(n40225), .X(n25687) );
  nand_x1_sg U56316 ( .A(n41144), .B(n25691), .X(n25690) );
  nand_x1_sg U56317 ( .A(n25696), .B(n50272), .X(n25695) );
  nand_x1_sg U56318 ( .A(n25699), .B(n38944), .X(n25694) );
  inv_x1_sg U56319 ( .A(n25697), .X(n50272) );
  nand_x1_sg U56320 ( .A(n26526), .B(n26527), .X(n26525) );
  nand_x1_sg U56321 ( .A(n26529), .B(n41311), .X(n26524) );
  nand_x1_sg U56322 ( .A(n39246), .B(n26528), .X(n26527) );
  nand_x1_sg U56323 ( .A(n26533), .B(n51133), .X(n26532) );
  nand_x1_sg U56324 ( .A(n26536), .B(n40225), .X(n26531) );
  inv_x1_sg U56325 ( .A(n26534), .X(n51133) );
  nor_x1_sg U56326 ( .A(n6950), .B(n47049), .X(n7573) );
  nor_x1_sg U56327 ( .A(n6949), .B(n47079), .X(n7572) );
  inv_x1_sg U56328 ( .A(n6949), .X(n47049) );
  nor_x1_sg U56329 ( .A(n7767), .B(n47336), .X(n8391) );
  nor_x1_sg U56330 ( .A(n7766), .B(n47365), .X(n8390) );
  inv_x1_sg U56331 ( .A(n7766), .X(n47336) );
  nor_x1_sg U56332 ( .A(n8585), .B(n47621), .X(n9209) );
  nor_x1_sg U56333 ( .A(n8584), .B(n47650), .X(n9208) );
  inv_x1_sg U56334 ( .A(n8584), .X(n47621) );
  nor_x1_sg U56335 ( .A(n9405), .B(n47906), .X(n10029) );
  nor_x1_sg U56336 ( .A(n9404), .B(n47935), .X(n10028) );
  inv_x1_sg U56337 ( .A(n9404), .X(n47906) );
  nor_x1_sg U56338 ( .A(n10224), .B(n48191), .X(n10848) );
  nor_x1_sg U56339 ( .A(n10223), .B(n48220), .X(n10847) );
  inv_x1_sg U56340 ( .A(n10223), .X(n48191) );
  nor_x1_sg U56341 ( .A(n11043), .B(n48476), .X(n11667) );
  nor_x1_sg U56342 ( .A(n11042), .B(n48505), .X(n11666) );
  inv_x1_sg U56343 ( .A(n11042), .X(n48476) );
  nor_x1_sg U56344 ( .A(n11862), .B(n48761), .X(n12486) );
  nor_x1_sg U56345 ( .A(n11861), .B(n48790), .X(n12485) );
  inv_x1_sg U56346 ( .A(n11861), .X(n48761) );
  nor_x1_sg U56347 ( .A(n12681), .B(n49047), .X(n13305) );
  nor_x1_sg U56348 ( .A(n12680), .B(n49077), .X(n13304) );
  inv_x1_sg U56349 ( .A(n12680), .X(n49047) );
  nor_x1_sg U56350 ( .A(n13500), .B(n49334), .X(n14124) );
  nor_x1_sg U56351 ( .A(n13499), .B(n49363), .X(n14123) );
  inv_x1_sg U56352 ( .A(n13499), .X(n49334) );
  nor_x1_sg U56353 ( .A(n14319), .B(n49620), .X(n14943) );
  nor_x1_sg U56354 ( .A(n14318), .B(n49649), .X(n14942) );
  inv_x1_sg U56355 ( .A(n14318), .X(n49620) );
  nor_x1_sg U56356 ( .A(n15138), .B(n49906), .X(n15762) );
  nor_x1_sg U56357 ( .A(n15137), .B(n49935), .X(n15761) );
  inv_x1_sg U56358 ( .A(n15137), .X(n49906) );
  nor_x1_sg U56359 ( .A(n15957), .B(n50192), .X(n16581) );
  nor_x1_sg U56360 ( .A(n15956), .B(n50221), .X(n16580) );
  inv_x1_sg U56361 ( .A(n15956), .X(n50192) );
  nor_x1_sg U56362 ( .A(n16774), .B(n50477), .X(n17398) );
  nor_x1_sg U56363 ( .A(n16773), .B(n50506), .X(n17397) );
  inv_x1_sg U56364 ( .A(n16773), .X(n50477) );
  nor_x1_sg U56365 ( .A(n17595), .B(n50766), .X(n18219) );
  nor_x1_sg U56366 ( .A(n17594), .B(n50795), .X(n18218) );
  inv_x1_sg U56367 ( .A(n17594), .X(n50766) );
  nor_x1_sg U56368 ( .A(n18416), .B(n51053), .X(n19040) );
  nor_x1_sg U56369 ( .A(n18415), .B(n51082), .X(n19039) );
  inv_x1_sg U56370 ( .A(n18415), .X(n51053) );
  nor_x1_sg U56371 ( .A(n39679), .B(n41724), .X(n17450) );
  nor_x1_sg U56372 ( .A(n6837), .B(n46855), .X(n6835) );
  nor_x1_sg U56373 ( .A(n6840), .B(n6839), .X(n6837) );
  nand_x1_sg U56374 ( .A(n6839), .B(n6840), .X(n6838) );
  nor_x1_sg U56375 ( .A(n7654), .B(n47148), .X(n7652) );
  nor_x1_sg U56376 ( .A(n7657), .B(n7656), .X(n7654) );
  nand_x1_sg U56377 ( .A(n7656), .B(n7657), .X(n7655) );
  nor_x1_sg U56378 ( .A(n8472), .B(n47433), .X(n8470) );
  nor_x1_sg U56379 ( .A(n8475), .B(n8474), .X(n8472) );
  nand_x1_sg U56380 ( .A(n8474), .B(n8475), .X(n8473) );
  nor_x1_sg U56381 ( .A(n9292), .B(n47718), .X(n9290) );
  nor_x1_sg U56382 ( .A(n9295), .B(n9294), .X(n9292) );
  nand_x1_sg U56383 ( .A(n9294), .B(n9295), .X(n9293) );
  nor_x1_sg U56384 ( .A(n10111), .B(n48003), .X(n10109) );
  nor_x1_sg U56385 ( .A(n10114), .B(n10113), .X(n10111) );
  nand_x1_sg U56386 ( .A(n10113), .B(n10114), .X(n10112) );
  nor_x1_sg U56387 ( .A(n10930), .B(n48288), .X(n10928) );
  nor_x1_sg U56388 ( .A(n10933), .B(n10932), .X(n10930) );
  nand_x1_sg U56389 ( .A(n10932), .B(n10933), .X(n10931) );
  nor_x1_sg U56390 ( .A(n11749), .B(n48573), .X(n11747) );
  nor_x1_sg U56391 ( .A(n11752), .B(n11751), .X(n11749) );
  nand_x1_sg U56392 ( .A(n11751), .B(n11752), .X(n11750) );
  nor_x1_sg U56393 ( .A(n12568), .B(n48859), .X(n12566) );
  nor_x1_sg U56394 ( .A(n12571), .B(n12570), .X(n12568) );
  nand_x1_sg U56395 ( .A(n12570), .B(n12571), .X(n12569) );
  nor_x1_sg U56396 ( .A(n13387), .B(n49146), .X(n13385) );
  nor_x1_sg U56397 ( .A(n13390), .B(n13389), .X(n13387) );
  nand_x1_sg U56398 ( .A(n13389), .B(n13390), .X(n13388) );
  nor_x1_sg U56399 ( .A(n14206), .B(n49432), .X(n14204) );
  nor_x1_sg U56400 ( .A(n14209), .B(n14208), .X(n14206) );
  nand_x1_sg U56401 ( .A(n14208), .B(n14209), .X(n14207) );
  nor_x1_sg U56402 ( .A(n15025), .B(n49717), .X(n15023) );
  nor_x1_sg U56403 ( .A(n15028), .B(n15027), .X(n15025) );
  nand_x1_sg U56404 ( .A(n15027), .B(n15028), .X(n15026) );
  nor_x1_sg U56405 ( .A(n15844), .B(n50004), .X(n15842) );
  nor_x1_sg U56406 ( .A(n15847), .B(n15846), .X(n15844) );
  nand_x1_sg U56407 ( .A(n15846), .B(n15847), .X(n15845) );
  nor_x1_sg U56408 ( .A(n16661), .B(n50287), .X(n16659) );
  nor_x1_sg U56409 ( .A(n16664), .B(n16663), .X(n16661) );
  nand_x1_sg U56410 ( .A(n16663), .B(n16664), .X(n16662) );
  nor_x1_sg U56411 ( .A(n17482), .B(n50578), .X(n17480) );
  nor_x1_sg U56412 ( .A(n17485), .B(n17484), .X(n17482) );
  nand_x1_sg U56413 ( .A(n17484), .B(n17485), .X(n17483) );
  nor_x1_sg U56414 ( .A(n18303), .B(n50865), .X(n18301) );
  nor_x1_sg U56415 ( .A(n18306), .B(n18305), .X(n18303) );
  nand_x1_sg U56416 ( .A(n18305), .B(n18306), .X(n18304) );
  nor_x1_sg U56417 ( .A(n46962), .B(n7275), .X(n7274) );
  nor_x1_sg U56418 ( .A(n46920), .B(n7276), .X(n7273) );
  inv_x1_sg U56419 ( .A(n7275), .X(n46920) );
  nor_x1_sg U56420 ( .A(n47253), .B(n8094), .X(n8093) );
  nor_x1_sg U56421 ( .A(n47212), .B(n8095), .X(n8092) );
  inv_x1_sg U56422 ( .A(n8094), .X(n47212) );
  nor_x1_sg U56423 ( .A(n47538), .B(n8912), .X(n8911) );
  nor_x1_sg U56424 ( .A(n47497), .B(n8913), .X(n8910) );
  inv_x1_sg U56425 ( .A(n8912), .X(n47497) );
  nor_x1_sg U56426 ( .A(n47823), .B(n9732), .X(n9731) );
  nor_x1_sg U56427 ( .A(n47782), .B(n9733), .X(n9730) );
  inv_x1_sg U56428 ( .A(n9732), .X(n47782) );
  nor_x1_sg U56429 ( .A(n48108), .B(n10551), .X(n10550) );
  nor_x1_sg U56430 ( .A(n48067), .B(n10552), .X(n10549) );
  inv_x1_sg U56431 ( .A(n10551), .X(n48067) );
  nor_x1_sg U56432 ( .A(n48393), .B(n11370), .X(n11369) );
  nor_x1_sg U56433 ( .A(n48352), .B(n11371), .X(n11368) );
  inv_x1_sg U56434 ( .A(n11370), .X(n48352) );
  nor_x1_sg U56435 ( .A(n48678), .B(n12189), .X(n12188) );
  nor_x1_sg U56436 ( .A(n48637), .B(n12190), .X(n12187) );
  inv_x1_sg U56437 ( .A(n12189), .X(n48637) );
  nor_x1_sg U56438 ( .A(n48964), .B(n13008), .X(n13007) );
  nor_x1_sg U56439 ( .A(n48923), .B(n13009), .X(n13006) );
  inv_x1_sg U56440 ( .A(n13008), .X(n48923) );
  nor_x1_sg U56441 ( .A(n49251), .B(n13827), .X(n13826) );
  nor_x1_sg U56442 ( .A(n49210), .B(n13828), .X(n13825) );
  inv_x1_sg U56443 ( .A(n13827), .X(n49210) );
  nor_x1_sg U56444 ( .A(n49537), .B(n14646), .X(n14645) );
  nor_x1_sg U56445 ( .A(n49496), .B(n14647), .X(n14644) );
  inv_x1_sg U56446 ( .A(n14646), .X(n49496) );
  nor_x1_sg U56447 ( .A(n49823), .B(n15465), .X(n15464) );
  nor_x1_sg U56448 ( .A(n49782), .B(n15466), .X(n15463) );
  inv_x1_sg U56449 ( .A(n15465), .X(n49782) );
  nor_x1_sg U56450 ( .A(n50109), .B(n16284), .X(n16283) );
  nor_x1_sg U56451 ( .A(n50068), .B(n16285), .X(n16282) );
  inv_x1_sg U56452 ( .A(n16284), .X(n50068) );
  nor_x1_sg U56453 ( .A(n50683), .B(n17922), .X(n17921) );
  nor_x1_sg U56454 ( .A(n50642), .B(n17923), .X(n17920) );
  inv_x1_sg U56455 ( .A(n17922), .X(n50642) );
  nor_x1_sg U56456 ( .A(n50970), .B(n18743), .X(n18742) );
  nor_x1_sg U56457 ( .A(n50929), .B(n18744), .X(n18741) );
  inv_x1_sg U56458 ( .A(n18743), .X(n50929) );
  nor_x1_sg U56459 ( .A(n6939), .B(n47080), .X(n6938) );
  nor_x1_sg U56460 ( .A(n6940), .B(n47101), .X(n6937) );
  inv_x1_sg U56461 ( .A(n6940), .X(n47080) );
  nor_x1_sg U56462 ( .A(n7756), .B(n47366), .X(n7755) );
  nor_x1_sg U56463 ( .A(n7757), .B(n47387), .X(n7754) );
  inv_x1_sg U56464 ( .A(n7757), .X(n47366) );
  nor_x1_sg U56465 ( .A(n8574), .B(n47651), .X(n8573) );
  nor_x1_sg U56466 ( .A(n8575), .B(n47672), .X(n8572) );
  inv_x1_sg U56467 ( .A(n8575), .X(n47651) );
  nor_x1_sg U56468 ( .A(n9394), .B(n47936), .X(n9393) );
  nor_x1_sg U56469 ( .A(n9395), .B(n47957), .X(n9392) );
  inv_x1_sg U56470 ( .A(n9395), .X(n47936) );
  nor_x1_sg U56471 ( .A(n10213), .B(n48221), .X(n10212) );
  nor_x1_sg U56472 ( .A(n10214), .B(n48242), .X(n10211) );
  inv_x1_sg U56473 ( .A(n10214), .X(n48221) );
  nor_x1_sg U56474 ( .A(n11032), .B(n48506), .X(n11031) );
  nor_x1_sg U56475 ( .A(n11033), .B(n48527), .X(n11030) );
  inv_x1_sg U56476 ( .A(n11033), .X(n48506) );
  nor_x1_sg U56477 ( .A(n11851), .B(n48791), .X(n11850) );
  nor_x1_sg U56478 ( .A(n11852), .B(n48812), .X(n11849) );
  inv_x1_sg U56479 ( .A(n11852), .X(n48791) );
  nor_x1_sg U56480 ( .A(n12670), .B(n49078), .X(n12669) );
  nor_x1_sg U56481 ( .A(n12671), .B(n49099), .X(n12668) );
  inv_x1_sg U56482 ( .A(n12671), .X(n49078) );
  nor_x1_sg U56483 ( .A(n13489), .B(n49364), .X(n13488) );
  nor_x1_sg U56484 ( .A(n13490), .B(n49385), .X(n13487) );
  inv_x1_sg U56485 ( .A(n13490), .X(n49364) );
  nor_x1_sg U56486 ( .A(n14308), .B(n49650), .X(n14307) );
  nor_x1_sg U56487 ( .A(n14309), .B(n49671), .X(n14306) );
  inv_x1_sg U56488 ( .A(n14309), .X(n49650) );
  nor_x1_sg U56489 ( .A(n15127), .B(n49936), .X(n15126) );
  nor_x1_sg U56490 ( .A(n15128), .B(n49957), .X(n15125) );
  inv_x1_sg U56491 ( .A(n15128), .X(n49936) );
  nor_x1_sg U56492 ( .A(n15946), .B(n50222), .X(n15945) );
  nor_x1_sg U56493 ( .A(n15947), .B(n50243), .X(n15944) );
  inv_x1_sg U56494 ( .A(n15947), .X(n50222) );
  nor_x1_sg U56495 ( .A(n16763), .B(n50507), .X(n16762) );
  nor_x1_sg U56496 ( .A(n16764), .B(n50528), .X(n16761) );
  inv_x1_sg U56497 ( .A(n16764), .X(n50507) );
  nor_x1_sg U56498 ( .A(n17584), .B(n50796), .X(n17583) );
  nor_x1_sg U56499 ( .A(n17585), .B(n50817), .X(n17582) );
  inv_x1_sg U56500 ( .A(n17585), .X(n50796) );
  nor_x1_sg U56501 ( .A(n18405), .B(n51083), .X(n18404) );
  nor_x1_sg U56502 ( .A(n18406), .B(n51104), .X(n18403) );
  inv_x1_sg U56503 ( .A(n18406), .X(n51083) );
  nand_x1_sg U56504 ( .A(n26236), .B(n26237), .X(n26235) );
  nand_x1_sg U56505 ( .A(n26239), .B(n39927), .X(n26234) );
  nand_x1_sg U56506 ( .A(n39244), .B(n26238), .X(n26237) );
  nand_x1_sg U56507 ( .A(n26244), .B(n50847), .X(n26243) );
  nand_x1_sg U56508 ( .A(n26247), .B(n39475), .X(n26242) );
  inv_x1_sg U56509 ( .A(n26245), .X(n50847) );
  nor_x1_sg U56510 ( .A(n47031), .B(n7530), .X(n7480) );
  inv_x1_sg U56511 ( .A(n7525), .X(n47031) );
  nor_x1_sg U56512 ( .A(n7531), .B(n7532), .X(n7530) );
  nor_x1_sg U56513 ( .A(n47318), .B(n8348), .X(n8298) );
  inv_x1_sg U56514 ( .A(n8343), .X(n47318) );
  nor_x1_sg U56515 ( .A(n8349), .B(n8350), .X(n8348) );
  nor_x1_sg U56516 ( .A(n47603), .B(n9166), .X(n9116) );
  inv_x1_sg U56517 ( .A(n9161), .X(n47603) );
  nor_x1_sg U56518 ( .A(n9167), .B(n9168), .X(n9166) );
  nor_x1_sg U56519 ( .A(n47888), .B(n9986), .X(n9936) );
  inv_x1_sg U56520 ( .A(n9981), .X(n47888) );
  nor_x1_sg U56521 ( .A(n9987), .B(n9988), .X(n9986) );
  nor_x1_sg U56522 ( .A(n48173), .B(n10805), .X(n10755) );
  inv_x1_sg U56523 ( .A(n10800), .X(n48173) );
  nor_x1_sg U56524 ( .A(n10806), .B(n10807), .X(n10805) );
  nor_x1_sg U56525 ( .A(n48458), .B(n11624), .X(n11574) );
  inv_x1_sg U56526 ( .A(n11619), .X(n48458) );
  nor_x1_sg U56527 ( .A(n11625), .B(n11626), .X(n11624) );
  nor_x1_sg U56528 ( .A(n48743), .B(n12443), .X(n12393) );
  inv_x1_sg U56529 ( .A(n12438), .X(n48743) );
  nor_x1_sg U56530 ( .A(n12444), .B(n12445), .X(n12443) );
  nor_x1_sg U56531 ( .A(n49029), .B(n13262), .X(n13212) );
  inv_x1_sg U56532 ( .A(n13257), .X(n49029) );
  nor_x1_sg U56533 ( .A(n13263), .B(n13264), .X(n13262) );
  nor_x1_sg U56534 ( .A(n49316), .B(n14081), .X(n14031) );
  inv_x1_sg U56535 ( .A(n14076), .X(n49316) );
  nor_x1_sg U56536 ( .A(n14082), .B(n14083), .X(n14081) );
  nor_x1_sg U56537 ( .A(n49602), .B(n14900), .X(n14850) );
  inv_x1_sg U56538 ( .A(n14895), .X(n49602) );
  nor_x1_sg U56539 ( .A(n14901), .B(n14902), .X(n14900) );
  nor_x1_sg U56540 ( .A(n49888), .B(n15719), .X(n15669) );
  inv_x1_sg U56541 ( .A(n15714), .X(n49888) );
  nor_x1_sg U56542 ( .A(n15720), .B(n15721), .X(n15719) );
  nor_x1_sg U56543 ( .A(n50174), .B(n16538), .X(n16488) );
  inv_x1_sg U56544 ( .A(n16533), .X(n50174) );
  nor_x1_sg U56545 ( .A(n16539), .B(n16540), .X(n16538) );
  nor_x1_sg U56546 ( .A(n50459), .B(n17355), .X(n17305) );
  inv_x1_sg U56547 ( .A(n17350), .X(n50459) );
  nor_x1_sg U56548 ( .A(n17356), .B(n17357), .X(n17355) );
  nor_x1_sg U56549 ( .A(n50748), .B(n18176), .X(n18126) );
  inv_x1_sg U56550 ( .A(n18171), .X(n50748) );
  nor_x1_sg U56551 ( .A(n18177), .B(n18178), .X(n18176) );
  nor_x1_sg U56552 ( .A(n51035), .B(n18997), .X(n18947) );
  inv_x1_sg U56553 ( .A(n18992), .X(n51035) );
  nor_x1_sg U56554 ( .A(n18998), .B(n18999), .X(n18997) );
  nor_x1_sg U56555 ( .A(n47012), .B(n7359), .X(n7320) );
  inv_x1_sg U56556 ( .A(n7362), .X(n47012) );
  nor_x1_sg U56557 ( .A(n7360), .B(n7361), .X(n7359) );
  nor_x1_sg U56558 ( .A(n47300), .B(n8177), .X(n8138) );
  inv_x1_sg U56559 ( .A(n8180), .X(n47300) );
  nor_x1_sg U56560 ( .A(n8178), .B(n8179), .X(n8177) );
  nor_x1_sg U56561 ( .A(n47585), .B(n8995), .X(n8956) );
  inv_x1_sg U56562 ( .A(n8998), .X(n47585) );
  nor_x1_sg U56563 ( .A(n8996), .B(n8997), .X(n8995) );
  nor_x1_sg U56564 ( .A(n47870), .B(n9815), .X(n9776) );
  inv_x1_sg U56565 ( .A(n9818), .X(n47870) );
  nor_x1_sg U56566 ( .A(n9816), .B(n9817), .X(n9815) );
  nor_x1_sg U56567 ( .A(n48155), .B(n10634), .X(n10595) );
  inv_x1_sg U56568 ( .A(n10637), .X(n48155) );
  nor_x1_sg U56569 ( .A(n10635), .B(n10636), .X(n10634) );
  nor_x1_sg U56570 ( .A(n48440), .B(n11453), .X(n11414) );
  inv_x1_sg U56571 ( .A(n11456), .X(n48440) );
  nor_x1_sg U56572 ( .A(n11454), .B(n11455), .X(n11453) );
  nor_x1_sg U56573 ( .A(n48725), .B(n12272), .X(n12233) );
  inv_x1_sg U56574 ( .A(n12275), .X(n48725) );
  nor_x1_sg U56575 ( .A(n12273), .B(n12274), .X(n12272) );
  nor_x1_sg U56576 ( .A(n49011), .B(n13091), .X(n13052) );
  inv_x1_sg U56577 ( .A(n13094), .X(n49011) );
  nor_x1_sg U56578 ( .A(n13092), .B(n13093), .X(n13091) );
  nor_x1_sg U56579 ( .A(n49298), .B(n13910), .X(n13871) );
  inv_x1_sg U56580 ( .A(n13913), .X(n49298) );
  nor_x1_sg U56581 ( .A(n13911), .B(n13912), .X(n13910) );
  nor_x1_sg U56582 ( .A(n49584), .B(n14729), .X(n14690) );
  inv_x1_sg U56583 ( .A(n14732), .X(n49584) );
  nor_x1_sg U56584 ( .A(n14730), .B(n14731), .X(n14729) );
  nor_x1_sg U56585 ( .A(n49870), .B(n15548), .X(n15509) );
  inv_x1_sg U56586 ( .A(n15551), .X(n49870) );
  nor_x1_sg U56587 ( .A(n15549), .B(n15550), .X(n15548) );
  nor_x1_sg U56588 ( .A(n50156), .B(n16367), .X(n16328) );
  inv_x1_sg U56589 ( .A(n16370), .X(n50156) );
  nor_x1_sg U56590 ( .A(n16368), .B(n16369), .X(n16367) );
  nor_x1_sg U56591 ( .A(n50441), .B(n17184), .X(n17145) );
  inv_x1_sg U56592 ( .A(n17187), .X(n50441) );
  nor_x1_sg U56593 ( .A(n17185), .B(n17186), .X(n17184) );
  nor_x1_sg U56594 ( .A(n50730), .B(n18005), .X(n17966) );
  inv_x1_sg U56595 ( .A(n18008), .X(n50730) );
  nor_x1_sg U56596 ( .A(n18006), .B(n18007), .X(n18005) );
  nor_x1_sg U56597 ( .A(n51017), .B(n18826), .X(n18787) );
  inv_x1_sg U56598 ( .A(n18829), .X(n51017) );
  nor_x1_sg U56599 ( .A(n18827), .B(n18828), .X(n18826) );
  nor_x1_sg U56600 ( .A(n47108), .B(n7024), .X(n7018) );
  nor_x1_sg U56601 ( .A(n7025), .B(n47107), .X(n7024) );
  nand_x1_sg U56602 ( .A(n47107), .B(n7025), .X(n7026) );
  nor_x1_sg U56603 ( .A(n47394), .B(n7842), .X(n7836) );
  nor_x1_sg U56604 ( .A(n7843), .B(n47393), .X(n7842) );
  nand_x1_sg U56605 ( .A(n47393), .B(n7843), .X(n7844) );
  nor_x1_sg U56606 ( .A(n47679), .B(n8660), .X(n8654) );
  nor_x1_sg U56607 ( .A(n8661), .B(n47678), .X(n8660) );
  nand_x1_sg U56608 ( .A(n47678), .B(n8661), .X(n8662) );
  nor_x1_sg U56609 ( .A(n47964), .B(n9480), .X(n9474) );
  nor_x1_sg U56610 ( .A(n9481), .B(n47963), .X(n9480) );
  nand_x1_sg U56611 ( .A(n47963), .B(n9481), .X(n9482) );
  nor_x1_sg U56612 ( .A(n48249), .B(n10299), .X(n10293) );
  nor_x1_sg U56613 ( .A(n10300), .B(n48248), .X(n10299) );
  nand_x1_sg U56614 ( .A(n48248), .B(n10300), .X(n10301) );
  nor_x1_sg U56615 ( .A(n48534), .B(n11118), .X(n11112) );
  nor_x1_sg U56616 ( .A(n11119), .B(n48533), .X(n11118) );
  nand_x1_sg U56617 ( .A(n48533), .B(n11119), .X(n11120) );
  nor_x1_sg U56618 ( .A(n48819), .B(n11937), .X(n11931) );
  nor_x1_sg U56619 ( .A(n11938), .B(n48818), .X(n11937) );
  nand_x1_sg U56620 ( .A(n48818), .B(n11938), .X(n11939) );
  nor_x1_sg U56621 ( .A(n49106), .B(n12756), .X(n12750) );
  nor_x1_sg U56622 ( .A(n12757), .B(n49105), .X(n12756) );
  nand_x1_sg U56623 ( .A(n49105), .B(n12757), .X(n12758) );
  nor_x1_sg U56624 ( .A(n49392), .B(n13575), .X(n13569) );
  nor_x1_sg U56625 ( .A(n13576), .B(n49391), .X(n13575) );
  nand_x1_sg U56626 ( .A(n49391), .B(n13576), .X(n13577) );
  nor_x1_sg U56627 ( .A(n49678), .B(n14394), .X(n14388) );
  nor_x1_sg U56628 ( .A(n14395), .B(n49677), .X(n14394) );
  nand_x1_sg U56629 ( .A(n49677), .B(n14395), .X(n14396) );
  nor_x1_sg U56630 ( .A(n49964), .B(n15213), .X(n15207) );
  nor_x1_sg U56631 ( .A(n15214), .B(n49963), .X(n15213) );
  nand_x1_sg U56632 ( .A(n49963), .B(n15214), .X(n15215) );
  nor_x1_sg U56633 ( .A(n50250), .B(n16032), .X(n16026) );
  nor_x1_sg U56634 ( .A(n16033), .B(n50249), .X(n16032) );
  nand_x1_sg U56635 ( .A(n50249), .B(n16033), .X(n16034) );
  nor_x1_sg U56636 ( .A(n50535), .B(n16851), .X(n16843) );
  nor_x1_sg U56637 ( .A(n16852), .B(n50534), .X(n16851) );
  nand_x1_sg U56638 ( .A(n50534), .B(n16852), .X(n16853) );
  nor_x1_sg U56639 ( .A(n50824), .B(n17670), .X(n17664) );
  nor_x1_sg U56640 ( .A(n17671), .B(n50823), .X(n17670) );
  nand_x1_sg U56641 ( .A(n50823), .B(n17671), .X(n17672) );
  nor_x1_sg U56642 ( .A(n51111), .B(n18491), .X(n18485) );
  nor_x1_sg U56643 ( .A(n18492), .B(n51110), .X(n18491) );
  nand_x1_sg U56644 ( .A(n51110), .B(n18492), .X(n18493) );
  nor_x1_sg U56645 ( .A(n46873), .B(n6851), .X(n6849) );
  nor_x1_sg U56646 ( .A(n6852), .B(n46872), .X(n6851) );
  nand_x1_sg U56647 ( .A(n46872), .B(n6852), .X(n6853) );
  nor_x1_sg U56648 ( .A(n46885), .B(n6857), .X(n6855) );
  nor_x1_sg U56649 ( .A(n6858), .B(n6859), .X(n6857) );
  nand_x1_sg U56650 ( .A(n6859), .B(n6858), .X(n6860) );
  nor_x1_sg U56651 ( .A(n46932), .B(n6875), .X(n6873) );
  nor_x1_sg U56652 ( .A(n6876), .B(n6877), .X(n6875) );
  nand_x1_sg U56653 ( .A(n6877), .B(n6876), .X(n6878) );
  nor_x1_sg U56654 ( .A(n46980), .B(n6887), .X(n6885) );
  nor_x1_sg U56655 ( .A(n6888), .B(n6889), .X(n6887) );
  nand_x1_sg U56656 ( .A(n6889), .B(n6888), .X(n6890) );
  nor_x1_sg U56657 ( .A(n47166), .B(n7668), .X(n7666) );
  nor_x1_sg U56658 ( .A(n7669), .B(n47165), .X(n7668) );
  nand_x1_sg U56659 ( .A(n47165), .B(n7669), .X(n7670) );
  nor_x1_sg U56660 ( .A(n47178), .B(n7674), .X(n7672) );
  nor_x1_sg U56661 ( .A(n7675), .B(n7676), .X(n7674) );
  nand_x1_sg U56662 ( .A(n7676), .B(n7675), .X(n7677) );
  nor_x1_sg U56663 ( .A(n47224), .B(n7692), .X(n7690) );
  nor_x1_sg U56664 ( .A(n7693), .B(n7694), .X(n7692) );
  nand_x1_sg U56665 ( .A(n7694), .B(n7693), .X(n7695) );
  nor_x1_sg U56666 ( .A(n47270), .B(n7704), .X(n7702) );
  nor_x1_sg U56667 ( .A(n7705), .B(n7706), .X(n7704) );
  nand_x1_sg U56668 ( .A(n7706), .B(n7705), .X(n7707) );
  nor_x1_sg U56669 ( .A(n47451), .B(n8486), .X(n8484) );
  nor_x1_sg U56670 ( .A(n8487), .B(n47450), .X(n8486) );
  nand_x1_sg U56671 ( .A(n47450), .B(n8487), .X(n8488) );
  nor_x1_sg U56672 ( .A(n47463), .B(n8492), .X(n8490) );
  nor_x1_sg U56673 ( .A(n8493), .B(n8494), .X(n8492) );
  nand_x1_sg U56674 ( .A(n8494), .B(n8493), .X(n8495) );
  nor_x1_sg U56675 ( .A(n47509), .B(n8510), .X(n8508) );
  nor_x1_sg U56676 ( .A(n8511), .B(n8512), .X(n8510) );
  nand_x1_sg U56677 ( .A(n8512), .B(n8511), .X(n8513) );
  nor_x1_sg U56678 ( .A(n47555), .B(n8522), .X(n8520) );
  nor_x1_sg U56679 ( .A(n8523), .B(n8524), .X(n8522) );
  nand_x1_sg U56680 ( .A(n8524), .B(n8523), .X(n8525) );
  nor_x1_sg U56681 ( .A(n47736), .B(n9306), .X(n9304) );
  nor_x1_sg U56682 ( .A(n9307), .B(n47735), .X(n9306) );
  nand_x1_sg U56683 ( .A(n47735), .B(n9307), .X(n9308) );
  nor_x1_sg U56684 ( .A(n47748), .B(n9312), .X(n9310) );
  nor_x1_sg U56685 ( .A(n9313), .B(n9314), .X(n9312) );
  nand_x1_sg U56686 ( .A(n9314), .B(n9313), .X(n9315) );
  nor_x1_sg U56687 ( .A(n47794), .B(n9330), .X(n9328) );
  nor_x1_sg U56688 ( .A(n9331), .B(n9332), .X(n9330) );
  nand_x1_sg U56689 ( .A(n9332), .B(n9331), .X(n9333) );
  nor_x1_sg U56690 ( .A(n47840), .B(n9342), .X(n9340) );
  nor_x1_sg U56691 ( .A(n9343), .B(n9344), .X(n9342) );
  nand_x1_sg U56692 ( .A(n9344), .B(n9343), .X(n9345) );
  nor_x1_sg U56693 ( .A(n48021), .B(n10125), .X(n10123) );
  nor_x1_sg U56694 ( .A(n10126), .B(n48020), .X(n10125) );
  nand_x1_sg U56695 ( .A(n48020), .B(n10126), .X(n10127) );
  nor_x1_sg U56696 ( .A(n48033), .B(n10131), .X(n10129) );
  nor_x1_sg U56697 ( .A(n10132), .B(n10133), .X(n10131) );
  nand_x1_sg U56698 ( .A(n10133), .B(n10132), .X(n10134) );
  nor_x1_sg U56699 ( .A(n48079), .B(n10149), .X(n10147) );
  nor_x1_sg U56700 ( .A(n10150), .B(n10151), .X(n10149) );
  nand_x1_sg U56701 ( .A(n10151), .B(n10150), .X(n10152) );
  nor_x1_sg U56702 ( .A(n48125), .B(n10161), .X(n10159) );
  nor_x1_sg U56703 ( .A(n10162), .B(n10163), .X(n10161) );
  nand_x1_sg U56704 ( .A(n10163), .B(n10162), .X(n10164) );
  nor_x1_sg U56705 ( .A(n48306), .B(n10944), .X(n10942) );
  nor_x1_sg U56706 ( .A(n10945), .B(n48305), .X(n10944) );
  nand_x1_sg U56707 ( .A(n48305), .B(n10945), .X(n10946) );
  nor_x1_sg U56708 ( .A(n48318), .B(n10950), .X(n10948) );
  nor_x1_sg U56709 ( .A(n10951), .B(n10952), .X(n10950) );
  nand_x1_sg U56710 ( .A(n10952), .B(n10951), .X(n10953) );
  nor_x1_sg U56711 ( .A(n48364), .B(n10968), .X(n10966) );
  nor_x1_sg U56712 ( .A(n10969), .B(n10970), .X(n10968) );
  nand_x1_sg U56713 ( .A(n10970), .B(n10969), .X(n10971) );
  nor_x1_sg U56714 ( .A(n48410), .B(n10980), .X(n10978) );
  nor_x1_sg U56715 ( .A(n10981), .B(n10982), .X(n10980) );
  nand_x1_sg U56716 ( .A(n10982), .B(n10981), .X(n10983) );
  nor_x1_sg U56717 ( .A(n48591), .B(n11763), .X(n11761) );
  nor_x1_sg U56718 ( .A(n11764), .B(n48590), .X(n11763) );
  nand_x1_sg U56719 ( .A(n48590), .B(n11764), .X(n11765) );
  nor_x1_sg U56720 ( .A(n48603), .B(n11769), .X(n11767) );
  nor_x1_sg U56721 ( .A(n11770), .B(n11771), .X(n11769) );
  nand_x1_sg U56722 ( .A(n11771), .B(n11770), .X(n11772) );
  nor_x1_sg U56723 ( .A(n48649), .B(n11787), .X(n11785) );
  nor_x1_sg U56724 ( .A(n11788), .B(n11789), .X(n11787) );
  nand_x1_sg U56725 ( .A(n11789), .B(n11788), .X(n11790) );
  nor_x1_sg U56726 ( .A(n48695), .B(n11799), .X(n11797) );
  nor_x1_sg U56727 ( .A(n11800), .B(n11801), .X(n11799) );
  nand_x1_sg U56728 ( .A(n11801), .B(n11800), .X(n11802) );
  nor_x1_sg U56729 ( .A(n48877), .B(n12582), .X(n12580) );
  nor_x1_sg U56730 ( .A(n12583), .B(n48876), .X(n12582) );
  nand_x1_sg U56731 ( .A(n48876), .B(n12583), .X(n12584) );
  nor_x1_sg U56732 ( .A(n48889), .B(n12588), .X(n12586) );
  nor_x1_sg U56733 ( .A(n12589), .B(n12590), .X(n12588) );
  nand_x1_sg U56734 ( .A(n12590), .B(n12589), .X(n12591) );
  nor_x1_sg U56735 ( .A(n48935), .B(n12606), .X(n12604) );
  nor_x1_sg U56736 ( .A(n12607), .B(n12608), .X(n12606) );
  nand_x1_sg U56737 ( .A(n12608), .B(n12607), .X(n12609) );
  nor_x1_sg U56738 ( .A(n48981), .B(n12618), .X(n12616) );
  nor_x1_sg U56739 ( .A(n12619), .B(n12620), .X(n12618) );
  nand_x1_sg U56740 ( .A(n12620), .B(n12619), .X(n12621) );
  nor_x1_sg U56741 ( .A(n49164), .B(n13401), .X(n13399) );
  nor_x1_sg U56742 ( .A(n13402), .B(n49163), .X(n13401) );
  nand_x1_sg U56743 ( .A(n49163), .B(n13402), .X(n13403) );
  nor_x1_sg U56744 ( .A(n49176), .B(n13407), .X(n13405) );
  nor_x1_sg U56745 ( .A(n13408), .B(n13409), .X(n13407) );
  nand_x1_sg U56746 ( .A(n13409), .B(n13408), .X(n13410) );
  nor_x1_sg U56747 ( .A(n49222), .B(n13425), .X(n13423) );
  nor_x1_sg U56748 ( .A(n13426), .B(n13427), .X(n13425) );
  nand_x1_sg U56749 ( .A(n13427), .B(n13426), .X(n13428) );
  nor_x1_sg U56750 ( .A(n49268), .B(n13437), .X(n13435) );
  nor_x1_sg U56751 ( .A(n13438), .B(n13439), .X(n13437) );
  nand_x1_sg U56752 ( .A(n13439), .B(n13438), .X(n13440) );
  nor_x1_sg U56753 ( .A(n49450), .B(n14220), .X(n14218) );
  nor_x1_sg U56754 ( .A(n14221), .B(n49449), .X(n14220) );
  nand_x1_sg U56755 ( .A(n49449), .B(n14221), .X(n14222) );
  nor_x1_sg U56756 ( .A(n49462), .B(n14226), .X(n14224) );
  nor_x1_sg U56757 ( .A(n14227), .B(n14228), .X(n14226) );
  nand_x1_sg U56758 ( .A(n14228), .B(n14227), .X(n14229) );
  nor_x1_sg U56759 ( .A(n49508), .B(n14244), .X(n14242) );
  nor_x1_sg U56760 ( .A(n14245), .B(n14246), .X(n14244) );
  nand_x1_sg U56761 ( .A(n14246), .B(n14245), .X(n14247) );
  nor_x1_sg U56762 ( .A(n49554), .B(n14256), .X(n14254) );
  nor_x1_sg U56763 ( .A(n14257), .B(n14258), .X(n14256) );
  nand_x1_sg U56764 ( .A(n14258), .B(n14257), .X(n14259) );
  nor_x1_sg U56765 ( .A(n49735), .B(n15039), .X(n15037) );
  nor_x1_sg U56766 ( .A(n15040), .B(n49734), .X(n15039) );
  nand_x1_sg U56767 ( .A(n49734), .B(n15040), .X(n15041) );
  nor_x1_sg U56768 ( .A(n49747), .B(n15045), .X(n15043) );
  nor_x1_sg U56769 ( .A(n15046), .B(n15047), .X(n15045) );
  nand_x1_sg U56770 ( .A(n15047), .B(n15046), .X(n15048) );
  nor_x1_sg U56771 ( .A(n49794), .B(n15063), .X(n15061) );
  nor_x1_sg U56772 ( .A(n15064), .B(n15065), .X(n15063) );
  nand_x1_sg U56773 ( .A(n15065), .B(n15064), .X(n15066) );
  nor_x1_sg U56774 ( .A(n49840), .B(n15075), .X(n15073) );
  nor_x1_sg U56775 ( .A(n15076), .B(n15077), .X(n15075) );
  nand_x1_sg U56776 ( .A(n15077), .B(n15076), .X(n15078) );
  nor_x1_sg U56777 ( .A(n50022), .B(n15858), .X(n15856) );
  nor_x1_sg U56778 ( .A(n15859), .B(n50021), .X(n15858) );
  nand_x1_sg U56779 ( .A(n50021), .B(n15859), .X(n15860) );
  nor_x1_sg U56780 ( .A(n50034), .B(n15864), .X(n15862) );
  nor_x1_sg U56781 ( .A(n15865), .B(n15866), .X(n15864) );
  nand_x1_sg U56782 ( .A(n15866), .B(n15865), .X(n15867) );
  nor_x1_sg U56783 ( .A(n50080), .B(n15882), .X(n15880) );
  nor_x1_sg U56784 ( .A(n15883), .B(n15884), .X(n15882) );
  nand_x1_sg U56785 ( .A(n15884), .B(n15883), .X(n15885) );
  nor_x1_sg U56786 ( .A(n50126), .B(n15894), .X(n15892) );
  nor_x1_sg U56787 ( .A(n15895), .B(n15896), .X(n15894) );
  nand_x1_sg U56788 ( .A(n15896), .B(n15895), .X(n15897) );
  nor_x1_sg U56789 ( .A(n50319), .B(n16681), .X(n16679) );
  nor_x1_sg U56790 ( .A(n16682), .B(n16683), .X(n16681) );
  nand_x1_sg U56791 ( .A(n16683), .B(n16682), .X(n16684) );
  nor_x1_sg U56792 ( .A(n50365), .B(n16699), .X(n16697) );
  nor_x1_sg U56793 ( .A(n16700), .B(n16701), .X(n16699) );
  nand_x1_sg U56794 ( .A(n16701), .B(n16700), .X(n16702) );
  nor_x1_sg U56795 ( .A(n50596), .B(n17496), .X(n17494) );
  nor_x1_sg U56796 ( .A(n17497), .B(n50595), .X(n17496) );
  nand_x1_sg U56797 ( .A(n50595), .B(n17497), .X(n17498) );
  nor_x1_sg U56798 ( .A(n50608), .B(n17502), .X(n17500) );
  nor_x1_sg U56799 ( .A(n17503), .B(n17504), .X(n17502) );
  nand_x1_sg U56800 ( .A(n17504), .B(n17503), .X(n17505) );
  nor_x1_sg U56801 ( .A(n50654), .B(n17520), .X(n17518) );
  nor_x1_sg U56802 ( .A(n17521), .B(n17522), .X(n17520) );
  nand_x1_sg U56803 ( .A(n17522), .B(n17521), .X(n17523) );
  nor_x1_sg U56804 ( .A(n50700), .B(n17532), .X(n17530) );
  nor_x1_sg U56805 ( .A(n17533), .B(n17534), .X(n17532) );
  nand_x1_sg U56806 ( .A(n17534), .B(n17533), .X(n17535) );
  nor_x1_sg U56807 ( .A(n50883), .B(n18317), .X(n18315) );
  nor_x1_sg U56808 ( .A(n18318), .B(n50882), .X(n18317) );
  nand_x1_sg U56809 ( .A(n50882), .B(n18318), .X(n18319) );
  nor_x1_sg U56810 ( .A(n50895), .B(n18323), .X(n18321) );
  nor_x1_sg U56811 ( .A(n18324), .B(n18325), .X(n18323) );
  nand_x1_sg U56812 ( .A(n18325), .B(n18324), .X(n18326) );
  nor_x1_sg U56813 ( .A(n50941), .B(n18341), .X(n18339) );
  nor_x1_sg U56814 ( .A(n18342), .B(n18343), .X(n18341) );
  nand_x1_sg U56815 ( .A(n18343), .B(n18342), .X(n18344) );
  nor_x1_sg U56816 ( .A(n50987), .B(n18353), .X(n18351) );
  nor_x1_sg U56817 ( .A(n18354), .B(n18355), .X(n18353) );
  nand_x1_sg U56818 ( .A(n18355), .B(n18354), .X(n18356) );
  nor_x1_sg U56819 ( .A(n47236), .B(n8070), .X(n8048) );
  nor_x1_sg U56820 ( .A(n8071), .B(n8072), .X(n8070) );
  nand_x1_sg U56821 ( .A(n8072), .B(n8071), .X(n8073) );
  nor_x1_sg U56822 ( .A(n47521), .B(n8888), .X(n8866) );
  nor_x1_sg U56823 ( .A(n8889), .B(n8890), .X(n8888) );
  nand_x1_sg U56824 ( .A(n8890), .B(n8889), .X(n8891) );
  nor_x1_sg U56825 ( .A(n47806), .B(n9708), .X(n9686) );
  nor_x1_sg U56826 ( .A(n9709), .B(n9710), .X(n9708) );
  nand_x1_sg U56827 ( .A(n9710), .B(n9709), .X(n9711) );
  nor_x1_sg U56828 ( .A(n48091), .B(n10527), .X(n10505) );
  nor_x1_sg U56829 ( .A(n10528), .B(n10529), .X(n10527) );
  nand_x1_sg U56830 ( .A(n10529), .B(n10528), .X(n10530) );
  nor_x1_sg U56831 ( .A(n48376), .B(n11346), .X(n11324) );
  nor_x1_sg U56832 ( .A(n11347), .B(n11348), .X(n11346) );
  nand_x1_sg U56833 ( .A(n11348), .B(n11347), .X(n11349) );
  nor_x1_sg U56834 ( .A(n48661), .B(n12165), .X(n12143) );
  nor_x1_sg U56835 ( .A(n12166), .B(n12167), .X(n12165) );
  nand_x1_sg U56836 ( .A(n12167), .B(n12166), .X(n12168) );
  nor_x1_sg U56837 ( .A(n48947), .B(n12984), .X(n12962) );
  nor_x1_sg U56838 ( .A(n12985), .B(n12986), .X(n12984) );
  nand_x1_sg U56839 ( .A(n12986), .B(n12985), .X(n12987) );
  nor_x1_sg U56840 ( .A(n49234), .B(n13803), .X(n13781) );
  nor_x1_sg U56841 ( .A(n13804), .B(n13805), .X(n13803) );
  nand_x1_sg U56842 ( .A(n13805), .B(n13804), .X(n13806) );
  nor_x1_sg U56843 ( .A(n49520), .B(n14622), .X(n14600) );
  nor_x1_sg U56844 ( .A(n14623), .B(n14624), .X(n14622) );
  nand_x1_sg U56845 ( .A(n14624), .B(n14623), .X(n14625) );
  nor_x1_sg U56846 ( .A(n49806), .B(n15441), .X(n15419) );
  nor_x1_sg U56847 ( .A(n15442), .B(n15443), .X(n15441) );
  nand_x1_sg U56848 ( .A(n15443), .B(n15442), .X(n15444) );
  nor_x1_sg U56849 ( .A(n50092), .B(n16260), .X(n16238) );
  nor_x1_sg U56850 ( .A(n16261), .B(n16262), .X(n16260) );
  nand_x1_sg U56851 ( .A(n16262), .B(n16261), .X(n16263) );
  nor_x1_sg U56852 ( .A(n50666), .B(n17898), .X(n17876) );
  nor_x1_sg U56853 ( .A(n17899), .B(n17900), .X(n17898) );
  nand_x1_sg U56854 ( .A(n17900), .B(n17899), .X(n17901) );
  nor_x1_sg U56855 ( .A(n50953), .B(n18719), .X(n18697) );
  nor_x1_sg U56856 ( .A(n18720), .B(n18721), .X(n18719) );
  nand_x1_sg U56857 ( .A(n18721), .B(n18720), .X(n18722) );
  nand_x1_sg U56858 ( .A(n16929), .B(n41603), .X(n16933) );
  nand_x1_sg U56859 ( .A(n8123), .B(n47158), .X(n8091) );
  nand_x1_sg U56860 ( .A(n8941), .B(n47443), .X(n8909) );
  nand_x1_sg U56861 ( .A(n9761), .B(n47728), .X(n9729) );
  nand_x1_sg U56862 ( .A(n10580), .B(n48013), .X(n10548) );
  nand_x1_sg U56863 ( .A(n11399), .B(n48298), .X(n11367) );
  nand_x1_sg U56864 ( .A(n12218), .B(n48583), .X(n12186) );
  nand_x1_sg U56865 ( .A(n13037), .B(n48869), .X(n13005) );
  nand_x1_sg U56866 ( .A(n13856), .B(n49156), .X(n13824) );
  nand_x1_sg U56867 ( .A(n14675), .B(n49442), .X(n14643) );
  nand_x1_sg U56868 ( .A(n15494), .B(n49727), .X(n15462) );
  nand_x1_sg U56869 ( .A(n16313), .B(n50014), .X(n16281) );
  nand_x1_sg U56870 ( .A(n17130), .B(n50298), .X(n17097) );
  nand_x1_sg U56871 ( .A(n17951), .B(n50588), .X(n17919) );
  nand_x1_sg U56872 ( .A(n18772), .B(n50875), .X(n18740) );
  nand_x1_sg U56873 ( .A(n6958), .B(n41604), .X(n7469) );
  nand_x1_sg U56874 ( .A(n7305), .B(n46865), .X(n7272) );
  nand_x1_sg U56875 ( .A(n16782), .B(n41603), .X(n17294) );
  nand_x1_sg U56876 ( .A(n7775), .B(n41605), .X(n8287) );
  nand_x1_sg U56877 ( .A(n8593), .B(n41606), .X(n9105) );
  nand_x1_sg U56878 ( .A(n9413), .B(n41607), .X(n9925) );
  nand_x1_sg U56879 ( .A(n10232), .B(n41608), .X(n10744) );
  nand_x1_sg U56880 ( .A(n11051), .B(n41609), .X(n11563) );
  nand_x1_sg U56881 ( .A(n11870), .B(n41610), .X(n12382) );
  nand_x1_sg U56882 ( .A(n12689), .B(n41611), .X(n13201) );
  nand_x1_sg U56883 ( .A(n13508), .B(n41612), .X(n14020) );
  nand_x1_sg U56884 ( .A(n14327), .B(n41613), .X(n14839) );
  nand_x1_sg U56885 ( .A(n15146), .B(n41614), .X(n15658) );
  nand_x1_sg U56886 ( .A(n15965), .B(n41615), .X(n16477) );
  nand_x1_sg U56887 ( .A(n17603), .B(n41616), .X(n18115) );
  nand_x1_sg U56888 ( .A(n18424), .B(n41617), .X(n18936) );
  nand_x1_sg U56889 ( .A(n22943), .B(n41578), .X(n22950) );
  nand_x1_sg U56890 ( .A(n23220), .B(n41577), .X(n23227) );
  nand_x1_sg U56891 ( .A(n23500), .B(n41576), .X(n23507) );
  nand_x1_sg U56892 ( .A(n23779), .B(n41575), .X(n23786) );
  nand_x1_sg U56893 ( .A(n24058), .B(n41582), .X(n24065) );
  nand_x1_sg U56894 ( .A(n24337), .B(n41581), .X(n24344) );
  nand_x1_sg U56895 ( .A(n24616), .B(n41580), .X(n24623) );
  nand_x1_sg U56896 ( .A(n24894), .B(n41579), .X(n24901) );
  nand_x1_sg U56897 ( .A(n25173), .B(n41586), .X(n25180) );
  nand_x1_sg U56898 ( .A(n25452), .B(n41585), .X(n25459) );
  nand_x1_sg U56899 ( .A(n25731), .B(n41584), .X(n25738) );
  nand_x1_sg U56900 ( .A(n25997), .B(n41693), .X(n26003) );
  nand_x1_sg U56901 ( .A(n26284), .B(n41587), .X(n26292) );
  nand_x1_sg U56902 ( .A(n26568), .B(n41583), .X(n26575) );
  nand_x1_sg U56903 ( .A(n22929), .B(n39730), .X(n22936) );
  nand_x1_sg U56904 ( .A(n23206), .B(n39733), .X(n23213) );
  nand_x1_sg U56905 ( .A(n23486), .B(n39736), .X(n23493) );
  nand_x1_sg U56906 ( .A(n23765), .B(n39739), .X(n23772) );
  nand_x1_sg U56907 ( .A(n24044), .B(n39742), .X(n24051) );
  nand_x1_sg U56908 ( .A(n24323), .B(n39745), .X(n24330) );
  nand_x1_sg U56909 ( .A(n24602), .B(n39748), .X(n24609) );
  nand_x1_sg U56910 ( .A(n24880), .B(n39751), .X(n24887) );
  nand_x1_sg U56911 ( .A(n25159), .B(n39754), .X(n25166) );
  nand_x1_sg U56912 ( .A(n25438), .B(n39757), .X(n25445) );
  nand_x1_sg U56913 ( .A(n25717), .B(n39760), .X(n25724) );
  nand_x1_sg U56914 ( .A(n25984), .B(n39603), .X(n25990) );
  nand_x1_sg U56915 ( .A(n26268), .B(n39763), .X(n26276) );
  nand_x1_sg U56916 ( .A(n26554), .B(n39766), .X(n26561) );
  nor_x1_sg U56917 ( .A(n41736), .B(n39035), .X(n8447) );
  nor_x1_sg U56918 ( .A(n41735), .B(n41630), .X(n9265) );
  nor_x1_sg U56919 ( .A(n41734), .B(n41628), .X(n10085) );
  nor_x1_sg U56920 ( .A(n41727), .B(n41626), .X(n10904) );
  nor_x1_sg U56921 ( .A(n41726), .B(n39033), .X(n11723) );
  nor_x1_sg U56922 ( .A(n41730), .B(n39031), .X(n12542) );
  nor_x1_sg U56923 ( .A(n41729), .B(n49055), .X(n13361) );
  nor_x1_sg U56924 ( .A(n41728), .B(n41624), .X(n14180) );
  nor_x1_sg U56925 ( .A(n41731), .B(n39029), .X(n14999) );
  nor_x1_sg U56926 ( .A(n41733), .B(n41621), .X(n15818) );
  nor_x1_sg U56927 ( .A(n41732), .B(n39028), .X(n16637) );
  nor_x1_sg U56928 ( .A(n41738), .B(n41619), .X(n18275) );
  nor_x1_sg U56929 ( .A(n41737), .B(n41620), .X(n19096) );
  nand_x1_sg U56930 ( .A(n22915), .B(n39612), .X(n22922) );
  nand_x1_sg U56931 ( .A(n23192), .B(n39609), .X(n23199) );
  nand_x1_sg U56932 ( .A(n23472), .B(n39626), .X(n23479) );
  nand_x1_sg U56933 ( .A(n23751), .B(n39623), .X(n23758) );
  nand_x1_sg U56934 ( .A(n24030), .B(n39620), .X(n24037) );
  nand_x1_sg U56935 ( .A(n24309), .B(n39617), .X(n24316) );
  nand_x1_sg U56936 ( .A(n24588), .B(n39638), .X(n24595) );
  nand_x1_sg U56937 ( .A(n24866), .B(n39636), .X(n24873) );
  nand_x1_sg U56938 ( .A(n25145), .B(n39633), .X(n25152) );
  nand_x1_sg U56939 ( .A(n25424), .B(n39630), .X(n25431) );
  nand_x1_sg U56940 ( .A(n25703), .B(n39648), .X(n25710) );
  nand_x1_sg U56941 ( .A(n25971), .B(n39614), .X(n25978) );
  nand_x1_sg U56942 ( .A(n26252), .B(n39645), .X(n26260) );
  nand_x1_sg U56943 ( .A(n26540), .B(n39642), .X(n26547) );
  nand_x1_sg U56944 ( .A(n22698), .B(n41983), .X(n22697) );
  nand_x1_sg U56945 ( .A(n22642), .B(n39725), .X(n22656) );
  nor_x1_sg U56946 ( .A(n40242), .B(n41195), .X(n22869) );
  nor_x1_sg U56947 ( .A(n40248), .B(n41187), .X(n23146) );
  nor_x1_sg U56948 ( .A(n40253), .B(n41182), .X(n23426) );
  nor_x1_sg U56949 ( .A(n40258), .B(n39228), .X(n23705) );
  nor_x1_sg U56950 ( .A(n40263), .B(n41174), .X(n23984) );
  nor_x1_sg U56951 ( .A(n40268), .B(n41168), .X(n24263) );
  nor_x1_sg U56952 ( .A(n40273), .B(n39234), .X(n24542) );
  nor_x1_sg U56953 ( .A(n40278), .B(n41869), .X(n24820) );
  nor_x1_sg U56954 ( .A(n40283), .B(n41153), .X(n25099) );
  nor_x1_sg U56955 ( .A(n40288), .B(n41149), .X(n25378) );
  nor_x1_sg U56956 ( .A(n40293), .B(n41144), .X(n25657) );
  nor_x1_sg U56957 ( .A(n40237), .B(n41140), .X(n26199) );
  nor_x1_sg U56958 ( .A(n40298), .B(n41132), .X(n26494) );
  nor_x1_sg U56959 ( .A(n7229), .B(n7230), .X(n7228) );
  nor_x1_sg U56960 ( .A(n17054), .B(n17055), .X(n17053) );
  nor_x1_sg U56961 ( .A(n7236), .B(n7237), .X(n7235) );
  nor_x1_sg U56962 ( .A(n8055), .B(n8056), .X(n8054) );
  nor_x1_sg U56963 ( .A(n8873), .B(n8874), .X(n8872) );
  nor_x1_sg U56964 ( .A(n9693), .B(n9694), .X(n9692) );
  nor_x1_sg U56965 ( .A(n10512), .B(n10513), .X(n10511) );
  nor_x1_sg U56966 ( .A(n11331), .B(n11332), .X(n11330) );
  nor_x1_sg U56967 ( .A(n12150), .B(n12151), .X(n12149) );
  nor_x1_sg U56968 ( .A(n12969), .B(n12970), .X(n12968) );
  nor_x1_sg U56969 ( .A(n13788), .B(n13789), .X(n13787) );
  nor_x1_sg U56970 ( .A(n14607), .B(n14608), .X(n14606) );
  nor_x1_sg U56971 ( .A(n15426), .B(n15427), .X(n15425) );
  nor_x1_sg U56972 ( .A(n16245), .B(n16246), .X(n16244) );
  nor_x1_sg U56973 ( .A(n17061), .B(n17062), .X(n17060) );
  nor_x1_sg U56974 ( .A(n17883), .B(n17884), .X(n17882) );
  nor_x1_sg U56975 ( .A(n18704), .B(n18705), .X(n18703) );
  nor_x1_sg U56976 ( .A(n7144), .B(n7145), .X(n7143) );
  nor_x1_sg U56977 ( .A(n7962), .B(n7963), .X(n7961) );
  nor_x1_sg U56978 ( .A(n8780), .B(n8781), .X(n8779) );
  nor_x1_sg U56979 ( .A(n9600), .B(n9601), .X(n9599) );
  nor_x1_sg U56980 ( .A(n10419), .B(n10420), .X(n10418) );
  nor_x1_sg U56981 ( .A(n11238), .B(n11239), .X(n11237) );
  nor_x1_sg U56982 ( .A(n12057), .B(n12058), .X(n12056) );
  nor_x1_sg U56983 ( .A(n12876), .B(n12877), .X(n12875) );
  nor_x1_sg U56984 ( .A(n13695), .B(n13696), .X(n13694) );
  nor_x1_sg U56985 ( .A(n14514), .B(n14515), .X(n14513) );
  nor_x1_sg U56986 ( .A(n15333), .B(n15334), .X(n15332) );
  nor_x1_sg U56987 ( .A(n16152), .B(n16153), .X(n16151) );
  nor_x1_sg U56988 ( .A(n16969), .B(n16970), .X(n16968) );
  nor_x1_sg U56989 ( .A(n17790), .B(n17791), .X(n17789) );
  nor_x1_sg U56990 ( .A(n18611), .B(n18612), .X(n18610) );
  nor_x1_sg U56991 ( .A(n8133), .B(n8134), .X(n8132) );
  nor_x1_sg U56992 ( .A(n8951), .B(n8952), .X(n8950) );
  nor_x1_sg U56993 ( .A(n9771), .B(n9772), .X(n9770) );
  nor_x1_sg U56994 ( .A(n10590), .B(n10591), .X(n10589) );
  nor_x1_sg U56995 ( .A(n11409), .B(n11410), .X(n11408) );
  nor_x1_sg U56996 ( .A(n12228), .B(n12229), .X(n12227) );
  nor_x1_sg U56997 ( .A(n13047), .B(n13048), .X(n13046) );
  nor_x1_sg U56998 ( .A(n13866), .B(n13867), .X(n13865) );
  nor_x1_sg U56999 ( .A(n14685), .B(n14686), .X(n14684) );
  nor_x1_sg U57000 ( .A(n15504), .B(n15505), .X(n15503) );
  nor_x1_sg U57001 ( .A(n16323), .B(n16324), .X(n16322) );
  nor_x1_sg U57002 ( .A(n17961), .B(n17962), .X(n17960) );
  nor_x1_sg U57003 ( .A(n18782), .B(n18783), .X(n18781) );
  nor_x1_sg U57004 ( .A(n8083), .B(n8084), .X(n8082) );
  nor_x1_sg U57005 ( .A(n8901), .B(n8902), .X(n8900) );
  nor_x1_sg U57006 ( .A(n9721), .B(n9722), .X(n9720) );
  nor_x1_sg U57007 ( .A(n10540), .B(n10541), .X(n10539) );
  nor_x1_sg U57008 ( .A(n11359), .B(n11360), .X(n11358) );
  nor_x1_sg U57009 ( .A(n12178), .B(n12179), .X(n12177) );
  nor_x1_sg U57010 ( .A(n12997), .B(n12998), .X(n12996) );
  nor_x1_sg U57011 ( .A(n13816), .B(n13817), .X(n13815) );
  nor_x1_sg U57012 ( .A(n14635), .B(n14636), .X(n14634) );
  nor_x1_sg U57013 ( .A(n15454), .B(n15455), .X(n15453) );
  nor_x1_sg U57014 ( .A(n16273), .B(n16274), .X(n16272) );
  nor_x1_sg U57015 ( .A(n17911), .B(n17912), .X(n17910) );
  nor_x1_sg U57016 ( .A(n18732), .B(n18733), .X(n18731) );
  nor_x1_sg U57017 ( .A(n7291), .B(n7292), .X(n7290) );
  nor_x1_sg U57018 ( .A(n7416), .B(n7417), .X(n7415) );
  nor_x1_sg U57019 ( .A(n8109), .B(n8110), .X(n8108) );
  nor_x1_sg U57020 ( .A(n8234), .B(n8235), .X(n8233) );
  nor_x1_sg U57021 ( .A(n8927), .B(n8928), .X(n8926) );
  nor_x1_sg U57022 ( .A(n9052), .B(n9053), .X(n9051) );
  nor_x1_sg U57023 ( .A(n9747), .B(n9748), .X(n9746) );
  nor_x1_sg U57024 ( .A(n9872), .B(n9873), .X(n9871) );
  nor_x1_sg U57025 ( .A(n10566), .B(n10567), .X(n10565) );
  nor_x1_sg U57026 ( .A(n10691), .B(n10692), .X(n10690) );
  nor_x1_sg U57027 ( .A(n11385), .B(n11386), .X(n11384) );
  nor_x1_sg U57028 ( .A(n11510), .B(n11511), .X(n11509) );
  nor_x1_sg U57029 ( .A(n12204), .B(n12205), .X(n12203) );
  nor_x1_sg U57030 ( .A(n12329), .B(n12330), .X(n12328) );
  nor_x1_sg U57031 ( .A(n13023), .B(n13024), .X(n13022) );
  nor_x1_sg U57032 ( .A(n13148), .B(n13149), .X(n13147) );
  nor_x1_sg U57033 ( .A(n13842), .B(n13843), .X(n13841) );
  nor_x1_sg U57034 ( .A(n13967), .B(n13968), .X(n13966) );
  nor_x1_sg U57035 ( .A(n14661), .B(n14662), .X(n14660) );
  nor_x1_sg U57036 ( .A(n14786), .B(n14787), .X(n14785) );
  nor_x1_sg U57037 ( .A(n15480), .B(n15481), .X(n15479) );
  nor_x1_sg U57038 ( .A(n15605), .B(n15606), .X(n15604) );
  nor_x1_sg U57039 ( .A(n16299), .B(n16300), .X(n16298) );
  nor_x1_sg U57040 ( .A(n16424), .B(n16425), .X(n16423) );
  nor_x1_sg U57041 ( .A(n17116), .B(n17117), .X(n17115) );
  nor_x1_sg U57042 ( .A(n17241), .B(n17242), .X(n17240) );
  nor_x1_sg U57043 ( .A(n17937), .B(n17938), .X(n17936) );
  nor_x1_sg U57044 ( .A(n18062), .B(n18063), .X(n18061) );
  nor_x1_sg U57045 ( .A(n18758), .B(n18759), .X(n18757) );
  nor_x1_sg U57046 ( .A(n18883), .B(n18884), .X(n18882) );
  nor_x1_sg U57047 ( .A(n7199), .B(n7200), .X(n7198) );
  nor_x1_sg U57048 ( .A(n8018), .B(n8019), .X(n8017) );
  nor_x1_sg U57049 ( .A(n8836), .B(n8837), .X(n8835) );
  nor_x1_sg U57050 ( .A(n9656), .B(n9657), .X(n9655) );
  nor_x1_sg U57051 ( .A(n10475), .B(n10476), .X(n10474) );
  nor_x1_sg U57052 ( .A(n11294), .B(n11295), .X(n11293) );
  nor_x1_sg U57053 ( .A(n12113), .B(n12114), .X(n12112) );
  nor_x1_sg U57054 ( .A(n12932), .B(n12933), .X(n12931) );
  nor_x1_sg U57055 ( .A(n13751), .B(n13752), .X(n13750) );
  nor_x1_sg U57056 ( .A(n14570), .B(n14571), .X(n14569) );
  nor_x1_sg U57057 ( .A(n15389), .B(n15390), .X(n15388) );
  nor_x1_sg U57058 ( .A(n16208), .B(n16209), .X(n16207) );
  nor_x1_sg U57059 ( .A(n17024), .B(n17025), .X(n17023) );
  nor_x1_sg U57060 ( .A(n17846), .B(n17847), .X(n17845) );
  nor_x1_sg U57061 ( .A(n18667), .B(n18668), .X(n18666) );
  nor_x1_sg U57062 ( .A(n47053), .B(n7616), .X(n7615) );
  nor_x1_sg U57063 ( .A(n47340), .B(n8434), .X(n8433) );
  nor_x1_sg U57064 ( .A(n47625), .B(n9252), .X(n9251) );
  nor_x1_sg U57065 ( .A(n47910), .B(n10072), .X(n10071) );
  nor_x1_sg U57066 ( .A(n48195), .B(n10891), .X(n10890) );
  nor_x1_sg U57067 ( .A(n48480), .B(n11710), .X(n11709) );
  nor_x1_sg U57068 ( .A(n48765), .B(n12529), .X(n12528) );
  nor_x1_sg U57069 ( .A(n49051), .B(n13348), .X(n13347) );
  nor_x1_sg U57070 ( .A(n49338), .B(n14167), .X(n14166) );
  nor_x1_sg U57071 ( .A(n49624), .B(n14986), .X(n14985) );
  nor_x1_sg U57072 ( .A(n49910), .B(n15805), .X(n15804) );
  nor_x1_sg U57073 ( .A(n50196), .B(n16624), .X(n16623) );
  nor_x1_sg U57074 ( .A(n50481), .B(n17441), .X(n17440) );
  nor_x1_sg U57075 ( .A(n50770), .B(n18262), .X(n18261) );
  nor_x1_sg U57076 ( .A(n51057), .B(n19083), .X(n19082) );
  nand_x1_sg U57077 ( .A(n7566), .B(n7565), .X(n7563) );
  nor_x1_sg U57078 ( .A(n7565), .B(n7566), .X(n7564) );
  nand_x1_sg U57079 ( .A(n17391), .B(n17390), .X(n17388) );
  nor_x1_sg U57080 ( .A(n17390), .B(n17391), .X(n17389) );
  nand_x1_sg U57081 ( .A(n8384), .B(n8383), .X(n8381) );
  nor_x1_sg U57082 ( .A(n8383), .B(n8384), .X(n8382) );
  nand_x1_sg U57083 ( .A(n9202), .B(n9201), .X(n9199) );
  nor_x1_sg U57084 ( .A(n9201), .B(n9202), .X(n9200) );
  nand_x1_sg U57085 ( .A(n10022), .B(n10021), .X(n10019) );
  nor_x1_sg U57086 ( .A(n10021), .B(n10022), .X(n10020) );
  nand_x1_sg U57087 ( .A(n10841), .B(n10840), .X(n10838) );
  nor_x1_sg U57088 ( .A(n10840), .B(n10841), .X(n10839) );
  nand_x1_sg U57089 ( .A(n11660), .B(n11659), .X(n11657) );
  nor_x1_sg U57090 ( .A(n11659), .B(n11660), .X(n11658) );
  nand_x1_sg U57091 ( .A(n12479), .B(n12478), .X(n12476) );
  nor_x1_sg U57092 ( .A(n12478), .B(n12479), .X(n12477) );
  nand_x1_sg U57093 ( .A(n13298), .B(n13297), .X(n13295) );
  nor_x1_sg U57094 ( .A(n13297), .B(n13298), .X(n13296) );
  nand_x1_sg U57095 ( .A(n14117), .B(n14116), .X(n14114) );
  nor_x1_sg U57096 ( .A(n14116), .B(n14117), .X(n14115) );
  nand_x1_sg U57097 ( .A(n14936), .B(n14935), .X(n14933) );
  nor_x1_sg U57098 ( .A(n14935), .B(n14936), .X(n14934) );
  nand_x1_sg U57099 ( .A(n15755), .B(n15754), .X(n15752) );
  nor_x1_sg U57100 ( .A(n15754), .B(n15755), .X(n15753) );
  nand_x1_sg U57101 ( .A(n16574), .B(n16573), .X(n16571) );
  nor_x1_sg U57102 ( .A(n16573), .B(n16574), .X(n16572) );
  nand_x1_sg U57103 ( .A(n18212), .B(n18211), .X(n18209) );
  nor_x1_sg U57104 ( .A(n18211), .B(n18212), .X(n18210) );
  nand_x1_sg U57105 ( .A(n19033), .B(n19032), .X(n19030) );
  nor_x1_sg U57106 ( .A(n19032), .B(n19033), .X(n19031) );
  nand_x1_sg U57107 ( .A(n17112), .B(n17113), .X(n17111) );
  nor_x1_sg U57108 ( .A(n17113), .B(n17112), .X(n17114) );
  nor_x1_sg U57109 ( .A(n39850), .B(n41304), .X(n22645) );
  nand_x1_sg U57110 ( .A(n40227), .B(n41193), .X(n22982) );
  nand_x1_sg U57111 ( .A(n39477), .B(n41175), .X(n24097) );
  nand_x1_sg U57112 ( .A(n41463), .B(n40486), .X(n24376) );
  nand_x1_sg U57113 ( .A(n40226), .B(n41165), .X(n24655) );
  nand_x1_sg U57114 ( .A(n40226), .B(n40478), .X(n24933) );
  nand_x1_sg U57115 ( .A(n40218), .B(n41155), .X(n25212) );
  nand_x1_sg U57116 ( .A(n39276), .B(n41147), .X(n25491) );
  nand_x1_sg U57117 ( .A(n41461), .B(n41142), .X(n25770) );
  nand_x1_sg U57118 ( .A(n41311), .B(n40458), .X(n26607) );
  nand_x1_sg U57119 ( .A(n39476), .B(n41188), .X(n23259) );
  nand_x1_sg U57120 ( .A(n39477), .B(n41185), .X(n23539) );
  nand_x1_sg U57121 ( .A(n40218), .B(n41178), .X(n23818) );
  nand_x1_sg U57122 ( .A(n39657), .B(n41137), .X(n26327) );
  nand_x1_sg U57123 ( .A(n6847), .B(n6848), .X(n7069) );
  nand_x1_sg U57124 ( .A(n7664), .B(n7665), .X(n7887) );
  nand_x1_sg U57125 ( .A(n8482), .B(n8483), .X(n8705) );
  nand_x1_sg U57126 ( .A(n9302), .B(n9303), .X(n9525) );
  nand_x1_sg U57127 ( .A(n10121), .B(n10122), .X(n10344) );
  nand_x1_sg U57128 ( .A(n10940), .B(n10941), .X(n11163) );
  nand_x1_sg U57129 ( .A(n11759), .B(n11760), .X(n11982) );
  nand_x1_sg U57130 ( .A(n12578), .B(n12579), .X(n12801) );
  nand_x1_sg U57131 ( .A(n13397), .B(n13398), .X(n13620) );
  nand_x1_sg U57132 ( .A(n14216), .B(n14217), .X(n14439) );
  nand_x1_sg U57133 ( .A(n15035), .B(n15036), .X(n15258) );
  nand_x1_sg U57134 ( .A(n15854), .B(n15855), .X(n16077) );
  nand_x1_sg U57135 ( .A(n17492), .B(n17493), .X(n17715) );
  nand_x1_sg U57136 ( .A(n18313), .B(n18314), .X(n18536) );
  nand_x1_sg U57137 ( .A(n16671), .B(n16672), .X(n16896) );
  nand_x1_sg U57138 ( .A(n7823), .B(n7949), .X(n8207) );
  nand_x1_sg U57139 ( .A(n8641), .B(n8767), .X(n9025) );
  nand_x1_sg U57140 ( .A(n9461), .B(n9587), .X(n9845) );
  nand_x1_sg U57141 ( .A(n10280), .B(n10406), .X(n10664) );
  nand_x1_sg U57142 ( .A(n11099), .B(n11225), .X(n11483) );
  nand_x1_sg U57143 ( .A(n11918), .B(n12044), .X(n12302) );
  nand_x1_sg U57144 ( .A(n12737), .B(n12863), .X(n13121) );
  nand_x1_sg U57145 ( .A(n13556), .B(n13682), .X(n13940) );
  nand_x1_sg U57146 ( .A(n14375), .B(n14501), .X(n14759) );
  nand_x1_sg U57147 ( .A(n15194), .B(n15320), .X(n15578) );
  nand_x1_sg U57148 ( .A(n16013), .B(n16139), .X(n16397) );
  nand_x1_sg U57149 ( .A(n17651), .B(n17777), .X(n18035) );
  nand_x1_sg U57150 ( .A(n18472), .B(n18598), .X(n18856) );
  nand_x1_sg U57151 ( .A(n8199), .B(n41605), .X(n8152) );
  nand_x1_sg U57152 ( .A(n9017), .B(n41606), .X(n8970) );
  nand_x1_sg U57153 ( .A(n9837), .B(n41607), .X(n9790) );
  nand_x1_sg U57154 ( .A(n10656), .B(n41608), .X(n10609) );
  nand_x1_sg U57155 ( .A(n11475), .B(n41609), .X(n11428) );
  nand_x1_sg U57156 ( .A(n12294), .B(n41610), .X(n12247) );
  nand_x1_sg U57157 ( .A(n13113), .B(n41611), .X(n13066) );
  nand_x1_sg U57158 ( .A(n13932), .B(n41612), .X(n13885) );
  nand_x1_sg U57159 ( .A(n14751), .B(n41613), .X(n14704) );
  nand_x1_sg U57160 ( .A(n15570), .B(n41614), .X(n15523) );
  nand_x1_sg U57161 ( .A(n16389), .B(n41615), .X(n16342) );
  nand_x1_sg U57162 ( .A(n17206), .B(n41603), .X(n17159) );
  nand_x1_sg U57163 ( .A(n18027), .B(n41616), .X(n17980) );
  nand_x1_sg U57164 ( .A(n18848), .B(n41617), .X(n18801) );
  nand_x1_sg U57165 ( .A(n17205), .B(n17042), .X(n17203) );
  nor_x1_sg U57166 ( .A(n17042), .B(n17205), .X(n17204) );
  nor_x1_sg U57167 ( .A(n41948), .B(n41808), .X(n22607) );
  nand_x1_sg U57168 ( .A(n46957), .B(n7333), .X(n7372) );
  nand_x1_sg U57169 ( .A(n46939), .B(n7374), .X(n7373) );
  nand_x1_sg U57170 ( .A(n47248), .B(n8151), .X(n8190) );
  nand_x1_sg U57171 ( .A(n47230), .B(n8192), .X(n8191) );
  nand_x1_sg U57172 ( .A(n47533), .B(n8969), .X(n9008) );
  nand_x1_sg U57173 ( .A(n47515), .B(n9010), .X(n9009) );
  nand_x1_sg U57174 ( .A(n47818), .B(n9789), .X(n9828) );
  nand_x1_sg U57175 ( .A(n47800), .B(n9830), .X(n9829) );
  nand_x1_sg U57176 ( .A(n48103), .B(n10608), .X(n10647) );
  nand_x1_sg U57177 ( .A(n48085), .B(n10649), .X(n10648) );
  nand_x1_sg U57178 ( .A(n48388), .B(n11427), .X(n11466) );
  nand_x1_sg U57179 ( .A(n48370), .B(n11468), .X(n11467) );
  nand_x1_sg U57180 ( .A(n48673), .B(n12246), .X(n12285) );
  nand_x1_sg U57181 ( .A(n48655), .B(n12287), .X(n12286) );
  nand_x1_sg U57182 ( .A(n48959), .B(n13065), .X(n13104) );
  nand_x1_sg U57183 ( .A(n48941), .B(n13106), .X(n13105) );
  nand_x1_sg U57184 ( .A(n49246), .B(n13884), .X(n13923) );
  nand_x1_sg U57185 ( .A(n49228), .B(n13925), .X(n13924) );
  nand_x1_sg U57186 ( .A(n49532), .B(n14703), .X(n14742) );
  nand_x1_sg U57187 ( .A(n49514), .B(n14744), .X(n14743) );
  nand_x1_sg U57188 ( .A(n49818), .B(n15522), .X(n15561) );
  nand_x1_sg U57189 ( .A(n49800), .B(n15563), .X(n15562) );
  nand_x1_sg U57190 ( .A(n50104), .B(n16341), .X(n16380) );
  nand_x1_sg U57191 ( .A(n50086), .B(n16382), .X(n16381) );
  nand_x1_sg U57192 ( .A(n50678), .B(n17979), .X(n18018) );
  nand_x1_sg U57193 ( .A(n50660), .B(n18020), .X(n18019) );
  nand_x1_sg U57194 ( .A(n50965), .B(n18800), .X(n18839) );
  nand_x1_sg U57195 ( .A(n50947), .B(n18841), .X(n18840) );
  nand_x1_sg U57196 ( .A(n50447), .B(n17247), .X(n17245) );
  nor_x1_sg U57197 ( .A(n17247), .B(n50447), .X(n17246) );
  nand_x1_sg U57198 ( .A(n46936), .B(n46958), .X(n7395) );
  nand_x1_sg U57199 ( .A(n7396), .B(n7397), .X(n7394) );
  nand_x1_sg U57200 ( .A(n47228), .B(n47249), .X(n8213) );
  nand_x1_sg U57201 ( .A(n8214), .B(n8215), .X(n8212) );
  nand_x1_sg U57202 ( .A(n47513), .B(n47534), .X(n9031) );
  nand_x1_sg U57203 ( .A(n9032), .B(n9033), .X(n9030) );
  nand_x1_sg U57204 ( .A(n47798), .B(n47819), .X(n9851) );
  nand_x1_sg U57205 ( .A(n9852), .B(n9853), .X(n9850) );
  nand_x1_sg U57206 ( .A(n48083), .B(n48104), .X(n10670) );
  nand_x1_sg U57207 ( .A(n10671), .B(n10672), .X(n10669) );
  nand_x1_sg U57208 ( .A(n48368), .B(n48389), .X(n11489) );
  nand_x1_sg U57209 ( .A(n11490), .B(n11491), .X(n11488) );
  nand_x1_sg U57210 ( .A(n48653), .B(n48674), .X(n12308) );
  nand_x1_sg U57211 ( .A(n12309), .B(n12310), .X(n12307) );
  nand_x1_sg U57212 ( .A(n48939), .B(n48960), .X(n13127) );
  nand_x1_sg U57213 ( .A(n13128), .B(n13129), .X(n13126) );
  nand_x1_sg U57214 ( .A(n49226), .B(n49247), .X(n13946) );
  nand_x1_sg U57215 ( .A(n13947), .B(n13948), .X(n13945) );
  nand_x1_sg U57216 ( .A(n49512), .B(n49533), .X(n14765) );
  nand_x1_sg U57217 ( .A(n14766), .B(n14767), .X(n14764) );
  nand_x1_sg U57218 ( .A(n49798), .B(n49819), .X(n15584) );
  nand_x1_sg U57219 ( .A(n15585), .B(n15586), .X(n15583) );
  nand_x1_sg U57220 ( .A(n50084), .B(n50105), .X(n16403) );
  nand_x1_sg U57221 ( .A(n16404), .B(n16405), .X(n16402) );
  nand_x1_sg U57222 ( .A(n50658), .B(n50679), .X(n18041) );
  nand_x1_sg U57223 ( .A(n18042), .B(n18043), .X(n18040) );
  nand_x1_sg U57224 ( .A(n50945), .B(n50966), .X(n18862) );
  nand_x1_sg U57225 ( .A(n18863), .B(n18864), .X(n18861) );
  nand_x1_sg U57226 ( .A(n46968), .B(n46939), .X(n7376) );
  nand_x1_sg U57227 ( .A(n7374), .B(n7377), .X(n7375) );
  nand_x1_sg U57228 ( .A(n47258), .B(n47230), .X(n8194) );
  nand_x1_sg U57229 ( .A(n8192), .B(n8195), .X(n8193) );
  nand_x1_sg U57230 ( .A(n47543), .B(n47515), .X(n9012) );
  nand_x1_sg U57231 ( .A(n9010), .B(n9013), .X(n9011) );
  nand_x1_sg U57232 ( .A(n47828), .B(n47800), .X(n9832) );
  nand_x1_sg U57233 ( .A(n9830), .B(n9833), .X(n9831) );
  nand_x1_sg U57234 ( .A(n48113), .B(n48085), .X(n10651) );
  nand_x1_sg U57235 ( .A(n10649), .B(n10652), .X(n10650) );
  nand_x1_sg U57236 ( .A(n48398), .B(n48370), .X(n11470) );
  nand_x1_sg U57237 ( .A(n11468), .B(n11471), .X(n11469) );
  nand_x1_sg U57238 ( .A(n48683), .B(n48655), .X(n12289) );
  nand_x1_sg U57239 ( .A(n12287), .B(n12290), .X(n12288) );
  nand_x1_sg U57240 ( .A(n48969), .B(n48941), .X(n13108) );
  nand_x1_sg U57241 ( .A(n13106), .B(n13109), .X(n13107) );
  nand_x1_sg U57242 ( .A(n49256), .B(n49228), .X(n13927) );
  nand_x1_sg U57243 ( .A(n13925), .B(n13928), .X(n13926) );
  nand_x1_sg U57244 ( .A(n49542), .B(n49514), .X(n14746) );
  nand_x1_sg U57245 ( .A(n14744), .B(n14747), .X(n14745) );
  nand_x1_sg U57246 ( .A(n49828), .B(n49800), .X(n15565) );
  nand_x1_sg U57247 ( .A(n15563), .B(n15566), .X(n15564) );
  nand_x1_sg U57248 ( .A(n50114), .B(n50086), .X(n16384) );
  nand_x1_sg U57249 ( .A(n16382), .B(n16385), .X(n16383) );
  nand_x1_sg U57250 ( .A(n50688), .B(n50660), .X(n18022) );
  nand_x1_sg U57251 ( .A(n18020), .B(n18023), .X(n18021) );
  nand_x1_sg U57252 ( .A(n50975), .B(n50947), .X(n18843) );
  nand_x1_sg U57253 ( .A(n18841), .B(n18844), .X(n18842) );
  nand_x1_sg U57254 ( .A(n50399), .B(n50371), .X(n17201) );
  nand_x1_sg U57255 ( .A(n17199), .B(n17202), .X(n17200) );
  nand_x1_sg U57256 ( .A(n50369), .B(n50390), .X(n17220) );
  nand_x1_sg U57257 ( .A(n17221), .B(n17222), .X(n17219) );
  nand_x1_sg U57258 ( .A(n7381), .B(n41604), .X(n7334) );
  nand_x1_sg U57259 ( .A(n7611), .B(n7612), .X(n7610) );
  nor_x1_sg U57260 ( .A(n7612), .B(n7611), .X(n7613) );
  nand_x1_sg U57261 ( .A(n17436), .B(n17437), .X(n17435) );
  nor_x1_sg U57262 ( .A(n17437), .B(n17436), .X(n17438) );
  nand_x1_sg U57263 ( .A(n17256), .B(n17257), .X(n17255) );
  nor_x1_sg U57264 ( .A(n17257), .B(n17256), .X(n17258) );
  nand_x1_sg U57265 ( .A(n7114), .B(n7116), .X(n7122) );
  nand_x1_sg U57266 ( .A(n7932), .B(n7934), .X(n7940) );
  nand_x1_sg U57267 ( .A(n8750), .B(n8752), .X(n8758) );
  nand_x1_sg U57268 ( .A(n9570), .B(n9572), .X(n9578) );
  nand_x1_sg U57269 ( .A(n10389), .B(n10391), .X(n10397) );
  nand_x1_sg U57270 ( .A(n11208), .B(n11210), .X(n11216) );
  nand_x1_sg U57271 ( .A(n12027), .B(n12029), .X(n12035) );
  nand_x1_sg U57272 ( .A(n12846), .B(n12848), .X(n12854) );
  nand_x1_sg U57273 ( .A(n13665), .B(n13667), .X(n13673) );
  nand_x1_sg U57274 ( .A(n14484), .B(n14486), .X(n14492) );
  nand_x1_sg U57275 ( .A(n15303), .B(n15305), .X(n15311) );
  nand_x1_sg U57276 ( .A(n16122), .B(n16124), .X(n16130) );
  nand_x1_sg U57277 ( .A(n16939), .B(n16941), .X(n16947) );
  nand_x1_sg U57278 ( .A(n17760), .B(n17762), .X(n17768) );
  nand_x1_sg U57279 ( .A(n18581), .B(n18583), .X(n18589) );
  nor_x1_sg U57280 ( .A(n22696), .B(n47099), .X(n22695) );
  inv_x1_sg U57281 ( .A(n22697), .X(n47099) );
  nor_x1_sg U57282 ( .A(n22698), .B(n41983), .X(n22696) );
  nor_x1_sg U57283 ( .A(n22971), .B(n47385), .X(n22970) );
  nor_x1_sg U57284 ( .A(n22972), .B(n41984), .X(n22971) );
  nor_x1_sg U57285 ( .A(n23248), .B(n47670), .X(n23247) );
  nor_x1_sg U57286 ( .A(n23249), .B(n41985), .X(n23248) );
  nor_x1_sg U57287 ( .A(n23528), .B(n47955), .X(n23527) );
  nor_x1_sg U57288 ( .A(n23529), .B(n41979), .X(n23528) );
  nor_x1_sg U57289 ( .A(n23807), .B(n48240), .X(n23806) );
  nor_x1_sg U57290 ( .A(n23808), .B(n41980), .X(n23807) );
  nor_x1_sg U57291 ( .A(n24086), .B(n48525), .X(n24085) );
  nor_x1_sg U57292 ( .A(n24087), .B(n41981), .X(n24086) );
  nor_x1_sg U57293 ( .A(n24365), .B(n48810), .X(n24364) );
  nor_x1_sg U57294 ( .A(n24366), .B(n41982), .X(n24365) );
  nor_x1_sg U57295 ( .A(n24644), .B(n49097), .X(n24643) );
  nor_x1_sg U57296 ( .A(n24645), .B(n41975), .X(n24644) );
  nor_x1_sg U57297 ( .A(n24922), .B(n49383), .X(n24921) );
  nor_x1_sg U57298 ( .A(n24923), .B(n41976), .X(n24922) );
  nor_x1_sg U57299 ( .A(n25201), .B(n49669), .X(n25200) );
  nor_x1_sg U57300 ( .A(n25202), .B(n41977), .X(n25201) );
  nor_x1_sg U57301 ( .A(n25480), .B(n49955), .X(n25479) );
  nor_x1_sg U57302 ( .A(n25481), .B(n41978), .X(n25480) );
  nor_x1_sg U57303 ( .A(n25759), .B(n50241), .X(n25758) );
  nor_x1_sg U57304 ( .A(n25760), .B(n41972), .X(n25759) );
  nor_x1_sg U57305 ( .A(n26316), .B(n50815), .X(n26315) );
  nor_x1_sg U57306 ( .A(n26317), .B(n41973), .X(n26316) );
  nor_x1_sg U57307 ( .A(n26596), .B(n51102), .X(n26595) );
  nor_x1_sg U57308 ( .A(n26597), .B(n41974), .X(n26596) );
  nand_x1_sg U57309 ( .A(n46958), .B(n7396), .X(n7429) );
  nand_x1_sg U57310 ( .A(n46940), .B(n7141), .X(n7428) );
  nand_x1_sg U57311 ( .A(n47249), .B(n8214), .X(n8247) );
  nand_x1_sg U57312 ( .A(n47231), .B(n7959), .X(n8246) );
  nand_x1_sg U57313 ( .A(n47534), .B(n9032), .X(n9065) );
  nand_x1_sg U57314 ( .A(n47516), .B(n8777), .X(n9064) );
  nand_x1_sg U57315 ( .A(n47819), .B(n9852), .X(n9885) );
  nand_x1_sg U57316 ( .A(n47801), .B(n9597), .X(n9884) );
  nand_x1_sg U57317 ( .A(n48104), .B(n10671), .X(n10704) );
  nand_x1_sg U57318 ( .A(n48086), .B(n10416), .X(n10703) );
  nand_x1_sg U57319 ( .A(n48389), .B(n11490), .X(n11523) );
  nand_x1_sg U57320 ( .A(n48371), .B(n11235), .X(n11522) );
  nand_x1_sg U57321 ( .A(n48674), .B(n12309), .X(n12342) );
  nand_x1_sg U57322 ( .A(n48656), .B(n12054), .X(n12341) );
  nand_x1_sg U57323 ( .A(n48960), .B(n13128), .X(n13161) );
  nand_x1_sg U57324 ( .A(n48942), .B(n12873), .X(n13160) );
  nand_x1_sg U57325 ( .A(n49247), .B(n13947), .X(n13980) );
  nand_x1_sg U57326 ( .A(n49229), .B(n13692), .X(n13979) );
  nand_x1_sg U57327 ( .A(n49533), .B(n14766), .X(n14799) );
  nand_x1_sg U57328 ( .A(n49515), .B(n14511), .X(n14798) );
  nand_x1_sg U57329 ( .A(n49819), .B(n15585), .X(n15618) );
  nand_x1_sg U57330 ( .A(n49801), .B(n15330), .X(n15617) );
  nand_x1_sg U57331 ( .A(n50105), .B(n16404), .X(n16437) );
  nand_x1_sg U57332 ( .A(n50087), .B(n16149), .X(n16436) );
  nand_x1_sg U57333 ( .A(n50679), .B(n18042), .X(n18075) );
  nand_x1_sg U57334 ( .A(n50661), .B(n17787), .X(n18074) );
  nand_x1_sg U57335 ( .A(n50966), .B(n18863), .X(n18896) );
  nand_x1_sg U57336 ( .A(n50948), .B(n18608), .X(n18895) );
  nand_x1_sg U57337 ( .A(n47086), .B(n7512), .X(n7517) );
  inv_x1_sg U57338 ( .A(n7511), .X(n47086) );
  nand_x1_sg U57339 ( .A(n47372), .B(n8330), .X(n8335) );
  inv_x1_sg U57340 ( .A(n8329), .X(n47372) );
  nand_x1_sg U57341 ( .A(n47657), .B(n9148), .X(n9153) );
  inv_x1_sg U57342 ( .A(n9147), .X(n47657) );
  nand_x1_sg U57343 ( .A(n47942), .B(n9968), .X(n9973) );
  inv_x1_sg U57344 ( .A(n9967), .X(n47942) );
  nand_x1_sg U57345 ( .A(n48227), .B(n10787), .X(n10792) );
  inv_x1_sg U57346 ( .A(n10786), .X(n48227) );
  nand_x1_sg U57347 ( .A(n48512), .B(n11606), .X(n11611) );
  inv_x1_sg U57348 ( .A(n11605), .X(n48512) );
  nand_x1_sg U57349 ( .A(n48797), .B(n12425), .X(n12430) );
  inv_x1_sg U57350 ( .A(n12424), .X(n48797) );
  nand_x1_sg U57351 ( .A(n49084), .B(n13244), .X(n13249) );
  inv_x1_sg U57352 ( .A(n13243), .X(n49084) );
  nand_x1_sg U57353 ( .A(n49370), .B(n14063), .X(n14068) );
  inv_x1_sg U57354 ( .A(n14062), .X(n49370) );
  nand_x1_sg U57355 ( .A(n49656), .B(n14882), .X(n14887) );
  inv_x1_sg U57356 ( .A(n14881), .X(n49656) );
  nand_x1_sg U57357 ( .A(n49942), .B(n15701), .X(n15706) );
  inv_x1_sg U57358 ( .A(n15700), .X(n49942) );
  nand_x1_sg U57359 ( .A(n50228), .B(n16520), .X(n16525) );
  inv_x1_sg U57360 ( .A(n16519), .X(n50228) );
  nand_x1_sg U57361 ( .A(n50513), .B(n17337), .X(n17342) );
  inv_x1_sg U57362 ( .A(n17336), .X(n50513) );
  nand_x1_sg U57363 ( .A(n50802), .B(n18158), .X(n18163) );
  inv_x1_sg U57364 ( .A(n18157), .X(n50802) );
  nand_x1_sg U57365 ( .A(n51089), .B(n18979), .X(n18984) );
  inv_x1_sg U57366 ( .A(n18978), .X(n51089) );
  inv_x1_sg U57367 ( .A(n6889), .X(n46979) );
  inv_x1_sg U57368 ( .A(n7706), .X(n47269) );
  inv_x1_sg U57369 ( .A(n8524), .X(n47554) );
  inv_x1_sg U57370 ( .A(n9344), .X(n47839) );
  inv_x1_sg U57371 ( .A(n10163), .X(n48124) );
  inv_x1_sg U57372 ( .A(n10982), .X(n48409) );
  inv_x1_sg U57373 ( .A(n11801), .X(n48694) );
  inv_x1_sg U57374 ( .A(n12620), .X(n48980) );
  inv_x1_sg U57375 ( .A(n13439), .X(n49267) );
  inv_x1_sg U57376 ( .A(n14258), .X(n49553) );
  inv_x1_sg U57377 ( .A(n15077), .X(n49839) );
  inv_x1_sg U57378 ( .A(n15896), .X(n50125) );
  inv_x1_sg U57379 ( .A(n17534), .X(n50699) );
  inv_x1_sg U57380 ( .A(n18355), .X(n50986) );
  nand_x1_sg U57381 ( .A(n47351), .B(n39563), .X(n8277) );
  nand_x1_sg U57382 ( .A(n47636), .B(n39566), .X(n9095) );
  nand_x1_sg U57383 ( .A(n47921), .B(n39570), .X(n9915) );
  nand_x1_sg U57384 ( .A(n48206), .B(n39572), .X(n10734) );
  nand_x1_sg U57385 ( .A(n48491), .B(n39575), .X(n11553) );
  nand_x1_sg U57386 ( .A(n48776), .B(n39579), .X(n12372) );
  nand_x1_sg U57387 ( .A(n49063), .B(n39581), .X(n13191) );
  nand_x1_sg U57388 ( .A(n49349), .B(n39584), .X(n14010) );
  nand_x1_sg U57389 ( .A(n49635), .B(n39588), .X(n14829) );
  nand_x1_sg U57390 ( .A(n49921), .B(n39590), .X(n15648) );
  nand_x1_sg U57391 ( .A(n50207), .B(n39593), .X(n16467) );
  nand_x1_sg U57392 ( .A(n50492), .B(n39561), .X(n17284) );
  nand_x1_sg U57393 ( .A(n50781), .B(n39600), .X(n18105) );
  nand_x1_sg U57394 ( .A(n51068), .B(n39597), .X(n18926) );
  nand_x1_sg U57395 ( .A(n47065), .B(n39851), .X(n7459) );
  inv_x1_sg U57396 ( .A(n7120), .X(n46910) );
  inv_x1_sg U57397 ( .A(n7938), .X(n47203) );
  inv_x1_sg U57398 ( .A(n8756), .X(n47488) );
  inv_x1_sg U57399 ( .A(n9576), .X(n47773) );
  inv_x1_sg U57400 ( .A(n10395), .X(n48058) );
  inv_x1_sg U57401 ( .A(n11214), .X(n48343) );
  inv_x1_sg U57402 ( .A(n12033), .X(n48628) );
  inv_x1_sg U57403 ( .A(n12852), .X(n48914) );
  inv_x1_sg U57404 ( .A(n13671), .X(n49201) );
  inv_x1_sg U57405 ( .A(n14490), .X(n49487) );
  inv_x1_sg U57406 ( .A(n15309), .X(n49773) );
  inv_x1_sg U57407 ( .A(n16128), .X(n50059) );
  inv_x1_sg U57408 ( .A(n16945), .X(n50344) );
  inv_x1_sg U57409 ( .A(n17766), .X(n50633) );
  inv_x1_sg U57410 ( .A(n18587), .X(n50920) );
  inv_x1_sg U57411 ( .A(n16999), .X(n50382) );
  nand_x1_sg U57412 ( .A(n7030), .B(n7029), .X(n7594) );
  nor_x1_sg U57413 ( .A(n7029), .B(n7030), .X(n7595) );
  nand_x1_sg U57414 ( .A(n7848), .B(n7847), .X(n8412) );
  nor_x1_sg U57415 ( .A(n7847), .B(n7848), .X(n8413) );
  nand_x1_sg U57416 ( .A(n8666), .B(n8665), .X(n9230) );
  nor_x1_sg U57417 ( .A(n8665), .B(n8666), .X(n9231) );
  nand_x1_sg U57418 ( .A(n9486), .B(n9485), .X(n10050) );
  nor_x1_sg U57419 ( .A(n9485), .B(n9486), .X(n10051) );
  nand_x1_sg U57420 ( .A(n10305), .B(n10304), .X(n10869) );
  nor_x1_sg U57421 ( .A(n10304), .B(n10305), .X(n10870) );
  nand_x1_sg U57422 ( .A(n11124), .B(n11123), .X(n11688) );
  nor_x1_sg U57423 ( .A(n11123), .B(n11124), .X(n11689) );
  nand_x1_sg U57424 ( .A(n11943), .B(n11942), .X(n12507) );
  nor_x1_sg U57425 ( .A(n11942), .B(n11943), .X(n12508) );
  nand_x1_sg U57426 ( .A(n12762), .B(n12761), .X(n13326) );
  nor_x1_sg U57427 ( .A(n12761), .B(n12762), .X(n13327) );
  nand_x1_sg U57428 ( .A(n13581), .B(n13580), .X(n14145) );
  nor_x1_sg U57429 ( .A(n13580), .B(n13581), .X(n14146) );
  nand_x1_sg U57430 ( .A(n14400), .B(n14399), .X(n14964) );
  nor_x1_sg U57431 ( .A(n14399), .B(n14400), .X(n14965) );
  nand_x1_sg U57432 ( .A(n15219), .B(n15218), .X(n15783) );
  nor_x1_sg U57433 ( .A(n15218), .B(n15219), .X(n15784) );
  nand_x1_sg U57434 ( .A(n16038), .B(n16037), .X(n16602) );
  nor_x1_sg U57435 ( .A(n16037), .B(n16038), .X(n16603) );
  nand_x1_sg U57436 ( .A(n16857), .B(n16856), .X(n17419) );
  nor_x1_sg U57437 ( .A(n16856), .B(n16857), .X(n17420) );
  nand_x1_sg U57438 ( .A(n17676), .B(n17675), .X(n18240) );
  nor_x1_sg U57439 ( .A(n17675), .B(n17676), .X(n18241) );
  nand_x1_sg U57440 ( .A(n18497), .B(n18496), .X(n19061) );
  nor_x1_sg U57441 ( .A(n18496), .B(n18497), .X(n19062) );
  nand_x1_sg U57442 ( .A(n7275), .B(n46962), .X(n7268) );
  nand_x1_sg U57443 ( .A(n8094), .B(n47253), .X(n8087) );
  nand_x1_sg U57444 ( .A(n8912), .B(n47538), .X(n8905) );
  nand_x1_sg U57445 ( .A(n9732), .B(n47823), .X(n9725) );
  nand_x1_sg U57446 ( .A(n10551), .B(n48108), .X(n10544) );
  nand_x1_sg U57447 ( .A(n11370), .B(n48393), .X(n11363) );
  nand_x1_sg U57448 ( .A(n12189), .B(n48678), .X(n12182) );
  nand_x1_sg U57449 ( .A(n13008), .B(n48964), .X(n13001) );
  nand_x1_sg U57450 ( .A(n13827), .B(n49251), .X(n13820) );
  nand_x1_sg U57451 ( .A(n14646), .B(n49537), .X(n14639) );
  nand_x1_sg U57452 ( .A(n15465), .B(n49823), .X(n15458) );
  nand_x1_sg U57453 ( .A(n16284), .B(n50109), .X(n16277) );
  nand_x1_sg U57454 ( .A(n17100), .B(n50394), .X(n17093) );
  nand_x1_sg U57455 ( .A(n17922), .B(n50683), .X(n17915) );
  nand_x1_sg U57456 ( .A(n18743), .B(n50970), .X(n18736) );
  nand_x1_sg U57457 ( .A(n47045), .B(n7592), .X(n7591) );
  nand_x1_sg U57458 ( .A(n46940), .B(n7593), .X(n7590) );
  nand_x1_sg U57459 ( .A(n47332), .B(n8410), .X(n8409) );
  nand_x1_sg U57460 ( .A(n47231), .B(n8411), .X(n8408) );
  nand_x1_sg U57461 ( .A(n47617), .B(n9228), .X(n9227) );
  nand_x1_sg U57462 ( .A(n47516), .B(n9229), .X(n9226) );
  nand_x1_sg U57463 ( .A(n47902), .B(n10048), .X(n10047) );
  nand_x1_sg U57464 ( .A(n47801), .B(n10049), .X(n10046) );
  nand_x1_sg U57465 ( .A(n48187), .B(n10867), .X(n10866) );
  nand_x1_sg U57466 ( .A(n48086), .B(n10868), .X(n10865) );
  nand_x1_sg U57467 ( .A(n48472), .B(n11686), .X(n11685) );
  nand_x1_sg U57468 ( .A(n48371), .B(n11687), .X(n11684) );
  nand_x1_sg U57469 ( .A(n48757), .B(n12505), .X(n12504) );
  nand_x1_sg U57470 ( .A(n48656), .B(n12506), .X(n12503) );
  nand_x1_sg U57471 ( .A(n49043), .B(n13324), .X(n13323) );
  nand_x1_sg U57472 ( .A(n48942), .B(n13325), .X(n13322) );
  nand_x1_sg U57473 ( .A(n49330), .B(n14143), .X(n14142) );
  nand_x1_sg U57474 ( .A(n49229), .B(n14144), .X(n14141) );
  nand_x1_sg U57475 ( .A(n49616), .B(n14962), .X(n14961) );
  nand_x1_sg U57476 ( .A(n49515), .B(n14963), .X(n14960) );
  nand_x1_sg U57477 ( .A(n49902), .B(n15781), .X(n15780) );
  nand_x1_sg U57478 ( .A(n49801), .B(n15782), .X(n15779) );
  nand_x1_sg U57479 ( .A(n50188), .B(n16600), .X(n16599) );
  nand_x1_sg U57480 ( .A(n50087), .B(n16601), .X(n16598) );
  nand_x1_sg U57481 ( .A(n50762), .B(n18238), .X(n18237) );
  nand_x1_sg U57482 ( .A(n50661), .B(n18239), .X(n18236) );
  nand_x1_sg U57483 ( .A(n51049), .B(n19059), .X(n19058) );
  nand_x1_sg U57484 ( .A(n50948), .B(n19060), .X(n19057) );
  nand_x1_sg U57485 ( .A(n47060), .B(n47032), .X(n7607) );
  nand_x1_sg U57486 ( .A(n7608), .B(n7609), .X(n7606) );
  nand_x1_sg U57487 ( .A(n47346), .B(n47319), .X(n8425) );
  nand_x1_sg U57488 ( .A(n8426), .B(n8427), .X(n8424) );
  nand_x1_sg U57489 ( .A(n47631), .B(n47604), .X(n9243) );
  nand_x1_sg U57490 ( .A(n9244), .B(n9245), .X(n9242) );
  nand_x1_sg U57491 ( .A(n47916), .B(n47889), .X(n10063) );
  nand_x1_sg U57492 ( .A(n10064), .B(n10065), .X(n10062) );
  nand_x1_sg U57493 ( .A(n48201), .B(n48174), .X(n10882) );
  nand_x1_sg U57494 ( .A(n10883), .B(n10884), .X(n10881) );
  nand_x1_sg U57495 ( .A(n48486), .B(n48459), .X(n11701) );
  nand_x1_sg U57496 ( .A(n11702), .B(n11703), .X(n11700) );
  nand_x1_sg U57497 ( .A(n48771), .B(n48744), .X(n12520) );
  nand_x1_sg U57498 ( .A(n12521), .B(n12522), .X(n12519) );
  nand_x1_sg U57499 ( .A(n49058), .B(n49030), .X(n13339) );
  nand_x1_sg U57500 ( .A(n13340), .B(n13341), .X(n13338) );
  nand_x1_sg U57501 ( .A(n49344), .B(n49317), .X(n14158) );
  nand_x1_sg U57502 ( .A(n14159), .B(n14160), .X(n14157) );
  nand_x1_sg U57503 ( .A(n49630), .B(n49603), .X(n14977) );
  nand_x1_sg U57504 ( .A(n14978), .B(n14979), .X(n14976) );
  nand_x1_sg U57505 ( .A(n49916), .B(n49889), .X(n15796) );
  nand_x1_sg U57506 ( .A(n15797), .B(n15798), .X(n15795) );
  nand_x1_sg U57507 ( .A(n50202), .B(n50175), .X(n16615) );
  nand_x1_sg U57508 ( .A(n16616), .B(n16617), .X(n16614) );
  nand_x1_sg U57509 ( .A(n50487), .B(n50460), .X(n17432) );
  nand_x1_sg U57510 ( .A(n17433), .B(n17434), .X(n17431) );
  nand_x1_sg U57511 ( .A(n50776), .B(n50749), .X(n18253) );
  nand_x1_sg U57512 ( .A(n18254), .B(n18255), .X(n18252) );
  nand_x1_sg U57513 ( .A(n51063), .B(n51036), .X(n19074) );
  nand_x1_sg U57514 ( .A(n19075), .B(n19076), .X(n19073) );
  nand_x1_sg U57515 ( .A(n50473), .B(n17417), .X(n17416) );
  nand_x1_sg U57516 ( .A(n50372), .B(n17418), .X(n17415) );
  nand_x1_sg U57517 ( .A(n7381), .B(n39347), .X(n7488) );
  nand_x1_sg U57518 ( .A(n7464), .B(n46956), .X(n7462) );
  nor_x1_sg U57519 ( .A(n46956), .B(n7464), .X(n7463) );
  nand_x1_sg U57520 ( .A(n8199), .B(n39345), .X(n8306) );
  nand_x1_sg U57521 ( .A(n8282), .B(n47247), .X(n8280) );
  nor_x1_sg U57522 ( .A(n47247), .B(n8282), .X(n8281) );
  nand_x1_sg U57523 ( .A(n9017), .B(n39343), .X(n9124) );
  nand_x1_sg U57524 ( .A(n9100), .B(n47532), .X(n9098) );
  nor_x1_sg U57525 ( .A(n47532), .B(n9100), .X(n9099) );
  nand_x1_sg U57526 ( .A(n9837), .B(n39341), .X(n9944) );
  nand_x1_sg U57527 ( .A(n9920), .B(n47817), .X(n9918) );
  nor_x1_sg U57528 ( .A(n47817), .B(n9920), .X(n9919) );
  nand_x1_sg U57529 ( .A(n10656), .B(n39339), .X(n10763) );
  nand_x1_sg U57530 ( .A(n10739), .B(n48102), .X(n10737) );
  nor_x1_sg U57531 ( .A(n48102), .B(n10739), .X(n10738) );
  nand_x1_sg U57532 ( .A(n11475), .B(n39337), .X(n11582) );
  nand_x1_sg U57533 ( .A(n11558), .B(n48387), .X(n11556) );
  nor_x1_sg U57534 ( .A(n48387), .B(n11558), .X(n11557) );
  nand_x1_sg U57535 ( .A(n12294), .B(n39335), .X(n12401) );
  nand_x1_sg U57536 ( .A(n12377), .B(n48672), .X(n12375) );
  nor_x1_sg U57537 ( .A(n48672), .B(n12377), .X(n12376) );
  nand_x1_sg U57538 ( .A(n13113), .B(n39333), .X(n13220) );
  nand_x1_sg U57539 ( .A(n13196), .B(n48958), .X(n13194) );
  nor_x1_sg U57540 ( .A(n48958), .B(n13196), .X(n13195) );
  nand_x1_sg U57541 ( .A(n13932), .B(n39331), .X(n14039) );
  nand_x1_sg U57542 ( .A(n14015), .B(n49245), .X(n14013) );
  nor_x1_sg U57543 ( .A(n49245), .B(n14015), .X(n14014) );
  nand_x1_sg U57544 ( .A(n14751), .B(n39329), .X(n14858) );
  nand_x1_sg U57545 ( .A(n14834), .B(n49531), .X(n14832) );
  nor_x1_sg U57546 ( .A(n49531), .B(n14834), .X(n14833) );
  nand_x1_sg U57547 ( .A(n15570), .B(n39327), .X(n15677) );
  nand_x1_sg U57548 ( .A(n15653), .B(n49817), .X(n15651) );
  nor_x1_sg U57549 ( .A(n49817), .B(n15653), .X(n15652) );
  nand_x1_sg U57550 ( .A(n16389), .B(n39325), .X(n16496) );
  nand_x1_sg U57551 ( .A(n16472), .B(n50103), .X(n16470) );
  nor_x1_sg U57552 ( .A(n50103), .B(n16472), .X(n16471) );
  nand_x1_sg U57553 ( .A(n17289), .B(n50388), .X(n17287) );
  nor_x1_sg U57554 ( .A(n50388), .B(n17289), .X(n17288) );
  nand_x1_sg U57555 ( .A(n18027), .B(n39323), .X(n18134) );
  nand_x1_sg U57556 ( .A(n18110), .B(n50677), .X(n18108) );
  nor_x1_sg U57557 ( .A(n50677), .B(n18110), .X(n18109) );
  nand_x1_sg U57558 ( .A(n18848), .B(n39321), .X(n18955) );
  nand_x1_sg U57559 ( .A(n18931), .B(n50964), .X(n18929) );
  nor_x1_sg U57560 ( .A(n50964), .B(n18931), .X(n18930) );
  nand_x1_sg U57561 ( .A(n17130), .B(n17386), .X(n17385) );
  nor_x1_sg U57562 ( .A(n17386), .B(n17130), .X(n17387) );
  nand_x1_sg U57563 ( .A(n7371), .B(n7504), .X(n7503) );
  nor_x1_sg U57564 ( .A(n7504), .B(n7371), .X(n7505) );
  nand_x1_sg U57565 ( .A(n8189), .B(n8322), .X(n8321) );
  nor_x1_sg U57566 ( .A(n8322), .B(n8189), .X(n8323) );
  nand_x1_sg U57567 ( .A(n9007), .B(n9140), .X(n9139) );
  nor_x1_sg U57568 ( .A(n9140), .B(n9007), .X(n9141) );
  nand_x1_sg U57569 ( .A(n9827), .B(n9960), .X(n9959) );
  nor_x1_sg U57570 ( .A(n9960), .B(n9827), .X(n9961) );
  nand_x1_sg U57571 ( .A(n10646), .B(n10779), .X(n10778) );
  nor_x1_sg U57572 ( .A(n10779), .B(n10646), .X(n10780) );
  nand_x1_sg U57573 ( .A(n11465), .B(n11598), .X(n11597) );
  nor_x1_sg U57574 ( .A(n11598), .B(n11465), .X(n11599) );
  nand_x1_sg U57575 ( .A(n12284), .B(n12417), .X(n12416) );
  nor_x1_sg U57576 ( .A(n12417), .B(n12284), .X(n12418) );
  nand_x1_sg U57577 ( .A(n13103), .B(n13236), .X(n13235) );
  nor_x1_sg U57578 ( .A(n13236), .B(n13103), .X(n13237) );
  nand_x1_sg U57579 ( .A(n13922), .B(n14055), .X(n14054) );
  nor_x1_sg U57580 ( .A(n14055), .B(n13922), .X(n14056) );
  nand_x1_sg U57581 ( .A(n14741), .B(n14874), .X(n14873) );
  nor_x1_sg U57582 ( .A(n14874), .B(n14741), .X(n14875) );
  nand_x1_sg U57583 ( .A(n15560), .B(n15693), .X(n15692) );
  nor_x1_sg U57584 ( .A(n15693), .B(n15560), .X(n15694) );
  nand_x1_sg U57585 ( .A(n16379), .B(n16512), .X(n16511) );
  nor_x1_sg U57586 ( .A(n16512), .B(n16379), .X(n16513) );
  nand_x1_sg U57587 ( .A(n17196), .B(n17329), .X(n17328) );
  nor_x1_sg U57588 ( .A(n17329), .B(n17196), .X(n17330) );
  nand_x1_sg U57589 ( .A(n18017), .B(n18150), .X(n18149) );
  nor_x1_sg U57590 ( .A(n18150), .B(n18017), .X(n18151) );
  nand_x1_sg U57591 ( .A(n18838), .B(n18971), .X(n18970) );
  nor_x1_sg U57592 ( .A(n18971), .B(n18838), .X(n18972) );
  nand_x1_sg U57593 ( .A(n7302), .B(n7303), .X(n7301) );
  nor_x1_sg U57594 ( .A(n7303), .B(n7302), .X(n7304) );
  nand_x1_sg U57595 ( .A(n8120), .B(n8121), .X(n8119) );
  nor_x1_sg U57596 ( .A(n8121), .B(n8120), .X(n8122) );
  nand_x1_sg U57597 ( .A(n8938), .B(n8939), .X(n8937) );
  nor_x1_sg U57598 ( .A(n8939), .B(n8938), .X(n8940) );
  nand_x1_sg U57599 ( .A(n9758), .B(n9759), .X(n9757) );
  nor_x1_sg U57600 ( .A(n9759), .B(n9758), .X(n9760) );
  nand_x1_sg U57601 ( .A(n10577), .B(n10578), .X(n10576) );
  nor_x1_sg U57602 ( .A(n10578), .B(n10577), .X(n10579) );
  nand_x1_sg U57603 ( .A(n11396), .B(n11397), .X(n11395) );
  nor_x1_sg U57604 ( .A(n11397), .B(n11396), .X(n11398) );
  nand_x1_sg U57605 ( .A(n12215), .B(n12216), .X(n12214) );
  nor_x1_sg U57606 ( .A(n12216), .B(n12215), .X(n12217) );
  nand_x1_sg U57607 ( .A(n13034), .B(n13035), .X(n13033) );
  nor_x1_sg U57608 ( .A(n13035), .B(n13034), .X(n13036) );
  nand_x1_sg U57609 ( .A(n13853), .B(n13854), .X(n13852) );
  nor_x1_sg U57610 ( .A(n13854), .B(n13853), .X(n13855) );
  nand_x1_sg U57611 ( .A(n14672), .B(n14673), .X(n14671) );
  nor_x1_sg U57612 ( .A(n14673), .B(n14672), .X(n14674) );
  nand_x1_sg U57613 ( .A(n15491), .B(n15492), .X(n15490) );
  nor_x1_sg U57614 ( .A(n15492), .B(n15491), .X(n15493) );
  nand_x1_sg U57615 ( .A(n16310), .B(n16311), .X(n16309) );
  nor_x1_sg U57616 ( .A(n16311), .B(n16310), .X(n16312) );
  nand_x1_sg U57617 ( .A(n17948), .B(n17949), .X(n17947) );
  nor_x1_sg U57618 ( .A(n17949), .B(n17948), .X(n17950) );
  nand_x1_sg U57619 ( .A(n18769), .B(n18770), .X(n18768) );
  nor_x1_sg U57620 ( .A(n18770), .B(n18769), .X(n18771) );
  nand_x1_sg U57621 ( .A(n22972), .B(n41984), .X(n22980) );
  nand_x1_sg U57622 ( .A(n23249), .B(n41985), .X(n23257) );
  nand_x1_sg U57623 ( .A(n23529), .B(n41979), .X(n23537) );
  nand_x1_sg U57624 ( .A(n23808), .B(n41980), .X(n23816) );
  nand_x1_sg U57625 ( .A(n24087), .B(n41981), .X(n24095) );
  nand_x1_sg U57626 ( .A(n24366), .B(n41982), .X(n24374) );
  nand_x1_sg U57627 ( .A(n24645), .B(n41975), .X(n24653) );
  nand_x1_sg U57628 ( .A(n24923), .B(n41976), .X(n24931) );
  nand_x1_sg U57629 ( .A(n25202), .B(n41977), .X(n25210) );
  nand_x1_sg U57630 ( .A(n25481), .B(n41978), .X(n25489) );
  nand_x1_sg U57631 ( .A(n25760), .B(n41972), .X(n25768) );
  nand_x1_sg U57632 ( .A(n26317), .B(n41973), .X(n26324) );
  nand_x1_sg U57633 ( .A(n26597), .B(n41974), .X(n26605) );
  nor_x1_sg U57634 ( .A(n22943), .B(n22944), .X(n22942) );
  nor_x1_sg U57635 ( .A(n22946), .B(n41469), .X(n22941) );
  nor_x1_sg U57636 ( .A(n41712), .B(n22945), .X(n22944) );
  nor_x1_sg U57637 ( .A(n23192), .B(n23193), .X(n23191) );
  nor_x1_sg U57638 ( .A(n23195), .B(n39152), .X(n23190) );
  nor_x1_sg U57639 ( .A(n41735), .B(n23194), .X(n23193) );
  nor_x1_sg U57640 ( .A(n23234), .B(n23235), .X(n23233) );
  nor_x1_sg U57641 ( .A(n23237), .B(n41466), .X(n23232) );
  nor_x1_sg U57642 ( .A(n39036), .B(n23236), .X(n23235) );
  nor_x1_sg U57643 ( .A(n23486), .B(n23487), .X(n23485) );
  nor_x1_sg U57644 ( .A(n23489), .B(n39654), .X(n23484) );
  nor_x1_sg U57645 ( .A(n39857), .B(n23488), .X(n23487) );
  nor_x1_sg U57646 ( .A(n23779), .B(n23780), .X(n23778) );
  nor_x1_sg U57647 ( .A(n23782), .B(n40019), .X(n23777) );
  nor_x1_sg U57648 ( .A(n41713), .B(n23781), .X(n23780) );
  nor_x1_sg U57649 ( .A(n24030), .B(n24031), .X(n24029) );
  nor_x1_sg U57650 ( .A(n24033), .B(n41410), .X(n24028) );
  nor_x1_sg U57651 ( .A(n41726), .B(n24032), .X(n24031) );
  nor_x1_sg U57652 ( .A(n24072), .B(n24073), .X(n24071) );
  nor_x1_sg U57653 ( .A(n24075), .B(n41467), .X(n24070) );
  nor_x1_sg U57654 ( .A(n41627), .B(n24074), .X(n24073) );
  nor_x1_sg U57655 ( .A(n24323), .B(n24324), .X(n24322) );
  nor_x1_sg U57656 ( .A(n24326), .B(n40021), .X(n24321) );
  nor_x1_sg U57657 ( .A(n39869), .B(n24325), .X(n24324) );
  nor_x1_sg U57658 ( .A(n24616), .B(n24617), .X(n24615) );
  nor_x1_sg U57659 ( .A(n24619), .B(n40371), .X(n24614) );
  nor_x1_sg U57660 ( .A(n41718), .B(n24618), .X(n24617) );
  nor_x1_sg U57661 ( .A(n24866), .B(n24867), .X(n24865) );
  nor_x1_sg U57662 ( .A(n24869), .B(n40371), .X(n24864) );
  nor_x1_sg U57663 ( .A(n41728), .B(n24868), .X(n24867) );
  nor_x1_sg U57664 ( .A(n24908), .B(n24909), .X(n24907) );
  nor_x1_sg U57665 ( .A(n24911), .B(n40456), .X(n24906) );
  nor_x1_sg U57666 ( .A(n39030), .B(n24910), .X(n24909) );
  nor_x1_sg U57667 ( .A(n25159), .B(n25160), .X(n25158) );
  nor_x1_sg U57668 ( .A(n25162), .B(n40370), .X(n25157) );
  nor_x1_sg U57669 ( .A(n39878), .B(n25161), .X(n25160) );
  nor_x1_sg U57670 ( .A(n25452), .B(n25453), .X(n25451) );
  nor_x1_sg U57671 ( .A(n25455), .B(n40020), .X(n25450) );
  nor_x1_sg U57672 ( .A(n41719), .B(n25454), .X(n25453) );
  nor_x1_sg U57673 ( .A(n25703), .B(n25704), .X(n25702) );
  nor_x1_sg U57674 ( .A(n25706), .B(n41310), .X(n25701) );
  nor_x1_sg U57675 ( .A(n41732), .B(n25705), .X(n25704) );
  nor_x1_sg U57676 ( .A(n25745), .B(n25746), .X(n25744) );
  nor_x1_sg U57677 ( .A(n25748), .B(n41404), .X(n25743) );
  nor_x1_sg U57678 ( .A(n41622), .B(n25747), .X(n25746) );
  nor_x1_sg U57679 ( .A(n26540), .B(n26541), .X(n26539) );
  nor_x1_sg U57680 ( .A(n26543), .B(n39152), .X(n26538) );
  nor_x1_sg U57681 ( .A(n41737), .B(n26542), .X(n26541) );
  nor_x1_sg U57682 ( .A(n26582), .B(n26583), .X(n26581) );
  nor_x1_sg U57683 ( .A(n26585), .B(n41407), .X(n26580) );
  nor_x1_sg U57684 ( .A(n39026), .B(n26584), .X(n26583) );
  nor_x1_sg U57685 ( .A(n22915), .B(n22916), .X(n22914) );
  nor_x1_sg U57686 ( .A(n22918), .B(n40015), .X(n22913) );
  nor_x1_sg U57687 ( .A(n41736), .B(n22917), .X(n22916) );
  nor_x1_sg U57688 ( .A(n22929), .B(n22930), .X(n22928) );
  nor_x1_sg U57689 ( .A(n22932), .B(n40018), .X(n22927) );
  nor_x1_sg U57690 ( .A(n41664), .B(n22931), .X(n22930) );
  nor_x1_sg U57691 ( .A(n22957), .B(n22958), .X(n22956) );
  nor_x1_sg U57692 ( .A(n22960), .B(n39436), .X(n22955) );
  nor_x1_sg U57693 ( .A(n41629), .B(n22959), .X(n22958) );
  nor_x1_sg U57694 ( .A(n23206), .B(n23207), .X(n23205) );
  nor_x1_sg U57695 ( .A(n23209), .B(n39274), .X(n23204) );
  nor_x1_sg U57696 ( .A(n39861), .B(n23208), .X(n23207) );
  nor_x1_sg U57697 ( .A(n23220), .B(n23221), .X(n23219) );
  nor_x1_sg U57698 ( .A(n23223), .B(n41469), .X(n23218) );
  nor_x1_sg U57699 ( .A(n41711), .B(n23222), .X(n23221) );
  nor_x1_sg U57700 ( .A(n23472), .B(n23473), .X(n23471) );
  nor_x1_sg U57701 ( .A(n23475), .B(n40373), .X(n23470) );
  nor_x1_sg U57702 ( .A(n41734), .B(n23474), .X(n23473) );
  nor_x1_sg U57703 ( .A(n23500), .B(n23501), .X(n23499) );
  nor_x1_sg U57704 ( .A(n23503), .B(n39436), .X(n23498) );
  nor_x1_sg U57705 ( .A(n41714), .B(n23502), .X(n23501) );
  nor_x1_sg U57706 ( .A(n23514), .B(n23515), .X(n23513) );
  nor_x1_sg U57707 ( .A(n23517), .B(n41404), .X(n23512) );
  nor_x1_sg U57708 ( .A(n39034), .B(n23516), .X(n23515) );
  nor_x1_sg U57709 ( .A(n23751), .B(n23752), .X(n23750) );
  nor_x1_sg U57710 ( .A(n23754), .B(n41399), .X(n23749) );
  nor_x1_sg U57711 ( .A(n41727), .B(n23753), .X(n23752) );
  nor_x1_sg U57712 ( .A(n23765), .B(n23766), .X(n23764) );
  nor_x1_sg U57713 ( .A(n23768), .B(n38813), .X(n23763) );
  nor_x1_sg U57714 ( .A(n39863), .B(n23767), .X(n23766) );
  nor_x1_sg U57715 ( .A(n23793), .B(n23794), .X(n23792) );
  nor_x1_sg U57716 ( .A(n23796), .B(n40454), .X(n23791) );
  nor_x1_sg U57717 ( .A(n39032), .B(n23795), .X(n23794) );
  nor_x1_sg U57718 ( .A(n24044), .B(n24045), .X(n24043) );
  nor_x1_sg U57719 ( .A(n24047), .B(n40370), .X(n24042) );
  nor_x1_sg U57720 ( .A(n39866), .B(n24046), .X(n24045) );
  nor_x1_sg U57721 ( .A(n24058), .B(n24059), .X(n24057) );
  nor_x1_sg U57722 ( .A(n24061), .B(n39284), .X(n24056) );
  nor_x1_sg U57723 ( .A(n41716), .B(n24060), .X(n24059) );
  nor_x1_sg U57724 ( .A(n24309), .B(n24310), .X(n24308) );
  nor_x1_sg U57725 ( .A(n24312), .B(n40014), .X(n24307) );
  nor_x1_sg U57726 ( .A(n41730), .B(n24311), .X(n24310) );
  nor_x1_sg U57727 ( .A(n24337), .B(n24338), .X(n24336) );
  nor_x1_sg U57728 ( .A(n24340), .B(n39155), .X(n24335) );
  nor_x1_sg U57729 ( .A(n41715), .B(n24339), .X(n24338) );
  nor_x1_sg U57730 ( .A(n24351), .B(n24352), .X(n24350) );
  nor_x1_sg U57731 ( .A(n24354), .B(n39154), .X(n24349) );
  nor_x1_sg U57732 ( .A(n41625), .B(n24353), .X(n24352) );
  nor_x1_sg U57733 ( .A(n24588), .B(n24589), .X(n24587) );
  nor_x1_sg U57734 ( .A(n24591), .B(n40021), .X(n24586) );
  nor_x1_sg U57735 ( .A(n41729), .B(n24590), .X(n24589) );
  nor_x1_sg U57736 ( .A(n24602), .B(n24603), .X(n24601) );
  nor_x1_sg U57737 ( .A(n24605), .B(n40454), .X(n24600) );
  nor_x1_sg U57738 ( .A(n39872), .B(n24604), .X(n24603) );
  nor_x1_sg U57739 ( .A(n24630), .B(n24631), .X(n24629) );
  nor_x1_sg U57740 ( .A(n24633), .B(n39284), .X(n24628) );
  nor_x1_sg U57741 ( .A(n49055), .B(n24632), .X(n24631) );
  nor_x1_sg U57742 ( .A(n24880), .B(n24881), .X(n24879) );
  nor_x1_sg U57743 ( .A(n24883), .B(n41408), .X(n24878) );
  nor_x1_sg U57744 ( .A(n39875), .B(n24882), .X(n24881) );
  nor_x1_sg U57745 ( .A(n24894), .B(n24895), .X(n24893) );
  nor_x1_sg U57746 ( .A(n24897), .B(n40015), .X(n24892) );
  nor_x1_sg U57747 ( .A(n41717), .B(n24896), .X(n24895) );
  nor_x1_sg U57748 ( .A(n25145), .B(n25146), .X(n25144) );
  nor_x1_sg U57749 ( .A(n25148), .B(n41410), .X(n25143) );
  nor_x1_sg U57750 ( .A(n41731), .B(n25147), .X(n25146) );
  nor_x1_sg U57751 ( .A(n25173), .B(n25174), .X(n25172) );
  nor_x1_sg U57752 ( .A(n25176), .B(n40374), .X(n25171) );
  nor_x1_sg U57753 ( .A(n41720), .B(n25175), .X(n25174) );
  nor_x1_sg U57754 ( .A(n25187), .B(n25188), .X(n25186) );
  nor_x1_sg U57755 ( .A(n25190), .B(n38981), .X(n25185) );
  nor_x1_sg U57756 ( .A(n41623), .B(n25189), .X(n25188) );
  nor_x1_sg U57757 ( .A(n25424), .B(n25425), .X(n25423) );
  nor_x1_sg U57758 ( .A(n25427), .B(n40376), .X(n25422) );
  nor_x1_sg U57759 ( .A(n41733), .B(n25426), .X(n25425) );
  nor_x1_sg U57760 ( .A(n25438), .B(n25439), .X(n25437) );
  nor_x1_sg U57761 ( .A(n25441), .B(n40020), .X(n25436) );
  nor_x1_sg U57762 ( .A(n39896), .B(n25440), .X(n25439) );
  nor_x1_sg U57763 ( .A(n25466), .B(n25467), .X(n25465) );
  nor_x1_sg U57764 ( .A(n25469), .B(n41404), .X(n25464) );
  nor_x1_sg U57765 ( .A(n39027), .B(n25468), .X(n25467) );
  nor_x1_sg U57766 ( .A(n25717), .B(n25718), .X(n25716) );
  nor_x1_sg U57767 ( .A(n25720), .B(n39275), .X(n25715) );
  nor_x1_sg U57768 ( .A(n39881), .B(n25719), .X(n25718) );
  nor_x1_sg U57769 ( .A(n25731), .B(n25732), .X(n25730) );
  nor_x1_sg U57770 ( .A(n25734), .B(n40016), .X(n25729) );
  nor_x1_sg U57771 ( .A(n41722), .B(n25733), .X(n25732) );
  nor_x1_sg U57772 ( .A(n26554), .B(n26555), .X(n26553) );
  nor_x1_sg U57773 ( .A(n26557), .B(n39653), .X(n26552) );
  nor_x1_sg U57774 ( .A(n39890), .B(n26556), .X(n26555) );
  nor_x1_sg U57775 ( .A(n26568), .B(n26569), .X(n26567) );
  nor_x1_sg U57776 ( .A(n26571), .B(n39151), .X(n26566) );
  nor_x1_sg U57777 ( .A(n41723), .B(n26570), .X(n26569) );
  inv_x1_sg U57778 ( .A(n16927), .X(n50288) );
  nand_x1_sg U57779 ( .A(n39222), .B(n47358), .X(n22965) );
  nand_x1_sg U57780 ( .A(n39224), .B(n47643), .X(n23242) );
  nand_x1_sg U57781 ( .A(n41184), .B(n47928), .X(n23522) );
  nand_x1_sg U57782 ( .A(n41177), .B(n48213), .X(n23801) );
  nand_x1_sg U57783 ( .A(n41173), .B(n48498), .X(n24080) );
  nand_x1_sg U57784 ( .A(n41170), .B(n48783), .X(n24359) );
  nand_x1_sg U57785 ( .A(n41164), .B(n49070), .X(n24638) );
  nand_x1_sg U57786 ( .A(n41160), .B(n49356), .X(n24916) );
  nand_x1_sg U57787 ( .A(n41153), .B(n49642), .X(n25195) );
  nand_x1_sg U57788 ( .A(n41147), .B(n49928), .X(n25474) );
  nand_x1_sg U57789 ( .A(n41145), .B(n50214), .X(n25753) );
  nand_x1_sg U57790 ( .A(n39244), .B(n50788), .X(n26309) );
  nand_x1_sg U57791 ( .A(n41133), .B(n51075), .X(n26590) );
  nand_x1_sg U57792 ( .A(n6949), .B(n6950), .X(n6948) );
  nand_x1_sg U57793 ( .A(n7766), .B(n7767), .X(n7765) );
  nand_x1_sg U57794 ( .A(n8584), .B(n8585), .X(n8583) );
  nand_x1_sg U57795 ( .A(n9404), .B(n9405), .X(n9403) );
  nand_x1_sg U57796 ( .A(n10223), .B(n10224), .X(n10222) );
  nand_x1_sg U57797 ( .A(n11042), .B(n11043), .X(n11041) );
  nand_x1_sg U57798 ( .A(n11861), .B(n11862), .X(n11860) );
  nand_x1_sg U57799 ( .A(n12680), .B(n12681), .X(n12679) );
  nand_x1_sg U57800 ( .A(n13499), .B(n13500), .X(n13498) );
  nand_x1_sg U57801 ( .A(n14318), .B(n14319), .X(n14317) );
  nand_x1_sg U57802 ( .A(n15137), .B(n15138), .X(n15136) );
  nand_x1_sg U57803 ( .A(n15956), .B(n15957), .X(n15955) );
  nand_x1_sg U57804 ( .A(n16773), .B(n16774), .X(n16772) );
  nand_x1_sg U57805 ( .A(n17594), .B(n17595), .X(n17593) );
  nand_x1_sg U57806 ( .A(n18415), .B(n18416), .X(n18414) );
  nand_x1_sg U57807 ( .A(n46875), .B(n7135), .X(n7121) );
  nand_x1_sg U57808 ( .A(n47168), .B(n7953), .X(n7939) );
  nand_x1_sg U57809 ( .A(n47453), .B(n8771), .X(n8757) );
  nand_x1_sg U57810 ( .A(n47738), .B(n9591), .X(n9577) );
  nand_x1_sg U57811 ( .A(n48023), .B(n10410), .X(n10396) );
  nand_x1_sg U57812 ( .A(n48308), .B(n11229), .X(n11215) );
  nand_x1_sg U57813 ( .A(n48593), .B(n12048), .X(n12034) );
  nand_x1_sg U57814 ( .A(n48879), .B(n12867), .X(n12853) );
  nand_x1_sg U57815 ( .A(n49166), .B(n13686), .X(n13672) );
  nand_x1_sg U57816 ( .A(n49452), .B(n14505), .X(n14491) );
  nand_x1_sg U57817 ( .A(n49737), .B(n15324), .X(n15310) );
  nand_x1_sg U57818 ( .A(n50024), .B(n16143), .X(n16129) );
  nand_x1_sg U57819 ( .A(n50309), .B(n16960), .X(n16946) );
  nand_x1_sg U57820 ( .A(n50598), .B(n17781), .X(n17767) );
  nand_x1_sg U57821 ( .A(n50885), .B(n18602), .X(n18588) );
  inv_x1_sg U57822 ( .A(n8410), .X(n47231) );
  inv_x1_sg U57823 ( .A(n9228), .X(n47516) );
  inv_x1_sg U57824 ( .A(n10048), .X(n47801) );
  inv_x1_sg U57825 ( .A(n10867), .X(n48086) );
  inv_x1_sg U57826 ( .A(n11686), .X(n48371) );
  inv_x1_sg U57827 ( .A(n12505), .X(n48656) );
  inv_x1_sg U57828 ( .A(n13324), .X(n48942) );
  inv_x1_sg U57829 ( .A(n14143), .X(n49229) );
  inv_x1_sg U57830 ( .A(n14962), .X(n49515) );
  inv_x1_sg U57831 ( .A(n15781), .X(n49801) );
  inv_x1_sg U57832 ( .A(n16600), .X(n50087) );
  inv_x1_sg U57833 ( .A(n17417), .X(n50372) );
  inv_x1_sg U57834 ( .A(n18238), .X(n50661) );
  inv_x1_sg U57835 ( .A(n19059), .X(n50948) );
  inv_x1_sg U57836 ( .A(n26010), .X(n50499) );
  inv_x1_sg U57837 ( .A(n7592), .X(n46940) );
  nand_x1_sg U57838 ( .A(n41305), .B(n47072), .X(n22691) );
  inv_x1_sg U57839 ( .A(n8369), .X(n47213) );
  inv_x1_sg U57840 ( .A(n9187), .X(n47498) );
  inv_x1_sg U57841 ( .A(n10007), .X(n47783) );
  inv_x1_sg U57842 ( .A(n10826), .X(n48068) );
  inv_x1_sg U57843 ( .A(n11645), .X(n48353) );
  inv_x1_sg U57844 ( .A(n12464), .X(n48638) );
  inv_x1_sg U57845 ( .A(n13283), .X(n48924) );
  inv_x1_sg U57846 ( .A(n14102), .X(n49211) );
  inv_x1_sg U57847 ( .A(n14921), .X(n49497) );
  inv_x1_sg U57848 ( .A(n15740), .X(n49783) );
  inv_x1_sg U57849 ( .A(n16559), .X(n50069) );
  inv_x1_sg U57850 ( .A(n18197), .X(n50643) );
  inv_x1_sg U57851 ( .A(n19018), .X(n50930) );
  nor_x1_sg U57852 ( .A(n7178), .B(n7179), .X(n7177) );
  nor_x1_sg U57853 ( .A(n7997), .B(n7998), .X(n7996) );
  nor_x1_sg U57854 ( .A(n8815), .B(n8816), .X(n8814) );
  nor_x1_sg U57855 ( .A(n9635), .B(n9636), .X(n9634) );
  nor_x1_sg U57856 ( .A(n10454), .B(n10455), .X(n10453) );
  nor_x1_sg U57857 ( .A(n11273), .B(n11274), .X(n11272) );
  nor_x1_sg U57858 ( .A(n12092), .B(n12093), .X(n12091) );
  nor_x1_sg U57859 ( .A(n12911), .B(n12912), .X(n12910) );
  nor_x1_sg U57860 ( .A(n13730), .B(n13731), .X(n13729) );
  nor_x1_sg U57861 ( .A(n14549), .B(n14550), .X(n14548) );
  nor_x1_sg U57862 ( .A(n15368), .B(n15369), .X(n15367) );
  nor_x1_sg U57863 ( .A(n16187), .B(n16188), .X(n16186) );
  nor_x1_sg U57864 ( .A(n17003), .B(n17004), .X(n17002) );
  nor_x1_sg U57865 ( .A(n17825), .B(n17826), .X(n17824) );
  nor_x1_sg U57866 ( .A(n18646), .B(n18647), .X(n18645) );
  nor_x1_sg U57867 ( .A(n22660), .B(n22661), .X(n22659) );
  nor_x1_sg U57868 ( .A(n22663), .B(n39155), .X(n22658) );
  nor_x1_sg U57869 ( .A(n39854), .B(n22662), .X(n22661) );
  nor_x1_sg U57870 ( .A(n22678), .B(n22679), .X(n22677) );
  nor_x1_sg U57871 ( .A(n22681), .B(n40375), .X(n22676) );
  nor_x1_sg U57872 ( .A(n41666), .B(n22680), .X(n22679) );
  nor_x1_sg U57873 ( .A(n25984), .B(n25985), .X(n25983) );
  nor_x1_sg U57874 ( .A(n25987), .B(n40016), .X(n25982) );
  nor_x1_sg U57875 ( .A(n39885), .B(n25986), .X(n25985) );
  nor_x1_sg U57876 ( .A(n26284), .B(n26285), .X(n26283) );
  nor_x1_sg U57877 ( .A(n26287), .B(n40019), .X(n26282) );
  nor_x1_sg U57878 ( .A(n41721), .B(n26286), .X(n26285) );
  nor_x1_sg U57879 ( .A(n46938), .B(n22648), .X(n22647) );
  nor_x1_sg U57880 ( .A(n22650), .B(n41466), .X(n22646) );
  nor_x1_sg U57881 ( .A(n39725), .B(n22649), .X(n22648) );
  nor_x1_sg U57882 ( .A(n22666), .B(n22667), .X(n22665) );
  nor_x1_sg U57883 ( .A(n22669), .B(n39284), .X(n22664) );
  nor_x1_sg U57884 ( .A(n39605), .B(n22668), .X(n22667) );
  nor_x1_sg U57885 ( .A(n22672), .B(n22673), .X(n22671) );
  nor_x1_sg U57886 ( .A(n22675), .B(n39283), .X(n22670) );
  nor_x1_sg U57887 ( .A(n41710), .B(n22674), .X(n22673) );
  nor_x1_sg U57888 ( .A(n22684), .B(n22685), .X(n22683) );
  nor_x1_sg U57889 ( .A(n22687), .B(n39283), .X(n22682) );
  nor_x1_sg U57890 ( .A(n41631), .B(n22686), .X(n22685) );
  nor_x1_sg U57891 ( .A(n25933), .B(n25934), .X(n25932) );
  nor_x1_sg U57892 ( .A(n25936), .B(n41402), .X(n25931) );
  nor_x1_sg U57893 ( .A(n39679), .B(n25935), .X(n25934) );
  nor_x1_sg U57894 ( .A(n25971), .B(n25972), .X(n25970) );
  nor_x1_sg U57895 ( .A(n25974), .B(n41469), .X(n25969) );
  nor_x1_sg U57896 ( .A(n41739), .B(n25973), .X(n25972) );
  nor_x1_sg U57897 ( .A(n25997), .B(n25998), .X(n25996) );
  nor_x1_sg U57898 ( .A(n26000), .B(n39282), .X(n25995) );
  nor_x1_sg U57899 ( .A(n41724), .B(n25999), .X(n25998) );
  nor_x1_sg U57900 ( .A(n26010), .B(n26011), .X(n26009) );
  nor_x1_sg U57901 ( .A(n26013), .B(n40018), .X(n26008) );
  nor_x1_sg U57902 ( .A(n41618), .B(n26012), .X(n26011) );
  nor_x1_sg U57903 ( .A(n26252), .B(n26253), .X(n26251) );
  nor_x1_sg U57904 ( .A(n26255), .B(n41407), .X(n26250) );
  nor_x1_sg U57905 ( .A(n41738), .B(n26254), .X(n26253) );
  nor_x1_sg U57906 ( .A(n26268), .B(n26269), .X(n26267) );
  nor_x1_sg U57907 ( .A(n26271), .B(n39653), .X(n26266) );
  nor_x1_sg U57908 ( .A(n39888), .B(n26270), .X(n26269) );
  nor_x1_sg U57909 ( .A(n26300), .B(n26301), .X(n26299) );
  nor_x1_sg U57910 ( .A(n26303), .B(n41399), .X(n26298) );
  nor_x1_sg U57911 ( .A(n41619), .B(n26302), .X(n26301) );
  nand_x1_sg U57912 ( .A(n38941), .B(n50499), .X(n26017) );
  nand_x1_sg U57913 ( .A(n16899), .B(n16895), .X(n16897) );
  nor_x1_sg U57914 ( .A(n16895), .B(n16899), .X(n16898) );
  nand_x1_sg U57915 ( .A(n7072), .B(n7068), .X(n7070) );
  nor_x1_sg U57916 ( .A(n7068), .B(n7072), .X(n7071) );
  nand_x1_sg U57917 ( .A(n7890), .B(n7886), .X(n7888) );
  nor_x1_sg U57918 ( .A(n7886), .B(n7890), .X(n7889) );
  nand_x1_sg U57919 ( .A(n8708), .B(n8704), .X(n8706) );
  nor_x1_sg U57920 ( .A(n8704), .B(n8708), .X(n8707) );
  nand_x1_sg U57921 ( .A(n9528), .B(n9524), .X(n9526) );
  nor_x1_sg U57922 ( .A(n9524), .B(n9528), .X(n9527) );
  nand_x1_sg U57923 ( .A(n10347), .B(n10343), .X(n10345) );
  nor_x1_sg U57924 ( .A(n10343), .B(n10347), .X(n10346) );
  nand_x1_sg U57925 ( .A(n11166), .B(n11162), .X(n11164) );
  nor_x1_sg U57926 ( .A(n11162), .B(n11166), .X(n11165) );
  nand_x1_sg U57927 ( .A(n11985), .B(n11981), .X(n11983) );
  nor_x1_sg U57928 ( .A(n11981), .B(n11985), .X(n11984) );
  nand_x1_sg U57929 ( .A(n12804), .B(n12800), .X(n12802) );
  nor_x1_sg U57930 ( .A(n12800), .B(n12804), .X(n12803) );
  nand_x1_sg U57931 ( .A(n13623), .B(n13619), .X(n13621) );
  nor_x1_sg U57932 ( .A(n13619), .B(n13623), .X(n13622) );
  nand_x1_sg U57933 ( .A(n14442), .B(n14438), .X(n14440) );
  nor_x1_sg U57934 ( .A(n14438), .B(n14442), .X(n14441) );
  nand_x1_sg U57935 ( .A(n15261), .B(n15257), .X(n15259) );
  nor_x1_sg U57936 ( .A(n15257), .B(n15261), .X(n15260) );
  nand_x1_sg U57937 ( .A(n16080), .B(n16076), .X(n16078) );
  nor_x1_sg U57938 ( .A(n16076), .B(n16080), .X(n16079) );
  nand_x1_sg U57939 ( .A(n17718), .B(n17714), .X(n17716) );
  nor_x1_sg U57940 ( .A(n17714), .B(n17718), .X(n17717) );
  nand_x1_sg U57941 ( .A(n18539), .B(n18535), .X(n18537) );
  nor_x1_sg U57942 ( .A(n18535), .B(n18539), .X(n18538) );
  nand_x1_sg U57943 ( .A(n46996), .B(n7312), .X(n7318) );
  inv_x1_sg U57944 ( .A(n7311), .X(n46996) );
  nand_x1_sg U57945 ( .A(n50426), .B(n17137), .X(n17143) );
  inv_x1_sg U57946 ( .A(n17136), .X(n50426) );
  nand_x1_sg U57947 ( .A(n8343), .B(n8296), .X(n8341) );
  nand_x1_sg U57948 ( .A(n9161), .B(n9114), .X(n9159) );
  nand_x1_sg U57949 ( .A(n9981), .B(n9934), .X(n9979) );
  nand_x1_sg U57950 ( .A(n10800), .B(n10753), .X(n10798) );
  nand_x1_sg U57951 ( .A(n11619), .B(n11572), .X(n11617) );
  nand_x1_sg U57952 ( .A(n12438), .B(n12391), .X(n12436) );
  nand_x1_sg U57953 ( .A(n13257), .B(n13210), .X(n13255) );
  nand_x1_sg U57954 ( .A(n14076), .B(n14029), .X(n14074) );
  nand_x1_sg U57955 ( .A(n14895), .B(n14848), .X(n14893) );
  nand_x1_sg U57956 ( .A(n15714), .B(n15667), .X(n15712) );
  nand_x1_sg U57957 ( .A(n16533), .B(n16486), .X(n16531) );
  nand_x1_sg U57958 ( .A(n18171), .B(n18124), .X(n18169) );
  nand_x1_sg U57959 ( .A(n18992), .B(n18945), .X(n18990) );
  nand_x1_sg U57960 ( .A(n7525), .B(n7478), .X(n7523) );
  nand_x1_sg U57961 ( .A(n17350), .B(n17303), .X(n17348) );
  nand_x1_sg U57962 ( .A(n17315), .B(n17316), .X(n17314) );
  nor_x1_sg U57963 ( .A(n17316), .B(n17315), .X(n17317) );
  inv_x1_sg U57964 ( .A(n22957), .X(n47358) );
  inv_x1_sg U57965 ( .A(n23234), .X(n47643) );
  inv_x1_sg U57966 ( .A(n23514), .X(n47928) );
  inv_x1_sg U57967 ( .A(n23793), .X(n48213) );
  inv_x1_sg U57968 ( .A(n24072), .X(n48498) );
  inv_x1_sg U57969 ( .A(n24351), .X(n48783) );
  inv_x1_sg U57970 ( .A(n24630), .X(n49070) );
  inv_x1_sg U57971 ( .A(n24908), .X(n49356) );
  inv_x1_sg U57972 ( .A(n25187), .X(n49642) );
  inv_x1_sg U57973 ( .A(n25466), .X(n49928) );
  inv_x1_sg U57974 ( .A(n25745), .X(n50214) );
  inv_x1_sg U57975 ( .A(n26300), .X(n50788) );
  inv_x1_sg U57976 ( .A(n26582), .X(n51075) );
  inv_x1_sg U57977 ( .A(n7166), .X(n46901) );
  inv_x1_sg U57978 ( .A(n16991), .X(n50334) );
  inv_x1_sg U57979 ( .A(n22653), .X(n46963) );
  inv_x1_sg U57980 ( .A(n7985), .X(n47186) );
  inv_x1_sg U57981 ( .A(n8803), .X(n47471) );
  inv_x1_sg U57982 ( .A(n9623), .X(n47756) );
  inv_x1_sg U57983 ( .A(n10442), .X(n48041) );
  inv_x1_sg U57984 ( .A(n11261), .X(n48326) );
  inv_x1_sg U57985 ( .A(n12080), .X(n48611) );
  inv_x1_sg U57986 ( .A(n12899), .X(n48897) );
  inv_x1_sg U57987 ( .A(n13718), .X(n49184) );
  inv_x1_sg U57988 ( .A(n14537), .X(n49470) );
  inv_x1_sg U57989 ( .A(n15356), .X(n49756) );
  inv_x1_sg U57990 ( .A(n16175), .X(n50042) );
  inv_x1_sg U57991 ( .A(n17813), .X(n50616) );
  inv_x1_sg U57992 ( .A(n18634), .X(n50903) );
  inv_x1_sg U57993 ( .A(n7276), .X(n46962) );
  inv_x1_sg U57994 ( .A(n8095), .X(n47253) );
  inv_x1_sg U57995 ( .A(n8913), .X(n47538) );
  inv_x1_sg U57996 ( .A(n9733), .X(n47823) );
  inv_x1_sg U57997 ( .A(n10552), .X(n48108) );
  inv_x1_sg U57998 ( .A(n11371), .X(n48393) );
  inv_x1_sg U57999 ( .A(n12190), .X(n48678) );
  inv_x1_sg U58000 ( .A(n13009), .X(n48964) );
  inv_x1_sg U58001 ( .A(n13828), .X(n49251) );
  inv_x1_sg U58002 ( .A(n14647), .X(n49537) );
  inv_x1_sg U58003 ( .A(n15466), .X(n49823) );
  inv_x1_sg U58004 ( .A(n16285), .X(n50109) );
  inv_x1_sg U58005 ( .A(n17923), .X(n50683) );
  inv_x1_sg U58006 ( .A(n18744), .X(n50970) );
  inv_x1_sg U58007 ( .A(n7082), .X(n46871) );
  inv_x1_sg U58008 ( .A(n7900), .X(n47164) );
  inv_x1_sg U58009 ( .A(n8718), .X(n47449) );
  inv_x1_sg U58010 ( .A(n9538), .X(n47734) );
  inv_x1_sg U58011 ( .A(n10357), .X(n48019) );
  inv_x1_sg U58012 ( .A(n11176), .X(n48304) );
  inv_x1_sg U58013 ( .A(n11995), .X(n48589) );
  inv_x1_sg U58014 ( .A(n12814), .X(n48875) );
  inv_x1_sg U58015 ( .A(n13633), .X(n49162) );
  inv_x1_sg U58016 ( .A(n14452), .X(n49448) );
  inv_x1_sg U58017 ( .A(n15271), .X(n49733) );
  inv_x1_sg U58018 ( .A(n16090), .X(n50020) );
  inv_x1_sg U58019 ( .A(n16909), .X(n50305) );
  inv_x1_sg U58020 ( .A(n17728), .X(n50594) );
  inv_x1_sg U58021 ( .A(n18549), .X(n50881) );
  inv_x1_sg U58022 ( .A(n22604), .X(n46849) );
  inv_x1_sg U58023 ( .A(n22866), .X(n47141) );
  inv_x1_sg U58024 ( .A(n23143), .X(n47426) );
  inv_x1_sg U58025 ( .A(n23423), .X(n47711) );
  inv_x1_sg U58026 ( .A(n23702), .X(n47996) );
  inv_x1_sg U58027 ( .A(n23981), .X(n48281) );
  inv_x1_sg U58028 ( .A(n24260), .X(n48566) );
  inv_x1_sg U58029 ( .A(n24539), .X(n48851) );
  inv_x1_sg U58030 ( .A(n24817), .X(n49138) );
  inv_x1_sg U58031 ( .A(n25096), .X(n49424) );
  inv_x1_sg U58032 ( .A(n25375), .X(n49710) );
  inv_x1_sg U58033 ( .A(n25654), .X(n49996) );
  inv_x1_sg U58034 ( .A(n26196), .X(n50571) );
  inv_x1_sg U58035 ( .A(n26491), .X(n50857) );
  inv_x1_sg U58036 ( .A(n22660), .X(n46982) );
  inv_x1_sg U58037 ( .A(n22684), .X(n47072) );
  inv_x1_sg U58038 ( .A(n22610), .X(n46853) );
  inv_x1_sg U58039 ( .A(n22666), .X(n47005) );
  inv_x1_sg U58040 ( .A(n22672), .X(n47024) );
  inv_x1_sg U58041 ( .A(n22678), .X(n47054) );
  inv_x1_sg U58042 ( .A(n22873), .X(n47146) );
  inv_x1_sg U58043 ( .A(n23150), .X(n47431) );
  inv_x1_sg U58044 ( .A(n23430), .X(n47716) );
  inv_x1_sg U58045 ( .A(n23709), .X(n48001) );
  inv_x1_sg U58046 ( .A(n23988), .X(n48286) );
  inv_x1_sg U58047 ( .A(n24267), .X(n48571) );
  inv_x1_sg U58048 ( .A(n24546), .X(n48857) );
  inv_x1_sg U58049 ( .A(n24824), .X(n49144) );
  inv_x1_sg U58050 ( .A(n25103), .X(n49430) );
  inv_x1_sg U58051 ( .A(n25382), .X(n49715) );
  inv_x1_sg U58052 ( .A(n25661), .X(n50002) );
  inv_x1_sg U58053 ( .A(n25933), .X(n50289) );
  inv_x1_sg U58054 ( .A(n25945), .X(n50302) );
  inv_x1_sg U58055 ( .A(n26204), .X(n50576) );
  inv_x1_sg U58056 ( .A(n26498), .X(n50863) );
  nor_x1_sg U58057 ( .A(n6883), .B(n6884), .X(n6882) );
  nor_x1_sg U58058 ( .A(n7700), .B(n7701), .X(n7699) );
  nor_x1_sg U58059 ( .A(n8518), .B(n8519), .X(n8517) );
  nor_x1_sg U58060 ( .A(n9338), .B(n9339), .X(n9337) );
  nor_x1_sg U58061 ( .A(n10157), .B(n10158), .X(n10156) );
  nor_x1_sg U58062 ( .A(n10976), .B(n10977), .X(n10975) );
  nor_x1_sg U58063 ( .A(n11795), .B(n11796), .X(n11794) );
  nor_x1_sg U58064 ( .A(n12614), .B(n12615), .X(n12613) );
  nor_x1_sg U58065 ( .A(n13433), .B(n13434), .X(n13432) );
  nor_x1_sg U58066 ( .A(n14252), .B(n14253), .X(n14251) );
  nor_x1_sg U58067 ( .A(n15071), .B(n15072), .X(n15070) );
  nor_x1_sg U58068 ( .A(n15890), .B(n15891), .X(n15889) );
  nor_x1_sg U58069 ( .A(n17528), .B(n17529), .X(n17527) );
  nor_x1_sg U58070 ( .A(n18349), .B(n18350), .X(n18348) );
  inv_x1_sg U58071 ( .A(n7449), .X(n47029) );
  inv_x1_sg U58072 ( .A(n8267), .X(n47316) );
  inv_x1_sg U58073 ( .A(n9085), .X(n47601) );
  inv_x1_sg U58074 ( .A(n9905), .X(n47886) );
  inv_x1_sg U58075 ( .A(n10724), .X(n48171) );
  inv_x1_sg U58076 ( .A(n11543), .X(n48456) );
  inv_x1_sg U58077 ( .A(n12362), .X(n48741) );
  inv_x1_sg U58078 ( .A(n13181), .X(n49027) );
  inv_x1_sg U58079 ( .A(n14000), .X(n49314) );
  inv_x1_sg U58080 ( .A(n14819), .X(n49600) );
  inv_x1_sg U58081 ( .A(n15638), .X(n49886) );
  inv_x1_sg U58082 ( .A(n16457), .X(n50172) );
  inv_x1_sg U58083 ( .A(n17274), .X(n50457) );
  inv_x1_sg U58084 ( .A(n18095), .X(n50746) );
  inv_x1_sg U58085 ( .A(n18916), .X(n51033) );
  inv_x1_sg U58086 ( .A(n6877), .X(n46931) );
  inv_x1_sg U58087 ( .A(n7694), .X(n47223) );
  inv_x1_sg U58088 ( .A(n8512), .X(n47508) );
  inv_x1_sg U58089 ( .A(n9332), .X(n47793) );
  inv_x1_sg U58090 ( .A(n10151), .X(n48078) );
  inv_x1_sg U58091 ( .A(n10970), .X(n48363) );
  inv_x1_sg U58092 ( .A(n11789), .X(n48648) );
  inv_x1_sg U58093 ( .A(n12608), .X(n48934) );
  inv_x1_sg U58094 ( .A(n13427), .X(n49221) );
  inv_x1_sg U58095 ( .A(n14246), .X(n49507) );
  inv_x1_sg U58096 ( .A(n15065), .X(n49793) );
  inv_x1_sg U58097 ( .A(n15884), .X(n50079) );
  inv_x1_sg U58098 ( .A(n16701), .X(n50364) );
  inv_x1_sg U58099 ( .A(n17522), .X(n50653) );
  inv_x1_sg U58100 ( .A(n18343), .X(n50940) );
  nand_x1_sg U58101 ( .A(n46884), .B(n6858), .X(n7065) );
  inv_x1_sg U58102 ( .A(n6859), .X(n46884) );
  nand_x1_sg U58103 ( .A(n47177), .B(n7675), .X(n7883) );
  inv_x1_sg U58104 ( .A(n7676), .X(n47177) );
  nand_x1_sg U58105 ( .A(n47462), .B(n8493), .X(n8701) );
  inv_x1_sg U58106 ( .A(n8494), .X(n47462) );
  nand_x1_sg U58107 ( .A(n47747), .B(n9313), .X(n9521) );
  inv_x1_sg U58108 ( .A(n9314), .X(n47747) );
  nand_x1_sg U58109 ( .A(n48032), .B(n10132), .X(n10340) );
  inv_x1_sg U58110 ( .A(n10133), .X(n48032) );
  nand_x1_sg U58111 ( .A(n48317), .B(n10951), .X(n11159) );
  inv_x1_sg U58112 ( .A(n10952), .X(n48317) );
  nand_x1_sg U58113 ( .A(n48602), .B(n11770), .X(n11978) );
  inv_x1_sg U58114 ( .A(n11771), .X(n48602) );
  nand_x1_sg U58115 ( .A(n48888), .B(n12589), .X(n12797) );
  inv_x1_sg U58116 ( .A(n12590), .X(n48888) );
  nand_x1_sg U58117 ( .A(n49175), .B(n13408), .X(n13616) );
  inv_x1_sg U58118 ( .A(n13409), .X(n49175) );
  nand_x1_sg U58119 ( .A(n49461), .B(n14227), .X(n14435) );
  inv_x1_sg U58120 ( .A(n14228), .X(n49461) );
  nand_x1_sg U58121 ( .A(n49746), .B(n15046), .X(n15254) );
  inv_x1_sg U58122 ( .A(n15047), .X(n49746) );
  nand_x1_sg U58123 ( .A(n50033), .B(n15865), .X(n16073) );
  inv_x1_sg U58124 ( .A(n15866), .X(n50033) );
  nand_x1_sg U58125 ( .A(n50318), .B(n16682), .X(n16892) );
  inv_x1_sg U58126 ( .A(n16683), .X(n50318) );
  nand_x1_sg U58127 ( .A(n50607), .B(n17503), .X(n17711) );
  inv_x1_sg U58128 ( .A(n17504), .X(n50607) );
  nand_x1_sg U58129 ( .A(n50894), .B(n18324), .X(n18532) );
  inv_x1_sg U58130 ( .A(n18325), .X(n50894) );
  inv_x1_sg U58131 ( .A(n7030), .X(n47105) );
  inv_x1_sg U58132 ( .A(n7848), .X(n47391) );
  inv_x1_sg U58133 ( .A(n8666), .X(n47676) );
  inv_x1_sg U58134 ( .A(n9486), .X(n47961) );
  inv_x1_sg U58135 ( .A(n10305), .X(n48246) );
  inv_x1_sg U58136 ( .A(n11124), .X(n48531) );
  inv_x1_sg U58137 ( .A(n11943), .X(n48816) );
  inv_x1_sg U58138 ( .A(n12762), .X(n49103) );
  inv_x1_sg U58139 ( .A(n13581), .X(n49389) );
  inv_x1_sg U58140 ( .A(n14400), .X(n49675) );
  inv_x1_sg U58141 ( .A(n15219), .X(n49961) );
  inv_x1_sg U58142 ( .A(n16038), .X(n50247) );
  inv_x1_sg U58143 ( .A(n16857), .X(n50532) );
  inv_x1_sg U58144 ( .A(n17676), .X(n50821) );
  inv_x1_sg U58145 ( .A(n18497), .X(n51108) );
  nand_x1_sg U58146 ( .A(n7309), .B(n7308), .X(n7306) );
  nor_x1_sg U58147 ( .A(n7308), .B(n7309), .X(n7307) );
  nand_x1_sg U58148 ( .A(n8127), .B(n8126), .X(n8124) );
  nor_x1_sg U58149 ( .A(n8126), .B(n8127), .X(n8125) );
  nand_x1_sg U58150 ( .A(n8945), .B(n8944), .X(n8942) );
  nor_x1_sg U58151 ( .A(n8944), .B(n8945), .X(n8943) );
  nand_x1_sg U58152 ( .A(n9765), .B(n9764), .X(n9762) );
  nor_x1_sg U58153 ( .A(n9764), .B(n9765), .X(n9763) );
  nand_x1_sg U58154 ( .A(n10584), .B(n10583), .X(n10581) );
  nor_x1_sg U58155 ( .A(n10583), .B(n10584), .X(n10582) );
  nand_x1_sg U58156 ( .A(n11403), .B(n11402), .X(n11400) );
  nor_x1_sg U58157 ( .A(n11402), .B(n11403), .X(n11401) );
  nand_x1_sg U58158 ( .A(n12222), .B(n12221), .X(n12219) );
  nor_x1_sg U58159 ( .A(n12221), .B(n12222), .X(n12220) );
  nand_x1_sg U58160 ( .A(n13041), .B(n13040), .X(n13038) );
  nor_x1_sg U58161 ( .A(n13040), .B(n13041), .X(n13039) );
  nand_x1_sg U58162 ( .A(n13860), .B(n13859), .X(n13857) );
  nor_x1_sg U58163 ( .A(n13859), .B(n13860), .X(n13858) );
  nand_x1_sg U58164 ( .A(n14679), .B(n14678), .X(n14676) );
  nor_x1_sg U58165 ( .A(n14678), .B(n14679), .X(n14677) );
  nand_x1_sg U58166 ( .A(n15498), .B(n15497), .X(n15495) );
  nor_x1_sg U58167 ( .A(n15497), .B(n15498), .X(n15496) );
  nand_x1_sg U58168 ( .A(n16317), .B(n16316), .X(n16314) );
  nor_x1_sg U58169 ( .A(n16316), .B(n16317), .X(n16315) );
  nand_x1_sg U58170 ( .A(n17955), .B(n17954), .X(n17952) );
  nor_x1_sg U58171 ( .A(n17954), .B(n17955), .X(n17953) );
  nand_x1_sg U58172 ( .A(n18776), .B(n18775), .X(n18773) );
  nor_x1_sg U58173 ( .A(n18775), .B(n18776), .X(n18774) );
  nand_x1_sg U58174 ( .A(n7980), .B(n47200), .X(n7967) );
  inv_x1_sg U58175 ( .A(n7979), .X(n47200) );
  nand_x1_sg U58176 ( .A(n8798), .B(n47485), .X(n8785) );
  inv_x1_sg U58177 ( .A(n8797), .X(n47485) );
  nand_x1_sg U58178 ( .A(n9618), .B(n47770), .X(n9605) );
  inv_x1_sg U58179 ( .A(n9617), .X(n47770) );
  nand_x1_sg U58180 ( .A(n10437), .B(n48055), .X(n10424) );
  inv_x1_sg U58181 ( .A(n10436), .X(n48055) );
  nand_x1_sg U58182 ( .A(n11256), .B(n48340), .X(n11243) );
  inv_x1_sg U58183 ( .A(n11255), .X(n48340) );
  nand_x1_sg U58184 ( .A(n12075), .B(n48625), .X(n12062) );
  inv_x1_sg U58185 ( .A(n12074), .X(n48625) );
  nand_x1_sg U58186 ( .A(n12894), .B(n48911), .X(n12881) );
  inv_x1_sg U58187 ( .A(n12893), .X(n48911) );
  nand_x1_sg U58188 ( .A(n13713), .B(n49198), .X(n13700) );
  inv_x1_sg U58189 ( .A(n13712), .X(n49198) );
  nand_x1_sg U58190 ( .A(n14532), .B(n49484), .X(n14519) );
  inv_x1_sg U58191 ( .A(n14531), .X(n49484) );
  nand_x1_sg U58192 ( .A(n15351), .B(n49770), .X(n15338) );
  inv_x1_sg U58193 ( .A(n15350), .X(n49770) );
  nand_x1_sg U58194 ( .A(n16170), .B(n50056), .X(n16157) );
  inv_x1_sg U58195 ( .A(n16169), .X(n50056) );
  nand_x1_sg U58196 ( .A(n18629), .B(n50917), .X(n18616) );
  inv_x1_sg U58197 ( .A(n18628), .X(n50917) );
  nand_x1_sg U58198 ( .A(n16986), .B(n50341), .X(n16974) );
  inv_x1_sg U58199 ( .A(n16985), .X(n50341) );
  nand_x1_sg U58200 ( .A(n17808), .B(n50630), .X(n17795) );
  inv_x1_sg U58201 ( .A(n17807), .X(n50630) );
  nand_x1_sg U58202 ( .A(n7161), .B(n46907), .X(n7149) );
  inv_x1_sg U58203 ( .A(n7160), .X(n46907) );
  nand_x1_sg U58204 ( .A(n7211), .B(n46916), .X(n7202) );
  inv_x1_sg U58205 ( .A(n7192), .X(n46918) );
  nand_x1_sg U58206 ( .A(n17036), .B(n50349), .X(n17027) );
  inv_x1_sg U58207 ( .A(n17017), .X(n50351) );
  nand_x1_sg U58208 ( .A(n8030), .B(n47208), .X(n8021) );
  inv_x1_sg U58209 ( .A(n8011), .X(n47210) );
  nand_x1_sg U58210 ( .A(n8848), .B(n47493), .X(n8839) );
  inv_x1_sg U58211 ( .A(n8829), .X(n47495) );
  nand_x1_sg U58212 ( .A(n9668), .B(n47778), .X(n9659) );
  inv_x1_sg U58213 ( .A(n9649), .X(n47780) );
  nand_x1_sg U58214 ( .A(n10487), .B(n48063), .X(n10478) );
  inv_x1_sg U58215 ( .A(n10468), .X(n48065) );
  nand_x1_sg U58216 ( .A(n11306), .B(n48348), .X(n11297) );
  inv_x1_sg U58217 ( .A(n11287), .X(n48350) );
  nand_x1_sg U58218 ( .A(n12125), .B(n48633), .X(n12116) );
  inv_x1_sg U58219 ( .A(n12106), .X(n48635) );
  nand_x1_sg U58220 ( .A(n12944), .B(n48919), .X(n12935) );
  inv_x1_sg U58221 ( .A(n12925), .X(n48921) );
  nand_x1_sg U58222 ( .A(n13763), .B(n49206), .X(n13754) );
  inv_x1_sg U58223 ( .A(n13744), .X(n49208) );
  nand_x1_sg U58224 ( .A(n14582), .B(n49492), .X(n14573) );
  inv_x1_sg U58225 ( .A(n14563), .X(n49494) );
  nand_x1_sg U58226 ( .A(n15401), .B(n49778), .X(n15392) );
  inv_x1_sg U58227 ( .A(n15382), .X(n49780) );
  nand_x1_sg U58228 ( .A(n16220), .B(n50064), .X(n16211) );
  inv_x1_sg U58229 ( .A(n16201), .X(n50066) );
  nand_x1_sg U58230 ( .A(n18679), .B(n50925), .X(n18670) );
  inv_x1_sg U58231 ( .A(n18660), .X(n50927) );
  nand_x1_sg U58232 ( .A(n17858), .B(n50638), .X(n17849) );
  inv_x1_sg U58233 ( .A(n17839), .X(n50640) );
  nand_x1_sg U58234 ( .A(n16785), .B(n16786), .X(n17413) );
  nor_x1_sg U58235 ( .A(n16785), .B(n16786), .X(n17414) );
  nand_x1_sg U58236 ( .A(n8069), .B(n8068), .X(n8065) );
  nand_x1_sg U58237 ( .A(n8887), .B(n8886), .X(n8883) );
  nand_x1_sg U58238 ( .A(n9707), .B(n9706), .X(n9703) );
  nand_x1_sg U58239 ( .A(n10526), .B(n10525), .X(n10522) );
  nand_x1_sg U58240 ( .A(n11345), .B(n11344), .X(n11341) );
  nand_x1_sg U58241 ( .A(n12164), .B(n12163), .X(n12160) );
  nand_x1_sg U58242 ( .A(n12983), .B(n12982), .X(n12979) );
  nand_x1_sg U58243 ( .A(n13802), .B(n13801), .X(n13798) );
  nand_x1_sg U58244 ( .A(n14621), .B(n14620), .X(n14617) );
  nand_x1_sg U58245 ( .A(n15440), .B(n15439), .X(n15436) );
  nand_x1_sg U58246 ( .A(n16259), .B(n16258), .X(n16255) );
  nand_x1_sg U58247 ( .A(n18718), .B(n18717), .X(n18714) );
  nand_x1_sg U58248 ( .A(n17075), .B(n17074), .X(n17071) );
  nand_x1_sg U58249 ( .A(n17897), .B(n17896), .X(n17893) );
  nand_x1_sg U58250 ( .A(n6961), .B(n6962), .X(n7588) );
  nor_x1_sg U58251 ( .A(n6961), .B(n6962), .X(n7589) );
  nand_x1_sg U58252 ( .A(n7250), .B(n7249), .X(n7246) );
  nand_x1_sg U58253 ( .A(n6979), .B(n6978), .X(n6976) );
  nor_x1_sg U58254 ( .A(n6978), .B(n6979), .X(n6977) );
  nand_x1_sg U58255 ( .A(n7796), .B(n7795), .X(n7793) );
  nor_x1_sg U58256 ( .A(n7795), .B(n7796), .X(n7794) );
  nand_x1_sg U58257 ( .A(n8614), .B(n8613), .X(n8611) );
  nor_x1_sg U58258 ( .A(n8613), .B(n8614), .X(n8612) );
  nand_x1_sg U58259 ( .A(n9434), .B(n9433), .X(n9431) );
  nor_x1_sg U58260 ( .A(n9433), .B(n9434), .X(n9432) );
  nand_x1_sg U58261 ( .A(n10253), .B(n10252), .X(n10250) );
  nor_x1_sg U58262 ( .A(n10252), .B(n10253), .X(n10251) );
  nand_x1_sg U58263 ( .A(n11072), .B(n11071), .X(n11069) );
  nor_x1_sg U58264 ( .A(n11071), .B(n11072), .X(n11070) );
  nand_x1_sg U58265 ( .A(n11891), .B(n11890), .X(n11888) );
  nor_x1_sg U58266 ( .A(n11890), .B(n11891), .X(n11889) );
  nand_x1_sg U58267 ( .A(n12710), .B(n12709), .X(n12707) );
  nor_x1_sg U58268 ( .A(n12709), .B(n12710), .X(n12708) );
  nand_x1_sg U58269 ( .A(n13529), .B(n13528), .X(n13526) );
  nor_x1_sg U58270 ( .A(n13528), .B(n13529), .X(n13527) );
  nand_x1_sg U58271 ( .A(n14348), .B(n14347), .X(n14345) );
  nor_x1_sg U58272 ( .A(n14347), .B(n14348), .X(n14346) );
  nand_x1_sg U58273 ( .A(n15167), .B(n15166), .X(n15164) );
  nor_x1_sg U58274 ( .A(n15166), .B(n15167), .X(n15165) );
  nand_x1_sg U58275 ( .A(n15986), .B(n15985), .X(n15983) );
  nor_x1_sg U58276 ( .A(n15985), .B(n15986), .X(n15984) );
  nand_x1_sg U58277 ( .A(n16803), .B(n16802), .X(n16800) );
  nor_x1_sg U58278 ( .A(n16802), .B(n16803), .X(n16801) );
  nand_x1_sg U58279 ( .A(n17624), .B(n17623), .X(n17621) );
  nor_x1_sg U58280 ( .A(n17623), .B(n17624), .X(n17622) );
  nand_x1_sg U58281 ( .A(n18445), .B(n18444), .X(n18442) );
  nor_x1_sg U58282 ( .A(n18444), .B(n18445), .X(n18443) );
  nand_x1_sg U58283 ( .A(n50423), .B(n17154), .X(n17150) );
  inv_x1_sg U58284 ( .A(n17133), .X(n50424) );
  inv_x1_sg U58285 ( .A(n7250), .X(n46922) );
  inv_x1_sg U58286 ( .A(n17075), .X(n50355) );
  inv_x1_sg U58287 ( .A(n8069), .X(n47214) );
  inv_x1_sg U58288 ( .A(n8887), .X(n47499) );
  inv_x1_sg U58289 ( .A(n9707), .X(n47784) );
  inv_x1_sg U58290 ( .A(n10526), .X(n48069) );
  inv_x1_sg U58291 ( .A(n11345), .X(n48354) );
  inv_x1_sg U58292 ( .A(n12164), .X(n48639) );
  inv_x1_sg U58293 ( .A(n12983), .X(n48925) );
  inv_x1_sg U58294 ( .A(n13802), .X(n49212) );
  inv_x1_sg U58295 ( .A(n14621), .X(n49498) );
  inv_x1_sg U58296 ( .A(n15440), .X(n49784) );
  inv_x1_sg U58297 ( .A(n16259), .X(n50070) );
  inv_x1_sg U58298 ( .A(n17897), .X(n50644) );
  inv_x1_sg U58299 ( .A(n18718), .X(n50931) );
  nand_x1_sg U58300 ( .A(n46959), .B(n46971), .X(n7387) );
  nand_x1_sg U58301 ( .A(n7388), .B(n7389), .X(n7386) );
  nand_x1_sg U58302 ( .A(n50391), .B(n50402), .X(n17212) );
  nand_x1_sg U58303 ( .A(n17213), .B(n17214), .X(n17211) );
  nand_x1_sg U58304 ( .A(n7401), .B(n7400), .X(n7419) );
  nand_x1_sg U58305 ( .A(n8219), .B(n8218), .X(n8237) );
  nand_x1_sg U58306 ( .A(n9037), .B(n9036), .X(n9055) );
  nand_x1_sg U58307 ( .A(n9857), .B(n9856), .X(n9875) );
  nand_x1_sg U58308 ( .A(n10676), .B(n10675), .X(n10694) );
  nand_x1_sg U58309 ( .A(n11495), .B(n11494), .X(n11513) );
  nand_x1_sg U58310 ( .A(n12314), .B(n12313), .X(n12332) );
  nand_x1_sg U58311 ( .A(n13133), .B(n13132), .X(n13151) );
  nand_x1_sg U58312 ( .A(n13952), .B(n13951), .X(n13970) );
  nand_x1_sg U58313 ( .A(n14771), .B(n14770), .X(n14789) );
  nand_x1_sg U58314 ( .A(n15590), .B(n15589), .X(n15608) );
  nand_x1_sg U58315 ( .A(n16409), .B(n16408), .X(n16427) );
  nand_x1_sg U58316 ( .A(n17226), .B(n17225), .X(n17244) );
  nand_x1_sg U58317 ( .A(n18047), .B(n18046), .X(n18065) );
  nand_x1_sg U58318 ( .A(n18868), .B(n18867), .X(n18886) );
  nand_x1_sg U58319 ( .A(n7221), .B(n7220), .X(n7218) );
  nor_x1_sg U58320 ( .A(n7220), .B(n7221), .X(n7219) );
  nand_x1_sg U58321 ( .A(n8040), .B(n8039), .X(n8037) );
  nor_x1_sg U58322 ( .A(n8039), .B(n8040), .X(n8038) );
  nand_x1_sg U58323 ( .A(n8858), .B(n8857), .X(n8855) );
  nor_x1_sg U58324 ( .A(n8857), .B(n8858), .X(n8856) );
  nand_x1_sg U58325 ( .A(n9678), .B(n9677), .X(n9675) );
  nor_x1_sg U58326 ( .A(n9677), .B(n9678), .X(n9676) );
  nand_x1_sg U58327 ( .A(n10497), .B(n10496), .X(n10494) );
  nor_x1_sg U58328 ( .A(n10496), .B(n10497), .X(n10495) );
  nand_x1_sg U58329 ( .A(n11316), .B(n11315), .X(n11313) );
  nor_x1_sg U58330 ( .A(n11315), .B(n11316), .X(n11314) );
  nand_x1_sg U58331 ( .A(n12135), .B(n12134), .X(n12132) );
  nor_x1_sg U58332 ( .A(n12134), .B(n12135), .X(n12133) );
  nand_x1_sg U58333 ( .A(n12954), .B(n12953), .X(n12951) );
  nor_x1_sg U58334 ( .A(n12953), .B(n12954), .X(n12952) );
  nand_x1_sg U58335 ( .A(n13773), .B(n13772), .X(n13770) );
  nor_x1_sg U58336 ( .A(n13772), .B(n13773), .X(n13771) );
  nand_x1_sg U58337 ( .A(n14592), .B(n14591), .X(n14589) );
  nor_x1_sg U58338 ( .A(n14591), .B(n14592), .X(n14590) );
  nand_x1_sg U58339 ( .A(n15411), .B(n15410), .X(n15408) );
  nor_x1_sg U58340 ( .A(n15410), .B(n15411), .X(n15409) );
  nand_x1_sg U58341 ( .A(n16230), .B(n16229), .X(n16227) );
  nor_x1_sg U58342 ( .A(n16229), .B(n16230), .X(n16228) );
  nand_x1_sg U58343 ( .A(n17046), .B(n17045), .X(n17043) );
  nor_x1_sg U58344 ( .A(n17045), .B(n17046), .X(n17044) );
  nand_x1_sg U58345 ( .A(n17868), .B(n17867), .X(n17865) );
  nor_x1_sg U58346 ( .A(n17867), .B(n17868), .X(n17866) );
  nand_x1_sg U58347 ( .A(n18689), .B(n18688), .X(n18686) );
  nor_x1_sg U58348 ( .A(n18688), .B(n18689), .X(n18687) );
  inv_x1_sg U58349 ( .A(n7221), .X(n46947) );
  inv_x1_sg U58350 ( .A(n8040), .X(n47238) );
  inv_x1_sg U58351 ( .A(n8858), .X(n47523) );
  inv_x1_sg U58352 ( .A(n9678), .X(n47808) );
  inv_x1_sg U58353 ( .A(n10497), .X(n48093) );
  inv_x1_sg U58354 ( .A(n11316), .X(n48378) );
  inv_x1_sg U58355 ( .A(n12135), .X(n48663) );
  inv_x1_sg U58356 ( .A(n12954), .X(n48949) );
  inv_x1_sg U58357 ( .A(n13773), .X(n49236) );
  inv_x1_sg U58358 ( .A(n14592), .X(n49522) );
  inv_x1_sg U58359 ( .A(n15411), .X(n49808) );
  inv_x1_sg U58360 ( .A(n16230), .X(n50094) );
  inv_x1_sg U58361 ( .A(n17046), .X(n50379) );
  inv_x1_sg U58362 ( .A(n17868), .X(n50668) );
  inv_x1_sg U58363 ( .A(n18689), .X(n50955) );
  nand_x1_sg U58364 ( .A(n16999), .B(n16998), .X(n16996) );
  nor_x1_sg U58365 ( .A(n16998), .B(n16999), .X(n16997) );
  nand_x1_sg U58366 ( .A(n8374), .B(n8373), .X(n8371) );
  nor_x1_sg U58367 ( .A(n8373), .B(n8374), .X(n8372) );
  nand_x1_sg U58368 ( .A(n9192), .B(n9191), .X(n9189) );
  nor_x1_sg U58369 ( .A(n9191), .B(n9192), .X(n9190) );
  nand_x1_sg U58370 ( .A(n10012), .B(n10011), .X(n10009) );
  nor_x1_sg U58371 ( .A(n10011), .B(n10012), .X(n10010) );
  nand_x1_sg U58372 ( .A(n10831), .B(n10830), .X(n10828) );
  nor_x1_sg U58373 ( .A(n10830), .B(n10831), .X(n10829) );
  nand_x1_sg U58374 ( .A(n11650), .B(n11649), .X(n11647) );
  nor_x1_sg U58375 ( .A(n11649), .B(n11650), .X(n11648) );
  nand_x1_sg U58376 ( .A(n12469), .B(n12468), .X(n12466) );
  nor_x1_sg U58377 ( .A(n12468), .B(n12469), .X(n12467) );
  nand_x1_sg U58378 ( .A(n13288), .B(n13287), .X(n13285) );
  nor_x1_sg U58379 ( .A(n13287), .B(n13288), .X(n13286) );
  nand_x1_sg U58380 ( .A(n14107), .B(n14106), .X(n14104) );
  nor_x1_sg U58381 ( .A(n14106), .B(n14107), .X(n14105) );
  nand_x1_sg U58382 ( .A(n14926), .B(n14925), .X(n14923) );
  nor_x1_sg U58383 ( .A(n14925), .B(n14926), .X(n14924) );
  nand_x1_sg U58384 ( .A(n15745), .B(n15744), .X(n15742) );
  nor_x1_sg U58385 ( .A(n15744), .B(n15745), .X(n15743) );
  nand_x1_sg U58386 ( .A(n16564), .B(n16563), .X(n16561) );
  nor_x1_sg U58387 ( .A(n16563), .B(n16564), .X(n16562) );
  nand_x1_sg U58388 ( .A(n17381), .B(n17380), .X(n17378) );
  nor_x1_sg U58389 ( .A(n17380), .B(n17381), .X(n17379) );
  nand_x1_sg U58390 ( .A(n18202), .B(n18201), .X(n18199) );
  nor_x1_sg U58391 ( .A(n18201), .B(n18202), .X(n18200) );
  nand_x1_sg U58392 ( .A(n19023), .B(n19022), .X(n19020) );
  nor_x1_sg U58393 ( .A(n19022), .B(n19023), .X(n19021) );
  inv_x1_sg U58394 ( .A(n8374), .X(n47338) );
  inv_x1_sg U58395 ( .A(n9192), .X(n47623) );
  inv_x1_sg U58396 ( .A(n10012), .X(n47908) );
  inv_x1_sg U58397 ( .A(n10831), .X(n48193) );
  inv_x1_sg U58398 ( .A(n11650), .X(n48478) );
  inv_x1_sg U58399 ( .A(n12469), .X(n48763) );
  inv_x1_sg U58400 ( .A(n13288), .X(n49049) );
  inv_x1_sg U58401 ( .A(n14107), .X(n49336) );
  inv_x1_sg U58402 ( .A(n14926), .X(n49622) );
  inv_x1_sg U58403 ( .A(n15745), .X(n49908) );
  inv_x1_sg U58404 ( .A(n16564), .X(n50194) );
  inv_x1_sg U58405 ( .A(n17381), .X(n50479) );
  inv_x1_sg U58406 ( .A(n18202), .X(n50768) );
  inv_x1_sg U58407 ( .A(n19023), .X(n51055) );
  nand_x1_sg U58408 ( .A(n7556), .B(n7555), .X(n7553) );
  nor_x1_sg U58409 ( .A(n7555), .B(n7556), .X(n7554) );
  inv_x1_sg U58410 ( .A(n7556), .X(n47051) );
  nand_x1_sg U58411 ( .A(n7449), .B(n7448), .X(n7446) );
  nor_x1_sg U58412 ( .A(n7448), .B(n7449), .X(n7447) );
  nand_x1_sg U58413 ( .A(n8267), .B(n8266), .X(n8264) );
  nor_x1_sg U58414 ( .A(n8266), .B(n8267), .X(n8265) );
  nand_x1_sg U58415 ( .A(n9085), .B(n9084), .X(n9082) );
  nor_x1_sg U58416 ( .A(n9084), .B(n9085), .X(n9083) );
  nand_x1_sg U58417 ( .A(n9905), .B(n9904), .X(n9902) );
  nor_x1_sg U58418 ( .A(n9904), .B(n9905), .X(n9903) );
  nand_x1_sg U58419 ( .A(n10724), .B(n10723), .X(n10721) );
  nor_x1_sg U58420 ( .A(n10723), .B(n10724), .X(n10722) );
  nand_x1_sg U58421 ( .A(n11543), .B(n11542), .X(n11540) );
  nor_x1_sg U58422 ( .A(n11542), .B(n11543), .X(n11541) );
  nand_x1_sg U58423 ( .A(n12362), .B(n12361), .X(n12359) );
  nor_x1_sg U58424 ( .A(n12361), .B(n12362), .X(n12360) );
  nand_x1_sg U58425 ( .A(n13181), .B(n13180), .X(n13178) );
  nor_x1_sg U58426 ( .A(n13180), .B(n13181), .X(n13179) );
  nand_x1_sg U58427 ( .A(n14000), .B(n13999), .X(n13997) );
  nor_x1_sg U58428 ( .A(n13999), .B(n14000), .X(n13998) );
  nand_x1_sg U58429 ( .A(n14819), .B(n14818), .X(n14816) );
  nor_x1_sg U58430 ( .A(n14818), .B(n14819), .X(n14817) );
  nand_x1_sg U58431 ( .A(n15638), .B(n15637), .X(n15635) );
  nor_x1_sg U58432 ( .A(n15637), .B(n15638), .X(n15636) );
  nand_x1_sg U58433 ( .A(n16457), .B(n16456), .X(n16454) );
  nor_x1_sg U58434 ( .A(n16456), .B(n16457), .X(n16455) );
  nand_x1_sg U58435 ( .A(n17274), .B(n17273), .X(n17271) );
  nor_x1_sg U58436 ( .A(n17273), .B(n17274), .X(n17272) );
  nand_x1_sg U58437 ( .A(n18095), .B(n18094), .X(n18092) );
  nor_x1_sg U58438 ( .A(n18094), .B(n18095), .X(n18093) );
  nand_x1_sg U58439 ( .A(n18916), .B(n18915), .X(n18913) );
  nor_x1_sg U58440 ( .A(n18915), .B(n18916), .X(n18914) );
  nand_x1_sg U58441 ( .A(n7540), .B(n47083), .X(n7538) );
  nor_x1_sg U58442 ( .A(n47083), .B(n7540), .X(n7539) );
  nand_x1_sg U58443 ( .A(n8358), .B(n47369), .X(n8356) );
  nor_x1_sg U58444 ( .A(n47369), .B(n8358), .X(n8357) );
  nand_x1_sg U58445 ( .A(n9176), .B(n47654), .X(n9174) );
  nor_x1_sg U58446 ( .A(n47654), .B(n9176), .X(n9175) );
  nand_x1_sg U58447 ( .A(n9996), .B(n47939), .X(n9994) );
  nor_x1_sg U58448 ( .A(n47939), .B(n9996), .X(n9995) );
  nand_x1_sg U58449 ( .A(n10815), .B(n48224), .X(n10813) );
  nor_x1_sg U58450 ( .A(n48224), .B(n10815), .X(n10814) );
  nand_x1_sg U58451 ( .A(n11634), .B(n48509), .X(n11632) );
  nor_x1_sg U58452 ( .A(n48509), .B(n11634), .X(n11633) );
  nand_x1_sg U58453 ( .A(n12453), .B(n48794), .X(n12451) );
  nor_x1_sg U58454 ( .A(n48794), .B(n12453), .X(n12452) );
  nand_x1_sg U58455 ( .A(n13272), .B(n49081), .X(n13270) );
  nor_x1_sg U58456 ( .A(n49081), .B(n13272), .X(n13271) );
  nand_x1_sg U58457 ( .A(n14091), .B(n49367), .X(n14089) );
  nor_x1_sg U58458 ( .A(n49367), .B(n14091), .X(n14090) );
  nand_x1_sg U58459 ( .A(n14910), .B(n49653), .X(n14908) );
  nor_x1_sg U58460 ( .A(n49653), .B(n14910), .X(n14909) );
  nand_x1_sg U58461 ( .A(n15729), .B(n49939), .X(n15727) );
  nor_x1_sg U58462 ( .A(n49939), .B(n15729), .X(n15728) );
  nand_x1_sg U58463 ( .A(n16548), .B(n50225), .X(n16546) );
  nor_x1_sg U58464 ( .A(n50225), .B(n16548), .X(n16547) );
  nand_x1_sg U58465 ( .A(n17365), .B(n50510), .X(n17363) );
  nor_x1_sg U58466 ( .A(n50510), .B(n17365), .X(n17364) );
  nand_x1_sg U58467 ( .A(n18186), .B(n50799), .X(n18184) );
  nor_x1_sg U58468 ( .A(n50799), .B(n18186), .X(n18185) );
  nand_x1_sg U58469 ( .A(n19007), .B(n51086), .X(n19005) );
  nor_x1_sg U58470 ( .A(n51086), .B(n19007), .X(n19006) );
  nand_x1_sg U58471 ( .A(n7249), .B(n46922), .X(n7247) );
  nor_x1_sg U58472 ( .A(n7249), .B(n46922), .X(n7248) );
  nand_x1_sg U58473 ( .A(n8068), .B(n47214), .X(n8066) );
  nor_x1_sg U58474 ( .A(n8068), .B(n47214), .X(n8067) );
  nand_x1_sg U58475 ( .A(n8886), .B(n47499), .X(n8884) );
  nor_x1_sg U58476 ( .A(n8886), .B(n47499), .X(n8885) );
  nand_x1_sg U58477 ( .A(n9706), .B(n47784), .X(n9704) );
  nor_x1_sg U58478 ( .A(n9706), .B(n47784), .X(n9705) );
  nand_x1_sg U58479 ( .A(n10525), .B(n48069), .X(n10523) );
  nor_x1_sg U58480 ( .A(n10525), .B(n48069), .X(n10524) );
  nand_x1_sg U58481 ( .A(n11344), .B(n48354), .X(n11342) );
  nor_x1_sg U58482 ( .A(n11344), .B(n48354), .X(n11343) );
  nand_x1_sg U58483 ( .A(n12163), .B(n48639), .X(n12161) );
  nor_x1_sg U58484 ( .A(n12163), .B(n48639), .X(n12162) );
  nand_x1_sg U58485 ( .A(n12982), .B(n48925), .X(n12980) );
  nor_x1_sg U58486 ( .A(n12982), .B(n48925), .X(n12981) );
  nand_x1_sg U58487 ( .A(n13801), .B(n49212), .X(n13799) );
  nor_x1_sg U58488 ( .A(n13801), .B(n49212), .X(n13800) );
  nand_x1_sg U58489 ( .A(n14620), .B(n49498), .X(n14618) );
  nor_x1_sg U58490 ( .A(n14620), .B(n49498), .X(n14619) );
  nand_x1_sg U58491 ( .A(n15439), .B(n49784), .X(n15437) );
  nor_x1_sg U58492 ( .A(n15439), .B(n49784), .X(n15438) );
  nand_x1_sg U58493 ( .A(n16258), .B(n50070), .X(n16256) );
  nor_x1_sg U58494 ( .A(n16258), .B(n50070), .X(n16257) );
  nand_x1_sg U58495 ( .A(n17074), .B(n50355), .X(n17072) );
  nor_x1_sg U58496 ( .A(n17074), .B(n50355), .X(n17073) );
  nand_x1_sg U58497 ( .A(n17896), .B(n50644), .X(n17894) );
  nor_x1_sg U58498 ( .A(n17896), .B(n50644), .X(n17895) );
  nand_x1_sg U58499 ( .A(n18717), .B(n50931), .X(n18715) );
  nor_x1_sg U58500 ( .A(n18717), .B(n50931), .X(n18716) );
  nand_x1_sg U58501 ( .A(n47045), .B(n46940), .X(n6959) );
  inv_x1_sg U58502 ( .A(n6962), .X(n46961) );
  nand_x1_sg U58503 ( .A(n50473), .B(n50372), .X(n16783) );
  inv_x1_sg U58504 ( .A(n16786), .X(n50393) );
  nand_x1_sg U58505 ( .A(n46970), .B(n47004), .X(n7355) );
  nand_x1_sg U58506 ( .A(n7357), .B(n7358), .X(n7356) );
  nand_x1_sg U58507 ( .A(n47260), .B(n47293), .X(n8173) );
  nand_x1_sg U58508 ( .A(n8175), .B(n8176), .X(n8174) );
  nand_x1_sg U58509 ( .A(n47545), .B(n47578), .X(n8991) );
  nand_x1_sg U58510 ( .A(n8993), .B(n8994), .X(n8992) );
  nand_x1_sg U58511 ( .A(n47830), .B(n47863), .X(n9811) );
  nand_x1_sg U58512 ( .A(n9813), .B(n9814), .X(n9812) );
  nand_x1_sg U58513 ( .A(n48115), .B(n48148), .X(n10630) );
  nand_x1_sg U58514 ( .A(n10632), .B(n10633), .X(n10631) );
  nand_x1_sg U58515 ( .A(n48400), .B(n48433), .X(n11449) );
  nand_x1_sg U58516 ( .A(n11451), .B(n11452), .X(n11450) );
  nand_x1_sg U58517 ( .A(n48685), .B(n48718), .X(n12268) );
  nand_x1_sg U58518 ( .A(n12270), .B(n12271), .X(n12269) );
  nand_x1_sg U58519 ( .A(n48971), .B(n49004), .X(n13087) );
  nand_x1_sg U58520 ( .A(n13089), .B(n13090), .X(n13088) );
  nand_x1_sg U58521 ( .A(n49258), .B(n49291), .X(n13906) );
  nand_x1_sg U58522 ( .A(n13908), .B(n13909), .X(n13907) );
  nand_x1_sg U58523 ( .A(n49544), .B(n49577), .X(n14725) );
  nand_x1_sg U58524 ( .A(n14727), .B(n14728), .X(n14726) );
  nand_x1_sg U58525 ( .A(n49830), .B(n49863), .X(n15544) );
  nand_x1_sg U58526 ( .A(n15546), .B(n15547), .X(n15545) );
  nand_x1_sg U58527 ( .A(n50116), .B(n50149), .X(n16363) );
  nand_x1_sg U58528 ( .A(n16365), .B(n16366), .X(n16364) );
  nand_x1_sg U58529 ( .A(n50401), .B(n50434), .X(n17180) );
  nand_x1_sg U58530 ( .A(n17182), .B(n17183), .X(n17181) );
  nand_x1_sg U58531 ( .A(n50690), .B(n50723), .X(n18001) );
  nand_x1_sg U58532 ( .A(n18003), .B(n18004), .X(n18002) );
  nand_x1_sg U58533 ( .A(n50977), .B(n51010), .X(n18822) );
  nand_x1_sg U58534 ( .A(n18824), .B(n18825), .X(n18823) );
  nand_x1_sg U58535 ( .A(n7160), .B(n7161), .X(n7159) );
  nor_x1_sg U58536 ( .A(n7160), .B(n7161), .X(n7162) );
  nand_x1_sg U58537 ( .A(n7979), .B(n7980), .X(n7978) );
  nor_x1_sg U58538 ( .A(n7979), .B(n7980), .X(n7981) );
  nand_x1_sg U58539 ( .A(n8797), .B(n8798), .X(n8796) );
  nor_x1_sg U58540 ( .A(n8797), .B(n8798), .X(n8799) );
  nand_x1_sg U58541 ( .A(n9617), .B(n9618), .X(n9616) );
  nor_x1_sg U58542 ( .A(n9617), .B(n9618), .X(n9619) );
  nand_x1_sg U58543 ( .A(n10436), .B(n10437), .X(n10435) );
  nor_x1_sg U58544 ( .A(n10436), .B(n10437), .X(n10438) );
  nand_x1_sg U58545 ( .A(n11255), .B(n11256), .X(n11254) );
  nor_x1_sg U58546 ( .A(n11255), .B(n11256), .X(n11257) );
  nand_x1_sg U58547 ( .A(n12074), .B(n12075), .X(n12073) );
  nor_x1_sg U58548 ( .A(n12074), .B(n12075), .X(n12076) );
  nand_x1_sg U58549 ( .A(n12893), .B(n12894), .X(n12892) );
  nor_x1_sg U58550 ( .A(n12893), .B(n12894), .X(n12895) );
  nand_x1_sg U58551 ( .A(n13712), .B(n13713), .X(n13711) );
  nor_x1_sg U58552 ( .A(n13712), .B(n13713), .X(n13714) );
  nand_x1_sg U58553 ( .A(n14531), .B(n14532), .X(n14530) );
  nor_x1_sg U58554 ( .A(n14531), .B(n14532), .X(n14533) );
  nand_x1_sg U58555 ( .A(n15350), .B(n15351), .X(n15349) );
  nor_x1_sg U58556 ( .A(n15350), .B(n15351), .X(n15352) );
  nand_x1_sg U58557 ( .A(n16169), .B(n16170), .X(n16168) );
  nor_x1_sg U58558 ( .A(n16169), .B(n16170), .X(n16171) );
  nand_x1_sg U58559 ( .A(n16985), .B(n16986), .X(n16984) );
  nor_x1_sg U58560 ( .A(n16985), .B(n16986), .X(n16987) );
  nand_x1_sg U58561 ( .A(n17807), .B(n17808), .X(n17806) );
  nor_x1_sg U58562 ( .A(n17807), .B(n17808), .X(n17809) );
  nand_x1_sg U58563 ( .A(n18628), .B(n18629), .X(n18627) );
  nor_x1_sg U58564 ( .A(n18628), .B(n18629), .X(n18630) );
  nand_x1_sg U58565 ( .A(n7191), .B(n7192), .X(n7190) );
  nor_x1_sg U58566 ( .A(n7192), .B(n7191), .X(n7193) );
  nand_x1_sg U58567 ( .A(n8010), .B(n8011), .X(n8009) );
  nor_x1_sg U58568 ( .A(n8011), .B(n8010), .X(n8012) );
  nand_x1_sg U58569 ( .A(n8828), .B(n8829), .X(n8827) );
  nor_x1_sg U58570 ( .A(n8829), .B(n8828), .X(n8830) );
  nand_x1_sg U58571 ( .A(n9648), .B(n9649), .X(n9647) );
  nor_x1_sg U58572 ( .A(n9649), .B(n9648), .X(n9650) );
  nand_x1_sg U58573 ( .A(n10467), .B(n10468), .X(n10466) );
  nor_x1_sg U58574 ( .A(n10468), .B(n10467), .X(n10469) );
  nand_x1_sg U58575 ( .A(n11286), .B(n11287), .X(n11285) );
  nor_x1_sg U58576 ( .A(n11287), .B(n11286), .X(n11288) );
  nand_x1_sg U58577 ( .A(n12105), .B(n12106), .X(n12104) );
  nor_x1_sg U58578 ( .A(n12106), .B(n12105), .X(n12107) );
  nand_x1_sg U58579 ( .A(n12924), .B(n12925), .X(n12923) );
  nor_x1_sg U58580 ( .A(n12925), .B(n12924), .X(n12926) );
  nand_x1_sg U58581 ( .A(n13743), .B(n13744), .X(n13742) );
  nor_x1_sg U58582 ( .A(n13744), .B(n13743), .X(n13745) );
  nand_x1_sg U58583 ( .A(n14562), .B(n14563), .X(n14561) );
  nor_x1_sg U58584 ( .A(n14563), .B(n14562), .X(n14564) );
  nand_x1_sg U58585 ( .A(n15381), .B(n15382), .X(n15380) );
  nor_x1_sg U58586 ( .A(n15382), .B(n15381), .X(n15383) );
  nand_x1_sg U58587 ( .A(n16200), .B(n16201), .X(n16199) );
  nor_x1_sg U58588 ( .A(n16201), .B(n16200), .X(n16202) );
  nand_x1_sg U58589 ( .A(n17016), .B(n17017), .X(n17015) );
  nor_x1_sg U58590 ( .A(n17017), .B(n17016), .X(n17018) );
  nand_x1_sg U58591 ( .A(n17838), .B(n17839), .X(n17837) );
  nor_x1_sg U58592 ( .A(n17839), .B(n17838), .X(n17840) );
  nand_x1_sg U58593 ( .A(n18659), .B(n18660), .X(n18658) );
  nor_x1_sg U58594 ( .A(n18660), .B(n18659), .X(n18661) );
  nand_x1_sg U58595 ( .A(n7511), .B(n7512), .X(n7510) );
  nor_x1_sg U58596 ( .A(n7512), .B(n7511), .X(n7513) );
  nand_x1_sg U58597 ( .A(n8329), .B(n8330), .X(n8328) );
  nor_x1_sg U58598 ( .A(n8330), .B(n8329), .X(n8331) );
  nand_x1_sg U58599 ( .A(n9147), .B(n9148), .X(n9146) );
  nor_x1_sg U58600 ( .A(n9148), .B(n9147), .X(n9149) );
  nand_x1_sg U58601 ( .A(n9967), .B(n9968), .X(n9966) );
  nor_x1_sg U58602 ( .A(n9968), .B(n9967), .X(n9969) );
  nand_x1_sg U58603 ( .A(n10786), .B(n10787), .X(n10785) );
  nor_x1_sg U58604 ( .A(n10787), .B(n10786), .X(n10788) );
  nand_x1_sg U58605 ( .A(n11605), .B(n11606), .X(n11604) );
  nor_x1_sg U58606 ( .A(n11606), .B(n11605), .X(n11607) );
  nand_x1_sg U58607 ( .A(n12424), .B(n12425), .X(n12423) );
  nor_x1_sg U58608 ( .A(n12425), .B(n12424), .X(n12426) );
  nand_x1_sg U58609 ( .A(n13243), .B(n13244), .X(n13242) );
  nor_x1_sg U58610 ( .A(n13244), .B(n13243), .X(n13245) );
  nand_x1_sg U58611 ( .A(n14062), .B(n14063), .X(n14061) );
  nor_x1_sg U58612 ( .A(n14063), .B(n14062), .X(n14064) );
  nand_x1_sg U58613 ( .A(n14881), .B(n14882), .X(n14880) );
  nor_x1_sg U58614 ( .A(n14882), .B(n14881), .X(n14883) );
  nand_x1_sg U58615 ( .A(n15700), .B(n15701), .X(n15699) );
  nor_x1_sg U58616 ( .A(n15701), .B(n15700), .X(n15702) );
  nand_x1_sg U58617 ( .A(n16519), .B(n16520), .X(n16518) );
  nor_x1_sg U58618 ( .A(n16520), .B(n16519), .X(n16521) );
  nand_x1_sg U58619 ( .A(n17336), .B(n17337), .X(n17335) );
  nor_x1_sg U58620 ( .A(n17337), .B(n17336), .X(n17338) );
  nand_x1_sg U58621 ( .A(n18157), .B(n18158), .X(n18156) );
  nor_x1_sg U58622 ( .A(n18158), .B(n18157), .X(n18159) );
  nand_x1_sg U58623 ( .A(n18978), .B(n18979), .X(n18977) );
  nor_x1_sg U58624 ( .A(n18979), .B(n18978), .X(n18980) );
  nand_x1_sg U58625 ( .A(n7311), .B(n7312), .X(n7310) );
  nor_x1_sg U58626 ( .A(n7312), .B(n7311), .X(n7313) );
  nand_x1_sg U58627 ( .A(n17136), .B(n17137), .X(n17135) );
  nor_x1_sg U58628 ( .A(n17137), .B(n17136), .X(n17138) );
  nand_x1_sg U58629 ( .A(n7021), .B(n7022), .X(n7020) );
  nor_x1_sg U58630 ( .A(n7022), .B(n7021), .X(n7023) );
  nand_x1_sg U58631 ( .A(n7839), .B(n7840), .X(n7838) );
  nor_x1_sg U58632 ( .A(n7840), .B(n7839), .X(n7841) );
  nand_x1_sg U58633 ( .A(n8657), .B(n8658), .X(n8656) );
  nor_x1_sg U58634 ( .A(n8658), .B(n8657), .X(n8659) );
  nand_x1_sg U58635 ( .A(n9477), .B(n9478), .X(n9476) );
  nor_x1_sg U58636 ( .A(n9478), .B(n9477), .X(n9479) );
  nand_x1_sg U58637 ( .A(n10296), .B(n10297), .X(n10295) );
  nor_x1_sg U58638 ( .A(n10297), .B(n10296), .X(n10298) );
  nand_x1_sg U58639 ( .A(n11115), .B(n11116), .X(n11114) );
  nor_x1_sg U58640 ( .A(n11116), .B(n11115), .X(n11117) );
  nand_x1_sg U58641 ( .A(n11934), .B(n11935), .X(n11933) );
  nor_x1_sg U58642 ( .A(n11935), .B(n11934), .X(n11936) );
  nand_x1_sg U58643 ( .A(n12753), .B(n12754), .X(n12752) );
  nor_x1_sg U58644 ( .A(n12754), .B(n12753), .X(n12755) );
  nand_x1_sg U58645 ( .A(n13572), .B(n13573), .X(n13571) );
  nor_x1_sg U58646 ( .A(n13573), .B(n13572), .X(n13574) );
  nand_x1_sg U58647 ( .A(n14391), .B(n14392), .X(n14390) );
  nor_x1_sg U58648 ( .A(n14392), .B(n14391), .X(n14393) );
  nand_x1_sg U58649 ( .A(n15210), .B(n15211), .X(n15209) );
  nor_x1_sg U58650 ( .A(n15211), .B(n15210), .X(n15212) );
  nand_x1_sg U58651 ( .A(n16029), .B(n16030), .X(n16028) );
  nor_x1_sg U58652 ( .A(n16030), .B(n16029), .X(n16031) );
  nand_x1_sg U58653 ( .A(n17667), .B(n17668), .X(n17666) );
  nor_x1_sg U58654 ( .A(n17668), .B(n17667), .X(n17669) );
  nand_x1_sg U58655 ( .A(n18488), .B(n18489), .X(n18487) );
  nor_x1_sg U58656 ( .A(n18489), .B(n18488), .X(n18490) );
  nand_x1_sg U58657 ( .A(n6845), .B(n46861), .X(n6844) );
  nor_x1_sg U58658 ( .A(n46861), .B(n6845), .X(n6846) );
  nand_x1_sg U58659 ( .A(n7662), .B(n47154), .X(n7661) );
  nor_x1_sg U58660 ( .A(n47154), .B(n7662), .X(n7663) );
  nand_x1_sg U58661 ( .A(n8480), .B(n47439), .X(n8479) );
  nor_x1_sg U58662 ( .A(n47439), .B(n8480), .X(n8481) );
  nand_x1_sg U58663 ( .A(n9300), .B(n47724), .X(n9299) );
  nor_x1_sg U58664 ( .A(n47724), .B(n9300), .X(n9301) );
  nand_x1_sg U58665 ( .A(n10119), .B(n48009), .X(n10118) );
  nor_x1_sg U58666 ( .A(n48009), .B(n10119), .X(n10120) );
  nand_x1_sg U58667 ( .A(n10938), .B(n48294), .X(n10937) );
  nor_x1_sg U58668 ( .A(n48294), .B(n10938), .X(n10939) );
  nand_x1_sg U58669 ( .A(n11757), .B(n48579), .X(n11756) );
  nor_x1_sg U58670 ( .A(n48579), .B(n11757), .X(n11758) );
  nand_x1_sg U58671 ( .A(n12576), .B(n48865), .X(n12575) );
  nor_x1_sg U58672 ( .A(n48865), .B(n12576), .X(n12577) );
  nand_x1_sg U58673 ( .A(n13395), .B(n49152), .X(n13394) );
  nor_x1_sg U58674 ( .A(n49152), .B(n13395), .X(n13396) );
  nand_x1_sg U58675 ( .A(n14214), .B(n49438), .X(n14213) );
  nor_x1_sg U58676 ( .A(n49438), .B(n14214), .X(n14215) );
  nand_x1_sg U58677 ( .A(n15033), .B(n49723), .X(n15032) );
  nor_x1_sg U58678 ( .A(n49723), .B(n15033), .X(n15034) );
  nand_x1_sg U58679 ( .A(n15852), .B(n50010), .X(n15851) );
  nor_x1_sg U58680 ( .A(n50010), .B(n15852), .X(n15853) );
  nand_x1_sg U58681 ( .A(n16669), .B(n50294), .X(n16668) );
  nor_x1_sg U58682 ( .A(n50294), .B(n16669), .X(n16670) );
  nand_x1_sg U58683 ( .A(n17490), .B(n50584), .X(n17489) );
  nor_x1_sg U58684 ( .A(n50584), .B(n17490), .X(n17491) );
  nand_x1_sg U58685 ( .A(n18311), .B(n50871), .X(n18310) );
  nor_x1_sg U58686 ( .A(n50871), .B(n18311), .X(n18312) );
  nand_x1_sg U58687 ( .A(n6968), .B(n6969), .X(n6967) );
  nor_x1_sg U58688 ( .A(n6969), .B(n6968), .X(n6970) );
  nand_x1_sg U58689 ( .A(n7785), .B(n7786), .X(n7784) );
  nor_x1_sg U58690 ( .A(n7786), .B(n7785), .X(n7787) );
  nand_x1_sg U58691 ( .A(n8603), .B(n8604), .X(n8602) );
  nor_x1_sg U58692 ( .A(n8604), .B(n8603), .X(n8605) );
  nand_x1_sg U58693 ( .A(n9423), .B(n9424), .X(n9422) );
  nor_x1_sg U58694 ( .A(n9424), .B(n9423), .X(n9425) );
  nand_x1_sg U58695 ( .A(n10242), .B(n10243), .X(n10241) );
  nor_x1_sg U58696 ( .A(n10243), .B(n10242), .X(n10244) );
  nand_x1_sg U58697 ( .A(n11061), .B(n11062), .X(n11060) );
  nor_x1_sg U58698 ( .A(n11062), .B(n11061), .X(n11063) );
  nand_x1_sg U58699 ( .A(n11880), .B(n11881), .X(n11879) );
  nor_x1_sg U58700 ( .A(n11881), .B(n11880), .X(n11882) );
  nand_x1_sg U58701 ( .A(n12699), .B(n12700), .X(n12698) );
  nor_x1_sg U58702 ( .A(n12700), .B(n12699), .X(n12701) );
  nand_x1_sg U58703 ( .A(n13518), .B(n13519), .X(n13517) );
  nor_x1_sg U58704 ( .A(n13519), .B(n13518), .X(n13520) );
  nand_x1_sg U58705 ( .A(n14337), .B(n14338), .X(n14336) );
  nor_x1_sg U58706 ( .A(n14338), .B(n14337), .X(n14339) );
  nand_x1_sg U58707 ( .A(n15156), .B(n15157), .X(n15155) );
  nor_x1_sg U58708 ( .A(n15157), .B(n15156), .X(n15158) );
  nand_x1_sg U58709 ( .A(n15975), .B(n15976), .X(n15974) );
  nor_x1_sg U58710 ( .A(n15976), .B(n15975), .X(n15977) );
  nand_x1_sg U58711 ( .A(n16792), .B(n16793), .X(n16791) );
  nor_x1_sg U58712 ( .A(n16793), .B(n16792), .X(n16794) );
  nand_x1_sg U58713 ( .A(n17613), .B(n17614), .X(n17612) );
  nor_x1_sg U58714 ( .A(n17614), .B(n17613), .X(n17615) );
  nand_x1_sg U58715 ( .A(n18434), .B(n18435), .X(n18433) );
  nor_x1_sg U58716 ( .A(n18435), .B(n18434), .X(n18436) );
  nand_x1_sg U58717 ( .A(n16842), .B(n16843), .X(n16841) );
  nor_x1_sg U58718 ( .A(n16843), .B(n16842), .X(n16844) );
  nand_x1_sg U58719 ( .A(n47076), .B(n6985), .X(n6984) );
  nor_x1_sg U58720 ( .A(n6985), .B(n47076), .X(n6986) );
  nand_x1_sg U58721 ( .A(n47362), .B(n7802), .X(n7801) );
  nor_x1_sg U58722 ( .A(n7802), .B(n47362), .X(n7803) );
  nand_x1_sg U58723 ( .A(n47647), .B(n8620), .X(n8619) );
  nor_x1_sg U58724 ( .A(n8620), .B(n47647), .X(n8621) );
  nand_x1_sg U58725 ( .A(n47932), .B(n9440), .X(n9439) );
  nor_x1_sg U58726 ( .A(n9440), .B(n47932), .X(n9441) );
  nand_x1_sg U58727 ( .A(n48217), .B(n10259), .X(n10258) );
  nor_x1_sg U58728 ( .A(n10259), .B(n48217), .X(n10260) );
  nand_x1_sg U58729 ( .A(n48502), .B(n11078), .X(n11077) );
  nor_x1_sg U58730 ( .A(n11078), .B(n48502), .X(n11079) );
  nand_x1_sg U58731 ( .A(n48787), .B(n11897), .X(n11896) );
  nor_x1_sg U58732 ( .A(n11897), .B(n48787), .X(n11898) );
  nand_x1_sg U58733 ( .A(n49074), .B(n12716), .X(n12715) );
  nor_x1_sg U58734 ( .A(n12716), .B(n49074), .X(n12717) );
  nand_x1_sg U58735 ( .A(n49360), .B(n13535), .X(n13534) );
  nor_x1_sg U58736 ( .A(n13535), .B(n49360), .X(n13536) );
  nand_x1_sg U58737 ( .A(n49646), .B(n14354), .X(n14353) );
  nor_x1_sg U58738 ( .A(n14354), .B(n49646), .X(n14355) );
  nand_x1_sg U58739 ( .A(n49932), .B(n15173), .X(n15172) );
  nor_x1_sg U58740 ( .A(n15173), .B(n49932), .X(n15174) );
  nand_x1_sg U58741 ( .A(n50218), .B(n15992), .X(n15991) );
  nor_x1_sg U58742 ( .A(n15992), .B(n50218), .X(n15993) );
  nand_x1_sg U58743 ( .A(n50503), .B(n16809), .X(n16808) );
  nor_x1_sg U58744 ( .A(n16809), .B(n50503), .X(n16810) );
  nand_x1_sg U58745 ( .A(n50792), .B(n17630), .X(n17629) );
  nor_x1_sg U58746 ( .A(n17630), .B(n50792), .X(n17631) );
  nand_x1_sg U58747 ( .A(n51079), .B(n18451), .X(n18450) );
  nor_x1_sg U58748 ( .A(n18451), .B(n51079), .X(n18452) );
  nand_x1_sg U58749 ( .A(n47297), .B(n7769), .X(n7768) );
  nor_x1_sg U58750 ( .A(n7769), .B(n47297), .X(n7770) );
  nand_x1_sg U58751 ( .A(n47582), .B(n8587), .X(n8586) );
  nor_x1_sg U58752 ( .A(n8587), .B(n47582), .X(n8588) );
  nand_x1_sg U58753 ( .A(n47867), .B(n9407), .X(n9406) );
  nor_x1_sg U58754 ( .A(n9407), .B(n47867), .X(n9408) );
  nand_x1_sg U58755 ( .A(n48152), .B(n10226), .X(n10225) );
  nor_x1_sg U58756 ( .A(n10226), .B(n48152), .X(n10227) );
  nand_x1_sg U58757 ( .A(n48437), .B(n11045), .X(n11044) );
  nor_x1_sg U58758 ( .A(n11045), .B(n48437), .X(n11046) );
  nand_x1_sg U58759 ( .A(n48722), .B(n11864), .X(n11863) );
  nor_x1_sg U58760 ( .A(n11864), .B(n48722), .X(n11865) );
  nand_x1_sg U58761 ( .A(n49008), .B(n12683), .X(n12682) );
  nor_x1_sg U58762 ( .A(n12683), .B(n49008), .X(n12684) );
  nand_x1_sg U58763 ( .A(n49295), .B(n13502), .X(n13501) );
  nor_x1_sg U58764 ( .A(n13502), .B(n49295), .X(n13503) );
  nand_x1_sg U58765 ( .A(n49581), .B(n14321), .X(n14320) );
  nor_x1_sg U58766 ( .A(n14321), .B(n49581), .X(n14322) );
  nand_x1_sg U58767 ( .A(n49867), .B(n15140), .X(n15139) );
  nor_x1_sg U58768 ( .A(n15140), .B(n49867), .X(n15141) );
  nand_x1_sg U58769 ( .A(n50153), .B(n15959), .X(n15958) );
  nor_x1_sg U58770 ( .A(n15959), .B(n50153), .X(n15960) );
  nand_x1_sg U58771 ( .A(n50727), .B(n17597), .X(n17596) );
  nor_x1_sg U58772 ( .A(n17597), .B(n50727), .X(n17598) );
  nand_x1_sg U58773 ( .A(n51014), .B(n18418), .X(n18417) );
  nor_x1_sg U58774 ( .A(n18418), .B(n51014), .X(n18419) );
  nor_x1_sg U58775 ( .A(n38893), .B(n16666), .X(\L2_0/n2552 ) );
  nor_x1_sg U58776 ( .A(n40927), .B(n16685), .X(\L2_0/n2540 ) );
  nor_x1_sg U58777 ( .A(n38893), .B(n16691), .X(\L2_0/n2536 ) );
  nor_x1_sg U58778 ( .A(n40925), .B(n16703), .X(\L2_0/n2528 ) );
  nor_x1_sg U58779 ( .A(n40967), .B(n17487), .X(\L2_0/n2472 ) );
  nor_x1_sg U58780 ( .A(n40965), .B(n17506), .X(\L2_0/n2460 ) );
  nor_x1_sg U58781 ( .A(n40966), .B(n17512), .X(\L2_0/n2456 ) );
  nor_x1_sg U58782 ( .A(n40967), .B(n17524), .X(\L2_0/n2448 ) );
  inv_x1_sg U58783 ( .A(n7600), .X(n46973) );
  inv_x1_sg U58784 ( .A(n8418), .X(n47263) );
  inv_x1_sg U58785 ( .A(n9236), .X(n47548) );
  inv_x1_sg U58786 ( .A(n10056), .X(n47833) );
  inv_x1_sg U58787 ( .A(n10875), .X(n48118) );
  inv_x1_sg U58788 ( .A(n11694), .X(n48403) );
  inv_x1_sg U58789 ( .A(n12513), .X(n48688) );
  inv_x1_sg U58790 ( .A(n13332), .X(n48974) );
  inv_x1_sg U58791 ( .A(n14151), .X(n49261) );
  inv_x1_sg U58792 ( .A(n14970), .X(n49547) );
  inv_x1_sg U58793 ( .A(n15789), .X(n49833) );
  inv_x1_sg U58794 ( .A(n16608), .X(n50119) );
  inv_x1_sg U58795 ( .A(n18246), .X(n50693) );
  inv_x1_sg U58796 ( .A(n19067), .X(n50980) );
  inv_x1_sg U58797 ( .A(n7582), .X(n46991) );
  inv_x1_sg U58798 ( .A(n8400), .X(n47280) );
  inv_x1_sg U58799 ( .A(n9218), .X(n47565) );
  inv_x1_sg U58800 ( .A(n10038), .X(n47850) );
  inv_x1_sg U58801 ( .A(n10857), .X(n48135) );
  inv_x1_sg U58802 ( .A(n11676), .X(n48420) );
  inv_x1_sg U58803 ( .A(n12495), .X(n48705) );
  inv_x1_sg U58804 ( .A(n13314), .X(n48991) );
  inv_x1_sg U58805 ( .A(n14133), .X(n49278) );
  inv_x1_sg U58806 ( .A(n14952), .X(n49564) );
  inv_x1_sg U58807 ( .A(n15771), .X(n49850) );
  inv_x1_sg U58808 ( .A(n16590), .X(n50136) );
  inv_x1_sg U58809 ( .A(n18228), .X(n50710) );
  inv_x1_sg U58810 ( .A(n19049), .X(n50997) );
  inv_x1_sg U58811 ( .A(n17425), .X(n50404) );
  inv_x1_sg U58812 ( .A(n17407), .X(n50421) );
  inv_x1_sg U58813 ( .A(n7357), .X(n47004) );
  inv_x1_sg U58814 ( .A(n8175), .X(n47293) );
  inv_x1_sg U58815 ( .A(n8993), .X(n47578) );
  inv_x1_sg U58816 ( .A(n9813), .X(n47863) );
  inv_x1_sg U58817 ( .A(n10632), .X(n48148) );
  inv_x1_sg U58818 ( .A(n11451), .X(n48433) );
  inv_x1_sg U58819 ( .A(n12270), .X(n48718) );
  inv_x1_sg U58820 ( .A(n13089), .X(n49004) );
  inv_x1_sg U58821 ( .A(n13908), .X(n49291) );
  inv_x1_sg U58822 ( .A(n14727), .X(n49577) );
  inv_x1_sg U58823 ( .A(n15546), .X(n49863) );
  inv_x1_sg U58824 ( .A(n16365), .X(n50149) );
  inv_x1_sg U58825 ( .A(n17182), .X(n50434) );
  inv_x1_sg U58826 ( .A(n18003), .X(n50723) );
  inv_x1_sg U58827 ( .A(n18824), .X(n51010) );
  nor_x1_sg U58828 ( .A(n38892), .B(n6861), .X(\L2_0/n3500 ) );
  nor_x1_sg U58829 ( .A(n40922), .B(n6867), .X(\L2_0/n3496 ) );
  nand_x1_sg U58830 ( .A(n41192), .B(n47141), .X(n22875) );
  nand_x1_sg U58831 ( .A(n41194), .B(n47159), .X(n22889) );
  nand_x1_sg U58832 ( .A(n39222), .B(n22908), .X(n22917) );
  nand_x1_sg U58833 ( .A(n41192), .B(n22922), .X(n22931) );
  nand_x1_sg U58834 ( .A(n41193), .B(n22936), .X(n22945) );
  nand_x1_sg U58835 ( .A(n40506), .B(n22950), .X(n22959) );
  nand_x1_sg U58836 ( .A(n41187), .B(n47426), .X(n23152) );
  nand_x1_sg U58837 ( .A(n41190), .B(n47444), .X(n23166) );
  nand_x1_sg U58838 ( .A(n41189), .B(n23185), .X(n23194) );
  nand_x1_sg U58839 ( .A(n41188), .B(n23199), .X(n23208) );
  nand_x1_sg U58840 ( .A(n41189), .B(n23213), .X(n23222) );
  nand_x1_sg U58841 ( .A(n41190), .B(n23227), .X(n23236) );
  nand_x1_sg U58842 ( .A(n41183), .B(n47711), .X(n23432) );
  nand_x1_sg U58843 ( .A(n41184), .B(n47729), .X(n23446) );
  nand_x1_sg U58844 ( .A(n41182), .B(n23465), .X(n23474) );
  nand_x1_sg U58845 ( .A(n40498), .B(n23479), .X(n23488) );
  nand_x1_sg U58846 ( .A(n41185), .B(n23493), .X(n23502) );
  nand_x1_sg U58847 ( .A(n39226), .B(n23507), .X(n23516) );
  nand_x1_sg U58848 ( .A(n39228), .B(n47996), .X(n23711) );
  nand_x1_sg U58849 ( .A(n41180), .B(n48014), .X(n23725) );
  nand_x1_sg U58850 ( .A(n40494), .B(n23744), .X(n23753) );
  nand_x1_sg U58851 ( .A(n41179), .B(n23758), .X(n23767) );
  nand_x1_sg U58852 ( .A(n41178), .B(n23772), .X(n23781) );
  nand_x1_sg U58853 ( .A(n41180), .B(n23786), .X(n23795) );
  nand_x1_sg U58854 ( .A(n39230), .B(n48281), .X(n23990) );
  nand_x1_sg U58855 ( .A(n41172), .B(n48299), .X(n24004) );
  nand_x1_sg U58856 ( .A(n41174), .B(n24023), .X(n24032) );
  nand_x1_sg U58857 ( .A(n41172), .B(n24037), .X(n24046) );
  nand_x1_sg U58858 ( .A(n41175), .B(n24051), .X(n24060) );
  nand_x1_sg U58859 ( .A(n41173), .B(n24065), .X(n24074) );
  nand_x1_sg U58860 ( .A(n41169), .B(n48566), .X(n24269) );
  nand_x1_sg U58861 ( .A(n41167), .B(n48584), .X(n24283) );
  nand_x1_sg U58862 ( .A(n41168), .B(n24302), .X(n24311) );
  nand_x1_sg U58863 ( .A(n41168), .B(n24316), .X(n24325) );
  nand_x1_sg U58864 ( .A(n39232), .B(n24330), .X(n24339) );
  nand_x1_sg U58865 ( .A(n41167), .B(n24344), .X(n24353) );
  nand_x1_sg U58866 ( .A(n41163), .B(n48851), .X(n24548) );
  nand_x1_sg U58867 ( .A(n41164), .B(n48870), .X(n24562) );
  nand_x1_sg U58868 ( .A(n39234), .B(n24581), .X(n24590) );
  nand_x1_sg U58869 ( .A(n41163), .B(n24595), .X(n24604) );
  nand_x1_sg U58870 ( .A(n41162), .B(n24609), .X(n24618) );
  nand_x1_sg U58871 ( .A(n41162), .B(n24623), .X(n24632) );
  nand_x1_sg U58872 ( .A(n39236), .B(n49138), .X(n24826) );
  nand_x1_sg U58873 ( .A(n41158), .B(n49157), .X(n24840) );
  nand_x1_sg U58874 ( .A(n39236), .B(n24859), .X(n24868) );
  nand_x1_sg U58875 ( .A(n41158), .B(n24873), .X(n24882) );
  nand_x1_sg U58876 ( .A(n41157), .B(n24887), .X(n24896) );
  nand_x1_sg U58877 ( .A(n41159), .B(n24901), .X(n24910) );
  nand_x1_sg U58878 ( .A(n41154), .B(n49424), .X(n25105) );
  nand_x1_sg U58879 ( .A(n41152), .B(n49443), .X(n25119) );
  nand_x1_sg U58880 ( .A(n41155), .B(n25138), .X(n25147) );
  nand_x1_sg U58881 ( .A(n41152), .B(n25152), .X(n25161) );
  nand_x1_sg U58882 ( .A(n41154), .B(n25166), .X(n25175) );
  nand_x1_sg U58883 ( .A(n41153), .B(n25180), .X(n25189) );
  nand_x1_sg U58884 ( .A(n41148), .B(n49710), .X(n25384) );
  nand_x1_sg U58885 ( .A(n41149), .B(n49728), .X(n25398) );
  nand_x1_sg U58886 ( .A(n39240), .B(n25417), .X(n25426) );
  nand_x1_sg U58887 ( .A(n41149), .B(n25431), .X(n25440) );
  nand_x1_sg U58888 ( .A(n41148), .B(n25445), .X(n25454) );
  nand_x1_sg U58889 ( .A(n40470), .B(n25459), .X(n25468) );
  nand_x1_sg U58890 ( .A(n41144), .B(n49996), .X(n25663) );
  nand_x1_sg U58891 ( .A(n40466), .B(n50015), .X(n25677) );
  nand_x1_sg U58892 ( .A(n41142), .B(n25696), .X(n25705) );
  nand_x1_sg U58893 ( .A(n41143), .B(n25710), .X(n25719) );
  nand_x1_sg U58894 ( .A(n39242), .B(n25724), .X(n25733) );
  nand_x1_sg U58895 ( .A(n39242), .B(n25738), .X(n25747) );
  nand_x1_sg U58896 ( .A(n41138), .B(n50571), .X(n26206) );
  nand_x1_sg U58897 ( .A(n41139), .B(n50589), .X(n26222) );
  nand_x1_sg U58898 ( .A(n41140), .B(n26244), .X(n26254) );
  nand_x1_sg U58899 ( .A(n40462), .B(n26260), .X(n26270) );
  nand_x1_sg U58900 ( .A(n41140), .B(n26276), .X(n26286) );
  nand_x1_sg U58901 ( .A(n41138), .B(n26292), .X(n26302) );
  nand_x1_sg U58902 ( .A(n41134), .B(n50857), .X(n26500) );
  nand_x1_sg U58903 ( .A(n41135), .B(n50876), .X(n26514) );
  nand_x1_sg U58904 ( .A(n41132), .B(n26533), .X(n26542) );
  nand_x1_sg U58905 ( .A(n41133), .B(n26547), .X(n26556) );
  nand_x1_sg U58906 ( .A(n41135), .B(n26561), .X(n26570) );
  nand_x1_sg U58907 ( .A(n41132), .B(n26575), .X(n26584) );
  nand_x1_sg U58908 ( .A(n39347), .B(n41604), .X(n7140) );
  nand_x1_sg U58909 ( .A(n39345), .B(n41605), .X(n7958) );
  nand_x1_sg U58910 ( .A(n39343), .B(n41606), .X(n8776) );
  nand_x1_sg U58911 ( .A(n39341), .B(n41607), .X(n9596) );
  nand_x1_sg U58912 ( .A(n39339), .B(n41608), .X(n10415) );
  nand_x1_sg U58913 ( .A(n39337), .B(n41609), .X(n11234) );
  nand_x1_sg U58914 ( .A(n39335), .B(n41610), .X(n12053) );
  nand_x1_sg U58915 ( .A(n39333), .B(n41611), .X(n12872) );
  nand_x1_sg U58916 ( .A(n39331), .B(n41612), .X(n13691) );
  nand_x1_sg U58917 ( .A(n39329), .B(n41613), .X(n14510) );
  nand_x1_sg U58918 ( .A(n39327), .B(n41614), .X(n15329) );
  nand_x1_sg U58919 ( .A(n39325), .B(n41615), .X(n16148) );
  nand_x1_sg U58920 ( .A(n39323), .B(n41616), .X(n17786) );
  nand_x1_sg U58921 ( .A(n39321), .B(n41617), .X(n18607) );
  inv_x1_sg U58922 ( .A(n7330), .X(n46993) );
  inv_x1_sg U58923 ( .A(n8148), .X(n47282) );
  inv_x1_sg U58924 ( .A(n8966), .X(n47567) );
  inv_x1_sg U58925 ( .A(n9786), .X(n47852) );
  inv_x1_sg U58926 ( .A(n10605), .X(n48137) );
  inv_x1_sg U58927 ( .A(n11424), .X(n48422) );
  inv_x1_sg U58928 ( .A(n12243), .X(n48707) );
  inv_x1_sg U58929 ( .A(n13062), .X(n48993) );
  inv_x1_sg U58930 ( .A(n13881), .X(n49280) );
  inv_x1_sg U58931 ( .A(n14700), .X(n49566) );
  inv_x1_sg U58932 ( .A(n15519), .X(n49852) );
  inv_x1_sg U58933 ( .A(n16338), .X(n50138) );
  inv_x1_sg U58934 ( .A(n17155), .X(n50423) );
  inv_x1_sg U58935 ( .A(n17976), .X(n50712) );
  inv_x1_sg U58936 ( .A(n18797), .X(n50999) );
  inv_x1_sg U58937 ( .A(n7423), .X(n47018) );
  inv_x1_sg U58938 ( .A(n8241), .X(n47306) );
  inv_x1_sg U58939 ( .A(n9059), .X(n47591) );
  inv_x1_sg U58940 ( .A(n9879), .X(n47876) );
  inv_x1_sg U58941 ( .A(n10698), .X(n48161) );
  inv_x1_sg U58942 ( .A(n11517), .X(n48446) );
  inv_x1_sg U58943 ( .A(n12336), .X(n48731) );
  inv_x1_sg U58944 ( .A(n13155), .X(n49017) );
  inv_x1_sg U58945 ( .A(n13974), .X(n49304) );
  inv_x1_sg U58946 ( .A(n14793), .X(n49590) );
  inv_x1_sg U58947 ( .A(n15612), .X(n49876) );
  inv_x1_sg U58948 ( .A(n16431), .X(n50162) );
  inv_x1_sg U58949 ( .A(n17248), .X(n50447) );
  inv_x1_sg U58950 ( .A(n18069), .X(n50736) );
  inv_x1_sg U58951 ( .A(n18890), .X(n51023) );
  inv_x1_sg U58952 ( .A(n7465), .X(n46956) );
  inv_x1_sg U58953 ( .A(n8283), .X(n47247) );
  inv_x1_sg U58954 ( .A(n9101), .X(n47532) );
  inv_x1_sg U58955 ( .A(n9921), .X(n47817) );
  inv_x1_sg U58956 ( .A(n10740), .X(n48102) );
  inv_x1_sg U58957 ( .A(n11559), .X(n48387) );
  inv_x1_sg U58958 ( .A(n12378), .X(n48672) );
  inv_x1_sg U58959 ( .A(n13197), .X(n48958) );
  inv_x1_sg U58960 ( .A(n14016), .X(n49245) );
  inv_x1_sg U58961 ( .A(n14835), .X(n49531) );
  inv_x1_sg U58962 ( .A(n15654), .X(n49817) );
  inv_x1_sg U58963 ( .A(n16473), .X(n50103) );
  inv_x1_sg U58964 ( .A(n18111), .X(n50677) );
  inv_x1_sg U58965 ( .A(n18932), .X(n50964) );
  inv_x1_sg U58966 ( .A(n7389), .X(n46971) );
  inv_x1_sg U58967 ( .A(n17214), .X(n50402) );
  nand_x1_sg U58968 ( .A(n39660), .B(n46849), .X(n22612) );
  nand_x1_sg U58969 ( .A(n41306), .B(n46853), .X(n22618) );
  nand_x1_sg U58970 ( .A(n41948), .B(n46866), .X(n22624) );
  nand_x1_sg U58971 ( .A(n39660), .B(n46876), .X(n22630) );
  nand_x1_sg U58972 ( .A(n39659), .B(n46914), .X(n22649) );
  inv_x1_sg U58973 ( .A(n22642), .X(n46914) );
  nand_x1_sg U58974 ( .A(n41948), .B(n46963), .X(n22662) );
  nand_x1_sg U58975 ( .A(n41305), .B(n46982), .X(n22668) );
  nand_x1_sg U58976 ( .A(n39137), .B(n47005), .X(n22674) );
  nand_x1_sg U58977 ( .A(n39137), .B(n47024), .X(n22680) );
  nand_x1_sg U58978 ( .A(n41307), .B(n47054), .X(n22686) );
  nand_x1_sg U58979 ( .A(n41304), .B(n22697), .X(n22703) );
  nand_x1_sg U58980 ( .A(n6958), .B(n41599), .X(n6955) );
  nand_x1_sg U58981 ( .A(n16782), .B(n41598), .X(n16779) );
  nand_x1_sg U58982 ( .A(n7775), .B(n41602), .X(n7772) );
  nand_x1_sg U58983 ( .A(n8593), .B(n41597), .X(n8590) );
  nand_x1_sg U58984 ( .A(n9413), .B(n41596), .X(n9410) );
  nand_x1_sg U58985 ( .A(n10232), .B(n41595), .X(n10229) );
  nand_x1_sg U58986 ( .A(n11051), .B(n41594), .X(n11048) );
  nand_x1_sg U58987 ( .A(n11870), .B(n41593), .X(n11867) );
  nand_x1_sg U58988 ( .A(n12689), .B(n41592), .X(n12686) );
  nand_x1_sg U58989 ( .A(n13508), .B(n41591), .X(n13505) );
  nand_x1_sg U58990 ( .A(n14327), .B(n41590), .X(n14324) );
  nand_x1_sg U58991 ( .A(n15146), .B(n41601), .X(n15143) );
  nand_x1_sg U58992 ( .A(n15965), .B(n41589), .X(n15962) );
  nand_x1_sg U58993 ( .A(n17603), .B(n41600), .X(n17600) );
  nand_x1_sg U58994 ( .A(n18424), .B(n41588), .X(n18421) );
  inv_x1_sg U58995 ( .A(n7593), .X(n47045) );
  inv_x1_sg U58996 ( .A(n17418), .X(n50473) );
  inv_x1_sg U58997 ( .A(n7397), .X(n46958) );
  inv_x1_sg U58998 ( .A(n8215), .X(n47249) );
  inv_x1_sg U58999 ( .A(n9033), .X(n47534) );
  inv_x1_sg U59000 ( .A(n9853), .X(n47819) );
  inv_x1_sg U59001 ( .A(n10672), .X(n48104) );
  inv_x1_sg U59002 ( .A(n11491), .X(n48389) );
  inv_x1_sg U59003 ( .A(n12310), .X(n48674) );
  inv_x1_sg U59004 ( .A(n13129), .X(n48960) );
  inv_x1_sg U59005 ( .A(n13948), .X(n49247) );
  inv_x1_sg U59006 ( .A(n14767), .X(n49533) );
  inv_x1_sg U59007 ( .A(n15586), .X(n49819) );
  inv_x1_sg U59008 ( .A(n16405), .X(n50105) );
  inv_x1_sg U59009 ( .A(n18043), .X(n50679) );
  inv_x1_sg U59010 ( .A(n18864), .X(n50966) );
  inv_x1_sg U59011 ( .A(n7377), .X(n46939) );
  inv_x1_sg U59012 ( .A(n8195), .X(n47230) );
  inv_x1_sg U59013 ( .A(n9013), .X(n47515) );
  inv_x1_sg U59014 ( .A(n9833), .X(n47800) );
  inv_x1_sg U59015 ( .A(n10652), .X(n48085) );
  inv_x1_sg U59016 ( .A(n11471), .X(n48370) );
  inv_x1_sg U59017 ( .A(n12290), .X(n48655) );
  inv_x1_sg U59018 ( .A(n13109), .X(n48941) );
  inv_x1_sg U59019 ( .A(n13928), .X(n49228) );
  inv_x1_sg U59020 ( .A(n14747), .X(n49514) );
  inv_x1_sg U59021 ( .A(n15566), .X(n49800) );
  inv_x1_sg U59022 ( .A(n16385), .X(n50086) );
  inv_x1_sg U59023 ( .A(n18023), .X(n50660) );
  inv_x1_sg U59024 ( .A(n18844), .X(n50947) );
  inv_x1_sg U59025 ( .A(n8411), .X(n47332) );
  inv_x1_sg U59026 ( .A(n9229), .X(n47617) );
  inv_x1_sg U59027 ( .A(n10049), .X(n47902) );
  inv_x1_sg U59028 ( .A(n10868), .X(n48187) );
  inv_x1_sg U59029 ( .A(n11687), .X(n48472) );
  inv_x1_sg U59030 ( .A(n12506), .X(n48757) );
  inv_x1_sg U59031 ( .A(n13325), .X(n49043) );
  inv_x1_sg U59032 ( .A(n14144), .X(n49330) );
  inv_x1_sg U59033 ( .A(n14963), .X(n49616) );
  inv_x1_sg U59034 ( .A(n15782), .X(n49902) );
  inv_x1_sg U59035 ( .A(n16601), .X(n50188) );
  inv_x1_sg U59036 ( .A(n18239), .X(n50762) );
  inv_x1_sg U59037 ( .A(n19060), .X(n51049) );
  inv_x1_sg U59038 ( .A(n17222), .X(n50390) );
  inv_x1_sg U59039 ( .A(n8427), .X(n47319) );
  inv_x1_sg U59040 ( .A(n9245), .X(n47604) );
  inv_x1_sg U59041 ( .A(n10065), .X(n47889) );
  inv_x1_sg U59042 ( .A(n10884), .X(n48174) );
  inv_x1_sg U59043 ( .A(n11703), .X(n48459) );
  inv_x1_sg U59044 ( .A(n12522), .X(n48744) );
  inv_x1_sg U59045 ( .A(n13341), .X(n49030) );
  inv_x1_sg U59046 ( .A(n14160), .X(n49317) );
  inv_x1_sg U59047 ( .A(n14979), .X(n49603) );
  inv_x1_sg U59048 ( .A(n15798), .X(n49889) );
  inv_x1_sg U59049 ( .A(n16617), .X(n50175) );
  inv_x1_sg U59050 ( .A(n18255), .X(n50749) );
  inv_x1_sg U59051 ( .A(n19076), .X(n51036) );
  inv_x1_sg U59052 ( .A(n7609), .X(n47032) );
  inv_x1_sg U59053 ( .A(n17434), .X(n50460) );
  inv_x1_sg U59054 ( .A(n17202), .X(n50371) );
  nor_x1_sg U59055 ( .A(n40984), .B(n5734), .X(\L1_0/n3464 ) );
  nor_x1_sg U59056 ( .A(n40985), .B(n5738), .X(\L1_0/n3460 ) );
  nor_x1_sg U59057 ( .A(n40982), .B(n5736), .X(\L1_0/n3452 ) );
  nor_x1_sg U59058 ( .A(n40984), .B(n5739), .X(n5131) );
  nor_x1_sg U59059 ( .A(n40985), .B(n5741), .X(\L1_0/n3440 ) );
  nor_x1_sg U59060 ( .A(n40982), .B(n5768), .X(\L1_0/n3432 ) );
  nor_x1_sg U59061 ( .A(n40983), .B(n5754), .X(n5127) );
  nor_x1_sg U59062 ( .A(n40985), .B(n5757), .X(\L1_0/n3424 ) );
  nor_x1_sg U59063 ( .A(n40983), .B(n5742), .X(n5130) );
  nor_x1_sg U59064 ( .A(n38939), .B(n5751), .X(\L1_0/n3416 ) );
  nor_x1_sg U59065 ( .A(n41944), .B(n5764), .X(\L1_0/n3412 ) );
  nor_x1_sg U59066 ( .A(n40983), .B(n5766), .X(\L1_0/n3404 ) );
  nand_x1_sg U59067 ( .A(n39481), .B(n50282), .X(n25935) );
  nand_x1_sg U59068 ( .A(n41296), .B(n50289), .X(n25941) );
  nand_x1_sg U59069 ( .A(n41296), .B(n50299), .X(n25947) );
  nand_x1_sg U59070 ( .A(n41295), .B(n50302), .X(n25953) );
  nand_x1_sg U59071 ( .A(n39481), .B(n25965), .X(n25973) );
  nand_x1_sg U59072 ( .A(n41297), .B(n25978), .X(n25986) );
  nand_x1_sg U59073 ( .A(n41297), .B(n25990), .X(n25999) );
  nand_x1_sg U59074 ( .A(n41947), .B(n26003), .X(n26012) );
  nand_x1_sg U59075 ( .A(n41295), .B(n42147), .X(n26028) );
  inv_x1_sg U59076 ( .A(n7477), .X(n47065) );
  inv_x1_sg U59077 ( .A(n8295), .X(n47351) );
  inv_x1_sg U59078 ( .A(n9113), .X(n47636) );
  inv_x1_sg U59079 ( .A(n9933), .X(n47921) );
  inv_x1_sg U59080 ( .A(n10752), .X(n48206) );
  inv_x1_sg U59081 ( .A(n11571), .X(n48491) );
  inv_x1_sg U59082 ( .A(n12390), .X(n48776) );
  inv_x1_sg U59083 ( .A(n13209), .X(n49063) );
  inv_x1_sg U59084 ( .A(n14028), .X(n49349) );
  inv_x1_sg U59085 ( .A(n14847), .X(n49635) );
  inv_x1_sg U59086 ( .A(n15666), .X(n49921) );
  inv_x1_sg U59087 ( .A(n16485), .X(n50207) );
  inv_x1_sg U59088 ( .A(n17302), .X(n50492) );
  inv_x1_sg U59089 ( .A(n18123), .X(n50781) );
  inv_x1_sg U59090 ( .A(n18944), .X(n51068) );
  nor_x1_sg U59091 ( .A(n22898), .B(n41387), .X(\L1_0/n4327 ) );
  nor_x1_sg U59092 ( .A(n22919), .B(n39900), .X(\L1_0/n4315 ) );
  nor_x1_sg U59093 ( .A(n22933), .B(n39142), .X(\L1_0/n4307 ) );
  nor_x1_sg U59094 ( .A(n22947), .B(n39143), .X(\L1_0/n4299 ) );
  nor_x1_sg U59095 ( .A(n22973), .B(n41385), .X(\L1_0/n4283 ) );
  nor_x1_sg U59096 ( .A(n40030), .B(n22884), .X(\L1_0/n4336 ) );
  nor_x1_sg U59097 ( .A(n8470), .B(n40843), .X(\L2_0/n3356 ) );
  nor_x1_sg U59098 ( .A(n16659), .B(n38893), .X(\L2_0/n2556 ) );
  nor_x1_sg U59099 ( .A(n17480), .B(n40967), .X(\L2_0/n2476 ) );
  nor_x1_sg U59100 ( .A(n8562), .B(n40844), .X(\L2_0/n3296 ) );
  nor_x1_sg U59101 ( .A(n16751), .B(n16646), .X(\L2_0/n2496 ) );
  nor_x1_sg U59102 ( .A(n17572), .B(n40966), .X(\L2_0/n2416 ) );
  inv_x1_sg U59103 ( .A(n8029), .X(n47208) );
  inv_x1_sg U59104 ( .A(n8847), .X(n47493) );
  inv_x1_sg U59105 ( .A(n9667), .X(n47778) );
  inv_x1_sg U59106 ( .A(n10486), .X(n48063) );
  inv_x1_sg U59107 ( .A(n11305), .X(n48348) );
  inv_x1_sg U59108 ( .A(n12124), .X(n48633) );
  inv_x1_sg U59109 ( .A(n12943), .X(n48919) );
  inv_x1_sg U59110 ( .A(n13762), .X(n49206) );
  inv_x1_sg U59111 ( .A(n14581), .X(n49492) );
  inv_x1_sg U59112 ( .A(n15400), .X(n49778) );
  inv_x1_sg U59113 ( .A(n16219), .X(n50064) );
  inv_x1_sg U59114 ( .A(n17035), .X(n50349) );
  inv_x1_sg U59115 ( .A(n17857), .X(n50638) );
  inv_x1_sg U59116 ( .A(n18678), .X(n50925) );
  nor_x1_sg U59117 ( .A(n8484), .B(n40844), .X(\L2_0/n3348 ) );
  nor_x1_sg U59118 ( .A(n8490), .B(n38861), .X(\L2_0/n3344 ) );
  nor_x1_sg U59119 ( .A(n8508), .B(n8456), .X(\L2_0/n3332 ) );
  nor_x1_sg U59120 ( .A(n8520), .B(n40842), .X(\L2_0/n3324 ) );
  nor_x1_sg U59121 ( .A(n8526), .B(n38861), .X(\L2_0/n3320 ) );
  nor_x1_sg U59122 ( .A(n8532), .B(n8456), .X(\L2_0/n3316 ) );
  nor_x1_sg U59123 ( .A(n8538), .B(n40843), .X(\L2_0/n3312 ) );
  nor_x1_sg U59124 ( .A(n8544), .B(n38861), .X(\L2_0/n3308 ) );
  nor_x1_sg U59125 ( .A(n8550), .B(n40843), .X(\L2_0/n3304 ) );
  nor_x1_sg U59126 ( .A(n8556), .B(n40842), .X(\L2_0/n3300 ) );
  nor_x1_sg U59127 ( .A(n16673), .B(n40926), .X(\L2_0/n2548 ) );
  nor_x1_sg U59128 ( .A(n16679), .B(n40925), .X(\L2_0/n2544 ) );
  nor_x1_sg U59129 ( .A(n16697), .B(n40925), .X(\L2_0/n2532 ) );
  nor_x1_sg U59130 ( .A(n16709), .B(n40926), .X(\L2_0/n2524 ) );
  nor_x1_sg U59131 ( .A(n16715), .B(n40926), .X(\L2_0/n2520 ) );
  nor_x1_sg U59132 ( .A(n16721), .B(n40925), .X(\L2_0/n2516 ) );
  nor_x1_sg U59133 ( .A(n16727), .B(n40926), .X(\L2_0/n2512 ) );
  nor_x1_sg U59134 ( .A(n16733), .B(n16646), .X(\L2_0/n2508 ) );
  nor_x1_sg U59135 ( .A(n16739), .B(n16646), .X(\L2_0/n2504 ) );
  nor_x1_sg U59136 ( .A(n16745), .B(n38893), .X(\L2_0/n2500 ) );
  nor_x1_sg U59137 ( .A(n17494), .B(n17466), .X(\L2_0/n2468 ) );
  nor_x1_sg U59138 ( .A(n17500), .B(n38903), .X(\L2_0/n2464 ) );
  nor_x1_sg U59139 ( .A(n17518), .B(n40965), .X(\L2_0/n2452 ) );
  nor_x1_sg U59140 ( .A(n17530), .B(n40966), .X(\L2_0/n2444 ) );
  nor_x1_sg U59141 ( .A(n17536), .B(n38903), .X(\L2_0/n2440 ) );
  nor_x1_sg U59142 ( .A(n17542), .B(n38903), .X(\L2_0/n2436 ) );
  nor_x1_sg U59143 ( .A(n17548), .B(n17466), .X(\L2_0/n2432 ) );
  nor_x1_sg U59144 ( .A(n17554), .B(n40967), .X(\L2_0/n2428 ) );
  nor_x1_sg U59145 ( .A(n17560), .B(n40965), .X(\L2_0/n2424 ) );
  nor_x1_sg U59146 ( .A(n17566), .B(n40965), .X(\L2_0/n2420 ) );
  nor_x1_sg U59147 ( .A(n41385), .B(n51326), .X(\L1_0/n4316 ) );
  inv_x1_sg U59148 ( .A(n22919), .X(n51326) );
  nor_x1_sg U59149 ( .A(n39142), .B(n51328), .X(\L1_0/n4300 ) );
  inv_x1_sg U59150 ( .A(n22947), .X(n51328) );
  nor_x1_sg U59151 ( .A(n39143), .B(n22961), .X(\L1_0/n4292 ) );
  nor_x1_sg U59152 ( .A(n39900), .B(n22966), .X(\L1_0/n4288 ) );
  nor_x1_sg U59153 ( .A(n40031), .B(n22863), .X(\L1_0/n4348 ) );
  nor_x1_sg U59154 ( .A(n41388), .B(n22877), .X(\L1_0/n4340 ) );
  nor_x1_sg U59155 ( .A(n41386), .B(n51331), .X(\L1_0/n4284 ) );
  inv_x1_sg U59156 ( .A(n22973), .X(n51331) );
  nand_x1_sg U59157 ( .A(n40912), .B(n6836), .X(\L2_0/n3515 ) );
  nand_x1_sg U59158 ( .A(n6835), .B(n39145), .X(n6836) );
  nand_x1_sg U59159 ( .A(n40912), .B(n6843), .X(\L2_0/n3511 ) );
  nand_x1_sg U59160 ( .A(n6842), .B(n41392), .X(n6843) );
  nand_x1_sg U59161 ( .A(n40913), .B(n6850), .X(\L2_0/n3507 ) );
  nand_x1_sg U59162 ( .A(n6849), .B(n40027), .X(n6850) );
  nand_x1_sg U59163 ( .A(n40911), .B(n6856), .X(\L2_0/n3503 ) );
  nand_x1_sg U59164 ( .A(n6855), .B(n39145), .X(n6856) );
  nand_x1_sg U59165 ( .A(n40913), .B(n6862), .X(\L2_0/n3499 ) );
  nand_x1_sg U59166 ( .A(n6861), .B(n40022), .X(n6862) );
  nand_x1_sg U59167 ( .A(n40911), .B(n6868), .X(\L2_0/n3495 ) );
  nand_x1_sg U59168 ( .A(n6867), .B(n40025), .X(n6868) );
  nand_x1_sg U59169 ( .A(n40912), .B(n6874), .X(\L2_0/n3491 ) );
  nand_x1_sg U59170 ( .A(n6873), .B(n40023), .X(n6874) );
  nand_x1_sg U59171 ( .A(n40912), .B(n6880), .X(\L2_0/n3487 ) );
  nand_x1_sg U59172 ( .A(n6879), .B(n40023), .X(n6880) );
  nand_x1_sg U59173 ( .A(n38889), .B(n6886), .X(\L2_0/n3483 ) );
  nand_x1_sg U59174 ( .A(n6885), .B(n41390), .X(n6886) );
  nand_x1_sg U59175 ( .A(n40914), .B(n6892), .X(\L2_0/n3479 ) );
  nand_x1_sg U59176 ( .A(n6891), .B(n40022), .X(n6892) );
  nand_x1_sg U59177 ( .A(n40914), .B(n6898), .X(\L2_0/n3475 ) );
  nand_x1_sg U59178 ( .A(n6897), .B(n39146), .X(n6898) );
  nand_x1_sg U59179 ( .A(n38889), .B(n6904), .X(\L2_0/n3471 ) );
  nand_x1_sg U59180 ( .A(n6903), .B(n39146), .X(n6904) );
  nand_x1_sg U59181 ( .A(n40911), .B(n6910), .X(\L2_0/n3467 ) );
  nand_x1_sg U59182 ( .A(n6909), .B(n41393), .X(n6910) );
  nand_x1_sg U59183 ( .A(n40914), .B(n6916), .X(\L2_0/n3463 ) );
  nand_x1_sg U59184 ( .A(n6915), .B(n41393), .X(n6916) );
  nand_x1_sg U59185 ( .A(n40914), .B(n6922), .X(\L2_0/n3459 ) );
  nand_x1_sg U59186 ( .A(n6921), .B(n40026), .X(n6922) );
  nand_x1_sg U59187 ( .A(n40913), .B(n6928), .X(\L2_0/n3455 ) );
  nand_x1_sg U59188 ( .A(n6927), .B(n40025), .X(n6928) );
  nor_x1_sg U59189 ( .A(n41386), .B(n22891), .X(\L1_0/n4332 ) );
  nor_x1_sg U59190 ( .A(n51203), .B(n41387), .X(\L1_0/n4347 ) );
  inv_x1_sg U59191 ( .A(n22863), .X(n51203) );
  nor_x1_sg U59192 ( .A(n51205), .B(n42000), .X(\L1_0/n4339 ) );
  inv_x1_sg U59193 ( .A(n22877), .X(n51205) );
  nor_x1_sg U59194 ( .A(n51329), .B(n41388), .X(\L1_0/n4291 ) );
  inv_x1_sg U59195 ( .A(n22961), .X(n51329) );
  nor_x1_sg U59196 ( .A(n51330), .B(n40029), .X(\L1_0/n4287 ) );
  inv_x1_sg U59197 ( .A(n22966), .X(n51330) );
  nor_x1_sg U59198 ( .A(n40842), .B(n8477), .X(\L2_0/n3352 ) );
  nor_x1_sg U59199 ( .A(n8456), .B(n8496), .X(\L2_0/n3340 ) );
  nor_x1_sg U59200 ( .A(n38861), .B(n8502), .X(\L2_0/n3336 ) );
  nor_x1_sg U59201 ( .A(n40844), .B(n8514), .X(\L2_0/n3328 ) );
  inv_x1_sg U59202 ( .A(n6950), .X(n47079) );
  inv_x1_sg U59203 ( .A(n7767), .X(n47365) );
  inv_x1_sg U59204 ( .A(n8585), .X(n47650) );
  inv_x1_sg U59205 ( .A(n9405), .X(n47935) );
  inv_x1_sg U59206 ( .A(n10224), .X(n48220) );
  inv_x1_sg U59207 ( .A(n11043), .X(n48505) );
  inv_x1_sg U59208 ( .A(n11862), .X(n48790) );
  inv_x1_sg U59209 ( .A(n12681), .X(n49077) );
  inv_x1_sg U59210 ( .A(n13500), .X(n49363) );
  inv_x1_sg U59211 ( .A(n14319), .X(n49649) );
  inv_x1_sg U59212 ( .A(n15138), .X(n49935) );
  inv_x1_sg U59213 ( .A(n15957), .X(n50221) );
  inv_x1_sg U59214 ( .A(n17595), .X(n50795) );
  inv_x1_sg U59215 ( .A(n18416), .X(n51082) );
  inv_x1_sg U59216 ( .A(n16774), .X(n50506) );
  nor_x1_sg U59217 ( .A(n51206), .B(n41387), .X(\L1_0/n4335 ) );
  inv_x1_sg U59218 ( .A(n22884), .X(n51206) );
  nor_x1_sg U59219 ( .A(n41385), .B(n51324), .X(\L1_0/n4328 ) );
  inv_x1_sg U59220 ( .A(n22898), .X(n51324) );
  nor_x1_sg U59221 ( .A(n41386), .B(n51327), .X(\L1_0/n4308 ) );
  inv_x1_sg U59222 ( .A(n22933), .X(n51327) );
  nor_x1_sg U59223 ( .A(n51207), .B(n40031), .X(\L1_0/n4331 ) );
  inv_x1_sg U59224 ( .A(n22891), .X(n51207) );
  inv_x1_sg U59225 ( .A(n6939), .X(n47101) );
  inv_x1_sg U59226 ( .A(n7756), .X(n47387) );
  inv_x1_sg U59227 ( .A(n8574), .X(n47672) );
  inv_x1_sg U59228 ( .A(n9394), .X(n47957) );
  inv_x1_sg U59229 ( .A(n10213), .X(n48242) );
  inv_x1_sg U59230 ( .A(n11032), .X(n48527) );
  inv_x1_sg U59231 ( .A(n11851), .X(n48812) );
  inv_x1_sg U59232 ( .A(n12670), .X(n49099) );
  inv_x1_sg U59233 ( .A(n13489), .X(n49385) );
  inv_x1_sg U59234 ( .A(n14308), .X(n49671) );
  inv_x1_sg U59235 ( .A(n15127), .X(n49957) );
  inv_x1_sg U59236 ( .A(n15946), .X(n50243) );
  inv_x1_sg U59237 ( .A(n16763), .X(n50528) );
  inv_x1_sg U59238 ( .A(n17584), .X(n50817) );
  inv_x1_sg U59239 ( .A(n18405), .X(n51104) );
  inv_x1_sg U59240 ( .A(n5945), .X(n51199) );
  nand_x1_sg U59241 ( .A(n40022), .B(n19106), .X(n19107) );
  nand_x1_sg U59242 ( .A(n41392), .B(n5952), .X(n5953) );
  nand_x1_sg U59243 ( .A(n40022), .B(n6150), .X(n6151) );
  nand_x1_sg U59244 ( .A(n41392), .B(n6243), .X(n6244) );
  nand_x1_sg U59245 ( .A(n40027), .B(n6332), .X(n6333) );
  nand_x1_sg U59246 ( .A(n40027), .B(n6421), .X(n6422) );
  nand_x1_sg U59247 ( .A(n39145), .B(n6510), .X(n6511) );
  nand_x1_sg U59248 ( .A(n41391), .B(n6599), .X(n6600) );
  nand_x1_sg U59249 ( .A(n41392), .B(n6692), .X(n6693) );
  nand_x1_sg U59250 ( .A(n40025), .B(n6008), .X(n6009) );
  nand_x1_sg U59251 ( .A(n41393), .B(n6105), .X(n6106) );
  nand_x1_sg U59252 ( .A(n41391), .B(n6196), .X(n6197) );
  nand_x1_sg U59253 ( .A(n39146), .B(n6288), .X(n6289) );
  nand_x1_sg U59254 ( .A(n40026), .B(n6377), .X(n6378) );
  nand_x1_sg U59255 ( .A(n41390), .B(n6466), .X(n6467) );
  nand_x1_sg U59256 ( .A(n41391), .B(n6555), .X(n6556) );
  nand_x1_sg U59257 ( .A(n39145), .B(n6644), .X(n6645) );
  nand_x1_sg U59258 ( .A(n41391), .B(n6732), .X(n6733) );
  nor_x1_sg U59259 ( .A(n39722), .B(n40232), .X(n7141) );
  nor_x1_sg U59260 ( .A(n41782), .B(n40180), .X(n7959) );
  nor_x1_sg U59261 ( .A(n41784), .B(n40212), .X(n8777) );
  nor_x1_sg U59262 ( .A(n41786), .B(n40206), .X(n9597) );
  nor_x1_sg U59263 ( .A(n41788), .B(n40204), .X(n10416) );
  nor_x1_sg U59264 ( .A(n39708), .B(n40198), .X(n11235) );
  nor_x1_sg U59265 ( .A(n39704), .B(n40194), .X(n12054) );
  nor_x1_sg U59266 ( .A(n41794), .B(n40190), .X(n12873) );
  nor_x1_sg U59267 ( .A(n39698), .B(n40174), .X(n13692) );
  nor_x1_sg U59268 ( .A(n41798), .B(n40186), .X(n14511) );
  nor_x1_sg U59269 ( .A(n41800), .B(n40170), .X(n15330) );
  nor_x1_sg U59270 ( .A(n41802), .B(n40167), .X(n16149) );
  nor_x1_sg U59271 ( .A(n39687), .B(n40214), .X(n17787) );
  nor_x1_sg U59272 ( .A(n41806), .B(n40182), .X(n18608) );
  nor_x1_sg U59273 ( .A(n39680), .B(n40088), .X(n16929) );
  nand_x1_sg U59274 ( .A(n41118), .B(n40583), .X(n17467) );
  nor_x1_sg U59275 ( .A(n22635), .B(n39851), .X(n22642) );
  nor_x1_sg U59276 ( .A(n39680), .B(n40301), .X(n16927) );
  nor_x1_sg U59277 ( .A(n26003), .B(n16821), .X(n26010) );
  nor_x1_sg U59278 ( .A(n8034), .B(n8033), .X(n8031) );
  nand_x1_sg U59279 ( .A(n8033), .B(n8034), .X(n8032) );
  nor_x1_sg U59280 ( .A(n8852), .B(n8851), .X(n8849) );
  nand_x1_sg U59281 ( .A(n8851), .B(n8852), .X(n8850) );
  nor_x1_sg U59282 ( .A(n9672), .B(n9671), .X(n9669) );
  nand_x1_sg U59283 ( .A(n9671), .B(n9672), .X(n9670) );
  nor_x1_sg U59284 ( .A(n10491), .B(n10490), .X(n10488) );
  nand_x1_sg U59285 ( .A(n10490), .B(n10491), .X(n10489) );
  nor_x1_sg U59286 ( .A(n11310), .B(n11309), .X(n11307) );
  nand_x1_sg U59287 ( .A(n11309), .B(n11310), .X(n11308) );
  nor_x1_sg U59288 ( .A(n12129), .B(n12128), .X(n12126) );
  nand_x1_sg U59289 ( .A(n12128), .B(n12129), .X(n12127) );
  nor_x1_sg U59290 ( .A(n12948), .B(n12947), .X(n12945) );
  nand_x1_sg U59291 ( .A(n12947), .B(n12948), .X(n12946) );
  nor_x1_sg U59292 ( .A(n13767), .B(n13766), .X(n13764) );
  nand_x1_sg U59293 ( .A(n13766), .B(n13767), .X(n13765) );
  nor_x1_sg U59294 ( .A(n14586), .B(n14585), .X(n14583) );
  nand_x1_sg U59295 ( .A(n14585), .B(n14586), .X(n14584) );
  nor_x1_sg U59296 ( .A(n15405), .B(n15404), .X(n15402) );
  nand_x1_sg U59297 ( .A(n15404), .B(n15405), .X(n15403) );
  nor_x1_sg U59298 ( .A(n16224), .B(n16223), .X(n16221) );
  nand_x1_sg U59299 ( .A(n16223), .B(n16224), .X(n16222) );
  nor_x1_sg U59300 ( .A(n17040), .B(n17039), .X(n17037) );
  nand_x1_sg U59301 ( .A(n17039), .B(n17040), .X(n17038) );
  nor_x1_sg U59302 ( .A(n17862), .B(n17861), .X(n17859) );
  nand_x1_sg U59303 ( .A(n17861), .B(n17862), .X(n17860) );
  nor_x1_sg U59304 ( .A(n18683), .B(n18682), .X(n18680) );
  nand_x1_sg U59305 ( .A(n18682), .B(n18683), .X(n18681) );
  nor_x1_sg U59306 ( .A(n46906), .B(n46901), .X(n7164) );
  nor_x1_sg U59307 ( .A(n7166), .B(n7165), .X(n7163) );
  inv_x1_sg U59308 ( .A(n7165), .X(n46906) );
  nor_x1_sg U59309 ( .A(n50340), .B(n50334), .X(n16989) );
  nor_x1_sg U59310 ( .A(n16991), .B(n16990), .X(n16988) );
  inv_x1_sg U59311 ( .A(n16990), .X(n50340) );
  nor_x1_sg U59312 ( .A(n47199), .B(n47186), .X(n7983) );
  nor_x1_sg U59313 ( .A(n7985), .B(n7984), .X(n7982) );
  inv_x1_sg U59314 ( .A(n7984), .X(n47199) );
  nor_x1_sg U59315 ( .A(n47484), .B(n47471), .X(n8801) );
  nor_x1_sg U59316 ( .A(n8803), .B(n8802), .X(n8800) );
  inv_x1_sg U59317 ( .A(n8802), .X(n47484) );
  nor_x1_sg U59318 ( .A(n47769), .B(n47756), .X(n9621) );
  nor_x1_sg U59319 ( .A(n9623), .B(n9622), .X(n9620) );
  inv_x1_sg U59320 ( .A(n9622), .X(n47769) );
  nor_x1_sg U59321 ( .A(n48054), .B(n48041), .X(n10440) );
  nor_x1_sg U59322 ( .A(n10442), .B(n10441), .X(n10439) );
  inv_x1_sg U59323 ( .A(n10441), .X(n48054) );
  nor_x1_sg U59324 ( .A(n48339), .B(n48326), .X(n11259) );
  nor_x1_sg U59325 ( .A(n11261), .B(n11260), .X(n11258) );
  inv_x1_sg U59326 ( .A(n11260), .X(n48339) );
  nor_x1_sg U59327 ( .A(n48624), .B(n48611), .X(n12078) );
  nor_x1_sg U59328 ( .A(n12080), .B(n12079), .X(n12077) );
  inv_x1_sg U59329 ( .A(n12079), .X(n48624) );
  nor_x1_sg U59330 ( .A(n48910), .B(n48897), .X(n12897) );
  nor_x1_sg U59331 ( .A(n12899), .B(n12898), .X(n12896) );
  inv_x1_sg U59332 ( .A(n12898), .X(n48910) );
  nor_x1_sg U59333 ( .A(n49197), .B(n49184), .X(n13716) );
  nor_x1_sg U59334 ( .A(n13718), .B(n13717), .X(n13715) );
  inv_x1_sg U59335 ( .A(n13717), .X(n49197) );
  nor_x1_sg U59336 ( .A(n49483), .B(n49470), .X(n14535) );
  nor_x1_sg U59337 ( .A(n14537), .B(n14536), .X(n14534) );
  inv_x1_sg U59338 ( .A(n14536), .X(n49483) );
  nor_x1_sg U59339 ( .A(n49769), .B(n49756), .X(n15354) );
  nor_x1_sg U59340 ( .A(n15356), .B(n15355), .X(n15353) );
  inv_x1_sg U59341 ( .A(n15355), .X(n49769) );
  nor_x1_sg U59342 ( .A(n50055), .B(n50042), .X(n16173) );
  nor_x1_sg U59343 ( .A(n16175), .B(n16174), .X(n16172) );
  inv_x1_sg U59344 ( .A(n16174), .X(n50055) );
  nor_x1_sg U59345 ( .A(n50629), .B(n50616), .X(n17811) );
  nor_x1_sg U59346 ( .A(n17813), .B(n17812), .X(n17810) );
  inv_x1_sg U59347 ( .A(n17812), .X(n50629) );
  nor_x1_sg U59348 ( .A(n50916), .B(n50903), .X(n18632) );
  nor_x1_sg U59349 ( .A(n18634), .B(n18633), .X(n18631) );
  inv_x1_sg U59350 ( .A(n18633), .X(n50916) );
  nor_x1_sg U59351 ( .A(n46993), .B(n46913), .X(n7327) );
  nor_x1_sg U59352 ( .A(n7329), .B(n7330), .X(n7328) );
  inv_x1_sg U59353 ( .A(n7329), .X(n46913) );
  nor_x1_sg U59354 ( .A(n47282), .B(n47206), .X(n8145) );
  nor_x1_sg U59355 ( .A(n8147), .B(n8148), .X(n8146) );
  inv_x1_sg U59356 ( .A(n8147), .X(n47206) );
  nor_x1_sg U59357 ( .A(n47567), .B(n47491), .X(n8963) );
  nor_x1_sg U59358 ( .A(n8965), .B(n8966), .X(n8964) );
  inv_x1_sg U59359 ( .A(n8965), .X(n47491) );
  nor_x1_sg U59360 ( .A(n47852), .B(n47776), .X(n9783) );
  nor_x1_sg U59361 ( .A(n9785), .B(n9786), .X(n9784) );
  inv_x1_sg U59362 ( .A(n9785), .X(n47776) );
  nor_x1_sg U59363 ( .A(n48137), .B(n48061), .X(n10602) );
  nor_x1_sg U59364 ( .A(n10604), .B(n10605), .X(n10603) );
  inv_x1_sg U59365 ( .A(n10604), .X(n48061) );
  nor_x1_sg U59366 ( .A(n48422), .B(n48346), .X(n11421) );
  nor_x1_sg U59367 ( .A(n11423), .B(n11424), .X(n11422) );
  inv_x1_sg U59368 ( .A(n11423), .X(n48346) );
  nor_x1_sg U59369 ( .A(n48707), .B(n48631), .X(n12240) );
  nor_x1_sg U59370 ( .A(n12242), .B(n12243), .X(n12241) );
  inv_x1_sg U59371 ( .A(n12242), .X(n48631) );
  nor_x1_sg U59372 ( .A(n48993), .B(n48917), .X(n13059) );
  nor_x1_sg U59373 ( .A(n13061), .B(n13062), .X(n13060) );
  inv_x1_sg U59374 ( .A(n13061), .X(n48917) );
  nor_x1_sg U59375 ( .A(n49280), .B(n49204), .X(n13878) );
  nor_x1_sg U59376 ( .A(n13880), .B(n13881), .X(n13879) );
  inv_x1_sg U59377 ( .A(n13880), .X(n49204) );
  nor_x1_sg U59378 ( .A(n49566), .B(n49490), .X(n14697) );
  nor_x1_sg U59379 ( .A(n14699), .B(n14700), .X(n14698) );
  inv_x1_sg U59380 ( .A(n14699), .X(n49490) );
  nor_x1_sg U59381 ( .A(n49852), .B(n49776), .X(n15516) );
  nor_x1_sg U59382 ( .A(n15518), .B(n15519), .X(n15517) );
  inv_x1_sg U59383 ( .A(n15518), .X(n49776) );
  nor_x1_sg U59384 ( .A(n50138), .B(n50062), .X(n16335) );
  nor_x1_sg U59385 ( .A(n16337), .B(n16338), .X(n16336) );
  inv_x1_sg U59386 ( .A(n16337), .X(n50062) );
  nor_x1_sg U59387 ( .A(n50712), .B(n50636), .X(n17973) );
  nor_x1_sg U59388 ( .A(n17975), .B(n17976), .X(n17974) );
  inv_x1_sg U59389 ( .A(n17975), .X(n50636) );
  nor_x1_sg U59390 ( .A(n50999), .B(n50923), .X(n18794) );
  nor_x1_sg U59391 ( .A(n18796), .B(n18797), .X(n18795) );
  inv_x1_sg U59392 ( .A(n18796), .X(n50923) );
  inv_x1_sg U59393 ( .A(n6947), .X(n47048) );
  nor_x1_sg U59394 ( .A(n7578), .B(n7579), .X(n7577) );
  inv_x1_sg U59395 ( .A(n7764), .X(n47335) );
  nor_x1_sg U59396 ( .A(n8396), .B(n8397), .X(n8395) );
  inv_x1_sg U59397 ( .A(n8582), .X(n47620) );
  nor_x1_sg U59398 ( .A(n9214), .B(n9215), .X(n9213) );
  inv_x1_sg U59399 ( .A(n9402), .X(n47905) );
  nor_x1_sg U59400 ( .A(n10034), .B(n10035), .X(n10033) );
  inv_x1_sg U59401 ( .A(n10221), .X(n48190) );
  nor_x1_sg U59402 ( .A(n10853), .B(n10854), .X(n10852) );
  inv_x1_sg U59403 ( .A(n11040), .X(n48475) );
  nor_x1_sg U59404 ( .A(n11672), .B(n11673), .X(n11671) );
  inv_x1_sg U59405 ( .A(n11859), .X(n48760) );
  nor_x1_sg U59406 ( .A(n12491), .B(n12492), .X(n12490) );
  inv_x1_sg U59407 ( .A(n12678), .X(n49046) );
  nor_x1_sg U59408 ( .A(n13310), .B(n13311), .X(n13309) );
  inv_x1_sg U59409 ( .A(n13497), .X(n49333) );
  nor_x1_sg U59410 ( .A(n14129), .B(n14130), .X(n14128) );
  inv_x1_sg U59411 ( .A(n14316), .X(n49619) );
  nor_x1_sg U59412 ( .A(n14948), .B(n14949), .X(n14947) );
  inv_x1_sg U59413 ( .A(n15135), .X(n49905) );
  nor_x1_sg U59414 ( .A(n15767), .B(n15768), .X(n15766) );
  inv_x1_sg U59415 ( .A(n15954), .X(n50191) );
  nor_x1_sg U59416 ( .A(n16586), .B(n16587), .X(n16585) );
  inv_x1_sg U59417 ( .A(n16771), .X(n50476) );
  nor_x1_sg U59418 ( .A(n17403), .B(n17404), .X(n17402) );
  inv_x1_sg U59419 ( .A(n17592), .X(n50765) );
  nor_x1_sg U59420 ( .A(n18224), .B(n18225), .X(n18223) );
  inv_x1_sg U59421 ( .A(n18413), .X(n51052) );
  nor_x1_sg U59422 ( .A(n19045), .B(n19046), .X(n19044) );
  nor_x1_sg U59423 ( .A(n8035), .B(n41777), .X(n8369) );
  nor_x1_sg U59424 ( .A(n40108), .B(n41776), .X(n9187) );
  nor_x1_sg U59425 ( .A(n9673), .B(n41775), .X(n10007) );
  nor_x1_sg U59426 ( .A(n10492), .B(n41774), .X(n10826) );
  nor_x1_sg U59427 ( .A(n40114), .B(n41773), .X(n11645) );
  nor_x1_sg U59428 ( .A(n12130), .B(n41772), .X(n12464) );
  nor_x1_sg U59429 ( .A(n12949), .B(n41771), .X(n13283) );
  nor_x1_sg U59430 ( .A(n40119), .B(n41770), .X(n14102) );
  nor_x1_sg U59431 ( .A(n14587), .B(n41769), .X(n14921) );
  nor_x1_sg U59432 ( .A(n15406), .B(n41768), .X(n15740) );
  nor_x1_sg U59433 ( .A(n40126), .B(n41767), .X(n16559) );
  nor_x1_sg U59434 ( .A(n40131), .B(n39390), .X(n18197) );
  nor_x1_sg U59435 ( .A(n18684), .B(n41766), .X(n19018) );
  nor_x1_sg U59436 ( .A(n39606), .B(n6834), .X(n7371) );
  nor_x1_sg U59437 ( .A(n39602), .B(n40303), .X(n17196) );
  nor_x1_sg U59438 ( .A(n22936), .B(n42319), .X(n22943) );
  nor_x1_sg U59439 ( .A(n23213), .B(n9081), .X(n23220) );
  nor_x1_sg U59440 ( .A(n23493), .B(n42318), .X(n23500) );
  nor_x1_sg U59441 ( .A(n23772), .B(n10720), .X(n23779) );
  nor_x1_sg U59442 ( .A(n24051), .B(n42317), .X(n24058) );
  nor_x1_sg U59443 ( .A(n24330), .B(n12358), .X(n24337) );
  nor_x1_sg U59444 ( .A(n24609), .B(n42316), .X(n24616) );
  nor_x1_sg U59445 ( .A(n24887), .B(n13996), .X(n24894) );
  nor_x1_sg U59446 ( .A(n25166), .B(n42315), .X(n25173) );
  nor_x1_sg U59447 ( .A(n25445), .B(n15634), .X(n25452) );
  nor_x1_sg U59448 ( .A(n25724), .B(n42314), .X(n25731) );
  nor_x1_sg U59449 ( .A(n25990), .B(n42235), .X(n25997) );
  nor_x1_sg U59450 ( .A(n26276), .B(n18091), .X(n26284) );
  nor_x1_sg U59451 ( .A(n26561), .B(n42313), .X(n26568) );
  nor_x1_sg U59452 ( .A(n22922), .B(n42161), .X(n22929) );
  nor_x1_sg U59453 ( .A(n23199), .B(n8936), .X(n23206) );
  nor_x1_sg U59454 ( .A(n23479), .B(n9756), .X(n23486) );
  nor_x1_sg U59455 ( .A(n23758), .B(n10575), .X(n23765) );
  nor_x1_sg U59456 ( .A(n24037), .B(n11394), .X(n24044) );
  nor_x1_sg U59457 ( .A(n24316), .B(n12213), .X(n24323) );
  nor_x1_sg U59458 ( .A(n24595), .B(n13032), .X(n24602) );
  nor_x1_sg U59459 ( .A(n24873), .B(n13851), .X(n24880) );
  nor_x1_sg U59460 ( .A(n25152), .B(n14670), .X(n25159) );
  nor_x1_sg U59461 ( .A(n25431), .B(n42160), .X(n25438) );
  nor_x1_sg U59462 ( .A(n25710), .B(n16308), .X(n25717) );
  nor_x1_sg U59463 ( .A(n25978), .B(n17125), .X(n25984) );
  nor_x1_sg U59464 ( .A(n26260), .B(n17946), .X(n26268) );
  nor_x1_sg U59465 ( .A(n26547), .B(n18767), .X(n26554) );
  nor_x1_sg U59466 ( .A(n39548), .B(n41915), .X(n8123) );
  nor_x1_sg U59467 ( .A(n41735), .B(n41916), .X(n8941) );
  nor_x1_sg U59468 ( .A(n39550), .B(n41907), .X(n9761) );
  nor_x1_sg U59469 ( .A(n41727), .B(n41909), .X(n10580) );
  nor_x1_sg U59470 ( .A(n39558), .B(n41913), .X(n11399) );
  nor_x1_sg U59471 ( .A(n41730), .B(n41914), .X(n12218) );
  nor_x1_sg U59472 ( .A(n39555), .B(n41908), .X(n13037) );
  nor_x1_sg U59473 ( .A(n39556), .B(n41911), .X(n13856) );
  nor_x1_sg U59474 ( .A(n39553), .B(n41917), .X(n14675) );
  nor_x1_sg U59475 ( .A(n39551), .B(n41904), .X(n15494) );
  nor_x1_sg U59476 ( .A(n41732), .B(n41905), .X(n16313) );
  nor_x1_sg U59477 ( .A(n41739), .B(n41860), .X(n17130) );
  nor_x1_sg U59478 ( .A(n39546), .B(n41912), .X(n17951) );
  nor_x1_sg U59479 ( .A(n39547), .B(n41906), .X(n18772) );
  nor_x1_sg U59480 ( .A(n41780), .B(n40368), .X(n7131) );
  nor_x1_sg U59481 ( .A(n39720), .B(n41847), .X(n7949) );
  nor_x1_sg U59482 ( .A(n39717), .B(n39069), .X(n8767) );
  nor_x1_sg U59483 ( .A(n39714), .B(n39073), .X(n9587) );
  nor_x1_sg U59484 ( .A(n39711), .B(n41855), .X(n10406) );
  nor_x1_sg U59485 ( .A(n41790), .B(n39072), .X(n11225) );
  nor_x1_sg U59486 ( .A(n39704), .B(n41857), .X(n12044) );
  nor_x1_sg U59487 ( .A(n39702), .B(n41859), .X(n12863) );
  nor_x1_sg U59488 ( .A(n41796), .B(n39071), .X(n13682) );
  nor_x1_sg U59489 ( .A(n39696), .B(n39066), .X(n14501) );
  nor_x1_sg U59490 ( .A(n39693), .B(n41765), .X(n15320) );
  nor_x1_sg U59491 ( .A(n39690), .B(n39067), .X(n16139) );
  nor_x1_sg U59492 ( .A(n39687), .B(n40365), .X(n17777) );
  nor_x1_sg U59493 ( .A(n39684), .B(n39068), .X(n18598) );
  nor_x1_sg U59494 ( .A(n22908), .B(n42324), .X(n22915) );
  nor_x1_sg U59495 ( .A(n23185), .B(n42323), .X(n23192) );
  nor_x1_sg U59496 ( .A(n23465), .B(n42322), .X(n23472) );
  nor_x1_sg U59497 ( .A(n23744), .B(n10311), .X(n23751) );
  nor_x1_sg U59498 ( .A(n24023), .B(n11130), .X(n24030) );
  nor_x1_sg U59499 ( .A(n24302), .B(n11949), .X(n24309) );
  nor_x1_sg U59500 ( .A(n24581), .B(n12768), .X(n24588) );
  nor_x1_sg U59501 ( .A(n24859), .B(n13587), .X(n24866) );
  nor_x1_sg U59502 ( .A(n25138), .B(n14406), .X(n25145) );
  nor_x1_sg U59503 ( .A(n25417), .B(n15225), .X(n25424) );
  nor_x1_sg U59504 ( .A(n25696), .B(n16044), .X(n25703) );
  nor_x1_sg U59505 ( .A(n25965), .B(n42236), .X(n25971) );
  nor_x1_sg U59506 ( .A(n26244), .B(n42321), .X(n26252) );
  nor_x1_sg U59507 ( .A(n26533), .B(n42320), .X(n26540) );
  nor_x1_sg U59508 ( .A(n50286), .B(n39316), .X(n16904) );
  nor_x1_sg U59509 ( .A(n39317), .B(n16906), .X(n16905) );
  nor_x1_sg U59510 ( .A(n46854), .B(n39289), .X(n7077) );
  nor_x1_sg U59511 ( .A(n39290), .B(n7079), .X(n7078) );
  nor_x1_sg U59512 ( .A(n47147), .B(n39314), .X(n7895) );
  nor_x1_sg U59513 ( .A(n39315), .B(n7897), .X(n7896) );
  nor_x1_sg U59514 ( .A(n47432), .B(n39023), .X(n8713) );
  nor_x1_sg U59515 ( .A(n39313), .B(n8715), .X(n8714) );
  nor_x1_sg U59516 ( .A(n47717), .B(n39311), .X(n9533) );
  nor_x1_sg U59517 ( .A(n39312), .B(n9535), .X(n9534) );
  nor_x1_sg U59518 ( .A(n48002), .B(n39309), .X(n10352) );
  nor_x1_sg U59519 ( .A(n39310), .B(n10354), .X(n10353) );
  nor_x1_sg U59520 ( .A(n48287), .B(n39307), .X(n11171) );
  nor_x1_sg U59521 ( .A(n39308), .B(n11173), .X(n11172) );
  nor_x1_sg U59522 ( .A(n48572), .B(n39305), .X(n11990) );
  nor_x1_sg U59523 ( .A(n39306), .B(n11992), .X(n11991) );
  nor_x1_sg U59524 ( .A(n48858), .B(n39303), .X(n12809) );
  nor_x1_sg U59525 ( .A(n39304), .B(n12811), .X(n12810) );
  nor_x1_sg U59526 ( .A(n49145), .B(n39301), .X(n13628) );
  nor_x1_sg U59527 ( .A(n39302), .B(n13630), .X(n13629) );
  nor_x1_sg U59528 ( .A(n49431), .B(n39299), .X(n14447) );
  nor_x1_sg U59529 ( .A(n39300), .B(n14449), .X(n14448) );
  nor_x1_sg U59530 ( .A(n49716), .B(n39297), .X(n15266) );
  nor_x1_sg U59531 ( .A(n39298), .B(n15268), .X(n15267) );
  nor_x1_sg U59532 ( .A(n50003), .B(n39295), .X(n16085) );
  nor_x1_sg U59533 ( .A(n39296), .B(n16087), .X(n16086) );
  nor_x1_sg U59534 ( .A(n50577), .B(n39291), .X(n17723) );
  nor_x1_sg U59535 ( .A(n39292), .B(n17725), .X(n17724) );
  nor_x1_sg U59536 ( .A(n50864), .B(n39293), .X(n18544) );
  nor_x1_sg U59537 ( .A(n39294), .B(n18546), .X(n18545) );
  nor_x1_sg U59538 ( .A(n17165), .B(n39018), .X(n17163) );
  nor_x1_sg U59539 ( .A(n16992), .B(n50331), .X(n17164) );
  nor_x1_sg U59540 ( .A(n7340), .B(n39019), .X(n7338) );
  nor_x1_sg U59541 ( .A(n7167), .B(n46898), .X(n7339) );
  nor_x1_sg U59542 ( .A(n8158), .B(n39022), .X(n8156) );
  nor_x1_sg U59543 ( .A(n7986), .B(n47193), .X(n8157) );
  nor_x1_sg U59544 ( .A(n8976), .B(n39017), .X(n8974) );
  nor_x1_sg U59545 ( .A(n8804), .B(n47478), .X(n8975) );
  nor_x1_sg U59546 ( .A(n9796), .B(n39016), .X(n9794) );
  nor_x1_sg U59547 ( .A(n9624), .B(n47763), .X(n9795) );
  nor_x1_sg U59548 ( .A(n10615), .B(n39015), .X(n10613) );
  nor_x1_sg U59549 ( .A(n10443), .B(n48048), .X(n10614) );
  nor_x1_sg U59550 ( .A(n11434), .B(n39014), .X(n11432) );
  nor_x1_sg U59551 ( .A(n11262), .B(n48333), .X(n11433) );
  nor_x1_sg U59552 ( .A(n12253), .B(n39013), .X(n12251) );
  nor_x1_sg U59553 ( .A(n12081), .B(n48618), .X(n12252) );
  nor_x1_sg U59554 ( .A(n13072), .B(n39012), .X(n13070) );
  nor_x1_sg U59555 ( .A(n12900), .B(n48904), .X(n13071) );
  nor_x1_sg U59556 ( .A(n13891), .B(n39011), .X(n13889) );
  nor_x1_sg U59557 ( .A(n13719), .B(n49191), .X(n13890) );
  nor_x1_sg U59558 ( .A(n14710), .B(n39010), .X(n14708) );
  nor_x1_sg U59559 ( .A(n14538), .B(n49477), .X(n14709) );
  nor_x1_sg U59560 ( .A(n15529), .B(n39021), .X(n15527) );
  nor_x1_sg U59561 ( .A(n15357), .B(n49763), .X(n15528) );
  nor_x1_sg U59562 ( .A(n16348), .B(n39009), .X(n16346) );
  nor_x1_sg U59563 ( .A(n16176), .B(n50049), .X(n16347) );
  nor_x1_sg U59564 ( .A(n17986), .B(n39020), .X(n17984) );
  nor_x1_sg U59565 ( .A(n17814), .B(n50623), .X(n17985) );
  nor_x1_sg U59566 ( .A(n18807), .B(n39008), .X(n18805) );
  nor_x1_sg U59567 ( .A(n18635), .B(n50910), .X(n18806) );
  nor_x1_sg U59568 ( .A(n46856), .B(n46865), .X(n7099) );
  nor_x1_sg U59569 ( .A(n7101), .B(n7102), .X(n7100) );
  nor_x1_sg U59570 ( .A(n47149), .B(n47158), .X(n7917) );
  nor_x1_sg U59571 ( .A(n7919), .B(n7920), .X(n7918) );
  nor_x1_sg U59572 ( .A(n47434), .B(n47443), .X(n8735) );
  nor_x1_sg U59573 ( .A(n8737), .B(n8738), .X(n8736) );
  nor_x1_sg U59574 ( .A(n47719), .B(n47728), .X(n9555) );
  nor_x1_sg U59575 ( .A(n9557), .B(n9558), .X(n9556) );
  nor_x1_sg U59576 ( .A(n48004), .B(n48013), .X(n10374) );
  nor_x1_sg U59577 ( .A(n10376), .B(n10377), .X(n10375) );
  nor_x1_sg U59578 ( .A(n48289), .B(n48298), .X(n11193) );
  nor_x1_sg U59579 ( .A(n11195), .B(n11196), .X(n11194) );
  nor_x1_sg U59580 ( .A(n48574), .B(n48583), .X(n12012) );
  nor_x1_sg U59581 ( .A(n12014), .B(n12015), .X(n12013) );
  nor_x1_sg U59582 ( .A(n48860), .B(n48869), .X(n12831) );
  nor_x1_sg U59583 ( .A(n12833), .B(n12834), .X(n12832) );
  nor_x1_sg U59584 ( .A(n49147), .B(n49156), .X(n13650) );
  nor_x1_sg U59585 ( .A(n13652), .B(n13653), .X(n13651) );
  nor_x1_sg U59586 ( .A(n49433), .B(n49442), .X(n14469) );
  nor_x1_sg U59587 ( .A(n14471), .B(n14472), .X(n14470) );
  nor_x1_sg U59588 ( .A(n49718), .B(n49727), .X(n15288) );
  nor_x1_sg U59589 ( .A(n15290), .B(n15291), .X(n15289) );
  nor_x1_sg U59590 ( .A(n50005), .B(n50014), .X(n16107) );
  nor_x1_sg U59591 ( .A(n16109), .B(n16110), .X(n16108) );
  nor_x1_sg U59592 ( .A(n50288), .B(n50298), .X(n16924) );
  nor_x1_sg U59593 ( .A(n16926), .B(n16927), .X(n16925) );
  nor_x1_sg U59594 ( .A(n50579), .B(n50588), .X(n17745) );
  nor_x1_sg U59595 ( .A(n17747), .B(n17748), .X(n17746) );
  nor_x1_sg U59596 ( .A(n50866), .B(n50875), .X(n18566) );
  nor_x1_sg U59597 ( .A(n18568), .B(n18569), .X(n18567) );
  nor_x1_sg U59598 ( .A(n39366), .B(n40308), .X(n8007) );
  nor_x1_sg U59599 ( .A(n39368), .B(n41754), .X(n8825) );
  nor_x1_sg U59600 ( .A(n39370), .B(n41852), .X(n9645) );
  nor_x1_sg U59601 ( .A(n39372), .B(n39074), .X(n10464) );
  nor_x1_sg U59602 ( .A(n39374), .B(n41850), .X(n11283) );
  nor_x1_sg U59603 ( .A(n39376), .B(n39075), .X(n12102) );
  nor_x1_sg U59604 ( .A(n39378), .B(n39076), .X(n12921) );
  nor_x1_sg U59605 ( .A(n39380), .B(n41848), .X(n13740) );
  nor_x1_sg U59606 ( .A(n39382), .B(n41759), .X(n14559) );
  nor_x1_sg U59607 ( .A(n39384), .B(n39070), .X(n15378) );
  nor_x1_sg U59608 ( .A(n39386), .B(n41764), .X(n16197) );
  nor_x1_sg U59609 ( .A(n39390), .B(n40363), .X(n17835) );
  nor_x1_sg U59610 ( .A(n39388), .B(n41762), .X(n18656) );
  nor_x1_sg U59611 ( .A(n39893), .B(n41777), .X(n7823) );
  nor_x1_sg U59612 ( .A(n39861), .B(n41776), .X(n8641) );
  nor_x1_sg U59613 ( .A(n41689), .B(n41775), .X(n9461) );
  nor_x1_sg U59614 ( .A(n41685), .B(n41774), .X(n10280) );
  nor_x1_sg U59615 ( .A(n41683), .B(n41773), .X(n11099) );
  nor_x1_sg U59616 ( .A(n41681), .B(n41772), .X(n11918) );
  nor_x1_sg U59617 ( .A(n41679), .B(n41771), .X(n12737) );
  nor_x1_sg U59618 ( .A(n41677), .B(n41770), .X(n13556) );
  nor_x1_sg U59619 ( .A(n41675), .B(n41769), .X(n14375) );
  nor_x1_sg U59620 ( .A(n41662), .B(n41768), .X(n15194) );
  nor_x1_sg U59621 ( .A(n41673), .B(n41767), .X(n16013) );
  nor_x1_sg U59622 ( .A(n41669), .B(n41755), .X(n17651) );
  nor_x1_sg U59623 ( .A(n41667), .B(n41766), .X(n18472) );
  nor_x1_sg U59624 ( .A(n41578), .B(n40306), .X(n8354) );
  nor_x1_sg U59625 ( .A(n41577), .B(n41754), .X(n9172) );
  nor_x1_sg U59626 ( .A(n41576), .B(n41756), .X(n9992) );
  nor_x1_sg U59627 ( .A(n41575), .B(n41757), .X(n10811) );
  nor_x1_sg U59628 ( .A(n41582), .B(n41758), .X(n11630) );
  nor_x1_sg U59629 ( .A(n41581), .B(n41763), .X(n12449) );
  nor_x1_sg U59630 ( .A(n41580), .B(n41760), .X(n13268) );
  nor_x1_sg U59631 ( .A(n41579), .B(n41761), .X(n14087) );
  nor_x1_sg U59632 ( .A(n41586), .B(n41837), .X(n14906) );
  nor_x1_sg U59633 ( .A(n41585), .B(n41765), .X(n15725) );
  nor_x1_sg U59634 ( .A(n41584), .B(n41839), .X(n16544) );
  nor_x1_sg U59635 ( .A(n41587), .B(n40363), .X(n18182) );
  nor_x1_sg U59636 ( .A(n41583), .B(n41841), .X(n19003) );
  nor_x1_sg U59637 ( .A(n39730), .B(n40559), .X(n8189) );
  nor_x1_sg U59638 ( .A(n39733), .B(n40555), .X(n9007) );
  nor_x1_sg U59639 ( .A(n39736), .B(n40553), .X(n9827) );
  nor_x1_sg U59640 ( .A(n41650), .B(n40547), .X(n10646) );
  nor_x1_sg U59641 ( .A(n39742), .B(n40543), .X(n11465) );
  nor_x1_sg U59642 ( .A(n39745), .B(n40539), .X(n12284) );
  nor_x1_sg U59643 ( .A(n39748), .B(n40535), .X(n13103) );
  nor_x1_sg U59644 ( .A(n39751), .B(n40533), .X(n13922) );
  nor_x1_sg U59645 ( .A(n41653), .B(n40527), .X(n14741) );
  nor_x1_sg U59646 ( .A(n39757), .B(n40524), .X(n15560) );
  nor_x1_sg U59647 ( .A(n39760), .B(n40519), .X(n16379) );
  nor_x1_sg U59648 ( .A(n41647), .B(n40515), .X(n18017) );
  nor_x1_sg U59649 ( .A(n39766), .B(n40511), .X(n18838) );
  nor_x1_sg U59650 ( .A(n41666), .B(n41903), .X(n7536) );
  nor_x1_sg U59651 ( .A(n41709), .B(n41861), .X(n7305) );
  nor_x1_sg U59652 ( .A(n41693), .B(n40312), .X(n17361) );
  nor_x1_sg U59653 ( .A(n22697), .B(n47127), .X(n5861) );
  nor_x1_sg U59654 ( .A(n16992), .B(n16820), .X(n16986) );
  nor_x1_sg U59655 ( .A(n7986), .B(n7813), .X(n7980) );
  nor_x1_sg U59656 ( .A(n8804), .B(n39313), .X(n8798) );
  nor_x1_sg U59657 ( .A(n9624), .B(n9451), .X(n9618) );
  nor_x1_sg U59658 ( .A(n10443), .B(n10270), .X(n10437) );
  nor_x1_sg U59659 ( .A(n11262), .B(n11089), .X(n11256) );
  nor_x1_sg U59660 ( .A(n12081), .B(n11908), .X(n12075) );
  nor_x1_sg U59661 ( .A(n12900), .B(n12727), .X(n12894) );
  nor_x1_sg U59662 ( .A(n13719), .B(n13546), .X(n13713) );
  nor_x1_sg U59663 ( .A(n14538), .B(n14365), .X(n14532) );
  nor_x1_sg U59664 ( .A(n15357), .B(n15184), .X(n15351) );
  nor_x1_sg U59665 ( .A(n16176), .B(n16003), .X(n16170) );
  nor_x1_sg U59666 ( .A(n17814), .B(n17641), .X(n17808) );
  nor_x1_sg U59667 ( .A(n18635), .B(n18462), .X(n18629) );
  nor_x1_sg U59668 ( .A(n7167), .B(n6996), .X(n7161) );
  nor_x1_sg U59669 ( .A(n7217), .B(n7075), .X(n7211) );
  nor_x1_sg U59670 ( .A(n17042), .B(n16902), .X(n17036) );
  nor_x1_sg U59671 ( .A(n8036), .B(n7893), .X(n8030) );
  nor_x1_sg U59672 ( .A(n8854), .B(n8711), .X(n8848) );
  nor_x1_sg U59673 ( .A(n9674), .B(n9531), .X(n9668) );
  nor_x1_sg U59674 ( .A(n10493), .B(n10350), .X(n10487) );
  nor_x1_sg U59675 ( .A(n11312), .B(n11169), .X(n11306) );
  nor_x1_sg U59676 ( .A(n12131), .B(n11988), .X(n12125) );
  nor_x1_sg U59677 ( .A(n12950), .B(n12807), .X(n12944) );
  nor_x1_sg U59678 ( .A(n13769), .B(n13626), .X(n13763) );
  nor_x1_sg U59679 ( .A(n14588), .B(n14445), .X(n14582) );
  nor_x1_sg U59680 ( .A(n15407), .B(n15264), .X(n15401) );
  nor_x1_sg U59681 ( .A(n16226), .B(n16083), .X(n16220) );
  nor_x1_sg U59682 ( .A(n17864), .B(n17721), .X(n17858) );
  nor_x1_sg U59683 ( .A(n18685), .B(n18542), .X(n18679) );
  inv_x1_sg U59684 ( .A(n7521), .X(n47058) );
  nor_x1_sg U59685 ( .A(n7519), .B(n7520), .X(n7518) );
  inv_x1_sg U59686 ( .A(n8339), .X(n47344) );
  nor_x1_sg U59687 ( .A(n8337), .B(n8338), .X(n8336) );
  inv_x1_sg U59688 ( .A(n9157), .X(n47629) );
  nor_x1_sg U59689 ( .A(n9155), .B(n9156), .X(n9154) );
  inv_x1_sg U59690 ( .A(n9977), .X(n47914) );
  nor_x1_sg U59691 ( .A(n9975), .B(n9976), .X(n9974) );
  inv_x1_sg U59692 ( .A(n10796), .X(n48199) );
  nor_x1_sg U59693 ( .A(n10794), .B(n10795), .X(n10793) );
  inv_x1_sg U59694 ( .A(n11615), .X(n48484) );
  nor_x1_sg U59695 ( .A(n11613), .B(n11614), .X(n11612) );
  inv_x1_sg U59696 ( .A(n12434), .X(n48769) );
  nor_x1_sg U59697 ( .A(n12432), .B(n12433), .X(n12431) );
  inv_x1_sg U59698 ( .A(n13253), .X(n49056) );
  nor_x1_sg U59699 ( .A(n13251), .B(n13252), .X(n13250) );
  inv_x1_sg U59700 ( .A(n14072), .X(n49342) );
  nor_x1_sg U59701 ( .A(n14070), .B(n14071), .X(n14069) );
  inv_x1_sg U59702 ( .A(n14891), .X(n49628) );
  nor_x1_sg U59703 ( .A(n14889), .B(n14890), .X(n14888) );
  inv_x1_sg U59704 ( .A(n15710), .X(n49914) );
  nor_x1_sg U59705 ( .A(n15708), .B(n15709), .X(n15707) );
  inv_x1_sg U59706 ( .A(n16529), .X(n50200) );
  nor_x1_sg U59707 ( .A(n16527), .B(n16528), .X(n16526) );
  inv_x1_sg U59708 ( .A(n17346), .X(n50485) );
  nor_x1_sg U59709 ( .A(n17344), .B(n17345), .X(n17343) );
  inv_x1_sg U59710 ( .A(n18167), .X(n50774) );
  nor_x1_sg U59711 ( .A(n18165), .B(n18166), .X(n18164) );
  inv_x1_sg U59712 ( .A(n18988), .X(n51061) );
  nor_x1_sg U59713 ( .A(n18986), .B(n18987), .X(n18985) );
  nand_x1_sg U59714 ( .A(n41419), .B(n42119), .X(n12551) );
  nand_x1_sg U59715 ( .A(n41420), .B(n42020), .X(n11732) );
  nor_x1_sg U59716 ( .A(n22950), .B(n7814), .X(n22957) );
  nor_x1_sg U59717 ( .A(n23227), .B(n8632), .X(n23234) );
  nor_x1_sg U59718 ( .A(n23507), .B(n9452), .X(n23514) );
  nor_x1_sg U59719 ( .A(n23786), .B(n10271), .X(n23793) );
  nor_x1_sg U59720 ( .A(n24065), .B(n11090), .X(n24072) );
  nor_x1_sg U59721 ( .A(n24344), .B(n11909), .X(n24351) );
  nor_x1_sg U59722 ( .A(n24623), .B(n12728), .X(n24630) );
  nor_x1_sg U59723 ( .A(n24901), .B(n13547), .X(n24908) );
  nor_x1_sg U59724 ( .A(n25180), .B(n14366), .X(n25187) );
  nor_x1_sg U59725 ( .A(n25459), .B(n15185), .X(n25466) );
  nor_x1_sg U59726 ( .A(n25738), .B(n16004), .X(n25745) );
  nor_x1_sg U59727 ( .A(n26292), .B(n17642), .X(n26300) );
  nor_x1_sg U59728 ( .A(n26575), .B(n18463), .X(n26582) );
  nor_x1_sg U59729 ( .A(n7186), .B(n46900), .X(n7166) );
  nor_x1_sg U59730 ( .A(n7189), .B(n7188), .X(n7186) );
  nand_x1_sg U59731 ( .A(n7188), .B(n7189), .X(n7187) );
  nor_x1_sg U59732 ( .A(n17011), .B(n50333), .X(n16991) );
  nor_x1_sg U59733 ( .A(n17014), .B(n17013), .X(n17011) );
  nand_x1_sg U59734 ( .A(n17013), .B(n17014), .X(n17012) );
  nor_x1_sg U59735 ( .A(n22656), .B(n6971), .X(n22653) );
  nor_x1_sg U59736 ( .A(n8005), .B(n47185), .X(n7985) );
  nor_x1_sg U59737 ( .A(n8008), .B(n8007), .X(n8005) );
  nand_x1_sg U59738 ( .A(n8007), .B(n8008), .X(n8006) );
  nor_x1_sg U59739 ( .A(n8823), .B(n47470), .X(n8803) );
  nor_x1_sg U59740 ( .A(n8826), .B(n8825), .X(n8823) );
  nand_x1_sg U59741 ( .A(n8825), .B(n8826), .X(n8824) );
  nor_x1_sg U59742 ( .A(n9643), .B(n47755), .X(n9623) );
  nor_x1_sg U59743 ( .A(n9646), .B(n9645), .X(n9643) );
  nand_x1_sg U59744 ( .A(n9645), .B(n9646), .X(n9644) );
  nor_x1_sg U59745 ( .A(n10462), .B(n48040), .X(n10442) );
  nor_x1_sg U59746 ( .A(n10465), .B(n10464), .X(n10462) );
  nand_x1_sg U59747 ( .A(n10464), .B(n10465), .X(n10463) );
  nor_x1_sg U59748 ( .A(n11281), .B(n48325), .X(n11261) );
  nor_x1_sg U59749 ( .A(n11284), .B(n11283), .X(n11281) );
  nand_x1_sg U59750 ( .A(n11283), .B(n11284), .X(n11282) );
  nor_x1_sg U59751 ( .A(n12100), .B(n48610), .X(n12080) );
  nor_x1_sg U59752 ( .A(n12103), .B(n12102), .X(n12100) );
  nand_x1_sg U59753 ( .A(n12102), .B(n12103), .X(n12101) );
  nor_x1_sg U59754 ( .A(n12919), .B(n48896), .X(n12899) );
  nor_x1_sg U59755 ( .A(n12922), .B(n12921), .X(n12919) );
  nand_x1_sg U59756 ( .A(n12921), .B(n12922), .X(n12920) );
  nor_x1_sg U59757 ( .A(n13738), .B(n49183), .X(n13718) );
  nor_x1_sg U59758 ( .A(n13741), .B(n13740), .X(n13738) );
  nand_x1_sg U59759 ( .A(n13740), .B(n13741), .X(n13739) );
  nor_x1_sg U59760 ( .A(n14557), .B(n49469), .X(n14537) );
  nor_x1_sg U59761 ( .A(n14560), .B(n14559), .X(n14557) );
  nand_x1_sg U59762 ( .A(n14559), .B(n14560), .X(n14558) );
  nor_x1_sg U59763 ( .A(n15376), .B(n49755), .X(n15356) );
  nor_x1_sg U59764 ( .A(n15379), .B(n15378), .X(n15376) );
  nand_x1_sg U59765 ( .A(n15378), .B(n15379), .X(n15377) );
  nor_x1_sg U59766 ( .A(n16195), .B(n50041), .X(n16175) );
  nor_x1_sg U59767 ( .A(n16198), .B(n16197), .X(n16195) );
  nand_x1_sg U59768 ( .A(n16197), .B(n16198), .X(n16196) );
  nor_x1_sg U59769 ( .A(n17833), .B(n50615), .X(n17813) );
  nor_x1_sg U59770 ( .A(n17836), .B(n17835), .X(n17833) );
  nand_x1_sg U59771 ( .A(n17835), .B(n17836), .X(n17834) );
  nor_x1_sg U59772 ( .A(n18654), .B(n50902), .X(n18634) );
  nor_x1_sg U59773 ( .A(n18657), .B(n18656), .X(n18654) );
  nand_x1_sg U59774 ( .A(n18656), .B(n18657), .X(n18655) );
  nand_x1_sg U59775 ( .A(n40220), .B(n51139), .X(n15827) );
  nor_x1_sg U59776 ( .A(n7279), .B(n42163), .X(n7278) );
  nor_x1_sg U59777 ( .A(n6962), .B(n46854), .X(n7277) );
  nand_x1_sg U59778 ( .A(n7252), .B(n40163), .X(n7279) );
  inv_x1_sg U59779 ( .A(n39358), .X(n49055) );
  nor_x1_sg U59780 ( .A(n8098), .B(n40105), .X(n8097) );
  nor_x1_sg U59781 ( .A(n7779), .B(n47147), .X(n8096) );
  nand_x1_sg U59782 ( .A(n8071), .B(n40243), .X(n8098) );
  nor_x1_sg U59783 ( .A(n8916), .B(n40107), .X(n8915) );
  nor_x1_sg U59784 ( .A(n8597), .B(n47432), .X(n8914) );
  nand_x1_sg U59785 ( .A(n8889), .B(n40248), .X(n8916) );
  nor_x1_sg U59786 ( .A(n9736), .B(n40109), .X(n9735) );
  nor_x1_sg U59787 ( .A(n9417), .B(n47717), .X(n9734) );
  nand_x1_sg U59788 ( .A(n9709), .B(n40254), .X(n9736) );
  nor_x1_sg U59789 ( .A(n10555), .B(n40112), .X(n10554) );
  nor_x1_sg U59790 ( .A(n10236), .B(n48002), .X(n10553) );
  nand_x1_sg U59791 ( .A(n10528), .B(n40257), .X(n10555) );
  nor_x1_sg U59792 ( .A(n11374), .B(n40113), .X(n11373) );
  nor_x1_sg U59793 ( .A(n11055), .B(n48287), .X(n11372) );
  nand_x1_sg U59794 ( .A(n11347), .B(n40265), .X(n11374) );
  nor_x1_sg U59795 ( .A(n12193), .B(n40115), .X(n12192) );
  nor_x1_sg U59796 ( .A(n11874), .B(n48572), .X(n12191) );
  nand_x1_sg U59797 ( .A(n12166), .B(n40269), .X(n12193) );
  nor_x1_sg U59798 ( .A(n13012), .B(n40118), .X(n13011) );
  nor_x1_sg U59799 ( .A(n12693), .B(n48858), .X(n13010) );
  nand_x1_sg U59800 ( .A(n12985), .B(n40272), .X(n13012) );
  nor_x1_sg U59801 ( .A(n13831), .B(n40120), .X(n13830) );
  nor_x1_sg U59802 ( .A(n13512), .B(n49145), .X(n13829) );
  nand_x1_sg U59803 ( .A(n13804), .B(n40278), .X(n13831) );
  nor_x1_sg U59804 ( .A(n14650), .B(n40121), .X(n14649) );
  nor_x1_sg U59805 ( .A(n14331), .B(n49431), .X(n14648) );
  nand_x1_sg U59806 ( .A(n14623), .B(n40283), .X(n14650) );
  nor_x1_sg U59807 ( .A(n15469), .B(n40123), .X(n15468) );
  nor_x1_sg U59808 ( .A(n15150), .B(n49716), .X(n15467) );
  nand_x1_sg U59809 ( .A(n15442), .B(n40287), .X(n15469) );
  nor_x1_sg U59810 ( .A(n16288), .B(n40125), .X(n16287) );
  nor_x1_sg U59811 ( .A(n15969), .B(n50003), .X(n16286) );
  nand_x1_sg U59812 ( .A(n16261), .B(n40295), .X(n16288) );
  nor_x1_sg U59813 ( .A(n17926), .B(n40132), .X(n17925) );
  nor_x1_sg U59814 ( .A(n17607), .B(n50577), .X(n17924) );
  nand_x1_sg U59815 ( .A(n17899), .B(n40240), .X(n17926) );
  nor_x1_sg U59816 ( .A(n18747), .B(n40127), .X(n18746) );
  nor_x1_sg U59817 ( .A(n18428), .B(n50864), .X(n18745) );
  nand_x1_sg U59818 ( .A(n18720), .B(n40299), .X(n18747) );
  nor_x1_sg U59819 ( .A(n46870), .B(n46863), .X(n7084) );
  nor_x1_sg U59820 ( .A(n7086), .B(n7087), .X(n7085) );
  inv_x1_sg U59821 ( .A(n7086), .X(n46870) );
  nor_x1_sg U59822 ( .A(n47163), .B(n47156), .X(n7902) );
  nor_x1_sg U59823 ( .A(n7904), .B(n7905), .X(n7903) );
  inv_x1_sg U59824 ( .A(n7904), .X(n47163) );
  nor_x1_sg U59825 ( .A(n47448), .B(n47441), .X(n8720) );
  nor_x1_sg U59826 ( .A(n8722), .B(n8723), .X(n8721) );
  inv_x1_sg U59827 ( .A(n8722), .X(n47448) );
  nor_x1_sg U59828 ( .A(n47733), .B(n47726), .X(n9540) );
  nor_x1_sg U59829 ( .A(n9542), .B(n9543), .X(n9541) );
  inv_x1_sg U59830 ( .A(n9542), .X(n47733) );
  nor_x1_sg U59831 ( .A(n48018), .B(n48011), .X(n10359) );
  nor_x1_sg U59832 ( .A(n10361), .B(n10362), .X(n10360) );
  inv_x1_sg U59833 ( .A(n10361), .X(n48018) );
  nor_x1_sg U59834 ( .A(n48303), .B(n48296), .X(n11178) );
  nor_x1_sg U59835 ( .A(n11180), .B(n11181), .X(n11179) );
  inv_x1_sg U59836 ( .A(n11180), .X(n48303) );
  nor_x1_sg U59837 ( .A(n48588), .B(n48581), .X(n11997) );
  nor_x1_sg U59838 ( .A(n11999), .B(n12000), .X(n11998) );
  inv_x1_sg U59839 ( .A(n11999), .X(n48588) );
  nor_x1_sg U59840 ( .A(n48874), .B(n48867), .X(n12816) );
  nor_x1_sg U59841 ( .A(n12818), .B(n12819), .X(n12817) );
  inv_x1_sg U59842 ( .A(n12818), .X(n48874) );
  nor_x1_sg U59843 ( .A(n49161), .B(n49154), .X(n13635) );
  nor_x1_sg U59844 ( .A(n13637), .B(n13638), .X(n13636) );
  inv_x1_sg U59845 ( .A(n13637), .X(n49161) );
  nor_x1_sg U59846 ( .A(n49447), .B(n49440), .X(n14454) );
  nor_x1_sg U59847 ( .A(n14456), .B(n14457), .X(n14455) );
  inv_x1_sg U59848 ( .A(n14456), .X(n49447) );
  nor_x1_sg U59849 ( .A(n49732), .B(n49725), .X(n15273) );
  nor_x1_sg U59850 ( .A(n15275), .B(n15276), .X(n15274) );
  inv_x1_sg U59851 ( .A(n15275), .X(n49732) );
  nor_x1_sg U59852 ( .A(n50019), .B(n50012), .X(n16092) );
  nor_x1_sg U59853 ( .A(n16094), .B(n16095), .X(n16093) );
  inv_x1_sg U59854 ( .A(n16094), .X(n50019) );
  nor_x1_sg U59855 ( .A(n50304), .B(n50296), .X(n16910) );
  nor_x1_sg U59856 ( .A(n16912), .B(n16913), .X(n16911) );
  inv_x1_sg U59857 ( .A(n16912), .X(n50304) );
  nor_x1_sg U59858 ( .A(n50593), .B(n50586), .X(n17730) );
  nor_x1_sg U59859 ( .A(n17732), .B(n17733), .X(n17731) );
  inv_x1_sg U59860 ( .A(n17732), .X(n50593) );
  nor_x1_sg U59861 ( .A(n50880), .B(n50873), .X(n18551) );
  nor_x1_sg U59862 ( .A(n18553), .B(n18554), .X(n18552) );
  inv_x1_sg U59863 ( .A(n18553), .X(n50880) );
  nor_x1_sg U59864 ( .A(n46845), .B(n40164), .X(n22604) );
  nor_x1_sg U59865 ( .A(n47136), .B(n40243), .X(n22866) );
  nor_x1_sg U59866 ( .A(n47421), .B(n40247), .X(n23143) );
  nor_x1_sg U59867 ( .A(n47706), .B(n40252), .X(n23423) );
  nor_x1_sg U59868 ( .A(n47991), .B(n40257), .X(n23702) );
  nor_x1_sg U59869 ( .A(n48276), .B(n40262), .X(n23981) );
  nor_x1_sg U59870 ( .A(n48561), .B(n40267), .X(n24260) );
  nor_x1_sg U59871 ( .A(n48846), .B(n40272), .X(n24539) );
  nor_x1_sg U59872 ( .A(n49133), .B(n40277), .X(n24817) );
  nor_x1_sg U59873 ( .A(n49419), .B(n40282), .X(n25096) );
  nor_x1_sg U59874 ( .A(n49705), .B(n40287), .X(n25375) );
  nor_x1_sg U59875 ( .A(n49991), .B(n40292), .X(n25654) );
  nor_x1_sg U59876 ( .A(n50852), .B(n40297), .X(n26491) );
  nor_x1_sg U59877 ( .A(n50566), .B(n40238), .X(n26196) );
  nor_x1_sg U59878 ( .A(n46963), .B(n7300), .X(n22660) );
  nor_x1_sg U59879 ( .A(n46849), .B(n41902), .X(n22610) );
  nor_x1_sg U59880 ( .A(n46982), .B(n39664), .X(n22666) );
  nor_x1_sg U59881 ( .A(n47005), .B(n7445), .X(n22672) );
  nor_x1_sg U59882 ( .A(n47024), .B(n7474), .X(n22678) );
  nor_x1_sg U59883 ( .A(n47054), .B(n6997), .X(n22684) );
  nor_x1_sg U59884 ( .A(n47141), .B(n39813), .X(n22873) );
  nor_x1_sg U59885 ( .A(n47426), .B(n39830), .X(n23150) );
  nor_x1_sg U59886 ( .A(n47711), .B(n41878), .X(n23430) );
  nor_x1_sg U59887 ( .A(n47996), .B(n39815), .X(n23709) );
  nor_x1_sg U59888 ( .A(n48281), .B(n39833), .X(n23988) );
  nor_x1_sg U59889 ( .A(n48566), .B(n41884), .X(n24267) );
  nor_x1_sg U59890 ( .A(n48851), .B(n39818), .X(n24546) );
  nor_x1_sg U59891 ( .A(n49138), .B(n39840), .X(n24824) );
  nor_x1_sg U59892 ( .A(n49424), .B(n41880), .X(n25103) );
  nor_x1_sg U59893 ( .A(n49710), .B(n39848), .X(n25382) );
  nor_x1_sg U59894 ( .A(n49996), .B(n41894), .X(n25661) );
  nor_x1_sg U59895 ( .A(n50282), .B(n40608), .X(n25933) );
  nor_x1_sg U59896 ( .A(n50299), .B(n40073), .X(n25945) );
  nor_x1_sg U59897 ( .A(n50571), .B(n41890), .X(n26204) );
  nor_x1_sg U59898 ( .A(n50857), .B(n39824), .X(n26498) );
  nand_x1_sg U59899 ( .A(n22922), .B(n22923), .X(n22921) );
  nand_x1_sg U59900 ( .A(n22925), .B(n39277), .X(n22920) );
  nand_x1_sg U59901 ( .A(n39519), .B(n22924), .X(n22923) );
  nand_x1_sg U59902 ( .A(n22936), .B(n22937), .X(n22935) );
  nand_x1_sg U59903 ( .A(n22939), .B(n41311), .X(n22934) );
  nand_x1_sg U59904 ( .A(n39532), .B(n22938), .X(n22937) );
  nand_x1_sg U59905 ( .A(n22950), .B(n22951), .X(n22949) );
  nand_x1_sg U59906 ( .A(n22953), .B(n38944), .X(n22948) );
  nand_x1_sg U59907 ( .A(n39506), .B(n22952), .X(n22951) );
  nand_x1_sg U59908 ( .A(n22976), .B(n47418), .X(n22975) );
  nand_x1_sg U59909 ( .A(n22981), .B(n39279), .X(n22974) );
  inv_x1_sg U59910 ( .A(n22977), .X(n47418) );
  nand_x1_sg U59911 ( .A(n23199), .B(n23200), .X(n23198) );
  nand_x1_sg U59912 ( .A(n23202), .B(n39657), .X(n23197) );
  nand_x1_sg U59913 ( .A(n42344), .B(n23201), .X(n23200) );
  nand_x1_sg U59914 ( .A(n23213), .B(n23214), .X(n23212) );
  nand_x1_sg U59915 ( .A(n23216), .B(n39475), .X(n23211) );
  nand_x1_sg U59916 ( .A(n39533), .B(n23215), .X(n23214) );
  nand_x1_sg U59917 ( .A(n23227), .B(n23228), .X(n23226) );
  nand_x1_sg U59918 ( .A(n23230), .B(n40224), .X(n23225) );
  nand_x1_sg U59919 ( .A(n39505), .B(n23229), .X(n23228) );
  nand_x1_sg U59920 ( .A(n23479), .B(n23480), .X(n23478) );
  nand_x1_sg U59921 ( .A(n23482), .B(n41309), .X(n23477) );
  nand_x1_sg U59922 ( .A(n42355), .B(n23481), .X(n23480) );
  nand_x1_sg U59923 ( .A(n23493), .B(n23494), .X(n23492) );
  nand_x1_sg U59924 ( .A(n23496), .B(n38943), .X(n23491) );
  nand_x1_sg U59925 ( .A(n39534), .B(n23495), .X(n23494) );
  nand_x1_sg U59926 ( .A(n23507), .B(n23508), .X(n23506) );
  nand_x1_sg U59927 ( .A(n23510), .B(n39926), .X(n23505) );
  nand_x1_sg U59928 ( .A(n39507), .B(n23509), .X(n23508) );
  nand_x1_sg U59929 ( .A(n23533), .B(n47988), .X(n23532) );
  nand_x1_sg U59930 ( .A(n23538), .B(n41464), .X(n23531) );
  inv_x1_sg U59931 ( .A(n23534), .X(n47988) );
  nand_x1_sg U59932 ( .A(n23758), .B(n23759), .X(n23757) );
  nand_x1_sg U59933 ( .A(n23761), .B(n39476), .X(n23756) );
  nand_x1_sg U59934 ( .A(n39523), .B(n23760), .X(n23759) );
  nand_x1_sg U59935 ( .A(n23772), .B(n23773), .X(n23771) );
  nand_x1_sg U59936 ( .A(n23775), .B(n41315), .X(n23770) );
  nand_x1_sg U59937 ( .A(n39535), .B(n23774), .X(n23773) );
  nand_x1_sg U59938 ( .A(n23786), .B(n23787), .X(n23785) );
  nand_x1_sg U59939 ( .A(n23789), .B(n41461), .X(n23784) );
  nand_x1_sg U59940 ( .A(n39509), .B(n23788), .X(n23787) );
  nand_x1_sg U59941 ( .A(n23812), .B(n48273), .X(n23811) );
  nand_x1_sg U59942 ( .A(n23817), .B(n39281), .X(n23810) );
  inv_x1_sg U59943 ( .A(n23813), .X(n48273) );
  nand_x1_sg U59944 ( .A(n24037), .B(n24038), .X(n24036) );
  nand_x1_sg U59945 ( .A(n24040), .B(n41315), .X(n24035) );
  nand_x1_sg U59946 ( .A(n39522), .B(n24039), .X(n24038) );
  nand_x1_sg U59947 ( .A(n24051), .B(n24052), .X(n24050) );
  nand_x1_sg U59948 ( .A(n24054), .B(n39657), .X(n24049) );
  nand_x1_sg U59949 ( .A(n39536), .B(n24053), .X(n24052) );
  nand_x1_sg U59950 ( .A(n24065), .B(n24066), .X(n24064) );
  nand_x1_sg U59951 ( .A(n24068), .B(n40224), .X(n24063) );
  nand_x1_sg U59952 ( .A(n39508), .B(n24067), .X(n24066) );
  nand_x1_sg U59953 ( .A(n24091), .B(n48558), .X(n24090) );
  nand_x1_sg U59954 ( .A(n24096), .B(n40227), .X(n24089) );
  inv_x1_sg U59955 ( .A(n24092), .X(n48558) );
  nand_x1_sg U59956 ( .A(n24316), .B(n24317), .X(n24315) );
  nand_x1_sg U59957 ( .A(n24319), .B(n41463), .X(n24314) );
  nand_x1_sg U59958 ( .A(n42352), .B(n24318), .X(n24317) );
  nand_x1_sg U59959 ( .A(n24330), .B(n24331), .X(n24329) );
  nand_x1_sg U59960 ( .A(n24333), .B(n41462), .X(n24328) );
  nand_x1_sg U59961 ( .A(n39537), .B(n24332), .X(n24331) );
  nand_x1_sg U59962 ( .A(n24344), .B(n24345), .X(n24343) );
  nand_x1_sg U59963 ( .A(n24347), .B(n39278), .X(n24342) );
  nand_x1_sg U59964 ( .A(n39511), .B(n24346), .X(n24345) );
  nand_x1_sg U59965 ( .A(n24370), .B(n48843), .X(n24369) );
  nand_x1_sg U59966 ( .A(n24375), .B(n41313), .X(n24368) );
  inv_x1_sg U59967 ( .A(n24371), .X(n48843) );
  nand_x1_sg U59968 ( .A(n24595), .B(n24596), .X(n24594) );
  nand_x1_sg U59969 ( .A(n24598), .B(n40225), .X(n24593) );
  nand_x1_sg U59970 ( .A(n42351), .B(n24597), .X(n24596) );
  nand_x1_sg U59971 ( .A(n24609), .B(n24610), .X(n24608) );
  nand_x1_sg U59972 ( .A(n24612), .B(n39277), .X(n24607) );
  nand_x1_sg U59973 ( .A(n39538), .B(n24611), .X(n24610) );
  nand_x1_sg U59974 ( .A(n24623), .B(n24624), .X(n24622) );
  nand_x1_sg U59975 ( .A(n24626), .B(n40218), .X(n24621) );
  nand_x1_sg U59976 ( .A(n39510), .B(n24625), .X(n24624) );
  nand_x1_sg U59977 ( .A(n24649), .B(n49130), .X(n24648) );
  nand_x1_sg U59978 ( .A(n24654), .B(n39281), .X(n24647) );
  inv_x1_sg U59979 ( .A(n24650), .X(n49130) );
  nand_x1_sg U59980 ( .A(n24873), .B(n24874), .X(n24872) );
  nand_x1_sg U59981 ( .A(n24876), .B(n41309), .X(n24871) );
  nand_x1_sg U59982 ( .A(n39527), .B(n24875), .X(n24874) );
  nand_x1_sg U59983 ( .A(n24887), .B(n24888), .X(n24886) );
  nand_x1_sg U59984 ( .A(n24890), .B(n39929), .X(n24885) );
  nand_x1_sg U59985 ( .A(n39539), .B(n24889), .X(n24888) );
  nand_x1_sg U59986 ( .A(n24901), .B(n24902), .X(n24900) );
  nand_x1_sg U59987 ( .A(n24904), .B(n40226), .X(n24899) );
  nand_x1_sg U59988 ( .A(n39513), .B(n24903), .X(n24902) );
  nand_x1_sg U59989 ( .A(n24927), .B(n49416), .X(n24926) );
  nand_x1_sg U59990 ( .A(n24932), .B(n39478), .X(n24925) );
  inv_x1_sg U59991 ( .A(n24928), .X(n49416) );
  nand_x1_sg U59992 ( .A(n25152), .B(n25153), .X(n25151) );
  nand_x1_sg U59993 ( .A(n25155), .B(n41317), .X(n25150) );
  nand_x1_sg U59994 ( .A(n39526), .B(n25154), .X(n25153) );
  nand_x1_sg U59995 ( .A(n25166), .B(n25167), .X(n25165) );
  nand_x1_sg U59996 ( .A(n25169), .B(n39478), .X(n25164) );
  nand_x1_sg U59997 ( .A(n39540), .B(n25168), .X(n25167) );
  nand_x1_sg U59998 ( .A(n25180), .B(n25181), .X(n25179) );
  nand_x1_sg U59999 ( .A(n25183), .B(n39476), .X(n25178) );
  nand_x1_sg U60000 ( .A(n39512), .B(n25182), .X(n25181) );
  nand_x1_sg U60001 ( .A(n25206), .B(n49702), .X(n25205) );
  nand_x1_sg U60002 ( .A(n25211), .B(n41317), .X(n25204) );
  inv_x1_sg U60003 ( .A(n25207), .X(n49702) );
  nand_x1_sg U60004 ( .A(n25431), .B(n25432), .X(n25430) );
  nand_x1_sg U60005 ( .A(n25434), .B(n41461), .X(n25429) );
  nand_x1_sg U60006 ( .A(n42348), .B(n25433), .X(n25432) );
  nand_x1_sg U60007 ( .A(n25445), .B(n25446), .X(n25444) );
  nand_x1_sg U60008 ( .A(n25448), .B(n39476), .X(n25443) );
  nand_x1_sg U60009 ( .A(n39541), .B(n25447), .X(n25446) );
  nand_x1_sg U60010 ( .A(n25459), .B(n25460), .X(n25458) );
  nand_x1_sg U60011 ( .A(n25462), .B(n39928), .X(n25457) );
  nand_x1_sg U60012 ( .A(n39515), .B(n25461), .X(n25460) );
  nand_x1_sg U60013 ( .A(n25485), .B(n49988), .X(n25484) );
  nand_x1_sg U60014 ( .A(n25490), .B(n39475), .X(n25483) );
  inv_x1_sg U60015 ( .A(n25486), .X(n49988) );
  nand_x1_sg U60016 ( .A(n25710), .B(n25711), .X(n25709) );
  nand_x1_sg U60017 ( .A(n25713), .B(n41462), .X(n25708) );
  nand_x1_sg U60018 ( .A(n42347), .B(n25712), .X(n25711) );
  nand_x1_sg U60019 ( .A(n25724), .B(n25725), .X(n25723) );
  nand_x1_sg U60020 ( .A(n25727), .B(n39926), .X(n25722) );
  nand_x1_sg U60021 ( .A(n39542), .B(n25726), .X(n25725) );
  nand_x1_sg U60022 ( .A(n25738), .B(n25739), .X(n25737) );
  nand_x1_sg U60023 ( .A(n25741), .B(n39278), .X(n25736) );
  nand_x1_sg U60024 ( .A(n39514), .B(n25740), .X(n25739) );
  nand_x1_sg U60025 ( .A(n25764), .B(n50274), .X(n25763) );
  nand_x1_sg U60026 ( .A(n25769), .B(n39278), .X(n25762) );
  inv_x1_sg U60027 ( .A(n25765), .X(n50274) );
  nand_x1_sg U60028 ( .A(n26547), .B(n26548), .X(n26546) );
  nand_x1_sg U60029 ( .A(n26550), .B(n41313), .X(n26545) );
  nand_x1_sg U60030 ( .A(n39529), .B(n26549), .X(n26548) );
  nand_x1_sg U60031 ( .A(n26561), .B(n26562), .X(n26560) );
  nand_x1_sg U60032 ( .A(n26564), .B(n39926), .X(n26559) );
  nand_x1_sg U60033 ( .A(n39544), .B(n26563), .X(n26562) );
  nand_x1_sg U60034 ( .A(n26575), .B(n26576), .X(n26574) );
  nand_x1_sg U60035 ( .A(n26578), .B(n39928), .X(n26573) );
  nand_x1_sg U60036 ( .A(n39517), .B(n26577), .X(n26576) );
  nand_x1_sg U60037 ( .A(n26601), .B(n51135), .X(n26600) );
  nand_x1_sg U60038 ( .A(n26606), .B(n39281), .X(n26599) );
  inv_x1_sg U60039 ( .A(n26602), .X(n51135) );
  nor_x1_sg U60040 ( .A(n39605), .B(n40085), .X(n7566) );
  nor_x1_sg U60041 ( .A(n39603), .B(n40088), .X(n17391) );
  nor_x1_sg U60042 ( .A(n39548), .B(n41750), .X(n8249) );
  nor_x1_sg U60043 ( .A(n39549), .B(n41742), .X(n9067) );
  nor_x1_sg U60044 ( .A(n39550), .B(n40206), .X(n9887) );
  nor_x1_sg U60045 ( .A(n39557), .B(n41744), .X(n10706) );
  nor_x1_sg U60046 ( .A(n39558), .B(n40198), .X(n11525) );
  nor_x1_sg U60047 ( .A(n39554), .B(n40194), .X(n12344) );
  nor_x1_sg U60048 ( .A(n39555), .B(n40192), .X(n13163) );
  nor_x1_sg U60049 ( .A(n39556), .B(n40176), .X(n13982) );
  nor_x1_sg U60050 ( .A(n39553), .B(n40188), .X(n14801) );
  nor_x1_sg U60051 ( .A(n39551), .B(n40170), .X(n15620) );
  nor_x1_sg U60052 ( .A(n39552), .B(n41753), .X(n16439) );
  nor_x1_sg U60053 ( .A(n41739), .B(n40087), .X(n17256) );
  nor_x1_sg U60054 ( .A(n39546), .B(n41741), .X(n18077) );
  nor_x1_sg U60055 ( .A(n39547), .B(n40182), .X(n18898) );
  nor_x1_sg U60056 ( .A(n41736), .B(n40308), .X(n8075) );
  nor_x1_sg U60057 ( .A(n39549), .B(n41843), .X(n8893) );
  nor_x1_sg U60058 ( .A(n41734), .B(n41756), .X(n9713) );
  nor_x1_sg U60059 ( .A(n39557), .B(n41854), .X(n10532) );
  nor_x1_sg U60060 ( .A(n41726), .B(n41758), .X(n11351) );
  nor_x1_sg U60061 ( .A(n39554), .B(n41856), .X(n12170) );
  nor_x1_sg U60062 ( .A(n41729), .B(n41858), .X(n12989) );
  nor_x1_sg U60063 ( .A(n39556), .B(n41761), .X(n13808) );
  nor_x1_sg U60064 ( .A(n41731), .B(n41837), .X(n14627) );
  nor_x1_sg U60065 ( .A(n39551), .B(n41845), .X(n15446) );
  nor_x1_sg U60066 ( .A(n39552), .B(n41839), .X(n16265) );
  nor_x1_sg U60067 ( .A(n39545), .B(n40311), .X(n17081) );
  nor_x1_sg U60068 ( .A(n39546), .B(n40365), .X(n17903) );
  nor_x1_sg U60069 ( .A(n41737), .B(n41841), .X(n18724) );
  nor_x1_sg U60070 ( .A(n41780), .B(n39605), .X(n7586) );
  nor_x1_sg U60071 ( .A(n41782), .B(n39730), .X(n8404) );
  nor_x1_sg U60072 ( .A(n39717), .B(n39734), .X(n9222) );
  nor_x1_sg U60073 ( .A(n41786), .B(n39737), .X(n10042) );
  nor_x1_sg U60074 ( .A(n41788), .B(n39739), .X(n10861) );
  nor_x1_sg U60075 ( .A(n41790), .B(n39743), .X(n11680) );
  nor_x1_sg U60076 ( .A(n41792), .B(n39745), .X(n12499) );
  nor_x1_sg U60077 ( .A(n41794), .B(n39749), .X(n13318) );
  nor_x1_sg U60078 ( .A(n39698), .B(n39752), .X(n14137) );
  nor_x1_sg U60079 ( .A(n39696), .B(n39754), .X(n14956) );
  nor_x1_sg U60080 ( .A(n41800), .B(n39758), .X(n15775) );
  nor_x1_sg U60081 ( .A(n41802), .B(n39760), .X(n16594) );
  nor_x1_sg U60082 ( .A(n39686), .B(n39763), .X(n18232) );
  nor_x1_sg U60083 ( .A(n41806), .B(n39767), .X(n19053) );
  nor_x1_sg U60084 ( .A(n39723), .B(n41691), .X(n7604) );
  nor_x1_sg U60085 ( .A(n39719), .B(n39894), .X(n8422) );
  nor_x1_sg U60086 ( .A(n41784), .B(n39860), .X(n9240) );
  nor_x1_sg U60087 ( .A(n39713), .B(n39858), .X(n10060) );
  nor_x1_sg U60088 ( .A(n39711), .B(n39864), .X(n10879) );
  nor_x1_sg U60089 ( .A(n39708), .B(n39867), .X(n11698) );
  nor_x1_sg U60090 ( .A(n39705), .B(n39870), .X(n12517) );
  nor_x1_sg U60091 ( .A(n39701), .B(n39873), .X(n13336) );
  nor_x1_sg U60092 ( .A(n39699), .B(n39876), .X(n14155) );
  nor_x1_sg U60093 ( .A(n41798), .B(n39879), .X(n14974) );
  nor_x1_sg U60094 ( .A(n39692), .B(n39896), .X(n15793) );
  nor_x1_sg U60095 ( .A(n39689), .B(n39882), .X(n16612) );
  nor_x1_sg U60096 ( .A(n41804), .B(n39887), .X(n18250) );
  nor_x1_sg U60097 ( .A(n39683), .B(n39891), .X(n19071) );
  nor_x1_sg U60098 ( .A(n39723), .B(n41710), .X(n7021) );
  nor_x1_sg U60099 ( .A(n39720), .B(n41712), .X(n7839) );
  nor_x1_sg U60100 ( .A(n41784), .B(n41711), .X(n8657) );
  nor_x1_sg U60101 ( .A(n39714), .B(n41714), .X(n9477) );
  nor_x1_sg U60102 ( .A(n41788), .B(n41713), .X(n10296) );
  nor_x1_sg U60103 ( .A(n39707), .B(n41716), .X(n11115) );
  nor_x1_sg U60104 ( .A(n39705), .B(n41715), .X(n11934) );
  nor_x1_sg U60105 ( .A(n39702), .B(n41718), .X(n12753) );
  nor_x1_sg U60106 ( .A(n39699), .B(n41717), .X(n13572) );
  nor_x1_sg U60107 ( .A(n41798), .B(n41720), .X(n14391) );
  nor_x1_sg U60108 ( .A(n39693), .B(n41719), .X(n15210) );
  nor_x1_sg U60109 ( .A(n39690), .B(n41722), .X(n16029) );
  nor_x1_sg U60110 ( .A(n41804), .B(n41721), .X(n17667) );
  nor_x1_sg U60111 ( .A(n39684), .B(n41723), .X(n18488) );
  nor_x1_sg U60112 ( .A(n39611), .B(n7651), .X(n8186) );
  nor_x1_sg U60113 ( .A(n39612), .B(n40178), .X(n8308) );
  nor_x1_sg U60114 ( .A(n39608), .B(n40557), .X(n9004) );
  nor_x1_sg U60115 ( .A(n39609), .B(n40210), .X(n9126) );
  nor_x1_sg U60116 ( .A(n39626), .B(n40553), .X(n9824) );
  nor_x1_sg U60117 ( .A(n39626), .B(n41743), .X(n9946) );
  nor_x1_sg U60118 ( .A(n39623), .B(n10108), .X(n10643) );
  nor_x1_sg U60119 ( .A(n39623), .B(n40202), .X(n10765) );
  nor_x1_sg U60120 ( .A(n39620), .B(n40543), .X(n11462) );
  nor_x1_sg U60121 ( .A(n39620), .B(n41745), .X(n11584) );
  nor_x1_sg U60122 ( .A(n39617), .B(n11746), .X(n12281) );
  nor_x1_sg U60123 ( .A(n39617), .B(n41746), .X(n12403) );
  nor_x1_sg U60124 ( .A(n39638), .B(n40537), .X(n13100) );
  nor_x1_sg U60125 ( .A(n39638), .B(n41747), .X(n13222) );
  nor_x1_sg U60126 ( .A(n39636), .B(n40532), .X(n13919) );
  nor_x1_sg U60127 ( .A(n39635), .B(n40176), .X(n14041) );
  nor_x1_sg U60128 ( .A(n39632), .B(n40529), .X(n14738) );
  nor_x1_sg U60129 ( .A(n39632), .B(n41748), .X(n14860) );
  nor_x1_sg U60130 ( .A(n39629), .B(n40523), .X(n15557) );
  nor_x1_sg U60131 ( .A(n39630), .B(n41752), .X(n15679) );
  nor_x1_sg U60132 ( .A(n39647), .B(n40519), .X(n16376) );
  nor_x1_sg U60133 ( .A(n39647), .B(n40166), .X(n16498) );
  nor_x1_sg U60134 ( .A(n39614), .B(n40303), .X(n17193) );
  nor_x1_sg U60135 ( .A(n39614), .B(n40087), .X(n17315) );
  nor_x1_sg U60136 ( .A(n39644), .B(n40515), .X(n18014) );
  nor_x1_sg U60137 ( .A(n39645), .B(n40214), .X(n18136) );
  nor_x1_sg U60138 ( .A(n39642), .B(n18300), .X(n18835) );
  nor_x1_sg U60139 ( .A(n39641), .B(n41749), .X(n18957) );
  nor_x1_sg U60140 ( .A(n39611), .B(n40306), .X(n8120) );
  nor_x1_sg U60141 ( .A(n39609), .B(n41754), .X(n8938) );
  nor_x1_sg U60142 ( .A(n39626), .B(n41756), .X(n9758) );
  nor_x1_sg U60143 ( .A(n39623), .B(n41855), .X(n10577) );
  nor_x1_sg U60144 ( .A(n39620), .B(n41758), .X(n11396) );
  nor_x1_sg U60145 ( .A(n39617), .B(n41857), .X(n12215) );
  nor_x1_sg U60146 ( .A(n39638), .B(n41859), .X(n13034) );
  nor_x1_sg U60147 ( .A(n39635), .B(n41761), .X(n13853) );
  nor_x1_sg U60148 ( .A(n39632), .B(n41759), .X(n14672) );
  nor_x1_sg U60149 ( .A(n39629), .B(n41765), .X(n15491) );
  nor_x1_sg U60150 ( .A(n39647), .B(n41764), .X(n16310) );
  nor_x1_sg U60151 ( .A(n39614), .B(n40311), .X(n17127) );
  nor_x1_sg U60152 ( .A(n39644), .B(n40365), .X(n17948) );
  nor_x1_sg U60153 ( .A(n39641), .B(n41762), .X(n18769) );
  nor_x1_sg U60154 ( .A(n6841), .B(n6847), .X(n6845) );
  nor_x1_sg U60155 ( .A(n7658), .B(n7664), .X(n7662) );
  nor_x1_sg U60156 ( .A(n8476), .B(n8482), .X(n8480) );
  nor_x1_sg U60157 ( .A(n9296), .B(n9302), .X(n9300) );
  nor_x1_sg U60158 ( .A(n10115), .B(n10121), .X(n10119) );
  nor_x1_sg U60159 ( .A(n10934), .B(n10940), .X(n10938) );
  nor_x1_sg U60160 ( .A(n11753), .B(n11759), .X(n11757) );
  nor_x1_sg U60161 ( .A(n12572), .B(n12578), .X(n12576) );
  nor_x1_sg U60162 ( .A(n13391), .B(n13397), .X(n13395) );
  nor_x1_sg U60163 ( .A(n14210), .B(n14216), .X(n14214) );
  nor_x1_sg U60164 ( .A(n15029), .B(n15035), .X(n15033) );
  nor_x1_sg U60165 ( .A(n15848), .B(n15854), .X(n15852) );
  nor_x1_sg U60166 ( .A(n17486), .B(n17492), .X(n17490) );
  nor_x1_sg U60167 ( .A(n18307), .B(n18313), .X(n18311) );
  nor_x1_sg U60168 ( .A(n16665), .B(n16671), .X(n16669) );
  nor_x1_sg U60169 ( .A(n7584), .B(n46990), .X(n7582) );
  nor_x1_sg U60170 ( .A(n7587), .B(n7586), .X(n7584) );
  nand_x1_sg U60171 ( .A(n7586), .B(n7587), .X(n7585) );
  nor_x1_sg U60172 ( .A(n8402), .B(n47279), .X(n8400) );
  nor_x1_sg U60173 ( .A(n8405), .B(n8404), .X(n8402) );
  nand_x1_sg U60174 ( .A(n8404), .B(n8405), .X(n8403) );
  nor_x1_sg U60175 ( .A(n9220), .B(n47564), .X(n9218) );
  nor_x1_sg U60176 ( .A(n9223), .B(n9222), .X(n9220) );
  nand_x1_sg U60177 ( .A(n9222), .B(n9223), .X(n9221) );
  nor_x1_sg U60178 ( .A(n10040), .B(n47849), .X(n10038) );
  nor_x1_sg U60179 ( .A(n10043), .B(n10042), .X(n10040) );
  nand_x1_sg U60180 ( .A(n10042), .B(n10043), .X(n10041) );
  nor_x1_sg U60181 ( .A(n10859), .B(n48134), .X(n10857) );
  nor_x1_sg U60182 ( .A(n10862), .B(n10861), .X(n10859) );
  nand_x1_sg U60183 ( .A(n10861), .B(n10862), .X(n10860) );
  nor_x1_sg U60184 ( .A(n11678), .B(n48419), .X(n11676) );
  nor_x1_sg U60185 ( .A(n11681), .B(n11680), .X(n11678) );
  nand_x1_sg U60186 ( .A(n11680), .B(n11681), .X(n11679) );
  nor_x1_sg U60187 ( .A(n12497), .B(n48704), .X(n12495) );
  nor_x1_sg U60188 ( .A(n12500), .B(n12499), .X(n12497) );
  nand_x1_sg U60189 ( .A(n12499), .B(n12500), .X(n12498) );
  nor_x1_sg U60190 ( .A(n13316), .B(n48990), .X(n13314) );
  nor_x1_sg U60191 ( .A(n13319), .B(n13318), .X(n13316) );
  nand_x1_sg U60192 ( .A(n13318), .B(n13319), .X(n13317) );
  nor_x1_sg U60193 ( .A(n14135), .B(n49277), .X(n14133) );
  nor_x1_sg U60194 ( .A(n14138), .B(n14137), .X(n14135) );
  nand_x1_sg U60195 ( .A(n14137), .B(n14138), .X(n14136) );
  nor_x1_sg U60196 ( .A(n14954), .B(n49563), .X(n14952) );
  nor_x1_sg U60197 ( .A(n14957), .B(n14956), .X(n14954) );
  nand_x1_sg U60198 ( .A(n14956), .B(n14957), .X(n14955) );
  nor_x1_sg U60199 ( .A(n15773), .B(n49849), .X(n15771) );
  nor_x1_sg U60200 ( .A(n15776), .B(n15775), .X(n15773) );
  nand_x1_sg U60201 ( .A(n15775), .B(n15776), .X(n15774) );
  nor_x1_sg U60202 ( .A(n16592), .B(n50135), .X(n16590) );
  nor_x1_sg U60203 ( .A(n16595), .B(n16594), .X(n16592) );
  nand_x1_sg U60204 ( .A(n16594), .B(n16595), .X(n16593) );
  nor_x1_sg U60205 ( .A(n18230), .B(n50709), .X(n18228) );
  nor_x1_sg U60206 ( .A(n18233), .B(n18232), .X(n18230) );
  nand_x1_sg U60207 ( .A(n18232), .B(n18233), .X(n18231) );
  nor_x1_sg U60208 ( .A(n19051), .B(n50996), .X(n19049) );
  nor_x1_sg U60209 ( .A(n19054), .B(n19053), .X(n19051) );
  nand_x1_sg U60210 ( .A(n19053), .B(n19054), .X(n19052) );
  nor_x1_sg U60211 ( .A(n7602), .B(n46972), .X(n7600) );
  nor_x1_sg U60212 ( .A(n7605), .B(n7604), .X(n7602) );
  nand_x1_sg U60213 ( .A(n7604), .B(n7605), .X(n7603) );
  nor_x1_sg U60214 ( .A(n8420), .B(n47262), .X(n8418) );
  nor_x1_sg U60215 ( .A(n8423), .B(n8422), .X(n8420) );
  nand_x1_sg U60216 ( .A(n8422), .B(n8423), .X(n8421) );
  nor_x1_sg U60217 ( .A(n9238), .B(n47547), .X(n9236) );
  nor_x1_sg U60218 ( .A(n9241), .B(n9240), .X(n9238) );
  nand_x1_sg U60219 ( .A(n9240), .B(n9241), .X(n9239) );
  nor_x1_sg U60220 ( .A(n10058), .B(n47832), .X(n10056) );
  nor_x1_sg U60221 ( .A(n10061), .B(n10060), .X(n10058) );
  nand_x1_sg U60222 ( .A(n10060), .B(n10061), .X(n10059) );
  nor_x1_sg U60223 ( .A(n10877), .B(n48117), .X(n10875) );
  nor_x1_sg U60224 ( .A(n10880), .B(n10879), .X(n10877) );
  nand_x1_sg U60225 ( .A(n10879), .B(n10880), .X(n10878) );
  nor_x1_sg U60226 ( .A(n11696), .B(n48402), .X(n11694) );
  nor_x1_sg U60227 ( .A(n11699), .B(n11698), .X(n11696) );
  nand_x1_sg U60228 ( .A(n11698), .B(n11699), .X(n11697) );
  nor_x1_sg U60229 ( .A(n12515), .B(n48687), .X(n12513) );
  nor_x1_sg U60230 ( .A(n12518), .B(n12517), .X(n12515) );
  nand_x1_sg U60231 ( .A(n12517), .B(n12518), .X(n12516) );
  nor_x1_sg U60232 ( .A(n13334), .B(n48973), .X(n13332) );
  nor_x1_sg U60233 ( .A(n13337), .B(n13336), .X(n13334) );
  nand_x1_sg U60234 ( .A(n13336), .B(n13337), .X(n13335) );
  nor_x1_sg U60235 ( .A(n14153), .B(n49260), .X(n14151) );
  nor_x1_sg U60236 ( .A(n14156), .B(n14155), .X(n14153) );
  nand_x1_sg U60237 ( .A(n14155), .B(n14156), .X(n14154) );
  nor_x1_sg U60238 ( .A(n14972), .B(n49546), .X(n14970) );
  nor_x1_sg U60239 ( .A(n14975), .B(n14974), .X(n14972) );
  nand_x1_sg U60240 ( .A(n14974), .B(n14975), .X(n14973) );
  nor_x1_sg U60241 ( .A(n15791), .B(n49832), .X(n15789) );
  nor_x1_sg U60242 ( .A(n15794), .B(n15793), .X(n15791) );
  nand_x1_sg U60243 ( .A(n15793), .B(n15794), .X(n15792) );
  nor_x1_sg U60244 ( .A(n16610), .B(n50118), .X(n16608) );
  nor_x1_sg U60245 ( .A(n16613), .B(n16612), .X(n16610) );
  nand_x1_sg U60246 ( .A(n16612), .B(n16613), .X(n16611) );
  nor_x1_sg U60247 ( .A(n18248), .B(n50692), .X(n18246) );
  nor_x1_sg U60248 ( .A(n18251), .B(n18250), .X(n18248) );
  nand_x1_sg U60249 ( .A(n18250), .B(n18251), .X(n18249) );
  nor_x1_sg U60250 ( .A(n19069), .B(n50979), .X(n19067) );
  nor_x1_sg U60251 ( .A(n19072), .B(n19071), .X(n19069) );
  nand_x1_sg U60252 ( .A(n19071), .B(n19072), .X(n19070) );
  nor_x1_sg U60253 ( .A(n17409), .B(n50420), .X(n17407) );
  nor_x1_sg U60254 ( .A(n17412), .B(n17411), .X(n17409) );
  nand_x1_sg U60255 ( .A(n17411), .B(n17412), .X(n17410) );
  nor_x1_sg U60256 ( .A(n17427), .B(n50403), .X(n17425) );
  nor_x1_sg U60257 ( .A(n17430), .B(n17429), .X(n17427) );
  nand_x1_sg U60258 ( .A(n17429), .B(n17430), .X(n17428) );
  nor_x1_sg U60259 ( .A(n40609), .B(n50305), .X(n16908) );
  nor_x1_sg U60260 ( .A(n16909), .B(n39681), .X(n16907) );
  nor_x1_sg U60261 ( .A(n16664), .B(n40304), .X(n16671) );
  nor_x1_sg U60262 ( .A(n6840), .B(n40614), .X(n6847) );
  nor_x1_sg U60263 ( .A(n7657), .B(n40559), .X(n7664) );
  nor_x1_sg U60264 ( .A(n8475), .B(n40556), .X(n8482) );
  nor_x1_sg U60265 ( .A(n9295), .B(n9289), .X(n9302) );
  nor_x1_sg U60266 ( .A(n10114), .B(n40547), .X(n10121) );
  nor_x1_sg U60267 ( .A(n10933), .B(n40544), .X(n10940) );
  nor_x1_sg U60268 ( .A(n11752), .B(n40541), .X(n11759) );
  nor_x1_sg U60269 ( .A(n12571), .B(n40535), .X(n12578) );
  nor_x1_sg U60270 ( .A(n13390), .B(n13384), .X(n13397) );
  nor_x1_sg U60271 ( .A(n14209), .B(n40528), .X(n14216) );
  nor_x1_sg U60272 ( .A(n15028), .B(n40524), .X(n15035) );
  nor_x1_sg U60273 ( .A(n15847), .B(n40520), .X(n15854) );
  nor_x1_sg U60274 ( .A(n17485), .B(n17479), .X(n17492) );
  nor_x1_sg U60275 ( .A(n18306), .B(n40513), .X(n18313) );
  nand_x1_sg U60276 ( .A(n39435), .B(n41125), .X(n19105) );
  nor_x1_sg U60277 ( .A(n40106), .B(n41847), .X(n8033) );
  nor_x1_sg U60278 ( .A(n8035), .B(n40179), .X(n8162) );
  nor_x1_sg U60279 ( .A(n40108), .B(n39069), .X(n8851) );
  nor_x1_sg U60280 ( .A(n40107), .B(n40211), .X(n8980) );
  nor_x1_sg U60281 ( .A(n40109), .B(n41852), .X(n9671) );
  nor_x1_sg U60282 ( .A(n9673), .B(n40208), .X(n9800) );
  nor_x1_sg U60283 ( .A(n40112), .B(n41757), .X(n10490) );
  nor_x1_sg U60284 ( .A(n10492), .B(n40203), .X(n10619) );
  nor_x1_sg U60285 ( .A(n40114), .B(n41850), .X(n11309) );
  nor_x1_sg U60286 ( .A(n40113), .B(n40200), .X(n11438) );
  nor_x1_sg U60287 ( .A(n40115), .B(n41763), .X(n12128) );
  nor_x1_sg U60288 ( .A(n12130), .B(n40196), .X(n12257) );
  nor_x1_sg U60289 ( .A(n40118), .B(n41760), .X(n12947) );
  nor_x1_sg U60290 ( .A(n12949), .B(n40190), .X(n13076) );
  nor_x1_sg U60291 ( .A(n40120), .B(n41848), .X(n13766) );
  nor_x1_sg U60292 ( .A(n40119), .B(n41751), .X(n13895) );
  nor_x1_sg U60293 ( .A(n40121), .B(n41836), .X(n14585) );
  nor_x1_sg U60294 ( .A(n14587), .B(n40186), .X(n14714) );
  nor_x1_sg U60295 ( .A(n40123), .B(n39070), .X(n15404) );
  nor_x1_sg U60296 ( .A(n40123), .B(n40172), .X(n15533) );
  nor_x1_sg U60297 ( .A(n40126), .B(n41838), .X(n16223) );
  nor_x1_sg U60298 ( .A(n40125), .B(n41753), .X(n16352) );
  nor_x1_sg U60299 ( .A(n17041), .B(n39679), .X(n17112) );
  nor_x1_sg U60300 ( .A(n17041), .B(n40311), .X(n17039) );
  nor_x1_sg U60301 ( .A(n40130), .B(n40087), .X(n17169) );
  nor_x1_sg U60302 ( .A(n40131), .B(n40365), .X(n17861) );
  nor_x1_sg U60303 ( .A(n40132), .B(n40216), .X(n17990) );
  nor_x1_sg U60304 ( .A(n40127), .B(n41840), .X(n18682) );
  nor_x1_sg U60305 ( .A(n18684), .B(n40184), .X(n18811) );
  nor_x1_sg U60306 ( .A(n40105), .B(n40561), .X(n8072) );
  nor_x1_sg U60307 ( .A(n8853), .B(n40555), .X(n8890) );
  nor_x1_sg U60308 ( .A(n40109), .B(n40551), .X(n9710) );
  nor_x1_sg U60309 ( .A(n40111), .B(n40549), .X(n10529) );
  nor_x1_sg U60310 ( .A(n11311), .B(n10927), .X(n11348) );
  nor_x1_sg U60311 ( .A(n40115), .B(n40541), .X(n12167) );
  nor_x1_sg U60312 ( .A(n40117), .B(n12565), .X(n12986) );
  nor_x1_sg U60313 ( .A(n40119), .B(n40531), .X(n13805) );
  nor_x1_sg U60314 ( .A(n40121), .B(n40527), .X(n14624) );
  nor_x1_sg U60315 ( .A(n15406), .B(n40525), .X(n15443) );
  nor_x1_sg U60316 ( .A(n16225), .B(n15841), .X(n16262) );
  nor_x1_sg U60317 ( .A(n40130), .B(n40302), .X(n17078) );
  nor_x1_sg U60318 ( .A(n17863), .B(n40517), .X(n17900) );
  nor_x1_sg U60319 ( .A(n40127), .B(n40513), .X(n18721) );
  nor_x1_sg U60320 ( .A(n41725), .B(n40615), .X(n7368) );
  nor_x1_sg U60321 ( .A(n39204), .B(n40084), .X(n7490) );
  nor_x1_sg U60322 ( .A(n39204), .B(n41903), .X(n7302) );
  nand_x1_sg U60323 ( .A(n38984), .B(n51181), .X(n10913) );
  nor_x1_sg U60324 ( .A(n46921), .B(n6996), .X(n7250) );
  nor_x1_sg U60325 ( .A(n50354), .B(n39317), .X(n17075) );
  nor_x1_sg U60326 ( .A(n47213), .B(n7813), .X(n8069) );
  nor_x1_sg U60327 ( .A(n47498), .B(n8631), .X(n8887) );
  nor_x1_sg U60328 ( .A(n47783), .B(n9451), .X(n9707) );
  nor_x1_sg U60329 ( .A(n48068), .B(n10270), .X(n10526) );
  nor_x1_sg U60330 ( .A(n48353), .B(n11089), .X(n11345) );
  nor_x1_sg U60331 ( .A(n48638), .B(n11908), .X(n12164) );
  nor_x1_sg U60332 ( .A(n48924), .B(n39304), .X(n12983) );
  nor_x1_sg U60333 ( .A(n49211), .B(n39302), .X(n13802) );
  nor_x1_sg U60334 ( .A(n49497), .B(n39300), .X(n14621) );
  nor_x1_sg U60335 ( .A(n49783), .B(n15184), .X(n15440) );
  nor_x1_sg U60336 ( .A(n50069), .B(n16003), .X(n16259) );
  nor_x1_sg U60337 ( .A(n50643), .B(n17641), .X(n17897) );
  nor_x1_sg U60338 ( .A(n50930), .B(n39294), .X(n18718) );
  nor_x1_sg U60339 ( .A(n39930), .B(n40368), .X(n7214) );
  nor_x1_sg U60340 ( .A(n39930), .B(n41779), .X(n7344) );
  nor_x1_sg U60341 ( .A(n39931), .B(n40614), .X(n7253) );
  nor_x1_sg U60342 ( .A(n46986), .B(n7363), .X(n7357) );
  nor_x1_sg U60343 ( .A(n7364), .B(n42163), .X(n7363) );
  nand_x1_sg U60344 ( .A(n7371), .B(n7283), .X(n7370) );
  nor_x1_sg U60345 ( .A(n47275), .B(n8181), .X(n8175) );
  nor_x1_sg U60346 ( .A(n8182), .B(n40106), .X(n8181) );
  nand_x1_sg U60347 ( .A(n8189), .B(n8102), .X(n8188) );
  nor_x1_sg U60348 ( .A(n47560), .B(n8999), .X(n8993) );
  nor_x1_sg U60349 ( .A(n9000), .B(n8853), .X(n8999) );
  nand_x1_sg U60350 ( .A(n9007), .B(n8920), .X(n9006) );
  nor_x1_sg U60351 ( .A(n47845), .B(n9819), .X(n9813) );
  nor_x1_sg U60352 ( .A(n9820), .B(n9673), .X(n9819) );
  nand_x1_sg U60353 ( .A(n9827), .B(n9740), .X(n9826) );
  nor_x1_sg U60354 ( .A(n48130), .B(n10638), .X(n10632) );
  nor_x1_sg U60355 ( .A(n10639), .B(n10492), .X(n10638) );
  nand_x1_sg U60356 ( .A(n10646), .B(n10559), .X(n10645) );
  nor_x1_sg U60357 ( .A(n48415), .B(n11457), .X(n11451) );
  nor_x1_sg U60358 ( .A(n11458), .B(n11311), .X(n11457) );
  nand_x1_sg U60359 ( .A(n11465), .B(n11378), .X(n11464) );
  nor_x1_sg U60360 ( .A(n48700), .B(n12276), .X(n12270) );
  nor_x1_sg U60361 ( .A(n12277), .B(n12130), .X(n12276) );
  nand_x1_sg U60362 ( .A(n12284), .B(n12197), .X(n12283) );
  nor_x1_sg U60363 ( .A(n48986), .B(n13095), .X(n13089) );
  nor_x1_sg U60364 ( .A(n13096), .B(n12949), .X(n13095) );
  nand_x1_sg U60365 ( .A(n13103), .B(n13016), .X(n13102) );
  nor_x1_sg U60366 ( .A(n49273), .B(n13914), .X(n13908) );
  nor_x1_sg U60367 ( .A(n13915), .B(n13768), .X(n13914) );
  nand_x1_sg U60368 ( .A(n13922), .B(n13835), .X(n13921) );
  nor_x1_sg U60369 ( .A(n49559), .B(n14733), .X(n14727) );
  nor_x1_sg U60370 ( .A(n14734), .B(n14587), .X(n14733) );
  nand_x1_sg U60371 ( .A(n14741), .B(n14654), .X(n14740) );
  nor_x1_sg U60372 ( .A(n49845), .B(n15552), .X(n15546) );
  nor_x1_sg U60373 ( .A(n15553), .B(n15406), .X(n15552) );
  nand_x1_sg U60374 ( .A(n15560), .B(n15473), .X(n15559) );
  nor_x1_sg U60375 ( .A(n50131), .B(n16371), .X(n16365) );
  nor_x1_sg U60376 ( .A(n16372), .B(n16225), .X(n16371) );
  nand_x1_sg U60377 ( .A(n16379), .B(n16292), .X(n16378) );
  nor_x1_sg U60378 ( .A(n50416), .B(n17188), .X(n17182) );
  nor_x1_sg U60379 ( .A(n17189), .B(n17041), .X(n17188) );
  nand_x1_sg U60380 ( .A(n17196), .B(n17108), .X(n17195) );
  nor_x1_sg U60381 ( .A(n50705), .B(n18009), .X(n18003) );
  nor_x1_sg U60382 ( .A(n18010), .B(n17863), .X(n18009) );
  nand_x1_sg U60383 ( .A(n18017), .B(n17930), .X(n18016) );
  nor_x1_sg U60384 ( .A(n50992), .B(n18830), .X(n18824) );
  nor_x1_sg U60385 ( .A(n18831), .B(n18684), .X(n18830) );
  nand_x1_sg U60386 ( .A(n18838), .B(n18751), .X(n18837) );
  nor_x1_sg U60387 ( .A(n39855), .B(n40369), .X(n7380) );
  nor_x1_sg U60388 ( .A(n41664), .B(n40306), .X(n8198) );
  nor_x1_sg U60389 ( .A(n39860), .B(n41754), .X(n9016) );
  nor_x1_sg U60390 ( .A(n39857), .B(n41853), .X(n9836) );
  nor_x1_sg U60391 ( .A(n39863), .B(n41854), .X(n10655) );
  nor_x1_sg U60392 ( .A(n39866), .B(n41851), .X(n11474) );
  nor_x1_sg U60393 ( .A(n39869), .B(n41856), .X(n12293) );
  nor_x1_sg U60394 ( .A(n39872), .B(n41858), .X(n13112) );
  nor_x1_sg U60395 ( .A(n39875), .B(n41849), .X(n13931) );
  nor_x1_sg U60396 ( .A(n39878), .B(n41759), .X(n14750) );
  nor_x1_sg U60397 ( .A(n41662), .B(n41846), .X(n15569) );
  nor_x1_sg U60398 ( .A(n39881), .B(n41764), .X(n16388) );
  nor_x1_sg U60399 ( .A(n41671), .B(n40312), .X(n17205) );
  nor_x1_sg U60400 ( .A(n41669), .B(n40364), .X(n18026) );
  nor_x1_sg U60401 ( .A(n39890), .B(n41762), .X(n18847) );
  nor_x1_sg U60402 ( .A(n39078), .B(n40369), .X(n7156) );
  nor_x1_sg U60403 ( .A(n39077), .B(n40310), .X(n16981) );
  nor_x1_sg U60404 ( .A(n39037), .B(n40369), .X(n7611) );
  nor_x1_sg U60405 ( .A(n41629), .B(n41847), .X(n8429) );
  nor_x1_sg U60406 ( .A(n41630), .B(n41844), .X(n9247) );
  nor_x1_sg U60407 ( .A(n41628), .B(n39073), .X(n10067) );
  nor_x1_sg U60408 ( .A(n41626), .B(n39074), .X(n10886) );
  nor_x1_sg U60409 ( .A(n41627), .B(n39072), .X(n11705) );
  nor_x1_sg U60410 ( .A(n41625), .B(n39075), .X(n12524) );
  nor_x1_sg U60411 ( .A(n49055), .B(n39076), .X(n13343) );
  nor_x1_sg U60412 ( .A(n41624), .B(n39071), .X(n14162) );
  nor_x1_sg U60413 ( .A(n41623), .B(n41836), .X(n14981) );
  nor_x1_sg U60414 ( .A(n41621), .B(n41845), .X(n15800) );
  nor_x1_sg U60415 ( .A(n41622), .B(n41838), .X(n16619) );
  nor_x1_sg U60416 ( .A(n41618), .B(n41842), .X(n17436) );
  nor_x1_sg U60417 ( .A(n41619), .B(n50565), .X(n18257) );
  nor_x1_sg U60418 ( .A(n41620), .B(n41840), .X(n19078) );
  nor_x1_sg U60419 ( .A(n41631), .B(n40615), .X(n7637) );
  nor_x1_sg U60420 ( .A(n41629), .B(n7651), .X(n8455) );
  nor_x1_sg U60421 ( .A(n41630), .B(n40556), .X(n9273) );
  nor_x1_sg U60422 ( .A(n41628), .B(n9289), .X(n10093) );
  nor_x1_sg U60423 ( .A(n41626), .B(n40547), .X(n10912) );
  nor_x1_sg U60424 ( .A(n41627), .B(n40544), .X(n11731) );
  nor_x1_sg U60425 ( .A(n41625), .B(n40541), .X(n12550) );
  nor_x1_sg U60426 ( .A(n49055), .B(n40536), .X(n13369) );
  nor_x1_sg U60427 ( .A(n41624), .B(n40532), .X(n14188) );
  nor_x1_sg U60428 ( .A(n41623), .B(n40528), .X(n15007) );
  nor_x1_sg U60429 ( .A(n41621), .B(n15022), .X(n15826) );
  nor_x1_sg U60430 ( .A(n41622), .B(n40520), .X(n16645) );
  nor_x1_sg U60431 ( .A(n39024), .B(n40301), .X(n17462) );
  nor_x1_sg U60432 ( .A(n41619), .B(n17479), .X(n18283) );
  nor_x1_sg U60433 ( .A(n41620), .B(n40513), .X(n19104) );
  nor_x1_sg U60434 ( .A(n41578), .B(n40178), .X(n7819) );
  nor_x1_sg U60435 ( .A(n41577), .B(n40210), .X(n8637) );
  nor_x1_sg U60436 ( .A(n41576), .B(n41743), .X(n9457) );
  nor_x1_sg U60437 ( .A(n41575), .B(n40202), .X(n10276) );
  nor_x1_sg U60438 ( .A(n41582), .B(n41745), .X(n11095) );
  nor_x1_sg U60439 ( .A(n41581), .B(n41746), .X(n11914) );
  nor_x1_sg U60440 ( .A(n41580), .B(n40191), .X(n12733) );
  nor_x1_sg U60441 ( .A(n41579), .B(n41751), .X(n13552) );
  nor_x1_sg U60442 ( .A(n41586), .B(n40187), .X(n14371) );
  nor_x1_sg U60443 ( .A(n41585), .B(n41752), .X(n15190) );
  nor_x1_sg U60444 ( .A(n41584), .B(n40167), .X(n16009) );
  nor_x1_sg U60445 ( .A(n41587), .B(n41741), .X(n17647) );
  nor_x1_sg U60446 ( .A(n41583), .B(n41749), .X(n18468) );
  nor_x1_sg U60447 ( .A(n39731), .B(n41750), .X(n8384) );
  nor_x1_sg U60448 ( .A(n41656), .B(n41742), .X(n9202) );
  nor_x1_sg U60449 ( .A(n41651), .B(n40208), .X(n10022) );
  nor_x1_sg U60450 ( .A(n39740), .B(n41744), .X(n10841) );
  nor_x1_sg U60451 ( .A(n41649), .B(n40200), .X(n11660) );
  nor_x1_sg U60452 ( .A(n39746), .B(n40196), .X(n12479) );
  nor_x1_sg U60453 ( .A(n41655), .B(n40190), .X(n13298) );
  nor_x1_sg U60454 ( .A(n41654), .B(n40174), .X(n14117) );
  nor_x1_sg U60455 ( .A(n39755), .B(n40186), .X(n14936) );
  nor_x1_sg U60456 ( .A(n41652), .B(n40172), .X(n15755) );
  nor_x1_sg U60457 ( .A(n39761), .B(n40166), .X(n16574) );
  nor_x1_sg U60458 ( .A(n39764), .B(n40216), .X(n18212) );
  nor_x1_sg U60459 ( .A(n39766), .B(n40184), .X(n19033) );
  nor_x1_sg U60460 ( .A(n40304), .B(n16665), .X(n16663) );
  nor_x1_sg U60461 ( .A(n41666), .B(n40084), .X(n7002) );
  nor_x1_sg U60462 ( .A(n41915), .B(n40308), .X(n7975) );
  nor_x1_sg U60463 ( .A(n41916), .B(n41844), .X(n8793) );
  nor_x1_sg U60464 ( .A(n41907), .B(n41852), .X(n9613) );
  nor_x1_sg U60465 ( .A(n41909), .B(n41854), .X(n10432) );
  nor_x1_sg U60466 ( .A(n41913), .B(n41850), .X(n11251) );
  nor_x1_sg U60467 ( .A(n41914), .B(n41856), .X(n12070) );
  nor_x1_sg U60468 ( .A(n41908), .B(n41858), .X(n12889) );
  nor_x1_sg U60469 ( .A(n41911), .B(n41848), .X(n13708) );
  nor_x1_sg U60470 ( .A(n41917), .B(n41837), .X(n14527) );
  nor_x1_sg U60471 ( .A(n41904), .B(n41845), .X(n15346) );
  nor_x1_sg U60472 ( .A(n41905), .B(n41839), .X(n16165) );
  nor_x1_sg U60473 ( .A(n41912), .B(n40364), .X(n17803) );
  nor_x1_sg U60474 ( .A(n41906), .B(n41841), .X(n18624) );
  nor_x1_sg U60475 ( .A(n39726), .B(n40084), .X(n7431) );
  nor_x1_sg U60476 ( .A(n39726), .B(n40368), .X(n7256) );
  nor_x1_sg U60477 ( .A(n41693), .B(n40228), .X(n16826) );
  nor_x1_sg U60478 ( .A(n8312), .B(n8314), .X(n8350) );
  nor_x1_sg U60479 ( .A(n9130), .B(n9132), .X(n9168) );
  nor_x1_sg U60480 ( .A(n9950), .B(n9952), .X(n9988) );
  nor_x1_sg U60481 ( .A(n10769), .B(n10771), .X(n10807) );
  nor_x1_sg U60482 ( .A(n11588), .B(n11590), .X(n11626) );
  nor_x1_sg U60483 ( .A(n12407), .B(n12409), .X(n12445) );
  nor_x1_sg U60484 ( .A(n13226), .B(n13228), .X(n13264) );
  nor_x1_sg U60485 ( .A(n14045), .B(n14047), .X(n14083) );
  nor_x1_sg U60486 ( .A(n14864), .B(n14866), .X(n14902) );
  nor_x1_sg U60487 ( .A(n15683), .B(n15685), .X(n15721) );
  nor_x1_sg U60488 ( .A(n16502), .B(n16504), .X(n16540) );
  nor_x1_sg U60489 ( .A(n17319), .B(n17321), .X(n17357) );
  nor_x1_sg U60490 ( .A(n42019), .B(n18142), .X(n18178) );
  nor_x1_sg U60491 ( .A(n18961), .B(n18963), .X(n18999) );
  nor_x1_sg U60492 ( .A(n41983), .B(n40367), .X(n6968) );
  nor_x1_sg U60493 ( .A(n41984), .B(n40308), .X(n7785) );
  nor_x1_sg U60494 ( .A(n41985), .B(n41843), .X(n8603) );
  nor_x1_sg U60495 ( .A(n41979), .B(n41853), .X(n9423) );
  nor_x1_sg U60496 ( .A(n41980), .B(n41757), .X(n10242) );
  nor_x1_sg U60497 ( .A(n41981), .B(n41851), .X(n11061) );
  nor_x1_sg U60498 ( .A(n41982), .B(n41763), .X(n11880) );
  nor_x1_sg U60499 ( .A(n41975), .B(n41760), .X(n12699) );
  nor_x1_sg U60500 ( .A(n41976), .B(n41849), .X(n13518) );
  nor_x1_sg U60501 ( .A(n41977), .B(n41836), .X(n14337) );
  nor_x1_sg U60502 ( .A(n41978), .B(n41846), .X(n15156) );
  nor_x1_sg U60503 ( .A(n41972), .B(n41838), .X(n15975) );
  nor_x1_sg U60504 ( .A(n41973), .B(n50565), .X(n17613) );
  nor_x1_sg U60505 ( .A(n41974), .B(n41840), .X(n18434) );
  nor_x1_sg U60506 ( .A(n6834), .B(n6841), .X(n6839) );
  nor_x1_sg U60507 ( .A(n7494), .B(n7496), .X(n7532) );
  nor_x1_sg U60508 ( .A(n40560), .B(n7658), .X(n7656) );
  nor_x1_sg U60509 ( .A(n40555), .B(n8476), .X(n8474) );
  nor_x1_sg U60510 ( .A(n40551), .B(n9296), .X(n9294) );
  nor_x1_sg U60511 ( .A(n40548), .B(n10115), .X(n10113) );
  nor_x1_sg U60512 ( .A(n40544), .B(n10934), .X(n10932) );
  nor_x1_sg U60513 ( .A(n40539), .B(n11753), .X(n11751) );
  nor_x1_sg U60514 ( .A(n40537), .B(n12572), .X(n12570) );
  nor_x1_sg U60515 ( .A(n40531), .B(n13391), .X(n13389) );
  nor_x1_sg U60516 ( .A(n40527), .B(n14210), .X(n14208) );
  nor_x1_sg U60517 ( .A(n40523), .B(n15029), .X(n15027) );
  nor_x1_sg U60518 ( .A(n40520), .B(n15848), .X(n15846) );
  nor_x1_sg U60519 ( .A(n40516), .B(n17486), .X(n17484) );
  nor_x1_sg U60520 ( .A(n40511), .B(n18307), .X(n18305) );
  nand_x1_sg U60521 ( .A(n39772), .B(n40082), .X(n6962) );
  nand_x1_sg U60522 ( .A(n39520), .B(n40078), .X(n16786) );
  nor_x1_sg U60523 ( .A(n50394), .B(n17100), .X(n17099) );
  nor_x1_sg U60524 ( .A(n50353), .B(n17101), .X(n17098) );
  inv_x1_sg U60525 ( .A(n17100), .X(n50353) );
  nor_x1_sg U60526 ( .A(n50525), .B(n40310), .X(n16792) );
  nor_x1_sg U60527 ( .A(n6980), .B(n47122), .X(n6978) );
  nor_x1_sg U60528 ( .A(n6983), .B(n6982), .X(n6980) );
  nand_x1_sg U60529 ( .A(n6982), .B(n6983), .X(n6981) );
  nor_x1_sg U60530 ( .A(n7797), .B(n47408), .X(n7795) );
  nor_x1_sg U60531 ( .A(n7800), .B(n7799), .X(n7797) );
  nand_x1_sg U60532 ( .A(n7799), .B(n7800), .X(n7798) );
  nor_x1_sg U60533 ( .A(n8615), .B(n47693), .X(n8613) );
  nor_x1_sg U60534 ( .A(n8618), .B(n8617), .X(n8615) );
  nand_x1_sg U60535 ( .A(n8617), .B(n8618), .X(n8616) );
  nor_x1_sg U60536 ( .A(n9435), .B(n47978), .X(n9433) );
  nor_x1_sg U60537 ( .A(n9438), .B(n9437), .X(n9435) );
  nand_x1_sg U60538 ( .A(n9437), .B(n9438), .X(n9436) );
  nor_x1_sg U60539 ( .A(n10254), .B(n48263), .X(n10252) );
  nor_x1_sg U60540 ( .A(n10257), .B(n10256), .X(n10254) );
  nand_x1_sg U60541 ( .A(n10256), .B(n10257), .X(n10255) );
  nor_x1_sg U60542 ( .A(n11073), .B(n48548), .X(n11071) );
  nor_x1_sg U60543 ( .A(n11076), .B(n11075), .X(n11073) );
  nand_x1_sg U60544 ( .A(n11075), .B(n11076), .X(n11074) );
  nor_x1_sg U60545 ( .A(n11892), .B(n48833), .X(n11890) );
  nor_x1_sg U60546 ( .A(n11895), .B(n11894), .X(n11892) );
  nand_x1_sg U60547 ( .A(n11894), .B(n11895), .X(n11893) );
  nor_x1_sg U60548 ( .A(n12711), .B(n49120), .X(n12709) );
  nor_x1_sg U60549 ( .A(n12714), .B(n12713), .X(n12711) );
  nand_x1_sg U60550 ( .A(n12713), .B(n12714), .X(n12712) );
  nor_x1_sg U60551 ( .A(n13530), .B(n49406), .X(n13528) );
  nor_x1_sg U60552 ( .A(n13533), .B(n13532), .X(n13530) );
  nand_x1_sg U60553 ( .A(n13532), .B(n13533), .X(n13531) );
  nor_x1_sg U60554 ( .A(n14349), .B(n49692), .X(n14347) );
  nor_x1_sg U60555 ( .A(n14352), .B(n14351), .X(n14349) );
  nand_x1_sg U60556 ( .A(n14351), .B(n14352), .X(n14350) );
  nor_x1_sg U60557 ( .A(n15168), .B(n49978), .X(n15166) );
  nor_x1_sg U60558 ( .A(n15171), .B(n15170), .X(n15168) );
  nand_x1_sg U60559 ( .A(n15170), .B(n15171), .X(n15169) );
  nor_x1_sg U60560 ( .A(n15987), .B(n50264), .X(n15985) );
  nor_x1_sg U60561 ( .A(n15990), .B(n15989), .X(n15987) );
  nand_x1_sg U60562 ( .A(n15989), .B(n15990), .X(n15988) );
  nor_x1_sg U60563 ( .A(n16804), .B(n50550), .X(n16802) );
  nor_x1_sg U60564 ( .A(n16807), .B(n16806), .X(n16804) );
  nand_x1_sg U60565 ( .A(n16806), .B(n16807), .X(n16805) );
  nor_x1_sg U60566 ( .A(n17625), .B(n50838), .X(n17623) );
  nor_x1_sg U60567 ( .A(n17628), .B(n17627), .X(n17625) );
  nand_x1_sg U60568 ( .A(n17627), .B(n17628), .X(n17626) );
  nor_x1_sg U60569 ( .A(n18446), .B(n51125), .X(n18444) );
  nor_x1_sg U60570 ( .A(n18449), .B(n18448), .X(n18446) );
  nand_x1_sg U60571 ( .A(n18448), .B(n18449), .X(n18447) );
  nor_x1_sg U60572 ( .A(n47358), .B(n42311), .X(n22972) );
  nor_x1_sg U60573 ( .A(n47643), .B(n42310), .X(n23249) );
  nor_x1_sg U60574 ( .A(n47928), .B(n42309), .X(n23529) );
  nor_x1_sg U60575 ( .A(n48213), .B(n10272), .X(n23808) );
  nor_x1_sg U60576 ( .A(n48498), .B(n42308), .X(n24087) );
  nor_x1_sg U60577 ( .A(n48783), .B(n42307), .X(n24366) );
  nor_x1_sg U60578 ( .A(n49070), .B(n42306), .X(n24645) );
  nor_x1_sg U60579 ( .A(n49356), .B(n13548), .X(n24923) );
  nor_x1_sg U60580 ( .A(n49642), .B(n42305), .X(n25202) );
  nor_x1_sg U60581 ( .A(n49928), .B(n42304), .X(n25481) );
  nor_x1_sg U60582 ( .A(n50214), .B(n42303), .X(n25760) );
  nor_x1_sg U60583 ( .A(n50788), .B(n17643), .X(n26317) );
  nor_x1_sg U60584 ( .A(n51075), .B(n18464), .X(n26597) );
  nor_x1_sg U60585 ( .A(n47072), .B(n42312), .X(n22698) );
  nor_x1_sg U60586 ( .A(n6995), .B(n39290), .X(n6992) );
  nand_x1_sg U60587 ( .A(n39350), .B(n39678), .X(n6995) );
  nor_x1_sg U60588 ( .A(n7812), .B(n39315), .X(n7809) );
  nand_x1_sg U60589 ( .A(n39352), .B(n39677), .X(n7812) );
  nor_x1_sg U60590 ( .A(n8630), .B(n8631), .X(n8627) );
  nand_x1_sg U60591 ( .A(n39351), .B(n39676), .X(n8630) );
  nor_x1_sg U60592 ( .A(n9450), .B(n39312), .X(n9447) );
  nand_x1_sg U60593 ( .A(n39353), .B(n39674), .X(n9450) );
  nor_x1_sg U60594 ( .A(n10269), .B(n39310), .X(n10266) );
  nand_x1_sg U60595 ( .A(n39355), .B(n10272), .X(n10269) );
  nor_x1_sg U60596 ( .A(n11088), .B(n11089), .X(n11085) );
  nand_x1_sg U60597 ( .A(n39354), .B(n39673), .X(n11088) );
  nor_x1_sg U60598 ( .A(n11907), .B(n39306), .X(n11904) );
  nand_x1_sg U60599 ( .A(n39356), .B(n39672), .X(n11907) );
  nor_x1_sg U60600 ( .A(n12726), .B(n12727), .X(n12723) );
  nand_x1_sg U60601 ( .A(n39358), .B(n39670), .X(n12726) );
  nor_x1_sg U60602 ( .A(n13545), .B(n13546), .X(n13542) );
  nand_x1_sg U60603 ( .A(n39357), .B(n13548), .X(n13545) );
  nor_x1_sg U60604 ( .A(n14364), .B(n14365), .X(n14361) );
  nand_x1_sg U60605 ( .A(n39359), .B(n39669), .X(n14364) );
  nor_x1_sg U60606 ( .A(n15183), .B(n15184), .X(n15180) );
  nand_x1_sg U60607 ( .A(n39361), .B(n39668), .X(n15183) );
  nor_x1_sg U60608 ( .A(n16002), .B(n39296), .X(n15999) );
  nand_x1_sg U60609 ( .A(n39360), .B(n39666), .X(n16002) );
  nor_x1_sg U60610 ( .A(n16819), .B(n16820), .X(n16816) );
  nand_x1_sg U60611 ( .A(n39364), .B(n39806), .X(n16819) );
  nor_x1_sg U60612 ( .A(n17640), .B(n39292), .X(n17637) );
  nand_x1_sg U60613 ( .A(n39363), .B(n17643), .X(n17640) );
  nor_x1_sg U60614 ( .A(n18461), .B(n18462), .X(n18458) );
  nand_x1_sg U60615 ( .A(n39362), .B(n18464), .X(n18461) );
  nand_x1_sg U60616 ( .A(n22635), .B(n22636), .X(n22634) );
  nand_x1_sg U60617 ( .A(n22639), .B(n40224), .X(n22633) );
  nand_x1_sg U60618 ( .A(n40081), .B(n22637), .X(n22636) );
  nand_x1_sg U60619 ( .A(n25965), .B(n50560), .X(n25964) );
  nand_x1_sg U60620 ( .A(n25968), .B(n41317), .X(n25963) );
  inv_x1_sg U60621 ( .A(n25966), .X(n50560) );
  nand_x1_sg U60622 ( .A(n26260), .B(n26261), .X(n26259) );
  nand_x1_sg U60623 ( .A(n26263), .B(n39276), .X(n26258) );
  nand_x1_sg U60624 ( .A(n39530), .B(n26262), .X(n26261) );
  nand_x1_sg U60625 ( .A(n26276), .B(n26277), .X(n26275) );
  nand_x1_sg U60626 ( .A(n26279), .B(n39278), .X(n26274) );
  nand_x1_sg U60627 ( .A(n39543), .B(n26278), .X(n26277) );
  nand_x1_sg U60628 ( .A(n26292), .B(n26293), .X(n26291) );
  nand_x1_sg U60629 ( .A(n26295), .B(n39927), .X(n26290) );
  nand_x1_sg U60630 ( .A(n39516), .B(n26294), .X(n26293) );
  nand_x1_sg U60631 ( .A(n25990), .B(n25991), .X(n25989) );
  nor_x1_sg U60632 ( .A(n25994), .B(n41405), .X(n25993) );
  nand_x1_sg U60633 ( .A(n26003), .B(n26004), .X(n26002) );
  nor_x1_sg U60634 ( .A(n26007), .B(n40456), .X(n26006) );
  nor_x1_sg U60635 ( .A(n46945), .B(n7251), .X(n7229) );
  nor_x1_sg U60636 ( .A(n7252), .B(n7253), .X(n7251) );
  nand_x1_sg U60637 ( .A(n7253), .B(n7252), .X(n7254) );
  nor_x1_sg U60638 ( .A(n50377), .B(n17076), .X(n17054) );
  nor_x1_sg U60639 ( .A(n17077), .B(n17078), .X(n17076) );
  nor_x1_sg U60640 ( .A(n46893), .B(n7136), .X(n7135) );
  inv_x1_sg U60641 ( .A(n7139), .X(n46893) );
  nor_x1_sg U60642 ( .A(n7137), .B(n7138), .X(n7136) );
  nor_x1_sg U60643 ( .A(n47188), .B(n7954), .X(n7953) );
  inv_x1_sg U60644 ( .A(n7957), .X(n47188) );
  nor_x1_sg U60645 ( .A(n7955), .B(n7956), .X(n7954) );
  nor_x1_sg U60646 ( .A(n47473), .B(n8772), .X(n8771) );
  inv_x1_sg U60647 ( .A(n8775), .X(n47473) );
  nor_x1_sg U60648 ( .A(n8773), .B(n8774), .X(n8772) );
  nor_x1_sg U60649 ( .A(n47758), .B(n9592), .X(n9591) );
  inv_x1_sg U60650 ( .A(n9595), .X(n47758) );
  nor_x1_sg U60651 ( .A(n9593), .B(n9594), .X(n9592) );
  nor_x1_sg U60652 ( .A(n48043), .B(n10411), .X(n10410) );
  inv_x1_sg U60653 ( .A(n10414), .X(n48043) );
  nor_x1_sg U60654 ( .A(n10412), .B(n10413), .X(n10411) );
  nor_x1_sg U60655 ( .A(n48328), .B(n11230), .X(n11229) );
  inv_x1_sg U60656 ( .A(n11233), .X(n48328) );
  nor_x1_sg U60657 ( .A(n11231), .B(n11232), .X(n11230) );
  nor_x1_sg U60658 ( .A(n48613), .B(n12049), .X(n12048) );
  inv_x1_sg U60659 ( .A(n12052), .X(n48613) );
  nor_x1_sg U60660 ( .A(n12050), .B(n12051), .X(n12049) );
  nor_x1_sg U60661 ( .A(n48899), .B(n12868), .X(n12867) );
  inv_x1_sg U60662 ( .A(n12871), .X(n48899) );
  nor_x1_sg U60663 ( .A(n12869), .B(n12870), .X(n12868) );
  nor_x1_sg U60664 ( .A(n49186), .B(n13687), .X(n13686) );
  inv_x1_sg U60665 ( .A(n13690), .X(n49186) );
  nor_x1_sg U60666 ( .A(n13688), .B(n13689), .X(n13687) );
  nor_x1_sg U60667 ( .A(n49472), .B(n14506), .X(n14505) );
  inv_x1_sg U60668 ( .A(n14509), .X(n49472) );
  nor_x1_sg U60669 ( .A(n14507), .B(n14508), .X(n14506) );
  nor_x1_sg U60670 ( .A(n49758), .B(n15325), .X(n15324) );
  inv_x1_sg U60671 ( .A(n15328), .X(n49758) );
  nor_x1_sg U60672 ( .A(n15326), .B(n15327), .X(n15325) );
  nor_x1_sg U60673 ( .A(n50044), .B(n16144), .X(n16143) );
  inv_x1_sg U60674 ( .A(n16147), .X(n50044) );
  nor_x1_sg U60675 ( .A(n16145), .B(n16146), .X(n16144) );
  nor_x1_sg U60676 ( .A(n50326), .B(n16961), .X(n16960) );
  inv_x1_sg U60677 ( .A(n16964), .X(n50326) );
  nor_x1_sg U60678 ( .A(n16962), .B(n16963), .X(n16961) );
  nor_x1_sg U60679 ( .A(n50618), .B(n17782), .X(n17781) );
  inv_x1_sg U60680 ( .A(n17785), .X(n50618) );
  nor_x1_sg U60681 ( .A(n17783), .B(n17784), .X(n17782) );
  nor_x1_sg U60682 ( .A(n50905), .B(n18603), .X(n18602) );
  inv_x1_sg U60683 ( .A(n18606), .X(n50905) );
  nor_x1_sg U60684 ( .A(n18604), .B(n18605), .X(n18603) );
  nor_x1_sg U60685 ( .A(n47011), .B(n7390), .X(n7360) );
  inv_x1_sg U60686 ( .A(n7393), .X(n47011) );
  nor_x1_sg U60687 ( .A(n7391), .B(n7392), .X(n7390) );
  nor_x1_sg U60688 ( .A(n47299), .B(n8208), .X(n8178) );
  inv_x1_sg U60689 ( .A(n8211), .X(n47299) );
  nor_x1_sg U60690 ( .A(n8209), .B(n8210), .X(n8208) );
  nor_x1_sg U60691 ( .A(n47584), .B(n9026), .X(n8996) );
  inv_x1_sg U60692 ( .A(n9029), .X(n47584) );
  nor_x1_sg U60693 ( .A(n9027), .B(n9028), .X(n9026) );
  nor_x1_sg U60694 ( .A(n47869), .B(n9846), .X(n9816) );
  inv_x1_sg U60695 ( .A(n9849), .X(n47869) );
  nor_x1_sg U60696 ( .A(n9847), .B(n9848), .X(n9846) );
  nor_x1_sg U60697 ( .A(n48154), .B(n10665), .X(n10635) );
  inv_x1_sg U60698 ( .A(n10668), .X(n48154) );
  nor_x1_sg U60699 ( .A(n10666), .B(n10667), .X(n10665) );
  nor_x1_sg U60700 ( .A(n48439), .B(n11484), .X(n11454) );
  inv_x1_sg U60701 ( .A(n11487), .X(n48439) );
  nor_x1_sg U60702 ( .A(n11485), .B(n11486), .X(n11484) );
  nor_x1_sg U60703 ( .A(n48724), .B(n12303), .X(n12273) );
  inv_x1_sg U60704 ( .A(n12306), .X(n48724) );
  nor_x1_sg U60705 ( .A(n12304), .B(n12305), .X(n12303) );
  nor_x1_sg U60706 ( .A(n49010), .B(n13122), .X(n13092) );
  inv_x1_sg U60707 ( .A(n13125), .X(n49010) );
  nor_x1_sg U60708 ( .A(n13123), .B(n13124), .X(n13122) );
  nor_x1_sg U60709 ( .A(n49297), .B(n13941), .X(n13911) );
  inv_x1_sg U60710 ( .A(n13944), .X(n49297) );
  nor_x1_sg U60711 ( .A(n13942), .B(n13943), .X(n13941) );
  nor_x1_sg U60712 ( .A(n49583), .B(n14760), .X(n14730) );
  inv_x1_sg U60713 ( .A(n14763), .X(n49583) );
  nor_x1_sg U60714 ( .A(n14761), .B(n14762), .X(n14760) );
  nor_x1_sg U60715 ( .A(n49869), .B(n15579), .X(n15549) );
  inv_x1_sg U60716 ( .A(n15582), .X(n49869) );
  nor_x1_sg U60717 ( .A(n15580), .B(n15581), .X(n15579) );
  nor_x1_sg U60718 ( .A(n50155), .B(n16398), .X(n16368) );
  inv_x1_sg U60719 ( .A(n16401), .X(n50155) );
  nor_x1_sg U60720 ( .A(n16399), .B(n16400), .X(n16398) );
  nor_x1_sg U60721 ( .A(n50440), .B(n17215), .X(n17185) );
  inv_x1_sg U60722 ( .A(n17218), .X(n50440) );
  nor_x1_sg U60723 ( .A(n17216), .B(n17217), .X(n17215) );
  nor_x1_sg U60724 ( .A(n50729), .B(n18036), .X(n18006) );
  inv_x1_sg U60725 ( .A(n18039), .X(n50729) );
  nor_x1_sg U60726 ( .A(n18037), .B(n18038), .X(n18036) );
  nor_x1_sg U60727 ( .A(n51016), .B(n18857), .X(n18827) );
  inv_x1_sg U60728 ( .A(n18860), .X(n51016) );
  nor_x1_sg U60729 ( .A(n18858), .B(n18859), .X(n18857) );
  nand_x1_sg U60730 ( .A(n7104), .B(n41604), .X(n7108) );
  nand_x1_sg U60731 ( .A(n7922), .B(n41605), .X(n7926) );
  nand_x1_sg U60732 ( .A(n8740), .B(n41606), .X(n8744) );
  nand_x1_sg U60733 ( .A(n9560), .B(n41607), .X(n9564) );
  nand_x1_sg U60734 ( .A(n10379), .B(n41608), .X(n10383) );
  nand_x1_sg U60735 ( .A(n11198), .B(n41609), .X(n11202) );
  nand_x1_sg U60736 ( .A(n12017), .B(n41610), .X(n12021) );
  nand_x1_sg U60737 ( .A(n12836), .B(n41611), .X(n12840) );
  nand_x1_sg U60738 ( .A(n13655), .B(n41612), .X(n13659) );
  nand_x1_sg U60739 ( .A(n14474), .B(n41613), .X(n14478) );
  nand_x1_sg U60740 ( .A(n15293), .B(n41614), .X(n15297) );
  nand_x1_sg U60741 ( .A(n16112), .B(n41615), .X(n16116) );
  nand_x1_sg U60742 ( .A(n17750), .B(n41616), .X(n17754) );
  nand_x1_sg U60743 ( .A(n18571), .B(n41617), .X(n18575) );
  nor_x1_sg U60744 ( .A(n40085), .B(n41710), .X(n6957) );
  nor_x1_sg U60745 ( .A(n40088), .B(n41724), .X(n16781) );
  nor_x1_sg U60746 ( .A(n40178), .B(n41712), .X(n7774) );
  nor_x1_sg U60747 ( .A(n40210), .B(n41711), .X(n8592) );
  nor_x1_sg U60748 ( .A(n40207), .B(n41714), .X(n9412) );
  nor_x1_sg U60749 ( .A(n40202), .B(n41713), .X(n10231) );
  nor_x1_sg U60750 ( .A(n40199), .B(n41716), .X(n11050) );
  nor_x1_sg U60751 ( .A(n40195), .B(n41715), .X(n11869) );
  nor_x1_sg U60752 ( .A(n41747), .B(n41718), .X(n12688) );
  nor_x1_sg U60753 ( .A(n40175), .B(n41717), .X(n13507) );
  nor_x1_sg U60754 ( .A(n41748), .B(n41720), .X(n14326) );
  nor_x1_sg U60755 ( .A(n40171), .B(n41719), .X(n15145) );
  nor_x1_sg U60756 ( .A(n41753), .B(n41722), .X(n15964) );
  nor_x1_sg U60757 ( .A(n40215), .B(n41721), .X(n17602) );
  nor_x1_sg U60758 ( .A(n40183), .B(n41723), .X(n18423) );
  nand_x1_sg U60759 ( .A(n40089), .B(n41740), .X(n21720) );
  nor_x1_sg U60760 ( .A(n39726), .B(n41631), .X(n7629) );
  nor_x1_sg U60761 ( .A(n39545), .B(n41618), .X(n17454) );
  nand_x1_sg U60762 ( .A(n22894), .B(n39366), .X(n22901) );
  nand_x1_sg U60763 ( .A(n23171), .B(n39368), .X(n23178) );
  nand_x1_sg U60764 ( .A(n23451), .B(n39370), .X(n23458) );
  nand_x1_sg U60765 ( .A(n23730), .B(n39372), .X(n23737) );
  nand_x1_sg U60766 ( .A(n24009), .B(n39374), .X(n24016) );
  nand_x1_sg U60767 ( .A(n24288), .B(n39376), .X(n24295) );
  nand_x1_sg U60768 ( .A(n24567), .B(n39378), .X(n24574) );
  nand_x1_sg U60769 ( .A(n24845), .B(n39380), .X(n24852) );
  nand_x1_sg U60770 ( .A(n25124), .B(n39382), .X(n25131) );
  nand_x1_sg U60771 ( .A(n25403), .B(n39384), .X(n25410) );
  nand_x1_sg U60772 ( .A(n25682), .B(n39386), .X(n25689) );
  nand_x1_sg U60773 ( .A(n26228), .B(n39390), .X(n26236) );
  nand_x1_sg U60774 ( .A(n26519), .B(n39388), .X(n26526) );
  nor_x1_sg U60775 ( .A(n39806), .B(n17458), .X(n26038) );
  nand_x1_sg U60776 ( .A(n16665), .B(n40609), .X(n16895) );
  nand_x1_sg U60777 ( .A(n6841), .B(n41902), .X(n7068) );
  nand_x1_sg U60778 ( .A(n7658), .B(n41900), .X(n7886) );
  nand_x1_sg U60779 ( .A(n8476), .B(n39830), .X(n8704) );
  nand_x1_sg U60780 ( .A(n9296), .B(n39846), .X(n9524) );
  nand_x1_sg U60781 ( .A(n10115), .B(n41898), .X(n10343) );
  nand_x1_sg U60782 ( .A(n10934), .B(n39833), .X(n11162) );
  nand_x1_sg U60783 ( .A(n11753), .B(n41884), .X(n11981) );
  nand_x1_sg U60784 ( .A(n12572), .B(n39818), .X(n12800) );
  nand_x1_sg U60785 ( .A(n13391), .B(n41882), .X(n13619) );
  nand_x1_sg U60786 ( .A(n14210), .B(n41880), .X(n14438) );
  nand_x1_sg U60787 ( .A(n15029), .B(n41875), .X(n15257) );
  nand_x1_sg U60788 ( .A(n15848), .B(n39822), .X(n16076) );
  nand_x1_sg U60789 ( .A(n17486), .B(n39827), .X(n17714) );
  nand_x1_sg U60790 ( .A(n18307), .B(n39824), .X(n18535) );
  nand_x1_sg U60791 ( .A(n40074), .B(n40077), .X(n17042) );
  nor_x1_sg U60792 ( .A(n42285), .B(n38923), .X(n6653) );
  nor_x1_sg U60793 ( .A(n40105), .B(n22910), .X(n22909) );
  nand_x1_sg U60794 ( .A(n41195), .B(n22901), .X(n22910) );
  nor_x1_sg U60795 ( .A(n40107), .B(n23187), .X(n23186) );
  nand_x1_sg U60796 ( .A(n40502), .B(n23178), .X(n23187) );
  nor_x1_sg U60797 ( .A(n40110), .B(n23467), .X(n23466) );
  nand_x1_sg U60798 ( .A(n39226), .B(n23458), .X(n23467) );
  nor_x1_sg U60799 ( .A(n40111), .B(n23746), .X(n23745) );
  nand_x1_sg U60800 ( .A(n39228), .B(n23737), .X(n23746) );
  nor_x1_sg U60801 ( .A(n40113), .B(n24025), .X(n24024) );
  nand_x1_sg U60802 ( .A(n41174), .B(n24016), .X(n24025) );
  nor_x1_sg U60803 ( .A(n40116), .B(n24304), .X(n24303) );
  nand_x1_sg U60804 ( .A(n41170), .B(n24295), .X(n24304) );
  nor_x1_sg U60805 ( .A(n40117), .B(n24583), .X(n24582) );
  nand_x1_sg U60806 ( .A(n40482), .B(n24574), .X(n24583) );
  nor_x1_sg U60807 ( .A(n13768), .B(n24861), .X(n24860) );
  nand_x1_sg U60808 ( .A(n41157), .B(n24852), .X(n24861) );
  nor_x1_sg U60809 ( .A(n40122), .B(n25140), .X(n25139) );
  nand_x1_sg U60810 ( .A(n39238), .B(n25131), .X(n25140) );
  nor_x1_sg U60811 ( .A(n40124), .B(n25419), .X(n25418) );
  nand_x1_sg U60812 ( .A(n41150), .B(n25410), .X(n25419) );
  nor_x1_sg U60813 ( .A(n40125), .B(n25698), .X(n25697) );
  nand_x1_sg U60814 ( .A(n41145), .B(n25689), .X(n25698) );
  nor_x1_sg U60815 ( .A(n40129), .B(n25967), .X(n25966) );
  nand_x1_sg U60816 ( .A(n41947), .B(n25958), .X(n25967) );
  nor_x1_sg U60817 ( .A(n40131), .B(n26246), .X(n26245) );
  nand_x1_sg U60818 ( .A(n41139), .B(n26236), .X(n26246) );
  nor_x1_sg U60819 ( .A(n40128), .B(n26535), .X(n26534) );
  nand_x1_sg U60820 ( .A(n41134), .B(n26526), .X(n26535) );
  nor_x1_sg U60821 ( .A(n22691), .B(n39678), .X(n22690) );
  nor_x1_sg U60822 ( .A(n22965), .B(n39677), .X(n22964) );
  nor_x1_sg U60823 ( .A(n23242), .B(n39676), .X(n23241) );
  nor_x1_sg U60824 ( .A(n23522), .B(n39674), .X(n23521) );
  nor_x1_sg U60825 ( .A(n23801), .B(n39675), .X(n23800) );
  nor_x1_sg U60826 ( .A(n24080), .B(n39673), .X(n24079) );
  nor_x1_sg U60827 ( .A(n24359), .B(n39672), .X(n24358) );
  nor_x1_sg U60828 ( .A(n24638), .B(n39670), .X(n24637) );
  nor_x1_sg U60829 ( .A(n24916), .B(n39671), .X(n24915) );
  nor_x1_sg U60830 ( .A(n25195), .B(n39669), .X(n25194) );
  nor_x1_sg U60831 ( .A(n25474), .B(n39668), .X(n25473) );
  nor_x1_sg U60832 ( .A(n25753), .B(n39666), .X(n25752) );
  nor_x1_sg U60833 ( .A(n26309), .B(n39667), .X(n26308) );
  nor_x1_sg U60834 ( .A(n26590), .B(n39665), .X(n26589) );
  nor_x1_sg U60835 ( .A(n6068), .B(n41004), .X(n6067) );
  nor_x1_sg U60836 ( .A(n6119), .B(n41008), .X(n6116) );
  nor_x1_sg U60837 ( .A(n39137), .B(n7300), .X(n22663) );
  nor_x1_sg U60838 ( .A(n41862), .B(n42161), .X(n22932) );
  nor_x1_sg U60839 ( .A(n41190), .B(n8936), .X(n23209) );
  nor_x1_sg U60840 ( .A(n41185), .B(n9756), .X(n23489) );
  nor_x1_sg U60841 ( .A(n41179), .B(n10575), .X(n23768) );
  nor_x1_sg U60842 ( .A(n39230), .B(n11394), .X(n24047) );
  nor_x1_sg U60843 ( .A(n41169), .B(n12213), .X(n24326) );
  nor_x1_sg U60844 ( .A(n41164), .B(n13032), .X(n24605) );
  nor_x1_sg U60845 ( .A(n41158), .B(n13851), .X(n24883) );
  nor_x1_sg U60846 ( .A(n41153), .B(n14670), .X(n25162) );
  nor_x1_sg U60847 ( .A(n41149), .B(n42160), .X(n25441) );
  nor_x1_sg U60848 ( .A(n41144), .B(n16308), .X(n25720) );
  nor_x1_sg U60849 ( .A(n41295), .B(n17125), .X(n25987) );
  nor_x1_sg U60850 ( .A(n41873), .B(n17946), .X(n26271) );
  nor_x1_sg U60851 ( .A(n41874), .B(n18767), .X(n26557) );
  nand_x1_sg U60852 ( .A(n40584), .B(n39095), .X(n16647) );
  nand_x1_sg U60853 ( .A(n47187), .B(n40106), .X(n22908) );
  inv_x1_sg U60854 ( .A(n22901), .X(n47187) );
  nand_x1_sg U60855 ( .A(n47472), .B(n40107), .X(n23185) );
  inv_x1_sg U60856 ( .A(n23178), .X(n47472) );
  nand_x1_sg U60857 ( .A(n47757), .B(n40109), .X(n23465) );
  inv_x1_sg U60858 ( .A(n23458), .X(n47757) );
  nand_x1_sg U60859 ( .A(n48042), .B(n40111), .X(n23744) );
  inv_x1_sg U60860 ( .A(n23737), .X(n48042) );
  nand_x1_sg U60861 ( .A(n48327), .B(n40113), .X(n24023) );
  inv_x1_sg U60862 ( .A(n24016), .X(n48327) );
  nand_x1_sg U60863 ( .A(n48612), .B(n40115), .X(n24302) );
  inv_x1_sg U60864 ( .A(n24295), .X(n48612) );
  nand_x1_sg U60865 ( .A(n48898), .B(n40117), .X(n24581) );
  inv_x1_sg U60866 ( .A(n24574), .X(n48898) );
  nand_x1_sg U60867 ( .A(n49185), .B(n40120), .X(n24859) );
  inv_x1_sg U60868 ( .A(n24852), .X(n49185) );
  nand_x1_sg U60869 ( .A(n49471), .B(n40121), .X(n25138) );
  inv_x1_sg U60870 ( .A(n25131), .X(n49471) );
  nand_x1_sg U60871 ( .A(n49757), .B(n40124), .X(n25417) );
  inv_x1_sg U60872 ( .A(n25410), .X(n49757) );
  nand_x1_sg U60873 ( .A(n50043), .B(n40125), .X(n25696) );
  inv_x1_sg U60874 ( .A(n25689), .X(n50043) );
  nand_x1_sg U60875 ( .A(n50335), .B(n40129), .X(n25965) );
  inv_x1_sg U60876 ( .A(n25958), .X(n50335) );
  nand_x1_sg U60877 ( .A(n50617), .B(n17863), .X(n26244) );
  inv_x1_sg U60878 ( .A(n26236), .X(n50617) );
  nand_x1_sg U60879 ( .A(n50904), .B(n40127), .X(n26533) );
  inv_x1_sg U60880 ( .A(n26526), .X(n50904) );
  inv_x1_sg U60881 ( .A(n6020), .X(n46567) );
  inv_x1_sg U60882 ( .A(n6119), .X(n46476) );
  inv_x1_sg U60883 ( .A(n6068), .X(n46518) );
  nor_x1_sg U60884 ( .A(n7324), .B(n40080), .X(n7323) );
  nor_x1_sg U60885 ( .A(n17149), .B(n40076), .X(n17148) );
  nand_x1_sg U60886 ( .A(n42311), .B(n22965), .X(n22963) );
  nand_x1_sg U60887 ( .A(n42310), .B(n23242), .X(n23240) );
  nand_x1_sg U60888 ( .A(n42308), .B(n24080), .X(n24078) );
  nand_x1_sg U60889 ( .A(n42307), .B(n24359), .X(n24357) );
  nand_x1_sg U60890 ( .A(n39671), .B(n24916), .X(n24914) );
  nand_x1_sg U60891 ( .A(n42305), .B(n25195), .X(n25193) );
  nand_x1_sg U60892 ( .A(n42304), .B(n25474), .X(n25472) );
  nand_x1_sg U60893 ( .A(n42303), .B(n25753), .X(n25751) );
  nand_x1_sg U60894 ( .A(n42309), .B(n23522), .X(n23520) );
  nand_x1_sg U60895 ( .A(n39675), .B(n23801), .X(n23799) );
  nand_x1_sg U60896 ( .A(n39665), .B(n26590), .X(n26588) );
  nand_x1_sg U60897 ( .A(n17162), .B(n39560), .X(n17161) );
  nand_x1_sg U60898 ( .A(n50332), .B(n16966), .X(n17160) );
  nor_x1_sg U60899 ( .A(n17113), .B(n39681), .X(n17162) );
  nor_x1_sg U60900 ( .A(n41305), .B(n6991), .X(n22669) );
  nor_x1_sg U60901 ( .A(n39659), .B(n39663), .X(n22681) );
  nor_x1_sg U60902 ( .A(n7498), .B(n7499), .X(n7497) );
  nor_x1_sg U60903 ( .A(n8316), .B(n8317), .X(n8315) );
  nor_x1_sg U60904 ( .A(n9134), .B(n9135), .X(n9133) );
  nor_x1_sg U60905 ( .A(n9954), .B(n9955), .X(n9953) );
  nor_x1_sg U60906 ( .A(n10773), .B(n10774), .X(n10772) );
  nor_x1_sg U60907 ( .A(n11592), .B(n11593), .X(n11591) );
  nor_x1_sg U60908 ( .A(n12411), .B(n12412), .X(n12410) );
  nor_x1_sg U60909 ( .A(n13230), .B(n13231), .X(n13229) );
  nor_x1_sg U60910 ( .A(n14049), .B(n14050), .X(n14048) );
  nor_x1_sg U60911 ( .A(n14868), .B(n14869), .X(n14867) );
  nor_x1_sg U60912 ( .A(n15687), .B(n15688), .X(n15686) );
  nor_x1_sg U60913 ( .A(n16506), .B(n16507), .X(n16505) );
  nor_x1_sg U60914 ( .A(n17323), .B(n17324), .X(n17322) );
  nor_x1_sg U60915 ( .A(n18144), .B(n18145), .X(n18143) );
  nor_x1_sg U60916 ( .A(n18965), .B(n18966), .X(n18964) );
  nor_x1_sg U60917 ( .A(n7147), .B(n7148), .X(n7146) );
  nor_x1_sg U60918 ( .A(n7965), .B(n7966), .X(n7964) );
  nor_x1_sg U60919 ( .A(n8783), .B(n8784), .X(n8782) );
  nor_x1_sg U60920 ( .A(n9603), .B(n9604), .X(n9602) );
  nor_x1_sg U60921 ( .A(n10422), .B(n10423), .X(n10421) );
  nor_x1_sg U60922 ( .A(n11241), .B(n11242), .X(n11240) );
  nor_x1_sg U60923 ( .A(n12060), .B(n12061), .X(n12059) );
  nor_x1_sg U60924 ( .A(n12879), .B(n12880), .X(n12878) );
  nor_x1_sg U60925 ( .A(n13698), .B(n13699), .X(n13697) );
  nor_x1_sg U60926 ( .A(n14517), .B(n14518), .X(n14516) );
  nor_x1_sg U60927 ( .A(n15336), .B(n15337), .X(n15335) );
  nor_x1_sg U60928 ( .A(n16155), .B(n16156), .X(n16154) );
  nor_x1_sg U60929 ( .A(n16972), .B(n16973), .X(n16971) );
  nor_x1_sg U60930 ( .A(n17793), .B(n17794), .X(n17792) );
  nor_x1_sg U60931 ( .A(n18614), .B(n18615), .X(n18613) );
  nor_x1_sg U60932 ( .A(n7089), .B(n7090), .X(n7088) );
  nor_x1_sg U60933 ( .A(n7907), .B(n7908), .X(n7906) );
  nor_x1_sg U60934 ( .A(n8725), .B(n8726), .X(n8724) );
  nor_x1_sg U60935 ( .A(n9545), .B(n9546), .X(n9544) );
  nor_x1_sg U60936 ( .A(n10364), .B(n10365), .X(n10363) );
  nor_x1_sg U60937 ( .A(n11183), .B(n11184), .X(n11182) );
  nor_x1_sg U60938 ( .A(n12002), .B(n12003), .X(n12001) );
  nor_x1_sg U60939 ( .A(n12821), .B(n12822), .X(n12820) );
  nor_x1_sg U60940 ( .A(n13640), .B(n13641), .X(n13639) );
  nor_x1_sg U60941 ( .A(n14459), .B(n14460), .X(n14458) );
  nor_x1_sg U60942 ( .A(n15278), .B(n15279), .X(n15277) );
  nor_x1_sg U60943 ( .A(n16097), .B(n16098), .X(n16096) );
  nor_x1_sg U60944 ( .A(n16915), .B(n16916), .X(n16914) );
  nor_x1_sg U60945 ( .A(n17735), .B(n17736), .X(n17734) );
  nor_x1_sg U60946 ( .A(n18556), .B(n18557), .X(n18555) );
  nor_x1_sg U60947 ( .A(n26017), .B(n39807), .X(n26016) );
  nor_x1_sg U60948 ( .A(n41296), .B(n16815), .X(n25994) );
  nor_x1_sg U60949 ( .A(n39481), .B(n17299), .X(n26007) );
  nand_x1_sg U60950 ( .A(n47078), .B(n46973), .X(n7574) );
  nand_x1_sg U60951 ( .A(n7576), .B(n41599), .X(n7575) );
  nor_x1_sg U60952 ( .A(n41725), .B(n39854), .X(n7576) );
  nand_x1_sg U60953 ( .A(n47364), .B(n47263), .X(n8392) );
  nand_x1_sg U60954 ( .A(n8394), .B(n41602), .X(n8393) );
  nor_x1_sg U60955 ( .A(n39612), .B(n39894), .X(n8394) );
  nand_x1_sg U60956 ( .A(n47649), .B(n47548), .X(n9210) );
  nand_x1_sg U60957 ( .A(n9212), .B(n41597), .X(n9211) );
  nor_x1_sg U60958 ( .A(n39608), .B(n41687), .X(n9212) );
  nand_x1_sg U60959 ( .A(n47934), .B(n47833), .X(n10030) );
  nand_x1_sg U60960 ( .A(n10032), .B(n41596), .X(n10031) );
  nor_x1_sg U60961 ( .A(n39627), .B(n41689), .X(n10032) );
  nand_x1_sg U60962 ( .A(n48219), .B(n48118), .X(n10849) );
  nand_x1_sg U60963 ( .A(n10851), .B(n41595), .X(n10850) );
  nor_x1_sg U60964 ( .A(n39624), .B(n41685), .X(n10851) );
  nand_x1_sg U60965 ( .A(n48504), .B(n48403), .X(n11668) );
  nand_x1_sg U60966 ( .A(n11670), .B(n41594), .X(n11669) );
  nor_x1_sg U60967 ( .A(n39621), .B(n41683), .X(n11670) );
  nand_x1_sg U60968 ( .A(n48789), .B(n48688), .X(n12487) );
  nand_x1_sg U60969 ( .A(n12489), .B(n41593), .X(n12488) );
  nor_x1_sg U60970 ( .A(n39618), .B(n41681), .X(n12489) );
  nand_x1_sg U60971 ( .A(n49076), .B(n48974), .X(n13306) );
  nand_x1_sg U60972 ( .A(n13308), .B(n41592), .X(n13307) );
  nor_x1_sg U60973 ( .A(n39639), .B(n41679), .X(n13308) );
  nand_x1_sg U60974 ( .A(n49362), .B(n49261), .X(n14125) );
  nand_x1_sg U60975 ( .A(n14127), .B(n41591), .X(n14126) );
  nor_x1_sg U60976 ( .A(n39636), .B(n41677), .X(n14127) );
  nand_x1_sg U60977 ( .A(n49648), .B(n49547), .X(n14944) );
  nand_x1_sg U60978 ( .A(n14946), .B(n41590), .X(n14945) );
  nor_x1_sg U60979 ( .A(n39633), .B(n41675), .X(n14946) );
  nand_x1_sg U60980 ( .A(n49934), .B(n49833), .X(n15763) );
  nand_x1_sg U60981 ( .A(n15765), .B(n41601), .X(n15764) );
  nor_x1_sg U60982 ( .A(n39630), .B(n39896), .X(n15765) );
  nand_x1_sg U60983 ( .A(n50220), .B(n50119), .X(n16582) );
  nand_x1_sg U60984 ( .A(n16584), .B(n41589), .X(n16583) );
  nor_x1_sg U60985 ( .A(n39648), .B(n41673), .X(n16584) );
  nand_x1_sg U60986 ( .A(n50505), .B(n50404), .X(n17399) );
  nand_x1_sg U60987 ( .A(n17401), .B(n41598), .X(n17400) );
  nor_x1_sg U60988 ( .A(n39615), .B(n39884), .X(n17401) );
  nand_x1_sg U60989 ( .A(n50794), .B(n50693), .X(n18220) );
  nand_x1_sg U60990 ( .A(n18222), .B(n41600), .X(n18221) );
  nor_x1_sg U60991 ( .A(n39645), .B(n39887), .X(n18222) );
  nand_x1_sg U60992 ( .A(n51081), .B(n50980), .X(n19041) );
  nand_x1_sg U60993 ( .A(n19043), .B(n41588), .X(n19042) );
  nor_x1_sg U60994 ( .A(n39642), .B(n41667), .X(n19043) );
  nor_x1_sg U60995 ( .A(n40304), .B(n39884), .X(n17265) );
  nand_x1_sg U60996 ( .A(n7287), .B(n7288), .X(n7286) );
  nor_x1_sg U60997 ( .A(n7288), .B(n7287), .X(n7289) );
  nand_x1_sg U60998 ( .A(n8105), .B(n8106), .X(n8104) );
  nor_x1_sg U60999 ( .A(n8106), .B(n8105), .X(n8107) );
  nand_x1_sg U61000 ( .A(n8923), .B(n8924), .X(n8922) );
  nor_x1_sg U61001 ( .A(n8924), .B(n8923), .X(n8925) );
  nand_x1_sg U61002 ( .A(n9743), .B(n9744), .X(n9742) );
  nor_x1_sg U61003 ( .A(n9744), .B(n9743), .X(n9745) );
  nand_x1_sg U61004 ( .A(n10562), .B(n10563), .X(n10561) );
  nor_x1_sg U61005 ( .A(n10563), .B(n10562), .X(n10564) );
  nand_x1_sg U61006 ( .A(n11381), .B(n11382), .X(n11380) );
  nor_x1_sg U61007 ( .A(n11382), .B(n11381), .X(n11383) );
  nand_x1_sg U61008 ( .A(n12200), .B(n12201), .X(n12199) );
  nor_x1_sg U61009 ( .A(n12201), .B(n12200), .X(n12202) );
  nand_x1_sg U61010 ( .A(n13019), .B(n13020), .X(n13018) );
  nor_x1_sg U61011 ( .A(n13020), .B(n13019), .X(n13021) );
  nand_x1_sg U61012 ( .A(n13838), .B(n13839), .X(n13837) );
  nor_x1_sg U61013 ( .A(n13839), .B(n13838), .X(n13840) );
  nand_x1_sg U61014 ( .A(n14657), .B(n14658), .X(n14656) );
  nor_x1_sg U61015 ( .A(n14658), .B(n14657), .X(n14659) );
  nand_x1_sg U61016 ( .A(n15476), .B(n15477), .X(n15475) );
  nor_x1_sg U61017 ( .A(n15477), .B(n15476), .X(n15478) );
  nand_x1_sg U61018 ( .A(n16295), .B(n16296), .X(n16294) );
  nor_x1_sg U61019 ( .A(n16296), .B(n16295), .X(n16297) );
  nand_x1_sg U61020 ( .A(n17933), .B(n17934), .X(n17932) );
  nor_x1_sg U61021 ( .A(n17934), .B(n17933), .X(n17935) );
  nand_x1_sg U61022 ( .A(n18754), .B(n18755), .X(n18753) );
  nor_x1_sg U61023 ( .A(n18755), .B(n18754), .X(n18756) );
  nand_x1_sg U61024 ( .A(n7097), .B(n7095), .X(n7096) );
  nor_x1_sg U61025 ( .A(n7095), .B(n7097), .X(n7098) );
  nand_x1_sg U61026 ( .A(n7915), .B(n7913), .X(n7914) );
  nor_x1_sg U61027 ( .A(n7913), .B(n7915), .X(n7916) );
  nand_x1_sg U61028 ( .A(n8733), .B(n8731), .X(n8732) );
  nor_x1_sg U61029 ( .A(n8731), .B(n8733), .X(n8734) );
  nand_x1_sg U61030 ( .A(n9553), .B(n9551), .X(n9552) );
  nor_x1_sg U61031 ( .A(n9551), .B(n9553), .X(n9554) );
  nand_x1_sg U61032 ( .A(n10372), .B(n10370), .X(n10371) );
  nor_x1_sg U61033 ( .A(n10370), .B(n10372), .X(n10373) );
  nand_x1_sg U61034 ( .A(n11191), .B(n11189), .X(n11190) );
  nor_x1_sg U61035 ( .A(n11189), .B(n11191), .X(n11192) );
  nand_x1_sg U61036 ( .A(n12010), .B(n12008), .X(n12009) );
  nor_x1_sg U61037 ( .A(n12008), .B(n12010), .X(n12011) );
  nand_x1_sg U61038 ( .A(n12829), .B(n12827), .X(n12828) );
  nor_x1_sg U61039 ( .A(n12827), .B(n12829), .X(n12830) );
  nand_x1_sg U61040 ( .A(n13648), .B(n13646), .X(n13647) );
  nor_x1_sg U61041 ( .A(n13646), .B(n13648), .X(n13649) );
  nand_x1_sg U61042 ( .A(n14467), .B(n14465), .X(n14466) );
  nor_x1_sg U61043 ( .A(n14465), .B(n14467), .X(n14468) );
  nand_x1_sg U61044 ( .A(n15286), .B(n15284), .X(n15285) );
  nor_x1_sg U61045 ( .A(n15284), .B(n15286), .X(n15287) );
  nand_x1_sg U61046 ( .A(n16105), .B(n16103), .X(n16104) );
  nor_x1_sg U61047 ( .A(n16103), .B(n16105), .X(n16106) );
  nand_x1_sg U61048 ( .A(n16922), .B(n16920), .X(n16921) );
  nor_x1_sg U61049 ( .A(n16920), .B(n16922), .X(n16923) );
  nand_x1_sg U61050 ( .A(n17743), .B(n17741), .X(n17742) );
  nor_x1_sg U61051 ( .A(n17741), .B(n17743), .X(n17744) );
  nand_x1_sg U61052 ( .A(n18564), .B(n18562), .X(n18563) );
  nor_x1_sg U61053 ( .A(n18562), .B(n18564), .X(n18565) );
  nor_x1_sg U61054 ( .A(n41194), .B(n42324), .X(n22918) );
  nor_x1_sg U61055 ( .A(n41192), .B(n39799), .X(n22946) );
  nor_x1_sg U61056 ( .A(n39222), .B(n7814), .X(n22960) );
  nor_x1_sg U61057 ( .A(n41189), .B(n42323), .X(n23195) );
  nor_x1_sg U61058 ( .A(n41187), .B(n39801), .X(n23223) );
  nor_x1_sg U61059 ( .A(n41190), .B(n8632), .X(n23237) );
  nor_x1_sg U61060 ( .A(n39226), .B(n42322), .X(n23475) );
  nor_x1_sg U61061 ( .A(n41184), .B(n39795), .X(n23503) );
  nor_x1_sg U61062 ( .A(n39226), .B(n9452), .X(n23517) );
  nor_x1_sg U61063 ( .A(n41179), .B(n10311), .X(n23754) );
  nor_x1_sg U61064 ( .A(n41177), .B(n39797), .X(n23782) );
  nor_x1_sg U61065 ( .A(n41178), .B(n10271), .X(n23796) );
  nor_x1_sg U61066 ( .A(n39230), .B(n11130), .X(n24033) );
  nor_x1_sg U61067 ( .A(n41175), .B(n39791), .X(n24061) );
  nor_x1_sg U61068 ( .A(n41173), .B(n11090), .X(n24075) );
  nor_x1_sg U61069 ( .A(n41867), .B(n11949), .X(n24312) );
  nor_x1_sg U61070 ( .A(n41170), .B(n39793), .X(n24340) );
  nor_x1_sg U61071 ( .A(n41169), .B(n11909), .X(n24354) );
  nor_x1_sg U61072 ( .A(n41162), .B(n12768), .X(n24591) );
  nor_x1_sg U61073 ( .A(n41164), .B(n39787), .X(n24619) );
  nor_x1_sg U61074 ( .A(n41868), .B(n12728), .X(n24633) );
  nor_x1_sg U61075 ( .A(n41157), .B(n13587), .X(n24869) );
  nor_x1_sg U61076 ( .A(n39236), .B(n39789), .X(n24897) );
  nor_x1_sg U61077 ( .A(n41159), .B(n13547), .X(n24911) );
  nor_x1_sg U61078 ( .A(n41154), .B(n14406), .X(n25148) );
  nor_x1_sg U61079 ( .A(n39238), .B(n39783), .X(n25176) );
  nor_x1_sg U61080 ( .A(n41154), .B(n14366), .X(n25190) );
  nor_x1_sg U61081 ( .A(n41147), .B(n15225), .X(n25427) );
  nor_x1_sg U61082 ( .A(n41148), .B(n39785), .X(n25455) );
  nor_x1_sg U61083 ( .A(n41148), .B(n15185), .X(n25469) );
  nor_x1_sg U61084 ( .A(n41142), .B(n16044), .X(n25706) );
  nor_x1_sg U61085 ( .A(n41143), .B(n39779), .X(n25734) );
  nor_x1_sg U61086 ( .A(n41142), .B(n16004), .X(n25748) );
  nor_x1_sg U61087 ( .A(n41138), .B(n42321), .X(n26255) );
  nor_x1_sg U61088 ( .A(n41138), .B(n39781), .X(n26287) );
  nor_x1_sg U61089 ( .A(n41137), .B(n17642), .X(n26303) );
  nor_x1_sg U61090 ( .A(n41134), .B(n42320), .X(n26543) );
  nor_x1_sg U61091 ( .A(n41135), .B(n39777), .X(n26571) );
  nor_x1_sg U61092 ( .A(n39246), .B(n18463), .X(n26585) );
  nor_x1_sg U61093 ( .A(n39809), .B(n41304), .X(n22613) );
  nor_x1_sg U61094 ( .A(n41900), .B(n41193), .X(n22876) );
  nor_x1_sg U61095 ( .A(n41888), .B(n41189), .X(n23153) );
  nor_x1_sg U61096 ( .A(n39846), .B(n41185), .X(n23433) );
  nor_x1_sg U61097 ( .A(n41898), .B(n41865), .X(n23712) );
  nor_x1_sg U61098 ( .A(n41886), .B(n41172), .X(n23991) );
  nor_x1_sg U61099 ( .A(n39836), .B(n41170), .X(n24270) );
  nor_x1_sg U61100 ( .A(n41896), .B(n39234), .X(n24549) );
  nor_x1_sg U61101 ( .A(n41882), .B(n39236), .X(n24827) );
  nor_x1_sg U61102 ( .A(n39843), .B(n41152), .X(n25106) );
  nor_x1_sg U61103 ( .A(n39849), .B(n41150), .X(n25385) );
  nor_x1_sg U61104 ( .A(n39822), .B(n41872), .X(n25664) );
  nor_x1_sg U61105 ( .A(n39827), .B(n41139), .X(n26207) );
  nor_x1_sg U61106 ( .A(n41892), .B(n39246), .X(n26501) );
  nand_x1_sg U61107 ( .A(n7006), .B(n7131), .X(n7389) );
  nand_x1_sg U61108 ( .A(n16830), .B(n16956), .X(n17214) );
  nand_x1_sg U61109 ( .A(n39564), .B(n39939), .X(n8410) );
  nand_x1_sg U61110 ( .A(n39567), .B(n39941), .X(n9228) );
  nand_x1_sg U61111 ( .A(n39569), .B(n39943), .X(n10048) );
  nand_x1_sg U61112 ( .A(n39573), .B(n39959), .X(n10867) );
  nand_x1_sg U61113 ( .A(n39576), .B(n39960), .X(n11686) );
  nand_x1_sg U61114 ( .A(n39578), .B(n39951), .X(n12505) );
  nand_x1_sg U61115 ( .A(n39582), .B(n39953), .X(n13324) );
  nand_x1_sg U61116 ( .A(n39585), .B(n39955), .X(n14143) );
  nand_x1_sg U61117 ( .A(n39587), .B(n39949), .X(n14962) );
  nand_x1_sg U61118 ( .A(n39591), .B(n39945), .X(n15781) );
  nand_x1_sg U61119 ( .A(n39594), .B(n39947), .X(n16600) );
  nand_x1_sg U61120 ( .A(n39560), .B(n39933), .X(n17417) );
  nand_x1_sg U61121 ( .A(n39599), .B(n39935), .X(n18238) );
  nand_x1_sg U61122 ( .A(n39596), .B(n39937), .X(n19059) );
  nor_x1_sg U61123 ( .A(n40613), .B(n41691), .X(n7440) );
  nor_x1_sg U61124 ( .A(n22968), .B(n22969), .X(n22967) );
  nor_x1_sg U61125 ( .A(n22970), .B(n40508), .X(n22968) );
  nor_x1_sg U61126 ( .A(n39222), .B(n8451), .X(n22969) );
  nor_x1_sg U61127 ( .A(n23245), .B(n23246), .X(n23244) );
  nor_x1_sg U61128 ( .A(n23247), .B(n40505), .X(n23245) );
  nor_x1_sg U61129 ( .A(n41188), .B(n9269), .X(n23246) );
  nand_x4_sg U61130 ( .A(n24082), .B(n41312), .X(n24081) );
  nor_x1_sg U61131 ( .A(n24083), .B(n24084), .X(n24082) );
  nor_x1_sg U61132 ( .A(n24085), .B(n40491), .X(n24083) );
  nor_x1_sg U61133 ( .A(n41174), .B(n11727), .X(n24084) );
  nand_x4_sg U61134 ( .A(n24361), .B(n41462), .X(n24360) );
  nor_x1_sg U61135 ( .A(n24362), .B(n24363), .X(n24361) );
  nor_x1_sg U61136 ( .A(n24364), .B(n40487), .X(n24362) );
  nor_x1_sg U61137 ( .A(n41167), .B(n12546), .X(n24363) );
  nor_x1_sg U61138 ( .A(n24641), .B(n24642), .X(n24640) );
  nor_x1_sg U61139 ( .A(n24643), .B(n24533), .X(n24641) );
  nor_x1_sg U61140 ( .A(n41162), .B(n13365), .X(n24642) );
  nand_x4_sg U61141 ( .A(n24918), .B(n39658), .X(n24917) );
  nor_x1_sg U61142 ( .A(n24919), .B(n24920), .X(n24918) );
  nor_x1_sg U61143 ( .A(n24921), .B(n40481), .X(n24919) );
  nor_x1_sg U61144 ( .A(n41160), .B(n14184), .X(n24920) );
  nor_x1_sg U61145 ( .A(n25198), .B(n25199), .X(n25197) );
  nor_x1_sg U61146 ( .A(n25200), .B(n25090), .X(n25198) );
  nor_x1_sg U61147 ( .A(n39238), .B(n15003), .X(n25199) );
  nand_x4_sg U61148 ( .A(n25476), .B(n41318), .X(n25475) );
  nor_x1_sg U61149 ( .A(n25477), .B(n25478), .X(n25476) );
  nor_x1_sg U61150 ( .A(n25479), .B(n40473), .X(n25477) );
  nor_x1_sg U61151 ( .A(n41147), .B(n15822), .X(n25478) );
  nor_x1_sg U61152 ( .A(n25756), .B(n25757), .X(n25755) );
  nor_x1_sg U61153 ( .A(n25758), .B(n40468), .X(n25756) );
  nor_x1_sg U61154 ( .A(n39242), .B(n16641), .X(n25757) );
  nand_x4_sg U61155 ( .A(n23524), .B(n39657), .X(n23523) );
  nor_x1_sg U61156 ( .A(n23525), .B(n23526), .X(n23524) );
  nor_x1_sg U61157 ( .A(n23527), .B(n40499), .X(n23525) );
  nor_x1_sg U61158 ( .A(n41864), .B(n10089), .X(n23526) );
  nand_x4_sg U61159 ( .A(n23803), .B(n41313), .X(n23802) );
  nor_x1_sg U61160 ( .A(n23804), .B(n23805), .X(n23803) );
  nor_x1_sg U61161 ( .A(n23806), .B(n40497), .X(n23804) );
  nor_x1_sg U61162 ( .A(n41178), .B(n10908), .X(n23805) );
  nor_x1_sg U61163 ( .A(n26593), .B(n26594), .X(n26592) );
  nor_x1_sg U61164 ( .A(n26595), .B(n40460), .X(n26593) );
  nor_x1_sg U61165 ( .A(n41133), .B(n19100), .X(n26594) );
  nor_x1_sg U61166 ( .A(n41777), .B(n22894), .X(n22903) );
  nor_x1_sg U61167 ( .A(n41776), .B(n23171), .X(n23180) );
  nor_x1_sg U61168 ( .A(n41775), .B(n23451), .X(n23460) );
  nor_x1_sg U61169 ( .A(n41774), .B(n23730), .X(n23739) );
  nor_x1_sg U61170 ( .A(n41773), .B(n24009), .X(n24018) );
  nor_x1_sg U61171 ( .A(n41772), .B(n24288), .X(n24297) );
  nor_x1_sg U61172 ( .A(n41771), .B(n24567), .X(n24576) );
  nor_x1_sg U61173 ( .A(n41770), .B(n24845), .X(n24854) );
  nor_x1_sg U61174 ( .A(n41769), .B(n25124), .X(n25133) );
  nor_x1_sg U61175 ( .A(n41768), .B(n25403), .X(n25412) );
  nor_x1_sg U61176 ( .A(n41767), .B(n25682), .X(n25691) );
  nor_x1_sg U61177 ( .A(n41755), .B(n26228), .X(n26238) );
  nor_x1_sg U61178 ( .A(n41766), .B(n26519), .X(n26528) );
  nor_x1_sg U61179 ( .A(n40561), .B(n39893), .X(n8258) );
  nor_x1_sg U61180 ( .A(n8469), .B(n39860), .X(n9076) );
  nor_x1_sg U61181 ( .A(n9289), .B(n39857), .X(n9896) );
  nor_x1_sg U61182 ( .A(n10108), .B(n39863), .X(n10715) );
  nor_x1_sg U61183 ( .A(n40543), .B(n39866), .X(n11534) );
  nor_x1_sg U61184 ( .A(n40540), .B(n39869), .X(n12353) );
  nor_x1_sg U61185 ( .A(n12565), .B(n39872), .X(n13172) );
  nor_x1_sg U61186 ( .A(n13384), .B(n39875), .X(n13991) );
  nor_x1_sg U61187 ( .A(n14203), .B(n39878), .X(n14810) );
  nor_x1_sg U61188 ( .A(n15022), .B(n41662), .X(n15629) );
  nor_x1_sg U61189 ( .A(n40519), .B(n39881), .X(n16448) );
  nor_x1_sg U61190 ( .A(n40515), .B(n39888), .X(n18086) );
  nor_x1_sg U61191 ( .A(n40512), .B(n39890), .X(n18907) );
  nand_x1_sg U61192 ( .A(n7380), .B(n7217), .X(n7378) );
  nor_x1_sg U61193 ( .A(n7217), .B(n7380), .X(n7379) );
  nand_x1_sg U61194 ( .A(n8198), .B(n8036), .X(n8196) );
  nor_x1_sg U61195 ( .A(n8036), .B(n8198), .X(n8197) );
  nand_x1_sg U61196 ( .A(n9016), .B(n8854), .X(n9014) );
  nor_x1_sg U61197 ( .A(n8854), .B(n9016), .X(n9015) );
  nand_x1_sg U61198 ( .A(n9836), .B(n9674), .X(n9834) );
  nor_x1_sg U61199 ( .A(n9674), .B(n9836), .X(n9835) );
  nand_x1_sg U61200 ( .A(n10655), .B(n10493), .X(n10653) );
  nor_x1_sg U61201 ( .A(n10493), .B(n10655), .X(n10654) );
  nand_x1_sg U61202 ( .A(n11474), .B(n11312), .X(n11472) );
  nor_x1_sg U61203 ( .A(n11312), .B(n11474), .X(n11473) );
  nand_x1_sg U61204 ( .A(n12293), .B(n12131), .X(n12291) );
  nor_x1_sg U61205 ( .A(n12131), .B(n12293), .X(n12292) );
  nand_x1_sg U61206 ( .A(n13112), .B(n12950), .X(n13110) );
  nor_x1_sg U61207 ( .A(n12950), .B(n13112), .X(n13111) );
  nand_x1_sg U61208 ( .A(n13931), .B(n13769), .X(n13929) );
  nor_x1_sg U61209 ( .A(n13769), .B(n13931), .X(n13930) );
  nand_x1_sg U61210 ( .A(n14750), .B(n14588), .X(n14748) );
  nor_x1_sg U61211 ( .A(n14588), .B(n14750), .X(n14749) );
  nand_x1_sg U61212 ( .A(n15569), .B(n15407), .X(n15567) );
  nor_x1_sg U61213 ( .A(n15407), .B(n15569), .X(n15568) );
  nand_x1_sg U61214 ( .A(n16388), .B(n16226), .X(n16386) );
  nor_x1_sg U61215 ( .A(n16226), .B(n16388), .X(n16387) );
  nand_x1_sg U61216 ( .A(n18026), .B(n17864), .X(n18024) );
  nor_x1_sg U61217 ( .A(n17864), .B(n18026), .X(n18025) );
  nand_x1_sg U61218 ( .A(n18847), .B(n18685), .X(n18845) );
  nor_x1_sg U61219 ( .A(n18685), .B(n18847), .X(n18846) );
  nor_x1_sg U61220 ( .A(n39137), .B(n6997), .X(n22687) );
  nor_x1_sg U61221 ( .A(n39482), .B(n16821), .X(n26013) );
  nor_x1_sg U61222 ( .A(n40072), .B(n38941), .X(n25948) );
  nor_x1_sg U61223 ( .A(n40610), .B(n40036), .X(n25936) );
  nor_x1_sg U61224 ( .A(n39348), .B(n39724), .X(n22650) );
  nor_x1_sg U61225 ( .A(n41306), .B(n39773), .X(n22657) );
  nor_x1_sg U61226 ( .A(n41307), .B(n39803), .X(n22675) );
  nand_x1_sg U61227 ( .A(n39347), .B(n7225), .X(n7224) );
  nor_x1_sg U61228 ( .A(n7225), .B(n7141), .X(n7226) );
  nand_x1_sg U61229 ( .A(n39345), .B(n8044), .X(n8043) );
  nor_x1_sg U61230 ( .A(n8044), .B(n7959), .X(n8045) );
  nand_x1_sg U61231 ( .A(n39343), .B(n8862), .X(n8861) );
  nor_x1_sg U61232 ( .A(n8862), .B(n8777), .X(n8863) );
  nand_x1_sg U61233 ( .A(n39341), .B(n9682), .X(n9681) );
  nor_x1_sg U61234 ( .A(n9682), .B(n9597), .X(n9683) );
  nand_x1_sg U61235 ( .A(n39339), .B(n10501), .X(n10500) );
  nor_x1_sg U61236 ( .A(n10501), .B(n10416), .X(n10502) );
  nand_x1_sg U61237 ( .A(n39337), .B(n11320), .X(n11319) );
  nor_x1_sg U61238 ( .A(n11320), .B(n11235), .X(n11321) );
  nand_x1_sg U61239 ( .A(n39335), .B(n12139), .X(n12138) );
  nor_x1_sg U61240 ( .A(n12139), .B(n12054), .X(n12140) );
  nand_x1_sg U61241 ( .A(n39333), .B(n12958), .X(n12957) );
  nor_x1_sg U61242 ( .A(n12958), .B(n12873), .X(n12959) );
  nand_x1_sg U61243 ( .A(n39331), .B(n13777), .X(n13776) );
  nor_x1_sg U61244 ( .A(n13777), .B(n13692), .X(n13778) );
  nand_x1_sg U61245 ( .A(n39329), .B(n14596), .X(n14595) );
  nor_x1_sg U61246 ( .A(n14596), .B(n14511), .X(n14597) );
  nand_x1_sg U61247 ( .A(n39327), .B(n15415), .X(n15414) );
  nor_x1_sg U61248 ( .A(n15415), .B(n15330), .X(n15416) );
  nand_x1_sg U61249 ( .A(n39325), .B(n16234), .X(n16233) );
  nor_x1_sg U61250 ( .A(n16234), .B(n16149), .X(n16235) );
  nand_x1_sg U61251 ( .A(n39323), .B(n17872), .X(n17871) );
  nor_x1_sg U61252 ( .A(n17872), .B(n17787), .X(n17873) );
  nand_x1_sg U61253 ( .A(n39321), .B(n18693), .X(n18692) );
  nor_x1_sg U61254 ( .A(n18693), .B(n18608), .X(n18694) );
  nand_x1_sg U61255 ( .A(n39319), .B(n17050), .X(n17049) );
  nor_x1_sg U61256 ( .A(n17050), .B(n16966), .X(n17051) );
  nand_x1_sg U61257 ( .A(n8429), .B(n8430), .X(n8428) );
  nor_x1_sg U61258 ( .A(n8430), .B(n8429), .X(n8431) );
  nand_x1_sg U61259 ( .A(n9247), .B(n9248), .X(n9246) );
  nor_x1_sg U61260 ( .A(n9248), .B(n9247), .X(n9249) );
  nand_x1_sg U61261 ( .A(n10067), .B(n10068), .X(n10066) );
  nor_x1_sg U61262 ( .A(n10068), .B(n10067), .X(n10069) );
  nand_x1_sg U61263 ( .A(n10886), .B(n10887), .X(n10885) );
  nor_x1_sg U61264 ( .A(n10887), .B(n10886), .X(n10888) );
  nand_x1_sg U61265 ( .A(n11705), .B(n11706), .X(n11704) );
  nor_x1_sg U61266 ( .A(n11706), .B(n11705), .X(n11707) );
  nand_x1_sg U61267 ( .A(n12524), .B(n12525), .X(n12523) );
  nor_x1_sg U61268 ( .A(n12525), .B(n12524), .X(n12526) );
  nand_x1_sg U61269 ( .A(n13343), .B(n13344), .X(n13342) );
  nor_x1_sg U61270 ( .A(n13344), .B(n13343), .X(n13345) );
  nand_x1_sg U61271 ( .A(n14162), .B(n14163), .X(n14161) );
  nor_x1_sg U61272 ( .A(n14163), .B(n14162), .X(n14164) );
  nand_x1_sg U61273 ( .A(n14981), .B(n14982), .X(n14980) );
  nor_x1_sg U61274 ( .A(n14982), .B(n14981), .X(n14983) );
  nand_x1_sg U61275 ( .A(n15800), .B(n15801), .X(n15799) );
  nor_x1_sg U61276 ( .A(n15801), .B(n15800), .X(n15802) );
  nand_x1_sg U61277 ( .A(n16619), .B(n16620), .X(n16618) );
  nor_x1_sg U61278 ( .A(n16620), .B(n16619), .X(n16621) );
  nand_x1_sg U61279 ( .A(n18257), .B(n18258), .X(n18256) );
  nor_x1_sg U61280 ( .A(n18258), .B(n18257), .X(n18259) );
  nand_x1_sg U61281 ( .A(n19078), .B(n19079), .X(n19077) );
  nor_x1_sg U61282 ( .A(n19079), .B(n19078), .X(n19080) );
  nand_x1_sg U61283 ( .A(n7431), .B(n7432), .X(n7430) );
  nor_x1_sg U61284 ( .A(n7432), .B(n7431), .X(n7433) );
  nand_x1_sg U61285 ( .A(n8249), .B(n8250), .X(n8248) );
  nor_x1_sg U61286 ( .A(n8250), .B(n8249), .X(n8251) );
  nand_x1_sg U61287 ( .A(n9067), .B(n9068), .X(n9066) );
  nor_x1_sg U61288 ( .A(n9068), .B(n9067), .X(n9069) );
  nand_x1_sg U61289 ( .A(n9887), .B(n9888), .X(n9886) );
  nor_x1_sg U61290 ( .A(n9888), .B(n9887), .X(n9889) );
  nand_x1_sg U61291 ( .A(n10706), .B(n10707), .X(n10705) );
  nor_x1_sg U61292 ( .A(n10707), .B(n10706), .X(n10708) );
  nand_x1_sg U61293 ( .A(n11525), .B(n11526), .X(n11524) );
  nor_x1_sg U61294 ( .A(n11526), .B(n11525), .X(n11527) );
  nand_x1_sg U61295 ( .A(n12344), .B(n12345), .X(n12343) );
  nor_x1_sg U61296 ( .A(n12345), .B(n12344), .X(n12346) );
  nand_x1_sg U61297 ( .A(n13163), .B(n13164), .X(n13162) );
  nor_x1_sg U61298 ( .A(n13164), .B(n13163), .X(n13165) );
  nand_x1_sg U61299 ( .A(n13982), .B(n13983), .X(n13981) );
  nor_x1_sg U61300 ( .A(n13983), .B(n13982), .X(n13984) );
  nand_x1_sg U61301 ( .A(n14801), .B(n14802), .X(n14800) );
  nor_x1_sg U61302 ( .A(n14802), .B(n14801), .X(n14803) );
  nand_x1_sg U61303 ( .A(n15620), .B(n15621), .X(n15619) );
  nor_x1_sg U61304 ( .A(n15621), .B(n15620), .X(n15622) );
  nand_x1_sg U61305 ( .A(n16439), .B(n16440), .X(n16438) );
  nor_x1_sg U61306 ( .A(n16440), .B(n16439), .X(n16441) );
  nand_x1_sg U61307 ( .A(n18077), .B(n18078), .X(n18076) );
  nor_x1_sg U61308 ( .A(n18078), .B(n18077), .X(n18079) );
  nand_x1_sg U61309 ( .A(n18898), .B(n18899), .X(n18897) );
  nor_x1_sg U61310 ( .A(n18899), .B(n18898), .X(n18900) );
  nor_x1_sg U61311 ( .A(n41970), .B(n38931), .X(n6163) );
  nand_x1_sg U61312 ( .A(n41901), .B(n39663), .X(n7593) );
  nor_x1_sg U61313 ( .A(n42259), .B(n41567), .X(n6103) );
  nor_x1_sg U61314 ( .A(n42262), .B(n41566), .X(n6114) );
  nor_x1_sg U61315 ( .A(n42257), .B(n41035), .X(n6148) );
  nor_x1_sg U61316 ( .A(n42256), .B(n41036), .X(n6194) );
  nor_x1_sg U61317 ( .A(n42214), .B(n41036), .X(n6241) );
  nor_x1_sg U61318 ( .A(n42213), .B(n41008), .X(n6256) );
  nor_x1_sg U61319 ( .A(n42212), .B(n41567), .X(n6286) );
  nor_x1_sg U61320 ( .A(n42211), .B(n41010), .X(n6301) );
  nor_x1_sg U61321 ( .A(n42210), .B(n41034), .X(n6330) );
  nor_x1_sg U61322 ( .A(n42209), .B(n41010), .X(n6345) );
  nor_x1_sg U61323 ( .A(n42152), .B(n41033), .X(n6375) );
  nor_x1_sg U61324 ( .A(n42208), .B(n41010), .X(n6390) );
  nor_x1_sg U61325 ( .A(n42207), .B(n41034), .X(n6419) );
  nor_x1_sg U61326 ( .A(n42206), .B(n41009), .X(n6434) );
  nor_x1_sg U61327 ( .A(n42151), .B(n38929), .X(n6464) );
  nor_x1_sg U61328 ( .A(n42205), .B(n41011), .X(n6479) );
  nor_x1_sg U61329 ( .A(n42150), .B(n41034), .X(n6508) );
  nor_x1_sg U61330 ( .A(n42149), .B(n41008), .X(n6523) );
  nor_x1_sg U61331 ( .A(n42204), .B(n41035), .X(n6553) );
  nor_x1_sg U61332 ( .A(n42203), .B(n41008), .X(n6568) );
  nor_x1_sg U61333 ( .A(n42148), .B(n41033), .X(n6597) );
  nor_x1_sg U61334 ( .A(n42202), .B(n41009), .X(n6612) );
  nor_x1_sg U61335 ( .A(n42201), .B(n38929), .X(n6642) );
  nor_x1_sg U61336 ( .A(n42227), .B(n38933), .X(n6704) );
  nor_x1_sg U61337 ( .A(n42229), .B(n41015), .X(n6731) );
  nand_x1_sg U61338 ( .A(n40080), .B(n40162), .X(n7215) );
  nand_x1_sg U61339 ( .A(n39560), .B(n40072), .X(n17257) );
  nand_x1_sg U61340 ( .A(n39563), .B(n42345), .X(n7786) );
  nand_x1_sg U61341 ( .A(n39566), .B(n39518), .X(n8604) );
  nand_x1_sg U61342 ( .A(n39569), .B(n39524), .X(n9424) );
  nand_x1_sg U61343 ( .A(n39572), .B(n42354), .X(n10243) );
  nand_x1_sg U61344 ( .A(n39575), .B(n42353), .X(n11062) );
  nand_x1_sg U61345 ( .A(n39578), .B(n39521), .X(n11881) );
  nand_x1_sg U61346 ( .A(n39581), .B(n39528), .X(n12700) );
  nand_x1_sg U61347 ( .A(n39584), .B(n42350), .X(n13519) );
  nand_x1_sg U61348 ( .A(n39587), .B(n42349), .X(n14338) );
  nand_x1_sg U61349 ( .A(n39590), .B(n39525), .X(n15157) );
  nand_x1_sg U61350 ( .A(n39593), .B(n39531), .X(n15976) );
  nand_x1_sg U61351 ( .A(n39561), .B(n42336), .X(n16793) );
  nand_x1_sg U61352 ( .A(n39599), .B(n42356), .X(n17614) );
  nand_x1_sg U61353 ( .A(n39596), .B(n42346), .X(n18435) );
  nand_x1_sg U61354 ( .A(n40611), .B(n39662), .X(n17418) );
  nor_x1_sg U61355 ( .A(n40507), .B(n22943), .X(n22952) );
  nor_x1_sg U61356 ( .A(n23137), .B(n23220), .X(n23229) );
  nor_x1_sg U61357 ( .A(n40500), .B(n23500), .X(n23509) );
  nor_x1_sg U61358 ( .A(n40495), .B(n23779), .X(n23788) );
  nor_x1_sg U61359 ( .A(n23975), .B(n24058), .X(n24067) );
  nor_x1_sg U61360 ( .A(n40487), .B(n24337), .X(n24346) );
  nor_x1_sg U61361 ( .A(n40483), .B(n24616), .X(n24625) );
  nor_x1_sg U61362 ( .A(n40480), .B(n24894), .X(n24903) );
  nor_x1_sg U61363 ( .A(n25090), .B(n25173), .X(n25182) );
  nor_x1_sg U61364 ( .A(n40471), .B(n25452), .X(n25461) );
  nor_x1_sg U61365 ( .A(n40469), .B(n25731), .X(n25740) );
  nor_x1_sg U61366 ( .A(n26189), .B(n26284), .X(n26294) );
  nor_x1_sg U61367 ( .A(n40461), .B(n26568), .X(n26577) );
  nor_x1_sg U61368 ( .A(n40507), .B(n22929), .X(n22938) );
  nor_x1_sg U61369 ( .A(n40503), .B(n23206), .X(n23215) );
  nor_x1_sg U61370 ( .A(n23417), .B(n23486), .X(n23495) );
  nor_x1_sg U61371 ( .A(n23696), .B(n23765), .X(n23774) );
  nor_x1_sg U61372 ( .A(n40491), .B(n24044), .X(n24053) );
  nor_x1_sg U61373 ( .A(n40488), .B(n24323), .X(n24332) );
  nor_x1_sg U61374 ( .A(n40483), .B(n24602), .X(n24611) );
  nor_x1_sg U61375 ( .A(n40480), .B(n24880), .X(n24889) );
  nor_x1_sg U61376 ( .A(n40477), .B(n25159), .X(n25168) );
  nor_x1_sg U61377 ( .A(n40472), .B(n25438), .X(n25447) );
  nor_x1_sg U61378 ( .A(n25648), .B(n25717), .X(n25726) );
  nor_x1_sg U61379 ( .A(n26189), .B(n26268), .X(n26278) );
  nor_x1_sg U61380 ( .A(n26485), .B(n26554), .X(n26563) );
  nor_x1_sg U61381 ( .A(n26022), .B(n50546), .X(n26021) );
  inv_x1_sg U61382 ( .A(n42147), .X(n50546) );
  nor_x1_sg U61383 ( .A(n26024), .B(n50525), .X(n26022) );
  nor_x1_sg U61384 ( .A(n16822), .B(n50499), .X(n26024) );
  nand_x1_sg U61385 ( .A(n42312), .B(n22691), .X(n22689) );
  nand_x1_sg U61386 ( .A(n39667), .B(n26309), .X(n26307) );
  nor_x1_sg U61387 ( .A(n40509), .B(n22915), .X(n22924) );
  nor_x1_sg U61388 ( .A(n40505), .B(n23192), .X(n23201) );
  nor_x1_sg U61389 ( .A(n40501), .B(n23472), .X(n23481) );
  nor_x1_sg U61390 ( .A(n40497), .B(n23751), .X(n23760) );
  nor_x1_sg U61391 ( .A(n40493), .B(n24030), .X(n24039) );
  nor_x1_sg U61392 ( .A(n40489), .B(n24309), .X(n24318) );
  nor_x1_sg U61393 ( .A(n40485), .B(n24588), .X(n24597) );
  nor_x1_sg U61394 ( .A(n40481), .B(n24866), .X(n24875) );
  nor_x1_sg U61395 ( .A(n40475), .B(n25145), .X(n25154) );
  nor_x1_sg U61396 ( .A(n40472), .B(n25424), .X(n25433) );
  nor_x1_sg U61397 ( .A(n40469), .B(n25703), .X(n25712) );
  nor_x1_sg U61398 ( .A(n40464), .B(n26252), .X(n26262) );
  nor_x1_sg U61399 ( .A(n40459), .B(n26540), .X(n26549) );
  nor_x1_sg U61400 ( .A(n39482), .B(n42236), .X(n25974) );
  nor_x1_sg U61401 ( .A(n41297), .B(n39775), .X(n26000) );
  nand_x1_sg U61402 ( .A(n50390), .B(n17221), .X(n17254) );
  nand_x1_sg U61403 ( .A(n50372), .B(n39319), .X(n17253) );
  inv_x1_sg U61404 ( .A(n42302), .X(n45922) );
  inv_x1_sg U61405 ( .A(n42298), .X(n45925) );
  inv_x1_sg U61406 ( .A(n42285), .X(n45928) );
  nand_x1_sg U61407 ( .A(n50362), .B(n40074), .X(n17001) );
  nand_x1_sg U61408 ( .A(n41599), .B(n38729), .X(n7222) );
  nand_x1_sg U61409 ( .A(n7206), .B(n7207), .X(n7223) );
  nand_x1_sg U61410 ( .A(n41602), .B(n38731), .X(n8041) );
  nand_x1_sg U61411 ( .A(n8025), .B(n8026), .X(n8042) );
  nand_x1_sg U61412 ( .A(n41597), .B(n38733), .X(n8859) );
  nand_x1_sg U61413 ( .A(n8843), .B(n8844), .X(n8860) );
  nand_x1_sg U61414 ( .A(n41596), .B(n38735), .X(n9679) );
  nand_x1_sg U61415 ( .A(n9663), .B(n9664), .X(n9680) );
  nand_x1_sg U61416 ( .A(n41595), .B(n38737), .X(n10498) );
  nand_x1_sg U61417 ( .A(n10482), .B(n10483), .X(n10499) );
  nand_x1_sg U61418 ( .A(n41594), .B(n38739), .X(n11317) );
  nand_x1_sg U61419 ( .A(n11301), .B(n11302), .X(n11318) );
  nand_x1_sg U61420 ( .A(n41593), .B(n38741), .X(n12136) );
  nand_x1_sg U61421 ( .A(n12120), .B(n12121), .X(n12137) );
  nand_x1_sg U61422 ( .A(n41592), .B(n38743), .X(n12955) );
  nand_x1_sg U61423 ( .A(n12939), .B(n12940), .X(n12956) );
  nand_x1_sg U61424 ( .A(n41591), .B(n38745), .X(n13774) );
  nand_x1_sg U61425 ( .A(n13758), .B(n13759), .X(n13775) );
  nand_x1_sg U61426 ( .A(n41590), .B(n38747), .X(n14593) );
  nand_x1_sg U61427 ( .A(n14577), .B(n14578), .X(n14594) );
  nand_x1_sg U61428 ( .A(n41601), .B(n38749), .X(n15412) );
  nand_x1_sg U61429 ( .A(n15396), .B(n15397), .X(n15413) );
  nand_x1_sg U61430 ( .A(n41589), .B(n38751), .X(n16231) );
  nand_x1_sg U61431 ( .A(n16215), .B(n16216), .X(n16232) );
  nand_x1_sg U61432 ( .A(n41600), .B(n38753), .X(n17869) );
  nand_x1_sg U61433 ( .A(n17853), .B(n17854), .X(n17870) );
  nand_x1_sg U61434 ( .A(n41588), .B(n38755), .X(n18690) );
  nand_x1_sg U61435 ( .A(n18674), .B(n18675), .X(n18691) );
  nand_x1_sg U61436 ( .A(n39809), .B(n41692), .X(n7504) );
  nand_x1_sg U61437 ( .A(n39812), .B(n41665), .X(n8322) );
  nand_x1_sg U61438 ( .A(n41888), .B(n41688), .X(n9140) );
  nand_x1_sg U61439 ( .A(n41877), .B(n41690), .X(n9960) );
  nand_x1_sg U61440 ( .A(n41897), .B(n41686), .X(n10779) );
  nand_x1_sg U61441 ( .A(n41886), .B(n41684), .X(n11598) );
  nand_x1_sg U61442 ( .A(n41883), .B(n41682), .X(n12417) );
  nand_x1_sg U61443 ( .A(n41895), .B(n41680), .X(n13236) );
  nand_x1_sg U61444 ( .A(n39839), .B(n41678), .X(n14055) );
  nand_x1_sg U61445 ( .A(n39843), .B(n41676), .X(n14874) );
  nand_x1_sg U61446 ( .A(n39848), .B(n41663), .X(n15693) );
  nand_x1_sg U61447 ( .A(n41894), .B(n41674), .X(n16512) );
  nand_x1_sg U61448 ( .A(n40609), .B(n41672), .X(n17329) );
  nand_x1_sg U61449 ( .A(n41890), .B(n41670), .X(n18150) );
  nand_x1_sg U61450 ( .A(n41891), .B(n41668), .X(n18971) );
  nand_x1_sg U61451 ( .A(n41598), .B(n38727), .X(n17047) );
  nand_x1_sg U61452 ( .A(n17031), .B(n17032), .X(n17048) );
  nor_x1_sg U61453 ( .A(n41539), .B(n38925), .X(n6002) );
  nor_x1_sg U61454 ( .A(n41534), .B(n41041), .X(n6701) );
  nor_x1_sg U61455 ( .A(n41536), .B(n41023), .X(n6724) );
  nand_x1_sg U61456 ( .A(n7552), .B(n46921), .X(n7549) );
  nand_x1_sg U61457 ( .A(n7551), .B(n46989), .X(n7550) );
  inv_x1_sg U61458 ( .A(n7552), .X(n46989) );
  nand_x1_sg U61459 ( .A(n17377), .B(n50354), .X(n17374) );
  nand_x1_sg U61460 ( .A(n17376), .B(n50419), .X(n17375) );
  inv_x1_sg U61461 ( .A(n17377), .X(n50419) );
  nor_x1_sg U61462 ( .A(n45881), .B(n41003), .X(n6702) );
  nor_x1_sg U61463 ( .A(n45878), .B(n40977), .X(n6729) );
  nand_x1_sg U61464 ( .A(n8369), .B(n47278), .X(n8368) );
  nand_x1_sg U61465 ( .A(n8370), .B(n47213), .X(n8367) );
  inv_x1_sg U61466 ( .A(n8370), .X(n47278) );
  nand_x1_sg U61467 ( .A(n9187), .B(n47563), .X(n9186) );
  nand_x1_sg U61468 ( .A(n9188), .B(n47498), .X(n9185) );
  inv_x1_sg U61469 ( .A(n9188), .X(n47563) );
  nand_x1_sg U61470 ( .A(n10007), .B(n47848), .X(n10006) );
  nand_x1_sg U61471 ( .A(n10008), .B(n47783), .X(n10005) );
  inv_x1_sg U61472 ( .A(n10008), .X(n47848) );
  nand_x1_sg U61473 ( .A(n10826), .B(n48133), .X(n10825) );
  nand_x1_sg U61474 ( .A(n10827), .B(n48068), .X(n10824) );
  inv_x1_sg U61475 ( .A(n10827), .X(n48133) );
  nand_x1_sg U61476 ( .A(n11645), .B(n48418), .X(n11644) );
  nand_x1_sg U61477 ( .A(n11646), .B(n48353), .X(n11643) );
  inv_x1_sg U61478 ( .A(n11646), .X(n48418) );
  nand_x1_sg U61479 ( .A(n12464), .B(n48703), .X(n12463) );
  nand_x1_sg U61480 ( .A(n12465), .B(n48638), .X(n12462) );
  inv_x1_sg U61481 ( .A(n12465), .X(n48703) );
  nand_x1_sg U61482 ( .A(n13283), .B(n48989), .X(n13282) );
  nand_x1_sg U61483 ( .A(n13284), .B(n48924), .X(n13281) );
  inv_x1_sg U61484 ( .A(n13284), .X(n48989) );
  nand_x1_sg U61485 ( .A(n14102), .B(n49276), .X(n14101) );
  nand_x1_sg U61486 ( .A(n14103), .B(n49211), .X(n14100) );
  inv_x1_sg U61487 ( .A(n14103), .X(n49276) );
  nand_x1_sg U61488 ( .A(n14921), .B(n49562), .X(n14920) );
  nand_x1_sg U61489 ( .A(n14922), .B(n49497), .X(n14919) );
  inv_x1_sg U61490 ( .A(n14922), .X(n49562) );
  nand_x1_sg U61491 ( .A(n15740), .B(n49848), .X(n15739) );
  nand_x1_sg U61492 ( .A(n15741), .B(n49783), .X(n15738) );
  inv_x1_sg U61493 ( .A(n15741), .X(n49848) );
  nand_x1_sg U61494 ( .A(n16559), .B(n50134), .X(n16558) );
  nand_x1_sg U61495 ( .A(n16560), .B(n50069), .X(n16557) );
  inv_x1_sg U61496 ( .A(n16560), .X(n50134) );
  nand_x1_sg U61497 ( .A(n18197), .B(n50708), .X(n18196) );
  nand_x1_sg U61498 ( .A(n18198), .B(n50643), .X(n18195) );
  inv_x1_sg U61499 ( .A(n18198), .X(n50708) );
  nand_x1_sg U61500 ( .A(n19018), .B(n50995), .X(n19017) );
  nand_x1_sg U61501 ( .A(n19019), .B(n50930), .X(n19016) );
  inv_x1_sg U61502 ( .A(n19019), .X(n50995) );
  nor_x1_sg U61503 ( .A(n47127), .B(n41305), .X(n22704) );
  nand_x1_sg U61504 ( .A(n8102), .B(n8103), .X(n8099) );
  nor_x1_sg U61505 ( .A(n8102), .B(n39366), .X(n8101) );
  nand_x1_sg U61506 ( .A(n8920), .B(n8921), .X(n8917) );
  nor_x1_sg U61507 ( .A(n8920), .B(n39368), .X(n8919) );
  nand_x1_sg U61508 ( .A(n9740), .B(n9741), .X(n9737) );
  nor_x1_sg U61509 ( .A(n9740), .B(n39370), .X(n9739) );
  nand_x1_sg U61510 ( .A(n10559), .B(n10560), .X(n10556) );
  nor_x1_sg U61511 ( .A(n10559), .B(n39372), .X(n10558) );
  nand_x1_sg U61512 ( .A(n11378), .B(n11379), .X(n11375) );
  nor_x1_sg U61513 ( .A(n11378), .B(n39374), .X(n11377) );
  nand_x1_sg U61514 ( .A(n12197), .B(n12198), .X(n12194) );
  nor_x1_sg U61515 ( .A(n12197), .B(n39376), .X(n12196) );
  nand_x1_sg U61516 ( .A(n13016), .B(n13017), .X(n13013) );
  nor_x1_sg U61517 ( .A(n13016), .B(n39378), .X(n13015) );
  nand_x1_sg U61518 ( .A(n13835), .B(n13836), .X(n13832) );
  nor_x1_sg U61519 ( .A(n13835), .B(n39380), .X(n13834) );
  nand_x1_sg U61520 ( .A(n14654), .B(n14655), .X(n14651) );
  nor_x1_sg U61521 ( .A(n14654), .B(n39382), .X(n14653) );
  nand_x1_sg U61522 ( .A(n15473), .B(n15474), .X(n15470) );
  nor_x1_sg U61523 ( .A(n15473), .B(n39384), .X(n15472) );
  nand_x1_sg U61524 ( .A(n16292), .B(n16293), .X(n16289) );
  nor_x1_sg U61525 ( .A(n16292), .B(n39386), .X(n16291) );
  nand_x1_sg U61526 ( .A(n17930), .B(n17931), .X(n17927) );
  nor_x1_sg U61527 ( .A(n17930), .B(n41755), .X(n17929) );
  nand_x1_sg U61528 ( .A(n18751), .B(n18752), .X(n18748) );
  nor_x1_sg U61529 ( .A(n18751), .B(n39388), .X(n18750) );
  nand_x1_sg U61530 ( .A(n8199), .B(n41602), .X(n8375) );
  nor_x1_sg U61531 ( .A(n40180), .B(n39893), .X(n8377) );
  nand_x1_sg U61532 ( .A(n9017), .B(n41597), .X(n9193) );
  nor_x1_sg U61533 ( .A(n40212), .B(n41687), .X(n9195) );
  nand_x1_sg U61534 ( .A(n9837), .B(n41596), .X(n10013) );
  nor_x1_sg U61535 ( .A(n40206), .B(n41689), .X(n10015) );
  nand_x1_sg U61536 ( .A(n10656), .B(n41595), .X(n10832) );
  nor_x1_sg U61537 ( .A(n40204), .B(n41685), .X(n10834) );
  nand_x1_sg U61538 ( .A(n11475), .B(n41594), .X(n11651) );
  nor_x1_sg U61539 ( .A(n40198), .B(n41683), .X(n11653) );
  nand_x1_sg U61540 ( .A(n12294), .B(n41593), .X(n12470) );
  nor_x1_sg U61541 ( .A(n40194), .B(n41681), .X(n12472) );
  nand_x1_sg U61542 ( .A(n13113), .B(n41592), .X(n13289) );
  nor_x1_sg U61543 ( .A(n41747), .B(n41679), .X(n13291) );
  nand_x1_sg U61544 ( .A(n13932), .B(n41591), .X(n14108) );
  nor_x1_sg U61545 ( .A(n40174), .B(n41677), .X(n14110) );
  nand_x1_sg U61546 ( .A(n14751), .B(n41590), .X(n14927) );
  nor_x1_sg U61547 ( .A(n41748), .B(n41675), .X(n14929) );
  nand_x1_sg U61548 ( .A(n15570), .B(n41601), .X(n15746) );
  nor_x1_sg U61549 ( .A(n40170), .B(n39897), .X(n15748) );
  nand_x1_sg U61550 ( .A(n16389), .B(n41589), .X(n16565) );
  nor_x1_sg U61551 ( .A(n40168), .B(n41673), .X(n16567) );
  nand_x1_sg U61552 ( .A(n17206), .B(n41598), .X(n17382) );
  nor_x1_sg U61553 ( .A(n41778), .B(n39885), .X(n17384) );
  nand_x1_sg U61554 ( .A(n18027), .B(n41600), .X(n18203) );
  nor_x1_sg U61555 ( .A(n40214), .B(n41669), .X(n18205) );
  nand_x1_sg U61556 ( .A(n18848), .B(n41588), .X(n19024) );
  nor_x1_sg U61557 ( .A(n40182), .B(n41667), .X(n19026) );
  nand_x1_sg U61558 ( .A(n7381), .B(n41599), .X(n7557) );
  nor_x1_sg U61559 ( .A(n40085), .B(n39854), .X(n7559) );
  nand_x1_sg U61560 ( .A(n7624), .B(n39663), .X(n7623) );
  nand_x1_sg U61561 ( .A(n7625), .B(n7626), .X(n7622) );
  nor_x1_sg U61562 ( .A(n7625), .B(n40614), .X(n7624) );
  nand_x1_sg U61563 ( .A(n8442), .B(n8292), .X(n8441) );
  nand_x1_sg U61564 ( .A(n8443), .B(n8444), .X(n8440) );
  nor_x1_sg U61565 ( .A(n8443), .B(n40559), .X(n8442) );
  nand_x1_sg U61566 ( .A(n9260), .B(n9110), .X(n9259) );
  nand_x1_sg U61567 ( .A(n9261), .B(n9262), .X(n9258) );
  nor_x1_sg U61568 ( .A(n9261), .B(n40557), .X(n9260) );
  nand_x1_sg U61569 ( .A(n10080), .B(n9930), .X(n10079) );
  nand_x1_sg U61570 ( .A(n10081), .B(n10082), .X(n10078) );
  nor_x1_sg U61571 ( .A(n10081), .B(n40551), .X(n10080) );
  nand_x1_sg U61572 ( .A(n10899), .B(n10749), .X(n10898) );
  nand_x1_sg U61573 ( .A(n10900), .B(n10901), .X(n10897) );
  nor_x1_sg U61574 ( .A(n10900), .B(n40549), .X(n10899) );
  nand_x1_sg U61575 ( .A(n11718), .B(n11568), .X(n11717) );
  nand_x1_sg U61576 ( .A(n11719), .B(n11720), .X(n11716) );
  nor_x1_sg U61577 ( .A(n11719), .B(n40545), .X(n11718) );
  nand_x1_sg U61578 ( .A(n12537), .B(n12387), .X(n12536) );
  nand_x1_sg U61579 ( .A(n12538), .B(n12539), .X(n12535) );
  nor_x1_sg U61580 ( .A(n12538), .B(n40540), .X(n12537) );
  nand_x1_sg U61581 ( .A(n13356), .B(n13206), .X(n13355) );
  nand_x1_sg U61582 ( .A(n13357), .B(n13358), .X(n13354) );
  nor_x1_sg U61583 ( .A(n13357), .B(n40536), .X(n13356) );
  nand_x1_sg U61584 ( .A(n14175), .B(n14025), .X(n14174) );
  nand_x1_sg U61585 ( .A(n14176), .B(n14177), .X(n14173) );
  nor_x1_sg U61586 ( .A(n14176), .B(n13384), .X(n14175) );
  nand_x1_sg U61587 ( .A(n14994), .B(n14844), .X(n14993) );
  nand_x1_sg U61588 ( .A(n14995), .B(n14996), .X(n14992) );
  nor_x1_sg U61589 ( .A(n14995), .B(n40529), .X(n14994) );
  nand_x1_sg U61590 ( .A(n15813), .B(n15663), .X(n15812) );
  nand_x1_sg U61591 ( .A(n15814), .B(n15815), .X(n15811) );
  nor_x1_sg U61592 ( .A(n15814), .B(n40525), .X(n15813) );
  nand_x1_sg U61593 ( .A(n16632), .B(n16482), .X(n16631) );
  nand_x1_sg U61594 ( .A(n16633), .B(n16634), .X(n16630) );
  nor_x1_sg U61595 ( .A(n16633), .B(n40521), .X(n16632) );
  nand_x1_sg U61596 ( .A(n18270), .B(n18120), .X(n18269) );
  nand_x1_sg U61597 ( .A(n18271), .B(n18272), .X(n18268) );
  nor_x1_sg U61598 ( .A(n18271), .B(n40515), .X(n18270) );
  nand_x1_sg U61599 ( .A(n19091), .B(n18941), .X(n19090) );
  nand_x1_sg U61600 ( .A(n19092), .B(n19093), .X(n19089) );
  nor_x1_sg U61601 ( .A(n19092), .B(n40512), .X(n19091) );
  nand_x1_sg U61602 ( .A(n17450), .B(n17451), .X(n17447) );
  nor_x1_sg U61603 ( .A(n17450), .B(n40302), .X(n17449) );
  nand_x1_sg U61604 ( .A(n7637), .B(n7636), .X(n7634) );
  nor_x1_sg U61605 ( .A(n7636), .B(n7637), .X(n7635) );
  nand_x1_sg U61606 ( .A(n8455), .B(n8454), .X(n8452) );
  nor_x1_sg U61607 ( .A(n8454), .B(n8455), .X(n8453) );
  nand_x1_sg U61608 ( .A(n9273), .B(n9272), .X(n9270) );
  nor_x1_sg U61609 ( .A(n9272), .B(n9273), .X(n9271) );
  nand_x1_sg U61610 ( .A(n10093), .B(n10092), .X(n10090) );
  nor_x1_sg U61611 ( .A(n10092), .B(n10093), .X(n10091) );
  nand_x1_sg U61612 ( .A(n10912), .B(n10911), .X(n10909) );
  nor_x1_sg U61613 ( .A(n10911), .B(n10912), .X(n10910) );
  nand_x1_sg U61614 ( .A(n11731), .B(n11730), .X(n11728) );
  nor_x1_sg U61615 ( .A(n11730), .B(n11731), .X(n11729) );
  nand_x1_sg U61616 ( .A(n12550), .B(n12549), .X(n12547) );
  nor_x1_sg U61617 ( .A(n12549), .B(n12550), .X(n12548) );
  nand_x1_sg U61618 ( .A(n13369), .B(n13368), .X(n13366) );
  nor_x1_sg U61619 ( .A(n13368), .B(n13369), .X(n13367) );
  nand_x1_sg U61620 ( .A(n14188), .B(n14187), .X(n14185) );
  nor_x1_sg U61621 ( .A(n14187), .B(n14188), .X(n14186) );
  nand_x1_sg U61622 ( .A(n15007), .B(n15006), .X(n15004) );
  nor_x1_sg U61623 ( .A(n15006), .B(n15007), .X(n15005) );
  nand_x1_sg U61624 ( .A(n15826), .B(n15825), .X(n15823) );
  nor_x1_sg U61625 ( .A(n15825), .B(n15826), .X(n15824) );
  nand_x1_sg U61626 ( .A(n16645), .B(n16644), .X(n16642) );
  nor_x1_sg U61627 ( .A(n16644), .B(n16645), .X(n16643) );
  nand_x1_sg U61628 ( .A(n17462), .B(n17461), .X(n17459) );
  nor_x1_sg U61629 ( .A(n17461), .B(n17462), .X(n17460) );
  nand_x1_sg U61630 ( .A(n18283), .B(n18282), .X(n18280) );
  nor_x1_sg U61631 ( .A(n18282), .B(n18283), .X(n18281) );
  nand_x1_sg U61632 ( .A(n19104), .B(n19103), .X(n19101) );
  nor_x1_sg U61633 ( .A(n19103), .B(n19104), .X(n19102) );
  nand_x1_sg U61634 ( .A(n39809), .B(n46871), .X(n7066) );
  nand_x1_sg U61635 ( .A(n39813), .B(n47164), .X(n7884) );
  nand_x1_sg U61636 ( .A(n39831), .B(n47449), .X(n8702) );
  nand_x1_sg U61637 ( .A(n39845), .B(n47734), .X(n9522) );
  nand_x1_sg U61638 ( .A(n39815), .B(n48019), .X(n10341) );
  nand_x1_sg U61639 ( .A(n41885), .B(n48304), .X(n11160) );
  nand_x1_sg U61640 ( .A(n39836), .B(n48589), .X(n11979) );
  nand_x1_sg U61641 ( .A(n39818), .B(n48875), .X(n12798) );
  nand_x1_sg U61642 ( .A(n41881), .B(n49162), .X(n13617) );
  nand_x1_sg U61643 ( .A(n39842), .B(n49448), .X(n14436) );
  nand_x1_sg U61644 ( .A(n41876), .B(n49733), .X(n15255) );
  nand_x1_sg U61645 ( .A(n41893), .B(n50020), .X(n16074) );
  nand_x1_sg U61646 ( .A(n39828), .B(n50594), .X(n17712) );
  nand_x1_sg U61647 ( .A(n39824), .B(n50881), .X(n18533) );
  nand_x1_sg U61648 ( .A(n47032), .B(n7608), .X(n7596) );
  nand_x1_sg U61649 ( .A(n47319), .B(n8426), .X(n8414) );
  nand_x1_sg U61650 ( .A(n47604), .B(n9244), .X(n9232) );
  nand_x1_sg U61651 ( .A(n47889), .B(n10064), .X(n10052) );
  nand_x1_sg U61652 ( .A(n48174), .B(n10883), .X(n10871) );
  nand_x1_sg U61653 ( .A(n48459), .B(n11702), .X(n11690) );
  nand_x1_sg U61654 ( .A(n48744), .B(n12521), .X(n12509) );
  nand_x1_sg U61655 ( .A(n49030), .B(n13340), .X(n13328) );
  nand_x1_sg U61656 ( .A(n49317), .B(n14159), .X(n14147) );
  nand_x1_sg U61657 ( .A(n49603), .B(n14978), .X(n14966) );
  nand_x1_sg U61658 ( .A(n49889), .B(n15797), .X(n15785) );
  nand_x1_sg U61659 ( .A(n50175), .B(n16616), .X(n16604) );
  nand_x1_sg U61660 ( .A(n50460), .B(n17433), .X(n17421) );
  nand_x1_sg U61661 ( .A(n50749), .B(n18254), .X(n18242) );
  nand_x1_sg U61662 ( .A(n51036), .B(n19075), .X(n19063) );
  inv_x1_sg U61663 ( .A(n7174), .X(n46950) );
  inv_x1_sg U61664 ( .A(n7993), .X(n47241) );
  inv_x1_sg U61665 ( .A(n8811), .X(n47526) );
  inv_x1_sg U61666 ( .A(n9631), .X(n47811) );
  inv_x1_sg U61667 ( .A(n10450), .X(n48096) );
  inv_x1_sg U61668 ( .A(n11269), .X(n48381) );
  inv_x1_sg U61669 ( .A(n12088), .X(n48666) );
  inv_x1_sg U61670 ( .A(n12907), .X(n48952) );
  inv_x1_sg U61671 ( .A(n13726), .X(n49239) );
  inv_x1_sg U61672 ( .A(n14545), .X(n49525) );
  inv_x1_sg U61673 ( .A(n15364), .X(n49811) );
  inv_x1_sg U61674 ( .A(n16183), .X(n50097) );
  inv_x1_sg U61675 ( .A(n17821), .X(n50671) );
  inv_x1_sg U61676 ( .A(n18642), .X(n50958) );
  nand_x1_sg U61677 ( .A(n40610), .B(n50305), .X(n16893) );
  nand_x1_sg U61678 ( .A(n16678), .B(n16676), .X(n16894) );
  nand_x1_sg U61679 ( .A(n7207), .B(n46926), .X(n7204) );
  nand_x1_sg U61680 ( .A(n46889), .B(n7206), .X(n7205) );
  inv_x1_sg U61681 ( .A(n7206), .X(n46926) );
  nand_x1_sg U61682 ( .A(n8026), .B(n47218), .X(n8023) );
  nand_x1_sg U61683 ( .A(n47182), .B(n8025), .X(n8024) );
  inv_x1_sg U61684 ( .A(n8025), .X(n47218) );
  nand_x1_sg U61685 ( .A(n8844), .B(n47503), .X(n8841) );
  nand_x1_sg U61686 ( .A(n47467), .B(n8843), .X(n8842) );
  inv_x1_sg U61687 ( .A(n8843), .X(n47503) );
  nand_x1_sg U61688 ( .A(n9664), .B(n47788), .X(n9661) );
  nand_x1_sg U61689 ( .A(n47752), .B(n9663), .X(n9662) );
  inv_x1_sg U61690 ( .A(n9663), .X(n47788) );
  nand_x1_sg U61691 ( .A(n10483), .B(n48073), .X(n10480) );
  nand_x1_sg U61692 ( .A(n48037), .B(n10482), .X(n10481) );
  inv_x1_sg U61693 ( .A(n10482), .X(n48073) );
  nand_x1_sg U61694 ( .A(n11302), .B(n48358), .X(n11299) );
  nand_x1_sg U61695 ( .A(n48322), .B(n11301), .X(n11300) );
  inv_x1_sg U61696 ( .A(n11301), .X(n48358) );
  nand_x1_sg U61697 ( .A(n12121), .B(n48643), .X(n12118) );
  nand_x1_sg U61698 ( .A(n48607), .B(n12120), .X(n12119) );
  inv_x1_sg U61699 ( .A(n12120), .X(n48643) );
  nand_x1_sg U61700 ( .A(n12940), .B(n48929), .X(n12937) );
  nand_x1_sg U61701 ( .A(n48893), .B(n12939), .X(n12938) );
  inv_x1_sg U61702 ( .A(n12939), .X(n48929) );
  nand_x1_sg U61703 ( .A(n13759), .B(n49216), .X(n13756) );
  nand_x1_sg U61704 ( .A(n49180), .B(n13758), .X(n13757) );
  inv_x1_sg U61705 ( .A(n13758), .X(n49216) );
  nand_x1_sg U61706 ( .A(n14578), .B(n49502), .X(n14575) );
  nand_x1_sg U61707 ( .A(n49466), .B(n14577), .X(n14576) );
  inv_x1_sg U61708 ( .A(n14577), .X(n49502) );
  nand_x1_sg U61709 ( .A(n15397), .B(n49788), .X(n15394) );
  nand_x1_sg U61710 ( .A(n49751), .B(n15396), .X(n15395) );
  inv_x1_sg U61711 ( .A(n15396), .X(n49788) );
  nand_x1_sg U61712 ( .A(n16216), .B(n50074), .X(n16213) );
  nand_x1_sg U61713 ( .A(n50038), .B(n16215), .X(n16214) );
  inv_x1_sg U61714 ( .A(n16215), .X(n50074) );
  nand_x1_sg U61715 ( .A(n17032), .B(n50359), .X(n17029) );
  nand_x1_sg U61716 ( .A(n50323), .B(n17031), .X(n17030) );
  inv_x1_sg U61717 ( .A(n17031), .X(n50359) );
  nand_x1_sg U61718 ( .A(n17854), .B(n50648), .X(n17851) );
  nand_x1_sg U61719 ( .A(n50612), .B(n17853), .X(n17852) );
  inv_x1_sg U61720 ( .A(n17853), .X(n50648) );
  nand_x1_sg U61721 ( .A(n18675), .B(n50935), .X(n18672) );
  nand_x1_sg U61722 ( .A(n50899), .B(n18674), .X(n18673) );
  inv_x1_sg U61723 ( .A(n18674), .X(n50935) );
  nand_x1_sg U61724 ( .A(n17206), .B(n39319), .X(n17313) );
  nand_x1_sg U61725 ( .A(n41899), .B(n39519), .X(n8215) );
  nand_x1_sg U61726 ( .A(n41888), .B(n39518), .X(n9033) );
  nand_x1_sg U61727 ( .A(n39845), .B(n39524), .X(n9853) );
  nand_x1_sg U61728 ( .A(n41897), .B(n39523), .X(n10672) );
  nand_x1_sg U61729 ( .A(n39833), .B(n39522), .X(n11491) );
  nand_x1_sg U61730 ( .A(n41883), .B(n39521), .X(n12310) );
  nand_x1_sg U61731 ( .A(n39819), .B(n39528), .X(n13129) );
  nand_x1_sg U61732 ( .A(n39839), .B(n39527), .X(n13948) );
  nand_x1_sg U61733 ( .A(n41879), .B(n39526), .X(n14767) );
  nand_x1_sg U61734 ( .A(n41875), .B(n39525), .X(n15586) );
  nand_x1_sg U61735 ( .A(n41893), .B(n39531), .X(n16405) );
  nand_x1_sg U61736 ( .A(n40611), .B(n39520), .X(n17222) );
  nand_x1_sg U61737 ( .A(n41890), .B(n39530), .X(n18043) );
  nand_x1_sg U61738 ( .A(n39825), .B(n39529), .X(n18864) );
  nand_x1_sg U61739 ( .A(n41899), .B(n39506), .X(n8411) );
  nand_x1_sg U61740 ( .A(n41887), .B(n39505), .X(n9229) );
  nand_x1_sg U61741 ( .A(n41877), .B(n39507), .X(n10049) );
  nand_x1_sg U61742 ( .A(n39815), .B(n39509), .X(n10868) );
  nand_x1_sg U61743 ( .A(n41885), .B(n39508), .X(n11687) );
  nand_x1_sg U61744 ( .A(n41884), .B(n39511), .X(n12506) );
  nand_x1_sg U61745 ( .A(n41895), .B(n39510), .X(n13325) );
  nand_x1_sg U61746 ( .A(n41881), .B(n39513), .X(n14144) );
  nand_x1_sg U61747 ( .A(n39843), .B(n39512), .X(n14963) );
  nand_x1_sg U61748 ( .A(n39848), .B(n39515), .X(n15782) );
  nand_x1_sg U61749 ( .A(n39822), .B(n39514), .X(n16601) );
  nand_x1_sg U61750 ( .A(n41889), .B(n39516), .X(n18239) );
  nand_x1_sg U61751 ( .A(n41891), .B(n39517), .X(n19060) );
  nand_x1_sg U61752 ( .A(n7305), .B(n7561), .X(n7560) );
  nor_x1_sg U61753 ( .A(n7561), .B(n7305), .X(n7562) );
  nand_x1_sg U61754 ( .A(n8123), .B(n8379), .X(n8378) );
  nor_x1_sg U61755 ( .A(n8379), .B(n8123), .X(n8380) );
  nand_x1_sg U61756 ( .A(n8941), .B(n9197), .X(n9196) );
  nor_x1_sg U61757 ( .A(n9197), .B(n8941), .X(n9198) );
  nand_x1_sg U61758 ( .A(n9761), .B(n10017), .X(n10016) );
  nor_x1_sg U61759 ( .A(n10017), .B(n9761), .X(n10018) );
  nand_x1_sg U61760 ( .A(n10580), .B(n10836), .X(n10835) );
  nor_x1_sg U61761 ( .A(n10836), .B(n10580), .X(n10837) );
  nand_x1_sg U61762 ( .A(n11399), .B(n11655), .X(n11654) );
  nor_x1_sg U61763 ( .A(n11655), .B(n11399), .X(n11656) );
  nand_x1_sg U61764 ( .A(n12218), .B(n12474), .X(n12473) );
  nor_x1_sg U61765 ( .A(n12474), .B(n12218), .X(n12475) );
  nand_x1_sg U61766 ( .A(n13037), .B(n13293), .X(n13292) );
  nor_x1_sg U61767 ( .A(n13293), .B(n13037), .X(n13294) );
  nand_x1_sg U61768 ( .A(n13856), .B(n14112), .X(n14111) );
  nor_x1_sg U61769 ( .A(n14112), .B(n13856), .X(n14113) );
  nand_x1_sg U61770 ( .A(n14675), .B(n14931), .X(n14930) );
  nor_x1_sg U61771 ( .A(n14931), .B(n14675), .X(n14932) );
  nand_x1_sg U61772 ( .A(n15494), .B(n15750), .X(n15749) );
  nor_x1_sg U61773 ( .A(n15750), .B(n15494), .X(n15751) );
  nand_x1_sg U61774 ( .A(n16313), .B(n16569), .X(n16568) );
  nor_x1_sg U61775 ( .A(n16569), .B(n16313), .X(n16570) );
  nand_x1_sg U61776 ( .A(n17951), .B(n18207), .X(n18206) );
  nor_x1_sg U61777 ( .A(n18207), .B(n17951), .X(n18208) );
  nand_x1_sg U61778 ( .A(n18772), .B(n19028), .X(n19027) );
  nor_x1_sg U61779 ( .A(n19028), .B(n18772), .X(n19029) );
  nand_x1_sg U61780 ( .A(n7256), .B(n7257), .X(n7255) );
  nor_x1_sg U61781 ( .A(n7257), .B(n7256), .X(n7258) );
  nand_x1_sg U61782 ( .A(n47021), .B(n7494), .X(n7493) );
  nor_x1_sg U61783 ( .A(n7494), .B(n47021), .X(n7495) );
  nand_x1_sg U61784 ( .A(n8075), .B(n8076), .X(n8074) );
  nor_x1_sg U61785 ( .A(n8076), .B(n8075), .X(n8077) );
  nand_x1_sg U61786 ( .A(n47309), .B(n8312), .X(n8311) );
  nor_x1_sg U61787 ( .A(n8312), .B(n47309), .X(n8313) );
  nand_x1_sg U61788 ( .A(n8893), .B(n8894), .X(n8892) );
  nor_x1_sg U61789 ( .A(n8894), .B(n8893), .X(n8895) );
  nand_x1_sg U61790 ( .A(n47594), .B(n9130), .X(n9129) );
  nor_x1_sg U61791 ( .A(n9130), .B(n47594), .X(n9131) );
  nand_x1_sg U61792 ( .A(n9713), .B(n9714), .X(n9712) );
  nor_x1_sg U61793 ( .A(n9714), .B(n9713), .X(n9715) );
  nand_x1_sg U61794 ( .A(n47879), .B(n9950), .X(n9949) );
  nor_x1_sg U61795 ( .A(n9950), .B(n47879), .X(n9951) );
  nand_x1_sg U61796 ( .A(n10532), .B(n10533), .X(n10531) );
  nor_x1_sg U61797 ( .A(n10533), .B(n10532), .X(n10534) );
  nand_x1_sg U61798 ( .A(n48164), .B(n10769), .X(n10768) );
  nor_x1_sg U61799 ( .A(n10769), .B(n48164), .X(n10770) );
  nand_x1_sg U61800 ( .A(n11351), .B(n11352), .X(n11350) );
  nor_x1_sg U61801 ( .A(n11352), .B(n11351), .X(n11353) );
  nand_x1_sg U61802 ( .A(n48449), .B(n11588), .X(n11587) );
  nor_x1_sg U61803 ( .A(n11588), .B(n48449), .X(n11589) );
  nand_x1_sg U61804 ( .A(n12170), .B(n12171), .X(n12169) );
  nor_x1_sg U61805 ( .A(n12171), .B(n12170), .X(n12172) );
  nand_x1_sg U61806 ( .A(n48734), .B(n12407), .X(n12406) );
  nor_x1_sg U61807 ( .A(n12407), .B(n48734), .X(n12408) );
  nand_x1_sg U61808 ( .A(n12989), .B(n12990), .X(n12988) );
  nor_x1_sg U61809 ( .A(n12990), .B(n12989), .X(n12991) );
  nand_x1_sg U61810 ( .A(n49020), .B(n13226), .X(n13225) );
  nor_x1_sg U61811 ( .A(n13226), .B(n49020), .X(n13227) );
  nand_x1_sg U61812 ( .A(n13808), .B(n13809), .X(n13807) );
  nor_x1_sg U61813 ( .A(n13809), .B(n13808), .X(n13810) );
  nand_x1_sg U61814 ( .A(n49307), .B(n14045), .X(n14044) );
  nor_x1_sg U61815 ( .A(n14045), .B(n49307), .X(n14046) );
  nand_x1_sg U61816 ( .A(n14627), .B(n14628), .X(n14626) );
  nor_x1_sg U61817 ( .A(n14628), .B(n14627), .X(n14629) );
  nand_x1_sg U61818 ( .A(n49593), .B(n14864), .X(n14863) );
  nor_x1_sg U61819 ( .A(n14864), .B(n49593), .X(n14865) );
  nand_x1_sg U61820 ( .A(n15446), .B(n15447), .X(n15445) );
  nor_x1_sg U61821 ( .A(n15447), .B(n15446), .X(n15448) );
  nand_x1_sg U61822 ( .A(n49879), .B(n15683), .X(n15682) );
  nor_x1_sg U61823 ( .A(n15683), .B(n49879), .X(n15684) );
  nand_x1_sg U61824 ( .A(n16265), .B(n16266), .X(n16264) );
  nor_x1_sg U61825 ( .A(n16266), .B(n16265), .X(n16267) );
  nand_x1_sg U61826 ( .A(n50165), .B(n16502), .X(n16501) );
  nor_x1_sg U61827 ( .A(n16502), .B(n50165), .X(n16503) );
  nand_x1_sg U61828 ( .A(n17081), .B(n17082), .X(n17080) );
  nor_x1_sg U61829 ( .A(n17082), .B(n17081), .X(n17083) );
  nand_x1_sg U61830 ( .A(n50450), .B(n17319), .X(n17318) );
  nor_x1_sg U61831 ( .A(n17319), .B(n50450), .X(n17320) );
  nand_x1_sg U61832 ( .A(n17903), .B(n17904), .X(n17902) );
  nor_x1_sg U61833 ( .A(n17904), .B(n17903), .X(n17905) );
  nand_x1_sg U61834 ( .A(n50739), .B(n42019), .X(n18139) );
  nor_x1_sg U61835 ( .A(n42019), .B(n50739), .X(n18141) );
  nand_x1_sg U61836 ( .A(n18724), .B(n18725), .X(n18723) );
  nor_x1_sg U61837 ( .A(n18725), .B(n18724), .X(n18726) );
  nand_x1_sg U61838 ( .A(n51026), .B(n18961), .X(n18960) );
  nor_x1_sg U61839 ( .A(n18961), .B(n51026), .X(n18962) );
  nand_x1_sg U61840 ( .A(n7131), .B(n7132), .X(n7130) );
  nor_x1_sg U61841 ( .A(n7132), .B(n7131), .X(n7133) );
  nand_x1_sg U61842 ( .A(n7949), .B(n7950), .X(n7948) );
  nor_x1_sg U61843 ( .A(n7950), .B(n7949), .X(n7951) );
  nand_x1_sg U61844 ( .A(n8767), .B(n8768), .X(n8766) );
  nor_x1_sg U61845 ( .A(n8768), .B(n8767), .X(n8769) );
  nand_x1_sg U61846 ( .A(n9587), .B(n9588), .X(n9586) );
  nor_x1_sg U61847 ( .A(n9588), .B(n9587), .X(n9589) );
  nand_x1_sg U61848 ( .A(n10406), .B(n10407), .X(n10405) );
  nor_x1_sg U61849 ( .A(n10407), .B(n10406), .X(n10408) );
  nand_x1_sg U61850 ( .A(n11225), .B(n11226), .X(n11224) );
  nor_x1_sg U61851 ( .A(n11226), .B(n11225), .X(n11227) );
  nand_x1_sg U61852 ( .A(n12044), .B(n12045), .X(n12043) );
  nor_x1_sg U61853 ( .A(n12045), .B(n12044), .X(n12046) );
  nand_x1_sg U61854 ( .A(n12863), .B(n12864), .X(n12862) );
  nor_x1_sg U61855 ( .A(n12864), .B(n12863), .X(n12865) );
  nand_x1_sg U61856 ( .A(n13682), .B(n13683), .X(n13681) );
  nor_x1_sg U61857 ( .A(n13683), .B(n13682), .X(n13684) );
  nand_x1_sg U61858 ( .A(n14501), .B(n14502), .X(n14500) );
  nor_x1_sg U61859 ( .A(n14502), .B(n14501), .X(n14503) );
  nand_x1_sg U61860 ( .A(n15320), .B(n15321), .X(n15319) );
  nor_x1_sg U61861 ( .A(n15321), .B(n15320), .X(n15322) );
  nand_x1_sg U61862 ( .A(n16139), .B(n16140), .X(n16138) );
  nor_x1_sg U61863 ( .A(n16140), .B(n16139), .X(n16141) );
  nand_x1_sg U61864 ( .A(n16956), .B(n16957), .X(n16955) );
  nor_x1_sg U61865 ( .A(n16957), .B(n16956), .X(n16958) );
  nand_x1_sg U61866 ( .A(n17777), .B(n17778), .X(n17776) );
  nor_x1_sg U61867 ( .A(n17778), .B(n17777), .X(n17779) );
  nand_x1_sg U61868 ( .A(n18598), .B(n18599), .X(n18597) );
  nor_x1_sg U61869 ( .A(n18599), .B(n18598), .X(n18600) );
  nand_x1_sg U61870 ( .A(n17127), .B(n17128), .X(n17126) );
  nor_x1_sg U61871 ( .A(n17128), .B(n17127), .X(n17129) );
  nor_x1_sg U61872 ( .A(n7809), .B(n41915), .X(n7807) );
  nor_x1_sg U61873 ( .A(n8627), .B(n41916), .X(n8625) );
  nor_x1_sg U61874 ( .A(n9447), .B(n41907), .X(n9445) );
  nor_x1_sg U61875 ( .A(n10266), .B(n41909), .X(n10264) );
  nor_x1_sg U61876 ( .A(n11085), .B(n41913), .X(n11083) );
  nor_x1_sg U61877 ( .A(n11904), .B(n41914), .X(n11902) );
  nor_x1_sg U61878 ( .A(n12723), .B(n41908), .X(n12721) );
  nor_x1_sg U61879 ( .A(n13542), .B(n41911), .X(n13540) );
  nor_x1_sg U61880 ( .A(n14361), .B(n41917), .X(n14359) );
  nor_x1_sg U61881 ( .A(n15180), .B(n41904), .X(n15178) );
  nor_x1_sg U61882 ( .A(n15999), .B(n41905), .X(n15997) );
  nor_x1_sg U61883 ( .A(n18458), .B(n41906), .X(n18456) );
  nor_x1_sg U61884 ( .A(n16816), .B(n41860), .X(n16814) );
  nor_x1_sg U61885 ( .A(n17637), .B(n41912), .X(n17635) );
  nor_x1_sg U61886 ( .A(n6992), .B(n41861), .X(n6990) );
  nand_x1_sg U61887 ( .A(n39804), .B(n40082), .X(n7612) );
  nand_x1_sg U61888 ( .A(n39933), .B(n40076), .X(n17437) );
  nand_x1_sg U61889 ( .A(n42306), .B(n24638), .X(n24636) );
  nand_x1_sg U61890 ( .A(n8432), .B(n8354), .X(n8427) );
  nor_x1_sg U61891 ( .A(n40560), .B(n41712), .X(n8432) );
  nand_x1_sg U61892 ( .A(n9250), .B(n9172), .X(n9245) );
  nor_x1_sg U61893 ( .A(n8469), .B(n41711), .X(n9250) );
  nand_x1_sg U61894 ( .A(n10070), .B(n9992), .X(n10065) );
  nor_x1_sg U61895 ( .A(n40552), .B(n41714), .X(n10070) );
  nand_x1_sg U61896 ( .A(n10889), .B(n10811), .X(n10884) );
  nor_x1_sg U61897 ( .A(n10108), .B(n41713), .X(n10889) );
  nand_x1_sg U61898 ( .A(n11708), .B(n11630), .X(n11703) );
  nor_x1_sg U61899 ( .A(n10927), .B(n41716), .X(n11708) );
  nand_x1_sg U61900 ( .A(n12527), .B(n12449), .X(n12522) );
  nor_x1_sg U61901 ( .A(n11746), .B(n41715), .X(n12527) );
  nand_x1_sg U61902 ( .A(n13346), .B(n13268), .X(n13341) );
  nor_x1_sg U61903 ( .A(n12565), .B(n41718), .X(n13346) );
  nand_x1_sg U61904 ( .A(n14165), .B(n14087), .X(n14160) );
  nor_x1_sg U61905 ( .A(n40533), .B(n41717), .X(n14165) );
  nand_x1_sg U61906 ( .A(n14984), .B(n14906), .X(n14979) );
  nor_x1_sg U61907 ( .A(n14203), .B(n41720), .X(n14984) );
  nand_x1_sg U61908 ( .A(n15803), .B(n15725), .X(n15798) );
  nor_x1_sg U61909 ( .A(n15022), .B(n41719), .X(n15803) );
  nand_x1_sg U61910 ( .A(n16622), .B(n16544), .X(n16617) );
  nor_x1_sg U61911 ( .A(n15841), .B(n41722), .X(n16622) );
  nand_x1_sg U61912 ( .A(n18260), .B(n18182), .X(n18255) );
  nor_x1_sg U61913 ( .A(n40516), .B(n41721), .X(n18260) );
  nand_x1_sg U61914 ( .A(n19081), .B(n19003), .X(n19076) );
  nor_x1_sg U61915 ( .A(n18300), .B(n41723), .X(n19081) );
  nand_x1_sg U61916 ( .A(n40081), .B(n7324), .X(n7317) );
  nand_x1_sg U61917 ( .A(n40078), .B(n17149), .X(n17142) );
  nand_x1_sg U61918 ( .A(n7614), .B(n7536), .X(n7609) );
  nor_x1_sg U61919 ( .A(n40613), .B(n41710), .X(n7614) );
  nand_x1_sg U61920 ( .A(n17439), .B(n17361), .X(n17434) );
  nor_x1_sg U61921 ( .A(n40301), .B(n41724), .X(n17439) );
  nand_x1_sg U61922 ( .A(n39852), .B(n39805), .X(n7592) );
  nand_x4_sg U61923 ( .A(n26312), .B(n41308), .X(n26310) );
  nor_x1_sg U61924 ( .A(n26313), .B(n26314), .X(n26312) );
  nor_x1_sg U61925 ( .A(n26315), .B(n40463), .X(n26313) );
  nor_x1_sg U61926 ( .A(n39244), .B(n18279), .X(n26314) );
  nand_x1_sg U61927 ( .A(n40072), .B(n39520), .X(n17386) );
  nor_x1_sg U61928 ( .A(n7438), .B(n40615), .X(n7437) );
  nor_x1_sg U61929 ( .A(n40367), .B(n39606), .X(n7438) );
  nor_x1_sg U61930 ( .A(n17263), .B(n40303), .X(n17262) );
  nor_x1_sg U61931 ( .A(n40310), .B(n39603), .X(n17263) );
  nand_x1_sg U61932 ( .A(n39810), .B(n39772), .X(n7397) );
  nand_x1_sg U61933 ( .A(n41902), .B(n39804), .X(n7377) );
  nand_x1_sg U61934 ( .A(n41899), .B(n39939), .X(n8195) );
  nand_x1_sg U61935 ( .A(n39830), .B(n39941), .X(n9013) );
  nand_x1_sg U61936 ( .A(n39845), .B(n39943), .X(n9833) );
  nand_x1_sg U61937 ( .A(n41898), .B(n39958), .X(n10652) );
  nand_x1_sg U61938 ( .A(n41885), .B(n39960), .X(n11471) );
  nand_x1_sg U61939 ( .A(n39837), .B(n39950), .X(n12290) );
  nand_x1_sg U61940 ( .A(n41896), .B(n39952), .X(n13109) );
  nand_x1_sg U61941 ( .A(n41882), .B(n39954), .X(n13928) );
  nand_x1_sg U61942 ( .A(n39842), .B(n39948), .X(n14747) );
  nand_x1_sg U61943 ( .A(n41875), .B(n39944), .X(n15566) );
  nand_x1_sg U61944 ( .A(n41894), .B(n39946), .X(n16385) );
  nand_x1_sg U61945 ( .A(n41889), .B(n39935), .X(n18023) );
  nand_x1_sg U61946 ( .A(n41892), .B(n39937), .X(n18844) );
  inv_x1_sg U61947 ( .A(n7102), .X(n46856) );
  inv_x1_sg U61948 ( .A(n7920), .X(n47149) );
  inv_x1_sg U61949 ( .A(n8738), .X(n47434) );
  inv_x1_sg U61950 ( .A(n9558), .X(n47719) );
  inv_x1_sg U61951 ( .A(n10377), .X(n48004) );
  inv_x1_sg U61952 ( .A(n11196), .X(n48289) );
  inv_x1_sg U61953 ( .A(n12015), .X(n48574) );
  inv_x1_sg U61954 ( .A(n12834), .X(n48860) );
  inv_x1_sg U61955 ( .A(n13653), .X(n49147) );
  inv_x1_sg U61956 ( .A(n14472), .X(n49433) );
  inv_x1_sg U61957 ( .A(n15291), .X(n49718) );
  inv_x1_sg U61958 ( .A(n16110), .X(n50005) );
  inv_x1_sg U61959 ( .A(n17748), .X(n50579) );
  inv_x1_sg U61960 ( .A(n18569), .X(n50866) );
  inv_x1_sg U61961 ( .A(n7079), .X(n46854) );
  inv_x1_sg U61962 ( .A(n7897), .X(n47147) );
  inv_x1_sg U61963 ( .A(n8715), .X(n47432) );
  inv_x1_sg U61964 ( .A(n9535), .X(n47717) );
  inv_x1_sg U61965 ( .A(n10354), .X(n48002) );
  inv_x1_sg U61966 ( .A(n11173), .X(n48287) );
  inv_x1_sg U61967 ( .A(n11992), .X(n48572) );
  inv_x1_sg U61968 ( .A(n12811), .X(n48858) );
  inv_x1_sg U61969 ( .A(n13630), .X(n49145) );
  inv_x1_sg U61970 ( .A(n14449), .X(n49431) );
  inv_x1_sg U61971 ( .A(n15268), .X(n49716) );
  inv_x1_sg U61972 ( .A(n16087), .X(n50003) );
  inv_x1_sg U61973 ( .A(n17725), .X(n50577) );
  inv_x1_sg U61974 ( .A(n18546), .X(n50864) );
  nor_x1_sg U61975 ( .A(n22894), .B(n22895), .X(n22893) );
  nor_x1_sg U61976 ( .A(n22897), .B(n41400), .X(n22892) );
  nor_x1_sg U61977 ( .A(n22860), .B(n22896), .X(n22895) );
  nor_x1_sg U61978 ( .A(n23157), .B(n23158), .X(n23156) );
  nor_x1_sg U61979 ( .A(n23160), .B(n41399), .X(n23155) );
  nor_x1_sg U61980 ( .A(n23137), .B(n23159), .X(n23158) );
  nor_x1_sg U61981 ( .A(n23423), .B(n23424), .X(n23422) );
  nor_x1_sg U61982 ( .A(n23426), .B(n40017), .X(n23421) );
  nor_x1_sg U61983 ( .A(n40499), .B(n23425), .X(n23424) );
  nor_x1_sg U61984 ( .A(n23444), .B(n23445), .X(n23443) );
  nor_x1_sg U61985 ( .A(n23447), .B(n41404), .X(n23442) );
  nor_x1_sg U61986 ( .A(n39713), .B(n23446), .X(n23445) );
  nor_x1_sg U61987 ( .A(n23730), .B(n23731), .X(n23729) );
  nor_x1_sg U61988 ( .A(n23733), .B(n41405), .X(n23728) );
  nor_x1_sg U61989 ( .A(n40496), .B(n23732), .X(n23731) );
  nor_x1_sg U61990 ( .A(n23995), .B(n23996), .X(n23994) );
  nor_x1_sg U61991 ( .A(n23998), .B(n39154), .X(n23993) );
  nor_x1_sg U61992 ( .A(n40492), .B(n23997), .X(n23996) );
  nor_x1_sg U61993 ( .A(n24260), .B(n24261), .X(n24259) );
  nor_x1_sg U61994 ( .A(n24263), .B(n39654), .X(n24258) );
  nor_x1_sg U61995 ( .A(n24254), .B(n24262), .X(n24261) );
  nor_x1_sg U61996 ( .A(n24281), .B(n24282), .X(n24280) );
  nor_x1_sg U61997 ( .A(n24284), .B(n39437), .X(n24279) );
  nor_x1_sg U61998 ( .A(n41792), .B(n24283), .X(n24282) );
  nor_x1_sg U61999 ( .A(n24567), .B(n24568), .X(n24566) );
  nor_x1_sg U62000 ( .A(n24570), .B(n40455), .X(n24565) );
  nor_x1_sg U62001 ( .A(n24533), .B(n24569), .X(n24568) );
  nor_x1_sg U62002 ( .A(n24831), .B(n24832), .X(n24830) );
  nor_x1_sg U62003 ( .A(n24834), .B(n40375), .X(n24829) );
  nor_x1_sg U62004 ( .A(n40479), .B(n24833), .X(n24832) );
  nor_x1_sg U62005 ( .A(n25096), .B(n25097), .X(n25095) );
  nor_x1_sg U62006 ( .A(n25099), .B(n39654), .X(n25094) );
  nor_x1_sg U62007 ( .A(n40476), .B(n25098), .X(n25097) );
  nor_x1_sg U62008 ( .A(n25117), .B(n25118), .X(n25116) );
  nor_x1_sg U62009 ( .A(n25120), .B(n39155), .X(n25115) );
  nor_x1_sg U62010 ( .A(n39695), .B(n25119), .X(n25118) );
  nor_x1_sg U62011 ( .A(n25403), .B(n25404), .X(n25402) );
  nor_x1_sg U62012 ( .A(n25406), .B(n40020), .X(n25401) );
  nor_x1_sg U62013 ( .A(n25369), .B(n25405), .X(n25404) );
  nor_x1_sg U62014 ( .A(n25668), .B(n25669), .X(n25667) );
  nor_x1_sg U62015 ( .A(n25671), .B(n40017), .X(n25666) );
  nor_x1_sg U62016 ( .A(n40467), .B(n25670), .X(n25669) );
  nor_x1_sg U62017 ( .A(n26505), .B(n26506), .X(n26504) );
  nor_x1_sg U62018 ( .A(n26508), .B(n40457), .X(n26503) );
  nor_x1_sg U62019 ( .A(n26485), .B(n26507), .X(n26506) );
  nor_x1_sg U62020 ( .A(n22866), .B(n22867), .X(n22865) );
  nor_x1_sg U62021 ( .A(n22869), .B(n39653), .X(n22864) );
  nor_x1_sg U62022 ( .A(n40509), .B(n22868), .X(n22867) );
  nor_x1_sg U62023 ( .A(n22880), .B(n22881), .X(n22879) );
  nor_x1_sg U62024 ( .A(n22883), .B(n40454), .X(n22878) );
  nor_x1_sg U62025 ( .A(n40508), .B(n22882), .X(n22881) );
  nor_x1_sg U62026 ( .A(n22887), .B(n22888), .X(n22886) );
  nor_x1_sg U62027 ( .A(n22890), .B(n39274), .X(n22885) );
  nor_x1_sg U62028 ( .A(n41782), .B(n22889), .X(n22888) );
  nor_x1_sg U62029 ( .A(n23143), .B(n23144), .X(n23142) );
  nor_x1_sg U62030 ( .A(n23146), .B(n39436), .X(n23141) );
  nor_x1_sg U62031 ( .A(n40504), .B(n23145), .X(n23144) );
  nor_x1_sg U62032 ( .A(n23164), .B(n23165), .X(n23163) );
  nor_x1_sg U62033 ( .A(n23167), .B(n41408), .X(n23162) );
  nor_x1_sg U62034 ( .A(n39716), .B(n23166), .X(n23165) );
  nor_x1_sg U62035 ( .A(n23171), .B(n23172), .X(n23170) );
  nor_x1_sg U62036 ( .A(n23174), .B(n41310), .X(n23169) );
  nor_x1_sg U62037 ( .A(n40503), .B(n23173), .X(n23172) );
  nor_x1_sg U62038 ( .A(n23437), .B(n23438), .X(n23436) );
  nor_x1_sg U62039 ( .A(n23440), .B(n39437), .X(n23435) );
  nor_x1_sg U62040 ( .A(n40500), .B(n23439), .X(n23438) );
  nor_x1_sg U62041 ( .A(n23451), .B(n23452), .X(n23450) );
  nor_x1_sg U62042 ( .A(n23454), .B(n40373), .X(n23449) );
  nor_x1_sg U62043 ( .A(n40501), .B(n23453), .X(n23452) );
  nor_x1_sg U62044 ( .A(n23702), .B(n23703), .X(n23701) );
  nor_x1_sg U62045 ( .A(n23705), .B(n41405), .X(n23700) );
  nor_x1_sg U62046 ( .A(n23696), .B(n23704), .X(n23703) );
  nor_x1_sg U62047 ( .A(n23716), .B(n23717), .X(n23715) );
  nor_x1_sg U62048 ( .A(n23719), .B(n40373), .X(n23714) );
  nor_x1_sg U62049 ( .A(n40495), .B(n23718), .X(n23717) );
  nor_x1_sg U62050 ( .A(n23723), .B(n23724), .X(n23722) );
  nor_x1_sg U62051 ( .A(n23726), .B(n38816), .X(n23721) );
  nor_x1_sg U62052 ( .A(n39710), .B(n23725), .X(n23724) );
  nor_x1_sg U62053 ( .A(n23981), .B(n23982), .X(n23980) );
  nor_x1_sg U62054 ( .A(n23984), .B(n39152), .X(n23979) );
  nor_x1_sg U62055 ( .A(n40493), .B(n23983), .X(n23982) );
  nor_x1_sg U62056 ( .A(n24002), .B(n24003), .X(n24001) );
  nor_x1_sg U62057 ( .A(n24005), .B(n41408), .X(n24000) );
  nor_x1_sg U62058 ( .A(n41790), .B(n24004), .X(n24003) );
  nor_x1_sg U62059 ( .A(n24009), .B(n24010), .X(n24008) );
  nor_x1_sg U62060 ( .A(n24012), .B(n41403), .X(n24007) );
  nor_x1_sg U62061 ( .A(n23975), .B(n24011), .X(n24010) );
  nor_x1_sg U62062 ( .A(n24274), .B(n24275), .X(n24273) );
  nor_x1_sg U62063 ( .A(n24277), .B(n40016), .X(n24272) );
  nor_x1_sg U62064 ( .A(n24254), .B(n24276), .X(n24275) );
  nor_x1_sg U62065 ( .A(n24288), .B(n24289), .X(n24287) );
  nor_x1_sg U62066 ( .A(n24291), .B(n41403), .X(n24286) );
  nor_x1_sg U62067 ( .A(n40488), .B(n24290), .X(n24289) );
  nor_x1_sg U62068 ( .A(n24539), .B(n24540), .X(n24538) );
  nor_x1_sg U62069 ( .A(n24542), .B(n41466), .X(n24537) );
  nor_x1_sg U62070 ( .A(n40485), .B(n24541), .X(n24540) );
  nor_x1_sg U62071 ( .A(n24553), .B(n24554), .X(n24552) );
  nor_x1_sg U62072 ( .A(n24556), .B(n40371), .X(n24551) );
  nor_x1_sg U62073 ( .A(n40484), .B(n24555), .X(n24554) );
  nor_x1_sg U62074 ( .A(n24560), .B(n24561), .X(n24559) );
  nor_x1_sg U62075 ( .A(n24563), .B(n41399), .X(n24558) );
  nor_x1_sg U62076 ( .A(n39701), .B(n24562), .X(n24561) );
  nor_x1_sg U62077 ( .A(n24817), .B(n24818), .X(n24816) );
  nor_x1_sg U62078 ( .A(n24820), .B(n38981), .X(n24815) );
  nor_x1_sg U62079 ( .A(n40479), .B(n24819), .X(n24818) );
  nor_x1_sg U62080 ( .A(n24838), .B(n24839), .X(n24837) );
  nor_x1_sg U62081 ( .A(n24841), .B(n41402), .X(n24836) );
  nor_x1_sg U62082 ( .A(n41796), .B(n24840), .X(n24839) );
  nor_x1_sg U62083 ( .A(n24845), .B(n24846), .X(n24844) );
  nor_x1_sg U62084 ( .A(n24848), .B(n39437), .X(n24843) );
  nor_x1_sg U62085 ( .A(n24811), .B(n24847), .X(n24846) );
  nor_x1_sg U62086 ( .A(n25110), .B(n25111), .X(n25109) );
  nor_x1_sg U62087 ( .A(n25113), .B(n41468), .X(n25108) );
  nor_x1_sg U62088 ( .A(n40477), .B(n25112), .X(n25111) );
  nor_x1_sg U62089 ( .A(n25124), .B(n25125), .X(n25123) );
  nor_x1_sg U62090 ( .A(n25127), .B(n41468), .X(n25122) );
  nor_x1_sg U62091 ( .A(n40475), .B(n25126), .X(n25125) );
  nor_x1_sg U62092 ( .A(n25375), .B(n25376), .X(n25374) );
  nor_x1_sg U62093 ( .A(n25378), .B(n39152), .X(n25373) );
  nor_x1_sg U62094 ( .A(n40473), .B(n25377), .X(n25376) );
  nor_x1_sg U62095 ( .A(n25389), .B(n25390), .X(n25388) );
  nor_x1_sg U62096 ( .A(n25392), .B(n40374), .X(n25387) );
  nor_x1_sg U62097 ( .A(n25369), .B(n25391), .X(n25390) );
  nor_x1_sg U62098 ( .A(n25396), .B(n25397), .X(n25395) );
  nor_x1_sg U62099 ( .A(n25399), .B(n40375), .X(n25394) );
  nor_x1_sg U62100 ( .A(n39692), .B(n25398), .X(n25397) );
  nor_x1_sg U62101 ( .A(n25654), .B(n25655), .X(n25653) );
  nor_x1_sg U62102 ( .A(n25657), .B(n41408), .X(n25652) );
  nor_x1_sg U62103 ( .A(n25648), .B(n25656), .X(n25655) );
  nor_x1_sg U62104 ( .A(n25675), .B(n25676), .X(n25674) );
  nor_x1_sg U62105 ( .A(n25678), .B(n40012), .X(n25673) );
  nor_x1_sg U62106 ( .A(n39689), .B(n25677), .X(n25676) );
  nor_x1_sg U62107 ( .A(n25682), .B(n25683), .X(n25681) );
  nor_x1_sg U62108 ( .A(n25685), .B(n40019), .X(n25680) );
  nor_x1_sg U62109 ( .A(n40468), .B(n25684), .X(n25683) );
  nor_x1_sg U62110 ( .A(n26491), .B(n26492), .X(n26490) );
  nor_x1_sg U62111 ( .A(n26494), .B(n40376), .X(n26489) );
  nor_x1_sg U62112 ( .A(n40460), .B(n26493), .X(n26492) );
  nor_x1_sg U62113 ( .A(n26512), .B(n26513), .X(n26511) );
  nor_x1_sg U62114 ( .A(n26515), .B(n40373), .X(n26510) );
  nor_x1_sg U62115 ( .A(n39683), .B(n26514), .X(n26513) );
  nor_x1_sg U62116 ( .A(n26519), .B(n26520), .X(n26518) );
  nor_x1_sg U62117 ( .A(n26522), .B(n41405), .X(n26517) );
  nor_x1_sg U62118 ( .A(n40459), .B(n26521), .X(n26520) );
  inv_x1_sg U62119 ( .A(n16906), .X(n50286) );
  nand_x1_sg U62120 ( .A(n39850), .B(n39773), .X(n6969) );
  nor_x1_sg U62121 ( .A(n8256), .B(n40561), .X(n8255) );
  nor_x1_sg U62122 ( .A(n40307), .B(n41657), .X(n8256) );
  nor_x1_sg U62123 ( .A(n9074), .B(n40557), .X(n9073) );
  nor_x1_sg U62124 ( .A(n41844), .B(n41656), .X(n9074) );
  nor_x1_sg U62125 ( .A(n9894), .B(n40552), .X(n9893) );
  nor_x1_sg U62126 ( .A(n41852), .B(n41651), .X(n9894) );
  nor_x1_sg U62127 ( .A(n10713), .B(n40548), .X(n10712) );
  nor_x1_sg U62128 ( .A(n41854), .B(n39740), .X(n10713) );
  nor_x1_sg U62129 ( .A(n11532), .B(n10927), .X(n11531) );
  nor_x1_sg U62130 ( .A(n41850), .B(n41649), .X(n11532) );
  nor_x1_sg U62131 ( .A(n12351), .B(n11746), .X(n12350) );
  nor_x1_sg U62132 ( .A(n41856), .B(n41648), .X(n12351) );
  nor_x1_sg U62133 ( .A(n13170), .B(n40537), .X(n13169) );
  nor_x1_sg U62134 ( .A(n41858), .B(n41655), .X(n13170) );
  nor_x1_sg U62135 ( .A(n13989), .B(n40532), .X(n13988) );
  nor_x1_sg U62136 ( .A(n41848), .B(n41654), .X(n13989) );
  nor_x1_sg U62137 ( .A(n14808), .B(n40529), .X(n14807) );
  nor_x1_sg U62138 ( .A(n41759), .B(n39755), .X(n14808) );
  nor_x1_sg U62139 ( .A(n15627), .B(n40523), .X(n15626) );
  nor_x1_sg U62140 ( .A(n41846), .B(n41652), .X(n15627) );
  nor_x1_sg U62141 ( .A(n16446), .B(n15841), .X(n16445) );
  nor_x1_sg U62142 ( .A(n41764), .B(n41659), .X(n16446) );
  nor_x1_sg U62143 ( .A(n18084), .B(n40517), .X(n18083) );
  nor_x1_sg U62144 ( .A(n40363), .B(n39764), .X(n18084) );
  nor_x1_sg U62145 ( .A(n18905), .B(n18300), .X(n18904) );
  nor_x1_sg U62146 ( .A(n41762), .B(n39767), .X(n18905) );
  nand_x1_sg U62147 ( .A(n39938), .B(n40243), .X(n8121) );
  nand_x1_sg U62148 ( .A(n39940), .B(n40248), .X(n8939) );
  nand_x1_sg U62149 ( .A(n39942), .B(n40252), .X(n9759) );
  nand_x1_sg U62150 ( .A(n39959), .B(n40259), .X(n10578) );
  nand_x1_sg U62151 ( .A(n39960), .B(n40262), .X(n11397) );
  nand_x1_sg U62152 ( .A(n39951), .B(n40269), .X(n12216) );
  nand_x1_sg U62153 ( .A(n39953), .B(n40274), .X(n13035) );
  nand_x1_sg U62154 ( .A(n39955), .B(n40280), .X(n13854) );
  nand_x1_sg U62155 ( .A(n39948), .B(n40283), .X(n14673) );
  nand_x1_sg U62156 ( .A(n39945), .B(n40289), .X(n15492) );
  nand_x1_sg U62157 ( .A(n39947), .B(n40292), .X(n16311) );
  nand_x1_sg U62158 ( .A(n39934), .B(n40238), .X(n17949) );
  nand_x1_sg U62159 ( .A(n39936), .B(n40299), .X(n18770) );
  nand_x1_sg U62160 ( .A(n40610), .B(n39932), .X(n17202) );
  nand_x1_sg U62161 ( .A(n39805), .B(n40162), .X(n7303) );
  nor_x1_sg U62162 ( .A(n5940), .B(n5941), .X(n5939) );
  nor_x1_sg U62163 ( .A(n5919), .B(n5920), .X(n5918) );
  nor_x1_sg U62164 ( .A(n5848), .B(n5849), .X(n5847) );
  nor_x1_sg U62165 ( .A(n5889), .B(n5890), .X(n5888) );
  nor_x1_sg U62166 ( .A(n5926), .B(n5927), .X(n5925) );
  nor_x1_sg U62167 ( .A(n5839), .B(n5840), .X(n5838) );
  nor_x1_sg U62168 ( .A(n5903), .B(n5904), .X(n5902) );
  nor_x1_sg U62169 ( .A(n5896), .B(n5897), .X(n5895) );
  nor_x1_sg U62170 ( .A(n5784), .B(n5785), .X(n5783) );
  nor_x1_sg U62171 ( .A(n5855), .B(n5856), .X(n5854) );
  nor_x1_sg U62172 ( .A(n5910), .B(n5911), .X(n5909) );
  nor_x1_sg U62173 ( .A(n5871), .B(n5872), .X(n5870) );
  nor_x1_sg U62174 ( .A(n5794), .B(n5795), .X(n5793) );
  nor_x1_sg U62175 ( .A(n5817), .B(n5818), .X(n5816) );
  nor_x1_sg U62176 ( .A(n5810), .B(n5811), .X(n5809) );
  nor_x1_sg U62177 ( .A(n5880), .B(n5881), .X(n5879) );
  nor_x1_sg U62178 ( .A(n5803), .B(n5804), .X(n5802) );
  nor_x1_sg U62179 ( .A(n5824), .B(n5825), .X(n5823) );
  nor_x1_sg U62180 ( .A(n5947), .B(n5948), .X(n5946) );
  inv_x1_sg U62181 ( .A(n7551), .X(n46921) );
  inv_x1_sg U62182 ( .A(n17376), .X(n50354) );
  nand_x1_sg U62183 ( .A(n41106), .B(n44981), .X(n22553) );
  nand_x1_sg U62184 ( .A(n41094), .B(n44990), .X(n22554) );
  inv_x1_sg U62185 ( .A(n7444), .X(n46899) );
  inv_x1_sg U62186 ( .A(n17269), .X(n50332) );
  nor_x1_sg U62187 ( .A(n26773), .B(n26774), .X(n26759) );
  nor_x1_sg U62188 ( .A(n21784), .B(n21785), .X(n21772) );
  nand_x1_sg U62189 ( .A(n21776), .B(n21777), .X(n21775) );
  nor_x1_sg U62190 ( .A(n21924), .B(n21925), .X(n21912) );
  nand_x1_sg U62191 ( .A(n21916), .B(n21917), .X(n21915) );
  nor_x1_sg U62192 ( .A(n22064), .B(n22065), .X(n22052) );
  nand_x1_sg U62193 ( .A(n22056), .B(n22057), .X(n22055) );
  nor_x1_sg U62194 ( .A(n22205), .B(n22206), .X(n22193) );
  nand_x1_sg U62195 ( .A(n22197), .B(n22198), .X(n22196) );
  nor_x1_sg U62196 ( .A(n22348), .B(n22349), .X(n22336) );
  nand_x1_sg U62197 ( .A(n22340), .B(n22341), .X(n22339) );
  nor_x1_sg U62198 ( .A(n22488), .B(n22489), .X(n22477) );
  nand_x1_sg U62199 ( .A(n22481), .B(n22482), .X(n22480) );
  nand_x1_sg U62200 ( .A(n39806), .B(n26017), .X(n26015) );
  nor_x1_sg U62201 ( .A(n21737), .B(n21738), .X(n21725) );
  nand_x1_sg U62202 ( .A(n21729), .B(n21730), .X(n21728) );
  nor_x1_sg U62203 ( .A(n21831), .B(n21832), .X(n21819) );
  nand_x1_sg U62204 ( .A(n21823), .B(n21824), .X(n21822) );
  nor_x1_sg U62205 ( .A(n21878), .B(n21879), .X(n21866) );
  nand_x1_sg U62206 ( .A(n21870), .B(n21871), .X(n21869) );
  nor_x1_sg U62207 ( .A(n21971), .B(n21972), .X(n21959) );
  nand_x1_sg U62208 ( .A(n21963), .B(n21964), .X(n21962) );
  nor_x1_sg U62209 ( .A(n22017), .B(n22018), .X(n22005) );
  nand_x1_sg U62210 ( .A(n22009), .B(n22010), .X(n22008) );
  nor_x1_sg U62211 ( .A(n22110), .B(n22111), .X(n22098) );
  nand_x1_sg U62212 ( .A(n22102), .B(n22103), .X(n22101) );
  nor_x1_sg U62213 ( .A(n22158), .B(n22159), .X(n22146) );
  nand_x1_sg U62214 ( .A(n22150), .B(n22151), .X(n22149) );
  nor_x1_sg U62215 ( .A(n22253), .B(n22254), .X(n22241) );
  nand_x1_sg U62216 ( .A(n22245), .B(n22246), .X(n22244) );
  nor_x1_sg U62217 ( .A(n22300), .B(n22301), .X(n22288) );
  nand_x1_sg U62218 ( .A(n22292), .B(n22293), .X(n22291) );
  nor_x1_sg U62219 ( .A(n22395), .B(n22396), .X(n22383) );
  nand_x1_sg U62220 ( .A(n22387), .B(n22388), .X(n22386) );
  nor_x1_sg U62221 ( .A(n22442), .B(n22443), .X(n22431) );
  nand_x1_sg U62222 ( .A(n22435), .B(n22436), .X(n22434) );
  nor_x1_sg U62223 ( .A(n22531), .B(n22532), .X(n22523) );
  nand_x1_sg U62224 ( .A(n22527), .B(n22528), .X(n22526) );
  nand_x1_sg U62225 ( .A(n8162), .B(n8161), .X(n8159) );
  nor_x1_sg U62226 ( .A(n8161), .B(n8162), .X(n8160) );
  nand_x1_sg U62227 ( .A(n8980), .B(n8979), .X(n8977) );
  nor_x1_sg U62228 ( .A(n8979), .B(n8980), .X(n8978) );
  nand_x1_sg U62229 ( .A(n9800), .B(n9799), .X(n9797) );
  nor_x1_sg U62230 ( .A(n9799), .B(n9800), .X(n9798) );
  nand_x1_sg U62231 ( .A(n10619), .B(n10618), .X(n10616) );
  nor_x1_sg U62232 ( .A(n10618), .B(n10619), .X(n10617) );
  nand_x1_sg U62233 ( .A(n11438), .B(n11437), .X(n11435) );
  nor_x1_sg U62234 ( .A(n11437), .B(n11438), .X(n11436) );
  nand_x1_sg U62235 ( .A(n12257), .B(n12256), .X(n12254) );
  nor_x1_sg U62236 ( .A(n12256), .B(n12257), .X(n12255) );
  nand_x1_sg U62237 ( .A(n13076), .B(n13075), .X(n13073) );
  nor_x1_sg U62238 ( .A(n13075), .B(n13076), .X(n13074) );
  nand_x1_sg U62239 ( .A(n13895), .B(n13894), .X(n13892) );
  nor_x1_sg U62240 ( .A(n13894), .B(n13895), .X(n13893) );
  nand_x1_sg U62241 ( .A(n14714), .B(n14713), .X(n14711) );
  nor_x1_sg U62242 ( .A(n14713), .B(n14714), .X(n14712) );
  nand_x1_sg U62243 ( .A(n15533), .B(n15532), .X(n15530) );
  nor_x1_sg U62244 ( .A(n15532), .B(n15533), .X(n15531) );
  nand_x1_sg U62245 ( .A(n16352), .B(n16351), .X(n16349) );
  nor_x1_sg U62246 ( .A(n16351), .B(n16352), .X(n16350) );
  nand_x1_sg U62247 ( .A(n17169), .B(n17168), .X(n17166) );
  nor_x1_sg U62248 ( .A(n17168), .B(n17169), .X(n17167) );
  nand_x1_sg U62249 ( .A(n17990), .B(n17989), .X(n17987) );
  nor_x1_sg U62250 ( .A(n17989), .B(n17990), .X(n17988) );
  nand_x1_sg U62251 ( .A(n18811), .B(n18810), .X(n18808) );
  nor_x1_sg U62252 ( .A(n18810), .B(n18811), .X(n18809) );
  inv_x1_sg U62253 ( .A(n27987), .X(n45081) );
  nand_x1_sg U62254 ( .A(n7344), .B(n7343), .X(n7341) );
  nor_x1_sg U62255 ( .A(n7343), .B(n7344), .X(n7342) );
  nand_x2_sg U62256 ( .A(n6943), .B(n6944), .X(n6942) );
  inv_x1_sg U62257 ( .A(n42074), .X(n47061) );
  nand_x2_sg U62258 ( .A(n7760), .B(n7761), .X(n7759) );
  inv_x1_sg U62259 ( .A(n42073), .X(n47347) );
  nand_x2_sg U62260 ( .A(n8578), .B(n8579), .X(n8577) );
  inv_x1_sg U62261 ( .A(n42071), .X(n47632) );
  nand_x2_sg U62262 ( .A(n9398), .B(n9399), .X(n9397) );
  inv_x1_sg U62263 ( .A(n42070), .X(n47917) );
  nand_x2_sg U62264 ( .A(n10217), .B(n10218), .X(n10216) );
  inv_x1_sg U62265 ( .A(n42069), .X(n48202) );
  nand_x2_sg U62266 ( .A(n11036), .B(n11037), .X(n11035) );
  inv_x1_sg U62267 ( .A(n42068), .X(n48487) );
  nand_x2_sg U62268 ( .A(n11855), .B(n11856), .X(n11854) );
  inv_x1_sg U62269 ( .A(n42067), .X(n48772) );
  nand_x2_sg U62270 ( .A(n12674), .B(n12675), .X(n12673) );
  inv_x1_sg U62271 ( .A(n42066), .X(n49059) );
  nand_x2_sg U62272 ( .A(n13493), .B(n13494), .X(n13492) );
  inv_x1_sg U62273 ( .A(n42065), .X(n49345) );
  nand_x2_sg U62274 ( .A(n14312), .B(n14313), .X(n14311) );
  inv_x1_sg U62275 ( .A(n42064), .X(n49631) );
  nand_x2_sg U62276 ( .A(n15131), .B(n15132), .X(n15130) );
  inv_x1_sg U62277 ( .A(n42072), .X(n49917) );
  nand_x2_sg U62278 ( .A(n15950), .B(n15951), .X(n15949) );
  inv_x1_sg U62279 ( .A(n42063), .X(n50203) );
  nand_x2_sg U62280 ( .A(n16767), .B(n16768), .X(n16766) );
  inv_x1_sg U62281 ( .A(n42088), .X(n50488) );
  nand_x2_sg U62282 ( .A(n17588), .B(n17589), .X(n17587) );
  inv_x1_sg U62283 ( .A(n42062), .X(n50777) );
  nand_x2_sg U62284 ( .A(n18409), .B(n18410), .X(n18408) );
  inv_x1_sg U62285 ( .A(n42061), .X(n51064) );
  nand_x1_sg U62286 ( .A(n40073), .B(n39933), .X(n17316) );
  inv_x1_sg U62287 ( .A(n8262), .X(n47194) );
  inv_x1_sg U62288 ( .A(n9080), .X(n47479) );
  inv_x1_sg U62289 ( .A(n9900), .X(n47764) );
  inv_x1_sg U62290 ( .A(n10719), .X(n48049) );
  inv_x1_sg U62291 ( .A(n11538), .X(n48334) );
  inv_x1_sg U62292 ( .A(n12357), .X(n48619) );
  inv_x1_sg U62293 ( .A(n13176), .X(n48905) );
  inv_x1_sg U62294 ( .A(n13995), .X(n49192) );
  inv_x1_sg U62295 ( .A(n14814), .X(n49478) );
  inv_x1_sg U62296 ( .A(n15633), .X(n49764) );
  inv_x1_sg U62297 ( .A(n16452), .X(n50050) );
  inv_x1_sg U62298 ( .A(n18090), .X(n50624) );
  inv_x1_sg U62299 ( .A(n18911), .X(n50911) );
  nand_x1_sg U62300 ( .A(n40072), .B(n40609), .X(n17014) );
  nand_x1_sg U62301 ( .A(n47010), .B(n46899), .X(n7434) );
  nand_x1_sg U62302 ( .A(n47298), .B(n47194), .X(n8252) );
  nand_x1_sg U62303 ( .A(n47583), .B(n47479), .X(n9070) );
  nand_x1_sg U62304 ( .A(n47868), .B(n47764), .X(n9890) );
  nand_x1_sg U62305 ( .A(n48153), .B(n48049), .X(n10709) );
  nand_x1_sg U62306 ( .A(n48438), .B(n48334), .X(n11528) );
  nand_x1_sg U62307 ( .A(n48723), .B(n48619), .X(n12347) );
  nand_x1_sg U62308 ( .A(n49009), .B(n48905), .X(n13166) );
  nand_x1_sg U62309 ( .A(n49296), .B(n49192), .X(n13985) );
  nand_x1_sg U62310 ( .A(n49582), .B(n49478), .X(n14804) );
  nand_x1_sg U62311 ( .A(n49868), .B(n49764), .X(n15623) );
  nand_x1_sg U62312 ( .A(n50154), .B(n50050), .X(n16442) );
  nand_x1_sg U62313 ( .A(n50439), .B(n50332), .X(n17259) );
  nand_x1_sg U62314 ( .A(n50728), .B(n50624), .X(n18080) );
  nand_x1_sg U62315 ( .A(n51015), .B(n50911), .X(n18901) );
  nor_x1_sg U62316 ( .A(n7480), .B(n7481), .X(n7479) );
  nor_x1_sg U62317 ( .A(n8298), .B(n8299), .X(n8297) );
  nor_x1_sg U62318 ( .A(n9116), .B(n9117), .X(n9115) );
  nor_x1_sg U62319 ( .A(n9936), .B(n9937), .X(n9935) );
  nor_x1_sg U62320 ( .A(n10755), .B(n10756), .X(n10754) );
  nor_x1_sg U62321 ( .A(n11574), .B(n11575), .X(n11573) );
  nor_x1_sg U62322 ( .A(n12393), .B(n12394), .X(n12392) );
  nor_x1_sg U62323 ( .A(n13212), .B(n13213), .X(n13211) );
  nor_x1_sg U62324 ( .A(n14031), .B(n14032), .X(n14030) );
  nor_x1_sg U62325 ( .A(n14850), .B(n14851), .X(n14849) );
  nor_x1_sg U62326 ( .A(n15669), .B(n15670), .X(n15668) );
  nor_x1_sg U62327 ( .A(n16488), .B(n16489), .X(n16487) );
  nor_x1_sg U62328 ( .A(n17305), .B(n17306), .X(n17304) );
  nor_x1_sg U62329 ( .A(n18126), .B(n18127), .X(n18125) );
  nor_x1_sg U62330 ( .A(n18947), .B(n18948), .X(n18946) );
  nor_x1_sg U62331 ( .A(n22616), .B(n22617), .X(n22615) );
  nor_x1_sg U62332 ( .A(n22619), .B(n41409), .X(n22614) );
  nor_x1_sg U62333 ( .A(n41779), .B(n22618), .X(n22617) );
  nor_x1_sg U62334 ( .A(n22642), .B(n22643), .X(n22641) );
  nor_x1_sg U62335 ( .A(n22645), .B(n40374), .X(n22640) );
  nor_x1_sg U62336 ( .A(n39930), .B(n22644), .X(n22643) );
  nor_x1_sg U62337 ( .A(n26228), .B(n26229), .X(n26227) );
  nor_x1_sg U62338 ( .A(n26231), .B(n40014), .X(n26226) );
  nor_x1_sg U62339 ( .A(n40465), .B(n26230), .X(n26229) );
  nor_x1_sg U62340 ( .A(n22604), .B(n22605), .X(n22603) );
  nor_x1_sg U62341 ( .A(n22607), .B(n41403), .X(n22602) );
  nor_x1_sg U62342 ( .A(n40161), .B(n22606), .X(n22605) );
  nor_x1_sg U62343 ( .A(n22622), .B(n22623), .X(n22621) );
  nor_x1_sg U62344 ( .A(n22625), .B(n41402), .X(n22620) );
  nor_x1_sg U62345 ( .A(n41780), .B(n22624), .X(n22623) );
  nor_x1_sg U62346 ( .A(n22628), .B(n22629), .X(n22627) );
  nor_x1_sg U62347 ( .A(n22631), .B(n40370), .X(n22626) );
  nor_x1_sg U62348 ( .A(n41861), .B(n22630), .X(n22629) );
  nor_x1_sg U62349 ( .A(n22653), .B(n47132), .X(n22652) );
  nor_x1_sg U62350 ( .A(n22657), .B(n40018), .X(n22651) );
  inv_x1_sg U62351 ( .A(n22654), .X(n47132) );
  nor_x1_sg U62352 ( .A(n25939), .B(n25940), .X(n25938) );
  nor_x1_sg U62353 ( .A(n25942), .B(n40374), .X(n25937) );
  nor_x1_sg U62354 ( .A(n41778), .B(n25941), .X(n25940) );
  nor_x1_sg U62355 ( .A(n25951), .B(n25952), .X(n25950) );
  nor_x1_sg U62356 ( .A(n25954), .B(n41402), .X(n25949) );
  nor_x1_sg U62357 ( .A(n41860), .B(n25953), .X(n25952) );
  nor_x1_sg U62358 ( .A(n5747), .B(n26027), .X(n26026) );
  nor_x1_sg U62359 ( .A(n26030), .B(n39155), .X(n26025) );
  nor_x1_sg U62360 ( .A(n50555), .B(n26028), .X(n26027) );
  nor_x1_sg U62361 ( .A(n26196), .B(n26197), .X(n26195) );
  nor_x1_sg U62362 ( .A(n26199), .B(n40020), .X(n26194) );
  nor_x1_sg U62363 ( .A(n40465), .B(n26198), .X(n26197) );
  nor_x1_sg U62364 ( .A(n26212), .B(n26213), .X(n26211) );
  nor_x1_sg U62365 ( .A(n26215), .B(n40017), .X(n26210) );
  nor_x1_sg U62366 ( .A(n40464), .B(n26214), .X(n26213) );
  nor_x1_sg U62367 ( .A(n26220), .B(n26221), .X(n26219) );
  nor_x1_sg U62368 ( .A(n26223), .B(n38816), .X(n26218) );
  nor_x1_sg U62369 ( .A(n39686), .B(n26222), .X(n26221) );
  nand_x1_sg U62370 ( .A(n39939), .B(n8389), .X(n8388) );
  nand_x1_sg U62371 ( .A(n47367), .B(n39548), .X(n8387) );
  nand_x1_sg U62372 ( .A(n39941), .B(n9207), .X(n9206) );
  nand_x1_sg U62373 ( .A(n47652), .B(n39549), .X(n9205) );
  nand_x1_sg U62374 ( .A(n39943), .B(n10027), .X(n10026) );
  nand_x1_sg U62375 ( .A(n47937), .B(n39550), .X(n10025) );
  nand_x1_sg U62376 ( .A(n39959), .B(n10846), .X(n10845) );
  nand_x1_sg U62377 ( .A(n48222), .B(n39557), .X(n10844) );
  nand_x1_sg U62378 ( .A(n39961), .B(n11665), .X(n11664) );
  nand_x1_sg U62379 ( .A(n48507), .B(n39558), .X(n11663) );
  nand_x1_sg U62380 ( .A(n39951), .B(n12484), .X(n12483) );
  nand_x1_sg U62381 ( .A(n48792), .B(n39554), .X(n12482) );
  nand_x1_sg U62382 ( .A(n39953), .B(n13303), .X(n13302) );
  nand_x1_sg U62383 ( .A(n49079), .B(n39555), .X(n13301) );
  nand_x1_sg U62384 ( .A(n39955), .B(n14122), .X(n14121) );
  nand_x1_sg U62385 ( .A(n49365), .B(n39556), .X(n14120) );
  nand_x1_sg U62386 ( .A(n39949), .B(n14941), .X(n14940) );
  nand_x1_sg U62387 ( .A(n49651), .B(n39553), .X(n14939) );
  nand_x1_sg U62388 ( .A(n39945), .B(n15760), .X(n15759) );
  nand_x1_sg U62389 ( .A(n49937), .B(n39551), .X(n15758) );
  nand_x1_sg U62390 ( .A(n39947), .B(n16579), .X(n16578) );
  nand_x1_sg U62391 ( .A(n50223), .B(n39552), .X(n16577) );
  nand_x1_sg U62392 ( .A(n39932), .B(n17396), .X(n17395) );
  nand_x1_sg U62393 ( .A(n50508), .B(n39545), .X(n17394) );
  nand_x1_sg U62394 ( .A(n39935), .B(n18217), .X(n18216) );
  nand_x1_sg U62395 ( .A(n50797), .B(n39546), .X(n18215) );
  nand_x1_sg U62396 ( .A(n39937), .B(n19038), .X(n19037) );
  nand_x1_sg U62397 ( .A(n51084), .B(n39547), .X(n19036) );
  nor_x1_sg U62398 ( .A(n39473), .B(n5771), .X(\L1_0/n4432 ) );
  nor_x1_sg U62399 ( .A(n41320), .B(n5788), .X(\L1_0/n4428 ) );
  nor_x1_sg U62400 ( .A(n39473), .B(n5913), .X(\L1_0/n4424 ) );
  nor_x1_sg U62401 ( .A(n39125), .B(n5865), .X(\L1_0/n4420 ) );
  nor_x1_sg U62402 ( .A(n41320), .B(n5842), .X(\L1_0/n4416 ) );
  nor_x1_sg U62403 ( .A(n41279), .B(n5773), .X(\L1_0/n4412 ) );
  nor_x1_sg U62404 ( .A(n41320), .B(n5786), .X(n5123) );
  nor_x1_sg U62405 ( .A(n38946), .B(n5874), .X(\L1_0/n4404 ) );
  nor_x1_sg U62406 ( .A(n39925), .B(n5829), .X(\L1_0/n4400 ) );
  nor_x1_sg U62407 ( .A(n39924), .B(n5777), .X(\L1_0/n4396 ) );
  nor_x1_sg U62408 ( .A(n41321), .B(n5863), .X(\L1_0/n4392 ) );
  nor_x1_sg U62409 ( .A(n41574), .B(n5827), .X(\L1_0/n4388 ) );
  nor_x1_sg U62410 ( .A(n39473), .B(n5775), .X(\L1_0/n4384 ) );
  nor_x1_sg U62411 ( .A(n39925), .B(n5833), .X(\L1_0/n4380 ) );
  nor_x1_sg U62412 ( .A(n41323), .B(n5883), .X(\L1_0/n4376 ) );
  nor_x1_sg U62413 ( .A(n38946), .B(n5950), .X(\L1_0/n4372 ) );
  nor_x1_sg U62414 ( .A(n41322), .B(n5797), .X(\L1_0/n4368 ) );
  nor_x1_sg U62415 ( .A(n41323), .B(n5831), .X(\L1_0/n4364 ) );
  nand_x1_sg U62416 ( .A(n47081), .B(n39726), .X(n7569) );
  nand_x1_sg U62417 ( .A(n39804), .B(n7571), .X(n7570) );
  nand_x1_sg U62418 ( .A(n7468), .B(n7469), .X(n7466) );
  nor_x1_sg U62419 ( .A(n7468), .B(n7469), .X(n7467) );
  nand_x1_sg U62420 ( .A(n17293), .B(n17294), .X(n17291) );
  nor_x1_sg U62421 ( .A(n17293), .B(n17294), .X(n17292) );
  nand_x1_sg U62422 ( .A(n8286), .B(n8287), .X(n8284) );
  nor_x1_sg U62423 ( .A(n8286), .B(n8287), .X(n8285) );
  nand_x1_sg U62424 ( .A(n9104), .B(n9105), .X(n9102) );
  nor_x1_sg U62425 ( .A(n9104), .B(n9105), .X(n9103) );
  nand_x1_sg U62426 ( .A(n9924), .B(n9925), .X(n9922) );
  nor_x1_sg U62427 ( .A(n9924), .B(n9925), .X(n9923) );
  nand_x1_sg U62428 ( .A(n10743), .B(n10744), .X(n10741) );
  nor_x1_sg U62429 ( .A(n10743), .B(n10744), .X(n10742) );
  nand_x1_sg U62430 ( .A(n11562), .B(n11563), .X(n11560) );
  nor_x1_sg U62431 ( .A(n11562), .B(n11563), .X(n11561) );
  nand_x1_sg U62432 ( .A(n12381), .B(n12382), .X(n12379) );
  nor_x1_sg U62433 ( .A(n12381), .B(n12382), .X(n12380) );
  nand_x1_sg U62434 ( .A(n13200), .B(n13201), .X(n13198) );
  nor_x1_sg U62435 ( .A(n13200), .B(n13201), .X(n13199) );
  nand_x1_sg U62436 ( .A(n14019), .B(n14020), .X(n14017) );
  nor_x1_sg U62437 ( .A(n14019), .B(n14020), .X(n14018) );
  nand_x1_sg U62438 ( .A(n14838), .B(n14839), .X(n14836) );
  nor_x1_sg U62439 ( .A(n14838), .B(n14839), .X(n14837) );
  nand_x1_sg U62440 ( .A(n15657), .B(n15658), .X(n15655) );
  nor_x1_sg U62441 ( .A(n15657), .B(n15658), .X(n15656) );
  nand_x1_sg U62442 ( .A(n16476), .B(n16477), .X(n16474) );
  nor_x1_sg U62443 ( .A(n16476), .B(n16477), .X(n16475) );
  nand_x1_sg U62444 ( .A(n18114), .B(n18115), .X(n18112) );
  nor_x1_sg U62445 ( .A(n18114), .B(n18115), .X(n18113) );
  nand_x1_sg U62446 ( .A(n18935), .B(n18936), .X(n18933) );
  nor_x1_sg U62447 ( .A(n18935), .B(n18936), .X(n18934) );
  inv_x1_sg U62448 ( .A(n7108), .X(n46864) );
  inv_x1_sg U62449 ( .A(n7926), .X(n47157) );
  inv_x1_sg U62450 ( .A(n8744), .X(n47442) );
  inv_x1_sg U62451 ( .A(n9564), .X(n47727) );
  inv_x1_sg U62452 ( .A(n10383), .X(n48012) );
  inv_x1_sg U62453 ( .A(n11202), .X(n48297) );
  inv_x1_sg U62454 ( .A(n12021), .X(n48582) );
  inv_x1_sg U62455 ( .A(n12840), .X(n48868) );
  inv_x1_sg U62456 ( .A(n13659), .X(n49155) );
  inv_x1_sg U62457 ( .A(n14478), .X(n49441) );
  inv_x1_sg U62458 ( .A(n15297), .X(n49726) );
  inv_x1_sg U62459 ( .A(n16116), .X(n50013) );
  inv_x1_sg U62460 ( .A(n16933), .X(n50297) );
  inv_x1_sg U62461 ( .A(n17754), .X(n50587) );
  inv_x1_sg U62462 ( .A(n18575), .X(n50874) );
  nand_x1_sg U62463 ( .A(n8052), .B(n47245), .X(n8058) );
  nand_x1_sg U62464 ( .A(n8870), .B(n47530), .X(n8876) );
  nand_x1_sg U62465 ( .A(n9690), .B(n47815), .X(n9696) );
  nand_x1_sg U62466 ( .A(n10509), .B(n48100), .X(n10515) );
  nand_x1_sg U62467 ( .A(n11328), .B(n48385), .X(n11334) );
  nand_x1_sg U62468 ( .A(n12147), .B(n48670), .X(n12153) );
  nand_x1_sg U62469 ( .A(n12966), .B(n48956), .X(n12972) );
  nand_x1_sg U62470 ( .A(n13785), .B(n49243), .X(n13791) );
  nand_x1_sg U62471 ( .A(n14604), .B(n49529), .X(n14610) );
  nand_x1_sg U62472 ( .A(n15423), .B(n49815), .X(n15429) );
  nand_x1_sg U62473 ( .A(n16242), .B(n50101), .X(n16248) );
  nand_x1_sg U62474 ( .A(n17880), .B(n50675), .X(n17886) );
  nand_x1_sg U62475 ( .A(n18701), .B(n50962), .X(n18707) );
  nand_x1_sg U62476 ( .A(n7233), .B(n46954), .X(n7239) );
  nand_x1_sg U62477 ( .A(n17058), .B(n50386), .X(n17064) );
  nand_x1_sg U62478 ( .A(n7490), .B(n7491), .X(n7489) );
  nor_x1_sg U62479 ( .A(n7491), .B(n7490), .X(n7492) );
  nand_x1_sg U62480 ( .A(n8308), .B(n8309), .X(n8307) );
  nor_x1_sg U62481 ( .A(n8309), .B(n8308), .X(n8310) );
  nand_x1_sg U62482 ( .A(n9126), .B(n9127), .X(n9125) );
  nor_x1_sg U62483 ( .A(n9127), .B(n9126), .X(n9128) );
  nand_x1_sg U62484 ( .A(n9946), .B(n9947), .X(n9945) );
  nor_x1_sg U62485 ( .A(n9947), .B(n9946), .X(n9948) );
  nand_x1_sg U62486 ( .A(n10765), .B(n10766), .X(n10764) );
  nor_x1_sg U62487 ( .A(n10766), .B(n10765), .X(n10767) );
  nand_x1_sg U62488 ( .A(n11584), .B(n11585), .X(n11583) );
  nor_x1_sg U62489 ( .A(n11585), .B(n11584), .X(n11586) );
  nand_x1_sg U62490 ( .A(n12403), .B(n12404), .X(n12402) );
  nor_x1_sg U62491 ( .A(n12404), .B(n12403), .X(n12405) );
  nand_x1_sg U62492 ( .A(n13222), .B(n13223), .X(n13221) );
  nor_x1_sg U62493 ( .A(n13223), .B(n13222), .X(n13224) );
  nand_x1_sg U62494 ( .A(n14041), .B(n14042), .X(n14040) );
  nor_x1_sg U62495 ( .A(n14042), .B(n14041), .X(n14043) );
  nand_x1_sg U62496 ( .A(n14860), .B(n14861), .X(n14859) );
  nor_x1_sg U62497 ( .A(n14861), .B(n14860), .X(n14862) );
  nand_x1_sg U62498 ( .A(n15679), .B(n15680), .X(n15678) );
  nor_x1_sg U62499 ( .A(n15680), .B(n15679), .X(n15681) );
  nand_x1_sg U62500 ( .A(n16498), .B(n16499), .X(n16497) );
  nor_x1_sg U62501 ( .A(n16499), .B(n16498), .X(n16500) );
  nand_x1_sg U62502 ( .A(n18136), .B(n18137), .X(n18135) );
  nor_x1_sg U62503 ( .A(n18137), .B(n18136), .X(n18138) );
  nand_x1_sg U62504 ( .A(n18957), .B(n18958), .X(n18956) );
  nor_x1_sg U62505 ( .A(n18958), .B(n18957), .X(n18959) );
  nand_x1_sg U62506 ( .A(n47285), .B(n8130), .X(n8136) );
  inv_x1_sg U62507 ( .A(n8129), .X(n47285) );
  nand_x1_sg U62508 ( .A(n47570), .B(n8948), .X(n8954) );
  inv_x1_sg U62509 ( .A(n8947), .X(n47570) );
  nand_x1_sg U62510 ( .A(n47855), .B(n9768), .X(n9774) );
  inv_x1_sg U62511 ( .A(n9767), .X(n47855) );
  nand_x1_sg U62512 ( .A(n48140), .B(n10587), .X(n10593) );
  inv_x1_sg U62513 ( .A(n10586), .X(n48140) );
  nand_x1_sg U62514 ( .A(n48425), .B(n11406), .X(n11412) );
  inv_x1_sg U62515 ( .A(n11405), .X(n48425) );
  nand_x1_sg U62516 ( .A(n48710), .B(n12225), .X(n12231) );
  inv_x1_sg U62517 ( .A(n12224), .X(n48710) );
  nand_x1_sg U62518 ( .A(n48996), .B(n13044), .X(n13050) );
  inv_x1_sg U62519 ( .A(n13043), .X(n48996) );
  nand_x1_sg U62520 ( .A(n49283), .B(n13863), .X(n13869) );
  inv_x1_sg U62521 ( .A(n13862), .X(n49283) );
  nand_x1_sg U62522 ( .A(n49569), .B(n14682), .X(n14688) );
  inv_x1_sg U62523 ( .A(n14681), .X(n49569) );
  nand_x1_sg U62524 ( .A(n49855), .B(n15501), .X(n15507) );
  inv_x1_sg U62525 ( .A(n15500), .X(n49855) );
  nand_x1_sg U62526 ( .A(n50141), .B(n16320), .X(n16326) );
  inv_x1_sg U62527 ( .A(n16319), .X(n50141) );
  nand_x1_sg U62528 ( .A(n50715), .B(n17958), .X(n17964) );
  inv_x1_sg U62529 ( .A(n17957), .X(n50715) );
  nand_x1_sg U62530 ( .A(n51002), .B(n18779), .X(n18785) );
  inv_x1_sg U62531 ( .A(n18778), .X(n51002) );
  nand_x1_sg U62532 ( .A(n46898), .B(n7079), .X(n7150) );
  nand_x1_sg U62533 ( .A(n47193), .B(n7897), .X(n7968) );
  nand_x1_sg U62534 ( .A(n47478), .B(n8715), .X(n8786) );
  nand_x1_sg U62535 ( .A(n47763), .B(n9535), .X(n9606) );
  nand_x1_sg U62536 ( .A(n48048), .B(n10354), .X(n10425) );
  nand_x1_sg U62537 ( .A(n48333), .B(n11173), .X(n11244) );
  nand_x1_sg U62538 ( .A(n48618), .B(n11992), .X(n12063) );
  nand_x1_sg U62539 ( .A(n48904), .B(n12811), .X(n12882) );
  nand_x1_sg U62540 ( .A(n49191), .B(n13630), .X(n13701) );
  nand_x1_sg U62541 ( .A(n49477), .B(n14449), .X(n14520) );
  nand_x1_sg U62542 ( .A(n49763), .B(n15268), .X(n15339) );
  nand_x1_sg U62543 ( .A(n50049), .B(n16087), .X(n16158) );
  nand_x1_sg U62544 ( .A(n50331), .B(n16906), .X(n16975) );
  nand_x1_sg U62545 ( .A(n50623), .B(n17725), .X(n17796) );
  nand_x1_sg U62546 ( .A(n50910), .B(n18546), .X(n18617) );
  inv_x1_sg U62547 ( .A(n17101), .X(n50394) );
  inv_x1_sg U62548 ( .A(n25927), .X(n50282) );
  inv_x1_sg U62549 ( .A(n22616), .X(n46866) );
  inv_x1_sg U62550 ( .A(n22622), .X(n46876) );
  inv_x1_sg U62551 ( .A(n22880), .X(n47159) );
  inv_x1_sg U62552 ( .A(n22887), .X(n47169) );
  inv_x1_sg U62553 ( .A(n23157), .X(n47444) );
  inv_x1_sg U62554 ( .A(n23164), .X(n47454) );
  inv_x1_sg U62555 ( .A(n23437), .X(n47729) );
  inv_x1_sg U62556 ( .A(n23444), .X(n47739) );
  inv_x1_sg U62557 ( .A(n23716), .X(n48014) );
  inv_x1_sg U62558 ( .A(n23723), .X(n48024) );
  inv_x1_sg U62559 ( .A(n23995), .X(n48299) );
  inv_x1_sg U62560 ( .A(n24002), .X(n48309) );
  inv_x1_sg U62561 ( .A(n24274), .X(n48584) );
  inv_x1_sg U62562 ( .A(n24281), .X(n48594) );
  inv_x1_sg U62563 ( .A(n24553), .X(n48870) );
  inv_x1_sg U62564 ( .A(n24560), .X(n48880) );
  inv_x1_sg U62565 ( .A(n24831), .X(n49157) );
  inv_x1_sg U62566 ( .A(n24838), .X(n49167) );
  inv_x1_sg U62567 ( .A(n25110), .X(n49443) );
  inv_x1_sg U62568 ( .A(n25117), .X(n49453) );
  inv_x1_sg U62569 ( .A(n25389), .X(n49728) );
  inv_x1_sg U62570 ( .A(n25396), .X(n49738) );
  inv_x1_sg U62571 ( .A(n25668), .X(n50015) );
  inv_x1_sg U62572 ( .A(n25675), .X(n50025) );
  inv_x1_sg U62573 ( .A(n25939), .X(n50299) );
  inv_x1_sg U62574 ( .A(n26212), .X(n50589) );
  inv_x1_sg U62575 ( .A(n26220), .X(n50599) );
  inv_x1_sg U62576 ( .A(n26505), .X(n50876) );
  inv_x1_sg U62577 ( .A(n26512), .X(n50886) );
  nor_x1_sg U62578 ( .A(n6865), .B(n6866), .X(n6864) );
  nor_x1_sg U62579 ( .A(n7682), .B(n7683), .X(n7681) );
  nor_x1_sg U62580 ( .A(n8500), .B(n8501), .X(n8499) );
  nor_x1_sg U62581 ( .A(n9320), .B(n9321), .X(n9319) );
  nor_x1_sg U62582 ( .A(n10139), .B(n10140), .X(n10138) );
  nor_x1_sg U62583 ( .A(n10958), .B(n10959), .X(n10957) );
  nor_x1_sg U62584 ( .A(n11777), .B(n11778), .X(n11776) );
  nor_x1_sg U62585 ( .A(n12596), .B(n12597), .X(n12595) );
  nor_x1_sg U62586 ( .A(n13415), .B(n13416), .X(n13414) );
  nor_x1_sg U62587 ( .A(n14234), .B(n14235), .X(n14233) );
  nor_x1_sg U62588 ( .A(n15053), .B(n15054), .X(n15052) );
  nor_x1_sg U62589 ( .A(n15872), .B(n15873), .X(n15871) );
  nor_x1_sg U62590 ( .A(n16689), .B(n16690), .X(n16688) );
  nor_x1_sg U62591 ( .A(n17510), .B(n17511), .X(n17509) );
  nor_x1_sg U62592 ( .A(n18331), .B(n18332), .X(n18330) );
  nor_x1_sg U62593 ( .A(n6871), .B(n6872), .X(n6870) );
  nor_x1_sg U62594 ( .A(n7688), .B(n7689), .X(n7687) );
  nor_x1_sg U62595 ( .A(n8506), .B(n8507), .X(n8505) );
  nor_x1_sg U62596 ( .A(n9326), .B(n9327), .X(n9325) );
  nor_x1_sg U62597 ( .A(n10145), .B(n10146), .X(n10144) );
  nor_x1_sg U62598 ( .A(n10964), .B(n10965), .X(n10963) );
  nor_x1_sg U62599 ( .A(n11783), .B(n11784), .X(n11782) );
  nor_x1_sg U62600 ( .A(n12602), .B(n12603), .X(n12601) );
  nor_x1_sg U62601 ( .A(n13421), .B(n13422), .X(n13420) );
  nor_x1_sg U62602 ( .A(n14240), .B(n14241), .X(n14239) );
  nor_x1_sg U62603 ( .A(n15059), .B(n15060), .X(n15058) );
  nor_x1_sg U62604 ( .A(n15878), .B(n15879), .X(n15877) );
  nor_x1_sg U62605 ( .A(n16695), .B(n16696), .X(n16694) );
  nor_x1_sg U62606 ( .A(n17516), .B(n17517), .X(n17515) );
  nor_x1_sg U62607 ( .A(n18337), .B(n18338), .X(n18336) );
  nand_x1_sg U62608 ( .A(n7439), .B(n6991), .X(n7435) );
  nand_x1_sg U62609 ( .A(n7437), .B(n41692), .X(n7436) );
  nor_x1_sg U62610 ( .A(n7440), .B(n40367), .X(n7439) );
  nand_x1_sg U62611 ( .A(n8257), .B(n39532), .X(n8253) );
  nand_x1_sg U62612 ( .A(n8255), .B(n41665), .X(n8254) );
  nor_x1_sg U62613 ( .A(n8258), .B(n40307), .X(n8257) );
  nand_x1_sg U62614 ( .A(n9075), .B(n39533), .X(n9071) );
  nand_x1_sg U62615 ( .A(n9073), .B(n41688), .X(n9072) );
  nor_x1_sg U62616 ( .A(n9076), .B(n41843), .X(n9075) );
  nand_x1_sg U62617 ( .A(n9895), .B(n39534), .X(n9891) );
  nand_x1_sg U62618 ( .A(n9893), .B(n41690), .X(n9892) );
  nor_x1_sg U62619 ( .A(n9896), .B(n41756), .X(n9895) );
  nand_x1_sg U62620 ( .A(n10714), .B(n39535), .X(n10710) );
  nand_x1_sg U62621 ( .A(n10712), .B(n41686), .X(n10711) );
  nor_x1_sg U62622 ( .A(n10715), .B(n41757), .X(n10714) );
  nand_x1_sg U62623 ( .A(n11533), .B(n39536), .X(n11529) );
  nand_x1_sg U62624 ( .A(n11531), .B(n41684), .X(n11530) );
  nor_x1_sg U62625 ( .A(n11534), .B(n41758), .X(n11533) );
  nand_x1_sg U62626 ( .A(n12352), .B(n39537), .X(n12348) );
  nand_x1_sg U62627 ( .A(n12350), .B(n41682), .X(n12349) );
  nor_x1_sg U62628 ( .A(n12353), .B(n41763), .X(n12352) );
  nand_x1_sg U62629 ( .A(n13171), .B(n39538), .X(n13167) );
  nand_x1_sg U62630 ( .A(n13169), .B(n41680), .X(n13168) );
  nor_x1_sg U62631 ( .A(n13172), .B(n41760), .X(n13171) );
  nand_x1_sg U62632 ( .A(n13990), .B(n39539), .X(n13986) );
  nand_x1_sg U62633 ( .A(n13988), .B(n41678), .X(n13987) );
  nor_x1_sg U62634 ( .A(n13991), .B(n41761), .X(n13990) );
  nand_x1_sg U62635 ( .A(n14809), .B(n39540), .X(n14805) );
  nand_x1_sg U62636 ( .A(n14807), .B(n41676), .X(n14806) );
  nor_x1_sg U62637 ( .A(n14810), .B(n39066), .X(n14809) );
  nand_x1_sg U62638 ( .A(n15628), .B(n39541), .X(n15624) );
  nand_x1_sg U62639 ( .A(n15626), .B(n41663), .X(n15625) );
  nor_x1_sg U62640 ( .A(n15629), .B(n41765), .X(n15628) );
  nand_x1_sg U62641 ( .A(n16447), .B(n39542), .X(n16443) );
  nand_x1_sg U62642 ( .A(n16445), .B(n41674), .X(n16444) );
  nor_x1_sg U62643 ( .A(n16448), .B(n39067), .X(n16447) );
  nand_x1_sg U62644 ( .A(n18085), .B(n17636), .X(n18081) );
  nand_x1_sg U62645 ( .A(n18083), .B(n41670), .X(n18082) );
  nor_x1_sg U62646 ( .A(n18086), .B(n40363), .X(n18085) );
  nand_x1_sg U62647 ( .A(n18906), .B(n39544), .X(n18902) );
  nand_x1_sg U62648 ( .A(n18904), .B(n41668), .X(n18903) );
  nor_x1_sg U62649 ( .A(n18907), .B(n39068), .X(n18906) );
  nand_x1_sg U62650 ( .A(n17264), .B(n39661), .X(n17260) );
  nand_x1_sg U62651 ( .A(n17262), .B(n41672), .X(n17261) );
  nor_x1_sg U62652 ( .A(n17265), .B(n41842), .X(n17264) );
  nor_x1_sg U62653 ( .A(n38905), .B(n7659), .X(\L2_0/n3432 ) );
  nor_x1_sg U62654 ( .A(n40975), .B(n7678), .X(\L2_0/n3420 ) );
  nor_x1_sg U62655 ( .A(n7638), .B(n7684), .X(\L2_0/n3416 ) );
  nor_x1_sg U62656 ( .A(n40974), .B(n7696), .X(\L2_0/n3408 ) );
  nand_x1_sg U62657 ( .A(n8295), .B(n39563), .X(n8293) );
  nand_x1_sg U62658 ( .A(n40105), .B(n47351), .X(n8294) );
  nand_x1_sg U62659 ( .A(n9113), .B(n39566), .X(n9111) );
  nand_x1_sg U62660 ( .A(n8853), .B(n47636), .X(n9112) );
  nand_x1_sg U62661 ( .A(n9933), .B(n39569), .X(n9931) );
  nand_x1_sg U62662 ( .A(n40110), .B(n47921), .X(n9932) );
  nand_x1_sg U62663 ( .A(n10752), .B(n39572), .X(n10750) );
  nand_x1_sg U62664 ( .A(n10492), .B(n48206), .X(n10751) );
  nand_x1_sg U62665 ( .A(n11571), .B(n39575), .X(n11569) );
  nand_x1_sg U62666 ( .A(n11311), .B(n48491), .X(n11570) );
  nand_x1_sg U62667 ( .A(n12390), .B(n39578), .X(n12388) );
  nand_x1_sg U62668 ( .A(n40116), .B(n48776), .X(n12389) );
  nand_x1_sg U62669 ( .A(n13209), .B(n39581), .X(n13207) );
  nand_x1_sg U62670 ( .A(n12949), .B(n49063), .X(n13208) );
  nand_x1_sg U62671 ( .A(n14028), .B(n39584), .X(n14026) );
  nand_x1_sg U62672 ( .A(n13768), .B(n49349), .X(n14027) );
  nand_x1_sg U62673 ( .A(n14847), .B(n39587), .X(n14845) );
  nand_x1_sg U62674 ( .A(n40122), .B(n49635), .X(n14846) );
  nand_x1_sg U62675 ( .A(n15666), .B(n39590), .X(n15664) );
  nand_x1_sg U62676 ( .A(n40123), .B(n49921), .X(n15665) );
  nand_x1_sg U62677 ( .A(n16485), .B(n39593), .X(n16483) );
  nand_x1_sg U62678 ( .A(n16225), .B(n50207), .X(n16484) );
  nand_x1_sg U62679 ( .A(n17302), .B(n39561), .X(n17300) );
  nand_x1_sg U62680 ( .A(n17041), .B(n50492), .X(n17301) );
  nand_x1_sg U62681 ( .A(n18123), .B(n39600), .X(n18121) );
  nand_x1_sg U62682 ( .A(n40132), .B(n50781), .X(n18122) );
  nand_x1_sg U62683 ( .A(n18944), .B(n39596), .X(n18942) );
  nand_x1_sg U62684 ( .A(n40128), .B(n51068), .X(n18943) );
  nand_x1_sg U62685 ( .A(n46977), .B(n46954), .X(n7232) );
  nand_x1_sg U62686 ( .A(n7234), .B(n7233), .X(n7231) );
  inv_x1_sg U62687 ( .A(n7233), .X(n46977) );
  nand_x1_sg U62688 ( .A(n47267), .B(n47245), .X(n8051) );
  nand_x1_sg U62689 ( .A(n8053), .B(n8052), .X(n8050) );
  inv_x1_sg U62690 ( .A(n8052), .X(n47267) );
  nand_x1_sg U62691 ( .A(n47552), .B(n47530), .X(n8869) );
  nand_x1_sg U62692 ( .A(n8871), .B(n8870), .X(n8868) );
  inv_x1_sg U62693 ( .A(n8870), .X(n47552) );
  nand_x1_sg U62694 ( .A(n47837), .B(n47815), .X(n9689) );
  nand_x1_sg U62695 ( .A(n9691), .B(n9690), .X(n9688) );
  inv_x1_sg U62696 ( .A(n9690), .X(n47837) );
  nand_x1_sg U62697 ( .A(n48122), .B(n48100), .X(n10508) );
  nand_x1_sg U62698 ( .A(n10510), .B(n10509), .X(n10507) );
  inv_x1_sg U62699 ( .A(n10509), .X(n48122) );
  nand_x1_sg U62700 ( .A(n48407), .B(n48385), .X(n11327) );
  nand_x1_sg U62701 ( .A(n11329), .B(n11328), .X(n11326) );
  inv_x1_sg U62702 ( .A(n11328), .X(n48407) );
  nand_x1_sg U62703 ( .A(n48692), .B(n48670), .X(n12146) );
  nand_x1_sg U62704 ( .A(n12148), .B(n12147), .X(n12145) );
  inv_x1_sg U62705 ( .A(n12147), .X(n48692) );
  nand_x1_sg U62706 ( .A(n48978), .B(n48956), .X(n12965) );
  nand_x1_sg U62707 ( .A(n12967), .B(n12966), .X(n12964) );
  inv_x1_sg U62708 ( .A(n12966), .X(n48978) );
  nand_x1_sg U62709 ( .A(n49265), .B(n49243), .X(n13784) );
  nand_x1_sg U62710 ( .A(n13786), .B(n13785), .X(n13783) );
  inv_x1_sg U62711 ( .A(n13785), .X(n49265) );
  nand_x1_sg U62712 ( .A(n49551), .B(n49529), .X(n14603) );
  nand_x1_sg U62713 ( .A(n14605), .B(n14604), .X(n14602) );
  inv_x1_sg U62714 ( .A(n14604), .X(n49551) );
  nand_x1_sg U62715 ( .A(n49837), .B(n49815), .X(n15422) );
  nand_x1_sg U62716 ( .A(n15424), .B(n15423), .X(n15421) );
  inv_x1_sg U62717 ( .A(n15423), .X(n49837) );
  nand_x1_sg U62718 ( .A(n50123), .B(n50101), .X(n16241) );
  nand_x1_sg U62719 ( .A(n16243), .B(n16242), .X(n16240) );
  inv_x1_sg U62720 ( .A(n16242), .X(n50123) );
  nand_x1_sg U62721 ( .A(n50408), .B(n50386), .X(n17057) );
  nand_x1_sg U62722 ( .A(n17059), .B(n17058), .X(n17056) );
  inv_x1_sg U62723 ( .A(n17058), .X(n50408) );
  nand_x1_sg U62724 ( .A(n50697), .B(n50675), .X(n17879) );
  nand_x1_sg U62725 ( .A(n17881), .B(n17880), .X(n17878) );
  inv_x1_sg U62726 ( .A(n17880), .X(n50697) );
  nand_x1_sg U62727 ( .A(n50984), .B(n50962), .X(n18700) );
  nand_x1_sg U62728 ( .A(n18702), .B(n18701), .X(n18699) );
  inv_x1_sg U62729 ( .A(n18701), .X(n50984) );
  nand_x1_sg U62730 ( .A(n8353), .B(n39799), .X(n8352) );
  nand_x1_sg U62731 ( .A(n8354), .B(n8355), .X(n8351) );
  nor_x1_sg U62732 ( .A(n8354), .B(n40560), .X(n8353) );
  nand_x1_sg U62733 ( .A(n9171), .B(n39801), .X(n9170) );
  nand_x1_sg U62734 ( .A(n9172), .B(n9173), .X(n9169) );
  nor_x1_sg U62735 ( .A(n9172), .B(n8469), .X(n9171) );
  nand_x1_sg U62736 ( .A(n9991), .B(n39795), .X(n9990) );
  nand_x1_sg U62737 ( .A(n9992), .B(n9993), .X(n9989) );
  nor_x1_sg U62738 ( .A(n9992), .B(n40551), .X(n9991) );
  nand_x1_sg U62739 ( .A(n10810), .B(n39797), .X(n10809) );
  nand_x1_sg U62740 ( .A(n10811), .B(n10812), .X(n10808) );
  nor_x1_sg U62741 ( .A(n10811), .B(n40549), .X(n10810) );
  nand_x1_sg U62742 ( .A(n11629), .B(n39791), .X(n11628) );
  nand_x1_sg U62743 ( .A(n11630), .B(n11631), .X(n11627) );
  nor_x1_sg U62744 ( .A(n11630), .B(n40543), .X(n11629) );
  nand_x1_sg U62745 ( .A(n12448), .B(n39793), .X(n12447) );
  nand_x1_sg U62746 ( .A(n12449), .B(n12450), .X(n12446) );
  nor_x1_sg U62747 ( .A(n12449), .B(n40540), .X(n12448) );
  nand_x1_sg U62748 ( .A(n13267), .B(n39787), .X(n13266) );
  nand_x1_sg U62749 ( .A(n13268), .B(n13269), .X(n13265) );
  nor_x1_sg U62750 ( .A(n13268), .B(n40536), .X(n13267) );
  nand_x1_sg U62751 ( .A(n14086), .B(n39789), .X(n14085) );
  nand_x1_sg U62752 ( .A(n14087), .B(n14088), .X(n14084) );
  nor_x1_sg U62753 ( .A(n14087), .B(n40533), .X(n14086) );
  nand_x1_sg U62754 ( .A(n14905), .B(n39783), .X(n14904) );
  nand_x1_sg U62755 ( .A(n14906), .B(n14907), .X(n14903) );
  nor_x1_sg U62756 ( .A(n14906), .B(n14203), .X(n14905) );
  nand_x1_sg U62757 ( .A(n15724), .B(n39785), .X(n15723) );
  nand_x1_sg U62758 ( .A(n15725), .B(n15726), .X(n15722) );
  nor_x1_sg U62759 ( .A(n15725), .B(n40525), .X(n15724) );
  nand_x1_sg U62760 ( .A(n16543), .B(n39779), .X(n16542) );
  nand_x1_sg U62761 ( .A(n16544), .B(n16545), .X(n16541) );
  nor_x1_sg U62762 ( .A(n16544), .B(n40519), .X(n16543) );
  nand_x1_sg U62763 ( .A(n18181), .B(n39781), .X(n18180) );
  nand_x1_sg U62764 ( .A(n18182), .B(n18183), .X(n18179) );
  nor_x1_sg U62765 ( .A(n18182), .B(n40516), .X(n18181) );
  nand_x1_sg U62766 ( .A(n19002), .B(n39776), .X(n19001) );
  nand_x1_sg U62767 ( .A(n19003), .B(n19004), .X(n19000) );
  nor_x1_sg U62768 ( .A(n19003), .B(n40512), .X(n19002) );
  nand_x1_sg U62769 ( .A(n7535), .B(n39803), .X(n7534) );
  nand_x1_sg U62770 ( .A(n7536), .B(n7537), .X(n7533) );
  nor_x1_sg U62771 ( .A(n7536), .B(n40613), .X(n7535) );
  nand_x1_sg U62772 ( .A(n17360), .B(n39775), .X(n17359) );
  nand_x1_sg U62773 ( .A(n17361), .B(n17362), .X(n17358) );
  nor_x1_sg U62774 ( .A(n17361), .B(n40301), .X(n17360) );
  nand_x1_sg U62775 ( .A(n7778), .B(n7779), .X(n8406) );
  nor_x1_sg U62776 ( .A(n7778), .B(n7779), .X(n8407) );
  nand_x1_sg U62777 ( .A(n8596), .B(n8597), .X(n9224) );
  nor_x1_sg U62778 ( .A(n8596), .B(n8597), .X(n9225) );
  nand_x1_sg U62779 ( .A(n9416), .B(n9417), .X(n10044) );
  nor_x1_sg U62780 ( .A(n9416), .B(n9417), .X(n10045) );
  nand_x1_sg U62781 ( .A(n10235), .B(n10236), .X(n10863) );
  nor_x1_sg U62782 ( .A(n10235), .B(n10236), .X(n10864) );
  nand_x1_sg U62783 ( .A(n11054), .B(n11055), .X(n11682) );
  nor_x1_sg U62784 ( .A(n11054), .B(n11055), .X(n11683) );
  nand_x1_sg U62785 ( .A(n11873), .B(n11874), .X(n12501) );
  nor_x1_sg U62786 ( .A(n11873), .B(n11874), .X(n12502) );
  nand_x1_sg U62787 ( .A(n12692), .B(n12693), .X(n13320) );
  nor_x1_sg U62788 ( .A(n12692), .B(n12693), .X(n13321) );
  nand_x1_sg U62789 ( .A(n13511), .B(n13512), .X(n14139) );
  nor_x1_sg U62790 ( .A(n13511), .B(n13512), .X(n14140) );
  nand_x1_sg U62791 ( .A(n14330), .B(n14331), .X(n14958) );
  nor_x1_sg U62792 ( .A(n14330), .B(n14331), .X(n14959) );
  nand_x1_sg U62793 ( .A(n15149), .B(n15150), .X(n15777) );
  nor_x1_sg U62794 ( .A(n15149), .B(n15150), .X(n15778) );
  nand_x1_sg U62795 ( .A(n15968), .B(n15969), .X(n16596) );
  nor_x1_sg U62796 ( .A(n15968), .B(n15969), .X(n16597) );
  nand_x1_sg U62797 ( .A(n17606), .B(n17607), .X(n18234) );
  nor_x1_sg U62798 ( .A(n17606), .B(n17607), .X(n18235) );
  nand_x1_sg U62799 ( .A(n18427), .B(n18428), .X(n19055) );
  nor_x1_sg U62800 ( .A(n18427), .B(n18428), .X(n19056) );
  nand_x1_sg U62801 ( .A(n7107), .B(n7108), .X(n7105) );
  nor_x1_sg U62802 ( .A(n7107), .B(n7108), .X(n7106) );
  nand_x1_sg U62803 ( .A(n7925), .B(n7926), .X(n7923) );
  nor_x1_sg U62804 ( .A(n7925), .B(n7926), .X(n7924) );
  nand_x1_sg U62805 ( .A(n8743), .B(n8744), .X(n8741) );
  nor_x1_sg U62806 ( .A(n8743), .B(n8744), .X(n8742) );
  nand_x1_sg U62807 ( .A(n9563), .B(n9564), .X(n9561) );
  nor_x1_sg U62808 ( .A(n9563), .B(n9564), .X(n9562) );
  nand_x1_sg U62809 ( .A(n10382), .B(n10383), .X(n10380) );
  nor_x1_sg U62810 ( .A(n10382), .B(n10383), .X(n10381) );
  nand_x1_sg U62811 ( .A(n11201), .B(n11202), .X(n11199) );
  nor_x1_sg U62812 ( .A(n11201), .B(n11202), .X(n11200) );
  nand_x1_sg U62813 ( .A(n12020), .B(n12021), .X(n12018) );
  nor_x1_sg U62814 ( .A(n12020), .B(n12021), .X(n12019) );
  nand_x1_sg U62815 ( .A(n12839), .B(n12840), .X(n12837) );
  nor_x1_sg U62816 ( .A(n12839), .B(n12840), .X(n12838) );
  nand_x1_sg U62817 ( .A(n13658), .B(n13659), .X(n13656) );
  nor_x1_sg U62818 ( .A(n13658), .B(n13659), .X(n13657) );
  nand_x1_sg U62819 ( .A(n14477), .B(n14478), .X(n14475) );
  nor_x1_sg U62820 ( .A(n14477), .B(n14478), .X(n14476) );
  nand_x1_sg U62821 ( .A(n15296), .B(n15297), .X(n15294) );
  nor_x1_sg U62822 ( .A(n15296), .B(n15297), .X(n15295) );
  nand_x1_sg U62823 ( .A(n16115), .B(n16116), .X(n16113) );
  nor_x1_sg U62824 ( .A(n16115), .B(n16116), .X(n16114) );
  nand_x1_sg U62825 ( .A(n17753), .B(n17754), .X(n17751) );
  nor_x1_sg U62826 ( .A(n17753), .B(n17754), .X(n17752) );
  nand_x1_sg U62827 ( .A(n18574), .B(n18575), .X(n18572) );
  nor_x1_sg U62828 ( .A(n18574), .B(n18575), .X(n18573) );
  nand_x1_sg U62829 ( .A(n16932), .B(n16933), .X(n16930) );
  nor_x1_sg U62830 ( .A(n16932), .B(n16933), .X(n16931) );
  nand_x1_sg U62831 ( .A(n7477), .B(n39850), .X(n7475) );
  nand_x1_sg U62832 ( .A(n39930), .B(n47065), .X(n7476) );
  inv_x1_sg U62833 ( .A(n6854), .X(n46872) );
  inv_x1_sg U62834 ( .A(n7671), .X(n47165) );
  inv_x1_sg U62835 ( .A(n8489), .X(n47450) );
  inv_x1_sg U62836 ( .A(n9309), .X(n47735) );
  inv_x1_sg U62837 ( .A(n10128), .X(n48020) );
  inv_x1_sg U62838 ( .A(n10947), .X(n48305) );
  inv_x1_sg U62839 ( .A(n11766), .X(n48590) );
  inv_x1_sg U62840 ( .A(n12585), .X(n48876) );
  inv_x1_sg U62841 ( .A(n13404), .X(n49163) );
  inv_x1_sg U62842 ( .A(n14223), .X(n49449) );
  inv_x1_sg U62843 ( .A(n15042), .X(n49734) );
  inv_x1_sg U62844 ( .A(n15861), .X(n50021) );
  inv_x1_sg U62845 ( .A(n17499), .X(n50595) );
  inv_x1_sg U62846 ( .A(n18320), .X(n50882) );
  nand_x1_sg U62847 ( .A(n8090), .B(n8091), .X(n8088) );
  nor_x1_sg U62848 ( .A(n8090), .B(n8091), .X(n8089) );
  nand_x1_sg U62849 ( .A(n8908), .B(n8909), .X(n8906) );
  nor_x1_sg U62850 ( .A(n8908), .B(n8909), .X(n8907) );
  nand_x1_sg U62851 ( .A(n9728), .B(n9729), .X(n9726) );
  nor_x1_sg U62852 ( .A(n9728), .B(n9729), .X(n9727) );
  nand_x1_sg U62853 ( .A(n10547), .B(n10548), .X(n10545) );
  nor_x1_sg U62854 ( .A(n10547), .B(n10548), .X(n10546) );
  nand_x1_sg U62855 ( .A(n11366), .B(n11367), .X(n11364) );
  nor_x1_sg U62856 ( .A(n11366), .B(n11367), .X(n11365) );
  nand_x1_sg U62857 ( .A(n12185), .B(n12186), .X(n12183) );
  nor_x1_sg U62858 ( .A(n12185), .B(n12186), .X(n12184) );
  nand_x1_sg U62859 ( .A(n13004), .B(n13005), .X(n13002) );
  nor_x1_sg U62860 ( .A(n13004), .B(n13005), .X(n13003) );
  nand_x1_sg U62861 ( .A(n13823), .B(n13824), .X(n13821) );
  nor_x1_sg U62862 ( .A(n13823), .B(n13824), .X(n13822) );
  nand_x1_sg U62863 ( .A(n14642), .B(n14643), .X(n14640) );
  nor_x1_sg U62864 ( .A(n14642), .B(n14643), .X(n14641) );
  nand_x1_sg U62865 ( .A(n15461), .B(n15462), .X(n15459) );
  nor_x1_sg U62866 ( .A(n15461), .B(n15462), .X(n15460) );
  nand_x1_sg U62867 ( .A(n16280), .B(n16281), .X(n16278) );
  nor_x1_sg U62868 ( .A(n16280), .B(n16281), .X(n16279) );
  nand_x1_sg U62869 ( .A(n17096), .B(n17097), .X(n17094) );
  nor_x1_sg U62870 ( .A(n17096), .B(n17097), .X(n17095) );
  nand_x1_sg U62871 ( .A(n17918), .B(n17919), .X(n17916) );
  nor_x1_sg U62872 ( .A(n17918), .B(n17919), .X(n17917) );
  nand_x1_sg U62873 ( .A(n18739), .B(n18740), .X(n18737) );
  nor_x1_sg U62874 ( .A(n18739), .B(n18740), .X(n18738) );
  nand_x1_sg U62875 ( .A(n7271), .B(n7272), .X(n7269) );
  nor_x1_sg U62876 ( .A(n7271), .B(n7272), .X(n7270) );
  nand_x1_sg U62877 ( .A(n7818), .B(n42311), .X(n7817) );
  nand_x1_sg U62878 ( .A(n7819), .B(n7820), .X(n7816) );
  nor_x1_sg U62879 ( .A(n7819), .B(n40559), .X(n7818) );
  nand_x1_sg U62880 ( .A(n8636), .B(n42310), .X(n8635) );
  nand_x1_sg U62881 ( .A(n8637), .B(n8638), .X(n8634) );
  nor_x1_sg U62882 ( .A(n8637), .B(n40555), .X(n8636) );
  nand_x1_sg U62883 ( .A(n9456), .B(n42309), .X(n9455) );
  nand_x1_sg U62884 ( .A(n9457), .B(n9458), .X(n9454) );
  nor_x1_sg U62885 ( .A(n9457), .B(n40553), .X(n9456) );
  nand_x1_sg U62886 ( .A(n10275), .B(n10272), .X(n10274) );
  nand_x1_sg U62887 ( .A(n10276), .B(n10277), .X(n10273) );
  nor_x1_sg U62888 ( .A(n10276), .B(n40547), .X(n10275) );
  nand_x1_sg U62889 ( .A(n11094), .B(n42308), .X(n11093) );
  nand_x1_sg U62890 ( .A(n11095), .B(n11096), .X(n11092) );
  nor_x1_sg U62891 ( .A(n11095), .B(n40545), .X(n11094) );
  nand_x1_sg U62892 ( .A(n11913), .B(n42307), .X(n11912) );
  nand_x1_sg U62893 ( .A(n11914), .B(n11915), .X(n11911) );
  nor_x1_sg U62894 ( .A(n11914), .B(n40539), .X(n11913) );
  nand_x1_sg U62895 ( .A(n12732), .B(n42306), .X(n12731) );
  nand_x1_sg U62896 ( .A(n12733), .B(n12734), .X(n12730) );
  nor_x1_sg U62897 ( .A(n12733), .B(n40535), .X(n12732) );
  nand_x1_sg U62898 ( .A(n13551), .B(n13548), .X(n13550) );
  nand_x1_sg U62899 ( .A(n13552), .B(n13553), .X(n13549) );
  nor_x1_sg U62900 ( .A(n13552), .B(n40531), .X(n13551) );
  nand_x1_sg U62901 ( .A(n14370), .B(n42305), .X(n14369) );
  nand_x1_sg U62902 ( .A(n14371), .B(n14372), .X(n14368) );
  nor_x1_sg U62903 ( .A(n14371), .B(n40527), .X(n14370) );
  nand_x1_sg U62904 ( .A(n15189), .B(n42304), .X(n15188) );
  nand_x1_sg U62905 ( .A(n15190), .B(n15191), .X(n15187) );
  nor_x1_sg U62906 ( .A(n15190), .B(n40523), .X(n15189) );
  nand_x1_sg U62907 ( .A(n16008), .B(n42303), .X(n16007) );
  nand_x1_sg U62908 ( .A(n16009), .B(n16010), .X(n16006) );
  nor_x1_sg U62909 ( .A(n16009), .B(n40521), .X(n16008) );
  nand_x1_sg U62910 ( .A(n17646), .B(n17643), .X(n17645) );
  nand_x1_sg U62911 ( .A(n17647), .B(n17648), .X(n17644) );
  nor_x1_sg U62912 ( .A(n17647), .B(n17479), .X(n17646) );
  nand_x1_sg U62913 ( .A(n18467), .B(n18464), .X(n18466) );
  nand_x1_sg U62914 ( .A(n18468), .B(n18469), .X(n18465) );
  nor_x1_sg U62915 ( .A(n18468), .B(n40511), .X(n18467) );
  nand_x1_sg U62916 ( .A(n7001), .B(n39678), .X(n7000) );
  nand_x1_sg U62917 ( .A(n7002), .B(n7003), .X(n6999) );
  nor_x1_sg U62918 ( .A(n7002), .B(n40613), .X(n7001) );
  nand_x1_sg U62919 ( .A(n16825), .B(n39807), .X(n16824) );
  nand_x1_sg U62920 ( .A(n16826), .B(n16827), .X(n16823) );
  nor_x1_sg U62921 ( .A(n16826), .B(n40302), .X(n16825) );
  nand_x1_sg U62922 ( .A(n6945), .B(n42074), .X(n7627) );
  nor_x1_sg U62923 ( .A(n6945), .B(n42074), .X(n7628) );
  nand_x1_sg U62924 ( .A(n16769), .B(n42088), .X(n17452) );
  nor_x1_sg U62925 ( .A(n16769), .B(n42088), .X(n17453) );
  nand_x1_sg U62926 ( .A(n7762), .B(n42073), .X(n8445) );
  nor_x1_sg U62927 ( .A(n7762), .B(n42073), .X(n8446) );
  nand_x1_sg U62928 ( .A(n8580), .B(n42071), .X(n9263) );
  nor_x1_sg U62929 ( .A(n8580), .B(n42071), .X(n9264) );
  nand_x1_sg U62930 ( .A(n9400), .B(n42070), .X(n10083) );
  nor_x1_sg U62931 ( .A(n9400), .B(n42070), .X(n10084) );
  nand_x1_sg U62932 ( .A(n10219), .B(n42069), .X(n10902) );
  nor_x1_sg U62933 ( .A(n10219), .B(n42069), .X(n10903) );
  nand_x1_sg U62934 ( .A(n11038), .B(n42068), .X(n11721) );
  nor_x1_sg U62935 ( .A(n11038), .B(n42068), .X(n11722) );
  nand_x1_sg U62936 ( .A(n11857), .B(n42067), .X(n12540) );
  nor_x1_sg U62937 ( .A(n11857), .B(n42067), .X(n12541) );
  nand_x1_sg U62938 ( .A(n12676), .B(n42066), .X(n13359) );
  nor_x1_sg U62939 ( .A(n12676), .B(n42066), .X(n13360) );
  nand_x1_sg U62940 ( .A(n13495), .B(n42065), .X(n14178) );
  nor_x1_sg U62941 ( .A(n13495), .B(n42065), .X(n14179) );
  nand_x1_sg U62942 ( .A(n14314), .B(n42064), .X(n14997) );
  nor_x1_sg U62943 ( .A(n14314), .B(n42064), .X(n14998) );
  nand_x1_sg U62944 ( .A(n15133), .B(n42072), .X(n15816) );
  nor_x1_sg U62945 ( .A(n15133), .B(n42072), .X(n15817) );
  nand_x1_sg U62946 ( .A(n15952), .B(n42063), .X(n16635) );
  nor_x1_sg U62947 ( .A(n15952), .B(n42063), .X(n16636) );
  nand_x1_sg U62948 ( .A(n17590), .B(n42062), .X(n18273) );
  nor_x1_sg U62949 ( .A(n17590), .B(n42062), .X(n18274) );
  nand_x1_sg U62950 ( .A(n18411), .B(n42061), .X(n19094) );
  nor_x1_sg U62951 ( .A(n18411), .B(n42061), .X(n19095) );
  nand_x1_sg U62952 ( .A(n46993), .B(n7329), .X(n7325) );
  inv_x1_sg U62953 ( .A(n7308), .X(n46994) );
  nand_x1_sg U62954 ( .A(n47282), .B(n8147), .X(n8143) );
  inv_x1_sg U62955 ( .A(n8126), .X(n47283) );
  nand_x1_sg U62956 ( .A(n47567), .B(n8965), .X(n8961) );
  inv_x1_sg U62957 ( .A(n8944), .X(n47568) );
  nand_x1_sg U62958 ( .A(n47852), .B(n9785), .X(n9781) );
  inv_x1_sg U62959 ( .A(n9764), .X(n47853) );
  nand_x1_sg U62960 ( .A(n48137), .B(n10604), .X(n10600) );
  inv_x1_sg U62961 ( .A(n10583), .X(n48138) );
  nand_x1_sg U62962 ( .A(n48422), .B(n11423), .X(n11419) );
  inv_x1_sg U62963 ( .A(n11402), .X(n48423) );
  nand_x1_sg U62964 ( .A(n48707), .B(n12242), .X(n12238) );
  inv_x1_sg U62965 ( .A(n12221), .X(n48708) );
  nand_x1_sg U62966 ( .A(n48993), .B(n13061), .X(n13057) );
  inv_x1_sg U62967 ( .A(n13040), .X(n48994) );
  nand_x1_sg U62968 ( .A(n49280), .B(n13880), .X(n13876) );
  inv_x1_sg U62969 ( .A(n13859), .X(n49281) );
  nand_x1_sg U62970 ( .A(n49566), .B(n14699), .X(n14695) );
  inv_x1_sg U62971 ( .A(n14678), .X(n49567) );
  nand_x1_sg U62972 ( .A(n49852), .B(n15518), .X(n15514) );
  inv_x1_sg U62973 ( .A(n15497), .X(n49853) );
  nand_x1_sg U62974 ( .A(n50138), .B(n16337), .X(n16333) );
  inv_x1_sg U62975 ( .A(n16316), .X(n50139) );
  nand_x1_sg U62976 ( .A(n50712), .B(n17975), .X(n17971) );
  inv_x1_sg U62977 ( .A(n17954), .X(n50713) );
  nand_x1_sg U62978 ( .A(n50999), .B(n18796), .X(n18792) );
  inv_x1_sg U62979 ( .A(n18775), .X(n51000) );
  nand_x1_sg U62980 ( .A(n46887), .B(n46905), .X(n7181) );
  nand_x1_sg U62981 ( .A(n46901), .B(n7165), .X(n7180) );
  nand_x1_sg U62982 ( .A(n47180), .B(n47198), .X(n8000) );
  nand_x1_sg U62983 ( .A(n47186), .B(n7984), .X(n7999) );
  nand_x1_sg U62984 ( .A(n47465), .B(n47483), .X(n8818) );
  nand_x1_sg U62985 ( .A(n47471), .B(n8802), .X(n8817) );
  nand_x1_sg U62986 ( .A(n47750), .B(n47768), .X(n9638) );
  nand_x1_sg U62987 ( .A(n47756), .B(n9622), .X(n9637) );
  nand_x1_sg U62988 ( .A(n48035), .B(n48053), .X(n10457) );
  nand_x1_sg U62989 ( .A(n48041), .B(n10441), .X(n10456) );
  nand_x1_sg U62990 ( .A(n48320), .B(n48338), .X(n11276) );
  nand_x1_sg U62991 ( .A(n48326), .B(n11260), .X(n11275) );
  nand_x1_sg U62992 ( .A(n48605), .B(n48623), .X(n12095) );
  nand_x1_sg U62993 ( .A(n48611), .B(n12079), .X(n12094) );
  nand_x1_sg U62994 ( .A(n48891), .B(n48909), .X(n12914) );
  nand_x1_sg U62995 ( .A(n48897), .B(n12898), .X(n12913) );
  nand_x1_sg U62996 ( .A(n49178), .B(n49196), .X(n13733) );
  nand_x1_sg U62997 ( .A(n49184), .B(n13717), .X(n13732) );
  nand_x1_sg U62998 ( .A(n49464), .B(n49482), .X(n14552) );
  nand_x1_sg U62999 ( .A(n49470), .B(n14536), .X(n14551) );
  nand_x1_sg U63000 ( .A(n49749), .B(n49768), .X(n15371) );
  nand_x1_sg U63001 ( .A(n49756), .B(n15355), .X(n15370) );
  nand_x1_sg U63002 ( .A(n50036), .B(n50054), .X(n16190) );
  nand_x1_sg U63003 ( .A(n50042), .B(n16174), .X(n16189) );
  nand_x1_sg U63004 ( .A(n50321), .B(n50339), .X(n17006) );
  nand_x1_sg U63005 ( .A(n50334), .B(n16990), .X(n17005) );
  nand_x1_sg U63006 ( .A(n50610), .B(n50628), .X(n17828) );
  nand_x1_sg U63007 ( .A(n50616), .B(n17812), .X(n17827) );
  nand_x1_sg U63008 ( .A(n50897), .B(n50915), .X(n18649) );
  nand_x1_sg U63009 ( .A(n50903), .B(n18633), .X(n18648) );
  nand_x1_sg U63010 ( .A(n7509), .B(n7508), .X(n7506) );
  nor_x1_sg U63011 ( .A(n7508), .B(n7509), .X(n7507) );
  nand_x1_sg U63012 ( .A(n8327), .B(n8326), .X(n8324) );
  nor_x1_sg U63013 ( .A(n8326), .B(n8327), .X(n8325) );
  nand_x1_sg U63014 ( .A(n9145), .B(n9144), .X(n9142) );
  nor_x1_sg U63015 ( .A(n9144), .B(n9145), .X(n9143) );
  nand_x1_sg U63016 ( .A(n9965), .B(n9964), .X(n9962) );
  nor_x1_sg U63017 ( .A(n9964), .B(n9965), .X(n9963) );
  nand_x1_sg U63018 ( .A(n10784), .B(n10783), .X(n10781) );
  nor_x1_sg U63019 ( .A(n10783), .B(n10784), .X(n10782) );
  nand_x1_sg U63020 ( .A(n11603), .B(n11602), .X(n11600) );
  nor_x1_sg U63021 ( .A(n11602), .B(n11603), .X(n11601) );
  nand_x1_sg U63022 ( .A(n12422), .B(n12421), .X(n12419) );
  nor_x1_sg U63023 ( .A(n12421), .B(n12422), .X(n12420) );
  nand_x1_sg U63024 ( .A(n13241), .B(n13240), .X(n13238) );
  nor_x1_sg U63025 ( .A(n13240), .B(n13241), .X(n13239) );
  nand_x1_sg U63026 ( .A(n14060), .B(n14059), .X(n14057) );
  nor_x1_sg U63027 ( .A(n14059), .B(n14060), .X(n14058) );
  nand_x1_sg U63028 ( .A(n14879), .B(n14878), .X(n14876) );
  nor_x1_sg U63029 ( .A(n14878), .B(n14879), .X(n14877) );
  nand_x1_sg U63030 ( .A(n15698), .B(n15697), .X(n15695) );
  nor_x1_sg U63031 ( .A(n15697), .B(n15698), .X(n15696) );
  nand_x1_sg U63032 ( .A(n16517), .B(n16516), .X(n16514) );
  nor_x1_sg U63033 ( .A(n16516), .B(n16517), .X(n16515) );
  nand_x1_sg U63034 ( .A(n17334), .B(n17333), .X(n17331) );
  nor_x1_sg U63035 ( .A(n17333), .B(n17334), .X(n17332) );
  nand_x1_sg U63036 ( .A(n18155), .B(n18154), .X(n18152) );
  nor_x1_sg U63037 ( .A(n18154), .B(n18155), .X(n18153) );
  nand_x1_sg U63038 ( .A(n18976), .B(n18975), .X(n18973) );
  nor_x1_sg U63039 ( .A(n18975), .B(n18976), .X(n18974) );
  nand_x1_sg U63040 ( .A(n7174), .B(n7173), .X(n7171) );
  nor_x1_sg U63041 ( .A(n7173), .B(n7174), .X(n7172) );
  nand_x1_sg U63042 ( .A(n7993), .B(n7992), .X(n7990) );
  nor_x1_sg U63043 ( .A(n7992), .B(n7993), .X(n7991) );
  nand_x1_sg U63044 ( .A(n8811), .B(n8810), .X(n8808) );
  nor_x1_sg U63045 ( .A(n8810), .B(n8811), .X(n8809) );
  nand_x1_sg U63046 ( .A(n9631), .B(n9630), .X(n9628) );
  nor_x1_sg U63047 ( .A(n9630), .B(n9631), .X(n9629) );
  nand_x1_sg U63048 ( .A(n10450), .B(n10449), .X(n10447) );
  nor_x1_sg U63049 ( .A(n10449), .B(n10450), .X(n10448) );
  nand_x1_sg U63050 ( .A(n11269), .B(n11268), .X(n11266) );
  nor_x1_sg U63051 ( .A(n11268), .B(n11269), .X(n11267) );
  nand_x1_sg U63052 ( .A(n12088), .B(n12087), .X(n12085) );
  nor_x1_sg U63053 ( .A(n12087), .B(n12088), .X(n12086) );
  nand_x1_sg U63054 ( .A(n12907), .B(n12906), .X(n12904) );
  nor_x1_sg U63055 ( .A(n12906), .B(n12907), .X(n12905) );
  nand_x1_sg U63056 ( .A(n13726), .B(n13725), .X(n13723) );
  nor_x1_sg U63057 ( .A(n13725), .B(n13726), .X(n13724) );
  nand_x1_sg U63058 ( .A(n14545), .B(n14544), .X(n14542) );
  nor_x1_sg U63059 ( .A(n14544), .B(n14545), .X(n14543) );
  nand_x1_sg U63060 ( .A(n15364), .B(n15363), .X(n15361) );
  nor_x1_sg U63061 ( .A(n15363), .B(n15364), .X(n15362) );
  nand_x1_sg U63062 ( .A(n16183), .B(n16182), .X(n16180) );
  nor_x1_sg U63063 ( .A(n16182), .B(n16183), .X(n16181) );
  nand_x1_sg U63064 ( .A(n17821), .B(n17820), .X(n17818) );
  nor_x1_sg U63065 ( .A(n17820), .B(n17821), .X(n17819) );
  nand_x1_sg U63066 ( .A(n18642), .B(n18641), .X(n18639) );
  nor_x1_sg U63067 ( .A(n18641), .B(n18642), .X(n18640) );
  inv_x1_sg U63068 ( .A(n7469), .X(n46988) );
  inv_x1_sg U63069 ( .A(n17294), .X(n50418) );
  nand_x2_sg U63070 ( .A(n7295), .B(n7296), .X(n7294) );
  inv_x1_sg U63071 ( .A(n7272), .X(n46937) );
  nand_x2_sg U63072 ( .A(n8113), .B(n8114), .X(n8112) );
  inv_x1_sg U63073 ( .A(n8091), .X(n47229) );
  nand_x2_sg U63074 ( .A(n8931), .B(n8932), .X(n8930) );
  inv_x1_sg U63075 ( .A(n8909), .X(n47514) );
  nand_x2_sg U63076 ( .A(n9751), .B(n9752), .X(n9750) );
  inv_x1_sg U63077 ( .A(n9729), .X(n47799) );
  nand_x2_sg U63078 ( .A(n10570), .B(n10571), .X(n10569) );
  inv_x1_sg U63079 ( .A(n10548), .X(n48084) );
  nand_x2_sg U63080 ( .A(n11389), .B(n11390), .X(n11388) );
  inv_x1_sg U63081 ( .A(n11367), .X(n48369) );
  nand_x2_sg U63082 ( .A(n12208), .B(n12209), .X(n12207) );
  inv_x1_sg U63083 ( .A(n12186), .X(n48654) );
  nand_x2_sg U63084 ( .A(n13027), .B(n13028), .X(n13026) );
  inv_x1_sg U63085 ( .A(n13005), .X(n48940) );
  nand_x2_sg U63086 ( .A(n13846), .B(n13847), .X(n13845) );
  inv_x1_sg U63087 ( .A(n13824), .X(n49227) );
  nand_x2_sg U63088 ( .A(n14665), .B(n14666), .X(n14664) );
  inv_x1_sg U63089 ( .A(n14643), .X(n49513) );
  nand_x2_sg U63090 ( .A(n15484), .B(n15485), .X(n15483) );
  inv_x1_sg U63091 ( .A(n15462), .X(n49799) );
  nand_x2_sg U63092 ( .A(n16303), .B(n16304), .X(n16302) );
  inv_x1_sg U63093 ( .A(n16281), .X(n50085) );
  nand_x2_sg U63094 ( .A(n17120), .B(n17121), .X(n17119) );
  inv_x1_sg U63095 ( .A(n17097), .X(n50370) );
  nand_x2_sg U63096 ( .A(n17941), .B(n17942), .X(n17940) );
  inv_x1_sg U63097 ( .A(n17919), .X(n50659) );
  nand_x2_sg U63098 ( .A(n18762), .B(n18763), .X(n18761) );
  inv_x1_sg U63099 ( .A(n18740), .X(n50946) );
  inv_x1_sg U63100 ( .A(n8287), .X(n47277) );
  inv_x1_sg U63101 ( .A(n9105), .X(n47562) );
  inv_x1_sg U63102 ( .A(n9925), .X(n47847) );
  inv_x1_sg U63103 ( .A(n10744), .X(n48132) );
  inv_x1_sg U63104 ( .A(n11563), .X(n48417) );
  inv_x1_sg U63105 ( .A(n12382), .X(n48702) );
  inv_x1_sg U63106 ( .A(n13201), .X(n48988) );
  inv_x1_sg U63107 ( .A(n14020), .X(n49275) );
  inv_x1_sg U63108 ( .A(n14839), .X(n49561) );
  inv_x1_sg U63109 ( .A(n15658), .X(n49847) );
  inv_x1_sg U63110 ( .A(n16477), .X(n50133) );
  inv_x1_sg U63111 ( .A(n18115), .X(n50707) );
  inv_x1_sg U63112 ( .A(n18936), .X(n50994) );
  nand_x1_sg U63113 ( .A(n47332), .B(n47231), .X(n7776) );
  inv_x1_sg U63114 ( .A(n7779), .X(n47252) );
  nand_x1_sg U63115 ( .A(n47617), .B(n47516), .X(n8594) );
  inv_x1_sg U63116 ( .A(n8597), .X(n47537) );
  nand_x1_sg U63117 ( .A(n47902), .B(n47801), .X(n9414) );
  inv_x1_sg U63118 ( .A(n9417), .X(n47822) );
  nand_x1_sg U63119 ( .A(n48187), .B(n48086), .X(n10233) );
  inv_x1_sg U63120 ( .A(n10236), .X(n48107) );
  nand_x1_sg U63121 ( .A(n48472), .B(n48371), .X(n11052) );
  inv_x1_sg U63122 ( .A(n11055), .X(n48392) );
  nand_x1_sg U63123 ( .A(n48757), .B(n48656), .X(n11871) );
  inv_x1_sg U63124 ( .A(n11874), .X(n48677) );
  nand_x1_sg U63125 ( .A(n49043), .B(n48942), .X(n12690) );
  inv_x1_sg U63126 ( .A(n12693), .X(n48963) );
  nand_x1_sg U63127 ( .A(n49330), .B(n49229), .X(n13509) );
  inv_x1_sg U63128 ( .A(n13512), .X(n49250) );
  nand_x1_sg U63129 ( .A(n49616), .B(n49515), .X(n14328) );
  inv_x1_sg U63130 ( .A(n14331), .X(n49536) );
  nand_x1_sg U63131 ( .A(n49902), .B(n49801), .X(n15147) );
  inv_x1_sg U63132 ( .A(n15150), .X(n49822) );
  nand_x1_sg U63133 ( .A(n50188), .B(n50087), .X(n15966) );
  inv_x1_sg U63134 ( .A(n15969), .X(n50108) );
  nand_x1_sg U63135 ( .A(n50762), .B(n50661), .X(n17604) );
  inv_x1_sg U63136 ( .A(n17607), .X(n50682) );
  nand_x1_sg U63137 ( .A(n51049), .B(n50948), .X(n18425) );
  inv_x1_sg U63138 ( .A(n18428), .X(n50969) );
  nand_x1_sg U63139 ( .A(n8129), .B(n8130), .X(n8128) );
  nor_x1_sg U63140 ( .A(n8130), .B(n8129), .X(n8131) );
  nand_x1_sg U63141 ( .A(n8947), .B(n8948), .X(n8946) );
  nor_x1_sg U63142 ( .A(n8948), .B(n8947), .X(n8949) );
  nand_x1_sg U63143 ( .A(n9767), .B(n9768), .X(n9766) );
  nor_x1_sg U63144 ( .A(n9768), .B(n9767), .X(n9769) );
  nand_x1_sg U63145 ( .A(n10586), .B(n10587), .X(n10585) );
  nor_x1_sg U63146 ( .A(n10587), .B(n10586), .X(n10588) );
  nand_x1_sg U63147 ( .A(n11405), .B(n11406), .X(n11404) );
  nor_x1_sg U63148 ( .A(n11406), .B(n11405), .X(n11407) );
  nand_x1_sg U63149 ( .A(n12224), .B(n12225), .X(n12223) );
  nor_x1_sg U63150 ( .A(n12225), .B(n12224), .X(n12226) );
  nand_x1_sg U63151 ( .A(n13043), .B(n13044), .X(n13042) );
  nor_x1_sg U63152 ( .A(n13044), .B(n13043), .X(n13045) );
  nand_x1_sg U63153 ( .A(n13862), .B(n13863), .X(n13861) );
  nor_x1_sg U63154 ( .A(n13863), .B(n13862), .X(n13864) );
  nand_x1_sg U63155 ( .A(n14681), .B(n14682), .X(n14680) );
  nor_x1_sg U63156 ( .A(n14682), .B(n14681), .X(n14683) );
  nand_x1_sg U63157 ( .A(n15500), .B(n15501), .X(n15499) );
  nor_x1_sg U63158 ( .A(n15501), .B(n15500), .X(n15502) );
  nand_x1_sg U63159 ( .A(n16319), .B(n16320), .X(n16318) );
  nor_x1_sg U63160 ( .A(n16320), .B(n16319), .X(n16321) );
  nand_x1_sg U63161 ( .A(n17957), .B(n17958), .X(n17956) );
  nor_x1_sg U63162 ( .A(n17958), .B(n17957), .X(n17959) );
  nand_x1_sg U63163 ( .A(n18778), .B(n18779), .X(n18777) );
  nor_x1_sg U63164 ( .A(n18779), .B(n18778), .X(n18780) );
  nand_x1_sg U63165 ( .A(n7156), .B(n7157), .X(n7155) );
  nor_x1_sg U63166 ( .A(n7157), .B(n7156), .X(n7158) );
  nand_x1_sg U63167 ( .A(n16846), .B(n16847), .X(n16845) );
  nor_x1_sg U63168 ( .A(n16847), .B(n16846), .X(n16848) );
  nand_x1_sg U63169 ( .A(n7975), .B(n7976), .X(n7974) );
  nor_x1_sg U63170 ( .A(n7976), .B(n7975), .X(n7977) );
  nand_x1_sg U63171 ( .A(n8793), .B(n8794), .X(n8792) );
  nor_x1_sg U63172 ( .A(n8794), .B(n8793), .X(n8795) );
  nand_x1_sg U63173 ( .A(n9613), .B(n9614), .X(n9612) );
  nor_x1_sg U63174 ( .A(n9614), .B(n9613), .X(n9615) );
  nand_x1_sg U63175 ( .A(n10432), .B(n10433), .X(n10431) );
  nor_x1_sg U63176 ( .A(n10433), .B(n10432), .X(n10434) );
  nand_x1_sg U63177 ( .A(n11251), .B(n11252), .X(n11250) );
  nor_x1_sg U63178 ( .A(n11252), .B(n11251), .X(n11253) );
  nand_x1_sg U63179 ( .A(n12070), .B(n12071), .X(n12069) );
  nor_x1_sg U63180 ( .A(n12071), .B(n12070), .X(n12072) );
  nand_x1_sg U63181 ( .A(n12889), .B(n12890), .X(n12888) );
  nor_x1_sg U63182 ( .A(n12890), .B(n12889), .X(n12891) );
  nand_x1_sg U63183 ( .A(n13708), .B(n13709), .X(n13707) );
  nor_x1_sg U63184 ( .A(n13709), .B(n13708), .X(n13710) );
  nand_x1_sg U63185 ( .A(n14527), .B(n14528), .X(n14526) );
  nor_x1_sg U63186 ( .A(n14528), .B(n14527), .X(n14529) );
  nand_x1_sg U63187 ( .A(n15346), .B(n15347), .X(n15345) );
  nor_x1_sg U63188 ( .A(n15347), .B(n15346), .X(n15348) );
  nand_x1_sg U63189 ( .A(n16165), .B(n16166), .X(n16164) );
  nor_x1_sg U63190 ( .A(n16166), .B(n16165), .X(n16167) );
  nand_x1_sg U63191 ( .A(n16981), .B(n16982), .X(n16980) );
  nor_x1_sg U63192 ( .A(n16982), .B(n16981), .X(n16983) );
  nand_x1_sg U63193 ( .A(n17803), .B(n17804), .X(n17802) );
  nor_x1_sg U63194 ( .A(n17804), .B(n17803), .X(n17805) );
  nand_x1_sg U63195 ( .A(n18624), .B(n18625), .X(n18623) );
  nor_x1_sg U63196 ( .A(n18625), .B(n18624), .X(n18626) );
  nand_x1_sg U63197 ( .A(n7074), .B(n7075), .X(n7073) );
  nor_x1_sg U63198 ( .A(n7075), .B(n7074), .X(n7076) );
  nand_x1_sg U63199 ( .A(n7892), .B(n7893), .X(n7891) );
  nor_x1_sg U63200 ( .A(n7893), .B(n7892), .X(n7894) );
  nand_x1_sg U63201 ( .A(n8710), .B(n8711), .X(n8709) );
  nor_x1_sg U63202 ( .A(n8711), .B(n8710), .X(n8712) );
  nand_x1_sg U63203 ( .A(n9530), .B(n9531), .X(n9529) );
  nor_x1_sg U63204 ( .A(n9531), .B(n9530), .X(n9532) );
  nand_x1_sg U63205 ( .A(n10349), .B(n10350), .X(n10348) );
  nor_x1_sg U63206 ( .A(n10350), .B(n10349), .X(n10351) );
  nand_x1_sg U63207 ( .A(n11168), .B(n11169), .X(n11167) );
  nor_x1_sg U63208 ( .A(n11169), .B(n11168), .X(n11170) );
  nand_x1_sg U63209 ( .A(n11987), .B(n11988), .X(n11986) );
  nor_x1_sg U63210 ( .A(n11988), .B(n11987), .X(n11989) );
  nand_x1_sg U63211 ( .A(n12806), .B(n12807), .X(n12805) );
  nor_x1_sg U63212 ( .A(n12807), .B(n12806), .X(n12808) );
  nand_x1_sg U63213 ( .A(n13625), .B(n13626), .X(n13624) );
  nor_x1_sg U63214 ( .A(n13626), .B(n13625), .X(n13627) );
  nand_x1_sg U63215 ( .A(n14444), .B(n14445), .X(n14443) );
  nor_x1_sg U63216 ( .A(n14445), .B(n14444), .X(n14446) );
  nand_x1_sg U63217 ( .A(n15263), .B(n15264), .X(n15262) );
  nor_x1_sg U63218 ( .A(n15264), .B(n15263), .X(n15265) );
  nand_x1_sg U63219 ( .A(n16082), .B(n16083), .X(n16081) );
  nor_x1_sg U63220 ( .A(n16083), .B(n16082), .X(n16084) );
  nand_x1_sg U63221 ( .A(n16901), .B(n16902), .X(n16900) );
  nor_x1_sg U63222 ( .A(n16902), .B(n16901), .X(n16903) );
  nand_x1_sg U63223 ( .A(n17720), .B(n17721), .X(n17719) );
  nor_x1_sg U63224 ( .A(n17721), .B(n17720), .X(n17722) );
  nand_x1_sg U63225 ( .A(n18541), .B(n18542), .X(n18540) );
  nor_x1_sg U63226 ( .A(n18542), .B(n18541), .X(n18543) );
  nand_x4_sg U63227 ( .A(n51412), .B(n26320), .X(n26318) );
  nor_x1_sg U63228 ( .A(n50843), .B(n26321), .X(n26320) );
  nand_x1_sg U63229 ( .A(n26326), .B(n40225), .X(n26325) );
  nand_x1_sg U63230 ( .A(n40242), .B(n47136), .X(n22868) );
  nand_x1_sg U63231 ( .A(n40249), .B(n47421), .X(n23145) );
  nand_x1_sg U63232 ( .A(n40253), .B(n47706), .X(n23425) );
  nand_x1_sg U63233 ( .A(n40257), .B(n47991), .X(n23704) );
  nand_x1_sg U63234 ( .A(n40263), .B(n48276), .X(n23983) );
  nand_x1_sg U63235 ( .A(n40267), .B(n48561), .X(n24262) );
  nand_x1_sg U63236 ( .A(n40272), .B(n48846), .X(n24541) );
  nand_x1_sg U63237 ( .A(n40278), .B(n49133), .X(n24819) );
  nand_x1_sg U63238 ( .A(n40284), .B(n49419), .X(n25098) );
  nand_x1_sg U63239 ( .A(n40287), .B(n49705), .X(n25377) );
  nand_x1_sg U63240 ( .A(n40293), .B(n49991), .X(n25656) );
  nand_x1_sg U63241 ( .A(n40237), .B(n50566), .X(n26198) );
  nand_x1_sg U63242 ( .A(n40297), .B(n50852), .X(n26493) );
  nor_x1_sg U63243 ( .A(n40927), .B(n16649), .X(\L2_0/n2564 ) );
  nand_x1_sg U63244 ( .A(n7474), .B(n40163), .X(n7626) );
  nand_x1_sg U63245 ( .A(n39366), .B(n41191), .X(n22904) );
  nand_x1_sg U63246 ( .A(n39368), .B(n40504), .X(n23181) );
  nand_x1_sg U63247 ( .A(n39370), .B(n40499), .X(n23461) );
  nand_x1_sg U63248 ( .A(n39372), .B(n40495), .X(n23740) );
  nand_x1_sg U63249 ( .A(n39374), .B(n40492), .X(n24019) );
  nand_x1_sg U63250 ( .A(n39376), .B(n40487), .X(n24298) );
  nand_x1_sg U63251 ( .A(n39378), .B(n40484), .X(n24577) );
  nand_x1_sg U63252 ( .A(n39380), .B(n40479), .X(n24855) );
  nand_x1_sg U63253 ( .A(n39382), .B(n40476), .X(n25134) );
  nand_x1_sg U63254 ( .A(n39384), .B(n41146), .X(n25413) );
  nand_x1_sg U63255 ( .A(n39386), .B(n40467), .X(n25692) );
  nand_x1_sg U63256 ( .A(n39390), .B(n40464), .X(n26239) );
  nand_x1_sg U63257 ( .A(n39388), .B(n40461), .X(n26529) );
  nor_x1_sg U63258 ( .A(n40955), .B(n15849), .X(\L2_0/n2632 ) );
  nor_x1_sg U63259 ( .A(n40955), .B(n15868), .X(\L2_0/n2620 ) );
  nor_x1_sg U63260 ( .A(n38900), .B(n15874), .X(\L2_0/n2616 ) );
  nor_x1_sg U63261 ( .A(n38900), .B(n15886), .X(\L2_0/n2608 ) );
  nor_x1_sg U63262 ( .A(n38904), .B(n9297), .X(\L2_0/n3272 ) );
  nor_x1_sg U63263 ( .A(n40971), .B(n9316), .X(\L2_0/n3260 ) );
  nor_x1_sg U63264 ( .A(n9276), .B(n9322), .X(\L2_0/n3256 ) );
  nor_x1_sg U63265 ( .A(n38904), .B(n9334), .X(\L2_0/n3248 ) );
  nor_x1_sg U63266 ( .A(n40963), .B(n10116), .X(\L2_0/n3192 ) );
  nor_x1_sg U63267 ( .A(n40962), .B(n10135), .X(\L2_0/n3180 ) );
  nor_x1_sg U63268 ( .A(n40961), .B(n10141), .X(\L2_0/n3176 ) );
  nor_x1_sg U63269 ( .A(n10095), .B(n10153), .X(\L2_0/n3168 ) );
  nor_x1_sg U63270 ( .A(n40931), .B(n10935), .X(\L2_0/n3112 ) );
  nor_x1_sg U63271 ( .A(n40931), .B(n10954), .X(\L2_0/n3100 ) );
  nor_x1_sg U63272 ( .A(n38894), .B(n10960), .X(\L2_0/n3096 ) );
  nor_x1_sg U63273 ( .A(n38894), .B(n10972), .X(\L2_0/n3088 ) );
  nor_x1_sg U63274 ( .A(n40935), .B(n11754), .X(\L2_0/n3032 ) );
  nor_x1_sg U63275 ( .A(n40933), .B(n11773), .X(\L2_0/n3020 ) );
  nor_x1_sg U63276 ( .A(n40933), .B(n11779), .X(\L2_0/n3016 ) );
  nor_x1_sg U63277 ( .A(n40935), .B(n11791), .X(\L2_0/n3008 ) );
  nor_x1_sg U63278 ( .A(n40938), .B(n12573), .X(\L2_0/n2952 ) );
  nor_x1_sg U63279 ( .A(n40939), .B(n12592), .X(\L2_0/n2940 ) );
  nor_x1_sg U63280 ( .A(n40939), .B(n12598), .X(\L2_0/n2936 ) );
  nor_x1_sg U63281 ( .A(n38896), .B(n12610), .X(\L2_0/n2928 ) );
  nor_x1_sg U63282 ( .A(n40943), .B(n13392), .X(\L2_0/n2872 ) );
  nor_x1_sg U63283 ( .A(n40941), .B(n13411), .X(\L2_0/n2860 ) );
  nor_x1_sg U63284 ( .A(n38897), .B(n13417), .X(\L2_0/n2856 ) );
  nor_x1_sg U63285 ( .A(n40943), .B(n13429), .X(\L2_0/n2848 ) );
  nor_x1_sg U63286 ( .A(n40947), .B(n14211), .X(\L2_0/n2792 ) );
  nor_x1_sg U63287 ( .A(n40947), .B(n14230), .X(\L2_0/n2780 ) );
  nor_x1_sg U63288 ( .A(n38898), .B(n14236), .X(\L2_0/n2776 ) );
  nor_x1_sg U63289 ( .A(n38898), .B(n14248), .X(\L2_0/n2768 ) );
  nor_x1_sg U63290 ( .A(n40951), .B(n15030), .X(\L2_0/n2712 ) );
  nor_x1_sg U63291 ( .A(n40949), .B(n15049), .X(\L2_0/n2700 ) );
  nor_x1_sg U63292 ( .A(n40949), .B(n15055), .X(\L2_0/n2696 ) );
  nor_x1_sg U63293 ( .A(n40951), .B(n15067), .X(\L2_0/n2688 ) );
  nor_x1_sg U63294 ( .A(n40959), .B(n18308), .X(\L2_0/n2392 ) );
  nor_x1_sg U63295 ( .A(n40957), .B(n18327), .X(\L2_0/n2380 ) );
  nor_x1_sg U63296 ( .A(n40957), .B(n18333), .X(\L2_0/n2376 ) );
  nor_x1_sg U63297 ( .A(n40959), .B(n18345), .X(\L2_0/n2368 ) );
  nor_x1_sg U63298 ( .A(n39901), .B(n25651), .X(\L1_0/n3548 ) );
  nor_x1_sg U63299 ( .A(n39140), .B(n25672), .X(\L1_0/n3536 ) );
  nor_x1_sg U63300 ( .A(n41380), .B(n51405), .X(\L1_0/n3524 ) );
  inv_x1_sg U63301 ( .A(n25693), .X(n51405) );
  nor_x1_sg U63302 ( .A(n41383), .B(n25714), .X(\L1_0/n3512 ) );
  nor_x1_sg U63303 ( .A(n40035), .B(n51408), .X(\L1_0/n3500 ) );
  inv_x1_sg U63304 ( .A(n25735), .X(n51408) );
  nor_x1_sg U63305 ( .A(n40033), .B(n25754), .X(\L1_0/n3488 ) );
  nand_x1_sg U63306 ( .A(n42312), .B(n40164), .X(n7003) );
  nand_x1_sg U63307 ( .A(n39677), .B(n40244), .X(n7820) );
  nand_x1_sg U63308 ( .A(n39676), .B(n40249), .X(n8638) );
  nand_x1_sg U63309 ( .A(n39674), .B(n40255), .X(n9458) );
  nand_x1_sg U63310 ( .A(n39675), .B(n40258), .X(n10277) );
  nand_x1_sg U63311 ( .A(n39673), .B(n40264), .X(n11096) );
  nand_x1_sg U63312 ( .A(n39672), .B(n40270), .X(n11915) );
  nand_x1_sg U63313 ( .A(n39670), .B(n40273), .X(n12734) );
  nand_x1_sg U63314 ( .A(n39671), .B(n40277), .X(n13553) );
  nand_x1_sg U63315 ( .A(n39669), .B(n40284), .X(n14372) );
  nand_x1_sg U63316 ( .A(n39668), .B(n40288), .X(n15191) );
  nand_x1_sg U63317 ( .A(n39666), .B(n40294), .X(n16010) );
  nand_x1_sg U63318 ( .A(n39667), .B(n40240), .X(n17648) );
  nand_x1_sg U63319 ( .A(n39665), .B(n40300), .X(n18469) );
  nand_x1_sg U63320 ( .A(n39803), .B(n39663), .X(n7620) );
  nand_x1_sg U63321 ( .A(n39774), .B(n17299), .X(n17445) );
  nor_x1_sg U63322 ( .A(n38892), .B(n6825), .X(\L2_0/n3524 ) );
  nand_x1_sg U63323 ( .A(n8292), .B(n40245), .X(n8444) );
  nand_x1_sg U63324 ( .A(n9110), .B(n40250), .X(n9262) );
  nand_x1_sg U63325 ( .A(n9930), .B(n40252), .X(n10082) );
  nand_x1_sg U63326 ( .A(n39509), .B(n40260), .X(n10901) );
  nand_x1_sg U63327 ( .A(n11568), .B(n40262), .X(n11720) );
  nand_x1_sg U63328 ( .A(n12387), .B(n40270), .X(n12539) );
  nand_x1_sg U63329 ( .A(n13206), .B(n40275), .X(n13358) );
  nand_x1_sg U63330 ( .A(n39513), .B(n40279), .X(n14177) );
  nand_x1_sg U63331 ( .A(n14844), .B(n40285), .X(n14996) );
  nand_x1_sg U63332 ( .A(n15663), .B(n40290), .X(n15815) );
  nand_x1_sg U63333 ( .A(n16482), .B(n40292), .X(n16634) );
  nand_x1_sg U63334 ( .A(n18120), .B(n40237), .X(n18272) );
  nand_x1_sg U63335 ( .A(n39517), .B(n40300), .X(n19093) );
  inv_x1_sg U63336 ( .A(n7919), .X(n47158) );
  inv_x1_sg U63337 ( .A(n8737), .X(n47443) );
  inv_x1_sg U63338 ( .A(n9557), .X(n47728) );
  inv_x1_sg U63339 ( .A(n10376), .X(n48013) );
  inv_x1_sg U63340 ( .A(n11195), .X(n48298) );
  inv_x1_sg U63341 ( .A(n12014), .X(n48583) );
  inv_x1_sg U63342 ( .A(n12833), .X(n48869) );
  inv_x1_sg U63343 ( .A(n13652), .X(n49156) );
  inv_x1_sg U63344 ( .A(n14471), .X(n49442) );
  inv_x1_sg U63345 ( .A(n15290), .X(n49727) );
  inv_x1_sg U63346 ( .A(n16109), .X(n50014) );
  inv_x1_sg U63347 ( .A(n17747), .X(n50588) );
  inv_x1_sg U63348 ( .A(n18568), .X(n50875) );
  inv_x1_sg U63349 ( .A(n7340), .X(n46898) );
  inv_x1_sg U63350 ( .A(n17165), .X(n50331) );
  inv_x1_sg U63351 ( .A(n7101), .X(n46865) );
  inv_x1_sg U63352 ( .A(n16926), .X(n50298) );
  nand_x1_sg U63353 ( .A(n40988), .B(n45012), .X(n22527) );
  inv_x1_sg U63354 ( .A(n7087), .X(n46863) );
  inv_x1_sg U63355 ( .A(n7905), .X(n47156) );
  inv_x1_sg U63356 ( .A(n8723), .X(n47441) );
  inv_x1_sg U63357 ( .A(n9543), .X(n47726) );
  inv_x1_sg U63358 ( .A(n10362), .X(n48011) );
  inv_x1_sg U63359 ( .A(n11181), .X(n48296) );
  inv_x1_sg U63360 ( .A(n12000), .X(n48581) );
  inv_x1_sg U63361 ( .A(n12819), .X(n48867) );
  inv_x1_sg U63362 ( .A(n13638), .X(n49154) );
  inv_x1_sg U63363 ( .A(n14457), .X(n49440) );
  inv_x1_sg U63364 ( .A(n15276), .X(n49725) );
  inv_x1_sg U63365 ( .A(n16095), .X(n50012) );
  inv_x1_sg U63366 ( .A(n17733), .X(n50586) );
  inv_x1_sg U63367 ( .A(n18554), .X(n50873) );
  nand_x1_sg U63368 ( .A(n39798), .B(n39506), .X(n8438) );
  nand_x1_sg U63369 ( .A(n39801), .B(n39505), .X(n9256) );
  nand_x1_sg U63370 ( .A(n39794), .B(n39507), .X(n10076) );
  nand_x1_sg U63371 ( .A(n39797), .B(n10749), .X(n10895) );
  nand_x1_sg U63372 ( .A(n39790), .B(n39508), .X(n11714) );
  nand_x1_sg U63373 ( .A(n39793), .B(n39511), .X(n12533) );
  nand_x1_sg U63374 ( .A(n39786), .B(n39510), .X(n13352) );
  nand_x1_sg U63375 ( .A(n39789), .B(n14025), .X(n14171) );
  nand_x1_sg U63376 ( .A(n39782), .B(n39512), .X(n14990) );
  nand_x1_sg U63377 ( .A(n39785), .B(n39515), .X(n15809) );
  nand_x1_sg U63378 ( .A(n39778), .B(n39514), .X(n16628) );
  nand_x1_sg U63379 ( .A(n39781), .B(n39516), .X(n18266) );
  nand_x1_sg U63380 ( .A(n39777), .B(n18941), .X(n19087) );
  nor_x1_sg U63381 ( .A(n39903), .B(n23147), .X(\L1_0/n4264 ) );
  nor_x1_sg U63382 ( .A(n38978), .B(n23168), .X(\L1_0/n4252 ) );
  nor_x1_sg U63383 ( .A(n41375), .B(n23189), .X(\L1_0/n4240 ) );
  nor_x1_sg U63384 ( .A(n41376), .B(n51335), .X(\L1_0/n4228 ) );
  inv_x1_sg U63385 ( .A(n23210), .X(n51335) );
  nor_x1_sg U63386 ( .A(n38978), .B(n23231), .X(\L1_0/n4216 ) );
  nor_x1_sg U63387 ( .A(n39439), .B(n51339), .X(\L1_0/n4204 ) );
  inv_x1_sg U63388 ( .A(n23250), .X(n51339) );
  nor_x1_sg U63389 ( .A(n39457), .B(n23427), .X(\L1_0/n4184 ) );
  nor_x1_sg U63390 ( .A(n39915), .B(n23448), .X(\L1_0/n4172 ) );
  nor_x1_sg U63391 ( .A(n41346), .B(n23469), .X(\L1_0/n4160 ) );
  nor_x1_sg U63392 ( .A(n39458), .B(n51343), .X(\L1_0/n4148 ) );
  inv_x1_sg U63393 ( .A(n23490), .X(n51343) );
  nor_x1_sg U63394 ( .A(n41345), .B(n23511), .X(\L1_0/n4136 ) );
  nor_x1_sg U63395 ( .A(n39457), .B(n51347), .X(\L1_0/n4124 ) );
  inv_x1_sg U63396 ( .A(n23530), .X(n51347) );
  nor_x1_sg U63397 ( .A(n39917), .B(n23706), .X(\L1_0/n4104 ) );
  nor_x1_sg U63398 ( .A(n38957), .B(n23727), .X(\L1_0/n4092 ) );
  nor_x1_sg U63399 ( .A(n41342), .B(n23748), .X(\L1_0/n4080 ) );
  nor_x1_sg U63400 ( .A(n41342), .B(n51351), .X(\L1_0/n4068 ) );
  inv_x1_sg U63401 ( .A(n23769), .X(n51351) );
  nor_x1_sg U63402 ( .A(n41340), .B(n23790), .X(\L1_0/n4056 ) );
  nor_x1_sg U63403 ( .A(n41343), .B(n51355), .X(\L1_0/n4044 ) );
  inv_x1_sg U63404 ( .A(n23809), .X(n51355) );
  nor_x1_sg U63405 ( .A(n39448), .B(n23985), .X(\L1_0/n4024 ) );
  nor_x1_sg U63406 ( .A(n41361), .B(n24006), .X(\L1_0/n4012 ) );
  nor_x1_sg U63407 ( .A(n39908), .B(n24027), .X(\L1_0/n4000 ) );
  nor_x1_sg U63408 ( .A(n41360), .B(n51359), .X(\L1_0/n3988 ) );
  inv_x1_sg U63409 ( .A(n24048), .X(n51359) );
  nor_x1_sg U63410 ( .A(n39909), .B(n24069), .X(\L1_0/n3976 ) );
  nor_x1_sg U63411 ( .A(n39449), .B(n51363), .X(\L1_0/n3964 ) );
  inv_x1_sg U63412 ( .A(n24088), .X(n51363) );
  nor_x1_sg U63413 ( .A(n41355), .B(n24264), .X(\L1_0/n3944 ) );
  nor_x1_sg U63414 ( .A(n39911), .B(n24285), .X(\L1_0/n3932 ) );
  nor_x1_sg U63415 ( .A(n41356), .B(n24306), .X(\L1_0/n3920 ) );
  nor_x1_sg U63416 ( .A(n39451), .B(n51367), .X(\L1_0/n3908 ) );
  inv_x1_sg U63417 ( .A(n24327), .X(n51367) );
  nor_x1_sg U63418 ( .A(n39910), .B(n24348), .X(\L1_0/n3896 ) );
  nor_x1_sg U63419 ( .A(n41358), .B(n51371), .X(\L1_0/n3884 ) );
  inv_x1_sg U63420 ( .A(n24367), .X(n51371) );
  nor_x1_sg U63421 ( .A(n38954), .B(n24543), .X(\L1_0/n3864 ) );
  nor_x1_sg U63422 ( .A(n38954), .B(n24564), .X(\L1_0/n3852 ) );
  nor_x1_sg U63423 ( .A(n41336), .B(n24585), .X(\L1_0/n3840 ) );
  nor_x1_sg U63424 ( .A(n41337), .B(n51375), .X(\L1_0/n3828 ) );
  inv_x1_sg U63425 ( .A(n24606), .X(n51375) );
  nor_x1_sg U63426 ( .A(n41338), .B(n24627), .X(\L1_0/n3816 ) );
  nor_x1_sg U63427 ( .A(n41338), .B(n51379), .X(\L1_0/n3804 ) );
  inv_x1_sg U63428 ( .A(n24646), .X(n51379) );
  nor_x1_sg U63429 ( .A(n41333), .B(n24821), .X(\L1_0/n3784 ) );
  nor_x1_sg U63430 ( .A(n38951), .B(n24842), .X(\L1_0/n3772 ) );
  nor_x1_sg U63431 ( .A(n41332), .B(n24863), .X(\L1_0/n3760 ) );
  nor_x1_sg U63432 ( .A(n39921), .B(n51383), .X(\L1_0/n3748 ) );
  inv_x1_sg U63433 ( .A(n24884), .X(n51383) );
  nor_x1_sg U63434 ( .A(n41332), .B(n24905), .X(\L1_0/n3736 ) );
  nor_x1_sg U63435 ( .A(n41332), .B(n51387), .X(\L1_0/n3724 ) );
  inv_x1_sg U63436 ( .A(n24924), .X(n51387) );
  nor_x1_sg U63437 ( .A(n41326), .B(n25100), .X(\L1_0/n3704 ) );
  nor_x1_sg U63438 ( .A(n41328), .B(n25121), .X(\L1_0/n3692 ) );
  nor_x1_sg U63439 ( .A(n38949), .B(n25142), .X(\L1_0/n3680 ) );
  nor_x1_sg U63440 ( .A(n38948), .B(n51391), .X(\L1_0/n3668 ) );
  inv_x1_sg U63441 ( .A(n25163), .X(n51391) );
  nor_x1_sg U63442 ( .A(n39470), .B(n25184), .X(\L1_0/n3656 ) );
  nor_x1_sg U63443 ( .A(n38949), .B(n51395), .X(\L1_0/n3644 ) );
  inv_x1_sg U63444 ( .A(n25203), .X(n51395) );
  nor_x1_sg U63445 ( .A(n39905), .B(n25379), .X(\L1_0/n3624 ) );
  nor_x1_sg U63446 ( .A(n39442), .B(n25400), .X(\L1_0/n3612 ) );
  nor_x1_sg U63447 ( .A(n41370), .B(n25421), .X(\L1_0/n3600 ) );
  nor_x1_sg U63448 ( .A(n41371), .B(n51399), .X(\L1_0/n3588 ) );
  inv_x1_sg U63449 ( .A(n25442), .X(n51399) );
  nor_x1_sg U63450 ( .A(n38975), .B(n25463), .X(\L1_0/n3576 ) );
  nor_x1_sg U63451 ( .A(n41371), .B(n51403), .X(\L1_0/n3564 ) );
  inv_x1_sg U63452 ( .A(n25482), .X(n51403) );
  nor_x1_sg U63453 ( .A(n41383), .B(n25658), .X(\L1_0/n3544 ) );
  nor_x1_sg U63454 ( .A(n41383), .B(n25679), .X(\L1_0/n3532 ) );
  nor_x1_sg U63455 ( .A(n40034), .B(n25700), .X(\L1_0/n3520 ) );
  nor_x1_sg U63456 ( .A(n41381), .B(n51407), .X(\L1_0/n3508 ) );
  inv_x1_sg U63457 ( .A(n25721), .X(n51407) );
  nor_x1_sg U63458 ( .A(n39139), .B(n25742), .X(\L1_0/n3496 ) );
  nor_x1_sg U63459 ( .A(n39140), .B(n51411), .X(\L1_0/n3484 ) );
  inv_x1_sg U63460 ( .A(n25761), .X(n51411) );
  nor_x1_sg U63461 ( .A(n39454), .B(n26495), .X(\L1_0/n3304 ) );
  nor_x1_sg U63462 ( .A(n38964), .B(n26516), .X(\L1_0/n3292 ) );
  nor_x1_sg U63463 ( .A(n39913), .B(n26537), .X(\L1_0/n3280 ) );
  nor_x1_sg U63464 ( .A(n38963), .B(n51416), .X(\L1_0/n3268 ) );
  inv_x1_sg U63465 ( .A(n26558), .X(n51416) );
  nor_x1_sg U63466 ( .A(n38964), .B(n26579), .X(\L1_0/n3256 ) );
  nor_x1_sg U63467 ( .A(n39912), .B(n51420), .X(\L1_0/n3244 ) );
  inv_x1_sg U63468 ( .A(n26598), .X(n51420) );
  inv_x1_sg U63469 ( .A(n16913), .X(n50296) );
  nor_x1_sg U63470 ( .A(n7618), .B(n7619), .X(n7617) );
  nor_x1_sg U63471 ( .A(n7620), .B(n46856), .X(n7619) );
  nor_x1_sg U63472 ( .A(n7621), .B(n39605), .X(n7618) );
  nor_x1_sg U63473 ( .A(n17443), .B(n17444), .X(n17442) );
  nor_x1_sg U63474 ( .A(n17445), .B(n50288), .X(n17444) );
  nor_x1_sg U63475 ( .A(n17446), .B(n39602), .X(n17443) );
  nand_x1_sg U63476 ( .A(n8035), .B(n40508), .X(n22911) );
  nand_x1_sg U63477 ( .A(n40108), .B(n41186), .X(n23188) );
  nand_x1_sg U63478 ( .A(n9673), .B(n41181), .X(n23468) );
  nand_x1_sg U63479 ( .A(n40112), .B(n40496), .X(n23747) );
  nand_x1_sg U63480 ( .A(n40114), .B(n40493), .X(n24026) );
  nand_x1_sg U63481 ( .A(n12130), .B(n39231), .X(n24305) );
  nand_x1_sg U63482 ( .A(n40118), .B(n40484), .X(n24584) );
  nand_x1_sg U63483 ( .A(n40119), .B(n40481), .X(n24862) );
  nand_x1_sg U63484 ( .A(n14587), .B(n40477), .X(n25141) );
  nand_x1_sg U63485 ( .A(n15406), .B(n40472), .X(n25420) );
  nand_x1_sg U63486 ( .A(n40126), .B(n40468), .X(n25699) );
  nand_x1_sg U63487 ( .A(n40131), .B(n41136), .X(n26247) );
  nand_x1_sg U63488 ( .A(n18684), .B(n40459), .X(n26536) );
  nor_x1_sg U63489 ( .A(n8436), .B(n8437), .X(n8435) );
  nor_x1_sg U63490 ( .A(n8438), .B(n47149), .X(n8437) );
  nor_x1_sg U63491 ( .A(n8439), .B(n41657), .X(n8436) );
  nor_x1_sg U63492 ( .A(n9254), .B(n9255), .X(n9253) );
  nor_x1_sg U63493 ( .A(n9256), .B(n47434), .X(n9255) );
  nor_x1_sg U63494 ( .A(n9257), .B(n39733), .X(n9254) );
  nor_x1_sg U63495 ( .A(n10074), .B(n10075), .X(n10073) );
  nor_x1_sg U63496 ( .A(n10076), .B(n47719), .X(n10075) );
  nor_x1_sg U63497 ( .A(n10077), .B(n39736), .X(n10074) );
  nor_x1_sg U63498 ( .A(n10893), .B(n10894), .X(n10892) );
  nor_x1_sg U63499 ( .A(n10895), .B(n48004), .X(n10894) );
  nor_x1_sg U63500 ( .A(n10896), .B(n41650), .X(n10893) );
  nor_x1_sg U63501 ( .A(n11712), .B(n11713), .X(n11711) );
  nor_x1_sg U63502 ( .A(n11714), .B(n48289), .X(n11713) );
  nor_x1_sg U63503 ( .A(n11715), .B(n39742), .X(n11712) );
  nor_x1_sg U63504 ( .A(n12531), .B(n12532), .X(n12530) );
  nor_x1_sg U63505 ( .A(n12533), .B(n48574), .X(n12532) );
  nor_x1_sg U63506 ( .A(n12534), .B(n41648), .X(n12531) );
  nor_x1_sg U63507 ( .A(n13350), .B(n13351), .X(n13349) );
  nor_x1_sg U63508 ( .A(n13352), .B(n48860), .X(n13351) );
  nor_x1_sg U63509 ( .A(n13353), .B(n39748), .X(n13350) );
  nor_x1_sg U63510 ( .A(n14169), .B(n14170), .X(n14168) );
  nor_x1_sg U63511 ( .A(n14171), .B(n49147), .X(n14170) );
  nor_x1_sg U63512 ( .A(n14172), .B(n39751), .X(n14169) );
  nor_x1_sg U63513 ( .A(n14988), .B(n14989), .X(n14987) );
  nor_x1_sg U63514 ( .A(n14990), .B(n49433), .X(n14989) );
  nor_x1_sg U63515 ( .A(n14991), .B(n41653), .X(n14988) );
  nor_x1_sg U63516 ( .A(n15807), .B(n15808), .X(n15806) );
  nor_x1_sg U63517 ( .A(n15809), .B(n49718), .X(n15808) );
  nor_x1_sg U63518 ( .A(n15810), .B(n39757), .X(n15807) );
  nor_x1_sg U63519 ( .A(n16626), .B(n16627), .X(n16625) );
  nor_x1_sg U63520 ( .A(n16628), .B(n50005), .X(n16627) );
  nor_x1_sg U63521 ( .A(n16629), .B(n41659), .X(n16626) );
  nor_x1_sg U63522 ( .A(n18264), .B(n18265), .X(n18263) );
  nor_x1_sg U63523 ( .A(n18266), .B(n50579), .X(n18265) );
  nor_x1_sg U63524 ( .A(n18267), .B(n41647), .X(n18264) );
  nor_x1_sg U63525 ( .A(n19085), .B(n19086), .X(n19084) );
  nor_x1_sg U63526 ( .A(n19087), .B(n50866), .X(n19086) );
  nor_x1_sg U63527 ( .A(n19088), .B(n41658), .X(n19085) );
  nand_x1_sg U63528 ( .A(n16966), .B(n41603), .X(n16965) );
  inv_x1_sg U63529 ( .A(n8158), .X(n47193) );
  inv_x1_sg U63530 ( .A(n8976), .X(n47478) );
  inv_x1_sg U63531 ( .A(n9796), .X(n47763) );
  inv_x1_sg U63532 ( .A(n10615), .X(n48048) );
  inv_x1_sg U63533 ( .A(n11434), .X(n48333) );
  inv_x1_sg U63534 ( .A(n12253), .X(n48618) );
  inv_x1_sg U63535 ( .A(n13072), .X(n48904) );
  inv_x1_sg U63536 ( .A(n13891), .X(n49191) );
  inv_x1_sg U63537 ( .A(n14710), .X(n49477) );
  inv_x1_sg U63538 ( .A(n15529), .X(n49763) );
  inv_x1_sg U63539 ( .A(n16348), .X(n50049) );
  inv_x1_sg U63540 ( .A(n17986), .X(n50623) );
  inv_x1_sg U63541 ( .A(n18807), .X(n50910) );
  nor_x1_sg U63542 ( .A(n39440), .B(n23132), .X(\L1_0/n4272 ) );
  nor_x1_sg U63543 ( .A(n38979), .B(n23140), .X(\L1_0/n4268 ) );
  nor_x1_sg U63544 ( .A(n39903), .B(n23154), .X(\L1_0/n4260 ) );
  nor_x1_sg U63545 ( .A(n41377), .B(n23161), .X(\L1_0/n4256 ) );
  nor_x1_sg U63546 ( .A(n39902), .B(n51332), .X(\L1_0/n4248 ) );
  inv_x1_sg U63547 ( .A(n23175), .X(n51332) );
  nor_x1_sg U63548 ( .A(n41378), .B(n51333), .X(\L1_0/n4244 ) );
  inv_x1_sg U63549 ( .A(n23182), .X(n51333) );
  nor_x1_sg U63550 ( .A(n41376), .B(n51334), .X(\L1_0/n4236 ) );
  inv_x1_sg U63551 ( .A(n23196), .X(n51334) );
  nor_x1_sg U63552 ( .A(n38979), .B(n23203), .X(\L1_0/n4232 ) );
  nor_x1_sg U63553 ( .A(n41375), .B(n23217), .X(\L1_0/n4224 ) );
  nor_x1_sg U63554 ( .A(n39902), .B(n51336), .X(\L1_0/n4220 ) );
  inv_x1_sg U63555 ( .A(n23224), .X(n51336) );
  nor_x1_sg U63556 ( .A(n41375), .B(n23238), .X(\L1_0/n4212 ) );
  nor_x1_sg U63557 ( .A(n38979), .B(n23243), .X(\L1_0/n4208 ) );
  nor_x1_sg U63558 ( .A(n41345), .B(n23412), .X(\L1_0/n4192 ) );
  nor_x1_sg U63559 ( .A(n39914), .B(n23420), .X(\L1_0/n4188 ) );
  nor_x1_sg U63560 ( .A(n39458), .B(n23434), .X(\L1_0/n4180 ) );
  nor_x1_sg U63561 ( .A(n39915), .B(n23441), .X(\L1_0/n4176 ) );
  nor_x1_sg U63562 ( .A(n41348), .B(n51340), .X(\L1_0/n4168 ) );
  inv_x1_sg U63563 ( .A(n23455), .X(n51340) );
  nor_x1_sg U63564 ( .A(n41345), .B(n51341), .X(\L1_0/n4164 ) );
  inv_x1_sg U63565 ( .A(n23462), .X(n51341) );
  nor_x1_sg U63566 ( .A(n39458), .B(n51342), .X(\L1_0/n4156 ) );
  inv_x1_sg U63567 ( .A(n23476), .X(n51342) );
  nor_x1_sg U63568 ( .A(n41346), .B(n23483), .X(\L1_0/n4152 ) );
  nor_x1_sg U63569 ( .A(n41346), .B(n23497), .X(\L1_0/n4144 ) );
  nor_x1_sg U63570 ( .A(n41345), .B(n51344), .X(\L1_0/n4140 ) );
  inv_x1_sg U63571 ( .A(n23504), .X(n51344) );
  nor_x1_sg U63572 ( .A(n38961), .B(n23518), .X(\L1_0/n4132 ) );
  nor_x1_sg U63573 ( .A(n39915), .B(n23523), .X(\L1_0/n4128 ) );
  nor_x1_sg U63574 ( .A(n39917), .B(n23691), .X(\L1_0/n4112 ) );
  nor_x1_sg U63575 ( .A(n39461), .B(n23699), .X(\L1_0/n4108 ) );
  nor_x1_sg U63576 ( .A(n38958), .B(n23713), .X(\L1_0/n4100 ) );
  nor_x1_sg U63577 ( .A(n41340), .B(n23720), .X(\L1_0/n4096 ) );
  nor_x1_sg U63578 ( .A(n41340), .B(n51348), .X(\L1_0/n4088 ) );
  inv_x1_sg U63579 ( .A(n23734), .X(n51348) );
  nor_x1_sg U63580 ( .A(n41342), .B(n51349), .X(\L1_0/n4084 ) );
  inv_x1_sg U63581 ( .A(n23741), .X(n51349) );
  nor_x1_sg U63582 ( .A(n41341), .B(n51350), .X(\L1_0/n4076 ) );
  inv_x1_sg U63583 ( .A(n23755), .X(n51350) );
  nor_x1_sg U63584 ( .A(n41341), .B(n23762), .X(\L1_0/n4072 ) );
  nor_x1_sg U63585 ( .A(n38958), .B(n23776), .X(\L1_0/n4064 ) );
  nor_x1_sg U63586 ( .A(n39916), .B(n51352), .X(\L1_0/n4060 ) );
  inv_x1_sg U63587 ( .A(n23783), .X(n51352) );
  nor_x1_sg U63588 ( .A(n39916), .B(n23797), .X(\L1_0/n4052 ) );
  nor_x1_sg U63589 ( .A(n38957), .B(n23802), .X(\L1_0/n4048 ) );
  nor_x1_sg U63590 ( .A(n38970), .B(n23970), .X(\L1_0/n4032 ) );
  nor_x1_sg U63591 ( .A(n41362), .B(n23978), .X(\L1_0/n4028 ) );
  nor_x1_sg U63592 ( .A(n39908), .B(n23992), .X(\L1_0/n4020 ) );
  nor_x1_sg U63593 ( .A(n38970), .B(n23999), .X(\L1_0/n4016 ) );
  nor_x1_sg U63594 ( .A(n41362), .B(n51356), .X(\L1_0/n4008 ) );
  inv_x1_sg U63595 ( .A(n24013), .X(n51356) );
  nor_x1_sg U63596 ( .A(n39909), .B(n51357), .X(\L1_0/n4004 ) );
  inv_x1_sg U63597 ( .A(n24020), .X(n51357) );
  nor_x1_sg U63598 ( .A(n38969), .B(n51358), .X(\L1_0/n3996 ) );
  inv_x1_sg U63599 ( .A(n24034), .X(n51358) );
  nor_x1_sg U63600 ( .A(n38970), .B(n24041), .X(\L1_0/n3992 ) );
  nor_x1_sg U63601 ( .A(n41363), .B(n24055), .X(\L1_0/n3984 ) );
  nor_x1_sg U63602 ( .A(n41363), .B(n51360), .X(\L1_0/n3980 ) );
  inv_x1_sg U63603 ( .A(n24062), .X(n51360) );
  nor_x1_sg U63604 ( .A(n41361), .B(n24076), .X(\L1_0/n3972 ) );
  nor_x1_sg U63605 ( .A(n41362), .B(n24081), .X(\L1_0/n3968 ) );
  nor_x1_sg U63606 ( .A(n38966), .B(n24249), .X(\L1_0/n3952 ) );
  nor_x1_sg U63607 ( .A(n39911), .B(n24257), .X(\L1_0/n3948 ) );
  nor_x1_sg U63608 ( .A(n41356), .B(n24271), .X(\L1_0/n3940 ) );
  nor_x1_sg U63609 ( .A(n39911), .B(n24278), .X(\L1_0/n3936 ) );
  nor_x1_sg U63610 ( .A(n38967), .B(n51364), .X(\L1_0/n3928 ) );
  inv_x1_sg U63611 ( .A(n24292), .X(n51364) );
  nor_x1_sg U63612 ( .A(n38967), .B(n51365), .X(\L1_0/n3924 ) );
  inv_x1_sg U63613 ( .A(n24299), .X(n51365) );
  nor_x1_sg U63614 ( .A(n39452), .B(n51366), .X(\L1_0/n3916 ) );
  inv_x1_sg U63615 ( .A(n24313), .X(n51366) );
  nor_x1_sg U63616 ( .A(n41355), .B(n24320), .X(\L1_0/n3912 ) );
  nor_x1_sg U63617 ( .A(n39452), .B(n24334), .X(\L1_0/n3904 ) );
  nor_x1_sg U63618 ( .A(n39452), .B(n51368), .X(\L1_0/n3900 ) );
  inv_x1_sg U63619 ( .A(n24341), .X(n51368) );
  nor_x1_sg U63620 ( .A(n39911), .B(n24355), .X(\L1_0/n3892 ) );
  nor_x1_sg U63621 ( .A(n41355), .B(n24360), .X(\L1_0/n3888 ) );
  nor_x1_sg U63622 ( .A(n39918), .B(n24528), .X(\L1_0/n3872 ) );
  nor_x1_sg U63623 ( .A(n41337), .B(n24536), .X(\L1_0/n3868 ) );
  nor_x1_sg U63624 ( .A(n39919), .B(n24550), .X(\L1_0/n3860 ) );
  nor_x1_sg U63625 ( .A(n39919), .B(n24557), .X(\L1_0/n3856 ) );
  nor_x1_sg U63626 ( .A(n38955), .B(n51372), .X(\L1_0/n3848 ) );
  inv_x1_sg U63627 ( .A(n24571), .X(n51372) );
  nor_x1_sg U63628 ( .A(n41336), .B(n51373), .X(\L1_0/n3844 ) );
  inv_x1_sg U63629 ( .A(n24578), .X(n51373) );
  nor_x1_sg U63630 ( .A(n39464), .B(n51374), .X(\L1_0/n3836 ) );
  inv_x1_sg U63631 ( .A(n24592), .X(n51374) );
  nor_x1_sg U63632 ( .A(n41337), .B(n24599), .X(\L1_0/n3832 ) );
  nor_x1_sg U63633 ( .A(n41335), .B(n24613), .X(\L1_0/n3824 ) );
  nor_x1_sg U63634 ( .A(n41336), .B(n51376), .X(\L1_0/n3820 ) );
  inv_x1_sg U63635 ( .A(n24620), .X(n51376) );
  nor_x1_sg U63636 ( .A(n38955), .B(n24634), .X(\L1_0/n3812 ) );
  nor_x1_sg U63637 ( .A(n41336), .B(n24639), .X(\L1_0/n3808 ) );
  nor_x1_sg U63638 ( .A(n39466), .B(n24806), .X(\L1_0/n3792 ) );
  nor_x1_sg U63639 ( .A(n39466), .B(n24814), .X(\L1_0/n3788 ) );
  nor_x1_sg U63640 ( .A(n39467), .B(n24828), .X(\L1_0/n3780 ) );
  nor_x1_sg U63641 ( .A(n41331), .B(n24835), .X(\L1_0/n3776 ) );
  nor_x1_sg U63642 ( .A(n38952), .B(n51380), .X(\L1_0/n3768 ) );
  inv_x1_sg U63643 ( .A(n24849), .X(n51380) );
  nor_x1_sg U63644 ( .A(n39920), .B(n51381), .X(\L1_0/n3764 ) );
  inv_x1_sg U63645 ( .A(n24856), .X(n51381) );
  nor_x1_sg U63646 ( .A(n41331), .B(n51382), .X(\L1_0/n3756 ) );
  inv_x1_sg U63647 ( .A(n24870), .X(n51382) );
  nor_x1_sg U63648 ( .A(n39467), .B(n24877), .X(\L1_0/n3752 ) );
  nor_x1_sg U63649 ( .A(n38952), .B(n24891), .X(\L1_0/n3744 ) );
  nor_x1_sg U63650 ( .A(n39920), .B(n51384), .X(\L1_0/n3740 ) );
  inv_x1_sg U63651 ( .A(n24898), .X(n51384) );
  nor_x1_sg U63652 ( .A(n39920), .B(n24912), .X(\L1_0/n3732 ) );
  nor_x1_sg U63653 ( .A(n39466), .B(n24917), .X(\L1_0/n3728 ) );
  nor_x1_sg U63654 ( .A(n41328), .B(n25085), .X(\L1_0/n3712 ) );
  nor_x1_sg U63655 ( .A(n41326), .B(n25093), .X(\L1_0/n3708 ) );
  nor_x1_sg U63656 ( .A(n41325), .B(n25107), .X(\L1_0/n3700 ) );
  nor_x1_sg U63657 ( .A(n39469), .B(n25114), .X(\L1_0/n3696 ) );
  nor_x1_sg U63658 ( .A(n39923), .B(n51388), .X(\L1_0/n3688 ) );
  inv_x1_sg U63659 ( .A(n25128), .X(n51388) );
  nor_x1_sg U63660 ( .A(n39470), .B(n51389), .X(\L1_0/n3684 ) );
  inv_x1_sg U63661 ( .A(n25135), .X(n51389) );
  nor_x1_sg U63662 ( .A(n41326), .B(n51390), .X(\L1_0/n3676 ) );
  inv_x1_sg U63663 ( .A(n25149), .X(n51390) );
  nor_x1_sg U63664 ( .A(n39470), .B(n25156), .X(\L1_0/n3672 ) );
  nor_x1_sg U63665 ( .A(n39470), .B(n25170), .X(\L1_0/n3664 ) );
  nor_x1_sg U63666 ( .A(n39922), .B(n51392), .X(\L1_0/n3660 ) );
  inv_x1_sg U63667 ( .A(n25177), .X(n51392) );
  nor_x1_sg U63668 ( .A(n39469), .B(n25191), .X(\L1_0/n3652 ) );
  nor_x1_sg U63669 ( .A(n39469), .B(n25196), .X(\L1_0/n3648 ) );
  nor_x1_sg U63670 ( .A(n38976), .B(n25364), .X(\L1_0/n3632 ) );
  nor_x1_sg U63671 ( .A(n39442), .B(n25372), .X(\L1_0/n3628 ) );
  nor_x1_sg U63672 ( .A(n41373), .B(n25386), .X(\L1_0/n3620 ) );
  nor_x1_sg U63673 ( .A(n38976), .B(n25393), .X(\L1_0/n3616 ) );
  nor_x1_sg U63674 ( .A(n39443), .B(n51396), .X(\L1_0/n3608 ) );
  inv_x1_sg U63675 ( .A(n25407), .X(n51396) );
  nor_x1_sg U63676 ( .A(n41372), .B(n51397), .X(\L1_0/n3604 ) );
  inv_x1_sg U63677 ( .A(n25414), .X(n51397) );
  nor_x1_sg U63678 ( .A(n39905), .B(n51398), .X(\L1_0/n3596 ) );
  inv_x1_sg U63679 ( .A(n25428), .X(n51398) );
  nor_x1_sg U63680 ( .A(n41370), .B(n25435), .X(\L1_0/n3592 ) );
  nor_x1_sg U63681 ( .A(n41371), .B(n25449), .X(\L1_0/n3584 ) );
  nor_x1_sg U63682 ( .A(n41370), .B(n51400), .X(\L1_0/n3580 ) );
  inv_x1_sg U63683 ( .A(n25456), .X(n51400) );
  nor_x1_sg U63684 ( .A(n41370), .B(n25470), .X(\L1_0/n3572 ) );
  nor_x1_sg U63685 ( .A(n39904), .B(n25475), .X(\L1_0/n3568 ) );
  nor_x1_sg U63686 ( .A(n25640), .B(n25643), .X(\L1_0/n3552 ) );
  nor_x1_sg U63687 ( .A(n41382), .B(n25665), .X(\L1_0/n3540 ) );
  nor_x1_sg U63688 ( .A(n40033), .B(n51404), .X(\L1_0/n3528 ) );
  inv_x1_sg U63689 ( .A(n25686), .X(n51404) );
  nor_x1_sg U63690 ( .A(n39140), .B(n51406), .X(\L1_0/n3516 ) );
  inv_x1_sg U63691 ( .A(n25707), .X(n51406) );
  nor_x1_sg U63692 ( .A(n41380), .B(n25728), .X(\L1_0/n3504 ) );
  nor_x1_sg U63693 ( .A(n25640), .B(n25749), .X(\L1_0/n3492 ) );
  nor_x1_sg U63694 ( .A(n38963), .B(n26480), .X(\L1_0/n3312 ) );
  nor_x1_sg U63695 ( .A(n41350), .B(n26488), .X(\L1_0/n3308 ) );
  nor_x1_sg U63696 ( .A(n38964), .B(n26502), .X(\L1_0/n3300 ) );
  nor_x1_sg U63697 ( .A(n39912), .B(n26509), .X(\L1_0/n3296 ) );
  nor_x1_sg U63698 ( .A(n39454), .B(n51413), .X(\L1_0/n3288 ) );
  inv_x1_sg U63699 ( .A(n26523), .X(n51413) );
  nor_x1_sg U63700 ( .A(n39454), .B(n51414), .X(\L1_0/n3284 ) );
  inv_x1_sg U63701 ( .A(n26530), .X(n51414) );
  nor_x1_sg U63702 ( .A(n39455), .B(n51415), .X(\L1_0/n3276 ) );
  inv_x1_sg U63703 ( .A(n26544), .X(n51415) );
  nor_x1_sg U63704 ( .A(n41350), .B(n26551), .X(\L1_0/n3272 ) );
  nor_x1_sg U63705 ( .A(n41353), .B(n26565), .X(\L1_0/n3264 ) );
  nor_x1_sg U63706 ( .A(n39913), .B(n51417), .X(\L1_0/n3260 ) );
  inv_x1_sg U63707 ( .A(n26572), .X(n51417) );
  nor_x1_sg U63708 ( .A(n41351), .B(n26586), .X(\L1_0/n3252 ) );
  nor_x1_sg U63709 ( .A(n39912), .B(n26591), .X(\L1_0/n3248 ) );
  inv_x1_sg U63710 ( .A(n7496), .X(n47021) );
  inv_x1_sg U63711 ( .A(n8314), .X(n47309) );
  inv_x1_sg U63712 ( .A(n9132), .X(n47594) );
  inv_x1_sg U63713 ( .A(n9952), .X(n47879) );
  inv_x1_sg U63714 ( .A(n10771), .X(n48164) );
  inv_x1_sg U63715 ( .A(n11590), .X(n48449) );
  inv_x1_sg U63716 ( .A(n12409), .X(n48734) );
  inv_x1_sg U63717 ( .A(n13228), .X(n49020) );
  inv_x1_sg U63718 ( .A(n14047), .X(n49307) );
  inv_x1_sg U63719 ( .A(n14866), .X(n49593) );
  inv_x1_sg U63720 ( .A(n15685), .X(n49879) );
  inv_x1_sg U63721 ( .A(n16504), .X(n50165) );
  inv_x1_sg U63722 ( .A(n17321), .X(n50450) );
  inv_x1_sg U63723 ( .A(n18142), .X(n50739) );
  inv_x1_sg U63724 ( .A(n18963), .X(n51026) );
  inv_x1_sg U63725 ( .A(n26329), .X(n50843) );
  nand_x1_sg U63726 ( .A(n40508), .B(n39611), .X(n22925) );
  nand_x1_sg U63727 ( .A(n39223), .B(n39608), .X(n23202) );
  nand_x1_sg U63728 ( .A(n40501), .B(n39627), .X(n23482) );
  nand_x1_sg U63729 ( .A(n39227), .B(n39624), .X(n23761) );
  nand_x1_sg U63730 ( .A(n40491), .B(n39621), .X(n24040) );
  nand_x1_sg U63731 ( .A(n40488), .B(n39618), .X(n24319) );
  nand_x1_sg U63732 ( .A(n39233), .B(n39639), .X(n24598) );
  nand_x1_sg U63733 ( .A(n39235), .B(n39635), .X(n24876) );
  nand_x1_sg U63734 ( .A(n40475), .B(n39632), .X(n25155) );
  nand_x1_sg U63735 ( .A(n39239), .B(n39629), .X(n25434) );
  nand_x1_sg U63736 ( .A(n40468), .B(n39647), .X(n25713) );
  nand_x1_sg U63737 ( .A(n40465), .B(n39644), .X(n26263) );
  nand_x1_sg U63738 ( .A(n41131), .B(n39641), .X(n26550) );
  nand_x1_sg U63739 ( .A(n41901), .B(n40081), .X(n7285) );
  nand_x1_sg U63740 ( .A(n40611), .B(n40077), .X(n17110) );
  nand_x1_sg U63741 ( .A(n41304), .B(n46845), .X(n22606) );
  nand_x1_sg U63742 ( .A(n41307), .B(n22635), .X(n22644) );
  inv_x1_sg U63743 ( .A(n8003), .X(n47180) );
  inv_x1_sg U63744 ( .A(n8821), .X(n47465) );
  inv_x1_sg U63745 ( .A(n9641), .X(n47750) );
  inv_x1_sg U63746 ( .A(n10460), .X(n48035) );
  inv_x1_sg U63747 ( .A(n11279), .X(n48320) );
  inv_x1_sg U63748 ( .A(n12098), .X(n48605) );
  inv_x1_sg U63749 ( .A(n12917), .X(n48891) );
  inv_x1_sg U63750 ( .A(n13736), .X(n49178) );
  inv_x1_sg U63751 ( .A(n14555), .X(n49464) );
  inv_x1_sg U63752 ( .A(n15374), .X(n49749) );
  inv_x1_sg U63753 ( .A(n16193), .X(n50036) );
  inv_x1_sg U63754 ( .A(n17831), .X(n50610) );
  inv_x1_sg U63755 ( .A(n18652), .X(n50897) );
  inv_x1_sg U63756 ( .A(n7184), .X(n46887) );
  inv_x1_sg U63757 ( .A(n17009), .X(n50321) );
  nand_x1_sg U63758 ( .A(n47081), .B(n39805), .X(n7032) );
  nand_x1_sg U63759 ( .A(n47367), .B(n39938), .X(n7850) );
  nand_x1_sg U63760 ( .A(n47652), .B(n39940), .X(n8668) );
  nand_x1_sg U63761 ( .A(n47937), .B(n39942), .X(n9488) );
  nand_x1_sg U63762 ( .A(n48222), .B(n39958), .X(n10307) );
  nand_x1_sg U63763 ( .A(n48507), .B(n39961), .X(n11126) );
  nand_x1_sg U63764 ( .A(n48792), .B(n39950), .X(n11945) );
  nand_x1_sg U63765 ( .A(n49079), .B(n39952), .X(n12764) );
  nand_x1_sg U63766 ( .A(n49365), .B(n39954), .X(n13583) );
  nand_x1_sg U63767 ( .A(n49651), .B(n39948), .X(n14402) );
  nand_x1_sg U63768 ( .A(n49937), .B(n39944), .X(n15221) );
  nand_x1_sg U63769 ( .A(n50223), .B(n39946), .X(n16040) );
  nand_x1_sg U63770 ( .A(n50508), .B(n39932), .X(n16859) );
  nand_x1_sg U63771 ( .A(n50797), .B(n39934), .X(n17678) );
  nand_x1_sg U63772 ( .A(n51084), .B(n39936), .X(n18499) );
  nand_x1_sg U63773 ( .A(n6990), .B(n39664), .X(n6989) );
  nand_x1_sg U63774 ( .A(n6992), .B(n6993), .X(n6988) );
  nand_x1_sg U63775 ( .A(n7807), .B(n42358), .X(n7806) );
  nand_x1_sg U63776 ( .A(n7809), .B(n7810), .X(n7805) );
  nand_x1_sg U63777 ( .A(n8625), .B(n42357), .X(n8624) );
  nand_x1_sg U63778 ( .A(n8627), .B(n8628), .X(n8623) );
  nand_x1_sg U63779 ( .A(n9445), .B(n42368), .X(n9444) );
  nand_x1_sg U63780 ( .A(n9447), .B(n9448), .X(n9443) );
  nand_x1_sg U63781 ( .A(n10264), .B(n42367), .X(n10263) );
  nand_x1_sg U63782 ( .A(n10266), .B(n10267), .X(n10262) );
  nand_x1_sg U63783 ( .A(n11083), .B(n42366), .X(n11082) );
  nand_x1_sg U63784 ( .A(n11085), .B(n11086), .X(n11081) );
  nand_x1_sg U63785 ( .A(n11902), .B(n42365), .X(n11901) );
  nand_x1_sg U63786 ( .A(n11904), .B(n11905), .X(n11900) );
  nand_x1_sg U63787 ( .A(n12721), .B(n42364), .X(n12720) );
  nand_x1_sg U63788 ( .A(n12723), .B(n12724), .X(n12719) );
  nand_x1_sg U63789 ( .A(n13540), .B(n42363), .X(n13539) );
  nand_x1_sg U63790 ( .A(n13542), .B(n13543), .X(n13538) );
  nand_x1_sg U63791 ( .A(n14359), .B(n42362), .X(n14358) );
  nand_x1_sg U63792 ( .A(n14361), .B(n14362), .X(n14357) );
  nand_x1_sg U63793 ( .A(n15178), .B(n42361), .X(n15177) );
  nand_x1_sg U63794 ( .A(n15180), .B(n15181), .X(n15176) );
  nand_x1_sg U63795 ( .A(n15997), .B(n42360), .X(n15996) );
  nand_x1_sg U63796 ( .A(n15999), .B(n16000), .X(n15995) );
  nand_x1_sg U63797 ( .A(n16814), .B(n39661), .X(n16813) );
  nand_x1_sg U63798 ( .A(n16816), .B(n16817), .X(n16812) );
  nand_x1_sg U63799 ( .A(n17635), .B(n39543), .X(n17634) );
  nand_x1_sg U63800 ( .A(n17637), .B(n17638), .X(n17633) );
  nand_x1_sg U63801 ( .A(n18456), .B(n42359), .X(n18455) );
  nand_x1_sg U63802 ( .A(n18458), .B(n18459), .X(n18454) );
  nand_x1_sg U63803 ( .A(n39802), .B(n40162), .X(n7537) );
  nand_x1_sg U63804 ( .A(n39799), .B(n40243), .X(n8355) );
  nand_x1_sg U63805 ( .A(n39801), .B(n40249), .X(n9173) );
  nand_x1_sg U63806 ( .A(n39795), .B(n40255), .X(n9993) );
  nand_x1_sg U63807 ( .A(n39797), .B(n40258), .X(n10812) );
  nand_x1_sg U63808 ( .A(n39791), .B(n40262), .X(n11631) );
  nand_x1_sg U63809 ( .A(n39793), .B(n40267), .X(n12450) );
  nand_x1_sg U63810 ( .A(n39787), .B(n40273), .X(n13269) );
  nand_x1_sg U63811 ( .A(n39789), .B(n40277), .X(n14088) );
  nand_x1_sg U63812 ( .A(n39783), .B(n40284), .X(n14907) );
  nand_x1_sg U63813 ( .A(n39785), .B(n40288), .X(n15726) );
  nand_x1_sg U63814 ( .A(n39779), .B(n40292), .X(n16545) );
  nand_x1_sg U63815 ( .A(n39781), .B(n40238), .X(n18183) );
  nand_x1_sg U63816 ( .A(n39777), .B(n40297), .X(n19004) );
  nor_x1_sg U63817 ( .A(n40984), .B(n5753), .X(\L1_0/n3472 ) );
  nor_x1_sg U63818 ( .A(n40985), .B(n5760), .X(\L1_0/n3468 ) );
  nor_x1_sg U63819 ( .A(n40984), .B(n5749), .X(\L1_0/n3456 ) );
  nor_x1_sg U63820 ( .A(n41944), .B(n5755), .X(n5126) );
  nor_x1_sg U63821 ( .A(n40982), .B(n5743), .X(n5129) );
  nor_x1_sg U63822 ( .A(n40983), .B(n5762), .X(\L1_0/n3408 ) );
  nor_x1_sg U63823 ( .A(n38939), .B(n5744), .X(n5128) );
  nor_x1_sg U63824 ( .A(n50556), .B(n5745), .X(n5744) );
  inv_x1_sg U63825 ( .A(n5747), .X(n50556) );
  nand_x1_sg U63826 ( .A(n41464), .B(n39482), .X(n5745) );
  inv_x1_sg U63827 ( .A(n8053), .X(n47245) );
  inv_x1_sg U63828 ( .A(n8871), .X(n47530) );
  inv_x1_sg U63829 ( .A(n9691), .X(n47815) );
  inv_x1_sg U63830 ( .A(n10510), .X(n48100) );
  inv_x1_sg U63831 ( .A(n11329), .X(n48385) );
  inv_x1_sg U63832 ( .A(n12148), .X(n48670) );
  inv_x1_sg U63833 ( .A(n12967), .X(n48956) );
  inv_x1_sg U63834 ( .A(n13786), .X(n49243) );
  inv_x1_sg U63835 ( .A(n14605), .X(n49529) );
  inv_x1_sg U63836 ( .A(n15424), .X(n49815) );
  inv_x1_sg U63837 ( .A(n16243), .X(n50101) );
  inv_x1_sg U63838 ( .A(n17881), .X(n50675) );
  inv_x1_sg U63839 ( .A(n18702), .X(n50962) );
  inv_x1_sg U63840 ( .A(n7234), .X(n46954) );
  inv_x1_sg U63841 ( .A(n17059), .X(n50386) );
  nor_x1_sg U63842 ( .A(n6017), .B(n6018), .X(n6016) );
  nor_x1_sg U63843 ( .A(n6021), .B(n6022), .X(n6015) );
  nor_x1_sg U63844 ( .A(n6020), .B(n41040), .X(n6017) );
  nor_x1_sg U63845 ( .A(n6205), .B(n6206), .X(n6204) );
  nor_x1_sg U63846 ( .A(n6208), .B(n6209), .X(n6203) );
  nor_x1_sg U63847 ( .A(n41538), .B(n38927), .X(n6206) );
  nor_x1_sg U63848 ( .A(n6005), .B(n6006), .X(n5999) );
  nor_x1_sg U63849 ( .A(n6001), .B(n6002), .X(n6000) );
  nor_x1_sg U63850 ( .A(n42023), .B(n41013), .X(n6006) );
  nor_x1_sg U63851 ( .A(n6066), .B(n6067), .X(n6065) );
  nor_x1_sg U63852 ( .A(n6069), .B(n6070), .X(n6064) );
  nor_x1_sg U63853 ( .A(n41953), .B(n41038), .X(n6066) );
  nor_x1_sg U63854 ( .A(n6114), .B(n6115), .X(n6113) );
  nor_x1_sg U63855 ( .A(n6116), .B(n6117), .X(n6112) );
  nor_x1_sg U63856 ( .A(n42226), .B(n41005), .X(n6115) );
  nor_x1_sg U63857 ( .A(n6053), .B(n6054), .X(n6047) );
  nor_x1_sg U63858 ( .A(n6049), .B(n6050), .X(n6048) );
  nor_x1_sg U63859 ( .A(n41525), .B(n41035), .X(n6053) );
  nor_x1_sg U63860 ( .A(n6103), .B(n6104), .X(n6097) );
  nor_x1_sg U63861 ( .A(n6099), .B(n6100), .X(n6098) );
  nor_x1_sg U63862 ( .A(n46506), .B(n41014), .X(n6104) );
  nor_x1_sg U63863 ( .A(n6148), .B(n6149), .X(n6143) );
  nor_x1_sg U63864 ( .A(n6145), .B(n6146), .X(n6144) );
  nor_x1_sg U63865 ( .A(n46469), .B(n41013), .X(n6149) );
  nor_x1_sg U63866 ( .A(n6163), .B(n6164), .X(n6157) );
  nor_x1_sg U63867 ( .A(n6159), .B(n6160), .X(n6158) );
  nor_x1_sg U63868 ( .A(n41537), .B(n41028), .X(n6164) );
  nor_x1_sg U63869 ( .A(n6194), .B(n6195), .X(n6189) );
  nor_x1_sg U63870 ( .A(n6191), .B(n6192), .X(n6190) );
  nor_x1_sg U63871 ( .A(n46422), .B(n41016), .X(n6195) );
  nor_x1_sg U63872 ( .A(n6241), .B(n6242), .X(n6235) );
  nor_x1_sg U63873 ( .A(n6237), .B(n6238), .X(n6236) );
  nor_x1_sg U63874 ( .A(n46374), .B(n38914), .X(n6242) );
  nor_x1_sg U63875 ( .A(n6256), .B(n6257), .X(n6250) );
  nor_x1_sg U63876 ( .A(n6252), .B(n6253), .X(n6251) );
  nor_x1_sg U63877 ( .A(n46336), .B(n41030), .X(n6257) );
  nor_x1_sg U63878 ( .A(n6286), .B(n6287), .X(n6280) );
  nor_x1_sg U63879 ( .A(n6282), .B(n6283), .X(n6281) );
  nor_x1_sg U63880 ( .A(n46333), .B(n38914), .X(n6287) );
  nor_x1_sg U63881 ( .A(n6301), .B(n6302), .X(n6295) );
  nor_x1_sg U63882 ( .A(n6297), .B(n6298), .X(n6296) );
  nor_x1_sg U63883 ( .A(n46290), .B(n38933), .X(n6302) );
  nor_x1_sg U63884 ( .A(n6330), .B(n6331), .X(n6324) );
  nor_x1_sg U63885 ( .A(n6326), .B(n6327), .X(n6325) );
  nor_x1_sg U63886 ( .A(n46287), .B(n41015), .X(n6331) );
  nor_x1_sg U63887 ( .A(n6345), .B(n6346), .X(n6339) );
  nor_x1_sg U63888 ( .A(n6341), .B(n6342), .X(n6340) );
  nor_x1_sg U63889 ( .A(n46245), .B(n41029), .X(n6346) );
  nor_x1_sg U63890 ( .A(n6375), .B(n6376), .X(n6369) );
  nor_x1_sg U63891 ( .A(n6371), .B(n6372), .X(n6370) );
  nor_x1_sg U63892 ( .A(n46242), .B(n41014), .X(n6376) );
  nor_x1_sg U63893 ( .A(n6390), .B(n6391), .X(n6384) );
  nor_x1_sg U63894 ( .A(n6386), .B(n6387), .X(n6385) );
  nor_x1_sg U63895 ( .A(n46199), .B(n41028), .X(n6391) );
  nor_x1_sg U63896 ( .A(n6419), .B(n6420), .X(n6413) );
  nor_x1_sg U63897 ( .A(n6415), .B(n6416), .X(n6414) );
  nor_x1_sg U63898 ( .A(n46196), .B(n41013), .X(n6420) );
  nor_x1_sg U63899 ( .A(n6434), .B(n6435), .X(n6428) );
  nor_x1_sg U63900 ( .A(n6430), .B(n6431), .X(n6429) );
  nor_x1_sg U63901 ( .A(n46154), .B(n41568), .X(n6435) );
  nor_x1_sg U63902 ( .A(n6464), .B(n6465), .X(n6458) );
  nor_x1_sg U63903 ( .A(n6460), .B(n6461), .X(n6459) );
  nor_x1_sg U63904 ( .A(n46151), .B(n41015), .X(n6465) );
  nor_x1_sg U63905 ( .A(n6479), .B(n6480), .X(n6473) );
  nor_x1_sg U63906 ( .A(n6475), .B(n6476), .X(n6474) );
  nor_x1_sg U63907 ( .A(n46108), .B(n41029), .X(n6480) );
  nor_x1_sg U63908 ( .A(n6508), .B(n6509), .X(n6502) );
  nor_x1_sg U63909 ( .A(n6504), .B(n6505), .X(n6503) );
  nor_x1_sg U63910 ( .A(n46105), .B(n41016), .X(n6509) );
  nor_x1_sg U63911 ( .A(n6523), .B(n6524), .X(n6517) );
  nor_x1_sg U63912 ( .A(n6519), .B(n6520), .X(n6518) );
  nor_x1_sg U63913 ( .A(n46063), .B(n41029), .X(n6524) );
  nor_x1_sg U63914 ( .A(n6553), .B(n6554), .X(n6547) );
  nor_x1_sg U63915 ( .A(n6549), .B(n6550), .X(n6548) );
  nor_x1_sg U63916 ( .A(n46060), .B(n41571), .X(n6554) );
  nor_x1_sg U63917 ( .A(n6568), .B(n6569), .X(n6562) );
  nor_x1_sg U63918 ( .A(n6564), .B(n6565), .X(n6563) );
  nor_x1_sg U63919 ( .A(n46017), .B(n41028), .X(n6569) );
  nor_x1_sg U63920 ( .A(n6597), .B(n6598), .X(n6591) );
  nor_x1_sg U63921 ( .A(n6593), .B(n6594), .X(n6592) );
  nor_x1_sg U63922 ( .A(n46014), .B(n41015), .X(n6598) );
  nor_x1_sg U63923 ( .A(n6612), .B(n6613), .X(n6606) );
  nor_x1_sg U63924 ( .A(n6608), .B(n6609), .X(n6607) );
  nor_x1_sg U63925 ( .A(n45972), .B(n41030), .X(n6613) );
  nor_x1_sg U63926 ( .A(n6642), .B(n6643), .X(n6636) );
  nor_x1_sg U63927 ( .A(n6638), .B(n6639), .X(n6637) );
  nor_x1_sg U63928 ( .A(n45969), .B(n41016), .X(n6643) );
  nor_x1_sg U63929 ( .A(n6657), .B(n6658), .X(n6651) );
  nor_x1_sg U63930 ( .A(n6653), .B(n6654), .X(n6652) );
  nor_x1_sg U63931 ( .A(n42200), .B(n41572), .X(n6657) );
  nor_x1_sg U63932 ( .A(n6689), .B(n6690), .X(n6683) );
  nor_x1_sg U63933 ( .A(n6685), .B(n6686), .X(n6684) );
  nor_x1_sg U63934 ( .A(n42199), .B(n41036), .X(n6689) );
  nor_x1_sg U63935 ( .A(n6703), .B(n6704), .X(n6699) );
  nor_x1_sg U63936 ( .A(n6701), .B(n6702), .X(n6700) );
  nor_x1_sg U63937 ( .A(n41528), .B(n41009), .X(n6703) );
  nor_x1_sg U63938 ( .A(n6730), .B(n6731), .X(n6726) );
  nor_x1_sg U63939 ( .A(n6728), .B(n6729), .X(n6727) );
  nor_x1_sg U63940 ( .A(n41529), .B(n41033), .X(n6730) );
  nand_x1_sg U63941 ( .A(n40509), .B(n39731), .X(n22939) );
  nand_x1_sg U63942 ( .A(n39221), .B(n41578), .X(n22953) );
  nand_x1_sg U63943 ( .A(n40504), .B(n39734), .X(n23216) );
  nand_x1_sg U63944 ( .A(n40503), .B(n41577), .X(n23230) );
  nand_x1_sg U63945 ( .A(n40500), .B(n39737), .X(n23496) );
  nand_x1_sg U63946 ( .A(n39225), .B(n41576), .X(n23510) );
  nand_x1_sg U63947 ( .A(n40496), .B(n39740), .X(n23775) );
  nand_x1_sg U63948 ( .A(n40497), .B(n41575), .X(n23789) );
  nand_x1_sg U63949 ( .A(n41171), .B(n39743), .X(n24054) );
  nand_x1_sg U63950 ( .A(n40492), .B(n41582), .X(n24068) );
  nand_x1_sg U63951 ( .A(n40488), .B(n39746), .X(n24333) );
  nand_x1_sg U63952 ( .A(n40489), .B(n41581), .X(n24347) );
  nand_x1_sg U63953 ( .A(n40485), .B(n39749), .X(n24612) );
  nand_x1_sg U63954 ( .A(n40483), .B(n41580), .X(n24626) );
  nand_x1_sg U63955 ( .A(n40480), .B(n39752), .X(n24890) );
  nand_x1_sg U63956 ( .A(n40480), .B(n41579), .X(n24904) );
  nand_x1_sg U63957 ( .A(n40476), .B(n39755), .X(n25169) );
  nand_x1_sg U63958 ( .A(n39237), .B(n41586), .X(n25183) );
  nand_x1_sg U63959 ( .A(n40472), .B(n39758), .X(n25448) );
  nand_x1_sg U63960 ( .A(n40473), .B(n41585), .X(n25462) );
  nand_x1_sg U63961 ( .A(n39241), .B(n39761), .X(n25727) );
  nand_x1_sg U63962 ( .A(n41141), .B(n41584), .X(n25741) );
  nand_x1_sg U63963 ( .A(n39243), .B(n39764), .X(n26279) );
  nand_x1_sg U63964 ( .A(n40463), .B(n41587), .X(n26295) );
  nand_x1_sg U63965 ( .A(n40460), .B(n39767), .X(n26564) );
  nand_x1_sg U63966 ( .A(n39245), .B(n41583), .X(n26578) );
  nor_x1_sg U63967 ( .A(n23175), .B(n39440), .X(\L1_0/n4247 ) );
  nor_x1_sg U63968 ( .A(n23182), .B(n41378), .X(\L1_0/n4243 ) );
  nor_x1_sg U63969 ( .A(n23196), .B(n39439), .X(\L1_0/n4235 ) );
  nor_x1_sg U63970 ( .A(n23210), .B(n41375), .X(\L1_0/n4227 ) );
  nor_x1_sg U63971 ( .A(n23224), .B(n41378), .X(\L1_0/n4219 ) );
  nor_x1_sg U63972 ( .A(n23455), .B(n41347), .X(\L1_0/n4167 ) );
  nor_x1_sg U63973 ( .A(n23462), .B(n39914), .X(\L1_0/n4163 ) );
  nor_x1_sg U63974 ( .A(n23476), .B(n38961), .X(\L1_0/n4155 ) );
  nor_x1_sg U63975 ( .A(n23490), .B(n41348), .X(\L1_0/n4147 ) );
  nor_x1_sg U63976 ( .A(n23504), .B(n38961), .X(\L1_0/n4139 ) );
  nor_x1_sg U63977 ( .A(n23530), .B(n39457), .X(\L1_0/n4123 ) );
  nor_x1_sg U63978 ( .A(n23734), .B(n41342), .X(\L1_0/n4087 ) );
  nor_x1_sg U63979 ( .A(n23741), .B(n41343), .X(\L1_0/n4083 ) );
  nor_x1_sg U63980 ( .A(n23755), .B(n41340), .X(\L1_0/n4075 ) );
  nor_x1_sg U63981 ( .A(n23769), .B(n38958), .X(\L1_0/n4067 ) );
  nor_x1_sg U63982 ( .A(n23783), .B(n39460), .X(\L1_0/n4059 ) );
  nor_x1_sg U63983 ( .A(n23809), .B(n41343), .X(\L1_0/n4043 ) );
  nor_x1_sg U63984 ( .A(n24013), .B(n39449), .X(\L1_0/n4007 ) );
  nor_x1_sg U63985 ( .A(n24020), .B(n41363), .X(\L1_0/n4003 ) );
  nor_x1_sg U63986 ( .A(n24034), .B(n41361), .X(\L1_0/n3995 ) );
  nor_x1_sg U63987 ( .A(n24048), .B(n41360), .X(\L1_0/n3987 ) );
  nor_x1_sg U63988 ( .A(n24062), .B(n41363), .X(\L1_0/n3979 ) );
  nor_x1_sg U63989 ( .A(n24088), .B(n39909), .X(\L1_0/n3963 ) );
  nor_x1_sg U63990 ( .A(n24292), .B(n38967), .X(\L1_0/n3927 ) );
  nor_x1_sg U63991 ( .A(n24299), .B(n41356), .X(\L1_0/n3923 ) );
  nor_x1_sg U63992 ( .A(n24313), .B(n38967), .X(\L1_0/n3915 ) );
  nor_x1_sg U63993 ( .A(n24327), .B(n41358), .X(\L1_0/n3907 ) );
  nor_x1_sg U63994 ( .A(n24341), .B(n39451), .X(\L1_0/n3899 ) );
  nor_x1_sg U63995 ( .A(n24367), .B(n38966), .X(\L1_0/n3883 ) );
  nor_x1_sg U63996 ( .A(n24571), .B(n39464), .X(\L1_0/n3847 ) );
  nor_x1_sg U63997 ( .A(n24578), .B(n39464), .X(\L1_0/n3843 ) );
  nor_x1_sg U63998 ( .A(n24592), .B(n39463), .X(\L1_0/n3835 ) );
  nor_x1_sg U63999 ( .A(n24606), .B(n39919), .X(\L1_0/n3827 ) );
  nor_x1_sg U64000 ( .A(n24620), .B(n41338), .X(\L1_0/n3819 ) );
  nor_x1_sg U64001 ( .A(n24646), .B(n39918), .X(\L1_0/n3803 ) );
  nor_x1_sg U64002 ( .A(n24849), .B(n39467), .X(\L1_0/n3767 ) );
  nor_x1_sg U64003 ( .A(n24856), .B(n41330), .X(\L1_0/n3763 ) );
  nor_x1_sg U64004 ( .A(n24870), .B(n41333), .X(\L1_0/n3755 ) );
  nor_x1_sg U64005 ( .A(n24884), .B(n38951), .X(\L1_0/n3747 ) );
  nor_x1_sg U64006 ( .A(n24898), .B(n39467), .X(\L1_0/n3739 ) );
  nor_x1_sg U64007 ( .A(n24924), .B(n41330), .X(\L1_0/n3723 ) );
  nor_x1_sg U64008 ( .A(n25128), .B(n39922), .X(\L1_0/n3687 ) );
  nor_x1_sg U64009 ( .A(n25135), .B(n39922), .X(\L1_0/n3683 ) );
  nor_x1_sg U64010 ( .A(n25149), .B(n41327), .X(\L1_0/n3675 ) );
  nor_x1_sg U64011 ( .A(n25163), .B(n41325), .X(\L1_0/n3667 ) );
  nor_x1_sg U64012 ( .A(n25177), .B(n38949), .X(\L1_0/n3659 ) );
  nor_x1_sg U64013 ( .A(n25203), .B(n41325), .X(\L1_0/n3643 ) );
  nor_x1_sg U64014 ( .A(n25407), .B(n39904), .X(\L1_0/n3607 ) );
  nor_x1_sg U64015 ( .A(n25414), .B(n38975), .X(\L1_0/n3603 ) );
  nor_x1_sg U64016 ( .A(n25428), .B(n41372), .X(\L1_0/n3595 ) );
  nor_x1_sg U64017 ( .A(n25442), .B(n41373), .X(\L1_0/n3587 ) );
  nor_x1_sg U64018 ( .A(n25456), .B(n38976), .X(\L1_0/n3579 ) );
  nor_x1_sg U64019 ( .A(n25482), .B(n41373), .X(\L1_0/n3563 ) );
  nor_x1_sg U64020 ( .A(n25686), .B(n40035), .X(\L1_0/n3527 ) );
  nor_x1_sg U64021 ( .A(n25693), .B(n39901), .X(\L1_0/n3523 ) );
  nor_x1_sg U64022 ( .A(n25707), .B(n40033), .X(\L1_0/n3515 ) );
  nor_x1_sg U64023 ( .A(n25721), .B(n41381), .X(\L1_0/n3507 ) );
  nor_x1_sg U64024 ( .A(n25735), .B(n41380), .X(\L1_0/n3499 ) );
  nor_x1_sg U64025 ( .A(n25761), .B(n41382), .X(\L1_0/n3483 ) );
  nor_x1_sg U64026 ( .A(n26523), .B(n39913), .X(\L1_0/n3287 ) );
  nor_x1_sg U64027 ( .A(n26530), .B(n38963), .X(\L1_0/n3283 ) );
  nor_x1_sg U64028 ( .A(n26544), .B(n41351), .X(\L1_0/n3275 ) );
  nor_x1_sg U64029 ( .A(n26558), .B(n39912), .X(\L1_0/n3267 ) );
  nor_x1_sg U64030 ( .A(n26572), .B(n39455), .X(\L1_0/n3259 ) );
  nor_x1_sg U64031 ( .A(n26598), .B(n38963), .X(\L1_0/n3243 ) );
  nor_x1_sg U64032 ( .A(n23250), .B(n39903), .X(\L1_0/n4203 ) );
  nand_x1_sg U64033 ( .A(n41110), .B(n44984), .X(n22541) );
  nand_x1_sg U64034 ( .A(n41087), .B(n44993), .X(n22540) );
  nor_x1_sg U64035 ( .A(n7652), .B(n40973), .X(\L2_0/n3436 ) );
  nor_x1_sg U64036 ( .A(n9290), .B(n40969), .X(\L2_0/n3276 ) );
  nor_x1_sg U64037 ( .A(n10109), .B(n40961), .X(\L2_0/n3196 ) );
  nor_x1_sg U64038 ( .A(n10928), .B(n40929), .X(\L2_0/n3116 ) );
  nor_x1_sg U64039 ( .A(n11747), .B(n40933), .X(\L2_0/n3036 ) );
  nor_x1_sg U64040 ( .A(n12566), .B(n40937), .X(\L2_0/n2956 ) );
  nor_x1_sg U64041 ( .A(n13385), .B(n40941), .X(\L2_0/n2876 ) );
  nor_x1_sg U64042 ( .A(n14204), .B(n40945), .X(\L2_0/n2796 ) );
  nor_x1_sg U64043 ( .A(n15023), .B(n40949), .X(\L2_0/n2716 ) );
  nor_x1_sg U64044 ( .A(n15842), .B(n40953), .X(\L2_0/n2636 ) );
  nor_x1_sg U64045 ( .A(n18301), .B(n40957), .X(\L2_0/n2396 ) );
  nor_x1_sg U64046 ( .A(n7744), .B(n40974), .X(\L2_0/n3376 ) );
  nor_x1_sg U64047 ( .A(n9382), .B(n40970), .X(\L2_0/n3216 ) );
  nor_x1_sg U64048 ( .A(n10201), .B(n40962), .X(\L2_0/n3136 ) );
  nor_x1_sg U64049 ( .A(n11020), .B(n40930), .X(\L2_0/n3056 ) );
  nor_x1_sg U64050 ( .A(n11839), .B(n40934), .X(\L2_0/n2976 ) );
  nor_x1_sg U64051 ( .A(n12658), .B(n40938), .X(\L2_0/n2896 ) );
  nor_x1_sg U64052 ( .A(n13477), .B(n40942), .X(\L2_0/n2816 ) );
  nor_x1_sg U64053 ( .A(n14296), .B(n40946), .X(\L2_0/n2736 ) );
  nor_x1_sg U64054 ( .A(n15115), .B(n40950), .X(\L2_0/n2656 ) );
  nor_x1_sg U64055 ( .A(n15934), .B(n40954), .X(\L2_0/n2576 ) );
  nor_x1_sg U64056 ( .A(n18393), .B(n40958), .X(\L2_0/n2336 ) );
  nor_x1_sg U64057 ( .A(n7666), .B(n38905), .X(\L2_0/n3428 ) );
  nor_x1_sg U64058 ( .A(n7672), .B(n38905), .X(\L2_0/n3424 ) );
  nor_x1_sg U64059 ( .A(n7690), .B(n40975), .X(\L2_0/n3412 ) );
  nor_x1_sg U64060 ( .A(n7702), .B(n40973), .X(\L2_0/n3404 ) );
  nor_x1_sg U64061 ( .A(n7708), .B(n7638), .X(\L2_0/n3400 ) );
  nor_x1_sg U64062 ( .A(n7714), .B(n40975), .X(\L2_0/n3396 ) );
  nor_x1_sg U64063 ( .A(n7720), .B(n40974), .X(\L2_0/n3392 ) );
  nor_x1_sg U64064 ( .A(n7726), .B(n40973), .X(\L2_0/n3388 ) );
  nor_x1_sg U64065 ( .A(n7732), .B(n40974), .X(\L2_0/n3384 ) );
  nor_x1_sg U64066 ( .A(n7738), .B(n38905), .X(\L2_0/n3380 ) );
  nor_x1_sg U64067 ( .A(n9304), .B(n40969), .X(\L2_0/n3268 ) );
  nor_x1_sg U64068 ( .A(n9310), .B(n40971), .X(\L2_0/n3264 ) );
  nor_x1_sg U64069 ( .A(n9328), .B(n40969), .X(\L2_0/n3252 ) );
  nor_x1_sg U64070 ( .A(n9340), .B(n40971), .X(\L2_0/n3244 ) );
  nor_x1_sg U64071 ( .A(n9346), .B(n40971), .X(\L2_0/n3240 ) );
  nor_x1_sg U64072 ( .A(n9352), .B(n38904), .X(\L2_0/n3236 ) );
  nor_x1_sg U64073 ( .A(n9358), .B(n40970), .X(\L2_0/n3232 ) );
  nor_x1_sg U64074 ( .A(n9364), .B(n9276), .X(\L2_0/n3228 ) );
  nor_x1_sg U64075 ( .A(n9370), .B(n40970), .X(\L2_0/n3224 ) );
  nor_x1_sg U64076 ( .A(n9376), .B(n9276), .X(\L2_0/n3220 ) );
  nor_x1_sg U64077 ( .A(n10123), .B(n40962), .X(\L2_0/n3188 ) );
  nor_x1_sg U64078 ( .A(n10129), .B(n40963), .X(\L2_0/n3184 ) );
  nor_x1_sg U64079 ( .A(n10147), .B(n38902), .X(\L2_0/n3172 ) );
  nor_x1_sg U64080 ( .A(n10159), .B(n40962), .X(\L2_0/n3164 ) );
  nor_x1_sg U64081 ( .A(n10165), .B(n38902), .X(\L2_0/n3160 ) );
  nor_x1_sg U64082 ( .A(n10171), .B(n40963), .X(\L2_0/n3156 ) );
  nor_x1_sg U64083 ( .A(n10177), .B(n10095), .X(\L2_0/n3152 ) );
  nor_x1_sg U64084 ( .A(n10183), .B(n40963), .X(\L2_0/n3148 ) );
  nor_x1_sg U64085 ( .A(n10189), .B(n10095), .X(\L2_0/n3144 ) );
  nor_x1_sg U64086 ( .A(n10195), .B(n38902), .X(\L2_0/n3140 ) );
  nor_x1_sg U64087 ( .A(n10942), .B(n38894), .X(\L2_0/n3108 ) );
  nor_x1_sg U64088 ( .A(n10948), .B(n40931), .X(\L2_0/n3104 ) );
  nor_x1_sg U64089 ( .A(n10966), .B(n40929), .X(\L2_0/n3092 ) );
  nor_x1_sg U64090 ( .A(n10978), .B(n40930), .X(\L2_0/n3084 ) );
  nor_x1_sg U64091 ( .A(n10984), .B(n38894), .X(\L2_0/n3080 ) );
  nor_x1_sg U64092 ( .A(n10990), .B(n40930), .X(\L2_0/n3076 ) );
  nor_x1_sg U64093 ( .A(n10996), .B(n10914), .X(\L2_0/n3072 ) );
  nor_x1_sg U64094 ( .A(n11002), .B(n40929), .X(\L2_0/n3068 ) );
  nor_x1_sg U64095 ( .A(n11008), .B(n10914), .X(\L2_0/n3064 ) );
  nor_x1_sg U64096 ( .A(n11014), .B(n40931), .X(\L2_0/n3060 ) );
  nor_x1_sg U64097 ( .A(n11761), .B(n38895), .X(\L2_0/n3028 ) );
  nor_x1_sg U64098 ( .A(n11767), .B(n38895), .X(\L2_0/n3024 ) );
  nor_x1_sg U64099 ( .A(n11785), .B(n11733), .X(\L2_0/n3012 ) );
  nor_x1_sg U64100 ( .A(n11797), .B(n40934), .X(\L2_0/n3004 ) );
  nor_x1_sg U64101 ( .A(n11803), .B(n40934), .X(\L2_0/n3000 ) );
  nor_x1_sg U64102 ( .A(n11809), .B(n40935), .X(\L2_0/n2996 ) );
  nor_x1_sg U64103 ( .A(n11815), .B(n40934), .X(\L2_0/n2992 ) );
  nor_x1_sg U64104 ( .A(n11821), .B(n11733), .X(\L2_0/n2988 ) );
  nor_x1_sg U64105 ( .A(n11827), .B(n40935), .X(\L2_0/n2984 ) );
  nor_x1_sg U64106 ( .A(n11833), .B(n11733), .X(\L2_0/n2980 ) );
  nor_x1_sg U64107 ( .A(n12580), .B(n12552), .X(\L2_0/n2948 ) );
  nor_x1_sg U64108 ( .A(n12586), .B(n40939), .X(\L2_0/n2944 ) );
  nor_x1_sg U64109 ( .A(n12604), .B(n40937), .X(\L2_0/n2932 ) );
  nor_x1_sg U64110 ( .A(n12616), .B(n12552), .X(\L2_0/n2924 ) );
  nor_x1_sg U64111 ( .A(n12622), .B(n38896), .X(\L2_0/n2920 ) );
  nor_x1_sg U64112 ( .A(n12628), .B(n12552), .X(\L2_0/n2916 ) );
  nor_x1_sg U64113 ( .A(n12634), .B(n38896), .X(\L2_0/n2912 ) );
  nor_x1_sg U64114 ( .A(n12640), .B(n40937), .X(\L2_0/n2908 ) );
  nor_x1_sg U64115 ( .A(n12646), .B(n40938), .X(\L2_0/n2904 ) );
  nor_x1_sg U64116 ( .A(n12652), .B(n40939), .X(\L2_0/n2900 ) );
  nor_x1_sg U64117 ( .A(n13399), .B(n40941), .X(\L2_0/n2868 ) );
  nor_x1_sg U64118 ( .A(n13405), .B(n38897), .X(\L2_0/n2864 ) );
  nor_x1_sg U64119 ( .A(n13423), .B(n38897), .X(\L2_0/n2852 ) );
  nor_x1_sg U64120 ( .A(n13435), .B(n13371), .X(\L2_0/n2844 ) );
  nor_x1_sg U64121 ( .A(n13441), .B(n38897), .X(\L2_0/n2840 ) );
  nor_x1_sg U64122 ( .A(n13447), .B(n40942), .X(\L2_0/n2836 ) );
  nor_x1_sg U64123 ( .A(n13453), .B(n40942), .X(\L2_0/n2832 ) );
  nor_x1_sg U64124 ( .A(n13459), .B(n40943), .X(\L2_0/n2828 ) );
  nor_x1_sg U64125 ( .A(n13465), .B(n40943), .X(\L2_0/n2824 ) );
  nor_x1_sg U64126 ( .A(n13471), .B(n13371), .X(\L2_0/n2820 ) );
  nor_x1_sg U64127 ( .A(n14218), .B(n14190), .X(\L2_0/n2788 ) );
  nor_x1_sg U64128 ( .A(n14224), .B(n40947), .X(\L2_0/n2784 ) );
  nor_x1_sg U64129 ( .A(n14242), .B(n40945), .X(\L2_0/n2772 ) );
  nor_x1_sg U64130 ( .A(n14254), .B(n40946), .X(\L2_0/n2764 ) );
  nor_x1_sg U64131 ( .A(n14260), .B(n38898), .X(\L2_0/n2760 ) );
  nor_x1_sg U64132 ( .A(n14266), .B(n40946), .X(\L2_0/n2756 ) );
  nor_x1_sg U64133 ( .A(n14272), .B(n14190), .X(\L2_0/n2752 ) );
  nor_x1_sg U64134 ( .A(n14278), .B(n40945), .X(\L2_0/n2748 ) );
  nor_x1_sg U64135 ( .A(n14284), .B(n14190), .X(\L2_0/n2744 ) );
  nor_x1_sg U64136 ( .A(n14290), .B(n40947), .X(\L2_0/n2740 ) );
  nor_x1_sg U64137 ( .A(n15037), .B(n38899), .X(\L2_0/n2708 ) );
  nor_x1_sg U64138 ( .A(n15043), .B(n38899), .X(\L2_0/n2704 ) );
  nor_x1_sg U64139 ( .A(n15061), .B(n15009), .X(\L2_0/n2692 ) );
  nor_x1_sg U64140 ( .A(n15073), .B(n40950), .X(\L2_0/n2684 ) );
  nor_x1_sg U64141 ( .A(n15079), .B(n40950), .X(\L2_0/n2680 ) );
  nor_x1_sg U64142 ( .A(n15085), .B(n40951), .X(\L2_0/n2676 ) );
  nor_x1_sg U64143 ( .A(n15091), .B(n40950), .X(\L2_0/n2672 ) );
  nor_x1_sg U64144 ( .A(n15097), .B(n15009), .X(\L2_0/n2668 ) );
  nor_x1_sg U64145 ( .A(n15103), .B(n40951), .X(\L2_0/n2664 ) );
  nor_x1_sg U64146 ( .A(n15109), .B(n15009), .X(\L2_0/n2660 ) );
  nor_x1_sg U64147 ( .A(n15856), .B(n38900), .X(\L2_0/n2628 ) );
  nor_x1_sg U64148 ( .A(n15862), .B(n40955), .X(\L2_0/n2624 ) );
  nor_x1_sg U64149 ( .A(n15880), .B(n40953), .X(\L2_0/n2612 ) );
  nor_x1_sg U64150 ( .A(n15892), .B(n40954), .X(\L2_0/n2604 ) );
  nor_x1_sg U64151 ( .A(n15898), .B(n38900), .X(\L2_0/n2600 ) );
  nor_x1_sg U64152 ( .A(n15904), .B(n40954), .X(\L2_0/n2596 ) );
  nor_x1_sg U64153 ( .A(n15910), .B(n15828), .X(\L2_0/n2592 ) );
  nor_x1_sg U64154 ( .A(n15916), .B(n40953), .X(\L2_0/n2588 ) );
  nor_x1_sg U64155 ( .A(n15922), .B(n15828), .X(\L2_0/n2584 ) );
  nor_x1_sg U64156 ( .A(n15928), .B(n40955), .X(\L2_0/n2580 ) );
  nor_x1_sg U64157 ( .A(n18315), .B(n38901), .X(\L2_0/n2388 ) );
  nor_x1_sg U64158 ( .A(n18321), .B(n38901), .X(\L2_0/n2384 ) );
  nor_x1_sg U64159 ( .A(n18339), .B(n18287), .X(\L2_0/n2372 ) );
  nor_x1_sg U64160 ( .A(n18351), .B(n40958), .X(\L2_0/n2364 ) );
  nor_x1_sg U64161 ( .A(n18357), .B(n40958), .X(\L2_0/n2360 ) );
  nor_x1_sg U64162 ( .A(n18363), .B(n40959), .X(\L2_0/n2356 ) );
  nor_x1_sg U64163 ( .A(n18369), .B(n40958), .X(\L2_0/n2352 ) );
  nor_x1_sg U64164 ( .A(n18375), .B(n18287), .X(\L2_0/n2348 ) );
  nor_x1_sg U64165 ( .A(n18381), .B(n40959), .X(\L2_0/n2344 ) );
  nor_x1_sg U64166 ( .A(n18387), .B(n18287), .X(\L2_0/n2340 ) );
  nand_x1_sg U64167 ( .A(n40909), .B(n17481), .X(\L2_0/n2475 ) );
  nand_x1_sg U64168 ( .A(n17480), .B(n39253), .X(n17481) );
  nand_x1_sg U64169 ( .A(n38887), .B(n17488), .X(\L2_0/n2471 ) );
  nand_x1_sg U64170 ( .A(n41117), .B(n17487), .X(n17488) );
  nand_x1_sg U64171 ( .A(n40908), .B(n17495), .X(\L2_0/n2467 ) );
  nand_x1_sg U64172 ( .A(n17494), .B(n41119), .X(n17495) );
  nand_x1_sg U64173 ( .A(n40907), .B(n17501), .X(\L2_0/n2463 ) );
  nand_x1_sg U64174 ( .A(n17500), .B(n41118), .X(n17501) );
  nand_x1_sg U64175 ( .A(n40908), .B(n17507), .X(\L2_0/n2459 ) );
  nand_x1_sg U64176 ( .A(n41120), .B(n17506), .X(n17507) );
  nand_x1_sg U64177 ( .A(n40906), .B(n17513), .X(\L2_0/n2455 ) );
  nand_x1_sg U64178 ( .A(n41118), .B(n17512), .X(n17513) );
  nand_x1_sg U64179 ( .A(n40908), .B(n17519), .X(\L2_0/n2451 ) );
  nand_x1_sg U64180 ( .A(n17518), .B(n41117), .X(n17519) );
  nand_x1_sg U64181 ( .A(n40906), .B(n17525), .X(\L2_0/n2447 ) );
  nand_x1_sg U64182 ( .A(n42328), .B(n17524), .X(n17525) );
  nand_x1_sg U64183 ( .A(n38887), .B(n17531), .X(\L2_0/n2443 ) );
  nand_x1_sg U64184 ( .A(n17530), .B(n41120), .X(n17531) );
  nand_x1_sg U64185 ( .A(n40909), .B(n17537), .X(\L2_0/n2439 ) );
  nand_x1_sg U64186 ( .A(n17536), .B(n39253), .X(n17537) );
  nand_x1_sg U64187 ( .A(n40909), .B(n17543), .X(\L2_0/n2435 ) );
  nand_x1_sg U64188 ( .A(n17542), .B(n41119), .X(n17543) );
  nand_x1_sg U64189 ( .A(n38887), .B(n17549), .X(\L2_0/n2431 ) );
  nand_x1_sg U64190 ( .A(n17548), .B(n39253), .X(n17549) );
  nand_x1_sg U64191 ( .A(n40909), .B(n17555), .X(\L2_0/n2427 ) );
  nand_x1_sg U64192 ( .A(n17554), .B(n39253), .X(n17555) );
  nand_x1_sg U64193 ( .A(n40907), .B(n17561), .X(\L2_0/n2423 ) );
  nand_x1_sg U64194 ( .A(n17560), .B(n41120), .X(n17561) );
  nand_x1_sg U64195 ( .A(n40906), .B(n17567), .X(\L2_0/n2419 ) );
  nand_x1_sg U64196 ( .A(n17566), .B(n41120), .X(n17567) );
  nand_x1_sg U64197 ( .A(n40907), .B(n17573), .X(\L2_0/n2415 ) );
  nand_x1_sg U64198 ( .A(n17572), .B(n41117), .X(n17573) );
  nor_x1_sg U64199 ( .A(n41385), .B(n22855), .X(\L1_0/n4352 ) );
  nor_x1_sg U64200 ( .A(n40029), .B(n22870), .X(\L1_0/n4344 ) );
  nand_x1_sg U64201 ( .A(n40911), .B(n6826), .X(\L2_0/n3523 ) );
  nand_x1_sg U64202 ( .A(n6825), .B(n40026), .X(n6826) );
  nor_x1_sg U64203 ( .A(n51304), .B(n39140), .X(\L1_0/n3543 ) );
  inv_x1_sg U64204 ( .A(n25658), .X(n51304) );
  nor_x1_sg U64205 ( .A(n51307), .B(n40033), .X(\L1_0/n3531 ) );
  inv_x1_sg U64206 ( .A(n25679), .X(n51307) );
  nor_x1_sg U64207 ( .A(n51308), .B(n41380), .X(\L1_0/n3519 ) );
  inv_x1_sg U64208 ( .A(n25700), .X(n51308) );
  nor_x1_sg U64209 ( .A(n51311), .B(n40034), .X(\L1_0/n3495 ) );
  inv_x1_sg U64210 ( .A(n25742), .X(n51311) );
  nor_x1_sg U64211 ( .A(n5940), .B(n41320), .X(n26758) );
  nor_x1_sg U64212 ( .A(n5896), .B(n41322), .X(n21724) );
  nor_x1_sg U64213 ( .A(n5919), .B(n41323), .X(n21771) );
  nor_x1_sg U64214 ( .A(n5784), .B(n39472), .X(n21818) );
  nor_x1_sg U64215 ( .A(n5855), .B(n41322), .X(n21865) );
  nor_x1_sg U64216 ( .A(n5848), .B(n39472), .X(n21911) );
  nor_x1_sg U64217 ( .A(n5910), .B(n39472), .X(n21958) );
  nor_x1_sg U64218 ( .A(n5871), .B(n39924), .X(n22004) );
  nor_x1_sg U64219 ( .A(n5889), .B(n41322), .X(n22051) );
  nor_x1_sg U64220 ( .A(n5794), .B(n39925), .X(n22097) );
  nor_x1_sg U64221 ( .A(n5817), .B(n38946), .X(n22145) );
  nor_x1_sg U64222 ( .A(n5926), .B(n39924), .X(n22192) );
  nor_x1_sg U64223 ( .A(n5810), .B(n41321), .X(n22240) );
  nor_x1_sg U64224 ( .A(n5880), .B(n39925), .X(n22287) );
  nor_x1_sg U64225 ( .A(n5839), .B(n41323), .X(n22335) );
  nor_x1_sg U64226 ( .A(n5803), .B(n41321), .X(n22382) );
  nor_x1_sg U64227 ( .A(n5824), .B(n39473), .X(n22430) );
  nor_x1_sg U64228 ( .A(n5903), .B(n39472), .X(n22476) );
  nor_x1_sg U64229 ( .A(n5947), .B(n41321), .X(n22522) );
  nor_x1_sg U64230 ( .A(n5933), .B(n39924), .X(n22558) );
  nor_x1_sg U64231 ( .A(n22982), .B(n51489), .X(\L1_0/n4280 ) );
  nor_x1_sg U64232 ( .A(n22976), .B(n40030), .X(n22983) );
  nor_x1_sg U64233 ( .A(n24097), .B(n51445), .X(\L1_0/n3960 ) );
  nor_x1_sg U64234 ( .A(n24091), .B(n41360), .X(n24098) );
  nor_x1_sg U64235 ( .A(n24376), .B(n51446), .X(\L1_0/n3880 ) );
  nor_x1_sg U64236 ( .A(n24370), .B(n41357), .X(n24377) );
  nor_x1_sg U64237 ( .A(n24655), .B(n51447), .X(\L1_0/n3800 ) );
  nor_x1_sg U64238 ( .A(n24649), .B(n41335), .X(n24656) );
  nor_x1_sg U64239 ( .A(n24933), .B(n51448), .X(\L1_0/n3720 ) );
  nor_x1_sg U64240 ( .A(n24927), .B(n41332), .X(n24934) );
  nor_x1_sg U64241 ( .A(n25212), .B(n51449), .X(\L1_0/n3640 ) );
  nor_x1_sg U64242 ( .A(n25206), .B(n39923), .X(n25213) );
  nor_x1_sg U64243 ( .A(n25491), .B(n51450), .X(\L1_0/n3560 ) );
  nor_x1_sg U64244 ( .A(n25485), .B(n41371), .X(n25492) );
  nor_x1_sg U64245 ( .A(n25770), .B(n51451), .X(\L1_0/n3480 ) );
  nor_x1_sg U64246 ( .A(n25764), .B(n25640), .X(n25771) );
  nor_x1_sg U64247 ( .A(n26607), .B(n51488), .X(\L1_0/n3240 ) );
  nor_x1_sg U64248 ( .A(n26601), .B(n41353), .X(n26608) );
  nor_x1_sg U64249 ( .A(n23259), .B(n51442), .X(\L1_0/n4200 ) );
  nor_x1_sg U64250 ( .A(n23253), .B(n39903), .X(n23260) );
  nor_x1_sg U64251 ( .A(n23539), .B(n51443), .X(\L1_0/n4120 ) );
  nor_x1_sg U64252 ( .A(n23533), .B(n38960), .X(n23540) );
  nor_x1_sg U64253 ( .A(n23818), .B(n51444), .X(\L1_0/n4040 ) );
  nor_x1_sg U64254 ( .A(n23812), .B(n39461), .X(n23819) );
  nor_x1_sg U64255 ( .A(n5935), .B(n39089), .X(n5103) );
  nand_x1_sg U64256 ( .A(n51201), .B(n51159), .X(n5937) );
  nand_x1_sg U64257 ( .A(n5939), .B(n51180), .X(n5936) );
  nor_x1_sg U64258 ( .A(n5891), .B(n41208), .X(n5109) );
  nand_x1_sg U64259 ( .A(n51182), .B(n51141), .X(n5893) );
  nand_x1_sg U64260 ( .A(n5895), .B(n51161), .X(n5892) );
  nor_x1_sg U64261 ( .A(n5914), .B(n41208), .X(n5106) );
  nand_x1_sg U64262 ( .A(n51183), .B(n51142), .X(n5916) );
  nand_x1_sg U64263 ( .A(n5918), .B(n51162), .X(n5915) );
  nor_x1_sg U64264 ( .A(n5778), .B(n5779), .X(n5124) );
  nand_x1_sg U64265 ( .A(n51184), .B(n51143), .X(n5781) );
  nand_x1_sg U64266 ( .A(n5783), .B(n51163), .X(n5780) );
  nor_x1_sg U64267 ( .A(n5850), .B(n39090), .X(n5115) );
  nand_x1_sg U64268 ( .A(n51185), .B(n51144), .X(n5852) );
  nand_x1_sg U64269 ( .A(n5854), .B(n51164), .X(n5851) );
  nor_x1_sg U64270 ( .A(n5843), .B(n41209), .X(n5116) );
  nand_x1_sg U64271 ( .A(n51186), .B(n51145), .X(n5845) );
  nand_x1_sg U64272 ( .A(n5847), .B(n51165), .X(n5844) );
  nor_x1_sg U64273 ( .A(n5905), .B(n41208), .X(n5107) );
  nand_x1_sg U64274 ( .A(n51187), .B(n51146), .X(n5907) );
  nand_x1_sg U64275 ( .A(n5909), .B(n51166), .X(n5906) );
  nor_x1_sg U64276 ( .A(n5866), .B(n39089), .X(n5112) );
  nand_x1_sg U64277 ( .A(n51188), .B(n51147), .X(n5868) );
  nand_x1_sg U64278 ( .A(n5870), .B(n51167), .X(n5867) );
  nor_x1_sg U64279 ( .A(n5884), .B(n41209), .X(n5110) );
  nand_x1_sg U64280 ( .A(n51189), .B(n51148), .X(n5886) );
  nand_x1_sg U64281 ( .A(n5888), .B(n51168), .X(n5885) );
  nor_x1_sg U64282 ( .A(n5789), .B(n41207), .X(n5122) );
  nand_x1_sg U64283 ( .A(n51190), .B(n51149), .X(n5791) );
  nand_x1_sg U64284 ( .A(n5793), .B(n51169), .X(n5790) );
  nor_x1_sg U64285 ( .A(n5812), .B(n41207), .X(n5119) );
  nand_x1_sg U64286 ( .A(n51191), .B(n51150), .X(n5814) );
  nand_x1_sg U64287 ( .A(n5816), .B(n51170), .X(n5813) );
  nor_x1_sg U64288 ( .A(n5921), .B(n5779), .X(n5105) );
  nand_x1_sg U64289 ( .A(n51192), .B(n51151), .X(n5923) );
  nand_x1_sg U64290 ( .A(n5925), .B(n51171), .X(n5922) );
  nor_x1_sg U64291 ( .A(n5805), .B(n41209), .X(n5120) );
  nand_x1_sg U64292 ( .A(n51193), .B(n51152), .X(n5807) );
  nand_x1_sg U64293 ( .A(n5809), .B(n51172), .X(n5806) );
  nor_x1_sg U64294 ( .A(n5875), .B(n41207), .X(n5111) );
  nand_x1_sg U64295 ( .A(n51194), .B(n51153), .X(n5877) );
  nand_x1_sg U64296 ( .A(n5879), .B(n51173), .X(n5876) );
  nor_x1_sg U64297 ( .A(n5834), .B(n39089), .X(n5117) );
  nand_x1_sg U64298 ( .A(n51195), .B(n51154), .X(n5836) );
  nand_x1_sg U64299 ( .A(n5838), .B(n51174), .X(n5835) );
  nor_x1_sg U64300 ( .A(n5798), .B(n39090), .X(n5121) );
  nand_x1_sg U64301 ( .A(n51196), .B(n51155), .X(n5800) );
  nand_x1_sg U64302 ( .A(n5802), .B(n51175), .X(n5799) );
  nor_x1_sg U64303 ( .A(n5819), .B(n39089), .X(n5118) );
  nand_x1_sg U64304 ( .A(n51197), .B(n51156), .X(n5821) );
  nand_x1_sg U64305 ( .A(n5823), .B(n51176), .X(n5820) );
  nor_x1_sg U64306 ( .A(n5898), .B(n39090), .X(n5108) );
  nand_x1_sg U64307 ( .A(n51198), .B(n51157), .X(n5900) );
  nand_x1_sg U64308 ( .A(n5902), .B(n51177), .X(n5899) );
  nor_x1_sg U64309 ( .A(n5942), .B(n41207), .X(n5102) );
  nand_x1_sg U64310 ( .A(n51199), .B(n51158), .X(n5944) );
  nand_x1_sg U64311 ( .A(n5946), .B(n51178), .X(n5943) );
  nor_x1_sg U64312 ( .A(n22984), .B(n39900), .X(\L1_0/n4279 ) );
  nor_x1_sg U64313 ( .A(n22976), .B(n22982), .X(n22984) );
  nor_x1_sg U64314 ( .A(n23261), .B(n41376), .X(\L1_0/n4199 ) );
  nor_x1_sg U64315 ( .A(n23253), .B(n23259), .X(n23261) );
  nor_x1_sg U64316 ( .A(n23541), .B(n41347), .X(\L1_0/n4119 ) );
  nor_x1_sg U64317 ( .A(n23533), .B(n23539), .X(n23541) );
  nor_x1_sg U64318 ( .A(n23820), .B(n39917), .X(\L1_0/n4039 ) );
  nor_x1_sg U64319 ( .A(n23812), .B(n23818), .X(n23820) );
  nor_x1_sg U64320 ( .A(n24099), .B(n39449), .X(\L1_0/n3959 ) );
  nor_x1_sg U64321 ( .A(n24091), .B(n24097), .X(n24099) );
  nor_x1_sg U64322 ( .A(n24378), .B(n41357), .X(\L1_0/n3879 ) );
  nor_x1_sg U64323 ( .A(n24370), .B(n24376), .X(n24378) );
  nor_x1_sg U64324 ( .A(n24657), .B(n38954), .X(\L1_0/n3799 ) );
  nor_x1_sg U64325 ( .A(n24649), .B(n24655), .X(n24657) );
  nor_x1_sg U64326 ( .A(n24935), .B(n41333), .X(\L1_0/n3719 ) );
  nor_x1_sg U64327 ( .A(n24927), .B(n24933), .X(n24935) );
  nor_x1_sg U64328 ( .A(n25214), .B(n38948), .X(\L1_0/n3639 ) );
  nor_x1_sg U64329 ( .A(n25206), .B(n25212), .X(n25214) );
  nor_x1_sg U64330 ( .A(n25493), .B(n39904), .X(\L1_0/n3559 ) );
  nor_x1_sg U64331 ( .A(n25485), .B(n25491), .X(n25493) );
  nor_x1_sg U64332 ( .A(n25772), .B(n41381), .X(\L1_0/n3479 ) );
  nor_x1_sg U64333 ( .A(n25764), .B(n25770), .X(n25772) );
  nor_x1_sg U64334 ( .A(n26609), .B(n38964), .X(\L1_0/n3239 ) );
  nor_x1_sg U64335 ( .A(n26601), .B(n26607), .X(n26609) );
  nor_x1_sg U64336 ( .A(n51262), .B(n38954), .X(\L1_0/n3871 ) );
  inv_x1_sg U64337 ( .A(n24528), .X(n51262) );
  nor_x1_sg U64338 ( .A(n51265), .B(n41338), .X(\L1_0/n3859 ) );
  inv_x1_sg U64339 ( .A(n24550), .X(n51265) );
  nor_x1_sg U64340 ( .A(n51270), .B(n41337), .X(\L1_0/n3823 ) );
  inv_x1_sg U64341 ( .A(n24613), .X(n51270) );
  nor_x1_sg U64342 ( .A(n51377), .B(n38955), .X(\L1_0/n3811 ) );
  inv_x1_sg U64343 ( .A(n24634), .X(n51377) );
  nor_x1_sg U64344 ( .A(n51212), .B(n38978), .X(\L1_0/n4271 ) );
  inv_x1_sg U64345 ( .A(n23132), .X(n51212) );
  nor_x1_sg U64346 ( .A(n51215), .B(n39902), .X(\L1_0/n4259 ) );
  inv_x1_sg U64347 ( .A(n23154), .X(n51215) );
  nor_x1_sg U64348 ( .A(n51220), .B(n41377), .X(\L1_0/n4223 ) );
  inv_x1_sg U64349 ( .A(n23217), .X(n51220) );
  nor_x1_sg U64350 ( .A(n51337), .B(n39439), .X(\L1_0/n4211 ) );
  inv_x1_sg U64351 ( .A(n23238), .X(n51337) );
  nor_x1_sg U64352 ( .A(n51232), .B(n39461), .X(\L1_0/n4111 ) );
  inv_x1_sg U64353 ( .A(n23691), .X(n51232) );
  nor_x1_sg U64354 ( .A(n51235), .B(n39461), .X(\L1_0/n4099 ) );
  inv_x1_sg U64355 ( .A(n23713), .X(n51235) );
  nor_x1_sg U64356 ( .A(n51240), .B(n41343), .X(\L1_0/n4063 ) );
  inv_x1_sg U64357 ( .A(n23776), .X(n51240) );
  nor_x1_sg U64358 ( .A(n51353), .B(n38958), .X(\L1_0/n4051 ) );
  inv_x1_sg U64359 ( .A(n23797), .X(n51353) );
  nor_x1_sg U64360 ( .A(n51242), .B(n39448), .X(\L1_0/n4031 ) );
  inv_x1_sg U64361 ( .A(n23970), .X(n51242) );
  nor_x1_sg U64362 ( .A(n51245), .B(n39908), .X(\L1_0/n4019 ) );
  inv_x1_sg U64363 ( .A(n23992), .X(n51245) );
  nor_x1_sg U64364 ( .A(n51250), .B(n39909), .X(\L1_0/n3983 ) );
  inv_x1_sg U64365 ( .A(n24055), .X(n51250) );
  nor_x1_sg U64366 ( .A(n51361), .B(n38970), .X(\L1_0/n3971 ) );
  inv_x1_sg U64367 ( .A(n24076), .X(n51361) );
  nor_x1_sg U64368 ( .A(n51252), .B(n41358), .X(\L1_0/n3951 ) );
  inv_x1_sg U64369 ( .A(n24249), .X(n51252) );
  nor_x1_sg U64370 ( .A(n51255), .B(n39910), .X(\L1_0/n3939 ) );
  inv_x1_sg U64371 ( .A(n24271), .X(n51255) );
  nor_x1_sg U64372 ( .A(n51260), .B(n41355), .X(\L1_0/n3903 ) );
  inv_x1_sg U64373 ( .A(n24334), .X(n51260) );
  nor_x1_sg U64374 ( .A(n51369), .B(n38966), .X(\L1_0/n3891 ) );
  inv_x1_sg U64375 ( .A(n24355), .X(n51369) );
  nor_x1_sg U64376 ( .A(n51272), .B(n39921), .X(\L1_0/n3791 ) );
  inv_x1_sg U64377 ( .A(n24806), .X(n51272) );
  nor_x1_sg U64378 ( .A(n51275), .B(n41330), .X(\L1_0/n3779 ) );
  inv_x1_sg U64379 ( .A(n24828), .X(n51275) );
  nor_x1_sg U64380 ( .A(n51280), .B(n38951), .X(\L1_0/n3743 ) );
  inv_x1_sg U64381 ( .A(n24891), .X(n51280) );
  nor_x1_sg U64382 ( .A(n51385), .B(n38952), .X(\L1_0/n3731 ) );
  inv_x1_sg U64383 ( .A(n24912), .X(n51385) );
  nor_x1_sg U64384 ( .A(n51282), .B(n41327), .X(\L1_0/n3711 ) );
  inv_x1_sg U64385 ( .A(n25085), .X(n51282) );
  nor_x1_sg U64386 ( .A(n51285), .B(n38948), .X(\L1_0/n3699 ) );
  inv_x1_sg U64387 ( .A(n25107), .X(n51285) );
  nor_x1_sg U64388 ( .A(n51290), .B(n38948), .X(\L1_0/n3663 ) );
  inv_x1_sg U64389 ( .A(n25170), .X(n51290) );
  nor_x1_sg U64390 ( .A(n51393), .B(n41328), .X(\L1_0/n3651 ) );
  inv_x1_sg U64391 ( .A(n25191), .X(n51393) );
  nor_x1_sg U64392 ( .A(n51292), .B(n41372), .X(\L1_0/n3631 ) );
  inv_x1_sg U64393 ( .A(n25364), .X(n51292) );
  nor_x1_sg U64394 ( .A(n51295), .B(n38975), .X(\L1_0/n3619 ) );
  inv_x1_sg U64395 ( .A(n25386), .X(n51295) );
  nor_x1_sg U64396 ( .A(n51300), .B(n39904), .X(\L1_0/n3583 ) );
  inv_x1_sg U64397 ( .A(n25449), .X(n51300) );
  nor_x1_sg U64398 ( .A(n51401), .B(n38976), .X(\L1_0/n3571 ) );
  inv_x1_sg U64399 ( .A(n25470), .X(n51401) );
  nor_x1_sg U64400 ( .A(n51302), .B(n41383), .X(\L1_0/n3551 ) );
  inv_x1_sg U64401 ( .A(n25643), .X(n51302) );
  nor_x1_sg U64402 ( .A(n51305), .B(n40034), .X(\L1_0/n3539 ) );
  inv_x1_sg U64403 ( .A(n25665), .X(n51305) );
  nor_x1_sg U64404 ( .A(n51310), .B(n40035), .X(\L1_0/n3503 ) );
  inv_x1_sg U64405 ( .A(n25728), .X(n51310) );
  nor_x1_sg U64406 ( .A(n51409), .B(n41381), .X(\L1_0/n3491 ) );
  inv_x1_sg U64407 ( .A(n25749), .X(n51409) );
  nor_x1_sg U64408 ( .A(n51314), .B(n41352), .X(\L1_0/n3311 ) );
  inv_x1_sg U64409 ( .A(n26480), .X(n51314) );
  nor_x1_sg U64410 ( .A(n51317), .B(n41351), .X(\L1_0/n3299 ) );
  inv_x1_sg U64411 ( .A(n26502), .X(n51317) );
  nor_x1_sg U64412 ( .A(n51322), .B(n41350), .X(\L1_0/n3263 ) );
  inv_x1_sg U64413 ( .A(n26565), .X(n51322) );
  nor_x1_sg U64414 ( .A(n51418), .B(n41352), .X(\L1_0/n3251 ) );
  inv_x1_sg U64415 ( .A(n26586), .X(n51418) );
  nor_x1_sg U64416 ( .A(n51222), .B(n39457), .X(\L1_0/n4191 ) );
  inv_x1_sg U64417 ( .A(n23412), .X(n51222) );
  nor_x1_sg U64418 ( .A(n51225), .B(n39914), .X(\L1_0/n4179 ) );
  inv_x1_sg U64419 ( .A(n23434), .X(n51225) );
  nor_x1_sg U64420 ( .A(n51230), .B(n41347), .X(\L1_0/n4143 ) );
  inv_x1_sg U64421 ( .A(n23497), .X(n51230) );
  nor_x1_sg U64422 ( .A(n51345), .B(n38961), .X(\L1_0/n4131 ) );
  inv_x1_sg U64423 ( .A(n23518), .X(n51345) );
  nor_x1_sg U64424 ( .A(n51204), .B(n40030), .X(\L1_0/n4343 ) );
  inv_x1_sg U64425 ( .A(n22870), .X(n51204) );
  nor_x1_sg U64426 ( .A(n51202), .B(n40031), .X(\L1_0/n4351 ) );
  inv_x1_sg U64427 ( .A(n22855), .X(n51202) );
  nor_x1_sg U64428 ( .A(n51263), .B(n41335), .X(\L1_0/n3867 ) );
  inv_x1_sg U64429 ( .A(n24536), .X(n51263) );
  nor_x1_sg U64430 ( .A(n51264), .B(n39464), .X(\L1_0/n3863 ) );
  inv_x1_sg U64431 ( .A(n24543), .X(n51264) );
  nor_x1_sg U64432 ( .A(n51266), .B(n39918), .X(\L1_0/n3855 ) );
  inv_x1_sg U64433 ( .A(n24557), .X(n51266) );
  nor_x1_sg U64434 ( .A(n51267), .B(n39463), .X(\L1_0/n3851 ) );
  inv_x1_sg U64435 ( .A(n24564), .X(n51267) );
  nor_x1_sg U64436 ( .A(n51268), .B(n41335), .X(\L1_0/n3839 ) );
  inv_x1_sg U64437 ( .A(n24585), .X(n51268) );
  nor_x1_sg U64438 ( .A(n51269), .B(n39919), .X(\L1_0/n3831 ) );
  inv_x1_sg U64439 ( .A(n24599), .X(n51269) );
  nor_x1_sg U64440 ( .A(n51271), .B(n39918), .X(\L1_0/n3815 ) );
  inv_x1_sg U64441 ( .A(n24627), .X(n51271) );
  nor_x1_sg U64442 ( .A(n51378), .B(n39463), .X(\L1_0/n3807 ) );
  inv_x1_sg U64443 ( .A(n24639), .X(n51378) );
  nor_x1_sg U64444 ( .A(n51213), .B(n38979), .X(\L1_0/n4267 ) );
  inv_x1_sg U64445 ( .A(n23140), .X(n51213) );
  nor_x1_sg U64446 ( .A(n51214), .B(n41377), .X(\L1_0/n4263 ) );
  inv_x1_sg U64447 ( .A(n23147), .X(n51214) );
  nor_x1_sg U64448 ( .A(n51216), .B(n41377), .X(\L1_0/n4255 ) );
  inv_x1_sg U64449 ( .A(n23161), .X(n51216) );
  nor_x1_sg U64450 ( .A(n51217), .B(n39440), .X(\L1_0/n4251 ) );
  inv_x1_sg U64451 ( .A(n23168), .X(n51217) );
  nor_x1_sg U64452 ( .A(n51218), .B(n39440), .X(\L1_0/n4239 ) );
  inv_x1_sg U64453 ( .A(n23189), .X(n51218) );
  nor_x1_sg U64454 ( .A(n51219), .B(n41378), .X(\L1_0/n4231 ) );
  inv_x1_sg U64455 ( .A(n23203), .X(n51219) );
  nor_x1_sg U64456 ( .A(n51221), .B(n39439), .X(\L1_0/n4215 ) );
  inv_x1_sg U64457 ( .A(n23231), .X(n51221) );
  nor_x1_sg U64458 ( .A(n51338), .B(n38978), .X(\L1_0/n4207 ) );
  inv_x1_sg U64459 ( .A(n23243), .X(n51338) );
  nor_x1_sg U64460 ( .A(n51233), .B(n39460), .X(\L1_0/n4107 ) );
  inv_x1_sg U64461 ( .A(n23699), .X(n51233) );
  nor_x1_sg U64462 ( .A(n51234), .B(n38957), .X(\L1_0/n4103 ) );
  inv_x1_sg U64463 ( .A(n23706), .X(n51234) );
  nor_x1_sg U64464 ( .A(n51236), .B(n41341), .X(\L1_0/n4095 ) );
  inv_x1_sg U64465 ( .A(n23720), .X(n51236) );
  nor_x1_sg U64466 ( .A(n51237), .B(n39916), .X(\L1_0/n4091 ) );
  inv_x1_sg U64467 ( .A(n23727), .X(n51237) );
  nor_x1_sg U64468 ( .A(n51238), .B(n38957), .X(\L1_0/n4079 ) );
  inv_x1_sg U64469 ( .A(n23748), .X(n51238) );
  nor_x1_sg U64470 ( .A(n51239), .B(n39916), .X(\L1_0/n4071 ) );
  inv_x1_sg U64471 ( .A(n23762), .X(n51239) );
  nor_x1_sg U64472 ( .A(n51241), .B(n39917), .X(\L1_0/n4055 ) );
  inv_x1_sg U64473 ( .A(n23790), .X(n51241) );
  nor_x1_sg U64474 ( .A(n51354), .B(n39460), .X(\L1_0/n4047 ) );
  inv_x1_sg U64475 ( .A(n23802), .X(n51354) );
  nor_x1_sg U64476 ( .A(n51243), .B(n41360), .X(\L1_0/n4027 ) );
  inv_x1_sg U64477 ( .A(n23978), .X(n51243) );
  nor_x1_sg U64478 ( .A(n51244), .B(n39908), .X(\L1_0/n4023 ) );
  inv_x1_sg U64479 ( .A(n23985), .X(n51244) );
  nor_x1_sg U64480 ( .A(n51246), .B(n41361), .X(\L1_0/n4015 ) );
  inv_x1_sg U64481 ( .A(n23999), .X(n51246) );
  nor_x1_sg U64482 ( .A(n51247), .B(n41362), .X(\L1_0/n4011 ) );
  inv_x1_sg U64483 ( .A(n24006), .X(n51247) );
  nor_x1_sg U64484 ( .A(n51248), .B(n38969), .X(\L1_0/n3999 ) );
  inv_x1_sg U64485 ( .A(n24027), .X(n51248) );
  nor_x1_sg U64486 ( .A(n51249), .B(n39448), .X(\L1_0/n3991 ) );
  inv_x1_sg U64487 ( .A(n24041), .X(n51249) );
  nor_x1_sg U64488 ( .A(n51251), .B(n39449), .X(\L1_0/n3975 ) );
  inv_x1_sg U64489 ( .A(n24069), .X(n51251) );
  nor_x1_sg U64490 ( .A(n51362), .B(n38969), .X(\L1_0/n3967 ) );
  inv_x1_sg U64491 ( .A(n24081), .X(n51362) );
  nor_x1_sg U64492 ( .A(n51253), .B(n39910), .X(\L1_0/n3947 ) );
  inv_x1_sg U64493 ( .A(n24257), .X(n51253) );
  nor_x1_sg U64494 ( .A(n51254), .B(n41357), .X(\L1_0/n3943 ) );
  inv_x1_sg U64495 ( .A(n24264), .X(n51254) );
  nor_x1_sg U64496 ( .A(n51256), .B(n41358), .X(\L1_0/n3935 ) );
  inv_x1_sg U64497 ( .A(n24278), .X(n51256) );
  nor_x1_sg U64498 ( .A(n51257), .B(n41357), .X(\L1_0/n3931 ) );
  inv_x1_sg U64499 ( .A(n24285), .X(n51257) );
  nor_x1_sg U64500 ( .A(n51258), .B(n41356), .X(\L1_0/n3919 ) );
  inv_x1_sg U64501 ( .A(n24306), .X(n51258) );
  nor_x1_sg U64502 ( .A(n51259), .B(n39451), .X(\L1_0/n3911 ) );
  inv_x1_sg U64503 ( .A(n24320), .X(n51259) );
  nor_x1_sg U64504 ( .A(n51261), .B(n39910), .X(\L1_0/n3895 ) );
  inv_x1_sg U64505 ( .A(n24348), .X(n51261) );
  nor_x1_sg U64506 ( .A(n51370), .B(n39451), .X(\L1_0/n3887 ) );
  inv_x1_sg U64507 ( .A(n24360), .X(n51370) );
  nor_x1_sg U64508 ( .A(n51273), .B(n41331), .X(\L1_0/n3787 ) );
  inv_x1_sg U64509 ( .A(n24814), .X(n51273) );
  nor_x1_sg U64510 ( .A(n51274), .B(n39921), .X(\L1_0/n3783 ) );
  inv_x1_sg U64511 ( .A(n24821), .X(n51274) );
  nor_x1_sg U64512 ( .A(n51276), .B(n39921), .X(\L1_0/n3775 ) );
  inv_x1_sg U64513 ( .A(n24835), .X(n51276) );
  nor_x1_sg U64514 ( .A(n51277), .B(n38952), .X(\L1_0/n3771 ) );
  inv_x1_sg U64515 ( .A(n24842), .X(n51277) );
  nor_x1_sg U64516 ( .A(n51278), .B(n41330), .X(\L1_0/n3759 ) );
  inv_x1_sg U64517 ( .A(n24863), .X(n51278) );
  nor_x1_sg U64518 ( .A(n51279), .B(n39920), .X(\L1_0/n3751 ) );
  inv_x1_sg U64519 ( .A(n24877), .X(n51279) );
  nor_x1_sg U64520 ( .A(n51281), .B(n39466), .X(\L1_0/n3735 ) );
  inv_x1_sg U64521 ( .A(n24905), .X(n51281) );
  nor_x1_sg U64522 ( .A(n51386), .B(n41333), .X(\L1_0/n3727 ) );
  inv_x1_sg U64523 ( .A(n24917), .X(n51386) );
  nor_x1_sg U64524 ( .A(n51283), .B(n41326), .X(\L1_0/n3707 ) );
  inv_x1_sg U64525 ( .A(n25093), .X(n51283) );
  nor_x1_sg U64526 ( .A(n51284), .B(n39923), .X(\L1_0/n3703 ) );
  inv_x1_sg U64527 ( .A(n25100), .X(n51284) );
  nor_x1_sg U64528 ( .A(n51286), .B(n38949), .X(\L1_0/n3695 ) );
  inv_x1_sg U64529 ( .A(n25114), .X(n51286) );
  nor_x1_sg U64530 ( .A(n51287), .B(n41327), .X(\L1_0/n3691 ) );
  inv_x1_sg U64531 ( .A(n25121), .X(n51287) );
  nor_x1_sg U64532 ( .A(n51288), .B(n41325), .X(\L1_0/n3679 ) );
  inv_x1_sg U64533 ( .A(n25142), .X(n51288) );
  nor_x1_sg U64534 ( .A(n51289), .B(n41328), .X(\L1_0/n3671 ) );
  inv_x1_sg U64535 ( .A(n25156), .X(n51289) );
  nor_x1_sg U64536 ( .A(n51291), .B(n39469), .X(\L1_0/n3655 ) );
  inv_x1_sg U64537 ( .A(n25184), .X(n51291) );
  nor_x1_sg U64538 ( .A(n51394), .B(n39922), .X(\L1_0/n3647 ) );
  inv_x1_sg U64539 ( .A(n25196), .X(n51394) );
  nor_x1_sg U64540 ( .A(n51293), .B(n39442), .X(\L1_0/n3627 ) );
  inv_x1_sg U64541 ( .A(n25372), .X(n51293) );
  nor_x1_sg U64542 ( .A(n51294), .B(n39905), .X(\L1_0/n3623 ) );
  inv_x1_sg U64543 ( .A(n25379), .X(n51294) );
  nor_x1_sg U64544 ( .A(n51296), .B(n39443), .X(\L1_0/n3615 ) );
  inv_x1_sg U64545 ( .A(n25393), .X(n51296) );
  nor_x1_sg U64546 ( .A(n51297), .B(n39443), .X(\L1_0/n3611 ) );
  inv_x1_sg U64547 ( .A(n25400), .X(n51297) );
  nor_x1_sg U64548 ( .A(n51298), .B(n39443), .X(\L1_0/n3599 ) );
  inv_x1_sg U64549 ( .A(n25421), .X(n51298) );
  nor_x1_sg U64550 ( .A(n51299), .B(n39442), .X(\L1_0/n3591 ) );
  inv_x1_sg U64551 ( .A(n25435), .X(n51299) );
  nor_x1_sg U64552 ( .A(n51301), .B(n41372), .X(\L1_0/n3575 ) );
  inv_x1_sg U64553 ( .A(n25463), .X(n51301) );
  nor_x1_sg U64554 ( .A(n51402), .B(n38975), .X(\L1_0/n3567 ) );
  inv_x1_sg U64555 ( .A(n25475), .X(n51402) );
  nor_x1_sg U64556 ( .A(n51303), .B(n41382), .X(\L1_0/n3547 ) );
  inv_x1_sg U64557 ( .A(n25651), .X(n51303) );
  nor_x1_sg U64558 ( .A(n51306), .B(n41382), .X(\L1_0/n3535 ) );
  inv_x1_sg U64559 ( .A(n25672), .X(n51306) );
  nor_x1_sg U64560 ( .A(n51309), .B(n39139), .X(\L1_0/n3511 ) );
  inv_x1_sg U64561 ( .A(n25714), .X(n51309) );
  nor_x1_sg U64562 ( .A(n51410), .B(n39901), .X(\L1_0/n3487 ) );
  inv_x1_sg U64563 ( .A(n25754), .X(n51410) );
  nor_x1_sg U64564 ( .A(n51315), .B(n41352), .X(\L1_0/n3307 ) );
  inv_x1_sg U64565 ( .A(n26488), .X(n51315) );
  nor_x1_sg U64566 ( .A(n51316), .B(n41353), .X(\L1_0/n3303 ) );
  inv_x1_sg U64567 ( .A(n26495), .X(n51316) );
  nor_x1_sg U64568 ( .A(n51318), .B(n39913), .X(\L1_0/n3295 ) );
  inv_x1_sg U64569 ( .A(n26509), .X(n51318) );
  nor_x1_sg U64570 ( .A(n51319), .B(n41352), .X(\L1_0/n3291 ) );
  inv_x1_sg U64571 ( .A(n26516), .X(n51319) );
  nor_x1_sg U64572 ( .A(n51320), .B(n41350), .X(\L1_0/n3279 ) );
  inv_x1_sg U64573 ( .A(n26537), .X(n51320) );
  nor_x1_sg U64574 ( .A(n51321), .B(n41353), .X(\L1_0/n3271 ) );
  inv_x1_sg U64575 ( .A(n26551), .X(n51321) );
  nor_x1_sg U64576 ( .A(n51323), .B(n39455), .X(\L1_0/n3255 ) );
  inv_x1_sg U64577 ( .A(n26579), .X(n51323) );
  nor_x1_sg U64578 ( .A(n51419), .B(n41351), .X(\L1_0/n3247 ) );
  inv_x1_sg U64579 ( .A(n26591), .X(n51419) );
  nor_x1_sg U64580 ( .A(n51223), .B(n38960), .X(\L1_0/n4187 ) );
  inv_x1_sg U64581 ( .A(n23420), .X(n51223) );
  nor_x1_sg U64582 ( .A(n51224), .B(n38960), .X(\L1_0/n4183 ) );
  inv_x1_sg U64583 ( .A(n23427), .X(n51224) );
  nor_x1_sg U64584 ( .A(n51226), .B(n39915), .X(\L1_0/n4175 ) );
  inv_x1_sg U64585 ( .A(n23441), .X(n51226) );
  nor_x1_sg U64586 ( .A(n51227), .B(n41348), .X(\L1_0/n4171 ) );
  inv_x1_sg U64587 ( .A(n23448), .X(n51227) );
  nor_x1_sg U64588 ( .A(n51228), .B(n39914), .X(\L1_0/n4159 ) );
  inv_x1_sg U64589 ( .A(n23469), .X(n51228) );
  nor_x1_sg U64590 ( .A(n51229), .B(n41346), .X(\L1_0/n4151 ) );
  inv_x1_sg U64591 ( .A(n23483), .X(n51229) );
  nor_x1_sg U64592 ( .A(n51231), .B(n41347), .X(\L1_0/n4135 ) );
  inv_x1_sg U64593 ( .A(n23511), .X(n51231) );
  nor_x1_sg U64594 ( .A(n51346), .B(n41348), .X(\L1_0/n4127 ) );
  inv_x1_sg U64595 ( .A(n23523), .X(n51346) );
  nand_x1_sg U64596 ( .A(n41211), .B(n26755), .X(\L1_0/n3195 ) );
  nor_x1_sg U64597 ( .A(n5941), .B(n51509), .X(n26757) );
  nor_x1_sg U64598 ( .A(n5938), .B(n26786), .X(n26756) );
  nand_x1_sg U64599 ( .A(n41211), .B(n21768), .X(\L1_0/n4507 ) );
  nor_x1_sg U64600 ( .A(n5920), .B(n51491), .X(n21770) );
  nor_x1_sg U64601 ( .A(n5917), .B(n21794), .X(n21769) );
  nand_x1_sg U64602 ( .A(n41211), .B(n21908), .X(\L1_0/n4495 ) );
  nor_x1_sg U64603 ( .A(n5849), .B(n51494), .X(n21910) );
  nor_x1_sg U64604 ( .A(n5846), .B(n21934), .X(n21909) );
  nand_x1_sg U64605 ( .A(n41213), .B(n22048), .X(\L1_0/n4483 ) );
  nor_x1_sg U64606 ( .A(n5890), .B(n51497), .X(n22050) );
  nor_x1_sg U64607 ( .A(n5887), .B(n22073), .X(n22049) );
  nand_x1_sg U64608 ( .A(n41211), .B(n22189), .X(\L1_0/n4471 ) );
  nor_x1_sg U64609 ( .A(n5927), .B(n51500), .X(n22191) );
  nor_x1_sg U64610 ( .A(n5924), .B(n22216), .X(n22190) );
  nand_x1_sg U64611 ( .A(n41214), .B(n22332), .X(\L1_0/n4459 ) );
  nor_x1_sg U64612 ( .A(n5840), .B(n51503), .X(n22334) );
  nor_x1_sg U64613 ( .A(n5837), .B(n22358), .X(n22333) );
  nand_x1_sg U64614 ( .A(n41212), .B(n22473), .X(\L1_0/n4447 ) );
  nor_x1_sg U64615 ( .A(n5904), .B(n51506), .X(n22475) );
  nor_x1_sg U64616 ( .A(n5901), .B(n22498), .X(n22474) );
  nor_x1_sg U64617 ( .A(n26031), .B(n26032), .X(\L1_0/n3400 ) );
  nand_x1_sg U64618 ( .A(n39482), .B(n38940), .X(n26031) );
  nand_x1_sg U64619 ( .A(n5747), .B(n41312), .X(n26032) );
  nand_x1_sg U64620 ( .A(n39093), .B(n21815), .X(\L1_0/n4503 ) );
  nor_x1_sg U64621 ( .A(n5785), .B(n51492), .X(n21817) );
  nor_x1_sg U64622 ( .A(n5782), .B(n21841), .X(n21816) );
  nand_x1_sg U64623 ( .A(n39093), .B(n21955), .X(\L1_0/n4491 ) );
  nor_x1_sg U64624 ( .A(n5911), .B(n51495), .X(n21957) );
  nor_x1_sg U64625 ( .A(n5908), .B(n21980), .X(n21956) );
  nand_x1_sg U64626 ( .A(n41213), .B(n22094), .X(\L1_0/n4479 ) );
  nor_x1_sg U64627 ( .A(n5795), .B(n51498), .X(n22096) );
  nor_x1_sg U64628 ( .A(n5792), .B(n22121), .X(n22095) );
  nand_x1_sg U64629 ( .A(n41212), .B(n22237), .X(\L1_0/n4467 ) );
  nor_x1_sg U64630 ( .A(n5811), .B(n51501), .X(n22239) );
  nor_x1_sg U64631 ( .A(n5808), .B(n22263), .X(n22238) );
  nand_x1_sg U64632 ( .A(n41213), .B(n22379), .X(\L1_0/n4455 ) );
  nor_x1_sg U64633 ( .A(n5804), .B(n51504), .X(n22381) );
  nor_x1_sg U64634 ( .A(n5801), .B(n22406), .X(n22380) );
  nand_x1_sg U64635 ( .A(n41213), .B(n22519), .X(\L1_0/n4443 ) );
  nor_x1_sg U64636 ( .A(n5948), .B(n51507), .X(n22521) );
  nor_x1_sg U64637 ( .A(n5945), .B(n22538), .X(n22520) );
  nand_x1_sg U64638 ( .A(n39092), .B(n21721), .X(\L1_0/n4511 ) );
  nor_x1_sg U64639 ( .A(n5897), .B(n51490), .X(n21723) );
  nor_x1_sg U64640 ( .A(n5894), .B(n21747), .X(n21722) );
  nand_x1_sg U64641 ( .A(n41214), .B(n21862), .X(\L1_0/n4499 ) );
  nor_x1_sg U64642 ( .A(n5856), .B(n51493), .X(n21864) );
  nor_x1_sg U64643 ( .A(n5853), .B(n21887), .X(n21863) );
  nand_x1_sg U64644 ( .A(n41214), .B(n22001), .X(\L1_0/n4487 ) );
  nor_x1_sg U64645 ( .A(n5872), .B(n51496), .X(n22003) );
  nor_x1_sg U64646 ( .A(n5869), .B(n22027), .X(n22002) );
  nand_x1_sg U64647 ( .A(n41212), .B(n22142), .X(\L1_0/n4475 ) );
  nor_x1_sg U64648 ( .A(n5818), .B(n51499), .X(n22144) );
  nor_x1_sg U64649 ( .A(n5815), .B(n22168), .X(n22143) );
  nand_x1_sg U64650 ( .A(n41212), .B(n22284), .X(\L1_0/n4463 ) );
  nor_x1_sg U64651 ( .A(n5881), .B(n51502), .X(n22286) );
  nor_x1_sg U64652 ( .A(n5878), .B(n22311), .X(n22285) );
  nand_x1_sg U64653 ( .A(n39092), .B(n22427), .X(\L1_0/n4451 ) );
  nor_x1_sg U64654 ( .A(n5825), .B(n51505), .X(n22429) );
  nor_x1_sg U64655 ( .A(n5822), .B(n22452), .X(n22428) );
  nand_x1_sg U64656 ( .A(n40902), .B(n16674), .X(\L2_0/n2547 ) );
  nand_x1_sg U64657 ( .A(n16673), .B(n41217), .X(n16674) );
  nand_x1_sg U64658 ( .A(n40901), .B(n16680), .X(\L2_0/n2543 ) );
  nand_x1_sg U64659 ( .A(n16679), .B(n41216), .X(n16680) );
  nand_x1_sg U64660 ( .A(n38885), .B(n16686), .X(\L2_0/n2539 ) );
  nand_x1_sg U64661 ( .A(n16685), .B(n41217), .X(n16686) );
  nand_x1_sg U64662 ( .A(n38885), .B(n16692), .X(\L2_0/n2535 ) );
  nand_x1_sg U64663 ( .A(n16691), .B(n41219), .X(n16692) );
  nand_x1_sg U64664 ( .A(n40903), .B(n16734), .X(\L2_0/n2507 ) );
  nand_x1_sg U64665 ( .A(n16733), .B(n39096), .X(n16734) );
  nand_x1_sg U64666 ( .A(n40903), .B(n16752), .X(\L2_0/n2495 ) );
  nand_x1_sg U64667 ( .A(n16751), .B(n41217), .X(n16752) );
  nand_x1_sg U64668 ( .A(n38885), .B(n16650), .X(\L2_0/n2563 ) );
  nand_x1_sg U64669 ( .A(n16649), .B(n41218), .X(n16650) );
  nand_x1_sg U64670 ( .A(n40902), .B(n16660), .X(\L2_0/n2555 ) );
  nand_x1_sg U64671 ( .A(n16659), .B(n39096), .X(n16660) );
  nand_x1_sg U64672 ( .A(n40903), .B(n16667), .X(\L2_0/n2551 ) );
  nand_x1_sg U64673 ( .A(n41219), .B(n16666), .X(n16667) );
  nand_x1_sg U64674 ( .A(n40901), .B(n16698), .X(\L2_0/n2531 ) );
  nand_x1_sg U64675 ( .A(n16697), .B(n41218), .X(n16698) );
  nand_x1_sg U64676 ( .A(n40901), .B(n16704), .X(\L2_0/n2527 ) );
  nand_x1_sg U64677 ( .A(n16703), .B(n41217), .X(n16704) );
  nand_x1_sg U64678 ( .A(n40904), .B(n16710), .X(\L2_0/n2523 ) );
  nand_x1_sg U64679 ( .A(n16709), .B(n41218), .X(n16710) );
  nand_x1_sg U64680 ( .A(n40902), .B(n16716), .X(\L2_0/n2519 ) );
  nand_x1_sg U64681 ( .A(n16715), .B(n39096), .X(n16716) );
  nand_x1_sg U64682 ( .A(n40904), .B(n16722), .X(\L2_0/n2515 ) );
  nand_x1_sg U64683 ( .A(n16721), .B(n41219), .X(n16722) );
  nand_x1_sg U64684 ( .A(n40902), .B(n16728), .X(\L2_0/n2511 ) );
  nand_x1_sg U64685 ( .A(n16727), .B(n41218), .X(n16728) );
  nand_x1_sg U64686 ( .A(n40903), .B(n16740), .X(\L2_0/n2503 ) );
  nand_x1_sg U64687 ( .A(n16739), .B(n41219), .X(n16740) );
  nand_x1_sg U64688 ( .A(n40904), .B(n16746), .X(\L2_0/n2499 ) );
  nand_x1_sg U64689 ( .A(n16745), .B(n41216), .X(n16746) );
  inv_x1_sg U64690 ( .A(n5894), .X(n51182) );
  inv_x1_sg U64691 ( .A(n5917), .X(n51183) );
  inv_x1_sg U64692 ( .A(n5782), .X(n51184) );
  inv_x1_sg U64693 ( .A(n5853), .X(n51185) );
  inv_x1_sg U64694 ( .A(n5846), .X(n51186) );
  inv_x1_sg U64695 ( .A(n5908), .X(n51187) );
  inv_x1_sg U64696 ( .A(n5869), .X(n51188) );
  inv_x1_sg U64697 ( .A(n5887), .X(n51189) );
  inv_x1_sg U64698 ( .A(n5792), .X(n51190) );
  inv_x1_sg U64699 ( .A(n5815), .X(n51191) );
  inv_x1_sg U64700 ( .A(n5924), .X(n51192) );
  inv_x1_sg U64701 ( .A(n5808), .X(n51193) );
  inv_x1_sg U64702 ( .A(n5878), .X(n51194) );
  inv_x1_sg U64703 ( .A(n5837), .X(n51195) );
  inv_x1_sg U64704 ( .A(n5801), .X(n51196) );
  inv_x1_sg U64705 ( .A(n5822), .X(n51197) );
  inv_x1_sg U64706 ( .A(n5901), .X(n51198) );
  inv_x1_sg U64707 ( .A(n5938), .X(n51201) );
  nand_x1_sg U64708 ( .A(n40025), .B(n6783), .X(n6784) );
  nand_x1_sg U64709 ( .A(n38940), .B(n5736), .X(n5735) );
  nand_x1_sg U64710 ( .A(n41113), .B(n5741), .X(n5740) );
  nand_x1_sg U64711 ( .A(n41115), .B(n5757), .X(n5756) );
  nand_x1_sg U64712 ( .A(n39254), .B(n5751), .X(n5750) );
  nand_x1_sg U64713 ( .A(n39254), .B(n5762), .X(n5761) );
  nand_x1_sg U64714 ( .A(n41115), .B(n5766), .X(n5765) );
  nand_x1_sg U64715 ( .A(n42372), .B(n5753), .X(n5752) );
  nand_x1_sg U64716 ( .A(n41115), .B(n5760), .X(n5759) );
  nand_x1_sg U64717 ( .A(n39254), .B(n5734), .X(n5732) );
  nand_x1_sg U64718 ( .A(n38940), .B(n5738), .X(n5737) );
  nand_x1_sg U64719 ( .A(n41114), .B(n5749), .X(n5748) );
  nand_x1_sg U64720 ( .A(n41114), .B(n5755), .X(n25955) );
  nand_x1_sg U64721 ( .A(n39254), .B(n5739), .X(n25962) );
  nand_x1_sg U64722 ( .A(n41114), .B(n5743), .X(n25975) );
  nand_x1_sg U64723 ( .A(n38940), .B(n5768), .X(n5767) );
  nand_x1_sg U64724 ( .A(n41115), .B(n5754), .X(n25988) );
  nand_x1_sg U64725 ( .A(n41113), .B(n5742), .X(n26001) );
  nand_x1_sg U64726 ( .A(n42372), .B(n5764), .X(n5763) );
  nor_x1_sg U64727 ( .A(n39728), .B(n41043), .X(n42388) );
  nor_x1_sg U64728 ( .A(n39770), .B(n40087), .X(n16966) );
  nor_x1_sg U64729 ( .A(n24101), .B(n42119), .X(n20575) );
  nor_x1_sg U64730 ( .A(n40040), .B(n40084), .X(n7104) );
  nor_x1_sg U64731 ( .A(n42089), .B(n40179), .X(n7922) );
  nor_x1_sg U64732 ( .A(n42130), .B(n40211), .X(n8740) );
  nor_x1_sg U64733 ( .A(n40044), .B(n40207), .X(n9560) );
  nor_x1_sg U64734 ( .A(n40046), .B(n40203), .X(n10379) );
  nor_x1_sg U64735 ( .A(n40048), .B(n40199), .X(n11198) );
  nor_x1_sg U64736 ( .A(n11996), .B(n40195), .X(n12017) );
  nor_x1_sg U64737 ( .A(n12815), .B(n40192), .X(n12836) );
  nor_x1_sg U64738 ( .A(n40066), .B(n40175), .X(n13655) );
  nor_x1_sg U64739 ( .A(n40053), .B(n40188), .X(n14474) );
  nor_x1_sg U64740 ( .A(n40056), .B(n40171), .X(n15293) );
  nor_x1_sg U64741 ( .A(n16091), .B(n40168), .X(n16112) );
  nor_x1_sg U64742 ( .A(n40060), .B(n40215), .X(n17750) );
  nor_x1_sg U64743 ( .A(n40062), .B(n40183), .X(n18571) );
  nor_x1_sg U64744 ( .A(n6687), .B(n20504), .X(n20503) );
  nand_x1_sg U64745 ( .A(n20504), .B(n38701), .X(n20505) );
  nor_x1_sg U64746 ( .A(n6655), .B(n19847), .X(n19846) );
  nand_x1_sg U64747 ( .A(n19847), .B(n38673), .X(n19848) );
  nor_x1_sg U64748 ( .A(n42343), .B(n21273), .X(n21272) );
  nand_x1_sg U64749 ( .A(n21273), .B(n38720), .X(n21274) );
  nand_x1_sg U64750 ( .A(n40104), .B(n24100), .X(n42374) );
  nand_x1_sg U64751 ( .A(n40103), .B(n24379), .X(n42373) );
  nand_x1_sg U64752 ( .A(n40102), .B(n26610), .X(n42371) );
  nor_x1_sg U64753 ( .A(n42340), .B(n28138), .X(n28137) );
  nand_x1_sg U64754 ( .A(n28138), .B(n38714), .X(n28139) );
  inv_x1_sg U64755 ( .A(n25495), .X(n51139) );
  nand_x1_sg U64756 ( .A(n40102), .B(n26332), .X(n25640) );
  nand_x1_sg U64757 ( .A(n40103), .B(n23542), .X(n23409) );
  nand_x1_sg U64758 ( .A(n40102), .B(n23821), .X(n42375) );
  nand_x1_sg U64759 ( .A(n40104), .B(n24658), .X(n24525) );
  nand_x1_sg U64760 ( .A(n40103), .B(n24936), .X(n24803) );
  nand_x1_sg U64761 ( .A(n40104), .B(n25215), .X(n25082) );
  nor_x1_sg U64762 ( .A(n39728), .B(n41052), .X(n42377) );
  nor_x1_sg U64763 ( .A(n39727), .B(n41274), .X(n5954) );
  nand_x1_sg U64764 ( .A(n46966), .B(n46942), .X(n22766) );
  nand_x1_sg U64765 ( .A(n22768), .B(n22767), .X(n22765) );
  inv_x1_sg U64766 ( .A(n22768), .X(n46966) );
  nand_x1_sg U64767 ( .A(n23045), .B(n23044), .X(n23042) );
  inv_x1_sg U64768 ( .A(n23045), .X(n47256) );
  nand_x1_sg U64769 ( .A(n47541), .B(n47518), .X(n23323) );
  nand_x1_sg U64770 ( .A(n23325), .B(n23324), .X(n23322) );
  inv_x1_sg U64771 ( .A(n23325), .X(n47541) );
  nand_x1_sg U64772 ( .A(n47826), .B(n47803), .X(n23602) );
  nand_x1_sg U64773 ( .A(n23604), .B(n23603), .X(n23601) );
  inv_x1_sg U64774 ( .A(n23604), .X(n47826) );
  nand_x1_sg U64775 ( .A(n48111), .B(n48088), .X(n23881) );
  nand_x1_sg U64776 ( .A(n23883), .B(n23882), .X(n23880) );
  inv_x1_sg U64777 ( .A(n23883), .X(n48111) );
  nand_x1_sg U64778 ( .A(n48396), .B(n48373), .X(n24160) );
  nand_x1_sg U64779 ( .A(n24162), .B(n24161), .X(n24159) );
  inv_x1_sg U64780 ( .A(n24162), .X(n48396) );
  nand_x1_sg U64781 ( .A(n48681), .B(n48658), .X(n24439) );
  nand_x1_sg U64782 ( .A(n24441), .B(n24440), .X(n24438) );
  inv_x1_sg U64783 ( .A(n24441), .X(n48681) );
  nand_x1_sg U64784 ( .A(n48967), .B(n48944), .X(n24717) );
  nand_x1_sg U64785 ( .A(n24719), .B(n24718), .X(n24716) );
  inv_x1_sg U64786 ( .A(n24719), .X(n48967) );
  nand_x1_sg U64787 ( .A(n49254), .B(n49231), .X(n24996) );
  nand_x1_sg U64788 ( .A(n24998), .B(n24997), .X(n24995) );
  inv_x1_sg U64789 ( .A(n24998), .X(n49254) );
  nand_x1_sg U64790 ( .A(n49540), .B(n49517), .X(n25275) );
  nand_x1_sg U64791 ( .A(n25277), .B(n25276), .X(n25274) );
  inv_x1_sg U64792 ( .A(n25277), .X(n49540) );
  nand_x1_sg U64793 ( .A(n25556), .B(n25555), .X(n25553) );
  inv_x1_sg U64794 ( .A(n25556), .X(n49826) );
  nand_x1_sg U64795 ( .A(n50112), .B(n50089), .X(n25831) );
  nand_x1_sg U64796 ( .A(n25833), .B(n25832), .X(n25830) );
  inv_x1_sg U64797 ( .A(n25833), .X(n50112) );
  nand_x1_sg U64798 ( .A(n50397), .B(n50395), .X(n26064) );
  nand_x1_sg U64799 ( .A(n26065), .B(n26066), .X(n26063) );
  inv_x1_sg U64800 ( .A(n26065), .X(n50397) );
  nand_x1_sg U64801 ( .A(n50686), .B(n50663), .X(n26391) );
  nand_x1_sg U64802 ( .A(n26393), .B(n26392), .X(n26390) );
  inv_x1_sg U64803 ( .A(n26393), .X(n50686) );
  nand_x1_sg U64804 ( .A(n50973), .B(n50950), .X(n26669) );
  nand_x1_sg U64805 ( .A(n26671), .B(n26670), .X(n26668) );
  inv_x1_sg U64806 ( .A(n26671), .X(n50973) );
  nor_x1_sg U64807 ( .A(n39502), .B(n40367), .X(n7188) );
  nor_x1_sg U64808 ( .A(n39504), .B(n40312), .X(n17013) );
  nor_x1_sg U64809 ( .A(n39931), .B(n42369), .X(n7551) );
  nor_x1_sg U64810 ( .A(n40129), .B(n42337), .X(n17376) );
  nor_x1_sg U64811 ( .A(n41691), .B(n42369), .X(n7006) );
  nor_x1_sg U64812 ( .A(n41671), .B(n42337), .X(n16830) );
  nor_x1_sg U64813 ( .A(n40039), .B(n6834), .X(n7102) );
  nor_x1_sg U64814 ( .A(n40063), .B(n7651), .X(n7920) );
  nor_x1_sg U64815 ( .A(n40041), .B(n40556), .X(n8738) );
  nor_x1_sg U64816 ( .A(n9539), .B(n40552), .X(n9558) );
  nor_x1_sg U64817 ( .A(n40046), .B(n40548), .X(n10377) );
  nor_x1_sg U64818 ( .A(n42126), .B(n40545), .X(n11196) );
  nor_x1_sg U64819 ( .A(n40049), .B(n40539), .X(n12015) );
  nor_x1_sg U64820 ( .A(n40051), .B(n40535), .X(n12834) );
  nor_x1_sg U64821 ( .A(n40066), .B(n40531), .X(n13653) );
  nor_x1_sg U64822 ( .A(n42124), .B(n40528), .X(n14472) );
  nor_x1_sg U64823 ( .A(n42122), .B(n40524), .X(n15291) );
  nor_x1_sg U64824 ( .A(n40058), .B(n40521), .X(n16110) );
  nor_x1_sg U64825 ( .A(n17729), .B(n40517), .X(n17748) );
  nor_x1_sg U64826 ( .A(n40061), .B(n40511), .X(n18569) );
  nor_x1_sg U64827 ( .A(n42325), .B(n41809), .X(n7079) );
  nor_x1_sg U64828 ( .A(n40063), .B(n41937), .X(n7897) );
  nor_x1_sg U64829 ( .A(n40042), .B(n41940), .X(n8715) );
  nor_x1_sg U64830 ( .A(n9539), .B(n39972), .X(n9535) );
  nor_x1_sg U64831 ( .A(n10358), .B(n41936), .X(n10354) );
  nor_x1_sg U64832 ( .A(n42126), .B(n39980), .X(n11173) );
  nor_x1_sg U64833 ( .A(n40049), .B(n39983), .X(n11992) );
  nor_x1_sg U64834 ( .A(n12815), .B(n39989), .X(n12811) );
  nor_x1_sg U64835 ( .A(n13634), .B(n41922), .X(n13630) );
  nor_x1_sg U64836 ( .A(n40053), .B(n41921), .X(n14449) );
  nor_x1_sg U64837 ( .A(n42122), .B(n40000), .X(n15268) );
  nor_x1_sg U64838 ( .A(n40057), .B(n41942), .X(n16087) );
  nor_x1_sg U64839 ( .A(n40059), .B(n41001), .X(n17725) );
  nor_x1_sg U64840 ( .A(n18550), .B(n40008), .X(n18546) );
  nor_x1_sg U64841 ( .A(n6118), .B(n20294), .X(n20293) );
  nand_x1_sg U64842 ( .A(n20294), .B(n38699), .X(n20295) );
  nor_x1_sg U64843 ( .A(n42331), .B(n20123), .X(n20122) );
  nand_x1_sg U64844 ( .A(n20123), .B(n38640), .X(n20124) );
  nor_x1_sg U64845 ( .A(n42330), .B(n19923), .X(n19922) );
  nand_x1_sg U64846 ( .A(n19923), .B(n38636), .X(n19924) );
  nand_x1_sg U64847 ( .A(n46965), .B(n22761), .X(n22758) );
  inv_x1_sg U64848 ( .A(n22761), .X(n46985) );
  nand_x1_sg U64849 ( .A(n47007), .B(n22747), .X(n22744) );
  inv_x1_sg U64850 ( .A(n22747), .X(n47027) );
  nand_x1_sg U64851 ( .A(n47255), .B(n23038), .X(n23035) );
  inv_x1_sg U64852 ( .A(n23038), .X(n47274) );
  nand_x1_sg U64853 ( .A(n47540), .B(n23318), .X(n23315) );
  inv_x1_sg U64854 ( .A(n23318), .X(n47559) );
  nand_x1_sg U64855 ( .A(n47825), .B(n23597), .X(n23594) );
  inv_x1_sg U64856 ( .A(n23597), .X(n47844) );
  nand_x1_sg U64857 ( .A(n48110), .B(n23876), .X(n23873) );
  inv_x1_sg U64858 ( .A(n23876), .X(n48129) );
  nand_x1_sg U64859 ( .A(n48395), .B(n24155), .X(n24152) );
  inv_x1_sg U64860 ( .A(n24155), .X(n48414) );
  nand_x1_sg U64861 ( .A(n48680), .B(n24434), .X(n24431) );
  inv_x1_sg U64862 ( .A(n24434), .X(n48699) );
  nand_x1_sg U64863 ( .A(n48966), .B(n24712), .X(n24709) );
  inv_x1_sg U64864 ( .A(n24712), .X(n48985) );
  nand_x1_sg U64865 ( .A(n49253), .B(n24991), .X(n24988) );
  inv_x1_sg U64866 ( .A(n24991), .X(n49272) );
  nand_x1_sg U64867 ( .A(n49539), .B(n25270), .X(n25267) );
  inv_x1_sg U64868 ( .A(n25270), .X(n49558) );
  nand_x1_sg U64869 ( .A(n49825), .B(n25549), .X(n25546) );
  inv_x1_sg U64870 ( .A(n25549), .X(n49844) );
  nand_x1_sg U64871 ( .A(n50111), .B(n25826), .X(n25823) );
  inv_x1_sg U64872 ( .A(n25826), .X(n50130) );
  nand_x1_sg U64873 ( .A(n50685), .B(n26386), .X(n26383) );
  inv_x1_sg U64874 ( .A(n26386), .X(n50704) );
  nand_x1_sg U64875 ( .A(n50972), .B(n26664), .X(n26661) );
  inv_x1_sg U64876 ( .A(n26664), .X(n50991) );
  nor_x1_sg U64877 ( .A(n39681), .B(n40993), .X(n16906) );
  nor_x1_sg U64878 ( .A(n42147), .B(n26029), .X(n5747) );
  nor_x1_sg U64879 ( .A(n39548), .B(n39965), .X(n8025) );
  nor_x1_sg U64880 ( .A(n39549), .B(n41940), .X(n8843) );
  nor_x1_sg U64881 ( .A(n39550), .B(n41927), .X(n9663) );
  nor_x1_sg U64882 ( .A(n39557), .B(n41936), .X(n10482) );
  nor_x1_sg U64883 ( .A(n39558), .B(n41939), .X(n11301) );
  nor_x1_sg U64884 ( .A(n39554), .B(n41943), .X(n12120) );
  nor_x1_sg U64885 ( .A(n39555), .B(n41935), .X(n12939) );
  nor_x1_sg U64886 ( .A(n41728), .B(n41938), .X(n13758) );
  nor_x1_sg U64887 ( .A(n39553), .B(n39995), .X(n14577) );
  nor_x1_sg U64888 ( .A(n41733), .B(n41934), .X(n15396) );
  nor_x1_sg U64889 ( .A(n39552), .B(n41919), .X(n16215) );
  nor_x1_sg U64890 ( .A(n39545), .B(n40995), .X(n17031) );
  nor_x1_sg U64891 ( .A(n41738), .B(n41000), .X(n17853) );
  nor_x1_sg U64892 ( .A(n39547), .B(n41941), .X(n18674) );
  nor_x1_sg U64893 ( .A(n16820), .B(n40995), .X(n16665) );
  nand_x1_sg U64894 ( .A(n50453), .B(n26048), .X(n26045) );
  inv_x1_sg U64895 ( .A(n26048), .X(n50455) );
  nand_x1_sg U64896 ( .A(n50413), .B(n26060), .X(n26057) );
  inv_x1_sg U64897 ( .A(n26060), .X(n50415) );
  nor_x1_sg U64898 ( .A(n6996), .B(n41060), .X(n6841) );
  nor_x1_sg U64899 ( .A(n7813), .B(n39964), .X(n7658) );
  nor_x1_sg U64900 ( .A(n8631), .B(n39967), .X(n8476) );
  nor_x1_sg U64901 ( .A(n9451), .B(n41933), .X(n9296) );
  nor_x1_sg U64902 ( .A(n10270), .B(n41936), .X(n10115) );
  nor_x1_sg U64903 ( .A(n39308), .B(n39981), .X(n10934) );
  nor_x1_sg U64904 ( .A(n11908), .B(n39985), .X(n11753) );
  nor_x1_sg U64905 ( .A(n12727), .B(n41935), .X(n12572) );
  nor_x1_sg U64906 ( .A(n13546), .B(n41938), .X(n13391) );
  nor_x1_sg U64907 ( .A(n14365), .B(n39995), .X(n14210) );
  nor_x1_sg U64908 ( .A(n39298), .B(n41934), .X(n15029) );
  nor_x1_sg U64909 ( .A(n16003), .B(n40005), .X(n15848) );
  nor_x1_sg U64910 ( .A(n17641), .B(n40999), .X(n17486) );
  nor_x1_sg U64911 ( .A(n18462), .B(n41941), .X(n18307) );
  nor_x1_sg U64912 ( .A(n40039), .B(n39606), .X(n7552) );
  nor_x1_sg U64913 ( .A(n40064), .B(n39731), .X(n8370) );
  nor_x1_sg U64914 ( .A(n40042), .B(n39734), .X(n9188) );
  nor_x1_sg U64915 ( .A(n9539), .B(n39737), .X(n10008) );
  nor_x1_sg U64916 ( .A(n40045), .B(n39739), .X(n10827) );
  nor_x1_sg U64917 ( .A(n40048), .B(n39743), .X(n11646) );
  nor_x1_sg U64918 ( .A(n40050), .B(n39746), .X(n12465) );
  nor_x1_sg U64919 ( .A(n40052), .B(n39749), .X(n13284) );
  nor_x1_sg U64920 ( .A(n13634), .B(n39752), .X(n14103) );
  nor_x1_sg U64921 ( .A(n42124), .B(n39754), .X(n14922) );
  nor_x1_sg U64922 ( .A(n40056), .B(n39758), .X(n15741) );
  nor_x1_sg U64923 ( .A(n16091), .B(n39761), .X(n16560) );
  nor_x1_sg U64924 ( .A(n40059), .B(n39763), .X(n18198) );
  nor_x1_sg U64925 ( .A(n18550), .B(n41658), .X(n19019) );
  nand_x1_sg U64926 ( .A(n47056), .B(n22733), .X(n22730) );
  inv_x1_sg U64927 ( .A(n22733), .X(n47075) );
  nand_x1_sg U64928 ( .A(n47342), .B(n23010), .X(n23007) );
  inv_x1_sg U64929 ( .A(n23010), .X(n47361) );
  nand_x1_sg U64930 ( .A(n47627), .B(n23290), .X(n23287) );
  inv_x1_sg U64931 ( .A(n23290), .X(n47646) );
  nand_x1_sg U64932 ( .A(n47912), .B(n23569), .X(n23566) );
  inv_x1_sg U64933 ( .A(n23569), .X(n47931) );
  nand_x1_sg U64934 ( .A(n48197), .B(n23848), .X(n23845) );
  inv_x1_sg U64935 ( .A(n23848), .X(n48216) );
  nand_x1_sg U64936 ( .A(n48482), .B(n24127), .X(n24124) );
  inv_x1_sg U64937 ( .A(n24127), .X(n48501) );
  nand_x1_sg U64938 ( .A(n48767), .B(n24406), .X(n24403) );
  inv_x1_sg U64939 ( .A(n24406), .X(n48786) );
  nand_x1_sg U64940 ( .A(n49053), .B(n24684), .X(n24681) );
  inv_x1_sg U64941 ( .A(n24684), .X(n49073) );
  nand_x1_sg U64942 ( .A(n49340), .B(n24963), .X(n24960) );
  inv_x1_sg U64943 ( .A(n24963), .X(n49359) );
  nand_x1_sg U64944 ( .A(n49626), .B(n25242), .X(n25239) );
  inv_x1_sg U64945 ( .A(n25242), .X(n49645) );
  nand_x1_sg U64946 ( .A(n49912), .B(n25521), .X(n25518) );
  inv_x1_sg U64947 ( .A(n25521), .X(n49931) );
  nand_x1_sg U64948 ( .A(n50198), .B(n25798), .X(n25795) );
  inv_x1_sg U64949 ( .A(n25798), .X(n50217) );
  nand_x1_sg U64950 ( .A(n50772), .B(n26358), .X(n26355) );
  inv_x1_sg U64951 ( .A(n26358), .X(n50791) );
  nand_x1_sg U64952 ( .A(n51059), .B(n26636), .X(n26633) );
  inv_x1_sg U64953 ( .A(n26636), .X(n51078) );
  nor_x1_sg U64954 ( .A(n39612), .B(n41937), .X(n8102) );
  nor_x1_sg U64955 ( .A(n39608), .B(n39968), .X(n8920) );
  nor_x1_sg U64956 ( .A(n39627), .B(n41933), .X(n9740) );
  nor_x1_sg U64957 ( .A(n39624), .B(n39976), .X(n10559) );
  nor_x1_sg U64958 ( .A(n39621), .B(n39979), .X(n11378) );
  nor_x1_sg U64959 ( .A(n39618), .B(n40710), .X(n12197) );
  nor_x1_sg U64960 ( .A(n39639), .B(n39987), .X(n13016) );
  nor_x1_sg U64961 ( .A(n39636), .B(n41938), .X(n13835) );
  nor_x1_sg U64962 ( .A(n39633), .B(n39996), .X(n14654) );
  nor_x1_sg U64963 ( .A(n39630), .B(n40730), .X(n15473) );
  nor_x1_sg U64964 ( .A(n39648), .B(n41942), .X(n16292) );
  nor_x1_sg U64965 ( .A(n39615), .B(n40996), .X(n17108) );
  nor_x1_sg U64966 ( .A(n39645), .B(n40998), .X(n17930) );
  nor_x1_sg U64967 ( .A(n39642), .B(n40007), .X(n18751) );
  nor_x1_sg U64968 ( .A(n39725), .B(n38913), .X(n7206) );
  nor_x1_sg U64969 ( .A(n46876), .B(n40573), .X(n22628) );
  nor_x1_sg U64970 ( .A(n47169), .B(n40633), .X(n22894) );
  nor_x1_sg U64971 ( .A(n47454), .B(n40628), .X(n23171) );
  nor_x1_sg U64972 ( .A(n47739), .B(n40667), .X(n23451) );
  nor_x1_sg U64973 ( .A(n48024), .B(n40657), .X(n23730) );
  nor_x1_sg U64974 ( .A(n48309), .B(n40644), .X(n24009) );
  nor_x1_sg U64975 ( .A(n48594), .B(n40639), .X(n24288) );
  nor_x1_sg U64976 ( .A(n48880), .B(n40662), .X(n24567) );
  nor_x1_sg U64977 ( .A(n49167), .B(n40652), .X(n24845) );
  nor_x1_sg U64978 ( .A(n49453), .B(n40622), .X(n25124) );
  nor_x1_sg U64979 ( .A(n49738), .B(n40684), .X(n25403) );
  nor_x1_sg U64980 ( .A(n50025), .B(n40678), .X(n25682) );
  nor_x1_sg U64981 ( .A(n50302), .B(n40579), .X(n25951) );
  nor_x1_sg U64982 ( .A(n50599), .B(n40646), .X(n26228) );
  nor_x1_sg U64983 ( .A(n50886), .B(n40673), .X(n26519) );
  nor_x1_sg U64984 ( .A(n39771), .B(n40312), .X(n16956) );
  nor_x1_sg U64985 ( .A(n41725), .B(n41059), .X(n7283) );
  nand_x1_sg U64986 ( .A(n40563), .B(n42092), .X(n16820) );
  nand_x1_sg U64987 ( .A(n40242), .B(n42105), .X(n7813) );
  nand_x1_sg U64988 ( .A(n40250), .B(n40361), .X(n8631) );
  nand_x1_sg U64989 ( .A(n40252), .B(n40355), .X(n9451) );
  nand_x1_sg U64990 ( .A(n40258), .B(n40351), .X(n10270) );
  nand_x1_sg U64991 ( .A(n40263), .B(n40347), .X(n11089) );
  nand_x1_sg U64992 ( .A(n40267), .B(n40327), .X(n11908) );
  nand_x1_sg U64993 ( .A(n40273), .B(n40339), .X(n12727) );
  nand_x1_sg U64994 ( .A(n40280), .B(n40335), .X(n13546) );
  nand_x1_sg U64995 ( .A(n40285), .B(n40343), .X(n14365) );
  nand_x1_sg U64996 ( .A(n40288), .B(n40319), .X(n15184) );
  nand_x1_sg U64997 ( .A(n40293), .B(n40323), .X(n16003) );
  nand_x1_sg U64998 ( .A(n40297), .B(n40331), .X(n18462) );
  nand_x1_sg U64999 ( .A(n40239), .B(n42091), .X(n17641) );
  nand_x1_sg U65000 ( .A(n40163), .B(n39957), .X(n6996) );
  nand_x1_sg U65001 ( .A(n39435), .B(n18286), .X(n18285) );
  nand_x1_sg U65002 ( .A(n50373), .B(n26072), .X(n26069) );
  inv_x1_sg U65003 ( .A(n26072), .X(n50375) );
  nand_x1_sg U65004 ( .A(n47216), .B(n23052), .X(n23049) );
  inv_x1_sg U65005 ( .A(n23052), .X(n47234) );
  inv_x1_sg U65006 ( .A(n23024), .X(n47314) );
  nand_x1_sg U65007 ( .A(n47501), .B(n23332), .X(n23329) );
  inv_x1_sg U65008 ( .A(n23332), .X(n47519) );
  inv_x1_sg U65009 ( .A(n23304), .X(n47599) );
  nand_x1_sg U65010 ( .A(n47786), .B(n23611), .X(n23608) );
  inv_x1_sg U65011 ( .A(n23611), .X(n47804) );
  inv_x1_sg U65012 ( .A(n23583), .X(n47884) );
  nand_x1_sg U65013 ( .A(n48071), .B(n23890), .X(n23887) );
  inv_x1_sg U65014 ( .A(n23890), .X(n48089) );
  inv_x1_sg U65015 ( .A(n23862), .X(n48169) );
  nand_x1_sg U65016 ( .A(n48356), .B(n24169), .X(n24166) );
  inv_x1_sg U65017 ( .A(n24169), .X(n48374) );
  inv_x1_sg U65018 ( .A(n24141), .X(n48454) );
  nand_x1_sg U65019 ( .A(n48641), .B(n24448), .X(n24445) );
  inv_x1_sg U65020 ( .A(n24448), .X(n48659) );
  inv_x1_sg U65021 ( .A(n24420), .X(n48739) );
  nand_x1_sg U65022 ( .A(n48927), .B(n24726), .X(n24723) );
  inv_x1_sg U65023 ( .A(n24726), .X(n48945) );
  inv_x1_sg U65024 ( .A(n24698), .X(n49025) );
  nand_x1_sg U65025 ( .A(n49214), .B(n25005), .X(n25002) );
  inv_x1_sg U65026 ( .A(n25005), .X(n49232) );
  inv_x1_sg U65027 ( .A(n24977), .X(n49312) );
  nand_x1_sg U65028 ( .A(n49500), .B(n25284), .X(n25281) );
  inv_x1_sg U65029 ( .A(n25284), .X(n49518) );
  inv_x1_sg U65030 ( .A(n25256), .X(n49598) );
  nand_x1_sg U65031 ( .A(n49786), .B(n25563), .X(n25560) );
  inv_x1_sg U65032 ( .A(n25563), .X(n49804) );
  inv_x1_sg U65033 ( .A(n25535), .X(n49884) );
  nand_x1_sg U65034 ( .A(n50072), .B(n25840), .X(n25837) );
  inv_x1_sg U65035 ( .A(n25840), .X(n50090) );
  inv_x1_sg U65036 ( .A(n25812), .X(n50170) );
  nand_x1_sg U65037 ( .A(n50646), .B(n26400), .X(n26397) );
  inv_x1_sg U65038 ( .A(n26400), .X(n50664) );
  inv_x1_sg U65039 ( .A(n26372), .X(n50744) );
  nand_x1_sg U65040 ( .A(n50933), .B(n26678), .X(n26675) );
  inv_x1_sg U65041 ( .A(n26678), .X(n50951) );
  inv_x1_sg U65042 ( .A(n26650), .X(n51031) );
  nand_x1_sg U65043 ( .A(n47057), .B(n47026), .X(n22738) );
  nand_x1_sg U65044 ( .A(n22740), .B(n22739), .X(n22737) );
  inv_x1_sg U65045 ( .A(n22740), .X(n47057) );
  nand_x1_sg U65046 ( .A(n47343), .B(n47313), .X(n23015) );
  nand_x1_sg U65047 ( .A(n23017), .B(n23016), .X(n23014) );
  inv_x1_sg U65048 ( .A(n23017), .X(n47343) );
  nand_x1_sg U65049 ( .A(n47628), .B(n47598), .X(n23295) );
  nand_x1_sg U65050 ( .A(n23297), .B(n23296), .X(n23294) );
  inv_x1_sg U65051 ( .A(n23297), .X(n47628) );
  nand_x1_sg U65052 ( .A(n47913), .B(n47883), .X(n23574) );
  nand_x1_sg U65053 ( .A(n23576), .B(n23575), .X(n23573) );
  inv_x1_sg U65054 ( .A(n23576), .X(n47913) );
  nand_x1_sg U65055 ( .A(n48198), .B(n48168), .X(n23853) );
  nand_x1_sg U65056 ( .A(n23855), .B(n23854), .X(n23852) );
  inv_x1_sg U65057 ( .A(n23855), .X(n48198) );
  nand_x1_sg U65058 ( .A(n48483), .B(n48453), .X(n24132) );
  nand_x1_sg U65059 ( .A(n24134), .B(n24133), .X(n24131) );
  inv_x1_sg U65060 ( .A(n24134), .X(n48483) );
  nand_x1_sg U65061 ( .A(n48768), .B(n48738), .X(n24411) );
  nand_x1_sg U65062 ( .A(n24413), .B(n24412), .X(n24410) );
  inv_x1_sg U65063 ( .A(n24413), .X(n48768) );
  nand_x1_sg U65064 ( .A(n49054), .B(n49024), .X(n24689) );
  nand_x1_sg U65065 ( .A(n24691), .B(n24690), .X(n24688) );
  inv_x1_sg U65066 ( .A(n24691), .X(n49054) );
  nand_x1_sg U65067 ( .A(n49341), .B(n49311), .X(n24968) );
  nand_x1_sg U65068 ( .A(n24970), .B(n24969), .X(n24967) );
  inv_x1_sg U65069 ( .A(n24970), .X(n49341) );
  nand_x1_sg U65070 ( .A(n49627), .B(n49597), .X(n25247) );
  nand_x1_sg U65071 ( .A(n25249), .B(n25248), .X(n25246) );
  inv_x1_sg U65072 ( .A(n25249), .X(n49627) );
  nand_x1_sg U65073 ( .A(n49913), .B(n49883), .X(n25526) );
  nand_x1_sg U65074 ( .A(n25528), .B(n25527), .X(n25525) );
  inv_x1_sg U65075 ( .A(n25528), .X(n49913) );
  nand_x1_sg U65076 ( .A(n50199), .B(n50169), .X(n25803) );
  nand_x1_sg U65077 ( .A(n25805), .B(n25804), .X(n25802) );
  inv_x1_sg U65078 ( .A(n25805), .X(n50199) );
  nand_x1_sg U65079 ( .A(n50484), .B(n50482), .X(n26040) );
  nand_x1_sg U65080 ( .A(n26041), .B(n26042), .X(n26039) );
  inv_x1_sg U65081 ( .A(n26041), .X(n50484) );
  nand_x1_sg U65082 ( .A(n50773), .B(n50743), .X(n26363) );
  nand_x1_sg U65083 ( .A(n26365), .B(n26364), .X(n26362) );
  inv_x1_sg U65084 ( .A(n26365), .X(n50773) );
  nand_x1_sg U65085 ( .A(n51060), .B(n51030), .X(n26641) );
  nand_x1_sg U65086 ( .A(n26643), .B(n26642), .X(n26640) );
  inv_x1_sg U65087 ( .A(n26643), .X(n51060) );
  nand_x1_sg U65088 ( .A(n47184), .B(n23066), .X(n23065) );
  nand_x1_sg U65089 ( .A(n47197), .B(n23063), .X(n23064) );
  nand_x1_sg U65090 ( .A(n47469), .B(n23346), .X(n23345) );
  nand_x1_sg U65091 ( .A(n47482), .B(n23343), .X(n23344) );
  nand_x1_sg U65092 ( .A(n47754), .B(n23625), .X(n23624) );
  nand_x1_sg U65093 ( .A(n47767), .B(n23622), .X(n23623) );
  nand_x1_sg U65094 ( .A(n48039), .B(n23904), .X(n23903) );
  nand_x1_sg U65095 ( .A(n48052), .B(n23901), .X(n23902) );
  nand_x1_sg U65096 ( .A(n48324), .B(n24183), .X(n24182) );
  nand_x1_sg U65097 ( .A(n48337), .B(n24180), .X(n24181) );
  nand_x1_sg U65098 ( .A(n48609), .B(n24462), .X(n24461) );
  nand_x1_sg U65099 ( .A(n48622), .B(n24459), .X(n24460) );
  nand_x1_sg U65100 ( .A(n48895), .B(n24740), .X(n24739) );
  nand_x1_sg U65101 ( .A(n48908), .B(n24737), .X(n24738) );
  nand_x1_sg U65102 ( .A(n49182), .B(n25019), .X(n25018) );
  nand_x1_sg U65103 ( .A(n49195), .B(n25016), .X(n25017) );
  nand_x1_sg U65104 ( .A(n49468), .B(n25298), .X(n25297) );
  nand_x1_sg U65105 ( .A(n49481), .B(n25295), .X(n25296) );
  nand_x1_sg U65106 ( .A(n49753), .B(n25577), .X(n25576) );
  nand_x1_sg U65107 ( .A(n49767), .B(n25574), .X(n25575) );
  nand_x1_sg U65108 ( .A(n50040), .B(n25854), .X(n25853) );
  nand_x1_sg U65109 ( .A(n50053), .B(n25851), .X(n25852) );
  nand_x1_sg U65110 ( .A(n50336), .B(n26083), .X(n26082) );
  nand_x1_sg U65111 ( .A(n50338), .B(n26084), .X(n26081) );
  nand_x1_sg U65112 ( .A(n50614), .B(n26414), .X(n26413) );
  nand_x1_sg U65113 ( .A(n50627), .B(n26411), .X(n26412) );
  nand_x1_sg U65114 ( .A(n50901), .B(n26692), .X(n26691) );
  nand_x1_sg U65115 ( .A(n50914), .B(n26689), .X(n26690) );
  nand_x1_sg U65116 ( .A(n40221), .B(n51138), .X(n15008) );
  nand_x1_sg U65117 ( .A(n40089), .B(n51140), .X(n14189) );
  nand_x1_sg U65118 ( .A(n46904), .B(n22786), .X(n22787) );
  nand_x1_sg U65119 ( .A(n38984), .B(n51137), .X(n10094) );
  nor_x1_sg U65120 ( .A(n17104), .B(n40129), .X(n17103) );
  nor_x1_sg U65121 ( .A(n16786), .B(n50286), .X(n17102) );
  nand_x1_sg U65122 ( .A(n17077), .B(n40564), .X(n17104) );
  nor_x1_sg U65123 ( .A(n50277), .B(n40564), .X(n25927) );
  nor_x1_sg U65124 ( .A(n46853), .B(n7111), .X(n22616) );
  nor_x1_sg U65125 ( .A(n46866), .B(n41781), .X(n22622) );
  nor_x1_sg U65126 ( .A(n47146), .B(n39065), .X(n22880) );
  nor_x1_sg U65127 ( .A(n47159), .B(n41783), .X(n22887) );
  nor_x1_sg U65128 ( .A(n47431), .B(n39064), .X(n23157) );
  nor_x1_sg U65129 ( .A(n47444), .B(n41785), .X(n23164) );
  nor_x1_sg U65130 ( .A(n47716), .B(n39063), .X(n23437) );
  nor_x1_sg U65131 ( .A(n47729), .B(n41787), .X(n23444) );
  nor_x1_sg U65132 ( .A(n48001), .B(n39062), .X(n23716) );
  nor_x1_sg U65133 ( .A(n48014), .B(n41789), .X(n23723) );
  nor_x1_sg U65134 ( .A(n48286), .B(n39061), .X(n23995) );
  nor_x1_sg U65135 ( .A(n48299), .B(n11188), .X(n24002) );
  nor_x1_sg U65136 ( .A(n48571), .B(n39060), .X(n24274) );
  nor_x1_sg U65137 ( .A(n48584), .B(n12007), .X(n24281) );
  nor_x1_sg U65138 ( .A(n48857), .B(n39059), .X(n24553) );
  nor_x1_sg U65139 ( .A(n48870), .B(n41795), .X(n24560) );
  nor_x1_sg U65140 ( .A(n49144), .B(n39058), .X(n24831) );
  nor_x1_sg U65141 ( .A(n49157), .B(n13645), .X(n24838) );
  nor_x1_sg U65142 ( .A(n49430), .B(n39057), .X(n25110) );
  nor_x1_sg U65143 ( .A(n49443), .B(n41799), .X(n25117) );
  nor_x1_sg U65144 ( .A(n49715), .B(n39056), .X(n25389) );
  nor_x1_sg U65145 ( .A(n49728), .B(n15283), .X(n25396) );
  nor_x1_sg U65146 ( .A(n50002), .B(n39055), .X(n25668) );
  nor_x1_sg U65147 ( .A(n50015), .B(n41803), .X(n25675) );
  nor_x1_sg U65148 ( .A(n50289), .B(n16936), .X(n25939) );
  nor_x1_sg U65149 ( .A(n50576), .B(n39053), .X(n26212) );
  nor_x1_sg U65150 ( .A(n50589), .B(n17740), .X(n26220) );
  nor_x1_sg U65151 ( .A(n50863), .B(n39054), .X(n26505) );
  nor_x1_sg U65152 ( .A(n50876), .B(n41807), .X(n26512) );
  nand_x1_sg U65153 ( .A(n23258), .B(n41316), .X(n23251) );
  nand_x1_sg U65154 ( .A(n23253), .B(n47703), .X(n23252) );
  nand_x1_sg U65155 ( .A(n23255), .B(n40505), .X(n23258) );
  nor_x1_sg U65156 ( .A(n39722), .B(n41060), .X(n7097) );
  nor_x1_sg U65157 ( .A(n39719), .B(n41929), .X(n7915) );
  nor_x1_sg U65158 ( .A(n39716), .B(n40690), .X(n8733) );
  nor_x1_sg U65159 ( .A(n41786), .B(n39972), .X(n9553) );
  nor_x1_sg U65160 ( .A(n39710), .B(n39975), .X(n10372) );
  nor_x1_sg U65161 ( .A(n39707), .B(n41939), .X(n11191) );
  nor_x1_sg U65162 ( .A(n41792), .B(n39985), .X(n12010) );
  nor_x1_sg U65163 ( .A(n41794), .B(n41935), .X(n12829) );
  nor_x1_sg U65164 ( .A(n41796), .B(n39992), .X(n13648) );
  nor_x1_sg U65165 ( .A(n39695), .B(n41921), .X(n14467) );
  nor_x1_sg U65166 ( .A(n41800), .B(n40001), .X(n15286) );
  nor_x1_sg U65167 ( .A(n41802), .B(n40003), .X(n16105) );
  nor_x1_sg U65168 ( .A(n41804), .B(n41001), .X(n17743) );
  nor_x1_sg U65169 ( .A(n41806), .B(n40009), .X(n18564) );
  nor_x1_sg U65170 ( .A(n40040), .B(n39038), .X(n7625) );
  nor_x1_sg U65171 ( .A(n42089), .B(n39040), .X(n8443) );
  nor_x1_sg U65172 ( .A(n40042), .B(n39039), .X(n9261) );
  nor_x1_sg U65173 ( .A(n40044), .B(n39042), .X(n10081) );
  nor_x1_sg U65174 ( .A(n40045), .B(n39041), .X(n10900) );
  nor_x1_sg U65175 ( .A(n42126), .B(n39044), .X(n11719) );
  nor_x1_sg U65176 ( .A(n40050), .B(n39043), .X(n12538) );
  nor_x1_sg U65177 ( .A(n40052), .B(n39046), .X(n13357) );
  nor_x1_sg U65178 ( .A(n40065), .B(n39045), .X(n14176) );
  nor_x1_sg U65179 ( .A(n42124), .B(n39048), .X(n14995) );
  nor_x1_sg U65180 ( .A(n40056), .B(n39047), .X(n15814) );
  nor_x1_sg U65181 ( .A(n40057), .B(n39050), .X(n16633) );
  nor_x1_sg U65182 ( .A(n17729), .B(n39049), .X(n18271) );
  nor_x1_sg U65183 ( .A(n40062), .B(n39051), .X(n19092) );
  nand_x1_sg U65184 ( .A(n41283), .B(n40456), .X(n42378) );
  nor_x1_sg U65185 ( .A(n39810), .B(n46871), .X(n7081) );
  nor_x1_sg U65186 ( .A(n7082), .B(n40040), .X(n7080) );
  nor_x1_sg U65187 ( .A(n39812), .B(n47164), .X(n7899) );
  nor_x1_sg U65188 ( .A(n7900), .B(n40064), .X(n7898) );
  nor_x1_sg U65189 ( .A(n39831), .B(n47449), .X(n8717) );
  nor_x1_sg U65190 ( .A(n8718), .B(n42130), .X(n8716) );
  nor_x1_sg U65191 ( .A(n39845), .B(n47734), .X(n9537) );
  nor_x1_sg U65192 ( .A(n9538), .B(n40044), .X(n9536) );
  nor_x1_sg U65193 ( .A(n39816), .B(n48019), .X(n10356) );
  nor_x1_sg U65194 ( .A(n10357), .B(n10358), .X(n10355) );
  nor_x1_sg U65195 ( .A(n39834), .B(n48304), .X(n11175) );
  nor_x1_sg U65196 ( .A(n11176), .B(n40047), .X(n11174) );
  nor_x1_sg U65197 ( .A(n39837), .B(n48589), .X(n11994) );
  nor_x1_sg U65198 ( .A(n11995), .B(n40050), .X(n11993) );
  nor_x1_sg U65199 ( .A(n39819), .B(n48875), .X(n12813) );
  nor_x1_sg U65200 ( .A(n12814), .B(n12815), .X(n12812) );
  nor_x1_sg U65201 ( .A(n39839), .B(n49162), .X(n13632) );
  nor_x1_sg U65202 ( .A(n13633), .B(n13634), .X(n13631) );
  nor_x1_sg U65203 ( .A(n39842), .B(n49448), .X(n14451) );
  nor_x1_sg U65204 ( .A(n14452), .B(n40054), .X(n14450) );
  nor_x1_sg U65205 ( .A(n41876), .B(n49733), .X(n15270) );
  nor_x1_sg U65206 ( .A(n15271), .B(n40055), .X(n15269) );
  nor_x1_sg U65207 ( .A(n39821), .B(n50020), .X(n16089) );
  nor_x1_sg U65208 ( .A(n16090), .B(n40058), .X(n16088) );
  nor_x1_sg U65209 ( .A(n39828), .B(n50594), .X(n17727) );
  nor_x1_sg U65210 ( .A(n17728), .B(n17729), .X(n17726) );
  nor_x1_sg U65211 ( .A(n39825), .B(n50881), .X(n18548) );
  nor_x1_sg U65212 ( .A(n18549), .B(n18550), .X(n18547) );
  nor_x1_sg U65213 ( .A(n39771), .B(n39602), .X(n17411) );
  nor_x1_sg U65214 ( .A(n39771), .B(n41671), .X(n17429) );
  nor_x1_sg U65215 ( .A(n39770), .B(n39052), .X(n16846) );
  nor_x1_sg U65216 ( .A(n39770), .B(n38908), .X(n16922) );
  nor_x1_sg U65217 ( .A(n8035), .B(n40064), .X(n8105) );
  nor_x1_sg U65218 ( .A(n8853), .B(n40041), .X(n8923) );
  nor_x1_sg U65219 ( .A(n40110), .B(n40043), .X(n9743) );
  nor_x1_sg U65220 ( .A(n40111), .B(n10358), .X(n10562) );
  nor_x1_sg U65221 ( .A(n11311), .B(n40048), .X(n11381) );
  nor_x1_sg U65222 ( .A(n40116), .B(n11996), .X(n12200) );
  nor_x1_sg U65223 ( .A(n40117), .B(n40052), .X(n13019) );
  nor_x1_sg U65224 ( .A(n13768), .B(n40066), .X(n13838) );
  nor_x1_sg U65225 ( .A(n40122), .B(n40054), .X(n14657) );
  nor_x1_sg U65226 ( .A(n40124), .B(n40055), .X(n15476) );
  nor_x1_sg U65227 ( .A(n16225), .B(n16091), .X(n16295) );
  nor_x1_sg U65228 ( .A(n17863), .B(n40060), .X(n17933) );
  nor_x1_sg U65229 ( .A(n40128), .B(n40062), .X(n18754) );
  nor_x1_sg U65230 ( .A(n42163), .B(n40039), .X(n7287) );
  nor_x1_sg U65231 ( .A(n40085), .B(n41058), .X(n7074) );
  nor_x1_sg U65232 ( .A(n40088), .B(n40995), .X(n16901) );
  nand_x1_sg U65233 ( .A(n17465), .B(n39279), .X(n26140) );
  nor_x1_sg U65234 ( .A(n41750), .B(n39963), .X(n7892) );
  nor_x1_sg U65235 ( .A(n41742), .B(n41940), .X(n8710) );
  nor_x1_sg U65236 ( .A(n41743), .B(n39972), .X(n9530) );
  nor_x1_sg U65237 ( .A(n41744), .B(n39977), .X(n10349) );
  nor_x1_sg U65238 ( .A(n41745), .B(n41925), .X(n11168) );
  nor_x1_sg U65239 ( .A(n41746), .B(n41943), .X(n11987) );
  nor_x1_sg U65240 ( .A(n40191), .B(n40715), .X(n12806) );
  nor_x1_sg U65241 ( .A(n41751), .B(n39991), .X(n13625) );
  nor_x1_sg U65242 ( .A(n40187), .B(n41932), .X(n14444) );
  nor_x1_sg U65243 ( .A(n41752), .B(n41934), .X(n15263) );
  nor_x1_sg U65244 ( .A(n40166), .B(n41942), .X(n16082) );
  nor_x1_sg U65245 ( .A(n41741), .B(n40999), .X(n17720) );
  nor_x1_sg U65246 ( .A(n41749), .B(n41941), .X(n18541) );
  nand_x1_sg U65247 ( .A(n25951), .B(n39504), .X(n25958) );
  nor_x1_sg U65248 ( .A(n7004), .B(n47121), .X(n6983) );
  nor_x1_sg U65249 ( .A(n42045), .B(n7006), .X(n7004) );
  nand_x1_sg U65250 ( .A(n7006), .B(n7007), .X(n7005) );
  nor_x1_sg U65251 ( .A(n16828), .B(n50549), .X(n16807) );
  nor_x1_sg U65252 ( .A(n16831), .B(n16830), .X(n16828) );
  nand_x1_sg U65253 ( .A(n16830), .B(n16831), .X(n16829) );
  nor_x1_sg U65254 ( .A(n7821), .B(n47407), .X(n7800) );
  nor_x1_sg U65255 ( .A(n7824), .B(n7823), .X(n7821) );
  nand_x1_sg U65256 ( .A(n7823), .B(n7824), .X(n7822) );
  nor_x1_sg U65257 ( .A(n8639), .B(n47692), .X(n8618) );
  nor_x1_sg U65258 ( .A(n8642), .B(n8641), .X(n8639) );
  nand_x1_sg U65259 ( .A(n8641), .B(n8642), .X(n8640) );
  nor_x1_sg U65260 ( .A(n9459), .B(n47977), .X(n9438) );
  nor_x1_sg U65261 ( .A(n9462), .B(n9461), .X(n9459) );
  nand_x1_sg U65262 ( .A(n9461), .B(n9462), .X(n9460) );
  nor_x1_sg U65263 ( .A(n10278), .B(n48262), .X(n10257) );
  nor_x1_sg U65264 ( .A(n10281), .B(n10280), .X(n10278) );
  nand_x1_sg U65265 ( .A(n10280), .B(n10281), .X(n10279) );
  nor_x1_sg U65266 ( .A(n11097), .B(n48547), .X(n11076) );
  nor_x1_sg U65267 ( .A(n11100), .B(n11099), .X(n11097) );
  nand_x1_sg U65268 ( .A(n11099), .B(n11100), .X(n11098) );
  nor_x1_sg U65269 ( .A(n11916), .B(n48832), .X(n11895) );
  nor_x1_sg U65270 ( .A(n11919), .B(n11918), .X(n11916) );
  nand_x1_sg U65271 ( .A(n11918), .B(n11919), .X(n11917) );
  nor_x1_sg U65272 ( .A(n12735), .B(n49119), .X(n12714) );
  nor_x1_sg U65273 ( .A(n12738), .B(n12737), .X(n12735) );
  nand_x1_sg U65274 ( .A(n12737), .B(n12738), .X(n12736) );
  nor_x1_sg U65275 ( .A(n13554), .B(n49405), .X(n13533) );
  nor_x1_sg U65276 ( .A(n13557), .B(n13556), .X(n13554) );
  nand_x1_sg U65277 ( .A(n13556), .B(n13557), .X(n13555) );
  nor_x1_sg U65278 ( .A(n14373), .B(n49691), .X(n14352) );
  nor_x1_sg U65279 ( .A(n14376), .B(n14375), .X(n14373) );
  nand_x1_sg U65280 ( .A(n14375), .B(n14376), .X(n14374) );
  nor_x1_sg U65281 ( .A(n15192), .B(n49977), .X(n15171) );
  nor_x1_sg U65282 ( .A(n15195), .B(n15194), .X(n15192) );
  nand_x1_sg U65283 ( .A(n15194), .B(n15195), .X(n15193) );
  nor_x1_sg U65284 ( .A(n16011), .B(n50263), .X(n15990) );
  nor_x1_sg U65285 ( .A(n16014), .B(n16013), .X(n16011) );
  nand_x1_sg U65286 ( .A(n16013), .B(n16014), .X(n16012) );
  nor_x1_sg U65287 ( .A(n17649), .B(n50837), .X(n17628) );
  nor_x1_sg U65288 ( .A(n17652), .B(n17651), .X(n17649) );
  nand_x1_sg U65289 ( .A(n17651), .B(n17652), .X(n17650) );
  nor_x1_sg U65290 ( .A(n18470), .B(n51124), .X(n18449) );
  nor_x1_sg U65291 ( .A(n18473), .B(n18472), .X(n18470) );
  nand_x1_sg U65292 ( .A(n18472), .B(n18473), .X(n18471) );
  inv_x1_sg U65293 ( .A(n40068), .X(n50565) );
  nand_x1_sg U65294 ( .A(n25961), .B(n39280), .X(n25956) );
  nand_x1_sg U65295 ( .A(n25958), .B(n25959), .X(n25957) );
  nand_x1_sg U65296 ( .A(n40038), .B(n39504), .X(n25961) );
  nand_x1_sg U65297 ( .A(n25978), .B(n25979), .X(n25977) );
  nand_x1_sg U65298 ( .A(n40037), .B(n39615), .X(n25981) );
  nand_x1_sg U65299 ( .A(n22628), .B(n39502), .X(n22635) );
  nand_x1_sg U65300 ( .A(n22782), .B(n22781), .X(n22779) );
  inv_x1_sg U65301 ( .A(n22782), .X(n46925) );
  nand_x1_sg U65302 ( .A(n39519), .B(n40134), .X(n7779) );
  nand_x1_sg U65303 ( .A(n39518), .B(n42183), .X(n8597) );
  nand_x1_sg U65304 ( .A(n39524), .B(n42181), .X(n9417) );
  nand_x1_sg U65305 ( .A(n39523), .B(n42179), .X(n10236) );
  nand_x1_sg U65306 ( .A(n39522), .B(n42177), .X(n11055) );
  nand_x1_sg U65307 ( .A(n39521), .B(n42175), .X(n11874) );
  nand_x1_sg U65308 ( .A(n39528), .B(n42173), .X(n12693) );
  nand_x1_sg U65309 ( .A(n39527), .B(n42171), .X(n13512) );
  nand_x1_sg U65310 ( .A(n39526), .B(n42169), .X(n14331) );
  nand_x1_sg U65311 ( .A(n39525), .B(n40152), .X(n15150) );
  nand_x1_sg U65312 ( .A(n39531), .B(n42166), .X(n15969) );
  nand_x1_sg U65313 ( .A(n39530), .B(n17800), .X(n17607) );
  nand_x1_sg U65314 ( .A(n39529), .B(n40156), .X(n18428) );
  nand_x1_sg U65315 ( .A(n23059), .B(n23058), .X(n23056) );
  inv_x1_sg U65316 ( .A(n23059), .X(n47217) );
  nand_x1_sg U65317 ( .A(n23339), .B(n23338), .X(n23336) );
  inv_x1_sg U65318 ( .A(n23339), .X(n47502) );
  nand_x1_sg U65319 ( .A(n23618), .B(n23617), .X(n23615) );
  inv_x1_sg U65320 ( .A(n23618), .X(n47787) );
  nand_x1_sg U65321 ( .A(n23897), .B(n23896), .X(n23894) );
  inv_x1_sg U65322 ( .A(n23897), .X(n48072) );
  nand_x1_sg U65323 ( .A(n24176), .B(n24175), .X(n24173) );
  inv_x1_sg U65324 ( .A(n24176), .X(n48357) );
  nand_x1_sg U65325 ( .A(n24455), .B(n24454), .X(n24452) );
  inv_x1_sg U65326 ( .A(n24455), .X(n48642) );
  nand_x1_sg U65327 ( .A(n24733), .B(n24732), .X(n24730) );
  inv_x1_sg U65328 ( .A(n24733), .X(n48928) );
  nand_x1_sg U65329 ( .A(n25012), .B(n25011), .X(n25009) );
  inv_x1_sg U65330 ( .A(n25012), .X(n49215) );
  nand_x1_sg U65331 ( .A(n25291), .B(n25290), .X(n25288) );
  inv_x1_sg U65332 ( .A(n25291), .X(n49501) );
  nand_x1_sg U65333 ( .A(n25570), .B(n25569), .X(n25567) );
  inv_x1_sg U65334 ( .A(n25570), .X(n49787) );
  nand_x1_sg U65335 ( .A(n25847), .B(n25846), .X(n25844) );
  inv_x1_sg U65336 ( .A(n25847), .X(n50073) );
  nand_x1_sg U65337 ( .A(n26077), .B(n26078), .X(n26075) );
  inv_x1_sg U65338 ( .A(n26077), .X(n50358) );
  nand_x1_sg U65339 ( .A(n26407), .B(n26406), .X(n26404) );
  inv_x1_sg U65340 ( .A(n26407), .X(n50647) );
  nand_x1_sg U65341 ( .A(n26685), .B(n26684), .X(n26682) );
  inv_x1_sg U65342 ( .A(n26685), .X(n50934) );
  nand_x1_sg U65343 ( .A(n41418), .B(n17465), .X(n17464) );
  nand_x1_sg U65344 ( .A(n50524), .B(n50522), .X(n26130) );
  nand_x1_sg U65345 ( .A(n26131), .B(n16840), .X(n26129) );
  inv_x1_sg U65346 ( .A(n26131), .X(n50524) );
  nand_x1_sg U65347 ( .A(n46924), .B(n22775), .X(n22772) );
  inv_x1_sg U65348 ( .A(n22775), .X(n46943) );
  nand_x1_sg U65349 ( .A(n22754), .B(n22753), .X(n22751) );
  inv_x1_sg U65350 ( .A(n22754), .X(n47008) );
  nand_x1_sg U65351 ( .A(n23031), .B(n23030), .X(n23028) );
  inv_x1_sg U65352 ( .A(n23031), .X(n47296) );
  nand_x1_sg U65353 ( .A(n23311), .B(n23310), .X(n23308) );
  inv_x1_sg U65354 ( .A(n23311), .X(n47581) );
  nand_x1_sg U65355 ( .A(n23590), .B(n23589), .X(n23587) );
  inv_x1_sg U65356 ( .A(n23590), .X(n47866) );
  nand_x1_sg U65357 ( .A(n23869), .B(n23868), .X(n23866) );
  inv_x1_sg U65358 ( .A(n23869), .X(n48151) );
  nand_x1_sg U65359 ( .A(n24148), .B(n24147), .X(n24145) );
  inv_x1_sg U65360 ( .A(n24148), .X(n48436) );
  nand_x1_sg U65361 ( .A(n24427), .B(n24426), .X(n24424) );
  inv_x1_sg U65362 ( .A(n24427), .X(n48721) );
  nand_x1_sg U65363 ( .A(n24705), .B(n24704), .X(n24702) );
  inv_x1_sg U65364 ( .A(n24705), .X(n49007) );
  nand_x1_sg U65365 ( .A(n24984), .B(n24983), .X(n24981) );
  inv_x1_sg U65366 ( .A(n24984), .X(n49294) );
  nand_x1_sg U65367 ( .A(n25263), .B(n25262), .X(n25260) );
  inv_x1_sg U65368 ( .A(n25263), .X(n49580) );
  nand_x1_sg U65369 ( .A(n25542), .B(n25541), .X(n25539) );
  inv_x1_sg U65370 ( .A(n25542), .X(n49866) );
  nand_x1_sg U65371 ( .A(n25819), .B(n25818), .X(n25816) );
  inv_x1_sg U65372 ( .A(n25819), .X(n50152) );
  nand_x1_sg U65373 ( .A(n26053), .B(n26054), .X(n26051) );
  inv_x1_sg U65374 ( .A(n26053), .X(n50437) );
  nand_x1_sg U65375 ( .A(n26379), .B(n26378), .X(n26376) );
  inv_x1_sg U65376 ( .A(n26379), .X(n50726) );
  nand_x1_sg U65377 ( .A(n26657), .B(n26656), .X(n26654) );
  inv_x1_sg U65378 ( .A(n26657), .X(n51013) );
  nor_x1_sg U65379 ( .A(n25495), .B(n18286), .X(n19120) );
  nand_x1_sg U65380 ( .A(n50500), .B(n26137), .X(n26134) );
  inv_x1_sg U65381 ( .A(n26137), .X(n50502) );
  nor_x1_sg U65382 ( .A(n42334), .B(n41079), .X(n5985) );
  nor_x1_sg U65383 ( .A(n41533), .B(n38922), .X(n6133) );
  nor_x1_sg U65384 ( .A(n46339), .B(n41079), .X(n6270) );
  nor_x1_sg U65385 ( .A(n46202), .B(n41076), .X(n6404) );
  nor_x1_sg U65386 ( .A(n46066), .B(n41077), .X(n6537) );
  nor_x1_sg U65387 ( .A(n6674), .B(n41078), .X(n6673) );
  nor_x1_sg U65388 ( .A(n39446), .B(n45804), .X(n6816) );
  nor_x1_sg U65389 ( .A(n38710), .B(n41010), .X(n6021) );
  nor_x1_sg U65390 ( .A(n38725), .B(n41254), .X(n6168) );
  nor_x1_sg U65391 ( .A(n38711), .B(n41011), .X(n6208) );
  nor_x1_sg U65392 ( .A(n38712), .B(n41031), .X(n6070) );
  nor_x1_sg U65393 ( .A(n46848), .B(n22837), .X(n6834) );
  inv_x1_sg U65394 ( .A(n22839), .X(n46848) );
  nor_x1_sg U65395 ( .A(n5964), .B(n41005), .X(n5963) );
  nor_x1_sg U65396 ( .A(n5965), .B(n41039), .X(n5962) );
  nor_x1_sg U65397 ( .A(n5968), .B(n41031), .X(n5967) );
  nor_x1_sg U65398 ( .A(n5974), .B(n41252), .X(n5973) );
  nor_x1_sg U65399 ( .A(n6077), .B(n41251), .X(n6076) );
  nand_x1_sg U65400 ( .A(n39564), .B(n40632), .X(n8312) );
  nand_x1_sg U65401 ( .A(n39567), .B(n40628), .X(n9130) );
  nand_x1_sg U65402 ( .A(n39570), .B(n40668), .X(n9950) );
  nand_x1_sg U65403 ( .A(n39573), .B(n40657), .X(n10769) );
  nand_x1_sg U65404 ( .A(n39576), .B(n40642), .X(n11588) );
  nand_x1_sg U65405 ( .A(n39579), .B(n40639), .X(n12407) );
  nand_x1_sg U65406 ( .A(n39582), .B(n40663), .X(n13226) );
  nand_x1_sg U65407 ( .A(n39585), .B(n40653), .X(n14045) );
  nand_x1_sg U65408 ( .A(n39588), .B(n40622), .X(n14864) );
  nand_x1_sg U65409 ( .A(n39591), .B(n40682), .X(n15683) );
  nand_x1_sg U65410 ( .A(n39594), .B(n40679), .X(n16502) );
  nand_x1_sg U65411 ( .A(n39561), .B(n40580), .X(n17319) );
  nand_x1_sg U65412 ( .A(n39597), .B(n40672), .X(n18961) );
  nor_x1_sg U65413 ( .A(n6003), .B(n39445), .X(n6001) );
  nor_x1_sg U65414 ( .A(n6087), .B(n41077), .X(n6086) );
  nor_x1_sg U65415 ( .A(n6161), .B(n41003), .X(n6160) );
  nor_x1_sg U65416 ( .A(n42342), .B(n41072), .X(n5984) );
  nor_x1_sg U65417 ( .A(n6134), .B(n41074), .X(n6132) );
  nor_x1_sg U65418 ( .A(n42224), .B(n39264), .X(n6269) );
  nor_x1_sg U65419 ( .A(n42221), .B(n38919), .X(n6403) );
  nor_x1_sg U65420 ( .A(n42219), .B(n41073), .X(n6536) );
  nor_x1_sg U65421 ( .A(n42217), .B(n41074), .X(n6672) );
  inv_x1_sg U65422 ( .A(n19156), .X(n46570) );
  nor_x1_sg U65423 ( .A(n42330), .B(n41573), .X(n6018) );
  nor_x1_sg U65424 ( .A(n42331), .B(n41011), .X(n6069) );
  nor_x1_sg U65425 ( .A(n42341), .B(n39264), .X(n6085) );
  nor_x1_sg U65426 ( .A(n6023), .B(n41031), .X(n6022) );
  nor_x1_sg U65427 ( .A(n6055), .B(n41571), .X(n6054) );
  nor_x1_sg U65428 ( .A(n6210), .B(n41030), .X(n6209) );
  nor_x1_sg U65429 ( .A(n6142), .B(n41026), .X(n6139) );
  nor_x1_sg U65430 ( .A(n6188), .B(n41023), .X(n6185) );
  nor_x1_sg U65431 ( .A(n6207), .B(n41566), .X(n6205) );
  nor_x1_sg U65432 ( .A(n6234), .B(n41024), .X(n6231) );
  nor_x1_sg U65433 ( .A(n6255), .B(n41040), .X(n6252) );
  nor_x1_sg U65434 ( .A(n6279), .B(n38937), .X(n6276) );
  nor_x1_sg U65435 ( .A(n6285), .B(n41365), .X(n6282) );
  nor_x1_sg U65436 ( .A(n6300), .B(n41038), .X(n6297) );
  nor_x1_sg U65437 ( .A(n6323), .B(n41025), .X(n6320) );
  nor_x1_sg U65438 ( .A(n6329), .B(n39906), .X(n6326) );
  nor_x1_sg U65439 ( .A(n6344), .B(n41038), .X(n6341) );
  nor_x1_sg U65440 ( .A(n6368), .B(n41026), .X(n6365) );
  nor_x1_sg U65441 ( .A(n6374), .B(n41368), .X(n6371) );
  nor_x1_sg U65442 ( .A(n6389), .B(n41041), .X(n6386) );
  nor_x1_sg U65443 ( .A(n6412), .B(n41026), .X(n6409) );
  nor_x1_sg U65444 ( .A(n6418), .B(n41367), .X(n6415) );
  nor_x1_sg U65445 ( .A(n6433), .B(n41041), .X(n6430) );
  nor_x1_sg U65446 ( .A(n6457), .B(n41025), .X(n6454) );
  nor_x1_sg U65447 ( .A(n6463), .B(n39446), .X(n6460) );
  nor_x1_sg U65448 ( .A(n6478), .B(n41039), .X(n6475) );
  nor_x1_sg U65449 ( .A(n6501), .B(n41023), .X(n6498) );
  nor_x1_sg U65450 ( .A(n6507), .B(n41366), .X(n6504) );
  nor_x1_sg U65451 ( .A(n6522), .B(n41041), .X(n6519) );
  nor_x1_sg U65452 ( .A(n6546), .B(n41025), .X(n6543) );
  nor_x1_sg U65453 ( .A(n6552), .B(n38973), .X(n6549) );
  nor_x1_sg U65454 ( .A(n6567), .B(n41039), .X(n6564) );
  nor_x1_sg U65455 ( .A(n6590), .B(n41024), .X(n6587) );
  nor_x1_sg U65456 ( .A(n6596), .B(n39446), .X(n6593) );
  nor_x1_sg U65457 ( .A(n6611), .B(n41038), .X(n6608) );
  nor_x1_sg U65458 ( .A(n6635), .B(n41026), .X(n6632) );
  nor_x1_sg U65459 ( .A(n6641), .B(n41368), .X(n6638) );
  nor_x1_sg U65460 ( .A(n42343), .B(n41020), .X(n6680) );
  nor_x1_sg U65461 ( .A(n5998), .B(n38937), .X(n5996) );
  nor_x1_sg U65462 ( .A(n6038), .B(n41074), .X(n6036) );
  nor_x1_sg U65463 ( .A(n6096), .B(n41569), .X(n6094) );
  nor_x1_sg U65464 ( .A(n6118), .B(n41030), .X(n6117) );
  nor_x1_sg U65465 ( .A(n6226), .B(n41072), .X(n6224) );
  nor_x1_sg U65466 ( .A(n6664), .B(n41252), .X(n6663) );
  nor_x1_sg U65467 ( .A(n6655), .B(n41004), .X(n6654) );
  nor_x1_sg U65468 ( .A(n6687), .B(n40978), .X(n6686) );
  nor_x1_sg U65469 ( .A(n42335), .B(n41034), .X(n6005) );
  nor_x1_sg U65470 ( .A(n42333), .B(n41074), .X(n6177) );
  nor_x1_sg U65471 ( .A(n42340), .B(n39906), .X(n22442) );
  nor_x1_sg U65472 ( .A(n41532), .B(n39907), .X(n6145) );
  nor_x1_sg U65473 ( .A(n42298), .B(n41367), .X(n6685) );
  nor_x1_sg U65474 ( .A(n26781), .B(n38973), .X(n26773) );
  nor_x1_sg U65475 ( .A(n42228), .B(n39445), .X(n21784) );
  nor_x1_sg U65476 ( .A(n42156), .B(n39907), .X(n21924) );
  nor_x1_sg U65477 ( .A(n42153), .B(n41367), .X(n22064) );
  nor_x1_sg U65478 ( .A(n22211), .B(n41366), .X(n22205) );
  nor_x1_sg U65479 ( .A(n22354), .B(n39906), .X(n22348) );
  nor_x1_sg U65480 ( .A(n41540), .B(n39445), .X(n22488) );
  nor_x1_sg U65481 ( .A(n22638), .B(n22628), .X(n22637) );
  nand_x1_sg U65482 ( .A(n39205), .B(n40082), .X(n7217) );
  inv_x1_sg U65483 ( .A(n42058), .X(n51181) );
  nor_x1_sg U65484 ( .A(n42283), .B(n39907), .X(n6049) );
  nor_x1_sg U65485 ( .A(n42295), .B(n41025), .X(n6044) );
  nor_x1_sg U65486 ( .A(n42284), .B(n40980), .X(n6238) );
  nor_x1_sg U65487 ( .A(n42282), .B(n41251), .X(n6261) );
  nor_x1_sg U65488 ( .A(n42294), .B(n41006), .X(n6253) );
  nor_x1_sg U65489 ( .A(n42296), .B(n40979), .X(n6283) );
  nor_x1_sg U65490 ( .A(n42281), .B(n41251), .X(n6306) );
  nor_x1_sg U65491 ( .A(n42293), .B(n41004), .X(n6298) );
  nor_x1_sg U65492 ( .A(n42297), .B(n38925), .X(n6327) );
  nor_x1_sg U65493 ( .A(n42280), .B(n41254), .X(n6350) );
  nor_x1_sg U65494 ( .A(n42292), .B(n41006), .X(n6342) );
  nor_x1_sg U65495 ( .A(n42231), .B(n40980), .X(n6372) );
  nor_x1_sg U65496 ( .A(n42279), .B(n39116), .X(n6395) );
  nor_x1_sg U65497 ( .A(n42291), .B(n41003), .X(n6387) );
  nor_x1_sg U65498 ( .A(n42299), .B(n40979), .X(n6416) );
  nor_x1_sg U65499 ( .A(n42268), .B(n39116), .X(n6439) );
  nor_x1_sg U65500 ( .A(n42286), .B(n41005), .X(n6431) );
  nor_x1_sg U65501 ( .A(n42232), .B(n40979), .X(n6461) );
  nor_x1_sg U65502 ( .A(n42278), .B(n42018), .X(n6484) );
  nor_x1_sg U65503 ( .A(n42290), .B(n41006), .X(n6476) );
  nor_x1_sg U65504 ( .A(n42234), .B(n40979), .X(n6505) );
  nor_x1_sg U65505 ( .A(n42277), .B(n42018), .X(n6528) );
  nor_x1_sg U65506 ( .A(n42289), .B(n41004), .X(n6520) );
  nor_x1_sg U65507 ( .A(n42301), .B(n40980), .X(n6550) );
  nor_x1_sg U65508 ( .A(n42230), .B(n41253), .X(n6573) );
  nor_x1_sg U65509 ( .A(n42288), .B(n38927), .X(n6565) );
  nor_x1_sg U65510 ( .A(n42233), .B(n40977), .X(n6594) );
  nor_x1_sg U65511 ( .A(n42276), .B(n41252), .X(n6617) );
  nor_x1_sg U65512 ( .A(n42287), .B(n41573), .X(n6609) );
  nor_x1_sg U65513 ( .A(n42300), .B(n40978), .X(n6639) );
  nand_x1_sg U65514 ( .A(n41900), .B(n40158), .X(n7893) );
  nand_x1_sg U65515 ( .A(n41887), .B(n40359), .X(n8711) );
  nand_x1_sg U65516 ( .A(n41878), .B(n40355), .X(n9531) );
  nand_x1_sg U65517 ( .A(n39816), .B(n40351), .X(n10350) );
  nand_x1_sg U65518 ( .A(n39834), .B(n40347), .X(n11169) );
  nand_x1_sg U65519 ( .A(n39837), .B(n40327), .X(n11988) );
  nand_x1_sg U65520 ( .A(n39819), .B(n40339), .X(n12807) );
  nand_x1_sg U65521 ( .A(n41881), .B(n40335), .X(n13626) );
  nand_x1_sg U65522 ( .A(n41879), .B(n40343), .X(n14445) );
  nand_x1_sg U65523 ( .A(n39849), .B(n40320), .X(n15264) );
  nand_x1_sg U65524 ( .A(n39821), .B(n40323), .X(n16083) );
  nand_x1_sg U65525 ( .A(n39825), .B(n40331), .X(n18542) );
  nor_x1_sg U65526 ( .A(n41071), .B(n45810), .X(n6805) );
  nor_x1_sg U65527 ( .A(n19527), .B(n39445), .X(n20572) );
  nor_x1_sg U65528 ( .A(n6102), .B(n41366), .X(n6099) );
  nor_x1_sg U65529 ( .A(n46424), .B(n38972), .X(n6191) );
  nor_x1_sg U65530 ( .A(n6240), .B(n38972), .X(n6237) );
  nor_x1_sg U65531 ( .A(n41535), .B(n38972), .X(n6728) );
  nor_x1_sg U65532 ( .A(n6778), .B(n38973), .X(n6775) );
  nor_x1_sg U65533 ( .A(n45753), .B(n39446), .X(n21737) );
  nor_x1_sg U65534 ( .A(n42158), .B(n38973), .X(n21831) );
  nor_x1_sg U65535 ( .A(n42157), .B(n39906), .X(n21878) );
  nor_x1_sg U65536 ( .A(n42155), .B(n41368), .X(n21971) );
  nor_x1_sg U65537 ( .A(n42154), .B(n39907), .X(n22017) );
  nor_x1_sg U65538 ( .A(n22116), .B(n41366), .X(n22110) );
  nor_x1_sg U65539 ( .A(n22164), .B(n41365), .X(n22158) );
  nor_x1_sg U65540 ( .A(n22259), .B(n38972), .X(n22253) );
  nor_x1_sg U65541 ( .A(n22306), .B(n41365), .X(n22300) );
  nor_x1_sg U65542 ( .A(n22401), .B(n41368), .X(n22395) );
  nor_x1_sg U65543 ( .A(n22535), .B(n41365), .X(n22531) );
  nor_x1_sg U65544 ( .A(n44969), .B(n41367), .X(n22570) );
  nor_x1_sg U65545 ( .A(n6162), .B(n41040), .X(n6159) );
  nor_x1_sg U65546 ( .A(n6216), .B(n41253), .X(n6215) );
  nor_x1_sg U65547 ( .A(n6659), .B(n41568), .X(n6658) );
  nor_x1_sg U65548 ( .A(n6691), .B(n41013), .X(n6690) );
  nor_x1_sg U65549 ( .A(n6051), .B(n40978), .X(n6050) );
  nor_x1_sg U65550 ( .A(n47140), .B(n23114), .X(n7651) );
  inv_x1_sg U65551 ( .A(n23116), .X(n47140) );
  nor_x1_sg U65552 ( .A(n47425), .B(n23394), .X(n8469) );
  inv_x1_sg U65553 ( .A(n23396), .X(n47425) );
  nor_x1_sg U65554 ( .A(n47710), .B(n23673), .X(n9289) );
  inv_x1_sg U65555 ( .A(n23675), .X(n47710) );
  nor_x1_sg U65556 ( .A(n47995), .B(n23952), .X(n10108) );
  inv_x1_sg U65557 ( .A(n23954), .X(n47995) );
  nor_x1_sg U65558 ( .A(n48280), .B(n24231), .X(n10927) );
  inv_x1_sg U65559 ( .A(n24233), .X(n48280) );
  nor_x1_sg U65560 ( .A(n48565), .B(n24510), .X(n11746) );
  inv_x1_sg U65561 ( .A(n24512), .X(n48565) );
  nor_x1_sg U65562 ( .A(n48850), .B(n24788), .X(n12565) );
  inv_x1_sg U65563 ( .A(n24790), .X(n48850) );
  nor_x1_sg U65564 ( .A(n49137), .B(n25067), .X(n13384) );
  inv_x1_sg U65565 ( .A(n25069), .X(n49137) );
  nor_x1_sg U65566 ( .A(n49423), .B(n25346), .X(n14203) );
  inv_x1_sg U65567 ( .A(n25348), .X(n49423) );
  nor_x1_sg U65568 ( .A(n49709), .B(n25625), .X(n15022) );
  inv_x1_sg U65569 ( .A(n25627), .X(n49709) );
  nor_x1_sg U65570 ( .A(n49995), .B(n25902), .X(n15841) );
  inv_x1_sg U65571 ( .A(n25904), .X(n49995) );
  nor_x1_sg U65572 ( .A(n50570), .B(n26462), .X(n17479) );
  inv_x1_sg U65573 ( .A(n26464), .X(n50570) );
  nor_x1_sg U65574 ( .A(n50856), .B(n26740), .X(n18300) );
  inv_x1_sg U65575 ( .A(n26742), .X(n50856) );
  nor_x1_sg U65576 ( .A(n6101), .B(n40978), .X(n6100) );
  nor_x1_sg U65577 ( .A(n6147), .B(n40977), .X(n6146) );
  nor_x1_sg U65578 ( .A(n6193), .B(n40977), .X(n6192) );
  nand_x1_sg U65579 ( .A(n40608), .B(n42092), .X(n16902) );
  nand_x1_sg U65580 ( .A(n39827), .B(n42091), .X(n17721) );
  nand_x1_sg U65581 ( .A(n39851), .B(n40574), .X(n7494) );
  nor_x1_sg U65582 ( .A(n40563), .B(n39481), .X(n25930) );
  nand_x1_sg U65583 ( .A(n41901), .B(n39956), .X(n7075) );
  nor_x1_sg U65584 ( .A(n39065), .B(n41193), .X(n22883) );
  nor_x1_sg U65585 ( .A(n39064), .B(n39224), .X(n23160) );
  nor_x1_sg U65586 ( .A(n39063), .B(n41183), .X(n23440) );
  nor_x1_sg U65587 ( .A(n39062), .B(n41180), .X(n23719) );
  nor_x1_sg U65588 ( .A(n39061), .B(n41866), .X(n23998) );
  nor_x1_sg U65589 ( .A(n39060), .B(n39232), .X(n24277) );
  nor_x1_sg U65590 ( .A(n39059), .B(n41165), .X(n24556) );
  nor_x1_sg U65591 ( .A(n39058), .B(n41157), .X(n24834) );
  nor_x1_sg U65592 ( .A(n39057), .B(n41870), .X(n25113) );
  nor_x1_sg U65593 ( .A(n39056), .B(n41150), .X(n25392) );
  nor_x1_sg U65594 ( .A(n39055), .B(n41143), .X(n25671) );
  nor_x1_sg U65595 ( .A(n39053), .B(n41140), .X(n26215) );
  nor_x1_sg U65596 ( .A(n39054), .B(n41135), .X(n26508) );
  nor_x1_sg U65597 ( .A(n19510), .B(n39263), .X(n19509) );
  nor_x1_sg U65598 ( .A(n41971), .B(n41078), .X(n6037) );
  nor_x1_sg U65599 ( .A(n42024), .B(n41078), .X(n6178) );
  nor_x1_sg U65600 ( .A(n41531), .B(n39263), .X(n6225) );
  nor_x1_sg U65601 ( .A(n46293), .B(n41079), .X(n6315) );
  nor_x1_sg U65602 ( .A(n46248), .B(n41079), .X(n6359) );
  nor_x1_sg U65603 ( .A(n46157), .B(n41077), .X(n6448) );
  nor_x1_sg U65604 ( .A(n46111), .B(n39263), .X(n6493) );
  nor_x1_sg U65605 ( .A(n46020), .B(n41078), .X(n6582) );
  nor_x1_sg U65606 ( .A(n45975), .B(n41077), .X(n6626) );
  nor_x1_sg U65607 ( .A(n42225), .B(n39263), .X(n6718) );
  nor_x1_sg U65608 ( .A(n6763), .B(n41076), .X(n6762) );
  nor_x1_sg U65609 ( .A(n42105), .B(n41192), .X(n22862) );
  nor_x1_sg U65610 ( .A(n40359), .B(n39224), .X(n23139) );
  nor_x1_sg U65611 ( .A(n40355), .B(n41182), .X(n23419) );
  nor_x1_sg U65612 ( .A(n40351), .B(n39228), .X(n23698) );
  nor_x1_sg U65613 ( .A(n40347), .B(n41172), .X(n23977) );
  nor_x1_sg U65614 ( .A(n40327), .B(n39232), .X(n24256) );
  nor_x1_sg U65615 ( .A(n40339), .B(n41163), .X(n24535) );
  nor_x1_sg U65616 ( .A(n40335), .B(n41160), .X(n24813) );
  nor_x1_sg U65617 ( .A(n40343), .B(n41152), .X(n25092) );
  nor_x1_sg U65618 ( .A(n40319), .B(n41871), .X(n25371) );
  nor_x1_sg U65619 ( .A(n40323), .B(n41145), .X(n25650) );
  nor_x1_sg U65620 ( .A(n40331), .B(n41133), .X(n26487) );
  nor_x1_sg U65621 ( .A(n40634), .B(n41194), .X(n22897) );
  nor_x1_sg U65622 ( .A(n40627), .B(n41863), .X(n23174) );
  nor_x1_sg U65623 ( .A(n40669), .B(n41184), .X(n23454) );
  nor_x1_sg U65624 ( .A(n40658), .B(n41180), .X(n23733) );
  nor_x1_sg U65625 ( .A(n40643), .B(n41173), .X(n24012) );
  nor_x1_sg U65626 ( .A(n40637), .B(n41167), .X(n24291) );
  nor_x1_sg U65627 ( .A(n40663), .B(n41165), .X(n24570) );
  nor_x1_sg U65628 ( .A(n40653), .B(n41159), .X(n24848) );
  nor_x1_sg U65629 ( .A(n40623), .B(n41155), .X(n25127) );
  nor_x1_sg U65630 ( .A(n40683), .B(n39240), .X(n25406) );
  nor_x1_sg U65631 ( .A(n40679), .B(n39242), .X(n25685) );
  nor_x1_sg U65632 ( .A(n40648), .B(n41139), .X(n26231) );
  nor_x1_sg U65633 ( .A(n40674), .B(n41134), .X(n26522) );
  nor_x1_sg U65634 ( .A(n26029), .B(n38941), .X(n26030) );
  nor_x1_sg U65635 ( .A(n6753), .B(n39116), .X(n6752) );
  nor_x1_sg U65636 ( .A(n6743), .B(n41005), .X(n6742) );
  nor_x1_sg U65637 ( .A(n6747), .B(n41031), .X(n6746) );
  nor_x1_sg U65638 ( .A(n6777), .B(n40980), .X(n6776) );
  nor_x1_sg U65639 ( .A(n6781), .B(n41014), .X(n6780) );
  nor_x1_sg U65640 ( .A(n6764), .B(n41073), .X(n6761) );
  nor_x1_sg U65641 ( .A(n6744), .B(n41040), .X(n6741) );
  nor_x1_sg U65642 ( .A(n6771), .B(n38935), .X(n6770) );
  nor_x1_sg U65643 ( .A(n40069), .B(n41947), .X(n25924) );
  nor_x1_sg U65644 ( .A(n42091), .B(n39244), .X(n26191) );
  nand_x1_sg U65645 ( .A(n41783), .B(n40134), .X(n8036) );
  nand_x1_sg U65646 ( .A(n39207), .B(n42183), .X(n8854) );
  nand_x1_sg U65647 ( .A(n41787), .B(n42181), .X(n9674) );
  nand_x1_sg U65648 ( .A(n41789), .B(n42179), .X(n10493) );
  nand_x1_sg U65649 ( .A(n39210), .B(n42177), .X(n11312) );
  nand_x1_sg U65650 ( .A(n41793), .B(n42175), .X(n12131) );
  nand_x1_sg U65651 ( .A(n39212), .B(n42173), .X(n12950) );
  nand_x1_sg U65652 ( .A(n39213), .B(n42171), .X(n13769) );
  nand_x1_sg U65653 ( .A(n39214), .B(n42169), .X(n14588) );
  nand_x1_sg U65654 ( .A(n39490), .B(n40152), .X(n15407) );
  nand_x1_sg U65655 ( .A(n39216), .B(n42166), .X(n16226) );
  nand_x1_sg U65656 ( .A(n39217), .B(n40160), .X(n17864) );
  nand_x1_sg U65657 ( .A(n39218), .B(n42164), .X(n18685) );
  nor_x1_sg U65658 ( .A(n22985), .B(n47415), .X(n22860) );
  inv_x1_sg U65659 ( .A(n22986), .X(n47415) );
  nor_x1_sg U65660 ( .A(n23265), .B(n47700), .X(n23137) );
  inv_x1_sg U65661 ( .A(n23266), .X(n47700) );
  nor_x1_sg U65662 ( .A(n23544), .B(n47985), .X(n23417) );
  inv_x1_sg U65663 ( .A(n23545), .X(n47985) );
  nor_x1_sg U65664 ( .A(n23823), .B(n48270), .X(n23696) );
  inv_x1_sg U65665 ( .A(n23824), .X(n48270) );
  nor_x1_sg U65666 ( .A(n24102), .B(n48555), .X(n23975) );
  inv_x1_sg U65667 ( .A(n24103), .X(n48555) );
  nor_x1_sg U65668 ( .A(n24381), .B(n48840), .X(n24254) );
  inv_x1_sg U65669 ( .A(n24382), .X(n48840) );
  nor_x1_sg U65670 ( .A(n24659), .B(n49127), .X(n24533) );
  inv_x1_sg U65671 ( .A(n24660), .X(n49127) );
  nor_x1_sg U65672 ( .A(n24938), .B(n49413), .X(n24811) );
  inv_x1_sg U65673 ( .A(n24939), .X(n49413) );
  nor_x1_sg U65674 ( .A(n25217), .B(n49699), .X(n25090) );
  inv_x1_sg U65675 ( .A(n25218), .X(n49699) );
  nor_x1_sg U65676 ( .A(n25496), .B(n49985), .X(n25369) );
  inv_x1_sg U65677 ( .A(n25497), .X(n49985) );
  nor_x1_sg U65678 ( .A(n25773), .B(n50271), .X(n25648) );
  inv_x1_sg U65679 ( .A(n25774), .X(n50271) );
  nor_x1_sg U65680 ( .A(n26333), .B(n50846), .X(n26189) );
  inv_x1_sg U65681 ( .A(n26334), .X(n50846) );
  nor_x1_sg U65682 ( .A(n26611), .B(n51132), .X(n26485) );
  inv_x1_sg U65683 ( .A(n26612), .X(n51132) );
  nand_x1_sg U65684 ( .A(n40586), .B(n41292), .X(n15829) );
  nand_x1_sg U65685 ( .A(n40584), .B(n39107), .X(n8457) );
  nand_x1_sg U65686 ( .A(n40584), .B(n39113), .X(n9277) );
  nand_x1_sg U65687 ( .A(n40584), .B(n41200), .X(n10096) );
  nand_x1_sg U65688 ( .A(n40583), .B(n41223), .X(n10915) );
  nand_x1_sg U65689 ( .A(n40585), .B(n41203), .X(n11734) );
  nand_x1_sg U65690 ( .A(n40586), .B(n39119), .X(n12553) );
  nand_x1_sg U65691 ( .A(n40586), .B(n41243), .X(n13372) );
  nand_x1_sg U65692 ( .A(n40585), .B(n41227), .X(n14191) );
  nand_x1_sg U65693 ( .A(n40585), .B(n41234), .X(n15010) );
  nand_x1_sg U65694 ( .A(n40583), .B(n41261), .X(n18288) );
  nor_x1_sg U65695 ( .A(n6827), .B(n39659), .X(n22601) );
  nor_x1_sg U65696 ( .A(n19137), .B(n39264), .X(n19508) );
  nor_x1_sg U65697 ( .A(n42223), .B(n41071), .X(n6314) );
  nor_x1_sg U65698 ( .A(n42222), .B(n41071), .X(n6358) );
  nor_x1_sg U65699 ( .A(n42216), .B(n41073), .X(n6447) );
  nor_x1_sg U65700 ( .A(n42220), .B(n39264), .X(n6492) );
  nor_x1_sg U65701 ( .A(n42261), .B(n41073), .X(n6581) );
  nor_x1_sg U65702 ( .A(n42218), .B(n41072), .X(n6625) );
  nor_x1_sg U65703 ( .A(n41527), .B(n41072), .X(n6717) );
  inv_x1_sg U65704 ( .A(n6240), .X(n46376) );
  nor_x1_sg U65705 ( .A(n50285), .B(n26111), .X(n16850) );
  inv_x1_sg U65706 ( .A(n26114), .X(n50285) );
  nor_x1_sg U65707 ( .A(n20566), .B(n41021), .X(n20565) );
  nor_x1_sg U65708 ( .A(n19131), .B(n41253), .X(n19130) );
  nor_x1_sg U65709 ( .A(n19117), .B(n41003), .X(n19116) );
  nor_x1_sg U65710 ( .A(n19119), .B(n41039), .X(n19115) );
  nor_x1_sg U65711 ( .A(n19123), .B(n41028), .X(n19122) );
  nor_x1_sg U65712 ( .A(n20574), .B(n42332), .X(n20573) );
  nor_x1_sg U65713 ( .A(n20960), .B(n41014), .X(n20959) );
  nand_x1_sg U65714 ( .A(n41835), .B(n40158), .X(n7919) );
  nand_x1_sg U65715 ( .A(n41833), .B(n40358), .X(n8737) );
  nand_x1_sg U65716 ( .A(n41831), .B(n40354), .X(n9557) );
  nand_x1_sg U65717 ( .A(n41829), .B(n40350), .X(n10376) );
  nand_x1_sg U65718 ( .A(n41827), .B(n40346), .X(n11195) );
  nand_x1_sg U65719 ( .A(n41825), .B(n40326), .X(n12014) );
  nand_x1_sg U65720 ( .A(n41822), .B(n40338), .X(n12833) );
  nand_x1_sg U65721 ( .A(n41821), .B(n40334), .X(n13652) );
  nand_x1_sg U65722 ( .A(n41818), .B(n40342), .X(n14471) );
  nand_x1_sg U65723 ( .A(n41817), .B(n42095), .X(n15290) );
  nand_x1_sg U65724 ( .A(n41814), .B(n40322), .X(n16109) );
  nand_x1_sg U65725 ( .A(n41810), .B(n42091), .X(n17747) );
  nand_x1_sg U65726 ( .A(n18578), .B(n40330), .X(n18568) );
  nor_x1_sg U65727 ( .A(n22978), .B(n22979), .X(n22977) );
  nand_x1_sg U65728 ( .A(n41195), .B(n22980), .X(n22979) );
  nor_x1_sg U65729 ( .A(n23535), .B(n23536), .X(n23534) );
  nand_x1_sg U65730 ( .A(n41182), .B(n23537), .X(n23536) );
  nor_x1_sg U65731 ( .A(n23814), .B(n23815), .X(n23813) );
  nand_x1_sg U65732 ( .A(n41177), .B(n23816), .X(n23815) );
  nor_x1_sg U65733 ( .A(n24093), .B(n24094), .X(n24092) );
  nand_x1_sg U65734 ( .A(n40490), .B(n24095), .X(n24094) );
  nor_x1_sg U65735 ( .A(n24372), .B(n24373), .X(n24371) );
  nand_x1_sg U65736 ( .A(n41169), .B(n24374), .X(n24373) );
  nor_x1_sg U65737 ( .A(n24651), .B(n24652), .X(n24650) );
  nand_x1_sg U65738 ( .A(n41165), .B(n24653), .X(n24652) );
  nor_x1_sg U65739 ( .A(n24929), .B(n24930), .X(n24928) );
  nand_x1_sg U65740 ( .A(n41159), .B(n24931), .X(n24930) );
  nor_x1_sg U65741 ( .A(n25208), .B(n25209), .X(n25207) );
  nand_x1_sg U65742 ( .A(n40474), .B(n25210), .X(n25209) );
  nor_x1_sg U65743 ( .A(n25487), .B(n25488), .X(n25486) );
  nand_x1_sg U65744 ( .A(n39240), .B(n25489), .X(n25488) );
  nor_x1_sg U65745 ( .A(n25766), .B(n25767), .X(n25765) );
  nand_x1_sg U65746 ( .A(n41143), .B(n25768), .X(n25767) );
  nor_x1_sg U65747 ( .A(n26603), .B(n26604), .X(n26602) );
  nand_x1_sg U65748 ( .A(n39246), .B(n26605), .X(n26604) );
  nand_x1_sg U65749 ( .A(n7103), .B(n7104), .X(n7087) );
  nor_x1_sg U65750 ( .A(n41809), .B(n41903), .X(n7103) );
  nand_x1_sg U65751 ( .A(n7921), .B(n7922), .X(n7905) );
  nor_x1_sg U65752 ( .A(n39965), .B(n40307), .X(n7921) );
  nand_x1_sg U65753 ( .A(n8739), .B(n8740), .X(n8723) );
  nor_x1_sg U65754 ( .A(n39968), .B(n41843), .X(n8739) );
  nand_x1_sg U65755 ( .A(n9559), .B(n9560), .X(n9543) );
  nor_x1_sg U65756 ( .A(n39973), .B(n41853), .X(n9559) );
  nand_x1_sg U65757 ( .A(n10378), .B(n10379), .X(n10362) );
  nor_x1_sg U65758 ( .A(n40700), .B(n41855), .X(n10378) );
  nand_x1_sg U65759 ( .A(n11197), .B(n11198), .X(n11181) );
  nor_x1_sg U65760 ( .A(n41925), .B(n41851), .X(n11197) );
  nand_x1_sg U65761 ( .A(n12016), .B(n12017), .X(n12000) );
  nor_x1_sg U65762 ( .A(n39985), .B(n41857), .X(n12016) );
  nand_x1_sg U65763 ( .A(n12835), .B(n12836), .X(n12819) );
  nor_x1_sg U65764 ( .A(n39988), .B(n41859), .X(n12835) );
  nand_x1_sg U65765 ( .A(n13654), .B(n13655), .X(n13638) );
  nor_x1_sg U65766 ( .A(n39993), .B(n41849), .X(n13654) );
  nand_x1_sg U65767 ( .A(n14473), .B(n14474), .X(n14457) );
  nor_x1_sg U65768 ( .A(n39996), .B(n41836), .X(n14473) );
  nand_x1_sg U65769 ( .A(n15292), .B(n15293), .X(n15276) );
  nor_x1_sg U65770 ( .A(n39999), .B(n41845), .X(n15292) );
  nand_x1_sg U65771 ( .A(n16111), .B(n16112), .X(n16095) );
  nor_x1_sg U65772 ( .A(n40004), .B(n41838), .X(n16111) );
  nand_x1_sg U65773 ( .A(n17749), .B(n17750), .X(n17733) );
  nor_x1_sg U65774 ( .A(n38910), .B(n50565), .X(n17749) );
  nand_x1_sg U65775 ( .A(n18570), .B(n18571), .X(n18554) );
  nor_x1_sg U65776 ( .A(n41910), .B(n41840), .X(n18570) );
  nor_x1_sg U65777 ( .A(n8142), .B(n42185), .X(n8141) );
  nor_x1_sg U65778 ( .A(n8960), .B(n42183), .X(n8959) );
  nor_x1_sg U65779 ( .A(n9780), .B(n42181), .X(n9779) );
  nor_x1_sg U65780 ( .A(n10599), .B(n42179), .X(n10598) );
  nor_x1_sg U65781 ( .A(n11418), .B(n42177), .X(n11417) );
  nor_x1_sg U65782 ( .A(n12237), .B(n42175), .X(n12236) );
  nor_x1_sg U65783 ( .A(n13056), .B(n42173), .X(n13055) );
  nor_x1_sg U65784 ( .A(n13875), .B(n42171), .X(n13874) );
  nor_x1_sg U65785 ( .A(n14694), .B(n42169), .X(n14693) );
  nor_x1_sg U65786 ( .A(n15513), .B(n42168), .X(n15512) );
  nor_x1_sg U65787 ( .A(n16332), .B(n42166), .X(n16331) );
  nor_x1_sg U65788 ( .A(n17970), .B(n17800), .X(n17969) );
  nor_x1_sg U65789 ( .A(n18791), .B(n42164), .X(n18790) );
  nand_x1_sg U65790 ( .A(n40080), .B(n40234), .X(n7340) );
  nand_x1_sg U65791 ( .A(n40077), .B(n40231), .X(n17165) );
  nand_x1_sg U65792 ( .A(n16928), .B(n16929), .X(n16913) );
  nor_x1_sg U65793 ( .A(n40996), .B(n41842), .X(n16928) );
  nand_x1_sg U65794 ( .A(n40233), .B(n39956), .X(n7101) );
  nand_x1_sg U65795 ( .A(n40231), .B(n40069), .X(n16926) );
  nand_x1_sg U65796 ( .A(n7337), .B(n39852), .X(n7336) );
  nand_x1_sg U65797 ( .A(n46899), .B(n7141), .X(n7335) );
  nor_x1_sg U65798 ( .A(n7288), .B(n42325), .X(n7337) );
  nand_x1_sg U65799 ( .A(n8155), .B(n39564), .X(n8154) );
  nand_x1_sg U65800 ( .A(n47194), .B(n7959), .X(n8153) );
  nor_x1_sg U65801 ( .A(n8106), .B(n42089), .X(n8155) );
  nand_x1_sg U65802 ( .A(n8973), .B(n39567), .X(n8972) );
  nand_x1_sg U65803 ( .A(n47479), .B(n8777), .X(n8971) );
  nor_x1_sg U65804 ( .A(n8924), .B(n42130), .X(n8973) );
  nand_x1_sg U65805 ( .A(n9793), .B(n39570), .X(n9792) );
  nand_x1_sg U65806 ( .A(n47764), .B(n9597), .X(n9791) );
  nor_x1_sg U65807 ( .A(n9744), .B(n40043), .X(n9793) );
  nand_x1_sg U65808 ( .A(n10612), .B(n39573), .X(n10611) );
  nand_x1_sg U65809 ( .A(n48049), .B(n10416), .X(n10610) );
  nor_x1_sg U65810 ( .A(n10563), .B(n40046), .X(n10612) );
  nand_x1_sg U65811 ( .A(n11431), .B(n39576), .X(n11430) );
  nand_x1_sg U65812 ( .A(n48334), .B(n11235), .X(n11429) );
  nor_x1_sg U65813 ( .A(n11382), .B(n40047), .X(n11431) );
  nand_x1_sg U65814 ( .A(n12250), .B(n39579), .X(n12249) );
  nand_x1_sg U65815 ( .A(n48619), .B(n12054), .X(n12248) );
  nor_x1_sg U65816 ( .A(n12201), .B(n11996), .X(n12250) );
  nand_x1_sg U65817 ( .A(n13069), .B(n39582), .X(n13068) );
  nand_x1_sg U65818 ( .A(n48905), .B(n12873), .X(n13067) );
  nor_x1_sg U65819 ( .A(n13020), .B(n40051), .X(n13069) );
  nand_x1_sg U65820 ( .A(n13888), .B(n39585), .X(n13887) );
  nand_x1_sg U65821 ( .A(n49192), .B(n13692), .X(n13886) );
  nor_x1_sg U65822 ( .A(n13839), .B(n40065), .X(n13888) );
  nand_x1_sg U65823 ( .A(n14707), .B(n39588), .X(n14706) );
  nand_x1_sg U65824 ( .A(n49478), .B(n14511), .X(n14705) );
  nor_x1_sg U65825 ( .A(n14658), .B(n40053), .X(n14707) );
  nand_x1_sg U65826 ( .A(n15526), .B(n39591), .X(n15525) );
  nand_x1_sg U65827 ( .A(n49764), .B(n15330), .X(n15524) );
  nor_x1_sg U65828 ( .A(n15477), .B(n40055), .X(n15526) );
  nand_x1_sg U65829 ( .A(n16345), .B(n39594), .X(n16344) );
  nand_x1_sg U65830 ( .A(n50050), .B(n16149), .X(n16343) );
  nor_x1_sg U65831 ( .A(n16296), .B(n40058), .X(n16345) );
  nand_x1_sg U65832 ( .A(n17983), .B(n39600), .X(n17982) );
  nand_x1_sg U65833 ( .A(n50624), .B(n17787), .X(n17981) );
  nor_x1_sg U65834 ( .A(n17934), .B(n40060), .X(n17983) );
  nand_x1_sg U65835 ( .A(n18804), .B(n39597), .X(n18803) );
  nand_x1_sg U65836 ( .A(n50911), .B(n18608), .X(n18802) );
  nor_x1_sg U65837 ( .A(n18755), .B(n40061), .X(n18804) );
  inv_x1_sg U65838 ( .A(n39770), .X(n50301) );
  nor_x1_sg U65839 ( .A(n41307), .B(n40235), .X(n22619) );
  nor_x1_sg U65840 ( .A(n41295), .B(n40231), .X(n25942) );
  nand_x1_sg U65841 ( .A(n47097), .B(n47074), .X(n22725) );
  nand_x1_sg U65842 ( .A(n22726), .B(n7015), .X(n22724) );
  inv_x1_sg U65843 ( .A(n22726), .X(n47097) );
  nand_x1_sg U65844 ( .A(n47383), .B(n47360), .X(n23002) );
  nand_x1_sg U65845 ( .A(n23003), .B(n7833), .X(n23001) );
  inv_x1_sg U65846 ( .A(n23003), .X(n47383) );
  nand_x1_sg U65847 ( .A(n47668), .B(n47645), .X(n23282) );
  nand_x1_sg U65848 ( .A(n23283), .B(n8651), .X(n23281) );
  inv_x1_sg U65849 ( .A(n23283), .X(n47668) );
  nand_x1_sg U65850 ( .A(n47953), .B(n47930), .X(n23561) );
  nand_x1_sg U65851 ( .A(n23562), .B(n9471), .X(n23560) );
  inv_x1_sg U65852 ( .A(n23562), .X(n47953) );
  nand_x1_sg U65853 ( .A(n48238), .B(n48215), .X(n23840) );
  nand_x1_sg U65854 ( .A(n23841), .B(n10290), .X(n23839) );
  inv_x1_sg U65855 ( .A(n23841), .X(n48238) );
  nand_x1_sg U65856 ( .A(n48523), .B(n48500), .X(n24119) );
  nand_x1_sg U65857 ( .A(n24120), .B(n11109), .X(n24118) );
  inv_x1_sg U65858 ( .A(n24120), .X(n48523) );
  nand_x1_sg U65859 ( .A(n48808), .B(n48785), .X(n24398) );
  nand_x1_sg U65860 ( .A(n24399), .B(n11928), .X(n24397) );
  inv_x1_sg U65861 ( .A(n24399), .X(n48808) );
  nand_x1_sg U65862 ( .A(n49095), .B(n49072), .X(n24676) );
  nand_x1_sg U65863 ( .A(n24677), .B(n12747), .X(n24675) );
  inv_x1_sg U65864 ( .A(n24677), .X(n49095) );
  nand_x1_sg U65865 ( .A(n49381), .B(n49358), .X(n24955) );
  nand_x1_sg U65866 ( .A(n24956), .B(n13566), .X(n24954) );
  inv_x1_sg U65867 ( .A(n24956), .X(n49381) );
  nand_x1_sg U65868 ( .A(n49667), .B(n49644), .X(n25234) );
  nand_x1_sg U65869 ( .A(n25235), .B(n14385), .X(n25233) );
  inv_x1_sg U65870 ( .A(n25235), .X(n49667) );
  nand_x1_sg U65871 ( .A(n49953), .B(n49930), .X(n25513) );
  nand_x1_sg U65872 ( .A(n25514), .B(n15204), .X(n25512) );
  inv_x1_sg U65873 ( .A(n25514), .X(n49953) );
  nand_x1_sg U65874 ( .A(n50239), .B(n50216), .X(n25790) );
  nand_x1_sg U65875 ( .A(n25791), .B(n16023), .X(n25789) );
  inv_x1_sg U65876 ( .A(n25791), .X(n50239) );
  nand_x1_sg U65877 ( .A(n50813), .B(n50790), .X(n26350) );
  nand_x1_sg U65878 ( .A(n26351), .B(n17661), .X(n26349) );
  inv_x1_sg U65879 ( .A(n26351), .X(n50813) );
  nand_x1_sg U65880 ( .A(n51100), .B(n51077), .X(n26628) );
  nand_x1_sg U65881 ( .A(n26629), .B(n18482), .X(n26627) );
  inv_x1_sg U65882 ( .A(n26629), .X(n51100) );
  nand_x1_sg U65883 ( .A(n47198), .B(n8003), .X(n8002) );
  nand_x1_sg U65884 ( .A(n47180), .B(n8004), .X(n8001) );
  nand_x1_sg U65885 ( .A(n47483), .B(n8821), .X(n8820) );
  nand_x1_sg U65886 ( .A(n47465), .B(n8822), .X(n8819) );
  nand_x1_sg U65887 ( .A(n47768), .B(n9641), .X(n9640) );
  nand_x1_sg U65888 ( .A(n47750), .B(n9642), .X(n9639) );
  nand_x1_sg U65889 ( .A(n48053), .B(n10460), .X(n10459) );
  nand_x1_sg U65890 ( .A(n48035), .B(n10461), .X(n10458) );
  nand_x1_sg U65891 ( .A(n48338), .B(n11279), .X(n11278) );
  nand_x1_sg U65892 ( .A(n48320), .B(n11280), .X(n11277) );
  nand_x1_sg U65893 ( .A(n48623), .B(n12098), .X(n12097) );
  nand_x1_sg U65894 ( .A(n48605), .B(n12099), .X(n12096) );
  nand_x1_sg U65895 ( .A(n48909), .B(n12917), .X(n12916) );
  nand_x1_sg U65896 ( .A(n48891), .B(n12918), .X(n12915) );
  nand_x1_sg U65897 ( .A(n49196), .B(n13736), .X(n13735) );
  nand_x1_sg U65898 ( .A(n49178), .B(n13737), .X(n13734) );
  nand_x1_sg U65899 ( .A(n49482), .B(n14555), .X(n14554) );
  nand_x1_sg U65900 ( .A(n49464), .B(n14556), .X(n14553) );
  nand_x1_sg U65901 ( .A(n49768), .B(n15374), .X(n15373) );
  nand_x1_sg U65902 ( .A(n49749), .B(n15375), .X(n15372) );
  nand_x1_sg U65903 ( .A(n50054), .B(n16193), .X(n16192) );
  nand_x1_sg U65904 ( .A(n50036), .B(n16194), .X(n16191) );
  nand_x1_sg U65905 ( .A(n50339), .B(n17009), .X(n17008) );
  nand_x1_sg U65906 ( .A(n50321), .B(n17010), .X(n17007) );
  nand_x1_sg U65907 ( .A(n50628), .B(n17831), .X(n17830) );
  nand_x1_sg U65908 ( .A(n50610), .B(n17832), .X(n17829) );
  nand_x1_sg U65909 ( .A(n50915), .B(n18652), .X(n18651) );
  nand_x1_sg U65910 ( .A(n50897), .B(n18653), .X(n18650) );
  nand_x1_sg U65911 ( .A(n46887), .B(n7185), .X(n7182) );
  nand_x1_sg U65912 ( .A(n46905), .B(n7184), .X(n7183) );
  nand_x1_sg U65913 ( .A(n40133), .B(n41835), .X(n8158) );
  nand_x1_sg U65914 ( .A(n40136), .B(n41833), .X(n8976) );
  nand_x1_sg U65915 ( .A(n40138), .B(n9567), .X(n9796) );
  nand_x1_sg U65916 ( .A(n40140), .B(n41828), .X(n10615) );
  nand_x1_sg U65917 ( .A(n40142), .B(n41826), .X(n11434) );
  nand_x1_sg U65918 ( .A(n40144), .B(n41824), .X(n12253) );
  nand_x1_sg U65919 ( .A(n40146), .B(n41823), .X(n13072) );
  nand_x1_sg U65920 ( .A(n40148), .B(n13662), .X(n13891) );
  nand_x1_sg U65921 ( .A(n40150), .B(n41819), .X(n14710) );
  nand_x1_sg U65922 ( .A(n42168), .B(n41816), .X(n15529) );
  nand_x1_sg U65923 ( .A(n40154), .B(n41815), .X(n16348) );
  nand_x1_sg U65924 ( .A(n40159), .B(n41811), .X(n17986) );
  nand_x1_sg U65925 ( .A(n42164), .B(n41813), .X(n18807) );
  nor_x1_sg U65926 ( .A(n19494), .B(n19490), .X(n19579) );
  nor_x1_sg U65927 ( .A(n38923), .B(n45808), .X(n6792) );
  nor_x1_sg U65928 ( .A(n41024), .B(n45800), .X(n6812) );
  nor_x1_sg U65929 ( .A(n39660), .B(n40574), .X(n22631) );
  nor_x1_sg U65930 ( .A(n41296), .B(n40580), .X(n25954) );
  nand_x1_sg U65931 ( .A(n41692), .B(n40576), .X(n7587) );
  nand_x1_sg U65932 ( .A(n41665), .B(n40634), .X(n8405) );
  nand_x1_sg U65933 ( .A(n41688), .B(n40628), .X(n9223) );
  nand_x1_sg U65934 ( .A(n41690), .B(n40669), .X(n10043) );
  nand_x1_sg U65935 ( .A(n41686), .B(n40656), .X(n10862) );
  nand_x1_sg U65936 ( .A(n41684), .B(n40644), .X(n11681) );
  nand_x1_sg U65937 ( .A(n41682), .B(n40636), .X(n12500) );
  nand_x1_sg U65938 ( .A(n41680), .B(n40661), .X(n13319) );
  nand_x1_sg U65939 ( .A(n41678), .B(n40654), .X(n14138) );
  nand_x1_sg U65940 ( .A(n41676), .B(n40621), .X(n14957) );
  nand_x1_sg U65941 ( .A(n41663), .B(n40681), .X(n15776) );
  nand_x1_sg U65942 ( .A(n41674), .B(n40678), .X(n16595) );
  nand_x1_sg U65943 ( .A(n41672), .B(n40579), .X(n17412) );
  nand_x1_sg U65944 ( .A(n17946), .B(n40646), .X(n18233) );
  nand_x1_sg U65945 ( .A(n41668), .B(n40673), .X(n19054) );
  nand_x1_sg U65946 ( .A(n41692), .B(n40233), .X(n7508) );
  nand_x1_sg U65947 ( .A(n41665), .B(n41834), .X(n8326) );
  nand_x1_sg U65948 ( .A(n41688), .B(n41832), .X(n9144) );
  nand_x1_sg U65949 ( .A(n41690), .B(n41830), .X(n9964) );
  nand_x1_sg U65950 ( .A(n41686), .B(n41828), .X(n10783) );
  nand_x1_sg U65951 ( .A(n41684), .B(n41826), .X(n11602) );
  nand_x1_sg U65952 ( .A(n41682), .B(n41824), .X(n12421) );
  nand_x1_sg U65953 ( .A(n41680), .B(n12843), .X(n13240) );
  nand_x1_sg U65954 ( .A(n41678), .B(n41820), .X(n14059) );
  nand_x1_sg U65955 ( .A(n41676), .B(n14481), .X(n14878) );
  nand_x1_sg U65956 ( .A(n41663), .B(n41816), .X(n15697) );
  nand_x1_sg U65957 ( .A(n41674), .B(n16119), .X(n16516) );
  nand_x1_sg U65958 ( .A(n41672), .B(n40230), .X(n17333) );
  nand_x1_sg U65959 ( .A(n41670), .B(n41810), .X(n18154) );
  nand_x1_sg U65960 ( .A(n41668), .B(n41812), .X(n18975) );
  nand_x1_sg U65961 ( .A(n40082), .B(n40574), .X(n7444) );
  nand_x1_sg U65962 ( .A(n40078), .B(n40579), .X(n17269) );
  nor_x1_sg U65963 ( .A(n20777), .B(n38600), .X(n20792) );
  nor_x1_sg U65964 ( .A(n19480), .B(n19478), .X(n19586) );
  nor_x1_sg U65965 ( .A(n19938), .B(n46552), .X(n20597) );
  nor_x1_sg U65966 ( .A(n20437), .B(n46376), .X(n20450) );
  nor_x1_sg U65967 ( .A(n6666), .B(n45930), .X(n6665) );
  nor_x1_sg U65968 ( .A(n6668), .B(n6664), .X(n6666) );
  nand_x1_sg U65969 ( .A(n38606), .B(n6668), .X(n6667) );
  nand_x1_sg U65970 ( .A(n39798), .B(n40158), .X(n8314) );
  nand_x1_sg U65971 ( .A(n39800), .B(n40358), .X(n9132) );
  nand_x1_sg U65972 ( .A(n39794), .B(n40354), .X(n9952) );
  nand_x1_sg U65973 ( .A(n39796), .B(n40350), .X(n10771) );
  nand_x1_sg U65974 ( .A(n39790), .B(n40346), .X(n11590) );
  nand_x1_sg U65975 ( .A(n39792), .B(n40326), .X(n12409) );
  nand_x1_sg U65976 ( .A(n39786), .B(n40338), .X(n13228) );
  nand_x1_sg U65977 ( .A(n39788), .B(n40334), .X(n14047) );
  nand_x1_sg U65978 ( .A(n39782), .B(n40342), .X(n14866) );
  nand_x1_sg U65979 ( .A(n39784), .B(n40318), .X(n15685) );
  nand_x1_sg U65980 ( .A(n39778), .B(n40322), .X(n16504) );
  nand_x1_sg U65981 ( .A(n39777), .B(n40330), .X(n18963) );
  nand_x1_sg U65982 ( .A(n21143), .B(n38660), .X(n21141) );
  nor_x1_sg U65983 ( .A(n6234), .B(n21143), .X(n21142) );
  nand_x1_sg U65984 ( .A(n21137), .B(n38658), .X(n21135) );
  nor_x1_sg U65985 ( .A(n6279), .B(n21137), .X(n21136) );
  nand_x1_sg U65986 ( .A(n21131), .B(n38656), .X(n21129) );
  nor_x1_sg U65987 ( .A(n6323), .B(n21131), .X(n21130) );
  nand_x1_sg U65988 ( .A(n21125), .B(n38654), .X(n21123) );
  nor_x1_sg U65989 ( .A(n6368), .B(n21125), .X(n21124) );
  nand_x1_sg U65990 ( .A(n21119), .B(n38652), .X(n21117) );
  nor_x1_sg U65991 ( .A(n6412), .B(n21119), .X(n21118) );
  nand_x1_sg U65992 ( .A(n21113), .B(n38650), .X(n21111) );
  nor_x1_sg U65993 ( .A(n6457), .B(n21113), .X(n21112) );
  nand_x1_sg U65994 ( .A(n21107), .B(n38648), .X(n21105) );
  nor_x1_sg U65995 ( .A(n6501), .B(n21107), .X(n21106) );
  nand_x1_sg U65996 ( .A(n21101), .B(n38646), .X(n21099) );
  nor_x1_sg U65997 ( .A(n6546), .B(n21101), .X(n21100) );
  nand_x1_sg U65998 ( .A(n21095), .B(n38644), .X(n21093) );
  nor_x1_sg U65999 ( .A(n6590), .B(n21095), .X(n21094) );
  nand_x1_sg U66000 ( .A(n21089), .B(n38642), .X(n21087) );
  nor_x1_sg U66001 ( .A(n6635), .B(n21089), .X(n21088) );
  nand_x1_sg U66002 ( .A(n21149), .B(n38662), .X(n21147) );
  nor_x1_sg U66003 ( .A(n6188), .B(n21149), .X(n21148) );
  nand_x1_sg U66004 ( .A(n21155), .B(n38664), .X(n21153) );
  nor_x1_sg U66005 ( .A(n6142), .B(n21155), .X(n21154) );
  nand_x1_sg U66006 ( .A(n20428), .B(n38709), .X(n20426) );
  nor_x1_sg U66007 ( .A(n6285), .B(n20428), .X(n20427) );
  nand_x1_sg U66008 ( .A(n20422), .B(n38724), .X(n20420) );
  nor_x1_sg U66009 ( .A(n6329), .B(n20422), .X(n20421) );
  nand_x1_sg U66010 ( .A(n20416), .B(n38610), .X(n20414) );
  nor_x1_sg U66011 ( .A(n6374), .B(n20416), .X(n20415) );
  nand_x1_sg U66012 ( .A(n20410), .B(n38707), .X(n20408) );
  nor_x1_sg U66013 ( .A(n6418), .B(n20410), .X(n20409) );
  nand_x1_sg U66014 ( .A(n20404), .B(n38612), .X(n20402) );
  nor_x1_sg U66015 ( .A(n6463), .B(n20404), .X(n20403) );
  nand_x1_sg U66016 ( .A(n20398), .B(n38616), .X(n20396) );
  nor_x1_sg U66017 ( .A(n6507), .B(n20398), .X(n20397) );
  nand_x1_sg U66018 ( .A(n20392), .B(n38705), .X(n20390) );
  nor_x1_sg U66019 ( .A(n6552), .B(n20392), .X(n20391) );
  nand_x1_sg U66020 ( .A(n20386), .B(n38614), .X(n20384) );
  nor_x1_sg U66021 ( .A(n6596), .B(n20386), .X(n20385) );
  nand_x1_sg U66022 ( .A(n20380), .B(n38722), .X(n20378) );
  nor_x1_sg U66023 ( .A(n6641), .B(n20380), .X(n20379) );
  nand_x1_sg U66024 ( .A(n19695), .B(n38697), .X(n19693) );
  nor_x1_sg U66025 ( .A(n6255), .B(n19695), .X(n19694) );
  nand_x1_sg U66026 ( .A(n19689), .B(n38691), .X(n19687) );
  nor_x1_sg U66027 ( .A(n6300), .B(n19689), .X(n19688) );
  nand_x1_sg U66028 ( .A(n19683), .B(n38687), .X(n19681) );
  nor_x1_sg U66029 ( .A(n6344), .B(n19683), .X(n19682) );
  nand_x1_sg U66030 ( .A(n19677), .B(n38685), .X(n19675) );
  nor_x1_sg U66031 ( .A(n6389), .B(n19677), .X(n19676) );
  nand_x1_sg U66032 ( .A(n19671), .B(n38683), .X(n19669) );
  nor_x1_sg U66033 ( .A(n6433), .B(n19671), .X(n19670) );
  nand_x1_sg U66034 ( .A(n19665), .B(n38681), .X(n19663) );
  nor_x1_sg U66035 ( .A(n6478), .B(n19665), .X(n19664) );
  nand_x1_sg U66036 ( .A(n19659), .B(n38679), .X(n19657) );
  nor_x1_sg U66037 ( .A(n6522), .B(n19659), .X(n19658) );
  nand_x1_sg U66038 ( .A(n19653), .B(n38677), .X(n19651) );
  nor_x1_sg U66039 ( .A(n6567), .B(n19653), .X(n19652) );
  nand_x1_sg U66040 ( .A(n19647), .B(n38689), .X(n19645) );
  nor_x1_sg U66041 ( .A(n6611), .B(n19647), .X(n19646) );
  nand_x1_sg U66042 ( .A(n21161), .B(n38666), .X(n21159) );
  nor_x1_sg U66043 ( .A(n6096), .B(n21161), .X(n21160) );
  nor_x1_sg U66044 ( .A(n46570), .B(n41253), .X(n6028) );
  nand_x1_sg U66045 ( .A(n39775), .B(n42092), .X(n17321) );
  nand_x1_sg U66046 ( .A(n39780), .B(n40067), .X(n18142) );
  nor_x1_sg U66047 ( .A(n41060), .B(n41861), .X(n7125) );
  nor_x1_sg U66048 ( .A(n41058), .B(n39855), .X(n7295) );
  nor_x1_sg U66049 ( .A(n41060), .B(n41983), .X(n6943) );
  nand_x1_sg U66050 ( .A(n40633), .B(n40244), .X(n8003) );
  nand_x1_sg U66051 ( .A(n40629), .B(n40247), .X(n8821) );
  nand_x1_sg U66052 ( .A(n40666), .B(n40254), .X(n9641) );
  nand_x1_sg U66053 ( .A(n40658), .B(n40259), .X(n10460) );
  nand_x1_sg U66054 ( .A(n40641), .B(n40264), .X(n11279) );
  nand_x1_sg U66055 ( .A(n40638), .B(n40268), .X(n12098) );
  nand_x1_sg U66056 ( .A(n40663), .B(n40274), .X(n12917) );
  nand_x1_sg U66057 ( .A(n40652), .B(n40280), .X(n13736) );
  nand_x1_sg U66058 ( .A(n40622), .B(n40282), .X(n14555) );
  nand_x1_sg U66059 ( .A(n40683), .B(n40289), .X(n15374) );
  nand_x1_sg U66060 ( .A(n40677), .B(n40294), .X(n16193) );
  nand_x1_sg U66061 ( .A(n40648), .B(n40238), .X(n17831) );
  nand_x1_sg U66062 ( .A(n40672), .B(n40298), .X(n18652) );
  nor_x1_sg U66063 ( .A(n39965), .B(n41915), .X(n7943) );
  nor_x1_sg U66064 ( .A(n39967), .B(n41916), .X(n8761) );
  nor_x1_sg U66065 ( .A(n39971), .B(n41907), .X(n9581) );
  nor_x1_sg U66066 ( .A(n39977), .B(n41909), .X(n10400) );
  nor_x1_sg U66067 ( .A(n41925), .B(n41913), .X(n11219) );
  nor_x1_sg U66068 ( .A(n39984), .B(n41914), .X(n12038) );
  nor_x1_sg U66069 ( .A(n39989), .B(n41908), .X(n12857) );
  nor_x1_sg U66070 ( .A(n39992), .B(n41911), .X(n13676) );
  nor_x1_sg U66071 ( .A(n39997), .B(n41917), .X(n14495) );
  nor_x1_sg U66072 ( .A(n40001), .B(n41904), .X(n15314) );
  nor_x1_sg U66073 ( .A(n40003), .B(n41905), .X(n16133) );
  nor_x1_sg U66074 ( .A(n38910), .B(n41912), .X(n17771) );
  nor_x1_sg U66075 ( .A(n40740), .B(n41906), .X(n18592) );
  nor_x1_sg U66076 ( .A(n39963), .B(n39894), .X(n8113) );
  nor_x1_sg U66077 ( .A(n39967), .B(n39861), .X(n8931) );
  nor_x1_sg U66078 ( .A(n41933), .B(n39858), .X(n9751) );
  nor_x1_sg U66079 ( .A(n41936), .B(n39864), .X(n10570) );
  nor_x1_sg U66080 ( .A(n39980), .B(n39867), .X(n11389) );
  nor_x1_sg U66081 ( .A(n39983), .B(n39870), .X(n12208) );
  nor_x1_sg U66082 ( .A(n41935), .B(n39873), .X(n13027) );
  nor_x1_sg U66083 ( .A(n41922), .B(n39876), .X(n13846) );
  nor_x1_sg U66084 ( .A(n39995), .B(n39879), .X(n14665) );
  nor_x1_sg U66085 ( .A(n41934), .B(n39897), .X(n15484) );
  nor_x1_sg U66086 ( .A(n40003), .B(n39882), .X(n16303) );
  nor_x1_sg U66087 ( .A(n40998), .B(n39887), .X(n17941) );
  nor_x1_sg U66088 ( .A(n40008), .B(n39891), .X(n18762) );
  nor_x1_sg U66089 ( .A(n39964), .B(n41984), .X(n7760) );
  nor_x1_sg U66090 ( .A(n39968), .B(n41985), .X(n8578) );
  nor_x1_sg U66091 ( .A(n41927), .B(n41979), .X(n9398) );
  nor_x1_sg U66092 ( .A(n39977), .B(n41980), .X(n10217) );
  nor_x1_sg U66093 ( .A(n39979), .B(n41981), .X(n11036) );
  nor_x1_sg U66094 ( .A(n39984), .B(n41982), .X(n11855) );
  nor_x1_sg U66095 ( .A(n39989), .B(n41975), .X(n12674) );
  nor_x1_sg U66096 ( .A(n41922), .B(n41976), .X(n13493) );
  nor_x1_sg U66097 ( .A(n39996), .B(n41977), .X(n14312) );
  nor_x1_sg U66098 ( .A(n40001), .B(n41978), .X(n15131) );
  nor_x1_sg U66099 ( .A(n41919), .B(n41972), .X(n15950) );
  nor_x1_sg U66100 ( .A(n41000), .B(n41973), .X(n17588) );
  nor_x1_sg U66101 ( .A(n41941), .B(n41974), .X(n18409) );
  nand_x1_sg U66102 ( .A(n39803), .B(n39957), .X(n7496) );
  nand_x1_sg U66103 ( .A(n40578), .B(n40565), .X(n17009) );
  nor_x1_sg U66104 ( .A(n38908), .B(n41860), .X(n16950) );
  nor_x1_sg U66105 ( .A(n38908), .B(n39885), .X(n17120) );
  nor_x1_sg U66106 ( .A(n40994), .B(n50525), .X(n16767) );
  nand_x1_sg U66107 ( .A(n7929), .B(n40245), .X(n7950) );
  nand_x1_sg U66108 ( .A(n8747), .B(n40247), .X(n8768) );
  nand_x1_sg U66109 ( .A(n41831), .B(n40254), .X(n9588) );
  nand_x1_sg U66110 ( .A(n10386), .B(n40260), .X(n10407) );
  nand_x1_sg U66111 ( .A(n11205), .B(n40264), .X(n11226) );
  nand_x1_sg U66112 ( .A(n12024), .B(n40269), .X(n12045) );
  nand_x1_sg U66113 ( .A(n41823), .B(n40275), .X(n12864) );
  nand_x1_sg U66114 ( .A(n41821), .B(n40278), .X(n13683) );
  nand_x1_sg U66115 ( .A(n41819), .B(n40282), .X(n14502) );
  nand_x1_sg U66116 ( .A(n15300), .B(n40290), .X(n15321) );
  nand_x1_sg U66117 ( .A(n41815), .B(n40294), .X(n16140) );
  nand_x1_sg U66118 ( .A(n17757), .B(n40240), .X(n17778) );
  nand_x1_sg U66119 ( .A(n18578), .B(n40299), .X(n18599) );
  nor_x1_sg U66120 ( .A(n26322), .B(n26323), .X(n26321) );
  nand_x1_sg U66121 ( .A(n41137), .B(n26324), .X(n26323) );
  nand_x1_sg U66122 ( .A(n40575), .B(n40164), .X(n7184) );
  nor_x1_sg U66123 ( .A(n42258), .B(n41254), .X(n6123) );
  nand_x1_sg U66124 ( .A(n40076), .B(n40566), .X(n17040) );
  nand_x1_sg U66125 ( .A(n39564), .B(n39206), .X(n8250) );
  nand_x1_sg U66126 ( .A(n39567), .B(n39498), .X(n9068) );
  nand_x1_sg U66127 ( .A(n39570), .B(n39208), .X(n9888) );
  nand_x1_sg U66128 ( .A(n39573), .B(n39209), .X(n10707) );
  nand_x1_sg U66129 ( .A(n39576), .B(n39495), .X(n11526) );
  nand_x1_sg U66130 ( .A(n39579), .B(n39211), .X(n12345) );
  nand_x1_sg U66131 ( .A(n39582), .B(n39493), .X(n13164) );
  nand_x1_sg U66132 ( .A(n39585), .B(n39492), .X(n13983) );
  nand_x1_sg U66133 ( .A(n39588), .B(n39491), .X(n14802) );
  nand_x1_sg U66134 ( .A(n39591), .B(n39215), .X(n15621) );
  nand_x1_sg U66135 ( .A(n39594), .B(n39489), .X(n16440) );
  nand_x1_sg U66136 ( .A(n39599), .B(n41805), .X(n18078) );
  nand_x1_sg U66137 ( .A(n39597), .B(n39487), .X(n18899) );
  nand_x1_sg U66138 ( .A(n40235), .B(n40163), .X(n7132) );
  nand_x1_sg U66139 ( .A(n40230), .B(n40565), .X(n16957) );
  inv_x1_sg U66140 ( .A(n42295), .X(n46549) );
  inv_x1_sg U66141 ( .A(n42284), .X(n46375) );
  inv_x1_sg U66142 ( .A(n42296), .X(n46334) );
  inv_x1_sg U66143 ( .A(n42297), .X(n46288) );
  inv_x1_sg U66144 ( .A(n42231), .X(n46243) );
  inv_x1_sg U66145 ( .A(n42299), .X(n46197) );
  inv_x1_sg U66146 ( .A(n42232), .X(n46152) );
  inv_x1_sg U66147 ( .A(n42234), .X(n46106) );
  inv_x1_sg U66148 ( .A(n42301), .X(n46061) );
  inv_x1_sg U66149 ( .A(n42233), .X(n46015) );
  inv_x1_sg U66150 ( .A(n42300), .X(n45970) );
  inv_x1_sg U66151 ( .A(n42294), .X(n46337) );
  inv_x1_sg U66152 ( .A(n42293), .X(n46291) );
  inv_x1_sg U66153 ( .A(n42292), .X(n46246) );
  inv_x1_sg U66154 ( .A(n42291), .X(n46200) );
  inv_x1_sg U66155 ( .A(n42286), .X(n46155) );
  inv_x1_sg U66156 ( .A(n42290), .X(n46109) );
  inv_x1_sg U66157 ( .A(n42289), .X(n46064) );
  inv_x1_sg U66158 ( .A(n42288), .X(n46018) );
  inv_x1_sg U66159 ( .A(n42287), .X(n45973) );
  inv_x1_sg U66160 ( .A(n42282), .X(n46340) );
  inv_x1_sg U66161 ( .A(n42281), .X(n46294) );
  inv_x1_sg U66162 ( .A(n42280), .X(n46249) );
  inv_x1_sg U66163 ( .A(n42279), .X(n46203) );
  inv_x1_sg U66164 ( .A(n42268), .X(n46158) );
  inv_x1_sg U66165 ( .A(n42278), .X(n46112) );
  inv_x1_sg U66166 ( .A(n42277), .X(n46067) );
  inv_x1_sg U66167 ( .A(n42230), .X(n46021) );
  inv_x1_sg U66168 ( .A(n42276), .X(n45976) );
  inv_x1_sg U66169 ( .A(n42269), .X(n46194) );
  inv_x1_sg U66170 ( .A(n42267), .X(n46149) );
  inv_x1_sg U66171 ( .A(n42266), .X(n46103) );
  inv_x1_sg U66172 ( .A(n42265), .X(n46058) );
  inv_x1_sg U66173 ( .A(n42264), .X(n46012) );
  inv_x1_sg U66174 ( .A(n42263), .X(n45967) );
  inv_x1_sg U66175 ( .A(n42270), .X(n46240) );
  inv_x1_sg U66176 ( .A(n42271), .X(n46285) );
  inv_x1_sg U66177 ( .A(n42272), .X(n46331) );
  inv_x1_sg U66178 ( .A(n42273), .X(n46372) );
  inv_x1_sg U66179 ( .A(n42274), .X(n46420) );
  inv_x1_sg U66180 ( .A(n42275), .X(n46467) );
  inv_x1_sg U66181 ( .A(n42283), .X(n46557) );
  nor_x1_sg U66182 ( .A(n7094), .B(n41306), .X(n22625) );
  nor_x1_sg U66183 ( .A(n7912), .B(n41195), .X(n22890) );
  nor_x1_sg U66184 ( .A(n8730), .B(n41188), .X(n23167) );
  nor_x1_sg U66185 ( .A(n9550), .B(n41183), .X(n23447) );
  nor_x1_sg U66186 ( .A(n10369), .B(n41177), .X(n23726) );
  nor_x1_sg U66187 ( .A(n41791), .B(n41175), .X(n24005) );
  nor_x1_sg U66188 ( .A(n41793), .B(n41168), .X(n24284) );
  nor_x1_sg U66189 ( .A(n12826), .B(n41163), .X(n24563) );
  nor_x1_sg U66190 ( .A(n41797), .B(n41158), .X(n24841) );
  nor_x1_sg U66191 ( .A(n14464), .B(n41155), .X(n25120) );
  nor_x1_sg U66192 ( .A(n41801), .B(n39240), .X(n25399) );
  nor_x1_sg U66193 ( .A(n16102), .B(n41145), .X(n25678) );
  nor_x1_sg U66194 ( .A(n41805), .B(n41137), .X(n26223) );
  nor_x1_sg U66195 ( .A(n18561), .B(n41132), .X(n26515) );
  nand_x1_sg U66196 ( .A(n46929), .B(n39205), .X(n7176) );
  nand_x1_sg U66197 ( .A(n47221), .B(n7912), .X(n7995) );
  nand_x1_sg U66198 ( .A(n47506), .B(n8730), .X(n8813) );
  nand_x1_sg U66199 ( .A(n47791), .B(n9550), .X(n9633) );
  nand_x1_sg U66200 ( .A(n48076), .B(n10369), .X(n10452) );
  nand_x1_sg U66201 ( .A(n48361), .B(n11188), .X(n11271) );
  nand_x1_sg U66202 ( .A(n48646), .B(n12007), .X(n12090) );
  nand_x1_sg U66203 ( .A(n48932), .B(n12826), .X(n12909) );
  nand_x1_sg U66204 ( .A(n49219), .B(n13645), .X(n13728) );
  nand_x1_sg U66205 ( .A(n49505), .B(n14464), .X(n14547) );
  nand_x1_sg U66206 ( .A(n49791), .B(n15283), .X(n15366) );
  nand_x1_sg U66207 ( .A(n50077), .B(n16102), .X(n16185) );
  nand_x1_sg U66208 ( .A(n50651), .B(n17740), .X(n17823) );
  nand_x1_sg U66209 ( .A(n50938), .B(n18561), .X(n18644) );
  nand_x1_sg U66210 ( .A(n39678), .B(n39956), .X(n7636) );
  nand_x1_sg U66211 ( .A(n42311), .B(n40157), .X(n8454) );
  nand_x1_sg U66212 ( .A(n42310), .B(n40359), .X(n9272) );
  nand_x1_sg U66213 ( .A(n42309), .B(n40355), .X(n10092) );
  nand_x1_sg U66214 ( .A(n10272), .B(n40351), .X(n10911) );
  nand_x1_sg U66215 ( .A(n42308), .B(n40347), .X(n11730) );
  nand_x1_sg U66216 ( .A(n42307), .B(n40327), .X(n12549) );
  nand_x1_sg U66217 ( .A(n42306), .B(n40339), .X(n13368) );
  nand_x1_sg U66218 ( .A(n13548), .B(n40335), .X(n14187) );
  nand_x1_sg U66219 ( .A(n42305), .B(n40343), .X(n15006) );
  nand_x1_sg U66220 ( .A(n42304), .B(n40319), .X(n15825) );
  nand_x1_sg U66221 ( .A(n42303), .B(n40323), .X(n16644) );
  nand_x1_sg U66222 ( .A(n17643), .B(n40068), .X(n18282) );
  nand_x1_sg U66223 ( .A(n18464), .B(n40331), .X(n19103) );
  nand_x1_sg U66224 ( .A(n40134), .B(n40634), .X(n8262) );
  nand_x1_sg U66225 ( .A(n40136), .B(n40627), .X(n9080) );
  nand_x1_sg U66226 ( .A(n40138), .B(n40666), .X(n9900) );
  nand_x1_sg U66227 ( .A(n40140), .B(n40659), .X(n10719) );
  nand_x1_sg U66228 ( .A(n40142), .B(n40644), .X(n11538) );
  nand_x1_sg U66229 ( .A(n40144), .B(n40636), .X(n12357) );
  nand_x1_sg U66230 ( .A(n40146), .B(n40662), .X(n13176) );
  nand_x1_sg U66231 ( .A(n40148), .B(n40651), .X(n13995) );
  nand_x1_sg U66232 ( .A(n40150), .B(n40623), .X(n14814) );
  nand_x1_sg U66233 ( .A(n40152), .B(n40684), .X(n15633) );
  nand_x1_sg U66234 ( .A(n40154), .B(n40676), .X(n16452) );
  nand_x1_sg U66235 ( .A(n40159), .B(n40648), .X(n18090) );
  nand_x1_sg U66236 ( .A(n40156), .B(n40671), .X(n18911) );
  nand_x1_sg U66237 ( .A(n41057), .B(n39956), .X(n6825) );
  nand_x1_sg U66238 ( .A(n17107), .B(n40608), .X(n17106) );
  nand_x1_sg U66239 ( .A(n17108), .B(n17110), .X(n17105) );
  nor_x1_sg U66240 ( .A(n17108), .B(n42337), .X(n17107) );
  nand_x1_sg U66241 ( .A(n7283), .B(n7285), .X(n7280) );
  nor_x1_sg U66242 ( .A(n7283), .B(n42369), .X(n7282) );
  inv_x1_sg U66243 ( .A(n27977), .X(n45000) );
  inv_x1_sg U66244 ( .A(n27808), .X(n45003) );
  inv_x1_sg U66245 ( .A(n27622), .X(n45006) );
  inv_x1_sg U66246 ( .A(n27419), .X(n45009) );
  inv_x1_sg U66247 ( .A(n21437), .X(n45814) );
  inv_x1_sg U66248 ( .A(n28468), .X(n44987) );
  inv_x1_sg U66249 ( .A(n28988), .X(n44978) );
  inv_x1_sg U66250 ( .A(n27197), .X(n45012) );
  inv_x1_sg U66251 ( .A(n28374), .X(n44990) );
  inv_x1_sg U66252 ( .A(n28817), .X(n44981) );
  inv_x1_sg U66253 ( .A(n26958), .X(n45015) );
  inv_x1_sg U66254 ( .A(n28261), .X(n44993) );
  inv_x1_sg U66255 ( .A(n28629), .X(n44984) );
  nand_x1_sg U66256 ( .A(n40631), .B(n7929), .X(n8076) );
  nand_x1_sg U66257 ( .A(n40628), .B(n8747), .X(n8894) );
  nand_x1_sg U66258 ( .A(n40669), .B(n9567), .X(n9714) );
  nand_x1_sg U66259 ( .A(n40658), .B(n10386), .X(n10533) );
  nand_x1_sg U66260 ( .A(n40641), .B(n11205), .X(n11352) );
  nand_x1_sg U66261 ( .A(n40639), .B(n12024), .X(n12171) );
  nand_x1_sg U66262 ( .A(n40663), .B(n41823), .X(n12990) );
  nand_x1_sg U66263 ( .A(n40651), .B(n13662), .X(n13809) );
  nand_x1_sg U66264 ( .A(n40621), .B(n41819), .X(n14628) );
  nand_x1_sg U66265 ( .A(n40683), .B(n15300), .X(n15447) );
  nand_x1_sg U66266 ( .A(n40676), .B(n41815), .X(n16266) );
  nand_x1_sg U66267 ( .A(n40647), .B(n17757), .X(n17904) );
  nand_x1_sg U66268 ( .A(n40671), .B(n41813), .X(n18725) );
  nand_x1_sg U66269 ( .A(n8185), .B(n39532), .X(n8184) );
  nand_x1_sg U66270 ( .A(n8186), .B(n8187), .X(n8183) );
  nor_x1_sg U66271 ( .A(n39963), .B(n8186), .X(n8185) );
  nand_x1_sg U66272 ( .A(n9003), .B(n39533), .X(n9002) );
  nand_x1_sg U66273 ( .A(n9004), .B(n9005), .X(n9001) );
  nor_x1_sg U66274 ( .A(n41940), .B(n9004), .X(n9003) );
  nand_x1_sg U66275 ( .A(n9823), .B(n39534), .X(n9822) );
  nand_x1_sg U66276 ( .A(n9824), .B(n9825), .X(n9821) );
  nor_x1_sg U66277 ( .A(n39973), .B(n9824), .X(n9823) );
  nand_x1_sg U66278 ( .A(n10642), .B(n39535), .X(n10641) );
  nand_x1_sg U66279 ( .A(n10643), .B(n10644), .X(n10640) );
  nor_x1_sg U66280 ( .A(n39975), .B(n10643), .X(n10642) );
  nand_x1_sg U66281 ( .A(n11461), .B(n39536), .X(n11460) );
  nand_x1_sg U66282 ( .A(n11462), .B(n11463), .X(n11459) );
  nor_x1_sg U66283 ( .A(n39979), .B(n11462), .X(n11461) );
  nand_x1_sg U66284 ( .A(n12280), .B(n39537), .X(n12279) );
  nand_x1_sg U66285 ( .A(n12281), .B(n12282), .X(n12278) );
  nor_x1_sg U66286 ( .A(n39983), .B(n12281), .X(n12280) );
  nand_x1_sg U66287 ( .A(n13099), .B(n39538), .X(n13098) );
  nand_x1_sg U66288 ( .A(n13100), .B(n13101), .X(n13097) );
  nor_x1_sg U66289 ( .A(n39987), .B(n13100), .X(n13099) );
  nand_x1_sg U66290 ( .A(n13918), .B(n39539), .X(n13917) );
  nand_x1_sg U66291 ( .A(n13919), .B(n13920), .X(n13916) );
  nor_x1_sg U66292 ( .A(n39991), .B(n13919), .X(n13918) );
  nand_x1_sg U66293 ( .A(n14737), .B(n39540), .X(n14736) );
  nand_x1_sg U66294 ( .A(n14738), .B(n14739), .X(n14735) );
  nor_x1_sg U66295 ( .A(n41932), .B(n14738), .X(n14737) );
  nand_x1_sg U66296 ( .A(n15556), .B(n39541), .X(n15555) );
  nand_x1_sg U66297 ( .A(n15557), .B(n15558), .X(n15554) );
  nor_x1_sg U66298 ( .A(n39999), .B(n15557), .X(n15556) );
  nand_x1_sg U66299 ( .A(n16375), .B(n39542), .X(n16374) );
  nand_x1_sg U66300 ( .A(n16376), .B(n16377), .X(n16373) );
  nor_x1_sg U66301 ( .A(n40005), .B(n16376), .X(n16375) );
  nand_x1_sg U66302 ( .A(n17193), .B(n17194), .X(n17190) );
  nor_x1_sg U66303 ( .A(n40995), .B(n17193), .X(n17192) );
  nand_x1_sg U66304 ( .A(n18013), .B(n39543), .X(n18012) );
  nand_x1_sg U66305 ( .A(n18014), .B(n18015), .X(n18011) );
  nor_x1_sg U66306 ( .A(n41001), .B(n18014), .X(n18013) );
  nand_x1_sg U66307 ( .A(n18834), .B(n39544), .X(n18833) );
  nand_x1_sg U66308 ( .A(n18835), .B(n18836), .X(n18832) );
  nor_x1_sg U66309 ( .A(n40009), .B(n18835), .X(n18834) );
  nand_x1_sg U66310 ( .A(n7367), .B(n6991), .X(n7366) );
  nand_x1_sg U66311 ( .A(n7368), .B(n7369), .X(n7365) );
  nor_x1_sg U66312 ( .A(n41059), .B(n7368), .X(n7367) );
  nand_x1_sg U66313 ( .A(n40993), .B(n40069), .X(n16649) );
  nand_x1_sg U66314 ( .A(n7296), .B(n7299), .X(n7297) );
  nor_x1_sg U66315 ( .A(n7299), .B(n7296), .X(n7298) );
  nand_x1_sg U66316 ( .A(n8114), .B(n8117), .X(n8115) );
  nor_x1_sg U66317 ( .A(n8117), .B(n8114), .X(n8116) );
  nand_x1_sg U66318 ( .A(n8932), .B(n8935), .X(n8933) );
  nor_x1_sg U66319 ( .A(n8935), .B(n8932), .X(n8934) );
  nand_x1_sg U66320 ( .A(n9752), .B(n9755), .X(n9753) );
  nor_x1_sg U66321 ( .A(n9755), .B(n9752), .X(n9754) );
  nand_x1_sg U66322 ( .A(n10571), .B(n10574), .X(n10572) );
  nor_x1_sg U66323 ( .A(n10574), .B(n10571), .X(n10573) );
  nand_x1_sg U66324 ( .A(n11390), .B(n11393), .X(n11391) );
  nor_x1_sg U66325 ( .A(n11393), .B(n11390), .X(n11392) );
  nand_x1_sg U66326 ( .A(n12209), .B(n12212), .X(n12210) );
  nor_x1_sg U66327 ( .A(n12212), .B(n12209), .X(n12211) );
  nand_x1_sg U66328 ( .A(n13028), .B(n13031), .X(n13029) );
  nor_x1_sg U66329 ( .A(n13031), .B(n13028), .X(n13030) );
  nand_x1_sg U66330 ( .A(n13847), .B(n13850), .X(n13848) );
  nor_x1_sg U66331 ( .A(n13850), .B(n13847), .X(n13849) );
  nand_x1_sg U66332 ( .A(n14666), .B(n14669), .X(n14667) );
  nor_x1_sg U66333 ( .A(n14669), .B(n14666), .X(n14668) );
  nand_x1_sg U66334 ( .A(n15485), .B(n15488), .X(n15486) );
  nor_x1_sg U66335 ( .A(n15488), .B(n15485), .X(n15487) );
  nand_x1_sg U66336 ( .A(n16304), .B(n16307), .X(n16305) );
  nor_x1_sg U66337 ( .A(n16307), .B(n16304), .X(n16306) );
  nand_x1_sg U66338 ( .A(n17121), .B(n17124), .X(n17122) );
  nor_x1_sg U66339 ( .A(n17124), .B(n17121), .X(n17123) );
  nand_x1_sg U66340 ( .A(n17942), .B(n17945), .X(n17943) );
  nor_x1_sg U66341 ( .A(n17945), .B(n17942), .X(n17944) );
  nand_x1_sg U66342 ( .A(n18763), .B(n18766), .X(n18764) );
  nor_x1_sg U66343 ( .A(n18766), .B(n18763), .X(n18765) );
  nand_x1_sg U66344 ( .A(n7473), .B(n7472), .X(n7470) );
  nor_x1_sg U66345 ( .A(n7472), .B(n7473), .X(n7471) );
  nand_x1_sg U66346 ( .A(n17298), .B(n17297), .X(n17295) );
  nor_x1_sg U66347 ( .A(n17297), .B(n17298), .X(n17296) );
  nor_x1_sg U66348 ( .A(n7947), .B(n7944), .X(n7946) );
  nor_x1_sg U66349 ( .A(n8765), .B(n8762), .X(n8764) );
  nor_x1_sg U66350 ( .A(n9585), .B(n9582), .X(n9584) );
  nor_x1_sg U66351 ( .A(n10404), .B(n10401), .X(n10403) );
  nor_x1_sg U66352 ( .A(n11223), .B(n11220), .X(n11222) );
  nor_x1_sg U66353 ( .A(n12042), .B(n12039), .X(n12041) );
  nor_x1_sg U66354 ( .A(n12861), .B(n12858), .X(n12860) );
  nor_x1_sg U66355 ( .A(n13680), .B(n13677), .X(n13679) );
  nand_x1_sg U66356 ( .A(n14496), .B(n14499), .X(n14497) );
  nor_x1_sg U66357 ( .A(n14499), .B(n14496), .X(n14498) );
  nand_x1_sg U66358 ( .A(n15315), .B(n15318), .X(n15316) );
  nor_x1_sg U66359 ( .A(n15318), .B(n15315), .X(n15317) );
  nand_x1_sg U66360 ( .A(n16134), .B(n16137), .X(n16135) );
  nor_x1_sg U66361 ( .A(n16137), .B(n16134), .X(n16136) );
  nand_x1_sg U66362 ( .A(n17772), .B(n17775), .X(n17773) );
  nor_x1_sg U66363 ( .A(n17775), .B(n17772), .X(n17774) );
  nand_x1_sg U66364 ( .A(n18593), .B(n18596), .X(n18594) );
  nor_x1_sg U66365 ( .A(n18596), .B(n18593), .X(n18595) );
  nand_x1_sg U66366 ( .A(n7126), .B(n7129), .X(n7127) );
  nor_x1_sg U66367 ( .A(n7129), .B(n7126), .X(n7128) );
  nand_x1_sg U66368 ( .A(n16951), .B(n16954), .X(n16952) );
  nor_x1_sg U66369 ( .A(n16954), .B(n16951), .X(n16953) );
  nand_x1_sg U66370 ( .A(n8291), .B(n8290), .X(n8288) );
  nor_x1_sg U66371 ( .A(n8290), .B(n8291), .X(n8289) );
  nand_x1_sg U66372 ( .A(n9109), .B(n9108), .X(n9106) );
  nor_x1_sg U66373 ( .A(n9108), .B(n9109), .X(n9107) );
  nand_x1_sg U66374 ( .A(n9929), .B(n9928), .X(n9926) );
  nor_x1_sg U66375 ( .A(n9928), .B(n9929), .X(n9927) );
  nand_x1_sg U66376 ( .A(n10748), .B(n10747), .X(n10745) );
  nor_x1_sg U66377 ( .A(n10747), .B(n10748), .X(n10746) );
  nand_x1_sg U66378 ( .A(n11567), .B(n11566), .X(n11564) );
  nor_x1_sg U66379 ( .A(n11566), .B(n11567), .X(n11565) );
  nand_x1_sg U66380 ( .A(n12386), .B(n12385), .X(n12383) );
  nor_x1_sg U66381 ( .A(n12385), .B(n12386), .X(n12384) );
  nand_x1_sg U66382 ( .A(n13205), .B(n13204), .X(n13202) );
  nor_x1_sg U66383 ( .A(n13204), .B(n13205), .X(n13203) );
  nand_x1_sg U66384 ( .A(n14024), .B(n14023), .X(n14021) );
  nor_x1_sg U66385 ( .A(n14023), .B(n14024), .X(n14022) );
  nand_x1_sg U66386 ( .A(n14843), .B(n14842), .X(n14840) );
  nor_x1_sg U66387 ( .A(n14842), .B(n14843), .X(n14841) );
  nand_x1_sg U66388 ( .A(n15662), .B(n15661), .X(n15659) );
  nor_x1_sg U66389 ( .A(n15661), .B(n15662), .X(n15660) );
  nand_x1_sg U66390 ( .A(n16481), .B(n16480), .X(n16478) );
  nor_x1_sg U66391 ( .A(n16480), .B(n16481), .X(n16479) );
  nand_x1_sg U66392 ( .A(n18119), .B(n18118), .X(n18116) );
  nor_x1_sg U66393 ( .A(n18118), .B(n18119), .X(n18117) );
  nand_x1_sg U66394 ( .A(n18940), .B(n18939), .X(n18937) );
  nor_x1_sg U66395 ( .A(n18939), .B(n18940), .X(n18938) );
  nand_x1_sg U66396 ( .A(n7761), .B(n8450), .X(n8448) );
  nor_x1_sg U66397 ( .A(n8450), .B(n7761), .X(n8449) );
  nand_x1_sg U66398 ( .A(n8579), .B(n9268), .X(n9266) );
  nor_x1_sg U66399 ( .A(n9268), .B(n8579), .X(n9267) );
  nand_x1_sg U66400 ( .A(n9399), .B(n10088), .X(n10086) );
  nor_x1_sg U66401 ( .A(n10088), .B(n9399), .X(n10087) );
  nand_x1_sg U66402 ( .A(n10218), .B(n10907), .X(n10905) );
  nor_x1_sg U66403 ( .A(n10907), .B(n10218), .X(n10906) );
  nand_x1_sg U66404 ( .A(n11037), .B(n11726), .X(n11724) );
  nor_x1_sg U66405 ( .A(n11726), .B(n11037), .X(n11725) );
  nand_x1_sg U66406 ( .A(n11856), .B(n12545), .X(n12543) );
  nor_x1_sg U66407 ( .A(n12545), .B(n11856), .X(n12544) );
  nand_x1_sg U66408 ( .A(n12675), .B(n13364), .X(n13362) );
  nor_x1_sg U66409 ( .A(n13364), .B(n12675), .X(n13363) );
  nand_x1_sg U66410 ( .A(n13494), .B(n14183), .X(n14181) );
  nor_x1_sg U66411 ( .A(n14183), .B(n13494), .X(n14182) );
  nand_x1_sg U66412 ( .A(n14313), .B(n15002), .X(n15000) );
  nor_x1_sg U66413 ( .A(n15002), .B(n14313), .X(n15001) );
  nand_x1_sg U66414 ( .A(n15132), .B(n15821), .X(n15819) );
  nor_x1_sg U66415 ( .A(n15821), .B(n15132), .X(n15820) );
  nand_x1_sg U66416 ( .A(n15951), .B(n16640), .X(n16638) );
  nor_x1_sg U66417 ( .A(n16640), .B(n15951), .X(n16639) );
  nand_x1_sg U66418 ( .A(n17589), .B(n18278), .X(n18276) );
  nor_x1_sg U66419 ( .A(n18278), .B(n17589), .X(n18277) );
  nand_x1_sg U66420 ( .A(n18410), .B(n19099), .X(n19097) );
  nor_x1_sg U66421 ( .A(n19099), .B(n18410), .X(n19098) );
  nand_x1_sg U66422 ( .A(n16768), .B(n17457), .X(n17455) );
  nor_x1_sg U66423 ( .A(n17457), .B(n16768), .X(n17456) );
  nand_x1_sg U66424 ( .A(n6944), .B(n7632), .X(n7630) );
  nor_x1_sg U66425 ( .A(n7632), .B(n6944), .X(n7631) );
  nand_x1_sg U66426 ( .A(n40073), .B(n40566), .X(n16982) );
  nand_x1_sg U66427 ( .A(n39932), .B(n40566), .X(n17128) );
  nand_x1_sg U66428 ( .A(n40573), .B(n40235), .X(n7257) );
  nand_x1_sg U66429 ( .A(n40579), .B(n40229), .X(n17082) );
  inv_x1_sg U66430 ( .A(n28123), .X(n44969) );
  nand_x1_sg U66431 ( .A(n39349), .B(n39502), .X(n22639) );
  nand_x1_sg U66432 ( .A(n42345), .B(n40633), .X(n8423) );
  nand_x1_sg U66433 ( .A(n42344), .B(n40626), .X(n9241) );
  nand_x1_sg U66434 ( .A(n42355), .B(n40669), .X(n10061) );
  nand_x1_sg U66435 ( .A(n42354), .B(n40659), .X(n10880) );
  nand_x1_sg U66436 ( .A(n42353), .B(n40644), .X(n11699) );
  nand_x1_sg U66437 ( .A(n42352), .B(n40637), .X(n12518) );
  nand_x1_sg U66438 ( .A(n42351), .B(n40664), .X(n13337) );
  nand_x1_sg U66439 ( .A(n42350), .B(n40654), .X(n14156) );
  nand_x1_sg U66440 ( .A(n42349), .B(n40623), .X(n14975) );
  nand_x1_sg U66441 ( .A(n42348), .B(n40684), .X(n15794) );
  nand_x1_sg U66442 ( .A(n42347), .B(n40679), .X(n16613) );
  nand_x1_sg U66443 ( .A(n42336), .B(n40580), .X(n17430) );
  nand_x1_sg U66444 ( .A(n42356), .B(n40647), .X(n18251) );
  nand_x1_sg U66445 ( .A(n42346), .B(n40674), .X(n19072) );
  nand_x1_sg U66446 ( .A(n39812), .B(n40634), .X(n8044) );
  nand_x1_sg U66447 ( .A(n39831), .B(n40629), .X(n8862) );
  nand_x1_sg U66448 ( .A(n41877), .B(n40667), .X(n9682) );
  nand_x1_sg U66449 ( .A(n39815), .B(n40656), .X(n10501) );
  nand_x1_sg U66450 ( .A(n39833), .B(n40643), .X(n11320) );
  nand_x1_sg U66451 ( .A(n41883), .B(n40637), .X(n12139) );
  nand_x1_sg U66452 ( .A(n41895), .B(n40661), .X(n12958) );
  nand_x1_sg U66453 ( .A(n39840), .B(n40654), .X(n13777) );
  nand_x1_sg U66454 ( .A(n41879), .B(n40624), .X(n14596) );
  nand_x1_sg U66455 ( .A(n39848), .B(n40681), .X(n15415) );
  nand_x1_sg U66456 ( .A(n39821), .B(n40679), .X(n16234) );
  nand_x1_sg U66457 ( .A(n41889), .B(n40649), .X(n17872) );
  nand_x1_sg U66458 ( .A(n41891), .B(n40674), .X(n18693) );
  nand_x1_sg U66459 ( .A(n39807), .B(n40070), .X(n17461) );
  nand_x1_sg U66460 ( .A(n39773), .B(n40573), .X(n7605) );
  nand_x1_sg U66461 ( .A(n39810), .B(n40576), .X(n7225) );
  nand_x1_sg U66462 ( .A(n40610), .B(n40580), .X(n17050) );
  nor_x1_sg U66463 ( .A(n22693), .B(n22694), .X(n22692) );
  nor_x1_sg U66464 ( .A(n39660), .B(n7633), .X(n22694) );
  nor_x1_sg U66465 ( .A(n22695), .B(n39349), .X(n22693) );
  nand_x1_sg U66466 ( .A(n38944), .B(n41283), .X(n5779) );
  nand_x1_sg U66467 ( .A(n40632), .B(n8060), .X(n8057) );
  nand_x1_sg U66468 ( .A(n40627), .B(n8878), .X(n8875) );
  nand_x1_sg U66469 ( .A(n40668), .B(n9698), .X(n9695) );
  nand_x1_sg U66470 ( .A(n40657), .B(n10517), .X(n10514) );
  nand_x1_sg U66471 ( .A(n40643), .B(n11336), .X(n11333) );
  nand_x1_sg U66472 ( .A(n40638), .B(n12155), .X(n12152) );
  nand_x1_sg U66473 ( .A(n40662), .B(n12974), .X(n12971) );
  nand_x1_sg U66474 ( .A(n40652), .B(n13793), .X(n13790) );
  nand_x1_sg U66475 ( .A(n40624), .B(n14612), .X(n14609) );
  nand_x1_sg U66476 ( .A(n40683), .B(n15431), .X(n15428) );
  nand_x1_sg U66477 ( .A(n40678), .B(n16250), .X(n16247) );
  nand_x1_sg U66478 ( .A(n40649), .B(n17888), .X(n17885) );
  nand_x1_sg U66479 ( .A(n40673), .B(n18709), .X(n18706) );
  nand_x1_sg U66480 ( .A(n39499), .B(n39519), .X(n8379) );
  nand_x1_sg U66481 ( .A(n8730), .B(n39518), .X(n9197) );
  nand_x1_sg U66482 ( .A(n9550), .B(n39524), .X(n10017) );
  nand_x1_sg U66483 ( .A(n10369), .B(n39523), .X(n10836) );
  nand_x1_sg U66484 ( .A(n39495), .B(n39522), .X(n11655) );
  nand_x1_sg U66485 ( .A(n39494), .B(n39521), .X(n12474) );
  nand_x1_sg U66486 ( .A(n12826), .B(n39528), .X(n13293) );
  nand_x1_sg U66487 ( .A(n13645), .B(n39527), .X(n14112) );
  nand_x1_sg U66488 ( .A(n14464), .B(n39526), .X(n14931) );
  nand_x1_sg U66489 ( .A(n41801), .B(n39525), .X(n15750) );
  nand_x1_sg U66490 ( .A(n16102), .B(n39531), .X(n16569) );
  nand_x1_sg U66491 ( .A(n39217), .B(n39530), .X(n18207) );
  nand_x1_sg U66492 ( .A(n18561), .B(n39529), .X(n19028) );
  inv_x1_sg U66493 ( .A(n7015), .X(n47074) );
  inv_x1_sg U66494 ( .A(n7833), .X(n47360) );
  inv_x1_sg U66495 ( .A(n8651), .X(n47645) );
  inv_x1_sg U66496 ( .A(n9471), .X(n47930) );
  inv_x1_sg U66497 ( .A(n10290), .X(n48215) );
  inv_x1_sg U66498 ( .A(n11109), .X(n48500) );
  inv_x1_sg U66499 ( .A(n11928), .X(n48785) );
  inv_x1_sg U66500 ( .A(n12747), .X(n49072) );
  inv_x1_sg U66501 ( .A(n13566), .X(n49358) );
  inv_x1_sg U66502 ( .A(n14385), .X(n49644) );
  inv_x1_sg U66503 ( .A(n15204), .X(n49930) );
  inv_x1_sg U66504 ( .A(n16023), .X(n50216) );
  inv_x1_sg U66505 ( .A(n16840), .X(n50522) );
  inv_x1_sg U66506 ( .A(n17661), .X(n50790) );
  inv_x1_sg U66507 ( .A(n18482), .X(n51077) );
  inv_x1_sg U66508 ( .A(n6051), .X(n46552) );
  inv_x1_sg U66509 ( .A(n6134), .X(n46479) );
  inv_x1_sg U66510 ( .A(n6193), .X(n46423) );
  inv_x1_sg U66511 ( .A(n6147), .X(n46470) );
  inv_x1_sg U66512 ( .A(n6101), .X(n46507) );
  inv_x1_sg U66513 ( .A(n6691), .X(n45923) );
  inv_x1_sg U66514 ( .A(n6102), .X(n46508) );
  inv_x1_sg U66515 ( .A(n6659), .X(n45926) );
  inv_x1_sg U66516 ( .A(n6674), .X(n45929) );
  inv_x1_sg U66517 ( .A(n22401), .X(n45127) );
  inv_x1_sg U66518 ( .A(n22354), .X(n45172) );
  inv_x1_sg U66519 ( .A(n22306), .X(n45218) );
  inv_x1_sg U66520 ( .A(n22259), .X(n45263) );
  inv_x1_sg U66521 ( .A(n22211), .X(n45308) );
  inv_x1_sg U66522 ( .A(n22164), .X(n45353) );
  inv_x1_sg U66523 ( .A(n22116), .X(n45399) );
  inv_x1_sg U66524 ( .A(n6162), .X(n46430) );
  inv_x1_sg U66525 ( .A(n6216), .X(n46385) );
  nand_x1_sg U66526 ( .A(n40575), .B(n7241), .X(n7238) );
  nand_x1_sg U66527 ( .A(n40581), .B(n17066), .X(n17063) );
  inv_x1_sg U66528 ( .A(n21170), .X(n46537) );
  nand_x1_sg U66529 ( .A(n38984), .B(n39108), .X(n8456) );
  nand_x1_sg U66530 ( .A(n42185), .B(n40244), .X(n8034) );
  nand_x1_sg U66531 ( .A(n40136), .B(n40247), .X(n8852) );
  nand_x1_sg U66532 ( .A(n40138), .B(n40253), .X(n9672) );
  nand_x1_sg U66533 ( .A(n40140), .B(n40259), .X(n10491) );
  nand_x1_sg U66534 ( .A(n40142), .B(n40265), .X(n11310) );
  nand_x1_sg U66535 ( .A(n40144), .B(n40268), .X(n12129) );
  nand_x1_sg U66536 ( .A(n40146), .B(n40274), .X(n12948) );
  nand_x1_sg U66537 ( .A(n40148), .B(n40277), .X(n13767) );
  nand_x1_sg U66538 ( .A(n40150), .B(n40282), .X(n14586) );
  nand_x1_sg U66539 ( .A(n40151), .B(n40289), .X(n15405) );
  nand_x1_sg U66540 ( .A(n40154), .B(n40295), .X(n16224) );
  nand_x1_sg U66541 ( .A(n40160), .B(n40239), .X(n17862) );
  nand_x1_sg U66542 ( .A(n42164), .B(n40298), .X(n18683) );
  nor_x1_sg U66543 ( .A(n22873), .B(n22874), .X(n22872) );
  nor_x1_sg U66544 ( .A(n22876), .B(n40370), .X(n22871) );
  nor_x1_sg U66545 ( .A(n40063), .B(n22875), .X(n22874) );
  nor_x1_sg U66546 ( .A(n23135), .B(n23136), .X(n23134) );
  nor_x1_sg U66547 ( .A(n23139), .B(n40457), .X(n23133) );
  nor_x1_sg U66548 ( .A(n40504), .B(n23138), .X(n23136) );
  nor_x1_sg U66549 ( .A(n23709), .B(n23710), .X(n23708) );
  nor_x1_sg U66550 ( .A(n23712), .B(n40015), .X(n23707) );
  nor_x1_sg U66551 ( .A(n40045), .B(n23711), .X(n23710) );
  nor_x1_sg U66552 ( .A(n23973), .B(n23974), .X(n23972) );
  nor_x1_sg U66553 ( .A(n23977), .B(n40455), .X(n23971) );
  nor_x1_sg U66554 ( .A(n40492), .B(n23976), .X(n23974) );
  nor_x1_sg U66555 ( .A(n24546), .B(n24547), .X(n24545) );
  nor_x1_sg U66556 ( .A(n24549), .B(n39151), .X(n24544) );
  nor_x1_sg U66557 ( .A(n40051), .B(n24548), .X(n24547) );
  nor_x1_sg U66558 ( .A(n24809), .B(n24810), .X(n24808) );
  nor_x1_sg U66559 ( .A(n24813), .B(n40014), .X(n24807) );
  nor_x1_sg U66560 ( .A(n24811), .B(n24812), .X(n24810) );
  nor_x1_sg U66561 ( .A(n25382), .B(n25383), .X(n25381) );
  nor_x1_sg U66562 ( .A(n25385), .B(n41467), .X(n25380) );
  nor_x1_sg U66563 ( .A(n42122), .B(n25384), .X(n25383) );
  nor_x1_sg U66564 ( .A(n25646), .B(n25647), .X(n25645) );
  nor_x1_sg U66565 ( .A(n25650), .B(n40012), .X(n25644) );
  nor_x1_sg U66566 ( .A(n40467), .B(n25649), .X(n25647) );
  nor_x1_sg U66567 ( .A(n26483), .B(n26484), .X(n26482) );
  nor_x1_sg U66568 ( .A(n26487), .B(n41467), .X(n26481) );
  nor_x1_sg U66569 ( .A(n40461), .B(n26486), .X(n26484) );
  nor_x1_sg U66570 ( .A(n22858), .B(n22859), .X(n22857) );
  nor_x1_sg U66571 ( .A(n22862), .B(n39282), .X(n22856) );
  nor_x1_sg U66572 ( .A(n22860), .B(n22861), .X(n22859) );
  nor_x1_sg U66573 ( .A(n23150), .B(n23151), .X(n23149) );
  nor_x1_sg U66574 ( .A(n23153), .B(n40456), .X(n23148) );
  nor_x1_sg U66575 ( .A(n40041), .B(n23152), .X(n23151) );
  nor_x1_sg U66576 ( .A(n23415), .B(n23416), .X(n23414) );
  nor_x1_sg U66577 ( .A(n23419), .B(n41410), .X(n23413) );
  nor_x1_sg U66578 ( .A(n23417), .B(n23418), .X(n23416) );
  nor_x1_sg U66579 ( .A(n23430), .B(n23431), .X(n23429) );
  nor_x1_sg U66580 ( .A(n23433), .B(n40376), .X(n23428) );
  nor_x1_sg U66581 ( .A(n40043), .B(n23432), .X(n23431) );
  nor_x1_sg U66582 ( .A(n23694), .B(n23695), .X(n23693) );
  nor_x1_sg U66583 ( .A(n23698), .B(n41409), .X(n23692) );
  nor_x1_sg U66584 ( .A(n40496), .B(n23697), .X(n23695) );
  nor_x1_sg U66585 ( .A(n23988), .B(n23989), .X(n23987) );
  nor_x1_sg U66586 ( .A(n23991), .B(n41469), .X(n23986) );
  nor_x1_sg U66587 ( .A(n40047), .B(n23990), .X(n23989) );
  nor_x1_sg U66588 ( .A(n24252), .B(n24253), .X(n24251) );
  nor_x1_sg U66589 ( .A(n24256), .B(n41400), .X(n24250) );
  nor_x1_sg U66590 ( .A(n40489), .B(n24255), .X(n24253) );
  nor_x1_sg U66591 ( .A(n24267), .B(n24268), .X(n24266) );
  nor_x1_sg U66592 ( .A(n24270), .B(n41468), .X(n24265) );
  nor_x1_sg U66593 ( .A(n40049), .B(n24269), .X(n24268) );
  nor_x1_sg U66594 ( .A(n24531), .B(n24532), .X(n24530) );
  nor_x1_sg U66595 ( .A(n24535), .B(n39151), .X(n24529) );
  nor_x1_sg U66596 ( .A(n40484), .B(n24534), .X(n24532) );
  nor_x1_sg U66597 ( .A(n24824), .B(n24825), .X(n24823) );
  nor_x1_sg U66598 ( .A(n24827), .B(n40455), .X(n24822) );
  nor_x1_sg U66599 ( .A(n40065), .B(n24826), .X(n24825) );
  nor_x1_sg U66600 ( .A(n25088), .B(n25089), .X(n25087) );
  nor_x1_sg U66601 ( .A(n25092), .B(n39653), .X(n25086) );
  nor_x1_sg U66602 ( .A(n40476), .B(n25091), .X(n25089) );
  nor_x1_sg U66603 ( .A(n25103), .B(n25104), .X(n25102) );
  nor_x1_sg U66604 ( .A(n25106), .B(n39154), .X(n25101) );
  nor_x1_sg U66605 ( .A(n40054), .B(n25105), .X(n25104) );
  nor_x1_sg U66606 ( .A(n25367), .B(n25368), .X(n25366) );
  nor_x1_sg U66607 ( .A(n25371), .B(n41409), .X(n25365) );
  nor_x1_sg U66608 ( .A(n40471), .B(n25370), .X(n25368) );
  nor_x1_sg U66609 ( .A(n25661), .B(n25662), .X(n25660) );
  nor_x1_sg U66610 ( .A(n25664), .B(n41400), .X(n25659) );
  nor_x1_sg U66611 ( .A(n40057), .B(n25663), .X(n25662) );
  nor_x1_sg U66612 ( .A(n26498), .B(n26499), .X(n26497) );
  nor_x1_sg U66613 ( .A(n26501), .B(n40014), .X(n26496) );
  nor_x1_sg U66614 ( .A(n40061), .B(n26500), .X(n26499) );
  nand_x1_sg U66615 ( .A(n39852), .B(n7094), .X(n7432) );
  nand_x1_sg U66616 ( .A(n39499), .B(n40245), .X(n7976) );
  nand_x1_sg U66617 ( .A(n39498), .B(n40250), .X(n8794) );
  nand_x1_sg U66618 ( .A(n39497), .B(n40253), .X(n9614) );
  nand_x1_sg U66619 ( .A(n39496), .B(n40260), .X(n10433) );
  nand_x1_sg U66620 ( .A(n11188), .B(n40263), .X(n11252) );
  nand_x1_sg U66621 ( .A(n12007), .B(n40270), .X(n12071) );
  nand_x1_sg U66622 ( .A(n39493), .B(n40275), .X(n12890) );
  nand_x1_sg U66623 ( .A(n39492), .B(n40279), .X(n13709) );
  nand_x1_sg U66624 ( .A(n39491), .B(n40285), .X(n14528) );
  nand_x1_sg U66625 ( .A(n39215), .B(n40290), .X(n15347) );
  nand_x1_sg U66626 ( .A(n39489), .B(n40293), .X(n16166) );
  nand_x1_sg U66627 ( .A(n39488), .B(n40239), .X(n17804) );
  nand_x1_sg U66628 ( .A(n39487), .B(n40300), .X(n18625) );
  nand_x1_sg U66629 ( .A(n39938), .B(n40134), .X(n8430) );
  nand_x1_sg U66630 ( .A(n39940), .B(n40136), .X(n9248) );
  nand_x1_sg U66631 ( .A(n39942), .B(n40138), .X(n10068) );
  nand_x1_sg U66632 ( .A(n39958), .B(n40140), .X(n10887) );
  nand_x1_sg U66633 ( .A(n39960), .B(n40142), .X(n11706) );
  nand_x1_sg U66634 ( .A(n39950), .B(n40144), .X(n12525) );
  nand_x1_sg U66635 ( .A(n39952), .B(n40146), .X(n13344) );
  nand_x1_sg U66636 ( .A(n39954), .B(n40148), .X(n14163) );
  nand_x1_sg U66637 ( .A(n39948), .B(n40150), .X(n14982) );
  nand_x1_sg U66638 ( .A(n39944), .B(n40152), .X(n15801) );
  nand_x1_sg U66639 ( .A(n39946), .B(n40154), .X(n16620) );
  nand_x1_sg U66640 ( .A(n39934), .B(n40160), .X(n18258) );
  nand_x1_sg U66641 ( .A(n39936), .B(n40155), .X(n19079) );
  nor_x1_sg U66642 ( .A(n5933), .B(n5934), .X(n5932) );
  nand_x1_sg U66643 ( .A(n5964), .B(n19557), .X(n19556) );
  nand_x1_sg U66644 ( .A(n5968), .B(n19543), .X(n19542) );
  nand_x1_sg U66645 ( .A(n7094), .B(n40164), .X(n7157) );
  nand_x1_sg U66646 ( .A(n39809), .B(n39500), .X(n7189) );
  nand_x1_sg U66647 ( .A(n38703), .B(n46578), .X(n20587) );
  inv_x1_sg U66648 ( .A(n22535), .X(n44996) );
  inv_x1_sg U66649 ( .A(n6772), .X(n45821) );
  inv_x1_sg U66650 ( .A(n6781), .X(n45825) );
  inv_x1_sg U66651 ( .A(n6782), .X(n45829) );
  inv_x1_sg U66652 ( .A(n6777), .X(n45833) );
  inv_x1_sg U66653 ( .A(n6778), .X(n45837) );
  inv_x1_sg U66654 ( .A(n6747), .X(n45841) );
  inv_x1_sg U66655 ( .A(n6748), .X(n45845) );
  inv_x1_sg U66656 ( .A(n6743), .X(n45849) );
  inv_x1_sg U66657 ( .A(n6744), .X(n45853) );
  inv_x1_sg U66658 ( .A(n6763), .X(n45857) );
  inv_x1_sg U66659 ( .A(n6771), .X(n45817) );
  inv_x1_sg U66660 ( .A(n6764), .X(n45861) );
  inv_x1_sg U66661 ( .A(n6753), .X(n45865) );
  nand_x1_sg U66662 ( .A(n40133), .B(n8142), .X(n8135) );
  nand_x1_sg U66663 ( .A(n40135), .B(n8960), .X(n8953) );
  nand_x1_sg U66664 ( .A(n40137), .B(n9780), .X(n9773) );
  nand_x1_sg U66665 ( .A(n40139), .B(n10599), .X(n10592) );
  nand_x1_sg U66666 ( .A(n40141), .B(n11418), .X(n11411) );
  nand_x1_sg U66667 ( .A(n40143), .B(n12237), .X(n12230) );
  nand_x1_sg U66668 ( .A(n40145), .B(n13056), .X(n13049) );
  nand_x1_sg U66669 ( .A(n40147), .B(n13875), .X(n13868) );
  nand_x1_sg U66670 ( .A(n40149), .B(n14694), .X(n14687) );
  nand_x1_sg U66671 ( .A(n40151), .B(n15513), .X(n15506) );
  nand_x1_sg U66672 ( .A(n40153), .B(n16332), .X(n16325) );
  nand_x1_sg U66673 ( .A(n17800), .B(n17970), .X(n17963) );
  nand_x1_sg U66674 ( .A(n40155), .B(n18791), .X(n18784) );
  nand_x1_sg U66675 ( .A(n39256), .B(n21767), .X(n21764) );
  nand_x1_sg U66676 ( .A(n41094), .B(n21766), .X(n21765) );
  nand_x1_sg U66677 ( .A(n38936), .B(n21814), .X(n21811) );
  nand_x1_sg U66678 ( .A(n41094), .B(n21813), .X(n21812) );
  nand_x1_sg U66679 ( .A(n38936), .B(n21861), .X(n21858) );
  nand_x1_sg U66680 ( .A(n41095), .B(n21860), .X(n21859) );
  nand_x1_sg U66681 ( .A(n41105), .B(n21907), .X(n21904) );
  nand_x1_sg U66682 ( .A(n39259), .B(n21906), .X(n21905) );
  nand_x1_sg U66683 ( .A(n38936), .B(n21954), .X(n21951) );
  nand_x1_sg U66684 ( .A(n41095), .B(n21953), .X(n21952) );
  nand_x1_sg U66685 ( .A(n39256), .B(n22000), .X(n21997) );
  nand_x1_sg U66686 ( .A(n41106), .B(n22047), .X(n22044) );
  nand_x1_sg U66687 ( .A(n41107), .B(n22093), .X(n22090) );
  nand_x1_sg U66688 ( .A(n41107), .B(n22141), .X(n22138) );
  nand_x1_sg U66689 ( .A(n41106), .B(n22188), .X(n22185) );
  nand_x1_sg U66690 ( .A(n41105), .B(n22236), .X(n22233) );
  nand_x1_sg U66691 ( .A(n39256), .B(n22283), .X(n22280) );
  nand_x1_sg U66692 ( .A(n41106), .B(n22331), .X(n22328) );
  nand_x1_sg U66693 ( .A(n20567), .B(n22378), .X(n22375) );
  nand_x1_sg U66694 ( .A(n41107), .B(n22426), .X(n22423) );
  nand_x1_sg U66695 ( .A(n41107), .B(n22472), .X(n22469) );
  nand_x1_sg U66696 ( .A(n38936), .B(n22518), .X(n22515) );
  nand_x1_sg U66697 ( .A(n22563), .B(n22564), .X(n22562) );
  inv_x1_sg U66698 ( .A(n21445), .X(n45919) );
  inv_x1_sg U66699 ( .A(n28997), .X(n45068) );
  inv_x1_sg U66700 ( .A(n21458), .X(n46010) );
  inv_x1_sg U66701 ( .A(n29010), .X(n45160) );
  inv_x1_sg U66702 ( .A(n21471), .X(n46101) );
  inv_x1_sg U66703 ( .A(n29023), .X(n45251) );
  inv_x1_sg U66704 ( .A(n21484), .X(n46192) );
  inv_x1_sg U66705 ( .A(n29036), .X(n45341) );
  inv_x1_sg U66706 ( .A(n21497), .X(n46283) );
  inv_x1_sg U66707 ( .A(n29049), .X(n45432) );
  inv_x1_sg U66708 ( .A(n21510), .X(n46370) );
  inv_x1_sg U66709 ( .A(n29062), .X(n45521) );
  inv_x1_sg U66710 ( .A(n21523), .X(n46465) );
  inv_x1_sg U66711 ( .A(n29075), .X(n45610) );
  inv_x1_sg U66712 ( .A(n27980), .X(n45037) );
  nand_x1_sg U66713 ( .A(n41781), .B(n39804), .X(n7491) );
  nand_x1_sg U66714 ( .A(n41783), .B(n39938), .X(n8309) );
  nand_x1_sg U66715 ( .A(n41785), .B(n39940), .X(n9127) );
  nand_x1_sg U66716 ( .A(n41787), .B(n39942), .X(n9947) );
  nand_x1_sg U66717 ( .A(n41789), .B(n39958), .X(n10766) );
  nand_x1_sg U66718 ( .A(n41791), .B(n39961), .X(n11585) );
  nand_x1_sg U66719 ( .A(n41793), .B(n39950), .X(n12404) );
  nand_x1_sg U66720 ( .A(n41795), .B(n39952), .X(n13223) );
  nand_x1_sg U66721 ( .A(n41797), .B(n39954), .X(n14042) );
  nand_x1_sg U66722 ( .A(n41799), .B(n39949), .X(n14861) );
  nand_x1_sg U66723 ( .A(n41801), .B(n39944), .X(n15680) );
  nand_x1_sg U66724 ( .A(n41803), .B(n39946), .X(n16499) );
  nand_x1_sg U66725 ( .A(n41805), .B(n39934), .X(n18137) );
  nand_x1_sg U66726 ( .A(n41807), .B(n39936), .X(n18958) );
  inv_x1_sg U66727 ( .A(n26096), .X(n50311) );
  nor_x1_sg U66728 ( .A(n8060), .B(n40632), .X(n8059) );
  nor_x1_sg U66729 ( .A(n8878), .B(n40629), .X(n8877) );
  nor_x1_sg U66730 ( .A(n9698), .B(n40668), .X(n9697) );
  nor_x1_sg U66731 ( .A(n10517), .B(n40659), .X(n10516) );
  nor_x1_sg U66732 ( .A(n11336), .B(n40642), .X(n11335) );
  nor_x1_sg U66733 ( .A(n12155), .B(n40638), .X(n12154) );
  nor_x1_sg U66734 ( .A(n12974), .B(n40664), .X(n12973) );
  nor_x1_sg U66735 ( .A(n13793), .B(n40654), .X(n13792) );
  nor_x1_sg U66736 ( .A(n14612), .B(n40624), .X(n14611) );
  nor_x1_sg U66737 ( .A(n15431), .B(n40682), .X(n15430) );
  nor_x1_sg U66738 ( .A(n16250), .B(n40677), .X(n16249) );
  nor_x1_sg U66739 ( .A(n17888), .B(n40647), .X(n17887) );
  nor_x1_sg U66740 ( .A(n18709), .B(n40672), .X(n18708) );
  nor_x1_sg U66741 ( .A(n7241), .B(n40575), .X(n7240) );
  nor_x1_sg U66742 ( .A(n17066), .B(n40578), .X(n17065) );
  nand_x1_sg U66743 ( .A(n39500), .B(n39773), .X(n7561) );
  nand_x1_sg U66744 ( .A(n7912), .B(n39813), .X(n8008) );
  nand_x1_sg U66745 ( .A(n41785), .B(n39830), .X(n8826) );
  nand_x1_sg U66746 ( .A(n39208), .B(n39846), .X(n9646) );
  nand_x1_sg U66747 ( .A(n39209), .B(n41897), .X(n10465) );
  nand_x1_sg U66748 ( .A(n41791), .B(n41886), .X(n11284) );
  nand_x1_sg U66749 ( .A(n39211), .B(n39836), .X(n12103) );
  nand_x1_sg U66750 ( .A(n41795), .B(n39818), .X(n12922) );
  nand_x1_sg U66751 ( .A(n41797), .B(n39840), .X(n13741) );
  nand_x1_sg U66752 ( .A(n41799), .B(n39842), .X(n14560) );
  nand_x1_sg U66753 ( .A(n15283), .B(n41876), .X(n15379) );
  nand_x1_sg U66754 ( .A(n41803), .B(n41893), .X(n16198) );
  nand_x1_sg U66755 ( .A(n17740), .B(n39828), .X(n17836) );
  nand_x1_sg U66756 ( .A(n41807), .B(n39824), .X(n18657) );
  nand_x1_sg U66757 ( .A(n41064), .B(n26784), .X(n26783) );
  nand_x1_sg U66758 ( .A(n40098), .B(n26785), .X(n26782) );
  nand_x1_sg U66759 ( .A(n41064), .B(n21839), .X(n21838) );
  nand_x1_sg U66760 ( .A(n40095), .B(n21840), .X(n21837) );
  nand_x1_sg U66761 ( .A(n38915), .B(n21886), .X(n21885) );
  nand_x1_sg U66762 ( .A(n40099), .B(n45610), .X(n21884) );
  nand_x1_sg U66763 ( .A(n41063), .B(n21932), .X(n21931) );
  nand_x1_sg U66764 ( .A(n40096), .B(n21933), .X(n21930) );
  nand_x1_sg U66765 ( .A(n41063), .B(n21979), .X(n21978) );
  nand_x1_sg U66766 ( .A(n41397), .B(n45521), .X(n21977) );
  nand_x1_sg U66767 ( .A(n20961), .B(n22025), .X(n22024) );
  nand_x1_sg U66768 ( .A(n41395), .B(n22026), .X(n22023) );
  nand_x1_sg U66769 ( .A(n41063), .B(n22072), .X(n22071) );
  nand_x1_sg U66770 ( .A(n41398), .B(n45432), .X(n22070) );
  nand_x1_sg U66771 ( .A(n41062), .B(n22119), .X(n22118) );
  nand_x1_sg U66772 ( .A(n41397), .B(n22120), .X(n22117) );
  nand_x1_sg U66773 ( .A(n38915), .B(n22167), .X(n22166) );
  nand_x1_sg U66774 ( .A(n40098), .B(n45341), .X(n22165) );
  nand_x1_sg U66775 ( .A(n39266), .B(n22214), .X(n22213) );
  nand_x1_sg U66776 ( .A(n41397), .B(n22215), .X(n22212) );
  nand_x1_sg U66777 ( .A(n41063), .B(n22262), .X(n22261) );
  nand_x1_sg U66778 ( .A(n39148), .B(n45251), .X(n22260) );
  nand_x1_sg U66779 ( .A(n20961), .B(n22309), .X(n22308) );
  nand_x1_sg U66780 ( .A(n41396), .B(n22310), .X(n22307) );
  nand_x1_sg U66781 ( .A(n38915), .B(n22357), .X(n22356) );
  nand_x1_sg U66782 ( .A(n39149), .B(n45160), .X(n22355) );
  nand_x1_sg U66783 ( .A(n41062), .B(n22404), .X(n22403) );
  nand_x1_sg U66784 ( .A(n40100), .B(n22405), .X(n22402) );
  nand_x1_sg U66785 ( .A(n38915), .B(n22451), .X(n22450) );
  nand_x1_sg U66786 ( .A(n40099), .B(n45068), .X(n22449) );
  nand_x1_sg U66787 ( .A(n41064), .B(n22496), .X(n22495) );
  nand_x1_sg U66788 ( .A(n40098), .B(n22497), .X(n22494) );
  nand_x1_sg U66789 ( .A(n39266), .B(n44987), .X(n22537) );
  nand_x1_sg U66790 ( .A(n40096), .B(n44978), .X(n22536) );
  nor_x1_sg U66791 ( .A(n25927), .B(n25928), .X(n25926) );
  nor_x1_sg U66792 ( .A(n25930), .B(n40454), .X(n25925) );
  nor_x1_sg U66793 ( .A(n40037), .B(n25929), .X(n25928) );
  nor_x1_sg U66794 ( .A(n25945), .B(n25946), .X(n25944) );
  nor_x1_sg U66795 ( .A(n25948), .B(n40457), .X(n25943) );
  nor_x1_sg U66796 ( .A(n40071), .B(n25947), .X(n25946) );
  nor_x1_sg U66797 ( .A(n26204), .B(n26205), .X(n26203) );
  nor_x1_sg U66798 ( .A(n26207), .B(n40012), .X(n26202) );
  nor_x1_sg U66799 ( .A(n40059), .B(n26206), .X(n26205) );
  nor_x1_sg U66800 ( .A(n22598), .B(n22599), .X(n22597) );
  nor_x1_sg U66801 ( .A(n22601), .B(n40017), .X(n22596) );
  nor_x1_sg U66802 ( .A(n40369), .B(n22600), .X(n22599) );
  nor_x1_sg U66803 ( .A(n22610), .B(n22611), .X(n22609) );
  nor_x1_sg U66804 ( .A(n22613), .B(n41409), .X(n22608) );
  nor_x1_sg U66805 ( .A(n42325), .B(n22612), .X(n22611) );
  nor_x1_sg U66806 ( .A(n5861), .B(n22701), .X(n22700) );
  nor_x1_sg U66807 ( .A(n22704), .B(n40012), .X(n22699) );
  nor_x1_sg U66808 ( .A(n22702), .B(n22703), .X(n22701) );
  nor_x1_sg U66809 ( .A(n25920), .B(n25921), .X(n25919) );
  nor_x1_sg U66810 ( .A(n25924), .B(n41466), .X(n25918) );
  nor_x1_sg U66811 ( .A(n42370), .B(n25923), .X(n25921) );
  nor_x1_sg U66812 ( .A(n26187), .B(n26188), .X(n26186) );
  nor_x1_sg U66813 ( .A(n26191), .B(n40019), .X(n26185) );
  nor_x1_sg U66814 ( .A(n40463), .B(n26190), .X(n26188) );
  nand_x1_sg U66815 ( .A(n39266), .B(n21745), .X(n21744) );
  nand_x1_sg U66816 ( .A(n41396), .B(n21746), .X(n21743) );
  nand_x1_sg U66817 ( .A(n41064), .B(n21792), .X(n21791) );
  nand_x1_sg U66818 ( .A(n40096), .B(n21793), .X(n21790) );
  nand_x1_sg U66819 ( .A(n46351), .B(n38632), .X(n20319) );
  nand_x1_sg U66820 ( .A(n46535), .B(n38693), .X(n21016) );
  nand_x1_sg U66821 ( .A(n46347), .B(n38638), .X(n19793) );
  nand_x1_sg U66822 ( .A(n46343), .B(n38604), .X(n19355) );
  inv_x1_sg U66823 ( .A(n25920), .X(n50277) );
  inv_x1_sg U66824 ( .A(n22598), .X(n46845) );
  nor_x1_sg U66825 ( .A(n26019), .B(n26020), .X(n26018) );
  nor_x1_sg U66826 ( .A(n41297), .B(n17458), .X(n26020) );
  nor_x1_sg U66827 ( .A(n26021), .B(n39134), .X(n26019) );
  nand_x1_sg U66828 ( .A(n40565), .B(n50277), .X(n25929) );
  nand_x1_sg U66829 ( .A(n46973), .B(n7601), .X(n7598) );
  nand_x1_sg U66830 ( .A(n7600), .B(n47078), .X(n7599) );
  nand_x1_sg U66831 ( .A(n47263), .B(n8419), .X(n8416) );
  nand_x1_sg U66832 ( .A(n8418), .B(n47364), .X(n8417) );
  nand_x1_sg U66833 ( .A(n47548), .B(n9237), .X(n9234) );
  nand_x1_sg U66834 ( .A(n9236), .B(n47649), .X(n9235) );
  nand_x1_sg U66835 ( .A(n47833), .B(n10057), .X(n10054) );
  nand_x1_sg U66836 ( .A(n10056), .B(n47934), .X(n10055) );
  nand_x1_sg U66837 ( .A(n48118), .B(n10876), .X(n10873) );
  nand_x1_sg U66838 ( .A(n10875), .B(n48219), .X(n10874) );
  nand_x1_sg U66839 ( .A(n48403), .B(n11695), .X(n11692) );
  nand_x1_sg U66840 ( .A(n11694), .B(n48504), .X(n11693) );
  nand_x1_sg U66841 ( .A(n48688), .B(n12514), .X(n12511) );
  nand_x1_sg U66842 ( .A(n12513), .B(n48789), .X(n12512) );
  nand_x1_sg U66843 ( .A(n48974), .B(n13333), .X(n13330) );
  nand_x1_sg U66844 ( .A(n13332), .B(n49076), .X(n13331) );
  nand_x1_sg U66845 ( .A(n49261), .B(n14152), .X(n14149) );
  nand_x1_sg U66846 ( .A(n14151), .B(n49362), .X(n14150) );
  nand_x1_sg U66847 ( .A(n49547), .B(n14971), .X(n14968) );
  nand_x1_sg U66848 ( .A(n14970), .B(n49648), .X(n14969) );
  nand_x1_sg U66849 ( .A(n49833), .B(n15790), .X(n15787) );
  nand_x1_sg U66850 ( .A(n15789), .B(n49934), .X(n15788) );
  nand_x1_sg U66851 ( .A(n50119), .B(n16609), .X(n16606) );
  nand_x1_sg U66852 ( .A(n16608), .B(n50220), .X(n16607) );
  nand_x1_sg U66853 ( .A(n50693), .B(n18247), .X(n18244) );
  nand_x1_sg U66854 ( .A(n18246), .B(n50794), .X(n18245) );
  nand_x1_sg U66855 ( .A(n50980), .B(n19068), .X(n19065) );
  nand_x1_sg U66856 ( .A(n19067), .B(n51081), .X(n19066) );
  inv_x1_sg U66857 ( .A(n22858), .X(n47136) );
  inv_x1_sg U66858 ( .A(n23135), .X(n47421) );
  inv_x1_sg U66859 ( .A(n23415), .X(n47706) );
  inv_x1_sg U66860 ( .A(n23694), .X(n47991) );
  inv_x1_sg U66861 ( .A(n23973), .X(n48276) );
  inv_x1_sg U66862 ( .A(n24252), .X(n48561) );
  inv_x1_sg U66863 ( .A(n24531), .X(n48846) );
  inv_x1_sg U66864 ( .A(n24809), .X(n49133) );
  inv_x1_sg U66865 ( .A(n25088), .X(n49419) );
  inv_x1_sg U66866 ( .A(n25367), .X(n49705) );
  inv_x1_sg U66867 ( .A(n25646), .X(n49991) );
  inv_x1_sg U66868 ( .A(n26483), .X(n50852) );
  nand_x1_sg U66869 ( .A(n50404), .B(n17426), .X(n17423) );
  nand_x1_sg U66870 ( .A(n17425), .B(n50505), .X(n17424) );
  inv_x1_sg U66871 ( .A(n26187), .X(n50566) );
  nand_x1_sg U66872 ( .A(n21116), .B(n38650), .X(n21233) );
  nand_x1_sg U66873 ( .A(n21110), .B(n38648), .X(n21236) );
  nand_x1_sg U66874 ( .A(n21104), .B(n38646), .X(n21239) );
  nand_x1_sg U66875 ( .A(n21098), .B(n38644), .X(n21242) );
  nand_x1_sg U66876 ( .A(n21122), .B(n38652), .X(n21230) );
  nand_x1_sg U66877 ( .A(n21128), .B(n38654), .X(n21227) );
  nand_x1_sg U66878 ( .A(n21134), .B(n38656), .X(n21224) );
  nand_x1_sg U66879 ( .A(n21140), .B(n38658), .X(n21221) );
  nand_x1_sg U66880 ( .A(n20431), .B(n38709), .X(n20452) );
  nand_x1_sg U66881 ( .A(n20425), .B(n38724), .X(n20456) );
  nand_x1_sg U66882 ( .A(n20419), .B(n38610), .X(n20459) );
  nand_x1_sg U66883 ( .A(n20413), .B(n38707), .X(n20462) );
  nand_x1_sg U66884 ( .A(n20407), .B(n38612), .X(n20465) );
  nand_x1_sg U66885 ( .A(n20401), .B(n38616), .X(n20468) );
  nand_x1_sg U66886 ( .A(n20395), .B(n38705), .X(n20471) );
  nand_x1_sg U66887 ( .A(n20389), .B(n38614), .X(n20474) );
  nand_x1_sg U66888 ( .A(n21146), .B(n38660), .X(n21218) );
  nand_x1_sg U66889 ( .A(n21152), .B(n38662), .X(n21215) );
  nand_x1_sg U66890 ( .A(n21158), .B(n38664), .X(n21212) );
  nand_x1_sg U66891 ( .A(n21164), .B(n38666), .X(n21209) );
  nand_x1_sg U66892 ( .A(n19698), .B(n38697), .X(n19795) );
  nand_x1_sg U66893 ( .A(n19692), .B(n38691), .X(n19799) );
  nand_x1_sg U66894 ( .A(n19686), .B(n38687), .X(n19802) );
  nand_x1_sg U66895 ( .A(n19680), .B(n38685), .X(n19805) );
  nand_x1_sg U66896 ( .A(n19674), .B(n38683), .X(n19808) );
  nand_x1_sg U66897 ( .A(n19668), .B(n38681), .X(n19811) );
  nand_x1_sg U66898 ( .A(n19662), .B(n38679), .X(n19814) );
  nand_x1_sg U66899 ( .A(n19656), .B(n38677), .X(n19817) );
  nand_x1_sg U66900 ( .A(n41834), .B(n47146), .X(n22882) );
  nand_x1_sg U66901 ( .A(n41832), .B(n47431), .X(n23159) );
  nand_x1_sg U66902 ( .A(n41830), .B(n47716), .X(n23439) );
  nand_x1_sg U66903 ( .A(n41828), .B(n48001), .X(n23718) );
  nand_x1_sg U66904 ( .A(n41826), .B(n48286), .X(n23997) );
  nand_x1_sg U66905 ( .A(n41824), .B(n48571), .X(n24276) );
  nand_x1_sg U66906 ( .A(n41822), .B(n48857), .X(n24555) );
  nand_x1_sg U66907 ( .A(n41820), .B(n49144), .X(n24833) );
  nand_x1_sg U66908 ( .A(n41818), .B(n49430), .X(n25112) );
  nand_x1_sg U66909 ( .A(n41816), .B(n49715), .X(n25391) );
  nand_x1_sg U66910 ( .A(n41814), .B(n50002), .X(n25670) );
  nand_x1_sg U66911 ( .A(n41810), .B(n50576), .X(n26214) );
  nand_x1_sg U66912 ( .A(n41812), .B(n50863), .X(n26507) );
  inv_x1_sg U66913 ( .A(n19557), .X(n46565) );
  inv_x1_sg U66914 ( .A(n19543), .X(n46560) );
  nand_x1_sg U66915 ( .A(n7153), .B(n40080), .X(n7152) );
  nand_x1_sg U66916 ( .A(n38729), .B(n7154), .X(n7151) );
  nor_x1_sg U66917 ( .A(n41058), .B(n7104), .X(n7153) );
  nand_x1_sg U66918 ( .A(n7971), .B(n40133), .X(n7970) );
  nand_x1_sg U66919 ( .A(n38731), .B(n7973), .X(n7969) );
  nor_x1_sg U66920 ( .A(n41937), .B(n7922), .X(n7971) );
  nand_x1_sg U66921 ( .A(n8789), .B(n40135), .X(n8788) );
  nand_x1_sg U66922 ( .A(n38733), .B(n8791), .X(n8787) );
  nor_x1_sg U66923 ( .A(n39967), .B(n8740), .X(n8789) );
  nand_x1_sg U66924 ( .A(n9609), .B(n40137), .X(n9608) );
  nand_x1_sg U66925 ( .A(n38735), .B(n9611), .X(n9607) );
  nor_x1_sg U66926 ( .A(n39971), .B(n9560), .X(n9609) );
  nand_x1_sg U66927 ( .A(n10428), .B(n40139), .X(n10427) );
  nand_x1_sg U66928 ( .A(n38737), .B(n10430), .X(n10426) );
  nor_x1_sg U66929 ( .A(n39976), .B(n10379), .X(n10428) );
  nand_x1_sg U66930 ( .A(n11247), .B(n40141), .X(n11246) );
  nand_x1_sg U66931 ( .A(n38739), .B(n11249), .X(n11245) );
  nor_x1_sg U66932 ( .A(n41939), .B(n11198), .X(n11247) );
  nand_x1_sg U66933 ( .A(n12066), .B(n40143), .X(n12065) );
  nand_x1_sg U66934 ( .A(n38741), .B(n12068), .X(n12064) );
  nor_x1_sg U66935 ( .A(n39984), .B(n12017), .X(n12066) );
  nand_x1_sg U66936 ( .A(n12885), .B(n40145), .X(n12884) );
  nand_x1_sg U66937 ( .A(n38743), .B(n12887), .X(n12883) );
  nor_x1_sg U66938 ( .A(n39988), .B(n12836), .X(n12885) );
  nand_x1_sg U66939 ( .A(n13704), .B(n40147), .X(n13703) );
  nand_x1_sg U66940 ( .A(n38745), .B(n13706), .X(n13702) );
  nor_x1_sg U66941 ( .A(n39993), .B(n13655), .X(n13704) );
  nand_x1_sg U66942 ( .A(n14523), .B(n40149), .X(n14522) );
  nand_x1_sg U66943 ( .A(n38747), .B(n14525), .X(n14521) );
  nor_x1_sg U66944 ( .A(n41932), .B(n14474), .X(n14523) );
  nand_x1_sg U66945 ( .A(n15342), .B(n42168), .X(n15341) );
  nand_x1_sg U66946 ( .A(n38749), .B(n15344), .X(n15340) );
  nor_x1_sg U66947 ( .A(n39999), .B(n15293), .X(n15342) );
  nand_x1_sg U66948 ( .A(n16161), .B(n40153), .X(n16160) );
  nand_x1_sg U66949 ( .A(n38751), .B(n16163), .X(n16159) );
  nor_x1_sg U66950 ( .A(n41942), .B(n16112), .X(n16161) );
  nand_x1_sg U66951 ( .A(n17799), .B(n40159), .X(n17798) );
  nand_x1_sg U66952 ( .A(n38753), .B(n17801), .X(n17797) );
  nor_x1_sg U66953 ( .A(n41001), .B(n17750), .X(n17799) );
  nand_x1_sg U66954 ( .A(n18620), .B(n40155), .X(n18619) );
  nand_x1_sg U66955 ( .A(n38755), .B(n18622), .X(n18618) );
  nor_x1_sg U66956 ( .A(n41910), .B(n18571), .X(n18620) );
  nand_x1_sg U66957 ( .A(n16978), .B(n40078), .X(n16977) );
  nand_x1_sg U66958 ( .A(n38727), .B(n16979), .X(n16976) );
  nor_x1_sg U66959 ( .A(n40996), .B(n16929), .X(n16978) );
  nand_x2_sg U66960 ( .A(n7548), .B(n7529), .X(n7547) );
  nand_x1_sg U66961 ( .A(n7552), .B(n7551), .X(n7546) );
  nor_x1_sg U66962 ( .A(n41059), .B(n41631), .X(n7548) );
  nand_x2_sg U66963 ( .A(n17373), .B(n17354), .X(n17372) );
  nand_x1_sg U66964 ( .A(n17377), .B(n17376), .X(n17371) );
  nor_x1_sg U66965 ( .A(n40994), .B(n41618), .X(n17373) );
  nand_x1_sg U66966 ( .A(n7930), .B(n7929), .X(n7881) );
  nand_x1_sg U66967 ( .A(n8748), .B(n8747), .X(n8699) );
  nand_x1_sg U66968 ( .A(n9568), .B(n9567), .X(n9519) );
  nand_x1_sg U66969 ( .A(n10387), .B(n10386), .X(n10338) );
  nand_x1_sg U66970 ( .A(n11206), .B(n11205), .X(n11157) );
  nand_x1_sg U66971 ( .A(n12025), .B(n12024), .X(n11976) );
  nand_x1_sg U66972 ( .A(n12844), .B(n41822), .X(n12795) );
  nand_x1_sg U66973 ( .A(n13663), .B(n13662), .X(n13614) );
  nand_x1_sg U66974 ( .A(n14482), .B(n41818), .X(n14433) );
  nand_x1_sg U66975 ( .A(n15301), .B(n15300), .X(n15252) );
  nand_x1_sg U66976 ( .A(n16120), .B(n41814), .X(n16071) );
  nand_x1_sg U66977 ( .A(n17758), .B(n41811), .X(n17709) );
  nand_x1_sg U66978 ( .A(n18579), .B(n41812), .X(n18530) );
  nand_x1_sg U66979 ( .A(n7112), .B(n40234), .X(n7063) );
  nand_x1_sg U66980 ( .A(n16937), .B(n40230), .X(n16890) );
  nor_x1_sg U66981 ( .A(n40975), .B(n7646), .X(\L2_0/n3440 ) );
  nand_x1_sg U66982 ( .A(n6958), .B(n7102), .X(n7500) );
  nor_x1_sg U66983 ( .A(n38913), .B(n41666), .X(n7502) );
  nand_x1_sg U66984 ( .A(n7775), .B(n7920), .X(n8318) );
  nor_x1_sg U66985 ( .A(n41937), .B(n38998), .X(n8320) );
  nand_x1_sg U66986 ( .A(n8593), .B(n8738), .X(n9136) );
  nor_x1_sg U66987 ( .A(n39969), .B(n38997), .X(n9138) );
  nand_x1_sg U66988 ( .A(n9413), .B(n9558), .X(n9956) );
  nor_x1_sg U66989 ( .A(n39973), .B(n38996), .X(n9958) );
  nand_x1_sg U66990 ( .A(n10232), .B(n10377), .X(n10775) );
  nor_x1_sg U66991 ( .A(n41926), .B(n38995), .X(n10777) );
  nand_x1_sg U66992 ( .A(n11051), .B(n11196), .X(n11594) );
  nor_x1_sg U66993 ( .A(n39980), .B(n39002), .X(n11596) );
  nand_x1_sg U66994 ( .A(n11870), .B(n12015), .X(n12413) );
  nor_x1_sg U66995 ( .A(n41924), .B(n39001), .X(n12415) );
  nand_x1_sg U66996 ( .A(n12689), .B(n12834), .X(n13232) );
  nor_x1_sg U66997 ( .A(n41923), .B(n39000), .X(n13234) );
  nand_x1_sg U66998 ( .A(n13508), .B(n13653), .X(n14051) );
  nor_x1_sg U66999 ( .A(n39991), .B(n38999), .X(n14053) );
  nand_x1_sg U67000 ( .A(n14327), .B(n14472), .X(n14870) );
  nor_x1_sg U67001 ( .A(n40725), .B(n39006), .X(n14872) );
  nand_x1_sg U67002 ( .A(n15146), .B(n15291), .X(n15689) );
  nor_x1_sg U67003 ( .A(n41920), .B(n39005), .X(n15691) );
  nand_x1_sg U67004 ( .A(n15965), .B(n16110), .X(n16508) );
  nor_x1_sg U67005 ( .A(n40004), .B(n39004), .X(n16510) );
  nand_x1_sg U67006 ( .A(n17603), .B(n17748), .X(n18146) );
  nor_x1_sg U67007 ( .A(n41000), .B(n39007), .X(n18148) );
  nand_x1_sg U67008 ( .A(n18424), .B(n18569), .X(n18967) );
  nor_x1_sg U67009 ( .A(n40007), .B(n39003), .X(n18969) );
  nand_x2_sg U67010 ( .A(n8366), .B(n8347), .X(n8365) );
  nand_x1_sg U67011 ( .A(n8370), .B(n8369), .X(n8364) );
  nor_x1_sg U67012 ( .A(n40685), .B(n41629), .X(n8366) );
  nand_x2_sg U67013 ( .A(n9184), .B(n9165), .X(n9183) );
  nand_x1_sg U67014 ( .A(n9188), .B(n9187), .X(n9182) );
  nor_x1_sg U67015 ( .A(n41928), .B(n41630), .X(n9184) );
  nand_x2_sg U67016 ( .A(n10004), .B(n9985), .X(n10003) );
  nand_x1_sg U67017 ( .A(n10008), .B(n10007), .X(n10002) );
  nor_x1_sg U67018 ( .A(n39971), .B(n41628), .X(n10004) );
  nand_x2_sg U67019 ( .A(n10823), .B(n10804), .X(n10822) );
  nand_x1_sg U67020 ( .A(n10827), .B(n10826), .X(n10821) );
  nor_x1_sg U67021 ( .A(n41926), .B(n41626), .X(n10823) );
  nand_x2_sg U67022 ( .A(n11642), .B(n11623), .X(n11641) );
  nand_x1_sg U67023 ( .A(n11646), .B(n11645), .X(n11640) );
  nor_x1_sg U67024 ( .A(n40705), .B(n41627), .X(n11642) );
  nand_x2_sg U67025 ( .A(n12461), .B(n12442), .X(n12460) );
  nand_x1_sg U67026 ( .A(n12465), .B(n12464), .X(n12459) );
  nor_x1_sg U67027 ( .A(n41924), .B(n41625), .X(n12461) );
  nand_x2_sg U67028 ( .A(n13280), .B(n13261), .X(n13279) );
  nand_x1_sg U67029 ( .A(n13284), .B(n13283), .X(n13278) );
  nor_x1_sg U67030 ( .A(n41923), .B(n39079), .X(n13280) );
  nand_x2_sg U67031 ( .A(n14099), .B(n14080), .X(n14098) );
  nand_x1_sg U67032 ( .A(n14103), .B(n14102), .X(n14097) );
  nor_x1_sg U67033 ( .A(n41938), .B(n41624), .X(n14099) );
  nand_x2_sg U67034 ( .A(n14918), .B(n14899), .X(n14917) );
  nand_x1_sg U67035 ( .A(n14922), .B(n14921), .X(n14916) );
  nor_x1_sg U67036 ( .A(n41932), .B(n41623), .X(n14918) );
  nand_x2_sg U67037 ( .A(n15737), .B(n15718), .X(n15736) );
  nand_x1_sg U67038 ( .A(n15741), .B(n15740), .X(n15735) );
  nor_x1_sg U67039 ( .A(n41920), .B(n41621), .X(n15737) );
  nand_x2_sg U67040 ( .A(n16556), .B(n16537), .X(n16555) );
  nand_x1_sg U67041 ( .A(n16560), .B(n16559), .X(n16554) );
  nor_x1_sg U67042 ( .A(n40735), .B(n41622), .X(n16556) );
  nand_x2_sg U67043 ( .A(n18194), .B(n18175), .X(n18193) );
  nand_x1_sg U67044 ( .A(n18198), .B(n18197), .X(n18192) );
  nor_x1_sg U67045 ( .A(n38910), .B(n39025), .X(n18194) );
  nand_x2_sg U67046 ( .A(n19015), .B(n18996), .X(n19014) );
  nand_x1_sg U67047 ( .A(n19019), .B(n19018), .X(n19013) );
  nor_x1_sg U67048 ( .A(n40008), .B(n41620), .X(n19015) );
  nand_x1_sg U67049 ( .A(n16782), .B(n16927), .X(n17325) );
  nor_x1_sg U67050 ( .A(n40993), .B(n41693), .X(n17327) );
  nand_x1_sg U67051 ( .A(n40633), .B(n47169), .X(n22896) );
  nand_x1_sg U67052 ( .A(n40629), .B(n47454), .X(n23173) );
  nand_x1_sg U67053 ( .A(n40667), .B(n47739), .X(n23453) );
  nand_x1_sg U67054 ( .A(n40659), .B(n48024), .X(n23732) );
  nand_x1_sg U67055 ( .A(n40643), .B(n48309), .X(n24011) );
  nand_x1_sg U67056 ( .A(n40639), .B(n48594), .X(n24290) );
  nand_x1_sg U67057 ( .A(n40664), .B(n48880), .X(n24569) );
  nand_x1_sg U67058 ( .A(n40653), .B(n49167), .X(n24847) );
  nand_x1_sg U67059 ( .A(n40623), .B(n49453), .X(n25126) );
  nand_x1_sg U67060 ( .A(n40682), .B(n49738), .X(n25405) );
  nand_x1_sg U67061 ( .A(n40677), .B(n50025), .X(n25684) );
  nand_x1_sg U67062 ( .A(n40647), .B(n50599), .X(n26230) );
  nand_x1_sg U67063 ( .A(n40674), .B(n50886), .X(n26521) );
  nand_x1_sg U67064 ( .A(n7112), .B(n41779), .X(n7109) );
  nand_x1_sg U67065 ( .A(n40233), .B(n46896), .X(n7110) );
  inv_x1_sg U67066 ( .A(n7112), .X(n46896) );
  nand_x1_sg U67067 ( .A(n16937), .B(n41778), .X(n16934) );
  nand_x1_sg U67068 ( .A(n40229), .B(n50329), .X(n16935) );
  inv_x1_sg U67069 ( .A(n16937), .X(n50329) );
  nand_x1_sg U67070 ( .A(n7930), .B(n40179), .X(n7927) );
  nand_x1_sg U67071 ( .A(n41835), .B(n47191), .X(n7928) );
  inv_x1_sg U67072 ( .A(n7930), .X(n47191) );
  nand_x1_sg U67073 ( .A(n8748), .B(n40211), .X(n8745) );
  nand_x1_sg U67074 ( .A(n41833), .B(n47476), .X(n8746) );
  inv_x1_sg U67075 ( .A(n8748), .X(n47476) );
  nand_x1_sg U67076 ( .A(n9568), .B(n40207), .X(n9565) );
  nand_x1_sg U67077 ( .A(n41830), .B(n47761), .X(n9566) );
  inv_x1_sg U67078 ( .A(n9568), .X(n47761) );
  nand_x1_sg U67079 ( .A(n10387), .B(n40203), .X(n10384) );
  nand_x1_sg U67080 ( .A(n41829), .B(n48046), .X(n10385) );
  inv_x1_sg U67081 ( .A(n10387), .X(n48046) );
  nand_x1_sg U67082 ( .A(n11206), .B(n40199), .X(n11203) );
  nand_x1_sg U67083 ( .A(n41827), .B(n48331), .X(n11204) );
  inv_x1_sg U67084 ( .A(n11206), .X(n48331) );
  nand_x1_sg U67085 ( .A(n12025), .B(n40195), .X(n12022) );
  nand_x1_sg U67086 ( .A(n41825), .B(n48616), .X(n12023) );
  inv_x1_sg U67087 ( .A(n12025), .X(n48616) );
  nand_x1_sg U67088 ( .A(n12844), .B(n40191), .X(n12841) );
  nand_x1_sg U67089 ( .A(n12843), .B(n48902), .X(n12842) );
  inv_x1_sg U67090 ( .A(n12844), .X(n48902) );
  nand_x1_sg U67091 ( .A(n13663), .B(n40175), .X(n13660) );
  nand_x1_sg U67092 ( .A(n41820), .B(n49189), .X(n13661) );
  inv_x1_sg U67093 ( .A(n13663), .X(n49189) );
  nand_x1_sg U67094 ( .A(n14482), .B(n40187), .X(n14479) );
  nand_x1_sg U67095 ( .A(n14481), .B(n49475), .X(n14480) );
  inv_x1_sg U67096 ( .A(n14482), .X(n49475) );
  nand_x1_sg U67097 ( .A(n15301), .B(n40171), .X(n15298) );
  nand_x1_sg U67098 ( .A(n41817), .B(n49761), .X(n15299) );
  inv_x1_sg U67099 ( .A(n15301), .X(n49761) );
  nand_x1_sg U67100 ( .A(n16120), .B(n40167), .X(n16117) );
  nand_x1_sg U67101 ( .A(n16119), .B(n50047), .X(n16118) );
  inv_x1_sg U67102 ( .A(n16120), .X(n50047) );
  nand_x1_sg U67103 ( .A(n17758), .B(n40215), .X(n17755) );
  nand_x1_sg U67104 ( .A(n17757), .B(n50621), .X(n17756) );
  inv_x1_sg U67105 ( .A(n17758), .X(n50621) );
  nand_x1_sg U67106 ( .A(n18579), .B(n40183), .X(n18576) );
  nand_x1_sg U67107 ( .A(n18578), .B(n50908), .X(n18577) );
  inv_x1_sg U67108 ( .A(n18579), .X(n50908) );
  nand_x1_sg U67109 ( .A(n16995), .B(n40074), .X(n16993) );
  nand_x1_sg U67110 ( .A(n39771), .B(n50362), .X(n16994) );
  nand_x1_sg U67111 ( .A(n46863), .B(n7086), .X(n7091) );
  nand_x1_sg U67112 ( .A(n7093), .B(n41781), .X(n7092) );
  nor_x1_sg U67113 ( .A(n41059), .B(n7095), .X(n7093) );
  nand_x1_sg U67114 ( .A(n47156), .B(n7904), .X(n7909) );
  nand_x1_sg U67115 ( .A(n7911), .B(n39206), .X(n7910) );
  nor_x1_sg U67116 ( .A(n39964), .B(n7913), .X(n7911) );
  nand_x1_sg U67117 ( .A(n47441), .B(n8722), .X(n8727) );
  nand_x1_sg U67118 ( .A(n8729), .B(n39207), .X(n8728) );
  nor_x1_sg U67119 ( .A(n39969), .B(n8731), .X(n8729) );
  nand_x1_sg U67120 ( .A(n47726), .B(n9542), .X(n9547) );
  nand_x1_sg U67121 ( .A(n9549), .B(n39497), .X(n9548) );
  nor_x1_sg U67122 ( .A(n41933), .B(n9551), .X(n9549) );
  nand_x1_sg U67123 ( .A(n48011), .B(n10361), .X(n10366) );
  nand_x1_sg U67124 ( .A(n10368), .B(n39496), .X(n10367) );
  nor_x1_sg U67125 ( .A(n39976), .B(n10370), .X(n10368) );
  nand_x1_sg U67126 ( .A(n48296), .B(n11180), .X(n11185) );
  nand_x1_sg U67127 ( .A(n11187), .B(n39210), .X(n11186) );
  nor_x1_sg U67128 ( .A(n39981), .B(n11189), .X(n11187) );
  nand_x1_sg U67129 ( .A(n48581), .B(n11999), .X(n12004) );
  nand_x1_sg U67130 ( .A(n12006), .B(n39494), .X(n12005) );
  nor_x1_sg U67131 ( .A(n41943), .B(n12008), .X(n12006) );
  nand_x1_sg U67132 ( .A(n48867), .B(n12818), .X(n12823) );
  nand_x1_sg U67133 ( .A(n12825), .B(n39212), .X(n12824) );
  nor_x1_sg U67134 ( .A(n39988), .B(n12827), .X(n12825) );
  nand_x1_sg U67135 ( .A(n49154), .B(n13637), .X(n13642) );
  nand_x1_sg U67136 ( .A(n13644), .B(n39213), .X(n13643) );
  nor_x1_sg U67137 ( .A(n39993), .B(n13646), .X(n13644) );
  nand_x1_sg U67138 ( .A(n49440), .B(n14456), .X(n14461) );
  nand_x1_sg U67139 ( .A(n14463), .B(n39214), .X(n14462) );
  nor_x1_sg U67140 ( .A(n39995), .B(n14465), .X(n14463) );
  nand_x1_sg U67141 ( .A(n49725), .B(n15275), .X(n15280) );
  nand_x1_sg U67142 ( .A(n15282), .B(n39490), .X(n15281) );
  nor_x1_sg U67143 ( .A(n40000), .B(n15284), .X(n15282) );
  nand_x1_sg U67144 ( .A(n50012), .B(n16094), .X(n16099) );
  nand_x1_sg U67145 ( .A(n16101), .B(n39216), .X(n16100) );
  nor_x1_sg U67146 ( .A(n40004), .B(n16103), .X(n16101) );
  nand_x1_sg U67147 ( .A(n50296), .B(n16912), .X(n16917) );
  nand_x1_sg U67148 ( .A(n16919), .B(n40073), .X(n16918) );
  nor_x1_sg U67149 ( .A(n40996), .B(n16920), .X(n16919) );
  nand_x1_sg U67150 ( .A(n50586), .B(n17732), .X(n17737) );
  nand_x1_sg U67151 ( .A(n17739), .B(n39488), .X(n17738) );
  nor_x1_sg U67152 ( .A(n40998), .B(n17741), .X(n17739) );
  nand_x1_sg U67153 ( .A(n50873), .B(n18553), .X(n18558) );
  nand_x1_sg U67154 ( .A(n18560), .B(n39218), .X(n18559) );
  nor_x1_sg U67155 ( .A(n41910), .B(n18562), .X(n18560) );
  nand_x1_sg U67156 ( .A(n47010), .B(n7444), .X(n7441) );
  nand_x1_sg U67157 ( .A(n46899), .B(n7443), .X(n7442) );
  nand_x1_sg U67158 ( .A(n50439), .B(n17269), .X(n17266) );
  nand_x1_sg U67159 ( .A(n50332), .B(n17268), .X(n17267) );
  nand_x1_sg U67160 ( .A(n47298), .B(n8262), .X(n8259) );
  nand_x1_sg U67161 ( .A(n47194), .B(n8261), .X(n8260) );
  nand_x1_sg U67162 ( .A(n47583), .B(n9080), .X(n9077) );
  nand_x1_sg U67163 ( .A(n47479), .B(n9079), .X(n9078) );
  nand_x1_sg U67164 ( .A(n47868), .B(n9900), .X(n9897) );
  nand_x1_sg U67165 ( .A(n47764), .B(n9899), .X(n9898) );
  nand_x1_sg U67166 ( .A(n48153), .B(n10719), .X(n10716) );
  nand_x1_sg U67167 ( .A(n48049), .B(n10718), .X(n10717) );
  nand_x1_sg U67168 ( .A(n48438), .B(n11538), .X(n11535) );
  nand_x1_sg U67169 ( .A(n48334), .B(n11537), .X(n11536) );
  nand_x1_sg U67170 ( .A(n48723), .B(n12357), .X(n12354) );
  nand_x1_sg U67171 ( .A(n48619), .B(n12356), .X(n12355) );
  nand_x1_sg U67172 ( .A(n49009), .B(n13176), .X(n13173) );
  nand_x1_sg U67173 ( .A(n48905), .B(n13175), .X(n13174) );
  nand_x1_sg U67174 ( .A(n49296), .B(n13995), .X(n13992) );
  nand_x1_sg U67175 ( .A(n49192), .B(n13994), .X(n13993) );
  nand_x1_sg U67176 ( .A(n49582), .B(n14814), .X(n14811) );
  nand_x1_sg U67177 ( .A(n49478), .B(n14813), .X(n14812) );
  nand_x1_sg U67178 ( .A(n49868), .B(n15633), .X(n15630) );
  nand_x1_sg U67179 ( .A(n49764), .B(n15632), .X(n15631) );
  nand_x1_sg U67180 ( .A(n50154), .B(n16452), .X(n16449) );
  nand_x1_sg U67181 ( .A(n50050), .B(n16451), .X(n16450) );
  nand_x1_sg U67182 ( .A(n50728), .B(n18090), .X(n18087) );
  nand_x1_sg U67183 ( .A(n50624), .B(n18089), .X(n18088) );
  nand_x1_sg U67184 ( .A(n51015), .B(n18911), .X(n18908) );
  nand_x1_sg U67185 ( .A(n50911), .B(n18910), .X(n18909) );
  nand_x1_sg U67186 ( .A(n7529), .B(n7528), .X(n7526) );
  nor_x1_sg U67187 ( .A(n7528), .B(n7529), .X(n7527) );
  nand_x1_sg U67188 ( .A(n8347), .B(n8346), .X(n8344) );
  nor_x1_sg U67189 ( .A(n8346), .B(n8347), .X(n8345) );
  nand_x1_sg U67190 ( .A(n9165), .B(n9164), .X(n9162) );
  nor_x1_sg U67191 ( .A(n9164), .B(n9165), .X(n9163) );
  nand_x1_sg U67192 ( .A(n9985), .B(n9984), .X(n9982) );
  nor_x1_sg U67193 ( .A(n9984), .B(n9985), .X(n9983) );
  nand_x1_sg U67194 ( .A(n10804), .B(n10803), .X(n10801) );
  nor_x1_sg U67195 ( .A(n10803), .B(n10804), .X(n10802) );
  nand_x1_sg U67196 ( .A(n11623), .B(n11622), .X(n11620) );
  nor_x1_sg U67197 ( .A(n11622), .B(n11623), .X(n11621) );
  nand_x1_sg U67198 ( .A(n12442), .B(n12441), .X(n12439) );
  nor_x1_sg U67199 ( .A(n12441), .B(n12442), .X(n12440) );
  nand_x1_sg U67200 ( .A(n13261), .B(n13260), .X(n13258) );
  nor_x1_sg U67201 ( .A(n13260), .B(n13261), .X(n13259) );
  nand_x1_sg U67202 ( .A(n14080), .B(n14079), .X(n14077) );
  nor_x1_sg U67203 ( .A(n14079), .B(n14080), .X(n14078) );
  nand_x1_sg U67204 ( .A(n14899), .B(n14898), .X(n14896) );
  nor_x1_sg U67205 ( .A(n14898), .B(n14899), .X(n14897) );
  nand_x1_sg U67206 ( .A(n15718), .B(n15717), .X(n15715) );
  nor_x1_sg U67207 ( .A(n15717), .B(n15718), .X(n15716) );
  nand_x1_sg U67208 ( .A(n16537), .B(n16536), .X(n16534) );
  nor_x1_sg U67209 ( .A(n16536), .B(n16537), .X(n16535) );
  nand_x1_sg U67210 ( .A(n17354), .B(n17353), .X(n17351) );
  nor_x1_sg U67211 ( .A(n17353), .B(n17354), .X(n17352) );
  nand_x1_sg U67212 ( .A(n18175), .B(n18174), .X(n18172) );
  nor_x1_sg U67213 ( .A(n18174), .B(n18175), .X(n18173) );
  nand_x1_sg U67214 ( .A(n18996), .B(n18995), .X(n18993) );
  nor_x1_sg U67215 ( .A(n18995), .B(n18996), .X(n18994) );
  nand_x1_sg U67216 ( .A(n7170), .B(n39500), .X(n7168) );
  nand_x1_sg U67217 ( .A(n39723), .B(n46929), .X(n7169) );
  nand_x1_sg U67218 ( .A(n7989), .B(n39499), .X(n7987) );
  nand_x1_sg U67219 ( .A(n39720), .B(n47221), .X(n7988) );
  nand_x1_sg U67220 ( .A(n8807), .B(n39498), .X(n8805) );
  nand_x1_sg U67221 ( .A(n39717), .B(n47506), .X(n8806) );
  nand_x1_sg U67222 ( .A(n9627), .B(n39497), .X(n9625) );
  nand_x1_sg U67223 ( .A(n39714), .B(n47791), .X(n9626) );
  nand_x1_sg U67224 ( .A(n10446), .B(n39496), .X(n10444) );
  nand_x1_sg U67225 ( .A(n39711), .B(n48076), .X(n10445) );
  nand_x1_sg U67226 ( .A(n11265), .B(n39495), .X(n11263) );
  nand_x1_sg U67227 ( .A(n39708), .B(n48361), .X(n11264) );
  nand_x1_sg U67228 ( .A(n12084), .B(n39494), .X(n12082) );
  nand_x1_sg U67229 ( .A(n39705), .B(n48646), .X(n12083) );
  nand_x1_sg U67230 ( .A(n12903), .B(n39493), .X(n12901) );
  nand_x1_sg U67231 ( .A(n39702), .B(n48932), .X(n12902) );
  nand_x1_sg U67232 ( .A(n13722), .B(n39492), .X(n13720) );
  nand_x1_sg U67233 ( .A(n39699), .B(n49219), .X(n13721) );
  nand_x1_sg U67234 ( .A(n14541), .B(n39491), .X(n14539) );
  nand_x1_sg U67235 ( .A(n39696), .B(n49505), .X(n14540) );
  nand_x1_sg U67236 ( .A(n15360), .B(n39490), .X(n15358) );
  nand_x1_sg U67237 ( .A(n39693), .B(n49791), .X(n15359) );
  nand_x1_sg U67238 ( .A(n16179), .B(n39489), .X(n16177) );
  nand_x1_sg U67239 ( .A(n39690), .B(n50077), .X(n16178) );
  nand_x1_sg U67240 ( .A(n17817), .B(n39488), .X(n17815) );
  nand_x1_sg U67241 ( .A(n39687), .B(n50651), .X(n17816) );
  nand_x1_sg U67242 ( .A(n18638), .B(n39487), .X(n18636) );
  nand_x1_sg U67243 ( .A(n39684), .B(n50938), .X(n18637) );
  nand_x1_sg U67244 ( .A(n46991), .B(n7583), .X(n7580) );
  nand_x1_sg U67245 ( .A(n6957), .B(n7582), .X(n7581) );
  nand_x1_sg U67246 ( .A(n39802), .B(n40234), .X(n7583) );
  nand_x1_sg U67247 ( .A(n47280), .B(n8401), .X(n8398) );
  nand_x1_sg U67248 ( .A(n7774), .B(n8400), .X(n8399) );
  nand_x1_sg U67249 ( .A(n39799), .B(n41834), .X(n8401) );
  nand_x1_sg U67250 ( .A(n47565), .B(n9219), .X(n9216) );
  nand_x1_sg U67251 ( .A(n8592), .B(n9218), .X(n9217) );
  nand_x1_sg U67252 ( .A(n39800), .B(n41832), .X(n9219) );
  nand_x1_sg U67253 ( .A(n47850), .B(n10039), .X(n10036) );
  nand_x1_sg U67254 ( .A(n9412), .B(n10038), .X(n10037) );
  nand_x1_sg U67255 ( .A(n39795), .B(n41830), .X(n10039) );
  nand_x1_sg U67256 ( .A(n48135), .B(n10858), .X(n10855) );
  nand_x1_sg U67257 ( .A(n10231), .B(n10857), .X(n10856) );
  nand_x1_sg U67258 ( .A(n39796), .B(n41829), .X(n10858) );
  nand_x1_sg U67259 ( .A(n48420), .B(n11677), .X(n11674) );
  nand_x1_sg U67260 ( .A(n11050), .B(n11676), .X(n11675) );
  nand_x1_sg U67261 ( .A(n39791), .B(n41827), .X(n11677) );
  nand_x1_sg U67262 ( .A(n48705), .B(n12496), .X(n12493) );
  nand_x1_sg U67263 ( .A(n11869), .B(n12495), .X(n12494) );
  nand_x1_sg U67264 ( .A(n39792), .B(n41825), .X(n12496) );
  nand_x1_sg U67265 ( .A(n48991), .B(n13315), .X(n13312) );
  nand_x1_sg U67266 ( .A(n12688), .B(n13314), .X(n13313) );
  nand_x1_sg U67267 ( .A(n39787), .B(n12843), .X(n13315) );
  nand_x1_sg U67268 ( .A(n49278), .B(n14134), .X(n14131) );
  nand_x1_sg U67269 ( .A(n13507), .B(n14133), .X(n14132) );
  nand_x1_sg U67270 ( .A(n39788), .B(n41820), .X(n14134) );
  nand_x1_sg U67271 ( .A(n49564), .B(n14953), .X(n14950) );
  nand_x1_sg U67272 ( .A(n14326), .B(n14952), .X(n14951) );
  nand_x1_sg U67273 ( .A(n39783), .B(n14481), .X(n14953) );
  nand_x1_sg U67274 ( .A(n49850), .B(n15772), .X(n15769) );
  nand_x1_sg U67275 ( .A(n15145), .B(n15771), .X(n15770) );
  nand_x1_sg U67276 ( .A(n39784), .B(n41817), .X(n15772) );
  nand_x1_sg U67277 ( .A(n50136), .B(n16591), .X(n16588) );
  nand_x1_sg U67278 ( .A(n15964), .B(n16590), .X(n16589) );
  nand_x1_sg U67279 ( .A(n39779), .B(n16119), .X(n16591) );
  nand_x1_sg U67280 ( .A(n50421), .B(n17408), .X(n17405) );
  nand_x1_sg U67281 ( .A(n16781), .B(n17407), .X(n17406) );
  nand_x1_sg U67282 ( .A(n39774), .B(n40231), .X(n17408) );
  nand_x1_sg U67283 ( .A(n50710), .B(n18229), .X(n18226) );
  nand_x1_sg U67284 ( .A(n17602), .B(n18228), .X(n18227) );
  nand_x1_sg U67285 ( .A(n39780), .B(n41811), .X(n18229) );
  nand_x1_sg U67286 ( .A(n50997), .B(n19050), .X(n19047) );
  nand_x1_sg U67287 ( .A(n18423), .B(n19049), .X(n19048) );
  nand_x1_sg U67288 ( .A(n39776), .B(n41812), .X(n19050) );
  inv_x1_sg U67289 ( .A(n22551), .X(n45018) );
  nand_x1_sg U67290 ( .A(n38932), .B(n21731), .X(n21730) );
  nand_x1_sg U67291 ( .A(n39258), .B(n21778), .X(n21777) );
  nand_x1_sg U67292 ( .A(n41099), .B(n21825), .X(n21824) );
  nand_x1_sg U67293 ( .A(n41099), .B(n21872), .X(n21871) );
  nand_x1_sg U67294 ( .A(n41097), .B(n21918), .X(n21917) );
  nand_x1_sg U67295 ( .A(n38932), .B(n21965), .X(n21964) );
  nand_x1_sg U67296 ( .A(n41099), .B(n22011), .X(n22010) );
  nand_x1_sg U67297 ( .A(n38932), .B(n22058), .X(n22057) );
  nand_x1_sg U67298 ( .A(n19126), .B(n22104), .X(n22103) );
  nand_x1_sg U67299 ( .A(n41098), .B(n22152), .X(n22151) );
  nand_x1_sg U67300 ( .A(n41097), .B(n22199), .X(n22198) );
  nand_x1_sg U67301 ( .A(n19126), .B(n22247), .X(n22246) );
  nand_x1_sg U67302 ( .A(n41098), .B(n22294), .X(n22293) );
  nand_x1_sg U67303 ( .A(n39258), .B(n22342), .X(n22341) );
  nand_x1_sg U67304 ( .A(n41098), .B(n22389), .X(n22388) );
  nand_x1_sg U67305 ( .A(n39258), .B(n22437), .X(n22436) );
  nand_x1_sg U67306 ( .A(n41098), .B(n22483), .X(n22482) );
  nand_x1_sg U67307 ( .A(n39258), .B(n45003), .X(n22528) );
  nand_x1_sg U67308 ( .A(n47120), .B(n22714), .X(n7009) );
  nor_x1_sg U67309 ( .A(n40927), .B(n16652), .X(\L2_0/n2560 ) );
  nand_x1_sg U67310 ( .A(n39664), .B(n40574), .X(n6993) );
  nand_x1_sg U67311 ( .A(n42358), .B(n40631), .X(n7810) );
  nand_x1_sg U67312 ( .A(n42357), .B(n40626), .X(n8628) );
  nand_x1_sg U67313 ( .A(n42368), .B(n40668), .X(n9448) );
  nand_x1_sg U67314 ( .A(n42367), .B(n40658), .X(n10267) );
  nand_x1_sg U67315 ( .A(n42366), .B(n40642), .X(n11086) );
  nand_x1_sg U67316 ( .A(n42365), .B(n40638), .X(n11905) );
  nand_x1_sg U67317 ( .A(n42364), .B(n40664), .X(n12724) );
  nand_x1_sg U67318 ( .A(n42363), .B(n40653), .X(n13543) );
  nand_x1_sg U67319 ( .A(n42362), .B(n40624), .X(n14362) );
  nand_x1_sg U67320 ( .A(n42361), .B(n40684), .X(n15181) );
  nand_x1_sg U67321 ( .A(n42360), .B(n40678), .X(n16000) );
  nand_x1_sg U67322 ( .A(n17636), .B(n40646), .X(n17638) );
  nand_x1_sg U67323 ( .A(n42359), .B(n40673), .X(n18459) );
  nand_x1_sg U67324 ( .A(n40076), .B(n25960), .X(n25959) );
  nor_x1_sg U67325 ( .A(n40038), .B(n25951), .X(n25960) );
  nor_x1_sg U67326 ( .A(n15828), .B(n15836), .X(\L2_0/n2640 ) );
  nor_x1_sg U67327 ( .A(n38904), .B(n9284), .X(\L2_0/n3280 ) );
  nor_x1_sg U67328 ( .A(n38902), .B(n10103), .X(\L2_0/n3200 ) );
  nor_x1_sg U67329 ( .A(n10914), .B(n10922), .X(\L2_0/n3120 ) );
  nor_x1_sg U67330 ( .A(n38895), .B(n11741), .X(\L2_0/n3040 ) );
  nor_x1_sg U67331 ( .A(n38896), .B(n12560), .X(\L2_0/n2960 ) );
  nor_x1_sg U67332 ( .A(n40942), .B(n13379), .X(\L2_0/n2880 ) );
  nor_x1_sg U67333 ( .A(n38898), .B(n14198), .X(\L2_0/n2800 ) );
  nor_x1_sg U67334 ( .A(n38899), .B(n15017), .X(\L2_0/n2720 ) );
  nor_x1_sg U67335 ( .A(n38901), .B(n18295), .X(\L2_0/n2400 ) );
  nand_x1_sg U67336 ( .A(n39662), .B(n40564), .X(n17451) );
  nand_x1_sg U67337 ( .A(n16815), .B(n40578), .X(n16817) );
  nand_x1_sg U67338 ( .A(n16815), .B(n25992), .X(n25991) );
  nor_x1_sg U67339 ( .A(n40038), .B(n25984), .X(n25992) );
  nand_x1_sg U67340 ( .A(n17299), .B(n26005), .X(n26004) );
  nor_x1_sg U67341 ( .A(n42370), .B(n25997), .X(n26005) );
  inv_x1_sg U67342 ( .A(n20310), .X(n46424) );
  nor_x1_sg U67343 ( .A(n40966), .B(n17474), .X(\L2_0/n2480 ) );
  inv_x1_sg U67344 ( .A(n21267), .X(n45875) );
  inv_x1_sg U67345 ( .A(n20498), .X(n45878) );
  inv_x1_sg U67346 ( .A(n19841), .X(n45881) );
  nand_x1_sg U67347 ( .A(n8383), .B(n41834), .X(n8439) );
  nand_x1_sg U67348 ( .A(n9201), .B(n41832), .X(n9257) );
  nand_x1_sg U67349 ( .A(n10021), .B(n41831), .X(n10077) );
  nand_x1_sg U67350 ( .A(n10840), .B(n41828), .X(n10896) );
  nand_x1_sg U67351 ( .A(n11659), .B(n41826), .X(n11715) );
  nand_x1_sg U67352 ( .A(n12478), .B(n41824), .X(n12534) );
  nand_x1_sg U67353 ( .A(n13297), .B(n41823), .X(n13353) );
  nand_x1_sg U67354 ( .A(n14116), .B(n41821), .X(n14172) );
  nand_x1_sg U67355 ( .A(n14935), .B(n41819), .X(n14991) );
  nand_x1_sg U67356 ( .A(n15754), .B(n41816), .X(n15810) );
  nand_x1_sg U67357 ( .A(n16573), .B(n41815), .X(n16629) );
  nand_x1_sg U67358 ( .A(n18211), .B(n41811), .X(n18267) );
  nand_x1_sg U67359 ( .A(n19032), .B(n41813), .X(n19088) );
  nand_x1_sg U67360 ( .A(n8161), .B(n41835), .X(n8182) );
  nand_x1_sg U67361 ( .A(n8979), .B(n41833), .X(n9000) );
  nand_x1_sg U67362 ( .A(n9799), .B(n41831), .X(n9820) );
  nand_x1_sg U67363 ( .A(n10618), .B(n41829), .X(n10639) );
  nand_x1_sg U67364 ( .A(n11437), .B(n41827), .X(n11458) );
  nand_x1_sg U67365 ( .A(n12256), .B(n41825), .X(n12277) );
  nand_x1_sg U67366 ( .A(n13075), .B(n41822), .X(n13096) );
  nand_x1_sg U67367 ( .A(n13894), .B(n41821), .X(n13915) );
  nand_x1_sg U67368 ( .A(n14713), .B(n41818), .X(n14734) );
  nand_x1_sg U67369 ( .A(n15532), .B(n41817), .X(n15553) );
  nand_x1_sg U67370 ( .A(n16351), .B(n41814), .X(n16372) );
  nand_x1_sg U67371 ( .A(n17989), .B(n41810), .X(n18010) );
  nand_x1_sg U67372 ( .A(n18810), .B(n41813), .X(n18831) );
  inv_x1_sg U67373 ( .A(n22702), .X(n47127) );
  nand_x1_sg U67374 ( .A(n17390), .B(n40229), .X(n17446) );
  nand_x1_sg U67375 ( .A(n17168), .B(n40229), .X(n17189) );
  nand_x1_sg U67376 ( .A(n7565), .B(n40235), .X(n7621) );
  nand_x1_sg U67377 ( .A(n7343), .B(n40233), .X(n7364) );
  nor_x1_sg U67378 ( .A(n6822), .B(n6828), .X(\L2_0/n3520 ) );
  inv_x1_sg U67379 ( .A(n22714), .X(n47096) );
  nand_x1_sg U67380 ( .A(n39520), .B(n25980), .X(n25979) );
  nor_x1_sg U67381 ( .A(n40037), .B(n25971), .X(n25980) );
  nand_x1_sg U67382 ( .A(n39772), .B(n22655), .X(n22654) );
  nor_x1_sg U67383 ( .A(n22638), .B(n46938), .X(n22655) );
  nand_x1_sg U67384 ( .A(n38921), .B(n26766), .X(n26763) );
  nand_x1_sg U67385 ( .A(n38906), .B(n21732), .X(n21729) );
  nand_x1_sg U67386 ( .A(n40986), .B(n21779), .X(n21776) );
  nand_x1_sg U67387 ( .A(n40988), .B(n21826), .X(n21823) );
  nand_x1_sg U67388 ( .A(n38906), .B(n21873), .X(n21870) );
  nand_x1_sg U67389 ( .A(n38906), .B(n21919), .X(n21916) );
  nand_x1_sg U67390 ( .A(n40986), .B(n21966), .X(n21963) );
  nand_x1_sg U67391 ( .A(n40988), .B(n22012), .X(n22009) );
  nand_x1_sg U67392 ( .A(n40986), .B(n22059), .X(n22056) );
  nand_x1_sg U67393 ( .A(n40987), .B(n22105), .X(n22102) );
  nand_x1_sg U67394 ( .A(n38920), .B(n22153), .X(n22150) );
  nand_x1_sg U67395 ( .A(n40987), .B(n22200), .X(n22197) );
  nand_x1_sg U67396 ( .A(n40986), .B(n22248), .X(n22245) );
  nand_x1_sg U67397 ( .A(n38921), .B(n22295), .X(n22292) );
  nand_x1_sg U67398 ( .A(n40987), .B(n22343), .X(n22340) );
  nand_x1_sg U67399 ( .A(n38906), .B(n22390), .X(n22387) );
  nand_x1_sg U67400 ( .A(n40987), .B(n22438), .X(n22435) );
  nand_x1_sg U67401 ( .A(n38920), .B(n22484), .X(n22481) );
  inv_x1_sg U67402 ( .A(n19507), .X(n46528) );
  inv_x1_sg U67403 ( .A(n19916), .X(n46445) );
  inv_x1_sg U67404 ( .A(n19951), .X(n46474) );
  inv_x1_sg U67405 ( .A(n19767), .X(n46516) );
  nand_x1_sg U67406 ( .A(n40130), .B(n39134), .X(n25968) );
  nand_x1_sg U67407 ( .A(n39775), .B(n40563), .X(n17362) );
  nand_x1_sg U67408 ( .A(n39806), .B(n40564), .X(n16827) );
  inv_x1_sg U67409 ( .A(n8004), .X(n47198) );
  inv_x1_sg U67410 ( .A(n8822), .X(n47483) );
  inv_x1_sg U67411 ( .A(n9642), .X(n47768) );
  inv_x1_sg U67412 ( .A(n10461), .X(n48053) );
  inv_x1_sg U67413 ( .A(n11280), .X(n48338) );
  inv_x1_sg U67414 ( .A(n12099), .X(n48623) );
  inv_x1_sg U67415 ( .A(n12918), .X(n48909) );
  inv_x1_sg U67416 ( .A(n13737), .X(n49196) );
  inv_x1_sg U67417 ( .A(n14556), .X(n49482) );
  inv_x1_sg U67418 ( .A(n15375), .X(n49768) );
  inv_x1_sg U67419 ( .A(n16194), .X(n50054) );
  inv_x1_sg U67420 ( .A(n17010), .X(n50339) );
  inv_x1_sg U67421 ( .A(n17832), .X(n50628) );
  inv_x1_sg U67422 ( .A(n18653), .X(n50915) );
  inv_x1_sg U67423 ( .A(n26029), .X(n50555) );
  inv_x1_sg U67424 ( .A(n7601), .X(n47078) );
  inv_x1_sg U67425 ( .A(n8419), .X(n47364) );
  inv_x1_sg U67426 ( .A(n9237), .X(n47649) );
  inv_x1_sg U67427 ( .A(n10057), .X(n47934) );
  inv_x1_sg U67428 ( .A(n10876), .X(n48219) );
  inv_x1_sg U67429 ( .A(n11695), .X(n48504) );
  inv_x1_sg U67430 ( .A(n12514), .X(n48789) );
  inv_x1_sg U67431 ( .A(n13333), .X(n49076) );
  inv_x1_sg U67432 ( .A(n14152), .X(n49362) );
  inv_x1_sg U67433 ( .A(n14971), .X(n49648) );
  inv_x1_sg U67434 ( .A(n15790), .X(n49934) );
  inv_x1_sg U67435 ( .A(n16609), .X(n50220) );
  inv_x1_sg U67436 ( .A(n18247), .X(n50794) );
  inv_x1_sg U67437 ( .A(n19068), .X(n51081) );
  inv_x1_sg U67438 ( .A(n8261), .X(n47298) );
  inv_x1_sg U67439 ( .A(n9079), .X(n47583) );
  inv_x1_sg U67440 ( .A(n9899), .X(n47868) );
  inv_x1_sg U67441 ( .A(n10718), .X(n48153) );
  inv_x1_sg U67442 ( .A(n11537), .X(n48438) );
  inv_x1_sg U67443 ( .A(n12356), .X(n48723) );
  inv_x1_sg U67444 ( .A(n13175), .X(n49009) );
  inv_x1_sg U67445 ( .A(n13994), .X(n49296) );
  inv_x1_sg U67446 ( .A(n14813), .X(n49582) );
  inv_x1_sg U67447 ( .A(n15632), .X(n49868) );
  inv_x1_sg U67448 ( .A(n16451), .X(n50154) );
  inv_x1_sg U67449 ( .A(n18089), .X(n50728) );
  inv_x1_sg U67450 ( .A(n18910), .X(n51015) );
  inv_x1_sg U67451 ( .A(n17426), .X(n50505) );
  inv_x1_sg U67452 ( .A(n17268), .X(n50439) );
  nor_x1_sg U67453 ( .A(n41057), .B(n38892), .X(\L2_0/n3532 ) );
  nor_x1_sg U67454 ( .A(n41057), .B(n39090), .X(\L1_0/n4436 ) );
  inv_x1_sg U67455 ( .A(n7443), .X(n47010) );
  inv_x1_sg U67456 ( .A(n7185), .X(n46905) );
  nor_x1_sg U67457 ( .A(n39963), .B(n7638), .X(\L2_0/n3452 ) );
  nor_x1_sg U67458 ( .A(n41928), .B(n40844), .X(\L2_0/n3372 ) );
  nor_x1_sg U67459 ( .A(n41927), .B(n40970), .X(\L2_0/n3292 ) );
  nor_x1_sg U67460 ( .A(n39975), .B(n40961), .X(\L2_0/n3212 ) );
  nor_x1_sg U67461 ( .A(n39979), .B(n40930), .X(\L2_0/n3132 ) );
  nor_x1_sg U67462 ( .A(n41924), .B(n38895), .X(\L2_0/n3052 ) );
  nor_x1_sg U67463 ( .A(n39987), .B(n40938), .X(\L2_0/n2972 ) );
  nor_x1_sg U67464 ( .A(n39992), .B(n13371), .X(\L2_0/n2892 ) );
  nor_x1_sg U67465 ( .A(n39997), .B(n40946), .X(\L2_0/n2812 ) );
  nor_x1_sg U67466 ( .A(n40000), .B(n38899), .X(\L2_0/n2732 ) );
  nor_x1_sg U67467 ( .A(n40003), .B(n40954), .X(\L2_0/n2652 ) );
  nor_x1_sg U67468 ( .A(n41000), .B(n38903), .X(\L2_0/n2492 ) );
  nor_x1_sg U67469 ( .A(n40009), .B(n38901), .X(\L2_0/n2412 ) );
  nor_x1_sg U67470 ( .A(n40993), .B(n40927), .X(\L2_0/n2572 ) );
  nand_x1_sg U67471 ( .A(n39812), .B(n42185), .X(n8103) );
  nand_x1_sg U67472 ( .A(n41887), .B(n42183), .X(n8921) );
  nand_x1_sg U67473 ( .A(n41878), .B(n42181), .X(n9741) );
  nand_x1_sg U67474 ( .A(n39816), .B(n42179), .X(n10560) );
  nand_x1_sg U67475 ( .A(n39834), .B(n42177), .X(n11379) );
  nand_x1_sg U67476 ( .A(n39836), .B(n42175), .X(n12198) );
  nand_x1_sg U67477 ( .A(n41896), .B(n42173), .X(n13017) );
  nand_x1_sg U67478 ( .A(n39839), .B(n42171), .X(n13836) );
  nand_x1_sg U67479 ( .A(n41880), .B(n42169), .X(n14655) );
  nand_x1_sg U67480 ( .A(n39849), .B(n42168), .X(n15474) );
  nand_x1_sg U67481 ( .A(n39821), .B(n42166), .X(n16293) );
  nand_x1_sg U67482 ( .A(n39827), .B(n17800), .X(n17931) );
  nand_x1_sg U67483 ( .A(n41892), .B(n40156), .X(n18752) );
  nor_x1_sg U67484 ( .A(n40982), .B(n5758), .X(n5125) );
  nor_x1_sg U67485 ( .A(n40994), .B(n39282), .X(n5758) );
  nor_x1_sg U67486 ( .A(n5972), .B(n5973), .X(n5971) );
  nor_x1_sg U67487 ( .A(n5984), .B(n5985), .X(n5970) );
  nor_x1_sg U67488 ( .A(n5976), .B(n39124), .X(n5972) );
  nor_x1_sg U67489 ( .A(n6122), .B(n6123), .X(n6121) );
  nor_x1_sg U67490 ( .A(n6132), .B(n6133), .X(n6120) );
  nor_x1_sg U67491 ( .A(n6124), .B(n41276), .X(n6122) );
  nor_x1_sg U67492 ( .A(n6260), .B(n6261), .X(n6259) );
  nor_x1_sg U67493 ( .A(n6269), .B(n6270), .X(n6258) );
  nor_x1_sg U67494 ( .A(n6263), .B(n41277), .X(n6260) );
  nor_x1_sg U67495 ( .A(n6394), .B(n6395), .X(n6393) );
  nor_x1_sg U67496 ( .A(n6403), .B(n6404), .X(n6392) );
  nor_x1_sg U67497 ( .A(n6397), .B(n5977), .X(n6394) );
  nor_x1_sg U67498 ( .A(n6527), .B(n6528), .X(n6526) );
  nor_x1_sg U67499 ( .A(n6536), .B(n6537), .X(n6525) );
  nor_x1_sg U67500 ( .A(n6530), .B(n5977), .X(n6527) );
  nor_x1_sg U67501 ( .A(n6662), .B(n6663), .X(n6661) );
  nor_x1_sg U67502 ( .A(n6672), .B(n6673), .X(n6660) );
  nor_x1_sg U67503 ( .A(n6665), .B(n39123), .X(n6662) );
  nor_x1_sg U67504 ( .A(n5966), .B(n5967), .X(n5960) );
  nor_x1_sg U67505 ( .A(n5962), .B(n5963), .X(n5961) );
  nor_x1_sg U67506 ( .A(n5969), .B(n41009), .X(n5966) );
  nand_x1_sg U67507 ( .A(n40100), .B(n5995), .X(n5993) );
  nor_x1_sg U67508 ( .A(n5996), .B(n5997), .X(n5992) );
  nor_x1_sg U67509 ( .A(n42260), .B(n41019), .X(n5997) );
  nor_x1_sg U67510 ( .A(n6027), .B(n6028), .X(n6026) );
  nor_x1_sg U67511 ( .A(n6036), .B(n6037), .X(n6025) );
  nor_x1_sg U67512 ( .A(n6029), .B(n5977), .X(n6027) );
  nor_x1_sg U67513 ( .A(n6075), .B(n6076), .X(n6074) );
  nor_x1_sg U67514 ( .A(n6085), .B(n6086), .X(n6073) );
  nor_x1_sg U67515 ( .A(n6078), .B(n39124), .X(n6075) );
  nand_x1_sg U67516 ( .A(n39149), .B(n6093), .X(n6092) );
  nor_x1_sg U67517 ( .A(n6094), .B(n6095), .X(n6091) );
  nor_x1_sg U67518 ( .A(n41969), .B(n41020), .X(n6095) );
  nand_x1_sg U67519 ( .A(n39148), .B(n46465), .X(n6138) );
  nor_x1_sg U67520 ( .A(n6139), .B(n6140), .X(n6137) );
  nor_x1_sg U67521 ( .A(n42275), .B(n41018), .X(n6140) );
  nor_x1_sg U67522 ( .A(n6167), .B(n6168), .X(n6166) );
  nor_x1_sg U67523 ( .A(n6177), .B(n6178), .X(n6165) );
  nor_x1_sg U67524 ( .A(n6170), .B(n41276), .X(n6167) );
  nand_x1_sg U67525 ( .A(n40095), .B(n6184), .X(n6183) );
  nor_x1_sg U67526 ( .A(n6185), .B(n6186), .X(n6182) );
  nor_x1_sg U67527 ( .A(n42274), .B(n41018), .X(n6186) );
  nor_x1_sg U67528 ( .A(n6214), .B(n6215), .X(n6213) );
  nor_x1_sg U67529 ( .A(n6224), .B(n6225), .X(n6212) );
  nor_x1_sg U67530 ( .A(n6217), .B(n41278), .X(n6214) );
  nand_x1_sg U67531 ( .A(n41398), .B(n46370), .X(n6230) );
  nor_x1_sg U67532 ( .A(n6231), .B(n6232), .X(n6229) );
  nor_x1_sg U67533 ( .A(n42273), .B(n41020), .X(n6232) );
  nand_x1_sg U67534 ( .A(n41395), .B(n6275), .X(n6274) );
  nor_x1_sg U67535 ( .A(n6276), .B(n6277), .X(n6273) );
  nor_x1_sg U67536 ( .A(n42272), .B(n41019), .X(n6277) );
  nand_x1_sg U67537 ( .A(n39148), .B(n46283), .X(n6319) );
  nor_x1_sg U67538 ( .A(n6320), .B(n6321), .X(n6318) );
  nor_x1_sg U67539 ( .A(n42271), .B(n38935), .X(n6321) );
  nand_x1_sg U67540 ( .A(n40095), .B(n6364), .X(n6363) );
  nor_x1_sg U67541 ( .A(n6365), .B(n6366), .X(n6362) );
  nor_x1_sg U67542 ( .A(n42270), .B(n41021), .X(n6366) );
  nand_x1_sg U67543 ( .A(n41397), .B(n46192), .X(n6408) );
  nor_x1_sg U67544 ( .A(n6409), .B(n6410), .X(n6407) );
  nor_x1_sg U67545 ( .A(n42269), .B(n41018), .X(n6410) );
  nand_x1_sg U67546 ( .A(n41396), .B(n6453), .X(n6452) );
  nor_x1_sg U67547 ( .A(n6454), .B(n6455), .X(n6451) );
  nor_x1_sg U67548 ( .A(n42267), .B(n41019), .X(n6455) );
  nand_x1_sg U67549 ( .A(n39149), .B(n46101), .X(n6497) );
  nor_x1_sg U67550 ( .A(n6498), .B(n6499), .X(n6496) );
  nor_x1_sg U67551 ( .A(n42266), .B(n41570), .X(n6499) );
  nand_x1_sg U67552 ( .A(n41396), .B(n6542), .X(n6541) );
  nor_x1_sg U67553 ( .A(n6543), .B(n6544), .X(n6540) );
  nor_x1_sg U67554 ( .A(n42265), .B(n41018), .X(n6544) );
  nand_x1_sg U67555 ( .A(n40099), .B(n46010), .X(n6586) );
  nor_x1_sg U67556 ( .A(n6587), .B(n6588), .X(n6585) );
  nor_x1_sg U67557 ( .A(n42264), .B(n41021), .X(n6588) );
  nand_x1_sg U67558 ( .A(n40100), .B(n6631), .X(n6630) );
  nor_x1_sg U67559 ( .A(n6632), .B(n6633), .X(n6629) );
  nor_x1_sg U67560 ( .A(n42263), .B(n41570), .X(n6633) );
  nand_x1_sg U67561 ( .A(n39148), .B(n6043), .X(n6042) );
  nor_x1_sg U67562 ( .A(n6044), .B(n6045), .X(n6041) );
  nor_x1_sg U67563 ( .A(n41968), .B(n41021), .X(n6045) );
  nand_x1_sg U67564 ( .A(n40100), .B(n45919), .X(n6678) );
  nor_x1_sg U67565 ( .A(n6679), .B(n6680), .X(n6677) );
  nor_x1_sg U67566 ( .A(n42302), .B(n41569), .X(n6679) );
  nor_x1_sg U67567 ( .A(n19129), .B(n19130), .X(n19128) );
  nor_x1_sg U67568 ( .A(n19508), .B(n19509), .X(n19127) );
  nor_x1_sg U67569 ( .A(n19132), .B(n41276), .X(n19129) );
  nor_x1_sg U67570 ( .A(n6305), .B(n6306), .X(n6304) );
  nor_x1_sg U67571 ( .A(n6314), .B(n6315), .X(n6303) );
  nor_x1_sg U67572 ( .A(n6308), .B(n41278), .X(n6305) );
  nor_x1_sg U67573 ( .A(n6349), .B(n6350), .X(n6348) );
  nor_x1_sg U67574 ( .A(n6358), .B(n6359), .X(n6347) );
  nor_x1_sg U67575 ( .A(n6352), .B(n41277), .X(n6349) );
  nor_x1_sg U67576 ( .A(n6438), .B(n6439), .X(n6437) );
  nor_x1_sg U67577 ( .A(n6447), .B(n6448), .X(n6436) );
  nor_x1_sg U67578 ( .A(n6441), .B(n39124), .X(n6438) );
  nor_x1_sg U67579 ( .A(n6483), .B(n6484), .X(n6482) );
  nor_x1_sg U67580 ( .A(n6492), .B(n6493), .X(n6481) );
  nor_x1_sg U67581 ( .A(n6486), .B(n41278), .X(n6483) );
  nor_x1_sg U67582 ( .A(n6572), .B(n6573), .X(n6571) );
  nor_x1_sg U67583 ( .A(n6581), .B(n6582), .X(n6570) );
  nor_x1_sg U67584 ( .A(n6575), .B(n41278), .X(n6572) );
  nor_x1_sg U67585 ( .A(n6616), .B(n6617), .X(n6615) );
  nor_x1_sg U67586 ( .A(n6625), .B(n6626), .X(n6614) );
  nor_x1_sg U67587 ( .A(n6619), .B(n41277), .X(n6616) );
  nor_x1_sg U67588 ( .A(n6707), .B(n6708), .X(n6706) );
  nor_x1_sg U67589 ( .A(n6717), .B(n6718), .X(n6705) );
  nor_x1_sg U67590 ( .A(n41530), .B(n41254), .X(n6708) );
  nor_x1_sg U67591 ( .A(n6751), .B(n6752), .X(n6750) );
  nor_x1_sg U67592 ( .A(n6761), .B(n6762), .X(n6749) );
  nor_x1_sg U67593 ( .A(n6754), .B(n39123), .X(n6751) );
  nor_x1_sg U67594 ( .A(n6745), .B(n6746), .X(n6739) );
  nor_x1_sg U67595 ( .A(n6741), .B(n6742), .X(n6740) );
  nor_x1_sg U67596 ( .A(n6748), .B(n38931), .X(n6745) );
  nand_x1_sg U67597 ( .A(n40098), .B(n45814), .X(n6768) );
  nor_x1_sg U67598 ( .A(n6769), .B(n6770), .X(n6767) );
  nor_x1_sg U67599 ( .A(n6772), .B(n41023), .X(n6769) );
  nor_x1_sg U67600 ( .A(n6779), .B(n6780), .X(n6773) );
  nor_x1_sg U67601 ( .A(n6775), .B(n6776), .X(n6774) );
  nor_x1_sg U67602 ( .A(n6782), .B(n41036), .X(n6779) );
  nor_x1_sg U67603 ( .A(n19121), .B(n19122), .X(n19113) );
  nor_x1_sg U67604 ( .A(n19115), .B(n19116), .X(n19114) );
  nor_x1_sg U67605 ( .A(n19125), .B(n41572), .X(n19121) );
  nand_x1_sg U67606 ( .A(n39149), .B(n20563), .X(n20562) );
  nor_x1_sg U67607 ( .A(n20564), .B(n20565), .X(n20561) );
  nor_x1_sg U67608 ( .A(n20568), .B(n41024), .X(n20564) );
  nor_x1_sg U67609 ( .A(n20958), .B(n20959), .X(n20570) );
  nor_x1_sg U67610 ( .A(n20572), .B(n20573), .X(n20571) );
  nor_x1_sg U67611 ( .A(n20580), .B(n41033), .X(n20958) );
  nand_x1_sg U67612 ( .A(n41395), .B(n6723), .X(n6722) );
  nor_x1_sg U67613 ( .A(n6724), .B(n6725), .X(n6721) );
  nor_x1_sg U67614 ( .A(n45875), .B(n41019), .X(n6725) );
  nor_x1_sg U67615 ( .A(n6795), .B(n6796), .X(n6790) );
  nor_x1_sg U67616 ( .A(n6792), .B(n6793), .X(n6791) );
  nor_x1_sg U67617 ( .A(n41011), .B(n45806), .X(n6795) );
  nand_x1_sg U67618 ( .A(n45798), .B(n41398), .X(n6811) );
  nor_x1_sg U67619 ( .A(n6812), .B(n6813), .X(n6810) );
  nor_x1_sg U67620 ( .A(n45799), .B(n41020), .X(n6813) );
  nor_x1_sg U67621 ( .A(n6819), .B(n6820), .X(n6814) );
  nor_x1_sg U67622 ( .A(n6816), .B(n6817), .X(n6815) );
  nor_x1_sg U67623 ( .A(n41035), .B(n45802), .X(n6819) );
  nor_x1_sg U67624 ( .A(n41127), .B(n26182), .X(\L1_0/n3392 ) );
  nor_x1_sg U67625 ( .A(n39248), .B(n26192), .X(\L1_0/n3388 ) );
  nor_x1_sg U67626 ( .A(n41128), .B(n26200), .X(\L1_0/n3384 ) );
  nor_x1_sg U67627 ( .A(n41127), .B(n26208), .X(\L1_0/n3380 ) );
  nor_x1_sg U67628 ( .A(n39249), .B(n26216), .X(\L1_0/n3376 ) );
  nor_x1_sg U67629 ( .A(n41127), .B(n26224), .X(\L1_0/n3372 ) );
  nor_x1_sg U67630 ( .A(n41128), .B(n26248), .X(\L1_0/n3360 ) );
  nor_x1_sg U67631 ( .A(n41130), .B(n26264), .X(\L1_0/n3352 ) );
  nor_x1_sg U67632 ( .A(n39248), .B(n26280), .X(\L1_0/n3344 ) );
  nor_x1_sg U67633 ( .A(n41129), .B(n26296), .X(\L1_0/n3336 ) );
  nor_x1_sg U67634 ( .A(n41130), .B(n26304), .X(\L1_0/n3332 ) );
  nor_x1_sg U67635 ( .A(n41129), .B(n26310), .X(\L1_0/n3328 ) );
  nor_x1_sg U67636 ( .A(n41129), .B(n26318), .X(\L1_0/n3324 ) );
  nand_x1_sg U67637 ( .A(n39255), .B(n21751), .X(n21750) );
  nand_x1_sg U67638 ( .A(n39261), .B(n21752), .X(n21749) );
  nand_x1_sg U67639 ( .A(n41110), .B(n21845), .X(n21844) );
  nand_x1_sg U67640 ( .A(n38926), .B(n21846), .X(n21843) );
  nand_x1_sg U67641 ( .A(n39255), .B(n21938), .X(n21937) );
  nand_x1_sg U67642 ( .A(n39261), .B(n21939), .X(n21936) );
  nand_x1_sg U67643 ( .A(n38938), .B(n22031), .X(n22030) );
  nand_x1_sg U67644 ( .A(n41086), .B(n22032), .X(n22029) );
  nand_x1_sg U67645 ( .A(n39255), .B(n22125), .X(n22124) );
  nand_x1_sg U67646 ( .A(n41085), .B(n22126), .X(n22123) );
  nand_x1_sg U67647 ( .A(n38938), .B(n22220), .X(n22219) );
  nand_x1_sg U67648 ( .A(n41087), .B(n22221), .X(n22218) );
  nand_x1_sg U67649 ( .A(n41109), .B(n22315), .X(n22314) );
  nand_x1_sg U67650 ( .A(n41087), .B(n22316), .X(n22313) );
  nand_x1_sg U67651 ( .A(n20569), .B(n22410), .X(n22409) );
  nand_x1_sg U67652 ( .A(n41085), .B(n22411), .X(n22408) );
  nand_x1_sg U67653 ( .A(n41086), .B(n22503), .X(n22500) );
  nand_x1_sg U67654 ( .A(n41110), .B(n26790), .X(n26789) );
  nand_x1_sg U67655 ( .A(n20575), .B(n26791), .X(n26788) );
  nand_x1_sg U67656 ( .A(n41109), .B(n21798), .X(n21797) );
  nand_x1_sg U67657 ( .A(n38926), .B(n21799), .X(n21796) );
  nand_x1_sg U67658 ( .A(n41111), .B(n21891), .X(n21890) );
  nand_x1_sg U67659 ( .A(n41086), .B(n21892), .X(n21889) );
  nand_x1_sg U67660 ( .A(n39255), .B(n21984), .X(n21983) );
  nand_x1_sg U67661 ( .A(n39261), .B(n21985), .X(n21982) );
  nand_x1_sg U67662 ( .A(n20569), .B(n22077), .X(n22076) );
  nand_x1_sg U67663 ( .A(n20575), .B(n22078), .X(n22075) );
  nand_x1_sg U67664 ( .A(n41111), .B(n22172), .X(n22171) );
  nand_x1_sg U67665 ( .A(n41087), .B(n22173), .X(n22170) );
  nand_x1_sg U67666 ( .A(n41111), .B(n22267), .X(n22266) );
  nand_x1_sg U67667 ( .A(n38926), .B(n22268), .X(n22265) );
  nand_x1_sg U67668 ( .A(n38938), .B(n22362), .X(n22361) );
  nand_x1_sg U67669 ( .A(n38926), .B(n22363), .X(n22360) );
  nand_x1_sg U67670 ( .A(n41086), .B(n22457), .X(n22454) );
  nand_x1_sg U67671 ( .A(n40746), .B(n26796), .X(n26795) );
  nand_x1_sg U67672 ( .A(n41122), .B(n26798), .X(n26794) );
  nand_x1_sg U67673 ( .A(n40746), .B(n21763), .X(n21754) );
  nand_x1_sg U67674 ( .A(n39251), .B(n21756), .X(n21755) );
  nand_x1_sg U67675 ( .A(n40747), .B(n21810), .X(n21801) );
  nand_x1_sg U67676 ( .A(n41123), .B(n21803), .X(n21802) );
  nand_x1_sg U67677 ( .A(n40748), .B(n21857), .X(n21848) );
  nand_x1_sg U67678 ( .A(n39252), .B(n21850), .X(n21849) );
  nand_x1_sg U67679 ( .A(n40747), .B(n21903), .X(n21894) );
  nand_x1_sg U67680 ( .A(n39252), .B(n21896), .X(n21895) );
  nand_x1_sg U67681 ( .A(n40746), .B(n21950), .X(n21941) );
  nand_x1_sg U67682 ( .A(n41123), .B(n21943), .X(n21942) );
  nand_x1_sg U67683 ( .A(n40749), .B(n21996), .X(n21987) );
  nand_x1_sg U67684 ( .A(n39252), .B(n21989), .X(n21988) );
  nand_x1_sg U67685 ( .A(n40746), .B(n22043), .X(n22034) );
  nand_x1_sg U67686 ( .A(n41122), .B(n22036), .X(n22035) );
  nand_x1_sg U67687 ( .A(n40747), .B(n22089), .X(n22080) );
  nand_x1_sg U67688 ( .A(n41125), .B(n22082), .X(n22081) );
  nand_x1_sg U67689 ( .A(n38829), .B(n22137), .X(n22128) );
  nand_x1_sg U67690 ( .A(n41123), .B(n22130), .X(n22129) );
  nand_x1_sg U67691 ( .A(n38829), .B(n22184), .X(n22175) );
  nand_x1_sg U67692 ( .A(n41122), .B(n22177), .X(n22176) );
  nand_x1_sg U67693 ( .A(n40748), .B(n22232), .X(n22223) );
  nand_x1_sg U67694 ( .A(n41123), .B(n22225), .X(n22224) );
  nand_x1_sg U67695 ( .A(n40747), .B(n22279), .X(n22270) );
  nand_x1_sg U67696 ( .A(n39251), .B(n22272), .X(n22271) );
  nand_x1_sg U67697 ( .A(n40748), .B(n22327), .X(n22318) );
  nand_x1_sg U67698 ( .A(n41125), .B(n22320), .X(n22319) );
  nand_x1_sg U67699 ( .A(n38829), .B(n22374), .X(n22365) );
  nand_x1_sg U67700 ( .A(n41125), .B(n22367), .X(n22366) );
  nand_x1_sg U67701 ( .A(n40749), .B(n22422), .X(n22413) );
  nand_x1_sg U67702 ( .A(n41124), .B(n22415), .X(n22414) );
  nand_x1_sg U67703 ( .A(n40748), .B(n22468), .X(n22459) );
  nand_x1_sg U67704 ( .A(n41124), .B(n22461), .X(n22460) );
  nand_x1_sg U67705 ( .A(n40749), .B(n22514), .X(n22505) );
  nand_x1_sg U67706 ( .A(n39251), .B(n22507), .X(n22506) );
  nand_x1_sg U67707 ( .A(n40749), .B(n22552), .X(n22543) );
  nand_x1_sg U67708 ( .A(n41124), .B(n22545), .X(n22544) );
  nand_x1_sg U67709 ( .A(n39262), .B(n26770), .X(n26769) );
  nand_x1_sg U67710 ( .A(n38924), .B(n21735), .X(n21734) );
  nand_x1_sg U67711 ( .A(n39257), .B(n21736), .X(n21733) );
  nand_x1_sg U67712 ( .A(n19120), .B(n21782), .X(n21781) );
  nand_x1_sg U67713 ( .A(n41102), .B(n21783), .X(n21780) );
  nand_x1_sg U67714 ( .A(n41081), .B(n21829), .X(n21828) );
  nand_x1_sg U67715 ( .A(n39257), .B(n21830), .X(n21827) );
  nand_x1_sg U67716 ( .A(n39262), .B(n21876), .X(n21875) );
  nand_x1_sg U67717 ( .A(n41082), .B(n21922), .X(n21921) );
  nand_x1_sg U67718 ( .A(n38924), .B(n21969), .X(n21968) );
  nand_x1_sg U67719 ( .A(n41082), .B(n22015), .X(n22014) );
  nand_x1_sg U67720 ( .A(n39262), .B(n22062), .X(n22061) );
  nand_x1_sg U67721 ( .A(n41081), .B(n22108), .X(n22107) );
  nand_x1_sg U67722 ( .A(n38924), .B(n22156), .X(n22155) );
  nand_x1_sg U67723 ( .A(n38924), .B(n22203), .X(n22202) );
  nand_x1_sg U67724 ( .A(n41083), .B(n22251), .X(n22250) );
  nand_x1_sg U67725 ( .A(n41083), .B(n22298), .X(n22297) );
  nand_x1_sg U67726 ( .A(n19120), .B(n22346), .X(n22345) );
  nand_x1_sg U67727 ( .A(n41083), .B(n22393), .X(n22392) );
  nand_x1_sg U67728 ( .A(n41082), .B(n22441), .X(n22440) );
  nand_x1_sg U67729 ( .A(n41103), .B(n45081), .X(n22439) );
  nand_x1_sg U67730 ( .A(n39262), .B(n22487), .X(n22486) );
  nand_x1_sg U67731 ( .A(n41103), .B(n45037), .X(n22485) );
  nand_x1_sg U67732 ( .A(n41082), .B(n45009), .X(n22530) );
  nand_x1_sg U67733 ( .A(n38934), .B(n45000), .X(n22529) );
  nand_x1_sg U67734 ( .A(n41083), .B(n38628), .X(n22568) );
  nand_x1_sg U67735 ( .A(n38934), .B(n42159), .X(n22567) );
  nor_x1_sg U67736 ( .A(n41068), .B(n19106), .X(\L2_0/n2292 ) );
  nor_x1_sg U67737 ( .A(n41067), .B(n5952), .X(\L2_0/n3608 ) );
  nor_x1_sg U67738 ( .A(n40024), .B(n6008), .X(\L2_0/n3604 ) );
  nor_x1_sg U67739 ( .A(n41067), .B(n6057), .X(\L2_0/n3600 ) );
  nor_x1_sg U67740 ( .A(n41069), .B(n6105), .X(\L2_0/n3596 ) );
  nor_x1_sg U67741 ( .A(n39265), .B(n6150), .X(\L2_0/n3592 ) );
  nor_x1_sg U67742 ( .A(n41068), .B(n6196), .X(\L2_0/n3588 ) );
  nor_x1_sg U67743 ( .A(n41068), .B(n6243), .X(\L2_0/n3584 ) );
  nor_x1_sg U67744 ( .A(n41069), .B(n6288), .X(\L2_0/n3580 ) );
  nor_x1_sg U67745 ( .A(n41068), .B(n6332), .X(\L2_0/n3576 ) );
  nor_x1_sg U67746 ( .A(n41069), .B(n6377), .X(\L2_0/n3572 ) );
  nor_x1_sg U67747 ( .A(n39265), .B(n6421), .X(\L2_0/n3568 ) );
  nor_x1_sg U67748 ( .A(n41066), .B(n6466), .X(\L2_0/n3564 ) );
  nor_x1_sg U67749 ( .A(n39265), .B(n6510), .X(\L2_0/n3560 ) );
  nor_x1_sg U67750 ( .A(n39265), .B(n6555), .X(\L2_0/n3556 ) );
  nor_x1_sg U67751 ( .A(n41067), .B(n6599), .X(\L2_0/n3552 ) );
  nor_x1_sg U67752 ( .A(n41067), .B(n6644), .X(\L2_0/n3548 ) );
  nor_x1_sg U67753 ( .A(n41066), .B(n6692), .X(\L2_0/n3544 ) );
  nor_x1_sg U67754 ( .A(n41066), .B(n6732), .X(\L2_0/n3540 ) );
  nor_x1_sg U67755 ( .A(n41069), .B(n6783), .X(\L2_0/n3536 ) );
  nand_x1_sg U67756 ( .A(n40918), .B(n7640), .X(\L2_0/n3451 ) );
  nand_x1_sg U67757 ( .A(n39965), .B(n41288), .X(n7640) );
  nand_x1_sg U67758 ( .A(n40917), .B(n7644), .X(\L2_0/n3443 ) );
  nand_x1_sg U67759 ( .A(n7645), .B(n41285), .X(n7644) );
  nand_x1_sg U67760 ( .A(n39964), .B(n40157), .X(n7645) );
  nand_x1_sg U67761 ( .A(n40919), .B(n7647), .X(\L2_0/n3439 ) );
  nand_x1_sg U67762 ( .A(n41285), .B(n7646), .X(n7647) );
  nand_x1_sg U67763 ( .A(n40916), .B(n7653), .X(\L2_0/n3435 ) );
  nand_x1_sg U67764 ( .A(n7652), .B(n41288), .X(n7653) );
  nand_x1_sg U67765 ( .A(n40919), .B(n7660), .X(\L2_0/n3431 ) );
  nand_x1_sg U67766 ( .A(n41288), .B(n7659), .X(n7660) );
  nand_x1_sg U67767 ( .A(n40918), .B(n7667), .X(\L2_0/n3427 ) );
  nand_x1_sg U67768 ( .A(n7666), .B(n41285), .X(n7667) );
  nand_x1_sg U67769 ( .A(n38891), .B(n7673), .X(\L2_0/n3423 ) );
  nand_x1_sg U67770 ( .A(n7672), .B(n39129), .X(n7673) );
  nand_x1_sg U67771 ( .A(n40917), .B(n7679), .X(\L2_0/n3419 ) );
  nand_x1_sg U67772 ( .A(n7678), .B(n41285), .X(n7679) );
  nand_x1_sg U67773 ( .A(n40919), .B(n7685), .X(\L2_0/n3415 ) );
  nand_x1_sg U67774 ( .A(n7684), .B(n41286), .X(n7685) );
  nand_x1_sg U67775 ( .A(n40917), .B(n7691), .X(\L2_0/n3411 ) );
  nand_x1_sg U67776 ( .A(n7690), .B(n39130), .X(n7691) );
  nand_x1_sg U67777 ( .A(n40917), .B(n7697), .X(\L2_0/n3407 ) );
  nand_x1_sg U67778 ( .A(n7696), .B(n41286), .X(n7697) );
  nand_x1_sg U67779 ( .A(n40918), .B(n7703), .X(\L2_0/n3403 ) );
  nand_x1_sg U67780 ( .A(n7702), .B(n41286), .X(n7703) );
  nand_x1_sg U67781 ( .A(n40916), .B(n7709), .X(\L2_0/n3399 ) );
  nand_x1_sg U67782 ( .A(n7708), .B(n41287), .X(n7709) );
  nand_x1_sg U67783 ( .A(n40919), .B(n7715), .X(\L2_0/n3395 ) );
  nand_x1_sg U67784 ( .A(n7714), .B(n39130), .X(n7715) );
  nand_x1_sg U67785 ( .A(n38891), .B(n7721), .X(\L2_0/n3391 ) );
  nand_x1_sg U67786 ( .A(n7720), .B(n41287), .X(n7721) );
  nand_x1_sg U67787 ( .A(n40916), .B(n7727), .X(\L2_0/n3387 ) );
  nand_x1_sg U67788 ( .A(n7726), .B(n41287), .X(n7727) );
  nand_x1_sg U67789 ( .A(n40916), .B(n7733), .X(\L2_0/n3383 ) );
  nand_x1_sg U67790 ( .A(n7732), .B(n39129), .X(n7733) );
  nand_x1_sg U67791 ( .A(n40918), .B(n7739), .X(\L2_0/n3379 ) );
  nand_x1_sg U67792 ( .A(n7738), .B(n39130), .X(n7739) );
  nand_x1_sg U67793 ( .A(n38891), .B(n7745), .X(\L2_0/n3375 ) );
  nand_x1_sg U67794 ( .A(n7744), .B(n41288), .X(n7745) );
  nand_x1_sg U67795 ( .A(n40990), .B(n26780), .X(n26775) );
  nand_x1_sg U67796 ( .A(n40991), .B(n21742), .X(n21739) );
  nand_x1_sg U67797 ( .A(n41091), .B(n21741), .X(n21740) );
  nand_x1_sg U67798 ( .A(n40989), .B(n21789), .X(n21786) );
  nand_x1_sg U67799 ( .A(n41091), .B(n21788), .X(n21787) );
  nand_x1_sg U67800 ( .A(n40989), .B(n21836), .X(n21833) );
  nand_x1_sg U67801 ( .A(n41089), .B(n21835), .X(n21834) );
  nand_x1_sg U67802 ( .A(n40991), .B(n21883), .X(n21880) );
  nand_x1_sg U67803 ( .A(n41090), .B(n21882), .X(n21881) );
  nand_x1_sg U67804 ( .A(n40989), .B(n21929), .X(n21926) );
  nand_x1_sg U67805 ( .A(n41089), .B(n21928), .X(n21927) );
  nand_x1_sg U67806 ( .A(n38918), .B(n21976), .X(n21973) );
  nand_x1_sg U67807 ( .A(n38917), .B(n22022), .X(n22019) );
  nand_x1_sg U67808 ( .A(n40991), .B(n22069), .X(n22066) );
  nand_x1_sg U67809 ( .A(n38907), .B(n22115), .X(n22112) );
  nand_x1_sg U67810 ( .A(n40990), .B(n22163), .X(n22160) );
  nand_x1_sg U67811 ( .A(n38907), .B(n22210), .X(n22207) );
  nand_x1_sg U67812 ( .A(n38907), .B(n22258), .X(n22255) );
  nand_x1_sg U67813 ( .A(n40989), .B(n22305), .X(n22302) );
  nand_x1_sg U67814 ( .A(n38907), .B(n22353), .X(n22350) );
  nand_x1_sg U67815 ( .A(n40990), .B(n22400), .X(n22397) );
  nand_x1_sg U67816 ( .A(n38918), .B(n22447), .X(n22444) );
  nand_x1_sg U67817 ( .A(n38917), .B(n22493), .X(n22490) );
  nand_x1_sg U67818 ( .A(n40991), .B(n45015), .X(n22533) );
  nand_x1_sg U67819 ( .A(n19118), .B(n45006), .X(n22534) );
  nand_x1_sg U67820 ( .A(n22978), .B(n40507), .X(n22981) );
  nand_x1_sg U67821 ( .A(n23535), .B(n40500), .X(n23538) );
  nand_x1_sg U67822 ( .A(n23814), .B(n41176), .X(n23817) );
  nand_x1_sg U67823 ( .A(n24093), .B(n39229), .X(n24096) );
  nand_x1_sg U67824 ( .A(n24372), .B(n41166), .X(n24375) );
  nand_x1_sg U67825 ( .A(n24651), .B(n41161), .X(n24654) );
  nand_x1_sg U67826 ( .A(n24929), .B(n41156), .X(n24932) );
  nand_x1_sg U67827 ( .A(n25208), .B(n41151), .X(n25211) );
  nand_x1_sg U67828 ( .A(n25487), .B(n40471), .X(n25490) );
  nand_x1_sg U67829 ( .A(n25766), .B(n40469), .X(n25769) );
  nand_x1_sg U67830 ( .A(n26322), .B(n40464), .X(n26326) );
  nand_x1_sg U67831 ( .A(n26603), .B(n40460), .X(n26606) );
  nor_x1_sg U67832 ( .A(n26233), .B(n41130), .X(\L1_0/n3367 ) );
  nor_x1_sg U67833 ( .A(n26241), .B(n41128), .X(\L1_0/n3363 ) );
  nor_x1_sg U67834 ( .A(n26257), .B(n39249), .X(\L1_0/n3355 ) );
  nor_x1_sg U67835 ( .A(n26273), .B(n41129), .X(\L1_0/n3347 ) );
  nor_x1_sg U67836 ( .A(n26289), .B(n39248), .X(\L1_0/n3339 ) );
  nor_x1_sg U67837 ( .A(n22854), .B(n39143), .X(\L1_0/n4355 ) );
  nor_x1_sg U67838 ( .A(n41929), .B(n41468), .X(n22854) );
  nor_x1_sg U67839 ( .A(n23690), .B(n39460), .X(\L1_0/n4115 ) );
  nor_x1_sg U67840 ( .A(n39975), .B(n39282), .X(n23690) );
  nor_x1_sg U67841 ( .A(n24527), .B(n39463), .X(\L1_0/n3875 ) );
  nor_x1_sg U67842 ( .A(n39987), .B(n40015), .X(n24527) );
  nor_x1_sg U67843 ( .A(n25363), .B(n41373), .X(\L1_0/n3635 ) );
  nor_x1_sg U67844 ( .A(n39999), .B(n40455), .X(n25363) );
  nor_x1_sg U67845 ( .A(n26181), .B(n41130), .X(\L1_0/n3395 ) );
  nor_x1_sg U67846 ( .A(n40999), .B(n39154), .X(n26181) );
  nor_x1_sg U67847 ( .A(n23131), .B(n39902), .X(\L1_0/n4275 ) );
  nor_x1_sg U67848 ( .A(n41928), .B(n41407), .X(n23131) );
  nor_x1_sg U67849 ( .A(n23411), .B(n38960), .X(\L1_0/n4195 ) );
  nor_x1_sg U67850 ( .A(n40695), .B(n39283), .X(n23411) );
  nor_x1_sg U67851 ( .A(n23969), .B(n39448), .X(\L1_0/n4035 ) );
  nor_x1_sg U67852 ( .A(n41939), .B(n39151), .X(n23969) );
  nor_x1_sg U67853 ( .A(n24248), .B(n38966), .X(\L1_0/n3955 ) );
  nor_x1_sg U67854 ( .A(n39983), .B(n40371), .X(n24248) );
  nor_x1_sg U67855 ( .A(n24805), .B(n41331), .X(\L1_0/n3795 ) );
  nor_x1_sg U67856 ( .A(n39991), .B(n41467), .X(n24805) );
  nor_x1_sg U67857 ( .A(n25084), .B(n39923), .X(\L1_0/n3715 ) );
  nor_x1_sg U67858 ( .A(n39997), .B(n41407), .X(n25084) );
  nor_x1_sg U67859 ( .A(n25642), .B(n40034), .X(\L1_0/n3555 ) );
  nor_x1_sg U67860 ( .A(n41919), .B(n41403), .X(n25642) );
  nor_x1_sg U67861 ( .A(n26479), .B(n39454), .X(\L1_0/n3315 ) );
  nor_x1_sg U67862 ( .A(n40007), .B(n39654), .X(n26479) );
  nand_x1_sg U67863 ( .A(n40906), .B(n17468), .X(\L2_0/n2491 ) );
  nand_x1_sg U67864 ( .A(n38910), .B(n41119), .X(n17468) );
  nand_x1_sg U67865 ( .A(n40908), .B(n17471), .X(\L2_0/n2483 ) );
  nand_x1_sg U67866 ( .A(n41119), .B(n17472), .X(n17471) );
  nand_x1_sg U67867 ( .A(n40998), .B(n40067), .X(n17472) );
  nand_x1_sg U67868 ( .A(n40907), .B(n17475), .X(\L2_0/n2479 ) );
  nand_x1_sg U67869 ( .A(n42328), .B(n17474), .X(n17475) );
  nand_x1_sg U67870 ( .A(n40913), .B(n6824), .X(\L2_0/n3531 ) );
  nand_x1_sg U67871 ( .A(n38913), .B(n41390), .X(n6824) );
  nand_x1_sg U67872 ( .A(n38889), .B(n6829), .X(\L2_0/n3519 ) );
  nand_x1_sg U67873 ( .A(n6828), .B(n41390), .X(n6829) );
  inv_x1_sg U67874 ( .A(n20108), .X(n46349) );
  inv_x1_sg U67875 ( .A(n6175), .X(n46386) );
  inv_x1_sg U67876 ( .A(n6034), .X(n46523) );
  nor_x1_sg U67877 ( .A(n5928), .B(n41208), .X(n5104) );
  nand_x1_sg U67878 ( .A(n51200), .B(n51160), .X(n5930) );
  nand_x1_sg U67879 ( .A(n5932), .B(n51179), .X(n5929) );
  nor_x1_sg U67880 ( .A(n40843), .B(n8464), .X(\L2_0/n3360 ) );
  nor_x1_sg U67881 ( .A(n26330), .B(n41127), .X(\L1_0/n3319 ) );
  nor_x1_sg U67882 ( .A(n26329), .B(n26327), .X(n26330) );
  nand_x1_sg U67883 ( .A(n39092), .B(n5858), .X(n5114) );
  nand_x1_sg U67884 ( .A(n41058), .B(n39127), .X(n5858) );
  nand_x1_sg U67885 ( .A(n39093), .B(n5859), .X(n5113) );
  nand_x1_sg U67886 ( .A(n5860), .B(n41281), .X(n5859) );
  nand_x1_sg U67887 ( .A(n5861), .B(n39659), .X(n5860) );
  nand_x1_sg U67888 ( .A(n41214), .B(n22555), .X(\L1_0/n4439 ) );
  nor_x1_sg U67889 ( .A(n5934), .B(n51508), .X(n22557) );
  nor_x1_sg U67890 ( .A(n5931), .B(n22579), .X(n22556) );
  nor_x1_sg U67891 ( .A(n23255), .B(n23256), .X(n23254) );
  nand_x1_sg U67892 ( .A(n41187), .B(n23257), .X(n23256) );
  nand_x1_sg U67893 ( .A(n38881), .B(n8458), .X(\L2_0/n3371 ) );
  nand_x1_sg U67894 ( .A(n39968), .B(n41238), .X(n8458) );
  nand_x1_sg U67895 ( .A(n40892), .B(n8462), .X(\L2_0/n3363 ) );
  nand_x1_sg U67896 ( .A(n8463), .B(n41237), .X(n8462) );
  nand_x1_sg U67897 ( .A(n39969), .B(n40360), .X(n8463) );
  nand_x1_sg U67898 ( .A(n38881), .B(n8465), .X(\L2_0/n3359 ) );
  nand_x1_sg U67899 ( .A(n41237), .B(n8464), .X(n8465) );
  nand_x1_sg U67900 ( .A(n40893), .B(n8471), .X(\L2_0/n3355 ) );
  nand_x1_sg U67901 ( .A(n8470), .B(n41237), .X(n8471) );
  nand_x1_sg U67902 ( .A(n38881), .B(n8478), .X(\L2_0/n3351 ) );
  nand_x1_sg U67903 ( .A(n41236), .B(n8477), .X(n8478) );
  nand_x1_sg U67904 ( .A(n40892), .B(n8485), .X(\L2_0/n3347 ) );
  nand_x1_sg U67905 ( .A(n8484), .B(n41238), .X(n8485) );
  nand_x1_sg U67906 ( .A(n40893), .B(n8491), .X(\L2_0/n3343 ) );
  nand_x1_sg U67907 ( .A(n8490), .B(n41239), .X(n8491) );
  nand_x1_sg U67908 ( .A(n40891), .B(n8497), .X(\L2_0/n3339 ) );
  nand_x1_sg U67909 ( .A(n8496), .B(n41239), .X(n8497) );
  nand_x1_sg U67910 ( .A(n40891), .B(n8503), .X(\L2_0/n3335 ) );
  nand_x1_sg U67911 ( .A(n8502), .B(n41236), .X(n8503) );
  nand_x1_sg U67912 ( .A(n40894), .B(n8509), .X(\L2_0/n3331 ) );
  nand_x1_sg U67913 ( .A(n8508), .B(n41239), .X(n8509) );
  nand_x1_sg U67914 ( .A(n40894), .B(n8515), .X(\L2_0/n3327 ) );
  nand_x1_sg U67915 ( .A(n8514), .B(n41236), .X(n8515) );
  nand_x1_sg U67916 ( .A(n40894), .B(n8521), .X(\L2_0/n3323 ) );
  nand_x1_sg U67917 ( .A(n8520), .B(n39107), .X(n8521) );
  nand_x1_sg U67918 ( .A(n40894), .B(n8527), .X(\L2_0/n3319 ) );
  nand_x1_sg U67919 ( .A(n8526), .B(n41238), .X(n8527) );
  nand_x1_sg U67920 ( .A(n40892), .B(n8533), .X(\L2_0/n3315 ) );
  nand_x1_sg U67921 ( .A(n8532), .B(n41238), .X(n8533) );
  nand_x1_sg U67922 ( .A(n40892), .B(n8539), .X(\L2_0/n3311 ) );
  nand_x1_sg U67923 ( .A(n8538), .B(n41239), .X(n8539) );
  nand_x1_sg U67924 ( .A(n40893), .B(n8545), .X(\L2_0/n3307 ) );
  nand_x1_sg U67925 ( .A(n8544), .B(n41237), .X(n8545) );
  nand_x1_sg U67926 ( .A(n40891), .B(n8551), .X(\L2_0/n3303 ) );
  nand_x1_sg U67927 ( .A(n8550), .B(n39108), .X(n8551) );
  nand_x1_sg U67928 ( .A(n40891), .B(n8557), .X(\L2_0/n3299 ) );
  nand_x1_sg U67929 ( .A(n8556), .B(n39108), .X(n8557) );
  nand_x1_sg U67930 ( .A(n40893), .B(n8563), .X(\L2_0/n3295 ) );
  nand_x1_sg U67931 ( .A(n8562), .B(n39107), .X(n8563) );
  nand_x1_sg U67932 ( .A(n38879), .B(n9278), .X(\L2_0/n3291 ) );
  nand_x1_sg U67933 ( .A(n39972), .B(n41248), .X(n9278) );
  nand_x1_sg U67934 ( .A(n40887), .B(n9282), .X(\L2_0/n3283 ) );
  nand_x1_sg U67935 ( .A(n9283), .B(n41247), .X(n9282) );
  nand_x1_sg U67936 ( .A(n39973), .B(n42103), .X(n9283) );
  nand_x1_sg U67937 ( .A(n38879), .B(n9285), .X(\L2_0/n3279 ) );
  nand_x1_sg U67938 ( .A(n39114), .B(n9284), .X(n9285) );
  nand_x1_sg U67939 ( .A(n40888), .B(n9291), .X(\L2_0/n3275 ) );
  nand_x1_sg U67940 ( .A(n9290), .B(n41246), .X(n9291) );
  nand_x1_sg U67941 ( .A(n38879), .B(n9298), .X(\L2_0/n3271 ) );
  nand_x1_sg U67942 ( .A(n41249), .B(n9297), .X(n9298) );
  nand_x1_sg U67943 ( .A(n40887), .B(n9305), .X(\L2_0/n3267 ) );
  nand_x1_sg U67944 ( .A(n9304), .B(n41249), .X(n9305) );
  nand_x1_sg U67945 ( .A(n40888), .B(n9311), .X(\L2_0/n3263 ) );
  nand_x1_sg U67946 ( .A(n9310), .B(n41249), .X(n9311) );
  nand_x1_sg U67947 ( .A(n40886), .B(n9317), .X(\L2_0/n3259 ) );
  nand_x1_sg U67948 ( .A(n9316), .B(n41247), .X(n9317) );
  nand_x1_sg U67949 ( .A(n40886), .B(n9323), .X(\L2_0/n3255 ) );
  nand_x1_sg U67950 ( .A(n9322), .B(n41247), .X(n9323) );
  nand_x1_sg U67951 ( .A(n40889), .B(n9329), .X(\L2_0/n3251 ) );
  nand_x1_sg U67952 ( .A(n9328), .B(n41246), .X(n9329) );
  nand_x1_sg U67953 ( .A(n40889), .B(n9335), .X(\L2_0/n3247 ) );
  nand_x1_sg U67954 ( .A(n9334), .B(n41247), .X(n9335) );
  nand_x1_sg U67955 ( .A(n40889), .B(n9341), .X(\L2_0/n3243 ) );
  nand_x1_sg U67956 ( .A(n9340), .B(n41248), .X(n9341) );
  nand_x1_sg U67957 ( .A(n40889), .B(n9347), .X(\L2_0/n3239 ) );
  nand_x1_sg U67958 ( .A(n9346), .B(n39113), .X(n9347) );
  nand_x1_sg U67959 ( .A(n40887), .B(n9353), .X(\L2_0/n3235 ) );
  nand_x1_sg U67960 ( .A(n9352), .B(n39114), .X(n9353) );
  nand_x1_sg U67961 ( .A(n40887), .B(n9359), .X(\L2_0/n3231 ) );
  nand_x1_sg U67962 ( .A(n9358), .B(n39113), .X(n9359) );
  nand_x1_sg U67963 ( .A(n40888), .B(n9365), .X(\L2_0/n3227 ) );
  nand_x1_sg U67964 ( .A(n9364), .B(n41249), .X(n9365) );
  nand_x1_sg U67965 ( .A(n40886), .B(n9371), .X(\L2_0/n3223 ) );
  nand_x1_sg U67966 ( .A(n9370), .B(n41248), .X(n9371) );
  nand_x1_sg U67967 ( .A(n40886), .B(n9377), .X(\L2_0/n3219 ) );
  nand_x1_sg U67968 ( .A(n9376), .B(n41246), .X(n9377) );
  nand_x1_sg U67969 ( .A(n40888), .B(n9383), .X(\L2_0/n3215 ) );
  nand_x1_sg U67970 ( .A(n9382), .B(n41248), .X(n9383) );
  nand_x1_sg U67971 ( .A(n40882), .B(n10097), .X(\L2_0/n3211 ) );
  nand_x1_sg U67972 ( .A(n39977), .B(n41197), .X(n10097) );
  nand_x1_sg U67973 ( .A(n40881), .B(n10101), .X(\L2_0/n3203 ) );
  nand_x1_sg U67974 ( .A(n10102), .B(n41197), .X(n10101) );
  nand_x1_sg U67975 ( .A(n39976), .B(n42102), .X(n10102) );
  nand_x1_sg U67976 ( .A(n38877), .B(n10104), .X(\L2_0/n3199 ) );
  nand_x1_sg U67977 ( .A(n39219), .B(n10103), .X(n10104) );
  nand_x1_sg U67978 ( .A(n38877), .B(n10110), .X(\L2_0/n3195 ) );
  nand_x1_sg U67979 ( .A(n10109), .B(n41198), .X(n10110) );
  nand_x1_sg U67980 ( .A(n40883), .B(n10117), .X(\L2_0/n3191 ) );
  nand_x1_sg U67981 ( .A(n41200), .B(n10116), .X(n10117) );
  nand_x1_sg U67982 ( .A(n40883), .B(n10124), .X(\L2_0/n3187 ) );
  nand_x1_sg U67983 ( .A(n10123), .B(n39220), .X(n10124) );
  nand_x1_sg U67984 ( .A(n38877), .B(n10130), .X(\L2_0/n3183 ) );
  nand_x1_sg U67985 ( .A(n10129), .B(n41200), .X(n10130) );
  nand_x1_sg U67986 ( .A(n40882), .B(n10136), .X(\L2_0/n3179 ) );
  nand_x1_sg U67987 ( .A(n10135), .B(n41200), .X(n10136) );
  nand_x1_sg U67988 ( .A(n40883), .B(n10148), .X(\L2_0/n3171 ) );
  nand_x1_sg U67989 ( .A(n10147), .B(n41199), .X(n10148) );
  nand_x1_sg U67990 ( .A(n40881), .B(n10154), .X(\L2_0/n3167 ) );
  nand_x1_sg U67991 ( .A(n10153), .B(n41198), .X(n10154) );
  nand_x1_sg U67992 ( .A(n40881), .B(n10160), .X(\L2_0/n3163 ) );
  nand_x1_sg U67993 ( .A(n10159), .B(n41197), .X(n10160) );
  nand_x1_sg U67994 ( .A(n40884), .B(n10166), .X(\L2_0/n3159 ) );
  nand_x1_sg U67995 ( .A(n10165), .B(n41199), .X(n10166) );
  nand_x1_sg U67996 ( .A(n40882), .B(n10172), .X(\L2_0/n3155 ) );
  nand_x1_sg U67997 ( .A(n10171), .B(n41199), .X(n10172) );
  nand_x1_sg U67998 ( .A(n40884), .B(n10178), .X(\L2_0/n3151 ) );
  nand_x1_sg U67999 ( .A(n10177), .B(n39219), .X(n10178) );
  nand_x1_sg U68000 ( .A(n40882), .B(n10184), .X(\L2_0/n3147 ) );
  nand_x1_sg U68001 ( .A(n10183), .B(n39220), .X(n10184) );
  nand_x1_sg U68002 ( .A(n40883), .B(n10190), .X(\L2_0/n3143 ) );
  nand_x1_sg U68003 ( .A(n10189), .B(n39219), .X(n10190) );
  nand_x1_sg U68004 ( .A(n40884), .B(n10196), .X(\L2_0/n3139 ) );
  nand_x1_sg U68005 ( .A(n10195), .B(n41198), .X(n10196) );
  nand_x1_sg U68006 ( .A(n40884), .B(n10202), .X(\L2_0/n3135 ) );
  nand_x1_sg U68007 ( .A(n10201), .B(n39220), .X(n10202) );
  nand_x1_sg U68008 ( .A(n38875), .B(n10916), .X(\L2_0/n3131 ) );
  nand_x1_sg U68009 ( .A(n39980), .B(n41224), .X(n10916) );
  nand_x1_sg U68010 ( .A(n40877), .B(n10920), .X(\L2_0/n3123 ) );
  nand_x1_sg U68011 ( .A(n10921), .B(n39099), .X(n10920) );
  nand_x1_sg U68012 ( .A(n39981), .B(n42101), .X(n10921) );
  nand_x1_sg U68013 ( .A(n38875), .B(n10923), .X(\L2_0/n3119 ) );
  nand_x1_sg U68014 ( .A(n41224), .B(n10922), .X(n10923) );
  nand_x1_sg U68015 ( .A(n40878), .B(n10929), .X(\L2_0/n3115 ) );
  nand_x1_sg U68016 ( .A(n10928), .B(n41222), .X(n10929) );
  nand_x1_sg U68017 ( .A(n38875), .B(n10936), .X(\L2_0/n3111 ) );
  nand_x1_sg U68018 ( .A(n41223), .B(n10935), .X(n10936) );
  nand_x1_sg U68019 ( .A(n40877), .B(n10943), .X(\L2_0/n3107 ) );
  nand_x1_sg U68020 ( .A(n10942), .B(n39099), .X(n10943) );
  nand_x1_sg U68021 ( .A(n40878), .B(n10949), .X(\L2_0/n3103 ) );
  nand_x1_sg U68022 ( .A(n10948), .B(n41222), .X(n10949) );
  nand_x1_sg U68023 ( .A(n40876), .B(n10955), .X(\L2_0/n3099 ) );
  nand_x1_sg U68024 ( .A(n10954), .B(n41223), .X(n10955) );
  nand_x1_sg U68025 ( .A(n40876), .B(n10961), .X(\L2_0/n3095 ) );
  nand_x1_sg U68026 ( .A(n10960), .B(n39098), .X(n10961) );
  nand_x1_sg U68027 ( .A(n40879), .B(n10967), .X(\L2_0/n3091 ) );
  nand_x1_sg U68028 ( .A(n10966), .B(n39098), .X(n10967) );
  nand_x1_sg U68029 ( .A(n40879), .B(n10973), .X(\L2_0/n3087 ) );
  nand_x1_sg U68030 ( .A(n10972), .B(n41224), .X(n10973) );
  nand_x1_sg U68031 ( .A(n40879), .B(n10979), .X(\L2_0/n3083 ) );
  nand_x1_sg U68032 ( .A(n10978), .B(n39099), .X(n10979) );
  nand_x1_sg U68033 ( .A(n40879), .B(n10985), .X(\L2_0/n3079 ) );
  nand_x1_sg U68034 ( .A(n10984), .B(n41221), .X(n10985) );
  nand_x1_sg U68035 ( .A(n40877), .B(n10991), .X(\L2_0/n3075 ) );
  nand_x1_sg U68036 ( .A(n10990), .B(n41221), .X(n10991) );
  nand_x1_sg U68037 ( .A(n40877), .B(n10997), .X(\L2_0/n3071 ) );
  nand_x1_sg U68038 ( .A(n10996), .B(n41221), .X(n10997) );
  nand_x1_sg U68039 ( .A(n40878), .B(n11003), .X(\L2_0/n3067 ) );
  nand_x1_sg U68040 ( .A(n11002), .B(n39098), .X(n11003) );
  nand_x1_sg U68041 ( .A(n40876), .B(n11009), .X(\L2_0/n3063 ) );
  nand_x1_sg U68042 ( .A(n11008), .B(n41223), .X(n11009) );
  nand_x1_sg U68043 ( .A(n40876), .B(n11015), .X(\L2_0/n3059 ) );
  nand_x1_sg U68044 ( .A(n11014), .B(n41224), .X(n11015) );
  nand_x1_sg U68045 ( .A(n40878), .B(n11021), .X(\L2_0/n3055 ) );
  nand_x1_sg U68046 ( .A(n11020), .B(n41222), .X(n11021) );
  nand_x1_sg U68047 ( .A(n38873), .B(n11735), .X(\L2_0/n3051 ) );
  nand_x1_sg U68048 ( .A(n39985), .B(n41205), .X(n11735) );
  nand_x1_sg U68049 ( .A(n40872), .B(n11739), .X(\L2_0/n3043 ) );
  nand_x1_sg U68050 ( .A(n11740), .B(n39086), .X(n11739) );
  nand_x1_sg U68051 ( .A(n39984), .B(n42100), .X(n11740) );
  nand_x1_sg U68052 ( .A(n38873), .B(n11742), .X(\L2_0/n3039 ) );
  nand_x1_sg U68053 ( .A(n41204), .B(n11741), .X(n11742) );
  nand_x1_sg U68054 ( .A(n40873), .B(n11748), .X(\L2_0/n3035 ) );
  nand_x1_sg U68055 ( .A(n11747), .B(n41203), .X(n11748) );
  nand_x1_sg U68056 ( .A(n38873), .B(n11755), .X(\L2_0/n3031 ) );
  nand_x1_sg U68057 ( .A(n39087), .B(n11754), .X(n11755) );
  nand_x1_sg U68058 ( .A(n40872), .B(n11762), .X(\L2_0/n3027 ) );
  nand_x1_sg U68059 ( .A(n11761), .B(n41202), .X(n11762) );
  nand_x1_sg U68060 ( .A(n40873), .B(n11768), .X(\L2_0/n3023 ) );
  nand_x1_sg U68061 ( .A(n11767), .B(n41205), .X(n11768) );
  nand_x1_sg U68062 ( .A(n40871), .B(n11774), .X(\L2_0/n3019 ) );
  nand_x1_sg U68063 ( .A(n11773), .B(n41202), .X(n11774) );
  nand_x1_sg U68064 ( .A(n40871), .B(n11780), .X(\L2_0/n3015 ) );
  nand_x1_sg U68065 ( .A(n11779), .B(n39086), .X(n11780) );
  nand_x1_sg U68066 ( .A(n40874), .B(n11786), .X(\L2_0/n3011 ) );
  nand_x1_sg U68067 ( .A(n11785), .B(n41203), .X(n11786) );
  nand_x1_sg U68068 ( .A(n40874), .B(n11792), .X(\L2_0/n3007 ) );
  nand_x1_sg U68069 ( .A(n11791), .B(n41205), .X(n11792) );
  nand_x1_sg U68070 ( .A(n40874), .B(n11798), .X(\L2_0/n3003 ) );
  nand_x1_sg U68071 ( .A(n11797), .B(n41204), .X(n11798) );
  nand_x1_sg U68072 ( .A(n40874), .B(n11804), .X(\L2_0/n2999 ) );
  nand_x1_sg U68073 ( .A(n11803), .B(n41202), .X(n11804) );
  nand_x1_sg U68074 ( .A(n40872), .B(n11810), .X(\L2_0/n2995 ) );
  nand_x1_sg U68075 ( .A(n11809), .B(n41205), .X(n11810) );
  nand_x1_sg U68076 ( .A(n40872), .B(n11816), .X(\L2_0/n2991 ) );
  nand_x1_sg U68077 ( .A(n11815), .B(n41204), .X(n11816) );
  nand_x1_sg U68078 ( .A(n40873), .B(n11822), .X(\L2_0/n2987 ) );
  nand_x1_sg U68079 ( .A(n11821), .B(n39086), .X(n11822) );
  nand_x1_sg U68080 ( .A(n40871), .B(n11828), .X(\L2_0/n2983 ) );
  nand_x1_sg U68081 ( .A(n11827), .B(n39087), .X(n11828) );
  nand_x1_sg U68082 ( .A(n40871), .B(n11834), .X(\L2_0/n2979 ) );
  nand_x1_sg U68083 ( .A(n11833), .B(n41204), .X(n11834) );
  nand_x1_sg U68084 ( .A(n40873), .B(n11840), .X(\L2_0/n2975 ) );
  nand_x1_sg U68085 ( .A(n11839), .B(n39087), .X(n11840) );
  nand_x1_sg U68086 ( .A(n40867), .B(n12554), .X(\L2_0/n2971 ) );
  nand_x1_sg U68087 ( .A(n39989), .B(n41259), .X(n12554) );
  nand_x1_sg U68088 ( .A(n40866), .B(n12558), .X(\L2_0/n2963 ) );
  nand_x1_sg U68089 ( .A(n12559), .B(n41258), .X(n12558) );
  nand_x1_sg U68090 ( .A(n39988), .B(n42099), .X(n12559) );
  nand_x1_sg U68091 ( .A(n38871), .B(n12561), .X(\L2_0/n2959 ) );
  nand_x1_sg U68092 ( .A(n41259), .B(n12560), .X(n12561) );
  nand_x1_sg U68093 ( .A(n38871), .B(n12567), .X(\L2_0/n2955 ) );
  nand_x1_sg U68094 ( .A(n12566), .B(n41257), .X(n12567) );
  nand_x1_sg U68095 ( .A(n40868), .B(n12574), .X(\L2_0/n2951 ) );
  nand_x1_sg U68096 ( .A(n41258), .B(n12573), .X(n12574) );
  nand_x1_sg U68097 ( .A(n40868), .B(n12581), .X(\L2_0/n2947 ) );
  nand_x1_sg U68098 ( .A(n12580), .B(n41258), .X(n12581) );
  nand_x1_sg U68099 ( .A(n38871), .B(n12587), .X(\L2_0/n2943 ) );
  nand_x1_sg U68100 ( .A(n12586), .B(n41258), .X(n12587) );
  nand_x1_sg U68101 ( .A(n40867), .B(n12593), .X(\L2_0/n2939 ) );
  nand_x1_sg U68102 ( .A(n12592), .B(n39118), .X(n12593) );
  nand_x1_sg U68103 ( .A(n40868), .B(n12599), .X(\L2_0/n2935 ) );
  nand_x1_sg U68104 ( .A(n12598), .B(n41256), .X(n12599) );
  nand_x1_sg U68105 ( .A(n40866), .B(n12605), .X(\L2_0/n2931 ) );
  nand_x1_sg U68106 ( .A(n12604), .B(n41257), .X(n12605) );
  nand_x1_sg U68107 ( .A(n40866), .B(n12611), .X(\L2_0/n2927 ) );
  nand_x1_sg U68108 ( .A(n12610), .B(n41257), .X(n12611) );
  nand_x1_sg U68109 ( .A(n40869), .B(n12617), .X(\L2_0/n2923 ) );
  nand_x1_sg U68110 ( .A(n12616), .B(n39119), .X(n12617) );
  nand_x1_sg U68111 ( .A(n40867), .B(n12623), .X(\L2_0/n2919 ) );
  nand_x1_sg U68112 ( .A(n12622), .B(n39118), .X(n12623) );
  nand_x1_sg U68113 ( .A(n40869), .B(n12629), .X(\L2_0/n2915 ) );
  nand_x1_sg U68114 ( .A(n12628), .B(n41256), .X(n12629) );
  nand_x1_sg U68115 ( .A(n40867), .B(n12635), .X(\L2_0/n2911 ) );
  nand_x1_sg U68116 ( .A(n12634), .B(n39118), .X(n12635) );
  nand_x1_sg U68117 ( .A(n40868), .B(n12641), .X(\L2_0/n2907 ) );
  nand_x1_sg U68118 ( .A(n12640), .B(n41259), .X(n12641) );
  nand_x1_sg U68119 ( .A(n40869), .B(n12653), .X(\L2_0/n2899 ) );
  nand_x1_sg U68120 ( .A(n12652), .B(n41259), .X(n12653) );
  nand_x1_sg U68121 ( .A(n40869), .B(n12659), .X(\L2_0/n2895 ) );
  nand_x1_sg U68122 ( .A(n12658), .B(n39119), .X(n12659) );
  nand_x1_sg U68123 ( .A(n40862), .B(n13373), .X(\L2_0/n2891 ) );
  nand_x1_sg U68124 ( .A(n39992), .B(n41243), .X(n13373) );
  nand_x1_sg U68125 ( .A(n40861), .B(n13377), .X(\L2_0/n2883 ) );
  nand_x1_sg U68126 ( .A(n13378), .B(n41242), .X(n13377) );
  nand_x1_sg U68127 ( .A(n39993), .B(n42098), .X(n13378) );
  nand_x1_sg U68128 ( .A(n38869), .B(n13380), .X(\L2_0/n2879 ) );
  nand_x1_sg U68129 ( .A(n39111), .B(n13379), .X(n13380) );
  nand_x1_sg U68130 ( .A(n38869), .B(n13386), .X(\L2_0/n2875 ) );
  nand_x1_sg U68131 ( .A(n13385), .B(n39110), .X(n13386) );
  nand_x1_sg U68132 ( .A(n40863), .B(n13393), .X(\L2_0/n2871 ) );
  nand_x1_sg U68133 ( .A(n41244), .B(n13392), .X(n13393) );
  nand_x1_sg U68134 ( .A(n40863), .B(n13400), .X(\L2_0/n2867 ) );
  nand_x1_sg U68135 ( .A(n13399), .B(n41244), .X(n13400) );
  nand_x1_sg U68136 ( .A(n38869), .B(n13406), .X(\L2_0/n2863 ) );
  nand_x1_sg U68137 ( .A(n13405), .B(n41244), .X(n13406) );
  nand_x1_sg U68138 ( .A(n40862), .B(n13412), .X(\L2_0/n2859 ) );
  nand_x1_sg U68139 ( .A(n13411), .B(n41242), .X(n13412) );
  nand_x1_sg U68140 ( .A(n40863), .B(n13418), .X(\L2_0/n2855 ) );
  nand_x1_sg U68141 ( .A(n13417), .B(n39110), .X(n13418) );
  nand_x1_sg U68142 ( .A(n40861), .B(n13424), .X(\L2_0/n2851 ) );
  nand_x1_sg U68143 ( .A(n13423), .B(n41243), .X(n13424) );
  nand_x1_sg U68144 ( .A(n40861), .B(n13430), .X(\L2_0/n2847 ) );
  nand_x1_sg U68145 ( .A(n13429), .B(n39111), .X(n13430) );
  nand_x1_sg U68146 ( .A(n40864), .B(n13436), .X(\L2_0/n2843 ) );
  nand_x1_sg U68147 ( .A(n13435), .B(n41241), .X(n13436) );
  nand_x1_sg U68148 ( .A(n40862), .B(n13442), .X(\L2_0/n2839 ) );
  nand_x1_sg U68149 ( .A(n13441), .B(n41242), .X(n13442) );
  nand_x1_sg U68150 ( .A(n40864), .B(n13448), .X(\L2_0/n2835 ) );
  nand_x1_sg U68151 ( .A(n13447), .B(n41242), .X(n13448) );
  nand_x1_sg U68152 ( .A(n40862), .B(n13454), .X(\L2_0/n2831 ) );
  nand_x1_sg U68153 ( .A(n13453), .B(n39110), .X(n13454) );
  nand_x1_sg U68154 ( .A(n40863), .B(n13460), .X(\L2_0/n2827 ) );
  nand_x1_sg U68155 ( .A(n13459), .B(n39111), .X(n13460) );
  nand_x1_sg U68156 ( .A(n40864), .B(n13472), .X(\L2_0/n2819 ) );
  nand_x1_sg U68157 ( .A(n13471), .B(n41243), .X(n13472) );
  nand_x1_sg U68158 ( .A(n40864), .B(n13478), .X(\L2_0/n2815 ) );
  nand_x1_sg U68159 ( .A(n13477), .B(n41241), .X(n13478) );
  nand_x1_sg U68160 ( .A(n38867), .B(n14192), .X(\L2_0/n2811 ) );
  nand_x1_sg U68161 ( .A(n39997), .B(n39101), .X(n14192) );
  nand_x1_sg U68162 ( .A(n40857), .B(n14196), .X(\L2_0/n2803 ) );
  nand_x1_sg U68163 ( .A(n14197), .B(n41227), .X(n14196) );
  nand_x1_sg U68164 ( .A(n39996), .B(n42097), .X(n14197) );
  nand_x1_sg U68165 ( .A(n38867), .B(n14199), .X(\L2_0/n2799 ) );
  nand_x1_sg U68166 ( .A(n39101), .B(n14198), .X(n14199) );
  nand_x1_sg U68167 ( .A(n40858), .B(n14205), .X(\L2_0/n2795 ) );
  nand_x1_sg U68168 ( .A(n14204), .B(n41226), .X(n14205) );
  nand_x1_sg U68169 ( .A(n38867), .B(n14212), .X(\L2_0/n2791 ) );
  nand_x1_sg U68170 ( .A(n41229), .B(n14211), .X(n14212) );
  nand_x1_sg U68171 ( .A(n40857), .B(n14219), .X(\L2_0/n2787 ) );
  nand_x1_sg U68172 ( .A(n14218), .B(n39102), .X(n14219) );
  nand_x1_sg U68173 ( .A(n40858), .B(n14225), .X(\L2_0/n2783 ) );
  nand_x1_sg U68174 ( .A(n14224), .B(n41228), .X(n14225) );
  nand_x1_sg U68175 ( .A(n40856), .B(n14231), .X(\L2_0/n2779 ) );
  nand_x1_sg U68176 ( .A(n14230), .B(n41227), .X(n14231) );
  nand_x1_sg U68177 ( .A(n40856), .B(n14237), .X(\L2_0/n2775 ) );
  nand_x1_sg U68178 ( .A(n14236), .B(n41226), .X(n14237) );
  nand_x1_sg U68179 ( .A(n40859), .B(n14243), .X(\L2_0/n2771 ) );
  nand_x1_sg U68180 ( .A(n14242), .B(n41228), .X(n14243) );
  nand_x1_sg U68181 ( .A(n40859), .B(n14249), .X(\L2_0/n2767 ) );
  nand_x1_sg U68182 ( .A(n14248), .B(n41229), .X(n14249) );
  nand_x1_sg U68183 ( .A(n40859), .B(n14255), .X(\L2_0/n2763 ) );
  nand_x1_sg U68184 ( .A(n14254), .B(n41229), .X(n14255) );
  nand_x1_sg U68185 ( .A(n40859), .B(n14261), .X(\L2_0/n2759 ) );
  nand_x1_sg U68186 ( .A(n14260), .B(n41227), .X(n14261) );
  nand_x1_sg U68187 ( .A(n40857), .B(n14267), .X(\L2_0/n2755 ) );
  nand_x1_sg U68188 ( .A(n14266), .B(n39102), .X(n14267) );
  nand_x1_sg U68189 ( .A(n40857), .B(n14273), .X(\L2_0/n2751 ) );
  nand_x1_sg U68190 ( .A(n14272), .B(n39101), .X(n14273) );
  nand_x1_sg U68191 ( .A(n40858), .B(n14279), .X(\L2_0/n2747 ) );
  nand_x1_sg U68192 ( .A(n14278), .B(n41229), .X(n14279) );
  nand_x1_sg U68193 ( .A(n40856), .B(n14285), .X(\L2_0/n2743 ) );
  nand_x1_sg U68194 ( .A(n14284), .B(n41226), .X(n14285) );
  nand_x1_sg U68195 ( .A(n40856), .B(n14291), .X(\L2_0/n2739 ) );
  nand_x1_sg U68196 ( .A(n14290), .B(n39102), .X(n14291) );
  nand_x1_sg U68197 ( .A(n40858), .B(n14297), .X(\L2_0/n2735 ) );
  nand_x1_sg U68198 ( .A(n14296), .B(n41228), .X(n14297) );
  nand_x1_sg U68199 ( .A(n38865), .B(n15011), .X(\L2_0/n2731 ) );
  nand_x1_sg U68200 ( .A(n40001), .B(n41234), .X(n15011) );
  nand_x1_sg U68201 ( .A(n40852), .B(n15015), .X(\L2_0/n2723 ) );
  nand_x1_sg U68202 ( .A(n15016), .B(n41234), .X(n15015) );
  nand_x1_sg U68203 ( .A(n40000), .B(n40320), .X(n15016) );
  nand_x1_sg U68204 ( .A(n38865), .B(n15018), .X(\L2_0/n2719 ) );
  nand_x1_sg U68205 ( .A(n39105), .B(n15017), .X(n15018) );
  nand_x1_sg U68206 ( .A(n40853), .B(n15024), .X(\L2_0/n2715 ) );
  nand_x1_sg U68207 ( .A(n15023), .B(n41232), .X(n15024) );
  nand_x1_sg U68208 ( .A(n38865), .B(n15031), .X(\L2_0/n2711 ) );
  nand_x1_sg U68209 ( .A(n39105), .B(n15030), .X(n15031) );
  nand_x1_sg U68210 ( .A(n40852), .B(n15038), .X(\L2_0/n2707 ) );
  nand_x1_sg U68211 ( .A(n15037), .B(n41233), .X(n15038) );
  nand_x1_sg U68212 ( .A(n40853), .B(n15044), .X(\L2_0/n2703 ) );
  nand_x1_sg U68213 ( .A(n15043), .B(n41231), .X(n15044) );
  nand_x1_sg U68214 ( .A(n40851), .B(n15050), .X(\L2_0/n2699 ) );
  nand_x1_sg U68215 ( .A(n15049), .B(n39104), .X(n15050) );
  nand_x1_sg U68216 ( .A(n40851), .B(n15056), .X(\L2_0/n2695 ) );
  nand_x1_sg U68217 ( .A(n15055), .B(n41233), .X(n15056) );
  nand_x1_sg U68218 ( .A(n40854), .B(n15062), .X(\L2_0/n2691 ) );
  nand_x1_sg U68219 ( .A(n15061), .B(n41233), .X(n15062) );
  nand_x1_sg U68220 ( .A(n40854), .B(n15068), .X(\L2_0/n2687 ) );
  nand_x1_sg U68221 ( .A(n15067), .B(n41232), .X(n15068) );
  nand_x1_sg U68222 ( .A(n40854), .B(n15074), .X(\L2_0/n2683 ) );
  nand_x1_sg U68223 ( .A(n15073), .B(n41231), .X(n15074) );
  nand_x1_sg U68224 ( .A(n40854), .B(n15080), .X(\L2_0/n2679 ) );
  nand_x1_sg U68225 ( .A(n15079), .B(n41232), .X(n15080) );
  nand_x1_sg U68226 ( .A(n40852), .B(n15086), .X(\L2_0/n2675 ) );
  nand_x1_sg U68227 ( .A(n15085), .B(n39104), .X(n15086) );
  nand_x1_sg U68228 ( .A(n40852), .B(n15092), .X(\L2_0/n2671 ) );
  nand_x1_sg U68229 ( .A(n15091), .B(n41233), .X(n15092) );
  nand_x1_sg U68230 ( .A(n40853), .B(n15098), .X(\L2_0/n2667 ) );
  nand_x1_sg U68231 ( .A(n15097), .B(n41234), .X(n15098) );
  nand_x1_sg U68232 ( .A(n40851), .B(n15104), .X(\L2_0/n2663 ) );
  nand_x1_sg U68233 ( .A(n15103), .B(n41231), .X(n15104) );
  nand_x1_sg U68234 ( .A(n40851), .B(n15110), .X(\L2_0/n2659 ) );
  nand_x1_sg U68235 ( .A(n15109), .B(n39105), .X(n15110) );
  nand_x1_sg U68236 ( .A(n40853), .B(n15116), .X(\L2_0/n2655 ) );
  nand_x1_sg U68237 ( .A(n15115), .B(n39104), .X(n15116) );
  nand_x1_sg U68238 ( .A(n38883), .B(n15830), .X(\L2_0/n2651 ) );
  nand_x1_sg U68239 ( .A(n40005), .B(n39132), .X(n15830) );
  nand_x1_sg U68240 ( .A(n40897), .B(n15834), .X(\L2_0/n2643 ) );
  nand_x1_sg U68241 ( .A(n15835), .B(n41293), .X(n15834) );
  nand_x1_sg U68242 ( .A(n40004), .B(n42094), .X(n15835) );
  nand_x1_sg U68243 ( .A(n38883), .B(n15837), .X(\L2_0/n2639 ) );
  nand_x1_sg U68244 ( .A(n41290), .B(n15836), .X(n15837) );
  nand_x1_sg U68245 ( .A(n40898), .B(n15843), .X(\L2_0/n2635 ) );
  nand_x1_sg U68246 ( .A(n15842), .B(n39132), .X(n15843) );
  nand_x1_sg U68247 ( .A(n38883), .B(n15850), .X(\L2_0/n2631 ) );
  nand_x1_sg U68248 ( .A(n41291), .B(n15849), .X(n15850) );
  nand_x1_sg U68249 ( .A(n40897), .B(n15857), .X(\L2_0/n2627 ) );
  nand_x1_sg U68250 ( .A(n15856), .B(n41291), .X(n15857) );
  nand_x1_sg U68251 ( .A(n40898), .B(n15863), .X(\L2_0/n2623 ) );
  nand_x1_sg U68252 ( .A(n15862), .B(n41291), .X(n15863) );
  nand_x1_sg U68253 ( .A(n40896), .B(n15869), .X(\L2_0/n2619 ) );
  nand_x1_sg U68254 ( .A(n15868), .B(n41293), .X(n15869) );
  nand_x1_sg U68255 ( .A(n40896), .B(n15875), .X(\L2_0/n2615 ) );
  nand_x1_sg U68256 ( .A(n15874), .B(n41290), .X(n15875) );
  nand_x1_sg U68257 ( .A(n40899), .B(n15881), .X(\L2_0/n2611 ) );
  nand_x1_sg U68258 ( .A(n15880), .B(n41292), .X(n15881) );
  nand_x1_sg U68259 ( .A(n40899), .B(n15887), .X(\L2_0/n2607 ) );
  nand_x1_sg U68260 ( .A(n15886), .B(n41293), .X(n15887) );
  nand_x1_sg U68261 ( .A(n40899), .B(n15893), .X(\L2_0/n2603 ) );
  nand_x1_sg U68262 ( .A(n15892), .B(n39133), .X(n15893) );
  nand_x1_sg U68263 ( .A(n40899), .B(n15899), .X(\L2_0/n2599 ) );
  nand_x1_sg U68264 ( .A(n15898), .B(n39132), .X(n15899) );
  nand_x1_sg U68265 ( .A(n40897), .B(n15905), .X(\L2_0/n2595 ) );
  nand_x1_sg U68266 ( .A(n15904), .B(n41290), .X(n15905) );
  nand_x1_sg U68267 ( .A(n40897), .B(n15911), .X(\L2_0/n2591 ) );
  nand_x1_sg U68268 ( .A(n15910), .B(n41292), .X(n15911) );
  nand_x1_sg U68269 ( .A(n40898), .B(n15917), .X(\L2_0/n2587 ) );
  nand_x1_sg U68270 ( .A(n15916), .B(n41293), .X(n15917) );
  nand_x1_sg U68271 ( .A(n40896), .B(n15923), .X(\L2_0/n2583 ) );
  nand_x1_sg U68272 ( .A(n15922), .B(n39133), .X(n15923) );
  nand_x1_sg U68273 ( .A(n40896), .B(n15929), .X(\L2_0/n2579 ) );
  nand_x1_sg U68274 ( .A(n15928), .B(n41290), .X(n15929) );
  nand_x1_sg U68275 ( .A(n40898), .B(n15935), .X(\L2_0/n2575 ) );
  nand_x1_sg U68276 ( .A(n15934), .B(n41292), .X(n15935) );
  nand_x1_sg U68277 ( .A(n40904), .B(n16648), .X(\L2_0/n2571 ) );
  nand_x1_sg U68278 ( .A(n38908), .B(n41216), .X(n16648) );
  nand_x1_sg U68279 ( .A(n40901), .B(n16653), .X(\L2_0/n2559 ) );
  nand_x1_sg U68280 ( .A(n39095), .B(n16652), .X(n16653) );
  nand_x1_sg U68281 ( .A(n40881), .B(n10142), .X(\L2_0/n3175 ) );
  nand_x1_sg U68282 ( .A(n10141), .B(n41199), .X(n10142) );
  nand_x1_sg U68283 ( .A(n40866), .B(n12647), .X(\L2_0/n2903 ) );
  nand_x1_sg U68284 ( .A(n12646), .B(n41256), .X(n12647) );
  nand_x1_sg U68285 ( .A(n40861), .B(n13466), .X(\L2_0/n2823 ) );
  nand_x1_sg U68286 ( .A(n13465), .B(n41244), .X(n13466) );
  nand_x1_sg U68287 ( .A(n38863), .B(n18289), .X(\L2_0/n2411 ) );
  nand_x1_sg U68288 ( .A(n40009), .B(n41264), .X(n18289) );
  nand_x1_sg U68289 ( .A(n40847), .B(n18293), .X(\L2_0/n2403 ) );
  nand_x1_sg U68290 ( .A(n18294), .B(n41262), .X(n18293) );
  nand_x1_sg U68291 ( .A(n40008), .B(n42093), .X(n18294) );
  nand_x1_sg U68292 ( .A(n38863), .B(n18296), .X(\L2_0/n2399 ) );
  nand_x1_sg U68293 ( .A(n41262), .B(n18295), .X(n18296) );
  nand_x1_sg U68294 ( .A(n40848), .B(n18302), .X(\L2_0/n2395 ) );
  nand_x1_sg U68295 ( .A(n18301), .B(n41263), .X(n18302) );
  nand_x1_sg U68296 ( .A(n38863), .B(n18309), .X(\L2_0/n2391 ) );
  nand_x1_sg U68297 ( .A(n41264), .B(n18308), .X(n18309) );
  nand_x1_sg U68298 ( .A(n40847), .B(n18316), .X(\L2_0/n2387 ) );
  nand_x1_sg U68299 ( .A(n18315), .B(n39121), .X(n18316) );
  nand_x1_sg U68300 ( .A(n40848), .B(n18322), .X(\L2_0/n2383 ) );
  nand_x1_sg U68301 ( .A(n18321), .B(n39121), .X(n18322) );
  nand_x1_sg U68302 ( .A(n40849), .B(n18328), .X(\L2_0/n2379 ) );
  nand_x1_sg U68303 ( .A(n18327), .B(n41262), .X(n18328) );
  nand_x1_sg U68304 ( .A(n40846), .B(n18334), .X(\L2_0/n2375 ) );
  nand_x1_sg U68305 ( .A(n18333), .B(n41261), .X(n18334) );
  nand_x1_sg U68306 ( .A(n40846), .B(n18340), .X(\L2_0/n2371 ) );
  nand_x1_sg U68307 ( .A(n18339), .B(n39122), .X(n18340) );
  nand_x1_sg U68308 ( .A(n40849), .B(n18346), .X(\L2_0/n2367 ) );
  nand_x1_sg U68309 ( .A(n18345), .B(n41264), .X(n18346) );
  nand_x1_sg U68310 ( .A(n40849), .B(n18352), .X(\L2_0/n2363 ) );
  nand_x1_sg U68311 ( .A(n18351), .B(n39121), .X(n18352) );
  nand_x1_sg U68312 ( .A(n40848), .B(n18358), .X(\L2_0/n2359 ) );
  nand_x1_sg U68313 ( .A(n18357), .B(n41264), .X(n18358) );
  nand_x1_sg U68314 ( .A(n40849), .B(n18364), .X(\L2_0/n2355 ) );
  nand_x1_sg U68315 ( .A(n18363), .B(n41263), .X(n18364) );
  nand_x1_sg U68316 ( .A(n40847), .B(n18370), .X(\L2_0/n2351 ) );
  nand_x1_sg U68317 ( .A(n18369), .B(n39122), .X(n18370) );
  nand_x1_sg U68318 ( .A(n40848), .B(n18376), .X(\L2_0/n2347 ) );
  nand_x1_sg U68319 ( .A(n18375), .B(n39122), .X(n18376) );
  nand_x1_sg U68320 ( .A(n40847), .B(n18382), .X(\L2_0/n2343 ) );
  nand_x1_sg U68321 ( .A(n18381), .B(n41262), .X(n18382) );
  nand_x1_sg U68322 ( .A(n40846), .B(n18388), .X(\L2_0/n2339 ) );
  nand_x1_sg U68323 ( .A(n18387), .B(n41263), .X(n18388) );
  nand_x1_sg U68324 ( .A(n40846), .B(n18394), .X(\L2_0/n2335 ) );
  nand_x1_sg U68325 ( .A(n18393), .B(n41263), .X(n18394) );
  inv_x1_sg U68326 ( .A(n23066), .X(n47197) );
  inv_x1_sg U68327 ( .A(n23346), .X(n47482) );
  inv_x1_sg U68328 ( .A(n23625), .X(n47767) );
  inv_x1_sg U68329 ( .A(n23904), .X(n48052) );
  inv_x1_sg U68330 ( .A(n24183), .X(n48337) );
  inv_x1_sg U68331 ( .A(n24462), .X(n48622) );
  inv_x1_sg U68332 ( .A(n24740), .X(n48908) );
  inv_x1_sg U68333 ( .A(n25019), .X(n49195) );
  inv_x1_sg U68334 ( .A(n25298), .X(n49481) );
  inv_x1_sg U68335 ( .A(n25577), .X(n49767) );
  inv_x1_sg U68336 ( .A(n25854), .X(n50053) );
  inv_x1_sg U68337 ( .A(n26083), .X(n50338) );
  inv_x1_sg U68338 ( .A(n26414), .X(n50627) );
  inv_x1_sg U68339 ( .A(n26692), .X(n50914) );
  inv_x1_sg U68340 ( .A(n22789), .X(n46904) );
  inv_x1_sg U68341 ( .A(n5931), .X(n51200) );
  nand_x1_sg U68342 ( .A(n5861), .B(n22706), .X(n22705) );
  nor_x1_sg U68343 ( .A(n41209), .B(n22638), .X(n22706) );
  nand_x1_sg U68344 ( .A(n41283), .B(n5913), .X(n5912) );
  nand_x1_sg U68345 ( .A(n41282), .B(n5773), .X(n5772) );
  nand_x1_sg U68346 ( .A(n41280), .B(n5786), .X(n22632) );
  nand_x1_sg U68347 ( .A(n41280), .B(n5874), .X(n5873) );
  nand_x1_sg U68348 ( .A(n41282), .B(n5829), .X(n5828) );
  nand_x1_sg U68349 ( .A(n39126), .B(n5777), .X(n5776) );
  nand_x1_sg U68350 ( .A(n39127), .B(n5863), .X(n5862) );
  nand_x1_sg U68351 ( .A(n41281), .B(n5833), .X(n5832) );
  nand_x1_sg U68352 ( .A(n41280), .B(n5771), .X(n5769) );
  nand_x1_sg U68353 ( .A(n39127), .B(n5788), .X(n5787) );
  nand_x1_sg U68354 ( .A(n39126), .B(n5842), .X(n5841) );
  nand_x1_sg U68355 ( .A(n39126), .B(n5827), .X(n5826) );
  nand_x1_sg U68356 ( .A(n41283), .B(n5775), .X(n5774) );
  nand_x1_sg U68357 ( .A(n41282), .B(n5883), .X(n5882) );
  nand_x1_sg U68358 ( .A(n41281), .B(n5950), .X(n5949) );
  nand_x1_sg U68359 ( .A(n41281), .B(n5831), .X(n5830) );
  nor_x1_sg U68360 ( .A(n36904), .B(n36905), .X(n1998) );
  nor_x1_sg U68361 ( .A(n36906), .B(n41522), .X(n36905) );
  nor_x1_sg U68362 ( .A(n39727), .B(n51530), .X(n36906) );
  nor_x1_sg U68363 ( .A(n36902), .B(n39728), .X(n42387) );
  inv_x1_sg U68364 ( .A(n36902), .X(n51529) );
  nor_x1_sg U68365 ( .A(n22796), .B(n22792), .X(n22794) );
  nand_x1_sg U68366 ( .A(n22792), .B(n22796), .X(n22795) );
  nor_x1_sg U68367 ( .A(n26090), .B(n26089), .X(n26087) );
  nand_x1_sg U68368 ( .A(n26089), .B(n26090), .X(n26088) );
  nor_x1_sg U68369 ( .A(n41632), .B(n42021), .X(n18286) );
  nor_x1_sg U68370 ( .A(n22710), .B(n22709), .X(n22707) );
  nand_x1_sg U68371 ( .A(n22709), .B(n22710), .X(n22708) );
  nand_x1_sg U68372 ( .A(n41299), .B(n38816), .X(n23262) );
  nand_x1_sg U68373 ( .A(n26767), .B(n18286), .X(n5987) );
  nor_x1_sg U68374 ( .A(n6210), .B(n20282), .X(n20281) );
  nand_x1_sg U68375 ( .A(n20282), .B(n38632), .X(n20283) );
  nor_x1_sg U68376 ( .A(n6102), .B(n20129), .X(n20128) );
  nand_x1_sg U68377 ( .A(n20129), .B(n6102), .X(n20130) );
  nor_x1_sg U68378 ( .A(n6023), .B(n19929), .X(n19928) );
  nand_x1_sg U68379 ( .A(n19929), .B(n38626), .X(n19930) );
  nor_x1_sg U68380 ( .A(n42333), .B(n19307), .X(n19306) );
  nand_x1_sg U68381 ( .A(n19307), .B(n38675), .X(n19308) );
  nor_x1_sg U68382 ( .A(n51136), .B(n42162), .X(n17465) );
  nor_x1_sg U68383 ( .A(n46555), .B(n19746), .X(n19743) );
  nor_x1_sg U68384 ( .A(n41539), .B(n19745), .X(n19744) );
  inv_x1_sg U68385 ( .A(n19745), .X(n46555) );
  nor_x1_sg U68386 ( .A(n46398), .B(n20113), .X(n20110) );
  nor_x1_sg U68387 ( .A(n41970), .B(n20112), .X(n20111) );
  inv_x1_sg U68388 ( .A(n20112), .X(n46398) );
  nor_x1_sg U68389 ( .A(n46485), .B(n19719), .X(n19716) );
  nor_x1_sg U68390 ( .A(n41953), .B(n19718), .X(n19717) );
  inv_x1_sg U68391 ( .A(n19718), .X(n46485) );
  nor_x1_sg U68392 ( .A(n38624), .B(n19735), .X(n19734) );
  nand_x1_sg U68393 ( .A(n19735), .B(n5969), .X(n19736) );
  nor_x1_sg U68394 ( .A(n38629), .B(n19732), .X(n19731) );
  nand_x1_sg U68395 ( .A(n19732), .B(n5964), .X(n19733) );
  nor_x1_sg U68396 ( .A(n42342), .B(n19330), .X(n19329) );
  nand_x1_sg U68397 ( .A(n19330), .B(n38718), .X(n19331) );
  nor_x1_sg U68398 ( .A(n38630), .B(n19741), .X(n19740) );
  nand_x1_sg U68399 ( .A(n19741), .B(n6003), .X(n19742) );
  nor_x1_sg U68400 ( .A(n42341), .B(n19318), .X(n19317) );
  nand_x1_sg U68401 ( .A(n19318), .B(n38716), .X(n19319) );
  nor_x1_sg U68402 ( .A(n38671), .B(n19738), .X(n19737) );
  nand_x1_sg U68403 ( .A(n19738), .B(n5968), .X(n19739) );
  inv_x1_sg U68404 ( .A(n25216), .X(n51138) );
  nor_x1_sg U68405 ( .A(n20434), .B(n46376), .X(n20432) );
  nor_x1_sg U68406 ( .A(n6240), .B(n46354), .X(n20433) );
  inv_x1_sg U68407 ( .A(n20434), .X(n46354) );
  nor_x1_sg U68408 ( .A(n21167), .B(n46549), .X(n21165) );
  nor_x1_sg U68409 ( .A(n42295), .B(n46538), .X(n21166) );
  inv_x1_sg U68410 ( .A(n21167), .X(n46538) );
  nor_x1_sg U68411 ( .A(n19933), .B(n46557), .X(n19931) );
  nor_x1_sg U68412 ( .A(n42283), .B(n46511), .X(n19932) );
  inv_x1_sg U68413 ( .A(n19933), .X(n46511) );
  nor_x1_sg U68414 ( .A(n19900), .B(n19899), .X(n19897) );
  nand_x1_sg U68415 ( .A(n19899), .B(n19900), .X(n19898) );
  nor_x1_sg U68416 ( .A(n46427), .B(n20143), .X(n20296) );
  nor_x1_sg U68417 ( .A(n41532), .B(n20298), .X(n20297) );
  inv_x1_sg U68418 ( .A(n20298), .X(n46427) );
  nor_x1_sg U68419 ( .A(n46345), .B(n19478), .X(n19475) );
  nor_x1_sg U68420 ( .A(n41531), .B(n19477), .X(n19476) );
  inv_x1_sg U68421 ( .A(n19477), .X(n46345) );
  nor_x1_sg U68422 ( .A(n46499), .B(n21341), .X(n21338) );
  nor_x1_sg U68423 ( .A(n41969), .B(n21340), .X(n21339) );
  inv_x1_sg U68424 ( .A(n21340), .X(n46499) );
  nor_x1_sg U68425 ( .A(n46529), .B(n19504), .X(n19501) );
  nor_x1_sg U68426 ( .A(n41971), .B(n19503), .X(n19502) );
  inv_x1_sg U68427 ( .A(n19503), .X(n46529) );
  nor_x1_sg U68428 ( .A(n45907), .B(n20677), .X(n20674) );
  nor_x1_sg U68429 ( .A(n42199), .B(n20676), .X(n20675) );
  inv_x1_sg U68430 ( .A(n20676), .X(n45907) );
  nor_x1_sg U68431 ( .A(n45897), .B(n20037), .X(n20034) );
  nor_x1_sg U68432 ( .A(n42200), .B(n20036), .X(n20035) );
  inv_x1_sg U68433 ( .A(n20036), .X(n45897) );
  nor_x1_sg U68434 ( .A(n45887), .B(n19233), .X(n19230) );
  nor_x1_sg U68435 ( .A(n42217), .B(n19232), .X(n19231) );
  inv_x1_sg U68436 ( .A(n19232), .X(n45887) );
  nor_x1_sg U68437 ( .A(n46548), .B(n20999), .X(n21174) );
  nor_x1_sg U68438 ( .A(n42260), .B(n21176), .X(n21175) );
  inv_x1_sg U68439 ( .A(n21176), .X(n46548) );
  nor_x1_sg U68440 ( .A(n46233), .B(n46240), .X(n21308) );
  nor_x1_sg U68441 ( .A(n42270), .B(n21310), .X(n21309) );
  inv_x1_sg U68442 ( .A(n21310), .X(n46233) );
  nor_x1_sg U68443 ( .A(n46188), .B(n46194), .X(n21303) );
  nor_x1_sg U68444 ( .A(n42269), .B(n21305), .X(n21304) );
  inv_x1_sg U68445 ( .A(n21305), .X(n46188) );
  nor_x1_sg U68446 ( .A(n46142), .B(n46149), .X(n21298) );
  nor_x1_sg U68447 ( .A(n42267), .B(n21300), .X(n21299) );
  inv_x1_sg U68448 ( .A(n21300), .X(n46142) );
  nor_x1_sg U68449 ( .A(n46097), .B(n46103), .X(n21293) );
  nor_x1_sg U68450 ( .A(n42266), .B(n21295), .X(n21294) );
  inv_x1_sg U68451 ( .A(n21295), .X(n46097) );
  nor_x1_sg U68452 ( .A(n46051), .B(n46058), .X(n21288) );
  nor_x1_sg U68453 ( .A(n42265), .B(n21290), .X(n21289) );
  inv_x1_sg U68454 ( .A(n21290), .X(n46051) );
  nor_x1_sg U68455 ( .A(n46006), .B(n46012), .X(n21283) );
  nor_x1_sg U68456 ( .A(n42264), .B(n21285), .X(n21284) );
  inv_x1_sg U68457 ( .A(n21285), .X(n46006) );
  nor_x1_sg U68458 ( .A(n45961), .B(n45967), .X(n21278) );
  nor_x1_sg U68459 ( .A(n42263), .B(n21280), .X(n21279) );
  inv_x1_sg U68460 ( .A(n21280), .X(n45961) );
  nor_x1_sg U68461 ( .A(n46279), .B(n46285), .X(n21313) );
  nor_x1_sg U68462 ( .A(n42271), .B(n21315), .X(n21314) );
  inv_x1_sg U68463 ( .A(n21315), .X(n46279) );
  nor_x1_sg U68464 ( .A(n46324), .B(n46331), .X(n21318) );
  nor_x1_sg U68465 ( .A(n42272), .B(n21320), .X(n21319) );
  inv_x1_sg U68466 ( .A(n21320), .X(n46324) );
  nor_x1_sg U68467 ( .A(n46366), .B(n46372), .X(n21323) );
  nor_x1_sg U68468 ( .A(n42273), .B(n21325), .X(n21324) );
  inv_x1_sg U68469 ( .A(n21325), .X(n46366) );
  nor_x1_sg U68470 ( .A(n46413), .B(n46420), .X(n21328) );
  nor_x1_sg U68471 ( .A(n42274), .B(n21330), .X(n21329) );
  inv_x1_sg U68472 ( .A(n21330), .X(n46413) );
  nor_x1_sg U68473 ( .A(n46315), .B(n46334), .X(n20549) );
  nor_x1_sg U68474 ( .A(n42296), .B(n20551), .X(n20550) );
  inv_x1_sg U68475 ( .A(n20551), .X(n46315) );
  nor_x1_sg U68476 ( .A(n46270), .B(n46288), .X(n20544) );
  nor_x1_sg U68477 ( .A(n42297), .B(n20546), .X(n20545) );
  inv_x1_sg U68478 ( .A(n20546), .X(n46270) );
  nor_x1_sg U68479 ( .A(n46224), .B(n46243), .X(n20539) );
  nor_x1_sg U68480 ( .A(n42231), .B(n20541), .X(n20540) );
  inv_x1_sg U68481 ( .A(n20541), .X(n46224) );
  nor_x1_sg U68482 ( .A(n46179), .B(n46197), .X(n20534) );
  nor_x1_sg U68483 ( .A(n42299), .B(n20536), .X(n20535) );
  inv_x1_sg U68484 ( .A(n20536), .X(n46179) );
  nor_x1_sg U68485 ( .A(n46133), .B(n46152), .X(n20529) );
  nor_x1_sg U68486 ( .A(n42232), .B(n20531), .X(n20530) );
  inv_x1_sg U68487 ( .A(n20531), .X(n46133) );
  nor_x1_sg U68488 ( .A(n46088), .B(n46106), .X(n20524) );
  nor_x1_sg U68489 ( .A(n42234), .B(n20526), .X(n20525) );
  inv_x1_sg U68490 ( .A(n20526), .X(n46088) );
  nor_x1_sg U68491 ( .A(n46042), .B(n46061), .X(n20519) );
  nor_x1_sg U68492 ( .A(n42301), .B(n20521), .X(n20520) );
  inv_x1_sg U68493 ( .A(n20521), .X(n46042) );
  nor_x1_sg U68494 ( .A(n45997), .B(n46015), .X(n20514) );
  nor_x1_sg U68495 ( .A(n42233), .B(n20516), .X(n20515) );
  inv_x1_sg U68496 ( .A(n20516), .X(n45997) );
  nor_x1_sg U68497 ( .A(n45952), .B(n45970), .X(n20509) );
  nor_x1_sg U68498 ( .A(n42300), .B(n20511), .X(n20510) );
  inv_x1_sg U68499 ( .A(n20511), .X(n45952) );
  nor_x1_sg U68500 ( .A(n46461), .B(n46467), .X(n21333) );
  nor_x1_sg U68501 ( .A(n42275), .B(n21335), .X(n21334) );
  inv_x1_sg U68502 ( .A(n21335), .X(n46461) );
  nor_x1_sg U68503 ( .A(n46306), .B(n46337), .X(n19892) );
  nor_x1_sg U68504 ( .A(n42294), .B(n19894), .X(n19893) );
  inv_x1_sg U68505 ( .A(n19894), .X(n46306) );
  nor_x1_sg U68506 ( .A(n46261), .B(n46291), .X(n19887) );
  nor_x1_sg U68507 ( .A(n42293), .B(n19889), .X(n19888) );
  inv_x1_sg U68508 ( .A(n19889), .X(n46261) );
  nor_x1_sg U68509 ( .A(n46215), .B(n46246), .X(n19882) );
  nor_x1_sg U68510 ( .A(n42292), .B(n19884), .X(n19883) );
  inv_x1_sg U68511 ( .A(n19884), .X(n46215) );
  nor_x1_sg U68512 ( .A(n46170), .B(n46200), .X(n19877) );
  nor_x1_sg U68513 ( .A(n42291), .B(n19879), .X(n19878) );
  inv_x1_sg U68514 ( .A(n19879), .X(n46170) );
  nor_x1_sg U68515 ( .A(n46124), .B(n46155), .X(n19872) );
  nor_x1_sg U68516 ( .A(n42286), .B(n19874), .X(n19873) );
  inv_x1_sg U68517 ( .A(n19874), .X(n46124) );
  nor_x1_sg U68518 ( .A(n46079), .B(n46109), .X(n19867) );
  nor_x1_sg U68519 ( .A(n42290), .B(n19869), .X(n19868) );
  inv_x1_sg U68520 ( .A(n19869), .X(n46079) );
  nor_x1_sg U68521 ( .A(n46033), .B(n46064), .X(n19862) );
  nor_x1_sg U68522 ( .A(n42289), .B(n19864), .X(n19863) );
  inv_x1_sg U68523 ( .A(n19864), .X(n46033) );
  nor_x1_sg U68524 ( .A(n45988), .B(n46018), .X(n19857) );
  nor_x1_sg U68525 ( .A(n42288), .B(n19859), .X(n19858) );
  inv_x1_sg U68526 ( .A(n19859), .X(n45988) );
  nor_x1_sg U68527 ( .A(n45943), .B(n45973), .X(n19852) );
  nor_x1_sg U68528 ( .A(n42287), .B(n19854), .X(n19853) );
  inv_x1_sg U68529 ( .A(n19854), .X(n45943) );
  nor_x1_sg U68530 ( .A(n6071), .B(n20126), .X(n20125) );
  nand_x1_sg U68531 ( .A(n20126), .B(n6071), .X(n20127) );
  nor_x1_sg U68532 ( .A(n38617), .B(n19729), .X(n19728) );
  nand_x1_sg U68533 ( .A(n19729), .B(n5965), .X(n19730) );
  nor_x1_sg U68534 ( .A(n42334), .B(n19333), .X(n19332) );
  nand_x1_sg U68535 ( .A(n19333), .B(n38695), .X(n19334) );
  nor_x1_sg U68536 ( .A(n38668), .B(n19496), .X(n19495) );
  nand_x1_sg U68537 ( .A(n19496), .B(n6087), .X(n19497) );
  nor_x1_sg U68538 ( .A(n6024), .B(n19926), .X(n19925) );
  nand_x1_sg U68539 ( .A(n19926), .B(n6024), .X(n19927) );
  nor_x1_sg U68540 ( .A(n21445), .B(n21446), .X(n21444) );
  nand_x1_sg U68541 ( .A(n21446), .B(n21445), .X(n21447) );
  nor_x1_sg U68542 ( .A(n45078), .B(n28269), .X(n28268) );
  nand_x1_sg U68543 ( .A(n28269), .B(n45078), .X(n28270) );
  nor_x1_sg U68544 ( .A(n42023), .B(n20782), .X(n20781) );
  nand_x1_sg U68545 ( .A(n20782), .B(n42023), .X(n20783) );
  nor_x1_sg U68546 ( .A(n42024), .B(n19483), .X(n19482) );
  nand_x1_sg U68547 ( .A(n19483), .B(n42024), .X(n19484) );
  inv_x1_sg U68548 ( .A(n24937), .X(n51140) );
  inv_x1_sg U68549 ( .A(n27616), .X(n44971) );
  nor_x1_sg U68550 ( .A(n38191), .B(n22574), .X(n27615) );
  inv_x1_sg U68551 ( .A(n28462), .X(n44966) );
  nor_x1_sg U68552 ( .A(n38192), .B(n22578), .X(n28461) );
  inv_x1_sg U68553 ( .A(n27191), .X(n44973) );
  nor_x1_sg U68554 ( .A(n38127), .B(n22566), .X(n27190) );
  nor_x1_sg U68555 ( .A(n46541), .B(n21200), .X(n21344) );
  nor_x1_sg U68556 ( .A(n41968), .B(n21346), .X(n21345) );
  inv_x1_sg U68557 ( .A(n21346), .X(n46541) );
  nor_x1_sg U68558 ( .A(n46359), .B(n20747), .X(n20744) );
  nor_x1_sg U68559 ( .A(n42214), .B(n20746), .X(n20745) );
  inv_x1_sg U68560 ( .A(n20746), .X(n46359) );
  nor_x1_sg U68561 ( .A(n46317), .B(n20740), .X(n20737) );
  nor_x1_sg U68562 ( .A(n42212), .B(n20739), .X(n20738) );
  inv_x1_sg U68563 ( .A(n20739), .X(n46317) );
  nor_x1_sg U68564 ( .A(n46272), .B(n20733), .X(n20730) );
  nor_x1_sg U68565 ( .A(n42210), .B(n20732), .X(n20731) );
  inv_x1_sg U68566 ( .A(n20732), .X(n46272) );
  nor_x1_sg U68567 ( .A(n46226), .B(n20726), .X(n20723) );
  nor_x1_sg U68568 ( .A(n42152), .B(n20725), .X(n20724) );
  inv_x1_sg U68569 ( .A(n20725), .X(n46226) );
  nor_x1_sg U68570 ( .A(n46181), .B(n20719), .X(n20716) );
  nor_x1_sg U68571 ( .A(n42207), .B(n20718), .X(n20717) );
  inv_x1_sg U68572 ( .A(n20718), .X(n46181) );
  nor_x1_sg U68573 ( .A(n46135), .B(n20712), .X(n20709) );
  nor_x1_sg U68574 ( .A(n42151), .B(n20711), .X(n20710) );
  inv_x1_sg U68575 ( .A(n20711), .X(n46135) );
  nor_x1_sg U68576 ( .A(n46090), .B(n20705), .X(n20702) );
  nor_x1_sg U68577 ( .A(n42150), .B(n20704), .X(n20703) );
  inv_x1_sg U68578 ( .A(n20704), .X(n46090) );
  nor_x1_sg U68579 ( .A(n46044), .B(n20698), .X(n20695) );
  nor_x1_sg U68580 ( .A(n42204), .B(n20697), .X(n20696) );
  inv_x1_sg U68581 ( .A(n20697), .X(n46044) );
  nor_x1_sg U68582 ( .A(n45999), .B(n20691), .X(n20688) );
  nor_x1_sg U68583 ( .A(n42148), .B(n20690), .X(n20689) );
  inv_x1_sg U68584 ( .A(n20690), .X(n45999) );
  nor_x1_sg U68585 ( .A(n45954), .B(n20684), .X(n20681) );
  nor_x1_sg U68586 ( .A(n42201), .B(n20683), .X(n20682) );
  inv_x1_sg U68587 ( .A(n20683), .X(n45954) );
  nor_x1_sg U68588 ( .A(n46308), .B(n20100), .X(n20097) );
  nor_x1_sg U68589 ( .A(n42213), .B(n20099), .X(n20098) );
  inv_x1_sg U68590 ( .A(n20099), .X(n46308) );
  nor_x1_sg U68591 ( .A(n46263), .B(n20093), .X(n20090) );
  nor_x1_sg U68592 ( .A(n42211), .B(n20092), .X(n20091) );
  inv_x1_sg U68593 ( .A(n20092), .X(n46263) );
  nor_x1_sg U68594 ( .A(n46217), .B(n20086), .X(n20083) );
  nor_x1_sg U68595 ( .A(n42209), .B(n20085), .X(n20084) );
  inv_x1_sg U68596 ( .A(n20085), .X(n46217) );
  nor_x1_sg U68597 ( .A(n46172), .B(n20079), .X(n20076) );
  nor_x1_sg U68598 ( .A(n42208), .B(n20078), .X(n20077) );
  inv_x1_sg U68599 ( .A(n20078), .X(n46172) );
  nor_x1_sg U68600 ( .A(n46126), .B(n20072), .X(n20069) );
  nor_x1_sg U68601 ( .A(n42206), .B(n20071), .X(n20070) );
  inv_x1_sg U68602 ( .A(n20071), .X(n46126) );
  nor_x1_sg U68603 ( .A(n46081), .B(n20065), .X(n20062) );
  nor_x1_sg U68604 ( .A(n42205), .B(n20064), .X(n20063) );
  inv_x1_sg U68605 ( .A(n20064), .X(n46081) );
  nor_x1_sg U68606 ( .A(n46035), .B(n20058), .X(n20055) );
  nor_x1_sg U68607 ( .A(n42149), .B(n20057), .X(n20056) );
  inv_x1_sg U68608 ( .A(n20057), .X(n46035) );
  nor_x1_sg U68609 ( .A(n45990), .B(n20051), .X(n20048) );
  nor_x1_sg U68610 ( .A(n42203), .B(n20050), .X(n20049) );
  inv_x1_sg U68611 ( .A(n20050), .X(n45990) );
  nor_x1_sg U68612 ( .A(n45945), .B(n20044), .X(n20041) );
  nor_x1_sg U68613 ( .A(n42202), .B(n20043), .X(n20042) );
  inv_x1_sg U68614 ( .A(n20043), .X(n45945) );
  nor_x1_sg U68615 ( .A(n46299), .B(n19296), .X(n19293) );
  nor_x1_sg U68616 ( .A(n42224), .B(n19295), .X(n19294) );
  inv_x1_sg U68617 ( .A(n19295), .X(n46299) );
  nor_x1_sg U68618 ( .A(n46254), .B(n19289), .X(n19286) );
  nor_x1_sg U68619 ( .A(n42223), .B(n19288), .X(n19287) );
  inv_x1_sg U68620 ( .A(n19288), .X(n46254) );
  nor_x1_sg U68621 ( .A(n46208), .B(n19282), .X(n19279) );
  nor_x1_sg U68622 ( .A(n42222), .B(n19281), .X(n19280) );
  inv_x1_sg U68623 ( .A(n19281), .X(n46208) );
  nor_x1_sg U68624 ( .A(n46163), .B(n19275), .X(n19272) );
  nor_x1_sg U68625 ( .A(n42221), .B(n19274), .X(n19273) );
  inv_x1_sg U68626 ( .A(n19274), .X(n46163) );
  nor_x1_sg U68627 ( .A(n46117), .B(n19268), .X(n19265) );
  nor_x1_sg U68628 ( .A(n42216), .B(n19267), .X(n19266) );
  inv_x1_sg U68629 ( .A(n19267), .X(n46117) );
  nor_x1_sg U68630 ( .A(n46072), .B(n19261), .X(n19258) );
  nor_x1_sg U68631 ( .A(n42220), .B(n19260), .X(n19259) );
  inv_x1_sg U68632 ( .A(n19260), .X(n46072) );
  nor_x1_sg U68633 ( .A(n46026), .B(n19254), .X(n19251) );
  nor_x1_sg U68634 ( .A(n42219), .B(n19253), .X(n19252) );
  inv_x1_sg U68635 ( .A(n19253), .X(n46026) );
  nor_x1_sg U68636 ( .A(n45981), .B(n19247), .X(n19244) );
  nor_x1_sg U68637 ( .A(n42261), .B(n19246), .X(n19245) );
  inv_x1_sg U68638 ( .A(n19246), .X(n45981) );
  nor_x1_sg U68639 ( .A(n45936), .B(n19240), .X(n19237) );
  nor_x1_sg U68640 ( .A(n42218), .B(n19239), .X(n19238) );
  inv_x1_sg U68641 ( .A(n19239), .X(n45936) );
  nor_x1_sg U68642 ( .A(n46418), .B(n21517), .X(n21516) );
  nand_x1_sg U68643 ( .A(n21517), .B(n46418), .X(n21518) );
  nor_x1_sg U68644 ( .A(n46329), .B(n21504), .X(n21503) );
  nand_x1_sg U68645 ( .A(n21504), .B(n46329), .X(n21505) );
  nor_x1_sg U68646 ( .A(n46238), .B(n21491), .X(n21490) );
  nand_x1_sg U68647 ( .A(n21491), .B(n46238), .X(n21492) );
  nor_x1_sg U68648 ( .A(n46147), .B(n21478), .X(n21477) );
  nand_x1_sg U68649 ( .A(n21478), .B(n46147), .X(n21479) );
  nor_x1_sg U68650 ( .A(n46056), .B(n21465), .X(n21464) );
  nand_x1_sg U68651 ( .A(n21465), .B(n46056), .X(n21466) );
  nor_x1_sg U68652 ( .A(n45965), .B(n21452), .X(n21451) );
  nand_x1_sg U68653 ( .A(n21452), .B(n45965), .X(n21453) );
  nor_x1_sg U68654 ( .A(n6051), .B(n19935), .X(n19934) );
  nand_x1_sg U68655 ( .A(n19935), .B(n6051), .X(n19936) );
  nor_x1_sg U68656 ( .A(n21523), .B(n21524), .X(n21522) );
  nand_x1_sg U68657 ( .A(n21524), .B(n21523), .X(n21525) );
  nor_x1_sg U68658 ( .A(n21510), .B(n21511), .X(n21509) );
  nand_x1_sg U68659 ( .A(n21511), .B(n21510), .X(n21512) );
  nor_x1_sg U68660 ( .A(n21497), .B(n21498), .X(n21496) );
  nand_x1_sg U68661 ( .A(n21498), .B(n21497), .X(n21499) );
  nor_x1_sg U68662 ( .A(n21484), .B(n21485), .X(n21483) );
  nand_x1_sg U68663 ( .A(n21485), .B(n21484), .X(n21486) );
  nor_x1_sg U68664 ( .A(n21471), .B(n21472), .X(n21470) );
  nand_x1_sg U68665 ( .A(n21472), .B(n21471), .X(n21473) );
  nor_x1_sg U68666 ( .A(n21458), .B(n21459), .X(n21457) );
  nand_x1_sg U68667 ( .A(n21459), .B(n21458), .X(n21460) );
  nand_x1_sg U68668 ( .A(n26767), .B(n39391), .X(n29271) );
  nor_x1_sg U68669 ( .A(n20774), .B(n42339), .X(n20772) );
  nand_x1_sg U68670 ( .A(n38600), .B(n20774), .X(n20773) );
  nor_x1_sg U68671 ( .A(n19491), .B(n19490), .X(n19488) );
  nand_x1_sg U68672 ( .A(n19490), .B(n19491), .X(n19489) );
  nor_x1_sg U68673 ( .A(n46406), .B(n20754), .X(n20751) );
  nor_x1_sg U68674 ( .A(n42256), .B(n20753), .X(n20752) );
  inv_x1_sg U68675 ( .A(n20753), .X(n46406) );
  nor_x1_sg U68676 ( .A(n46454), .B(n20761), .X(n20758) );
  nor_x1_sg U68677 ( .A(n42257), .B(n20760), .X(n20759) );
  inv_x1_sg U68678 ( .A(n20760), .X(n46454) );
  nor_x1_sg U68679 ( .A(n46492), .B(n20768), .X(n20765) );
  nor_x1_sg U68680 ( .A(n42259), .B(n20767), .X(n20766) );
  inv_x1_sg U68681 ( .A(n20767), .X(n46492) );
  nor_x1_sg U68682 ( .A(n45913), .B(n45922), .X(n21082) );
  nor_x1_sg U68683 ( .A(n42302), .B(n21084), .X(n21083) );
  inv_x1_sg U68684 ( .A(n21084), .X(n45913) );
  nor_x1_sg U68685 ( .A(n45903), .B(n45925), .X(n20373) );
  nor_x1_sg U68686 ( .A(n42298), .B(n20375), .X(n20374) );
  inv_x1_sg U68687 ( .A(n20375), .X(n45903) );
  nor_x1_sg U68688 ( .A(n45893), .B(n45928), .X(n19640) );
  nor_x1_sg U68689 ( .A(n42285), .B(n19642), .X(n19641) );
  inv_x1_sg U68690 ( .A(n19642), .X(n45893) );
  nor_x1_sg U68691 ( .A(n46490), .B(n46507), .X(n20131) );
  nor_x1_sg U68692 ( .A(n6101), .B(n20133), .X(n20132) );
  inv_x1_sg U68693 ( .A(n20133), .X(n46490) );
  nor_x1_sg U68694 ( .A(n45125), .B(n28275), .X(n28274) );
  nand_x1_sg U68695 ( .A(n28275), .B(n45125), .X(n28276) );
  nor_x1_sg U68696 ( .A(n45170), .B(n28281), .X(n28280) );
  nand_x1_sg U68697 ( .A(n28281), .B(n45170), .X(n28282) );
  nor_x1_sg U68698 ( .A(n45216), .B(n28287), .X(n28286) );
  nand_x1_sg U68699 ( .A(n28287), .B(n45216), .X(n28288) );
  nor_x1_sg U68700 ( .A(n45261), .B(n28293), .X(n28292) );
  nand_x1_sg U68701 ( .A(n28293), .B(n45261), .X(n28294) );
  nor_x1_sg U68702 ( .A(n45306), .B(n28299), .X(n28298) );
  nand_x1_sg U68703 ( .A(n28299), .B(n45306), .X(n28300) );
  nor_x1_sg U68704 ( .A(n45351), .B(n28305), .X(n28304) );
  nand_x1_sg U68705 ( .A(n28305), .B(n45351), .X(n28306) );
  nor_x1_sg U68706 ( .A(n45397), .B(n28311), .X(n28310) );
  nand_x1_sg U68707 ( .A(n28311), .B(n45397), .X(n28312) );
  nor_x1_sg U68708 ( .A(n38670), .B(n19905), .X(n19904) );
  nand_x1_sg U68709 ( .A(n19905), .B(n6161), .X(n19906) );
  nor_x1_sg U68710 ( .A(n6226), .B(n19301), .X(n19300) );
  nand_x1_sg U68711 ( .A(n19301), .B(n38604), .X(n19302) );
  nor_x1_sg U68712 ( .A(n45067), .B(n29154), .X(n29153) );
  nor_x1_sg U68713 ( .A(n29155), .B(n45022), .X(n29152) );
  inv_x1_sg U68714 ( .A(n29155), .X(n45067) );
  nor_x1_sg U68715 ( .A(n45159), .B(n29166), .X(n29165) );
  nor_x1_sg U68716 ( .A(n29167), .B(n45112), .X(n29164) );
  inv_x1_sg U68717 ( .A(n29167), .X(n45159) );
  nor_x1_sg U68718 ( .A(n45250), .B(n29178), .X(n29177) );
  nor_x1_sg U68719 ( .A(n29179), .B(n45203), .X(n29176) );
  inv_x1_sg U68720 ( .A(n29179), .X(n45250) );
  nor_x1_sg U68721 ( .A(n45340), .B(n29190), .X(n29189) );
  nor_x1_sg U68722 ( .A(n29191), .B(n45294), .X(n29188) );
  inv_x1_sg U68723 ( .A(n29191), .X(n45340) );
  nor_x1_sg U68724 ( .A(n45431), .B(n29202), .X(n29201) );
  nor_x1_sg U68725 ( .A(n29203), .B(n45384), .X(n29200) );
  inv_x1_sg U68726 ( .A(n29203), .X(n45431) );
  nor_x1_sg U68727 ( .A(n45520), .B(n29214), .X(n29213) );
  nor_x1_sg U68728 ( .A(n29215), .B(n45474), .X(n29212) );
  inv_x1_sg U68729 ( .A(n29215), .X(n45520) );
  nor_x1_sg U68730 ( .A(n45609), .B(n29089), .X(n29225) );
  nor_x1_sg U68731 ( .A(n29226), .B(n45563), .X(n29224) );
  inv_x1_sg U68732 ( .A(n29226), .X(n45609) );
  nor_x1_sg U68733 ( .A(n45918), .B(n21603), .X(n21602) );
  nor_x1_sg U68734 ( .A(n21604), .B(n45870), .X(n21601) );
  inv_x1_sg U68735 ( .A(n21604), .X(n45918) );
  nor_x1_sg U68736 ( .A(n46464), .B(n21538), .X(n21674) );
  nor_x1_sg U68737 ( .A(n21675), .B(n46415), .X(n21673) );
  inv_x1_sg U68738 ( .A(n21675), .X(n46464) );
  nor_x1_sg U68739 ( .A(n46369), .B(n21663), .X(n21662) );
  nor_x1_sg U68740 ( .A(n21664), .B(n46326), .X(n21661) );
  inv_x1_sg U68741 ( .A(n21664), .X(n46369) );
  nor_x1_sg U68742 ( .A(n46282), .B(n21651), .X(n21650) );
  nor_x1_sg U68743 ( .A(n21652), .B(n46235), .X(n21649) );
  inv_x1_sg U68744 ( .A(n21652), .X(n46282) );
  nor_x1_sg U68745 ( .A(n46191), .B(n21639), .X(n21638) );
  nor_x1_sg U68746 ( .A(n21640), .B(n46144), .X(n21637) );
  inv_x1_sg U68747 ( .A(n21640), .X(n46191) );
  nor_x1_sg U68748 ( .A(n46100), .B(n21627), .X(n21626) );
  nor_x1_sg U68749 ( .A(n21628), .B(n46053), .X(n21625) );
  inv_x1_sg U68750 ( .A(n21628), .X(n46100) );
  nor_x1_sg U68751 ( .A(n46009), .B(n21615), .X(n21614) );
  nor_x1_sg U68752 ( .A(n21616), .B(n45963), .X(n21613) );
  inv_x1_sg U68753 ( .A(n21616), .X(n46009) );
  nor_x1_sg U68754 ( .A(n44998), .B(n28133), .X(n28130) );
  nor_x1_sg U68755 ( .A(n41540), .B(n28132), .X(n28131) );
  inv_x1_sg U68756 ( .A(n28132), .X(n44998) );
  inv_x1_sg U68757 ( .A(n28255), .X(n44968) );
  nor_x1_sg U68758 ( .A(n38193), .B(n22584), .X(n28254) );
  inv_x1_sg U68759 ( .A(n23543), .X(n51137) );
  nor_x1_sg U68760 ( .A(n6457), .B(n21116), .X(n21231) );
  nand_x1_sg U68761 ( .A(n21233), .B(n38568), .X(n21232) );
  nor_x1_sg U68762 ( .A(n6501), .B(n21110), .X(n21234) );
  nand_x1_sg U68763 ( .A(n21236), .B(n38569), .X(n21235) );
  nor_x1_sg U68764 ( .A(n6546), .B(n21104), .X(n21237) );
  nand_x1_sg U68765 ( .A(n21239), .B(n38570), .X(n21238) );
  nor_x1_sg U68766 ( .A(n6590), .B(n21098), .X(n21240) );
  nand_x1_sg U68767 ( .A(n21242), .B(n38571), .X(n21241) );
  nor_x1_sg U68768 ( .A(n6635), .B(n21092), .X(n21243) );
  nand_x1_sg U68769 ( .A(n21245), .B(n38591), .X(n21244) );
  nor_x1_sg U68770 ( .A(n6412), .B(n21122), .X(n21228) );
  nand_x1_sg U68771 ( .A(n21230), .B(n38567), .X(n21229) );
  nor_x1_sg U68772 ( .A(n6368), .B(n21128), .X(n21225) );
  nand_x1_sg U68773 ( .A(n21227), .B(n38566), .X(n21226) );
  nor_x1_sg U68774 ( .A(n6323), .B(n21134), .X(n21222) );
  nand_x1_sg U68775 ( .A(n21224), .B(n38565), .X(n21223) );
  nor_x1_sg U68776 ( .A(n6279), .B(n21140), .X(n21219) );
  nand_x1_sg U68777 ( .A(n21221), .B(n38564), .X(n21220) );
  nor_x1_sg U68778 ( .A(n6329), .B(n20425), .X(n20454) );
  nand_x1_sg U68779 ( .A(n20456), .B(n38576), .X(n20455) );
  nor_x1_sg U68780 ( .A(n6374), .B(n20419), .X(n20457) );
  nand_x1_sg U68781 ( .A(n20459), .B(n38577), .X(n20458) );
  nor_x1_sg U68782 ( .A(n6418), .B(n20413), .X(n20460) );
  nand_x1_sg U68783 ( .A(n20462), .B(n38578), .X(n20461) );
  nor_x1_sg U68784 ( .A(n6463), .B(n20407), .X(n20463) );
  nand_x1_sg U68785 ( .A(n20465), .B(n38579), .X(n20464) );
  nor_x1_sg U68786 ( .A(n6507), .B(n20401), .X(n20466) );
  nand_x1_sg U68787 ( .A(n20468), .B(n38580), .X(n20467) );
  nor_x1_sg U68788 ( .A(n6552), .B(n20395), .X(n20469) );
  nand_x1_sg U68789 ( .A(n20471), .B(n38581), .X(n20470) );
  nor_x1_sg U68790 ( .A(n6596), .B(n20389), .X(n20472) );
  nand_x1_sg U68791 ( .A(n20474), .B(n38582), .X(n20473) );
  nor_x1_sg U68792 ( .A(n6641), .B(n20383), .X(n20475) );
  nand_x1_sg U68793 ( .A(n20477), .B(n38592), .X(n20476) );
  nor_x1_sg U68794 ( .A(n6234), .B(n21146), .X(n21216) );
  nand_x1_sg U68795 ( .A(n21218), .B(n38563), .X(n21217) );
  nor_x1_sg U68796 ( .A(n6188), .B(n21152), .X(n21213) );
  nand_x1_sg U68797 ( .A(n21215), .B(n38572), .X(n21214) );
  nor_x1_sg U68798 ( .A(n6142), .B(n21158), .X(n21210) );
  nand_x1_sg U68799 ( .A(n21212), .B(n38573), .X(n21211) );
  nor_x1_sg U68800 ( .A(n6300), .B(n19692), .X(n19797) );
  nand_x1_sg U68801 ( .A(n19799), .B(n38584), .X(n19798) );
  nor_x1_sg U68802 ( .A(n6344), .B(n19686), .X(n19800) );
  nand_x1_sg U68803 ( .A(n19802), .B(n38585), .X(n19801) );
  nor_x1_sg U68804 ( .A(n6389), .B(n19680), .X(n19803) );
  nand_x1_sg U68805 ( .A(n19805), .B(n38586), .X(n19804) );
  nor_x1_sg U68806 ( .A(n6433), .B(n19674), .X(n19806) );
  nand_x1_sg U68807 ( .A(n19808), .B(n38587), .X(n19807) );
  nor_x1_sg U68808 ( .A(n6478), .B(n19668), .X(n19809) );
  nand_x1_sg U68809 ( .A(n19811), .B(n38588), .X(n19810) );
  nor_x1_sg U68810 ( .A(n6522), .B(n19662), .X(n19812) );
  nand_x1_sg U68811 ( .A(n19814), .B(n38589), .X(n19813) );
  nor_x1_sg U68812 ( .A(n6567), .B(n19656), .X(n19815) );
  nand_x1_sg U68813 ( .A(n19817), .B(n38590), .X(n19816) );
  nor_x1_sg U68814 ( .A(n6611), .B(n19650), .X(n19818) );
  nand_x1_sg U68815 ( .A(n19820), .B(n38593), .X(n19819) );
  nand_x1_sg U68816 ( .A(n17465), .B(n41660), .X(n42385) );
  nand_x1_sg U68817 ( .A(n26119), .B(n26120), .X(n26117) );
  nor_x1_sg U68818 ( .A(n26119), .B(n26120), .X(n26118) );
  nor_x1_sg U68819 ( .A(n6096), .B(n21164), .X(n21207) );
  nand_x1_sg U68820 ( .A(n21209), .B(n38574), .X(n21208) );
  nor_x1_sg U68821 ( .A(n50548), .B(n16834), .X(n26034) );
  nor_x1_sg U68822 ( .A(n26035), .B(n41526), .X(n26033) );
  nor_x1_sg U68823 ( .A(n28255), .B(n28258), .X(n28256) );
  nand_x1_sg U68824 ( .A(n28258), .B(n28255), .X(n28257) );
  nor_x1_sg U68825 ( .A(n21072), .B(n21071), .X(n21069) );
  nand_x1_sg U68826 ( .A(n21071), .B(n21072), .X(n21070) );
  nor_x1_sg U68827 ( .A(n20664), .B(n20663), .X(n20661) );
  nand_x1_sg U68828 ( .A(n20663), .B(n20664), .X(n20662) );
  nor_x1_sg U68829 ( .A(n20493), .B(n20492), .X(n20490) );
  nand_x1_sg U68830 ( .A(n20492), .B(n20493), .X(n20491) );
  nor_x1_sg U68831 ( .A(n20024), .B(n20023), .X(n20021) );
  nand_x1_sg U68832 ( .A(n20023), .B(n20024), .X(n20022) );
  nor_x1_sg U68833 ( .A(n20363), .B(n20362), .X(n20360) );
  nand_x1_sg U68834 ( .A(n20362), .B(n20363), .X(n20361) );
  nor_x1_sg U68835 ( .A(n19836), .B(n19835), .X(n19833) );
  nand_x1_sg U68836 ( .A(n19835), .B(n19836), .X(n19834) );
  nor_x1_sg U68837 ( .A(n19630), .B(n19629), .X(n19627) );
  nand_x1_sg U68838 ( .A(n19629), .B(n19630), .X(n19628) );
  nor_x1_sg U68839 ( .A(n19397), .B(n19396), .X(n19394) );
  nand_x1_sg U68840 ( .A(n19396), .B(n19397), .X(n19395) );
  nor_x1_sg U68841 ( .A(n21434), .B(n21433), .X(n21431) );
  nand_x1_sg U68842 ( .A(n21433), .B(n21434), .X(n21432) );
  nor_x1_sg U68843 ( .A(n19220), .B(n19219), .X(n19217) );
  nand_x1_sg U68844 ( .A(n19219), .B(n19220), .X(n19218) );
  nor_x1_sg U68845 ( .A(n20203), .B(n20202), .X(n20200) );
  nand_x1_sg U68846 ( .A(n20202), .B(n20203), .X(n20201) );
  nor_x1_sg U68847 ( .A(n21262), .B(n21261), .X(n21259) );
  nand_x1_sg U68848 ( .A(n21261), .B(n21262), .X(n21260) );
  nor_x1_sg U68849 ( .A(n20846), .B(n20845), .X(n20843) );
  nand_x1_sg U68850 ( .A(n20845), .B(n20846), .X(n20844) );
  nor_x1_sg U68851 ( .A(n46357), .B(n46375), .X(n20554) );
  nor_x1_sg U68852 ( .A(n42284), .B(n20556), .X(n20555) );
  inv_x1_sg U68853 ( .A(n20556), .X(n46357) );
  nand_x1_sg U68854 ( .A(n41302), .B(n41660), .X(n18284) );
  nand_x1_sg U68855 ( .A(n23098), .B(n47143), .X(n23097) );
  inv_x1_sg U68856 ( .A(n23098), .X(n47151) );
  nand_x1_sg U68857 ( .A(n23378), .B(n47428), .X(n23377) );
  inv_x1_sg U68858 ( .A(n23378), .X(n47436) );
  nand_x1_sg U68859 ( .A(n23657), .B(n47713), .X(n23656) );
  inv_x1_sg U68860 ( .A(n23657), .X(n47721) );
  nand_x1_sg U68861 ( .A(n23936), .B(n47998), .X(n23935) );
  inv_x1_sg U68862 ( .A(n23936), .X(n48006) );
  nand_x1_sg U68863 ( .A(n24215), .B(n48283), .X(n24214) );
  inv_x1_sg U68864 ( .A(n24215), .X(n48291) );
  nand_x1_sg U68865 ( .A(n24494), .B(n48568), .X(n24493) );
  inv_x1_sg U68866 ( .A(n24494), .X(n48576) );
  nand_x1_sg U68867 ( .A(n24772), .B(n48853), .X(n24771) );
  inv_x1_sg U68868 ( .A(n24772), .X(n48862) );
  nand_x1_sg U68869 ( .A(n25051), .B(n49140), .X(n25050) );
  inv_x1_sg U68870 ( .A(n25051), .X(n49149) );
  nand_x1_sg U68871 ( .A(n25330), .B(n49426), .X(n25329) );
  inv_x1_sg U68872 ( .A(n25330), .X(n49435) );
  nand_x1_sg U68873 ( .A(n25609), .B(n49712), .X(n25608) );
  inv_x1_sg U68874 ( .A(n25609), .X(n49720) );
  nand_x1_sg U68875 ( .A(n25886), .B(n49998), .X(n25885) );
  inv_x1_sg U68876 ( .A(n25886), .X(n50007) );
  nand_x1_sg U68877 ( .A(n26446), .B(n50573), .X(n26445) );
  inv_x1_sg U68878 ( .A(n26446), .X(n50581) );
  nand_x1_sg U68879 ( .A(n26724), .B(n50859), .X(n26723) );
  inv_x1_sg U68880 ( .A(n26724), .X(n50868) );
  nand_x1_sg U68881 ( .A(n41299), .B(n41632), .X(n24658) );
  nor_x1_sg U68882 ( .A(n46802), .B(n26102), .X(n26162) );
  nand_x1_sg U68883 ( .A(n26164), .B(n50300), .X(n26163) );
  nand_x1_sg U68884 ( .A(n26106), .B(n26107), .X(n26105) );
  nor_x1_sg U68885 ( .A(n26106), .B(n26107), .X(n26108) );
  nand_x1_sg U68886 ( .A(n46858), .B(n46850), .X(n22819) );
  nand_x1_sg U68887 ( .A(n22821), .B(n22816), .X(n22820) );
  inv_x1_sg U68888 ( .A(n22821), .X(n46858) );
  nor_x1_sg U68889 ( .A(n26144), .B(n26143), .X(n26141) );
  nand_x1_sg U68890 ( .A(n26143), .B(n26144), .X(n26142) );
  nor_x1_sg U68891 ( .A(n26825), .B(n26791), .X(n26823) );
  nand_x1_sg U68892 ( .A(n26791), .B(n26825), .X(n26824) );
  nor_x1_sg U68893 ( .A(n20974), .B(n20563), .X(n20972) );
  nand_x1_sg U68894 ( .A(n20563), .B(n20974), .X(n20973) );
  nor_x1_sg U68895 ( .A(n6023), .B(n19761), .X(n19758) );
  nand_x1_sg U68896 ( .A(n19760), .B(n38268), .X(n19759) );
  nor_x1_sg U68897 ( .A(n42330), .B(n19773), .X(n19770) );
  nand_x1_sg U68898 ( .A(n19772), .B(n38595), .X(n19771) );
  nand_x1_sg U68899 ( .A(n39479), .B(n42162), .X(n26332) );
  nand_x1_sg U68900 ( .A(n39480), .B(n42058), .X(n23821) );
  nand_x1_sg U68901 ( .A(n39480), .B(n24101), .X(n24100) );
  nand_x1_sg U68902 ( .A(n38942), .B(n24380), .X(n24379) );
  nand_x1_sg U68903 ( .A(n41301), .B(n24937), .X(n24936) );
  nand_x1_sg U68904 ( .A(n41302), .B(n25216), .X(n25215) );
  nand_x1_sg U68905 ( .A(n41300), .B(n25495), .X(n25494) );
  nand_x1_sg U68906 ( .A(n41301), .B(n39123), .X(n26610) );
  nor_x1_sg U68907 ( .A(n19125), .B(n19521), .X(n19520) );
  nand_x1_sg U68908 ( .A(n19521), .B(n19125), .X(n19522) );
  nor_x1_sg U68909 ( .A(n19117), .B(n19518), .X(n19517) );
  nand_x1_sg U68910 ( .A(n19518), .B(n19117), .X(n19519) );
  nor_x1_sg U68911 ( .A(n19119), .B(n19515), .X(n19514) );
  nand_x1_sg U68912 ( .A(n19515), .B(n19119), .X(n19516) );
  nor_x1_sg U68913 ( .A(n20580), .B(n20581), .X(n20579) );
  nand_x1_sg U68914 ( .A(n20581), .B(n20580), .X(n20582) );
  nor_x1_sg U68915 ( .A(n19510), .B(n19512), .X(n19511) );
  nand_x1_sg U68916 ( .A(n19512), .B(n19510), .X(n19513) );
  nor_x1_sg U68917 ( .A(n20574), .B(n20577), .X(n20576) );
  nand_x1_sg U68918 ( .A(n20577), .B(n20574), .X(n20578) );
  nor_x1_sg U68919 ( .A(n19137), .B(n19138), .X(n19136) );
  nand_x1_sg U68920 ( .A(n19138), .B(n19137), .X(n19139) );
  nor_x1_sg U68921 ( .A(n19527), .B(n19528), .X(n19526) );
  nand_x1_sg U68922 ( .A(n19528), .B(n19527), .X(n19529) );
  nor_x1_sg U68923 ( .A(n20568), .B(n20967), .X(n20966) );
  nand_x1_sg U68924 ( .A(n20967), .B(n20568), .X(n20968) );
  nor_x1_sg U68925 ( .A(n19123), .B(n19524), .X(n19523) );
  nand_x1_sg U68926 ( .A(n19524), .B(n19123), .X(n19525) );
  nor_x1_sg U68927 ( .A(n20566), .B(n20970), .X(n20969) );
  nand_x1_sg U68928 ( .A(n20970), .B(n20566), .X(n20971) );
  nor_x1_sg U68929 ( .A(n20960), .B(n20964), .X(n20963) );
  nand_x1_sg U68930 ( .A(n20964), .B(n20960), .X(n20965) );
  nor_x1_sg U68931 ( .A(n23126), .B(n47134), .X(n23125) );
  nand_x1_sg U68932 ( .A(n23406), .B(n42057), .X(n23404) );
  nor_x1_sg U68933 ( .A(n23406), .B(n42057), .X(n23405) );
  nand_x1_sg U68934 ( .A(n23685), .B(n42056), .X(n23683) );
  nor_x1_sg U68935 ( .A(n23685), .B(n42056), .X(n23684) );
  nand_x1_sg U68936 ( .A(n23964), .B(n42055), .X(n23962) );
  nor_x1_sg U68937 ( .A(n23964), .B(n42055), .X(n23963) );
  nand_x1_sg U68938 ( .A(n24243), .B(n42054), .X(n24241) );
  nor_x1_sg U68939 ( .A(n24243), .B(n42054), .X(n24242) );
  nand_x1_sg U68940 ( .A(n24522), .B(n42053), .X(n24520) );
  nor_x1_sg U68941 ( .A(n24522), .B(n42053), .X(n24521) );
  nand_x1_sg U68942 ( .A(n24800), .B(n42052), .X(n24798) );
  nor_x1_sg U68943 ( .A(n24800), .B(n42052), .X(n24799) );
  nand_x1_sg U68944 ( .A(n25079), .B(n42051), .X(n25077) );
  nor_x1_sg U68945 ( .A(n25079), .B(n42051), .X(n25078) );
  nand_x1_sg U68946 ( .A(n25358), .B(n42050), .X(n25356) );
  nor_x1_sg U68947 ( .A(n25358), .B(n42050), .X(n25357) );
  nand_x1_sg U68948 ( .A(n25637), .B(n42049), .X(n25635) );
  nor_x1_sg U68949 ( .A(n25637), .B(n42049), .X(n25636) );
  nand_x1_sg U68950 ( .A(n25914), .B(n42048), .X(n25912) );
  nor_x1_sg U68951 ( .A(n25914), .B(n42048), .X(n25913) );
  nand_x1_sg U68952 ( .A(n26752), .B(n50850), .X(n26750) );
  nor_x1_sg U68953 ( .A(n26752), .B(n50850), .X(n26751) );
  nand_x1_sg U68954 ( .A(n47172), .B(n47170), .X(n23078) );
  nand_x1_sg U68955 ( .A(n23080), .B(n23077), .X(n23079) );
  inv_x1_sg U68956 ( .A(n23080), .X(n47172) );
  nand_x1_sg U68957 ( .A(n47457), .B(n47455), .X(n23358) );
  nand_x1_sg U68958 ( .A(n23360), .B(n23357), .X(n23359) );
  inv_x1_sg U68959 ( .A(n23360), .X(n47457) );
  nand_x1_sg U68960 ( .A(n47742), .B(n47740), .X(n23637) );
  nand_x1_sg U68961 ( .A(n23639), .B(n23636), .X(n23638) );
  inv_x1_sg U68962 ( .A(n23639), .X(n47742) );
  nand_x1_sg U68963 ( .A(n48027), .B(n48025), .X(n23916) );
  nand_x1_sg U68964 ( .A(n23918), .B(n23915), .X(n23917) );
  inv_x1_sg U68965 ( .A(n23918), .X(n48027) );
  nand_x1_sg U68966 ( .A(n48312), .B(n48310), .X(n24195) );
  nand_x1_sg U68967 ( .A(n24197), .B(n24194), .X(n24196) );
  inv_x1_sg U68968 ( .A(n24197), .X(n48312) );
  nand_x1_sg U68969 ( .A(n48597), .B(n48595), .X(n24474) );
  nand_x1_sg U68970 ( .A(n24476), .B(n24473), .X(n24475) );
  inv_x1_sg U68971 ( .A(n24476), .X(n48597) );
  nand_x1_sg U68972 ( .A(n48883), .B(n48881), .X(n24752) );
  nand_x1_sg U68973 ( .A(n24754), .B(n24751), .X(n24753) );
  inv_x1_sg U68974 ( .A(n24754), .X(n48883) );
  nand_x1_sg U68975 ( .A(n49170), .B(n49168), .X(n25031) );
  nand_x1_sg U68976 ( .A(n25033), .B(n25030), .X(n25032) );
  inv_x1_sg U68977 ( .A(n25033), .X(n49170) );
  nand_x1_sg U68978 ( .A(n49456), .B(n49454), .X(n25310) );
  nand_x1_sg U68979 ( .A(n25312), .B(n25309), .X(n25311) );
  inv_x1_sg U68980 ( .A(n25312), .X(n49456) );
  nand_x1_sg U68981 ( .A(n49741), .B(n49739), .X(n25589) );
  nand_x1_sg U68982 ( .A(n25591), .B(n25588), .X(n25590) );
  inv_x1_sg U68983 ( .A(n25591), .X(n49741) );
  nand_x1_sg U68984 ( .A(n50028), .B(n50026), .X(n25866) );
  nand_x1_sg U68985 ( .A(n25868), .B(n25865), .X(n25867) );
  inv_x1_sg U68986 ( .A(n25868), .X(n50028) );
  nand_x1_sg U68987 ( .A(n50602), .B(n50600), .X(n26426) );
  nand_x1_sg U68988 ( .A(n26428), .B(n26425), .X(n26427) );
  inv_x1_sg U68989 ( .A(n26428), .X(n50602) );
  nand_x1_sg U68990 ( .A(n50889), .B(n50887), .X(n26704) );
  nand_x1_sg U68991 ( .A(n26706), .B(n26703), .X(n26705) );
  inv_x1_sg U68992 ( .A(n26706), .X(n50889) );
  nand_x1_sg U68993 ( .A(n22829), .B(n22824), .X(n22828) );
  nor_x1_sg U68994 ( .A(n22829), .B(n22824), .X(n22830) );
  nand_x1_sg U68995 ( .A(n23106), .B(n23102), .X(n23105) );
  nor_x1_sg U68996 ( .A(n23106), .B(n23102), .X(n23107) );
  nand_x1_sg U68997 ( .A(n23386), .B(n23382), .X(n23385) );
  nor_x1_sg U68998 ( .A(n23386), .B(n23382), .X(n23387) );
  nand_x1_sg U68999 ( .A(n23665), .B(n23661), .X(n23664) );
  nor_x1_sg U69000 ( .A(n23665), .B(n23661), .X(n23666) );
  nand_x1_sg U69001 ( .A(n23944), .B(n23940), .X(n23943) );
  nor_x1_sg U69002 ( .A(n23944), .B(n23940), .X(n23945) );
  nand_x1_sg U69003 ( .A(n24223), .B(n24219), .X(n24222) );
  nor_x1_sg U69004 ( .A(n24223), .B(n24219), .X(n24224) );
  nand_x1_sg U69005 ( .A(n24502), .B(n24498), .X(n24501) );
  nor_x1_sg U69006 ( .A(n24502), .B(n24498), .X(n24503) );
  nand_x1_sg U69007 ( .A(n24780), .B(n24776), .X(n24779) );
  nor_x1_sg U69008 ( .A(n24780), .B(n24776), .X(n24781) );
  nand_x1_sg U69009 ( .A(n25059), .B(n25055), .X(n25058) );
  nor_x1_sg U69010 ( .A(n25059), .B(n25055), .X(n25060) );
  nand_x1_sg U69011 ( .A(n25338), .B(n25334), .X(n25337) );
  nor_x1_sg U69012 ( .A(n25338), .B(n25334), .X(n25339) );
  nand_x1_sg U69013 ( .A(n25617), .B(n25613), .X(n25616) );
  nor_x1_sg U69014 ( .A(n25617), .B(n25613), .X(n25618) );
  nand_x1_sg U69015 ( .A(n25894), .B(n25890), .X(n25893) );
  nor_x1_sg U69016 ( .A(n25894), .B(n25890), .X(n25895) );
  nand_x1_sg U69017 ( .A(n26454), .B(n26450), .X(n26453) );
  nor_x1_sg U69018 ( .A(n26454), .B(n26450), .X(n26455) );
  nand_x1_sg U69019 ( .A(n26732), .B(n26728), .X(n26731) );
  nor_x1_sg U69020 ( .A(n26732), .B(n26728), .X(n26733) );
  nand_x1_sg U69021 ( .A(n41660), .B(n39391), .X(n29270) );
  nand_x1_sg U69022 ( .A(n23543), .B(n38942), .X(n23542) );
  nand_x1_sg U69023 ( .A(n26125), .B(n42043), .X(n26123) );
  nor_x1_sg U69024 ( .A(n26125), .B(n42043), .X(n26124) );
  nand_x1_sg U69025 ( .A(n26474), .B(n42047), .X(n26472) );
  nor_x1_sg U69026 ( .A(n26474), .B(n42047), .X(n26473) );
  nand_x1_sg U69027 ( .A(n46879), .B(n46877), .X(n22801) );
  nand_x1_sg U69028 ( .A(n22803), .B(n22800), .X(n22802) );
  inv_x1_sg U69029 ( .A(n22803), .X(n46879) );
  nand_x1_sg U69030 ( .A(n50313), .B(n50311), .X(n26093) );
  nand_x1_sg U69031 ( .A(n26095), .B(n26096), .X(n26094) );
  inv_x1_sg U69032 ( .A(n26095), .X(n50313) );
  nand_x1_sg U69033 ( .A(n26101), .B(n26102), .X(n26099) );
  nor_x1_sg U69034 ( .A(n26101), .B(n26102), .X(n26100) );
  nor_x1_sg U69035 ( .A(n22848), .B(n42046), .X(n22847) );
  nor_x1_sg U69036 ( .A(n40568), .B(n42092), .X(n25920) );
  nor_x1_sg U69037 ( .A(n40314), .B(n6827), .X(n22598) );
  nand_x1_sg U69038 ( .A(n23543), .B(n51136), .X(n28520) );
  nor_x1_sg U69039 ( .A(n40157), .B(n40688), .X(n22858) );
  nor_x1_sg U69040 ( .A(n40358), .B(n40693), .X(n23135) );
  nor_x1_sg U69041 ( .A(n40354), .B(n40698), .X(n23415) );
  nor_x1_sg U69042 ( .A(n40350), .B(n39974), .X(n23694) );
  nor_x1_sg U69043 ( .A(n40346), .B(n39978), .X(n23973) );
  nor_x1_sg U69044 ( .A(n40326), .B(n40713), .X(n24252) );
  nor_x1_sg U69045 ( .A(n40338), .B(n39986), .X(n24531) );
  nor_x1_sg U69046 ( .A(n40334), .B(n39990), .X(n24809) );
  nor_x1_sg U69047 ( .A(n40342), .B(n40728), .X(n25088) );
  nor_x1_sg U69048 ( .A(n40318), .B(n39998), .X(n25367) );
  nor_x1_sg U69049 ( .A(n40322), .B(n40002), .X(n25646) );
  nor_x1_sg U69050 ( .A(n40330), .B(n40006), .X(n26483) );
  nor_x1_sg U69051 ( .A(n40067), .B(n40618), .X(n26187) );
  nand_x1_sg U69052 ( .A(n39479), .B(n12551), .X(\L2_0/n3047 ) );
  nor_x1_sg U69053 ( .A(n28982), .B(n44980), .X(n28817) );
  nor_x1_sg U69054 ( .A(n28985), .B(n28984), .X(n28982) );
  nand_x1_sg U69055 ( .A(n28984), .B(n28985), .X(n28983) );
  nor_x1_sg U69056 ( .A(n28811), .B(n44983), .X(n28629) );
  nor_x1_sg U69057 ( .A(n28814), .B(n28813), .X(n28811) );
  nand_x1_sg U69058 ( .A(n28813), .B(n28814), .X(n28812) );
  nor_x1_sg U69059 ( .A(n28623), .B(n44986), .X(n28468) );
  nor_x1_sg U69060 ( .A(n28626), .B(n28625), .X(n28623) );
  nand_x1_sg U69061 ( .A(n28625), .B(n28626), .X(n28624) );
  nor_x1_sg U69062 ( .A(n28463), .B(n44989), .X(n28374) );
  nor_x1_sg U69063 ( .A(n28462), .B(n28465), .X(n28463) );
  nand_x1_sg U69064 ( .A(n28465), .B(n28462), .X(n28464) );
  nor_x1_sg U69065 ( .A(n28368), .B(n44992), .X(n28261) );
  nor_x1_sg U69066 ( .A(n28371), .B(n28370), .X(n28368) );
  nand_x1_sg U69067 ( .A(n28370), .B(n28371), .X(n28369) );
  nor_x1_sg U69068 ( .A(n27971), .B(n45002), .X(n27808) );
  nor_x1_sg U69069 ( .A(n27974), .B(n27973), .X(n27971) );
  nand_x1_sg U69070 ( .A(n27973), .B(n27974), .X(n27972) );
  nor_x1_sg U69071 ( .A(n27802), .B(n45005), .X(n27622) );
  nor_x1_sg U69072 ( .A(n27805), .B(n27804), .X(n27802) );
  nand_x1_sg U69073 ( .A(n27804), .B(n27805), .X(n27803) );
  nor_x1_sg U69074 ( .A(n27617), .B(n45008), .X(n27419) );
  nor_x1_sg U69075 ( .A(n27616), .B(n27619), .X(n27617) );
  nand_x1_sg U69076 ( .A(n27619), .B(n27616), .X(n27618) );
  nor_x1_sg U69077 ( .A(n27413), .B(n45011), .X(n27197) );
  nor_x1_sg U69078 ( .A(n27416), .B(n27415), .X(n27413) );
  nand_x1_sg U69079 ( .A(n27415), .B(n27416), .X(n27414) );
  nor_x1_sg U69080 ( .A(n27192), .B(n45014), .X(n26958) );
  nor_x1_sg U69081 ( .A(n27191), .B(n27194), .X(n27192) );
  nand_x1_sg U69082 ( .A(n27194), .B(n27191), .X(n27193) );
  nor_x1_sg U69083 ( .A(n29141), .B(n44977), .X(n28988) );
  nor_x1_sg U69084 ( .A(n29140), .B(n29143), .X(n29141) );
  nand_x1_sg U69085 ( .A(n29143), .B(n29140), .X(n29142) );
  nor_x1_sg U69086 ( .A(n28124), .B(n44999), .X(n27977) );
  nor_x1_sg U69087 ( .A(n28127), .B(n28126), .X(n28124) );
  nand_x1_sg U69088 ( .A(n28126), .B(n28127), .X(n28125) );
  nor_x1_sg U69089 ( .A(n21590), .B(n45813), .X(n21437) );
  nor_x1_sg U69090 ( .A(n21589), .B(n21592), .X(n21590) );
  nand_x1_sg U69091 ( .A(n21592), .B(n21589), .X(n21591) );
  nand_x1_sg U69092 ( .A(n39083), .B(n42021), .X(n26778) );
  nor_x1_sg U69093 ( .A(n38559), .B(n22552), .X(n22551) );
  nand_x1_sg U69094 ( .A(n41302), .B(n10913), .X(n42383) );
  nand_x1_sg U69095 ( .A(n23069), .B(n23072), .X(n23071) );
  nor_x1_sg U69096 ( .A(n23072), .B(n23069), .X(n23073) );
  nand_x1_sg U69097 ( .A(n23349), .B(n23352), .X(n23351) );
  nor_x1_sg U69098 ( .A(n23352), .B(n23349), .X(n23353) );
  nand_x1_sg U69099 ( .A(n23628), .B(n23631), .X(n23630) );
  nor_x1_sg U69100 ( .A(n23631), .B(n23628), .X(n23632) );
  nand_x1_sg U69101 ( .A(n23907), .B(n23910), .X(n23909) );
  nor_x1_sg U69102 ( .A(n23910), .B(n23907), .X(n23911) );
  nand_x1_sg U69103 ( .A(n24186), .B(n24189), .X(n24188) );
  nor_x1_sg U69104 ( .A(n24189), .B(n24186), .X(n24190) );
  nand_x1_sg U69105 ( .A(n24465), .B(n24468), .X(n24467) );
  nor_x1_sg U69106 ( .A(n24468), .B(n24465), .X(n24469) );
  nand_x1_sg U69107 ( .A(n24743), .B(n24746), .X(n24745) );
  nor_x1_sg U69108 ( .A(n24746), .B(n24743), .X(n24747) );
  nand_x1_sg U69109 ( .A(n25022), .B(n25025), .X(n25024) );
  nor_x1_sg U69110 ( .A(n25025), .B(n25022), .X(n25026) );
  nand_x1_sg U69111 ( .A(n25301), .B(n25304), .X(n25303) );
  nor_x1_sg U69112 ( .A(n25304), .B(n25301), .X(n25305) );
  nand_x1_sg U69113 ( .A(n25580), .B(n25583), .X(n25582) );
  nor_x1_sg U69114 ( .A(n25583), .B(n25580), .X(n25584) );
  nand_x1_sg U69115 ( .A(n25857), .B(n25860), .X(n25859) );
  nor_x1_sg U69116 ( .A(n25860), .B(n25857), .X(n25861) );
  nand_x1_sg U69117 ( .A(n26417), .B(n26420), .X(n26419) );
  nor_x1_sg U69118 ( .A(n26420), .B(n26417), .X(n26421) );
  nand_x1_sg U69119 ( .A(n26695), .B(n26698), .X(n26697) );
  nor_x1_sg U69120 ( .A(n26698), .B(n26695), .X(n26699) );
  nor_x1_sg U69121 ( .A(n22812), .B(n42146), .X(n22810) );
  nor_x1_sg U69122 ( .A(n23089), .B(n42145), .X(n23087) );
  nor_x1_sg U69123 ( .A(n23369), .B(n42144), .X(n23367) );
  nor_x1_sg U69124 ( .A(n23648), .B(n42143), .X(n23646) );
  nor_x1_sg U69125 ( .A(n23927), .B(n42142), .X(n23925) );
  nor_x1_sg U69126 ( .A(n24206), .B(n42141), .X(n24204) );
  nor_x1_sg U69127 ( .A(n24485), .B(n42140), .X(n24483) );
  nor_x1_sg U69128 ( .A(n24763), .B(n42139), .X(n24761) );
  nor_x1_sg U69129 ( .A(n25042), .B(n42138), .X(n25040) );
  nor_x1_sg U69130 ( .A(n25321), .B(n42137), .X(n25319) );
  nor_x1_sg U69131 ( .A(n25600), .B(n42060), .X(n25598) );
  nor_x1_sg U69132 ( .A(n25877), .B(n42136), .X(n25875) );
  nor_x1_sg U69133 ( .A(n26437), .B(n42135), .X(n26435) );
  nor_x1_sg U69134 ( .A(n26715), .B(n42134), .X(n26713) );
  nor_x1_sg U69135 ( .A(n22988), .B(n22987), .X(n22985) );
  nor_x1_sg U69136 ( .A(n23268), .B(n23267), .X(n23265) );
  nor_x1_sg U69137 ( .A(n23547), .B(n23546), .X(n23544) );
  nor_x1_sg U69138 ( .A(n23826), .B(n23825), .X(n23823) );
  nor_x1_sg U69139 ( .A(n24105), .B(n24104), .X(n24102) );
  nor_x1_sg U69140 ( .A(n24384), .B(n24383), .X(n24381) );
  nor_x1_sg U69141 ( .A(n24662), .B(n24661), .X(n24659) );
  nor_x1_sg U69142 ( .A(n24941), .B(n24940), .X(n24938) );
  nor_x1_sg U69143 ( .A(n25220), .B(n25219), .X(n25217) );
  nor_x1_sg U69144 ( .A(n25499), .B(n25498), .X(n25496) );
  nor_x1_sg U69145 ( .A(n25776), .B(n25775), .X(n25773) );
  nor_x1_sg U69146 ( .A(n26336), .B(n26335), .X(n26333) );
  nor_x1_sg U69147 ( .A(n26614), .B(n26613), .X(n26611) );
  nor_x1_sg U69148 ( .A(n38176), .B(n44993), .X(n28259) );
  nor_x1_sg U69149 ( .A(n38168), .B(n44996), .X(n28128) );
  nor_x1_sg U69150 ( .A(n38177), .B(n45000), .X(n27975) );
  nor_x1_sg U69151 ( .A(n38178), .B(n45003), .X(n27806) );
  nor_x1_sg U69152 ( .A(n38179), .B(n45006), .X(n27620) );
  nor_x1_sg U69153 ( .A(n38180), .B(n44984), .X(n28627) );
  nor_x1_sg U69154 ( .A(n38181), .B(n45009), .X(n27417) );
  nor_x1_sg U69155 ( .A(n38182), .B(n45814), .X(n21435) );
  nor_x1_sg U69156 ( .A(n38183), .B(n44987), .X(n28466) );
  nor_x1_sg U69157 ( .A(n38184), .B(n44978), .X(n28986) );
  nor_x1_sg U69158 ( .A(n38185), .B(n45012), .X(n27195) );
  nor_x1_sg U69159 ( .A(n38186), .B(n44990), .X(n28372) );
  nor_x1_sg U69160 ( .A(n38187), .B(n44981), .X(n28815) );
  nor_x1_sg U69161 ( .A(n38188), .B(n45015), .X(n26956) );
  nor_x1_sg U69162 ( .A(n38148), .B(n45821), .X(n21073) );
  nor_x1_sg U69163 ( .A(n38173), .B(n45825), .X(n20847) );
  nor_x1_sg U69164 ( .A(n38149), .B(n45829), .X(n20665) );
  nor_x1_sg U69165 ( .A(n38169), .B(n45833), .X(n20494) );
  nor_x1_sg U69166 ( .A(n38150), .B(n45837), .X(n20364) );
  nor_x1_sg U69167 ( .A(n38174), .B(n45841), .X(n20204) );
  nor_x1_sg U69168 ( .A(n38151), .B(n45845), .X(n20025) );
  nor_x1_sg U69169 ( .A(n38170), .B(n45849), .X(n19837) );
  nor_x1_sg U69170 ( .A(n38152), .B(n45853), .X(n19631) );
  nor_x1_sg U69171 ( .A(n38175), .B(n45857), .X(n19398) );
  nor_x1_sg U69172 ( .A(n38171), .B(n45817), .X(n21263) );
  nor_x1_sg U69173 ( .A(n38153), .B(n45861), .X(n19221) );
  nor_x1_sg U69174 ( .A(n38172), .B(n45865), .X(n6759) );
  nand_x1_sg U69175 ( .A(n20954), .B(n38693), .X(n20952) );
  nor_x1_sg U69176 ( .A(n6055), .B(n20954), .X(n20953) );
  nand_x1_sg U69177 ( .A(n40099), .B(n39479), .X(n29273) );
  nor_x1_sg U69178 ( .A(n23115), .B(n23111), .X(n23114) );
  nor_x1_sg U69179 ( .A(n23395), .B(n23391), .X(n23394) );
  nor_x1_sg U69180 ( .A(n23674), .B(n23670), .X(n23673) );
  nor_x1_sg U69181 ( .A(n23953), .B(n23949), .X(n23952) );
  nor_x1_sg U69182 ( .A(n24232), .B(n24228), .X(n24231) );
  nor_x1_sg U69183 ( .A(n24511), .B(n24507), .X(n24510) );
  nor_x1_sg U69184 ( .A(n24789), .B(n24785), .X(n24788) );
  nor_x1_sg U69185 ( .A(n25068), .B(n25064), .X(n25067) );
  nor_x1_sg U69186 ( .A(n25347), .B(n25343), .X(n25346) );
  nor_x1_sg U69187 ( .A(n25626), .B(n25622), .X(n25625) );
  nor_x1_sg U69188 ( .A(n25903), .B(n25899), .X(n25902) );
  nor_x1_sg U69189 ( .A(n26463), .B(n26459), .X(n26462) );
  nor_x1_sg U69190 ( .A(n26741), .B(n26737), .X(n26740) );
  nor_x1_sg U69191 ( .A(n22838), .B(n22834), .X(n22837) );
  nor_x1_sg U69192 ( .A(n26112), .B(n26113), .X(n26111) );
  nor_x1_sg U69193 ( .A(n41951), .B(n44976), .X(n29143) );
  inv_x1_sg U69194 ( .A(n29145), .X(n44976) );
  nor_x1_sg U69195 ( .A(n41952), .B(n45812), .X(n21592) );
  inv_x1_sg U69196 ( .A(n21594), .X(n45812) );
  nor_x1_sg U69197 ( .A(n21719), .B(n41287), .X(n5951) );
  nor_x1_sg U69198 ( .A(n40583), .B(n51136), .X(n21719) );
  inv_x1_sg U69199 ( .A(n23120), .X(n47134) );
  inv_x1_sg U69200 ( .A(n26746), .X(n50850) );
  nand_x1_sg U69201 ( .A(n50522), .B(n26132), .X(n26148) );
  nand_x1_sg U69202 ( .A(n20106), .B(n6211), .X(n20104) );
  nor_x1_sg U69203 ( .A(n6211), .B(n20106), .X(n20105) );
  nand_x1_sg U69204 ( .A(n19701), .B(n38638), .X(n19699) );
  nor_x1_sg U69205 ( .A(n6207), .B(n19701), .X(n19700) );
  nand_x1_sg U69206 ( .A(n20780), .B(n38703), .X(n20778) );
  nor_x1_sg U69207 ( .A(n42335), .B(n20780), .X(n20779) );
  nand_x1_sg U69208 ( .A(n46470), .B(n46452), .X(n20300) );
  nand_x1_sg U69209 ( .A(n20301), .B(n6147), .X(n20299) );
  nand_x1_sg U69210 ( .A(n20100), .B(n20103), .X(n20162) );
  nand_x1_sg U69211 ( .A(n46307), .B(n42213), .X(n20164) );
  nand_x1_sg U69212 ( .A(n46391), .B(n42024), .X(n19582) );
  nand_x1_sg U69213 ( .A(n41545), .B(n6084), .X(n19157) );
  nand_x1_sg U69214 ( .A(n46480), .B(n6077), .X(n19159) );
  nand_x1_sg U69215 ( .A(n20852), .B(n42229), .X(n20849) );
  nand_x1_sg U69216 ( .A(n20851), .B(n45827), .X(n20850) );
  nand_x1_sg U69217 ( .A(n20209), .B(n42227), .X(n20206) );
  nand_x1_sg U69218 ( .A(n20208), .B(n45843), .X(n20207) );
  nand_x1_sg U69219 ( .A(n19713), .B(n42262), .X(n19710) );
  nand_x1_sg U69220 ( .A(n19712), .B(n46444), .X(n19711) );
  nand_x1_sg U69221 ( .A(n19403), .B(n42225), .X(n19400) );
  nand_x1_sg U69222 ( .A(n19402), .B(n45859), .X(n19401) );
  nand_x1_sg U69223 ( .A(n28264), .B(n45035), .X(n28262) );
  nor_x1_sg U69224 ( .A(n45035), .B(n28264), .X(n28263) );
  nand_x1_sg U69225 ( .A(n46385), .B(n46341), .X(n19166) );
  nand_x1_sg U69226 ( .A(n6223), .B(n6216), .X(n19168) );
  nand_x1_sg U69227 ( .A(n21268), .B(n45875), .X(n21265) );
  nand_x1_sg U69228 ( .A(n21267), .B(n45819), .X(n21266) );
  nand_x1_sg U69229 ( .A(n20440), .B(n46424), .X(n20438) );
  nand_x1_sg U69230 ( .A(n20310), .B(n46379), .X(n20439) );
  nand_x1_sg U69231 ( .A(n20499), .B(n45878), .X(n20496) );
  nand_x1_sg U69232 ( .A(n20498), .B(n45835), .X(n20497) );
  nand_x1_sg U69233 ( .A(n19842), .B(n45881), .X(n19839) );
  nand_x1_sg U69234 ( .A(n19841), .B(n45851), .X(n19840) );
  nand_x1_sg U69235 ( .A(n19224), .B(n19225), .X(n19223) );
  nor_x1_sg U69236 ( .A(n19225), .B(n19224), .X(n19226) );
  nor_x1_sg U69237 ( .A(n23543), .B(n51181), .X(n20961) );
  nand_x1_sg U69238 ( .A(n47360), .B(n22998), .X(n22997) );
  nand_x1_sg U69239 ( .A(n47645), .B(n23278), .X(n23277) );
  nand_x1_sg U69240 ( .A(n47930), .B(n23557), .X(n23556) );
  nand_x1_sg U69241 ( .A(n48215), .B(n23836), .X(n23835) );
  nand_x1_sg U69242 ( .A(n48500), .B(n24115), .X(n24114) );
  nand_x1_sg U69243 ( .A(n48785), .B(n24394), .X(n24393) );
  nand_x1_sg U69244 ( .A(n49072), .B(n24672), .X(n24671) );
  nand_x1_sg U69245 ( .A(n49358), .B(n24951), .X(n24950) );
  nand_x1_sg U69246 ( .A(n49644), .B(n25230), .X(n25229) );
  nand_x1_sg U69247 ( .A(n49930), .B(n25509), .X(n25508) );
  nand_x1_sg U69248 ( .A(n50216), .B(n25786), .X(n25785) );
  nand_x1_sg U69249 ( .A(n50790), .B(n26346), .X(n26345) );
  nand_x1_sg U69250 ( .A(n51077), .B(n26624), .X(n26623) );
  nand_x1_sg U69251 ( .A(n46423), .B(n46404), .X(n20442) );
  nand_x1_sg U69252 ( .A(n20443), .B(n6193), .X(n20441) );
  nand_x1_sg U69253 ( .A(n21440), .B(n45873), .X(n21438) );
  nor_x1_sg U69254 ( .A(n45873), .B(n21440), .X(n21439) );
  nand_x1_sg U69255 ( .A(n20668), .B(n20669), .X(n20667) );
  nor_x1_sg U69256 ( .A(n20669), .B(n20668), .X(n20670) );
  nand_x1_sg U69257 ( .A(n20028), .B(n20029), .X(n20027) );
  nor_x1_sg U69258 ( .A(n20029), .B(n20028), .X(n20030) );
  nand_x1_sg U69259 ( .A(n20768), .B(n20771), .X(n20793) );
  nand_x1_sg U69260 ( .A(n46491), .B(n42259), .X(n20795) );
  nand_x1_sg U69261 ( .A(n19470), .B(n19474), .X(n19587) );
  nand_x1_sg U69262 ( .A(n46300), .B(n46339), .X(n19589) );
  nand_x1_sg U69263 ( .A(n46507), .B(n46489), .X(n20598) );
  nand_x1_sg U69264 ( .A(n20136), .B(n6101), .X(n20600) );
  nand_x1_sg U69265 ( .A(n20452), .B(n38575), .X(n20451) );
  nor_x1_sg U69266 ( .A(n6285), .B(n20431), .X(n20453) );
  nand_x1_sg U69267 ( .A(n42020), .B(n26792), .X(n24380) );
  nand_x1_sg U69268 ( .A(n39083), .B(n39391), .X(n26792) );
  nor_x1_sg U69269 ( .A(n6807), .B(n41076), .X(n6806) );
  nand_x1_sg U69270 ( .A(n47074), .B(n22721), .X(n22720) );
  nand_x1_sg U69271 ( .A(n22566), .B(n38127), .X(n27191) );
  nor_x1_sg U69272 ( .A(n6794), .B(n41006), .X(n6793) );
  nor_x1_sg U69273 ( .A(n6797), .B(n41029), .X(n6796) );
  nor_x1_sg U69274 ( .A(n6818), .B(n42332), .X(n6817) );
  nor_x1_sg U69275 ( .A(n6821), .B(n41016), .X(n6820) );
  nor_x1_sg U69276 ( .A(n28920), .B(n38126), .X(n28919) );
  nand_x1_sg U69277 ( .A(n47056), .B(n22729), .X(n22728) );
  nand_x1_sg U69278 ( .A(n47342), .B(n23006), .X(n23005) );
  nand_x1_sg U69279 ( .A(n47627), .B(n23286), .X(n23285) );
  nand_x1_sg U69280 ( .A(n47912), .B(n23565), .X(n23564) );
  nand_x1_sg U69281 ( .A(n48197), .B(n23844), .X(n23843) );
  nand_x1_sg U69282 ( .A(n48482), .B(n24123), .X(n24122) );
  nand_x1_sg U69283 ( .A(n48767), .B(n24402), .X(n24401) );
  nand_x1_sg U69284 ( .A(n49053), .B(n24680), .X(n24679) );
  nand_x1_sg U69285 ( .A(n49340), .B(n24959), .X(n24958) );
  nand_x1_sg U69286 ( .A(n49626), .B(n25238), .X(n25237) );
  nand_x1_sg U69287 ( .A(n49912), .B(n25517), .X(n25516) );
  nand_x1_sg U69288 ( .A(n50198), .B(n25794), .X(n25793) );
  nand_x1_sg U69289 ( .A(n50500), .B(n26138), .X(n26149) );
  nand_x1_sg U69290 ( .A(n50772), .B(n26354), .X(n26353) );
  nand_x1_sg U69291 ( .A(n51059), .B(n26632), .X(n26631) );
  nand_x1_sg U69292 ( .A(n21531), .B(n46503), .X(n21529) );
  nor_x1_sg U69293 ( .A(n46503), .B(n21531), .X(n21530) );
  nand_x1_sg U69294 ( .A(n21349), .B(n46545), .X(n21347) );
  nor_x1_sg U69295 ( .A(n46545), .B(n21349), .X(n21348) );
  nor_x1_sg U69296 ( .A(n6802), .B(n41252), .X(n6801) );
  nand_x1_sg U69297 ( .A(n20288), .B(n20289), .X(n20287) );
  nor_x1_sg U69298 ( .A(n20289), .B(n20288), .X(n20290) );
  nand_x1_sg U69299 ( .A(n46567), .B(n19724), .X(n19723) );
  nor_x1_sg U69300 ( .A(n19724), .B(n46567), .X(n19725) );
  nand_x1_sg U69301 ( .A(n46518), .B(n19918), .X(n19917) );
  nor_x1_sg U69302 ( .A(n19918), .B(n46518), .X(n19919) );
  nor_x1_sg U69303 ( .A(n38121), .B(n29197), .X(n29241) );
  nor_x1_sg U69304 ( .A(n38122), .B(n29209), .X(n29235) );
  nor_x1_sg U69305 ( .A(n38124), .B(n29221), .X(n29229) );
  nor_x1_sg U69306 ( .A(n38125), .B(n21356), .X(n21355) );
  nor_x1_sg U69307 ( .A(n38123), .B(n21670), .X(n21678) );
  nand_x1_sg U69308 ( .A(n45923), .B(n45910), .X(n20857) );
  nand_x1_sg U69309 ( .A(n20858), .B(n6691), .X(n20856) );
  nand_x1_sg U69310 ( .A(n45926), .B(n45900), .X(n20214) );
  nand_x1_sg U69311 ( .A(n20215), .B(n6659), .X(n20213) );
  nand_x1_sg U69312 ( .A(n45929), .B(n45890), .X(n19408) );
  nand_x1_sg U69313 ( .A(n19409), .B(n6674), .X(n19407) );
  nand_x1_sg U69314 ( .A(n46479), .B(n19314), .X(n19313) );
  nand_x1_sg U69315 ( .A(n46439), .B(n6134), .X(n19312) );
  inv_x1_sg U69316 ( .A(n19314), .X(n46439) );
  nand_x1_sg U69317 ( .A(n20660), .B(n38141), .X(n20664) );
  nand_x1_sg U69318 ( .A(n20020), .B(n38143), .X(n20024) );
  nand_x1_sg U69319 ( .A(n20359), .B(n38142), .X(n20363) );
  nand_x1_sg U69320 ( .A(n19626), .B(n38144), .X(n19630) );
  nand_x1_sg U69321 ( .A(n19216), .B(n38146), .X(n19220) );
  nand_x1_sg U69322 ( .A(n21068), .B(n38145), .X(n21072) );
  nand_x1_sg U69323 ( .A(n28123), .B(n38147), .X(n28127) );
  nand_x1_sg U69324 ( .A(n23069), .B(n23070), .X(n23068) );
  nand_x1_sg U69325 ( .A(n23349), .B(n23350), .X(n23348) );
  nand_x1_sg U69326 ( .A(n23628), .B(n23629), .X(n23627) );
  nand_x1_sg U69327 ( .A(n23907), .B(n23908), .X(n23906) );
  nand_x1_sg U69328 ( .A(n24186), .B(n24187), .X(n24185) );
  nand_x1_sg U69329 ( .A(n24465), .B(n24466), .X(n24464) );
  nand_x1_sg U69330 ( .A(n24743), .B(n24744), .X(n24742) );
  nand_x1_sg U69331 ( .A(n25022), .B(n25023), .X(n25021) );
  nand_x1_sg U69332 ( .A(n25301), .B(n25302), .X(n25300) );
  nand_x1_sg U69333 ( .A(n25580), .B(n25581), .X(n25579) );
  nand_x1_sg U69334 ( .A(n25857), .B(n25858), .X(n25856) );
  nand_x1_sg U69335 ( .A(n26089), .B(n26091), .X(n26158) );
  nand_x1_sg U69336 ( .A(n26417), .B(n26418), .X(n26416) );
  nand_x1_sg U69337 ( .A(n26695), .B(n26696), .X(n26694) );
  nand_x1_sg U69338 ( .A(n22792), .B(n22793), .X(n22791) );
  inv_x1_sg U69339 ( .A(n6821), .X(n45801) );
  inv_x1_sg U69340 ( .A(n6818), .X(n45803) );
  inv_x1_sg U69341 ( .A(n6797), .X(n45805) );
  inv_x1_sg U69342 ( .A(n6794), .X(n45807) );
  inv_x1_sg U69343 ( .A(n6807), .X(n45809) );
  nand_x1_sg U69344 ( .A(n19913), .B(n42226), .X(n19910) );
  nand_x1_sg U69345 ( .A(n19912), .B(n46446), .X(n19911) );
  nand_x1_sg U69346 ( .A(n20927), .B(n46374), .X(n20924) );
  nand_x1_sg U69347 ( .A(n20926), .B(n46361), .X(n20925) );
  nand_x1_sg U69348 ( .A(n20920), .B(n46333), .X(n20917) );
  nand_x1_sg U69349 ( .A(n20919), .B(n46319), .X(n20918) );
  nand_x1_sg U69350 ( .A(n20913), .B(n46287), .X(n20910) );
  nand_x1_sg U69351 ( .A(n20912), .B(n46274), .X(n20911) );
  nand_x1_sg U69352 ( .A(n20906), .B(n46242), .X(n20903) );
  nand_x1_sg U69353 ( .A(n20905), .B(n46228), .X(n20904) );
  nand_x1_sg U69354 ( .A(n20899), .B(n46196), .X(n20896) );
  nand_x1_sg U69355 ( .A(n20898), .B(n46183), .X(n20897) );
  nand_x1_sg U69356 ( .A(n20892), .B(n46151), .X(n20889) );
  nand_x1_sg U69357 ( .A(n20891), .B(n46137), .X(n20890) );
  nand_x1_sg U69358 ( .A(n20885), .B(n46105), .X(n20882) );
  nand_x1_sg U69359 ( .A(n20884), .B(n46092), .X(n20883) );
  nand_x1_sg U69360 ( .A(n20878), .B(n46060), .X(n20875) );
  nand_x1_sg U69361 ( .A(n20877), .B(n46046), .X(n20876) );
  nand_x1_sg U69362 ( .A(n20871), .B(n46014), .X(n20868) );
  nand_x1_sg U69363 ( .A(n20870), .B(n46001), .X(n20869) );
  nand_x1_sg U69364 ( .A(n20864), .B(n45969), .X(n20861) );
  nand_x1_sg U69365 ( .A(n20863), .B(n45956), .X(n20862) );
  nand_x1_sg U69366 ( .A(n20934), .B(n46422), .X(n20931) );
  nand_x1_sg U69367 ( .A(n20933), .B(n46408), .X(n20932) );
  nand_x1_sg U69368 ( .A(n20941), .B(n46469), .X(n20938) );
  nand_x1_sg U69369 ( .A(n20940), .B(n46456), .X(n20939) );
  nand_x1_sg U69370 ( .A(n20948), .B(n46506), .X(n20945) );
  nand_x1_sg U69371 ( .A(n20947), .B(n46494), .X(n20946) );
  nand_x1_sg U69372 ( .A(n20277), .B(n46336), .X(n20274) );
  nand_x1_sg U69373 ( .A(n20276), .B(n46310), .X(n20275) );
  nand_x1_sg U69374 ( .A(n20270), .B(n46290), .X(n20267) );
  nand_x1_sg U69375 ( .A(n20269), .B(n46265), .X(n20268) );
  nand_x1_sg U69376 ( .A(n20263), .B(n46245), .X(n20260) );
  nand_x1_sg U69377 ( .A(n20262), .B(n46219), .X(n20261) );
  nand_x1_sg U69378 ( .A(n20256), .B(n46199), .X(n20253) );
  nand_x1_sg U69379 ( .A(n20255), .B(n46174), .X(n20254) );
  nand_x1_sg U69380 ( .A(n20249), .B(n46154), .X(n20246) );
  nand_x1_sg U69381 ( .A(n20248), .B(n46128), .X(n20247) );
  nand_x1_sg U69382 ( .A(n20242), .B(n46108), .X(n20239) );
  nand_x1_sg U69383 ( .A(n20241), .B(n46083), .X(n20240) );
  nand_x1_sg U69384 ( .A(n20235), .B(n46063), .X(n20232) );
  nand_x1_sg U69385 ( .A(n20234), .B(n46037), .X(n20233) );
  nand_x1_sg U69386 ( .A(n20228), .B(n46017), .X(n20225) );
  nand_x1_sg U69387 ( .A(n20227), .B(n45992), .X(n20226) );
  nand_x1_sg U69388 ( .A(n20221), .B(n45972), .X(n20218) );
  nand_x1_sg U69389 ( .A(n20220), .B(n45947), .X(n20219) );
  nand_x1_sg U69390 ( .A(n28318), .B(n45442), .X(n28316) );
  nor_x1_sg U69391 ( .A(n45442), .B(n28318), .X(n28317) );
  nand_x1_sg U69392 ( .A(n28189), .B(n45487), .X(n28187) );
  nor_x1_sg U69393 ( .A(n45487), .B(n28189), .X(n28188) );
  nand_x1_sg U69394 ( .A(n28054), .B(n45531), .X(n28052) );
  nor_x1_sg U69395 ( .A(n45531), .B(n28054), .X(n28053) );
  nand_x1_sg U69396 ( .A(n27892), .B(n45576), .X(n27890) );
  nor_x1_sg U69397 ( .A(n45576), .B(n27892), .X(n27891) );
  nand_x1_sg U69398 ( .A(n27715), .B(n45620), .X(n27713) );
  nor_x1_sg U69399 ( .A(n45620), .B(n27715), .X(n27714) );
  nand_x1_sg U69400 ( .A(n27521), .B(n45664), .X(n27519) );
  nor_x1_sg U69401 ( .A(n45664), .B(n27521), .X(n27520) );
  nand_x1_sg U69402 ( .A(n27308), .B(n45708), .X(n27306) );
  nor_x1_sg U69403 ( .A(n45708), .B(n27308), .X(n27307) );
  nand_x1_sg U69404 ( .A(n21179), .B(n46585), .X(n21177) );
  nor_x1_sg U69405 ( .A(n46585), .B(n21179), .X(n21178) );
  nand_x1_sg U69406 ( .A(n19471), .B(n46339), .X(n19468) );
  nand_x1_sg U69407 ( .A(n19470), .B(n46301), .X(n19469) );
  nand_x1_sg U69408 ( .A(n19464), .B(n46293), .X(n19461) );
  nand_x1_sg U69409 ( .A(n19463), .B(n46256), .X(n19462) );
  nand_x1_sg U69410 ( .A(n19457), .B(n46248), .X(n19454) );
  nand_x1_sg U69411 ( .A(n19456), .B(n46210), .X(n19455) );
  nand_x1_sg U69412 ( .A(n19450), .B(n46202), .X(n19447) );
  nand_x1_sg U69413 ( .A(n19449), .B(n46165), .X(n19448) );
  nand_x1_sg U69414 ( .A(n19443), .B(n46157), .X(n19440) );
  nand_x1_sg U69415 ( .A(n19442), .B(n46119), .X(n19441) );
  nand_x1_sg U69416 ( .A(n19436), .B(n46111), .X(n19433) );
  nand_x1_sg U69417 ( .A(n19435), .B(n46074), .X(n19434) );
  nand_x1_sg U69418 ( .A(n19429), .B(n46066), .X(n19426) );
  nand_x1_sg U69419 ( .A(n19428), .B(n46028), .X(n19427) );
  nand_x1_sg U69420 ( .A(n19422), .B(n46020), .X(n19419) );
  nand_x1_sg U69421 ( .A(n19421), .B(n45983), .X(n19420) );
  nand_x1_sg U69422 ( .A(n19415), .B(n45975), .X(n19412) );
  nand_x1_sg U69423 ( .A(n19414), .B(n45938), .X(n19413) );
  nand_x1_sg U69424 ( .A(n41548), .B(n46396), .X(n19967) );
  nand_x1_sg U69425 ( .A(n19969), .B(n38194), .X(n19968) );
  nand_x1_sg U69426 ( .A(n41546), .B(n46483), .X(n19574) );
  nand_x1_sg U69427 ( .A(n19576), .B(n38195), .X(n19575) );
  nand_x1_sg U69428 ( .A(n20147), .B(n38596), .X(n20146) );
  nor_x1_sg U69429 ( .A(n6118), .B(n20148), .X(n20149) );
  nand_x1_sg U69430 ( .A(n19955), .B(n38594), .X(n19954) );
  nor_x1_sg U69431 ( .A(n42331), .B(n19956), .X(n19957) );
  nand_x1_sg U69432 ( .A(n21076), .B(n21077), .X(n21075) );
  nor_x1_sg U69433 ( .A(n21077), .B(n21076), .X(n21078) );
  nand_x1_sg U69434 ( .A(n20367), .B(n20368), .X(n20366) );
  nor_x1_sg U69435 ( .A(n20368), .B(n20367), .X(n20369) );
  nand_x1_sg U69436 ( .A(n46476), .B(n20118), .X(n20117) );
  nor_x1_sg U69437 ( .A(n20118), .B(n46476), .X(n20119) );
  nand_x1_sg U69438 ( .A(n19634), .B(n19635), .X(n19633) );
  nor_x1_sg U69439 ( .A(n19635), .B(n19634), .X(n19636) );
  inv_x1_sg U69440 ( .A(n21430), .X(n45798) );
  inv_x1_sg U69441 ( .A(n28981), .X(n44964) );
  nor_x1_sg U69442 ( .A(n19746), .B(n19748), .X(n20594) );
  nor_x1_sg U69443 ( .A(n20673), .B(n20668), .X(n20837) );
  nor_x1_sg U69444 ( .A(n20033), .B(n20028), .X(n20194) );
  nor_x1_sg U69445 ( .A(n19229), .B(n19224), .X(n19388) );
  nor_x1_sg U69446 ( .A(n21081), .B(n21076), .X(n21252) );
  nor_x1_sg U69447 ( .A(n20372), .B(n20367), .X(n20484) );
  nor_x1_sg U69448 ( .A(n19639), .B(n19634), .X(n19827) );
  nand_x1_sg U69449 ( .A(n7300), .B(n40316), .X(n7299) );
  nand_x1_sg U69450 ( .A(n42161), .B(n40688), .X(n8117) );
  nand_x1_sg U69451 ( .A(n8936), .B(n40691), .X(n8935) );
  nand_x1_sg U69452 ( .A(n9756), .B(n40696), .X(n9755) );
  nand_x1_sg U69453 ( .A(n10575), .B(n40703), .X(n10574) );
  nand_x1_sg U69454 ( .A(n11394), .B(n40706), .X(n11393) );
  nand_x1_sg U69455 ( .A(n12213), .B(n40714), .X(n12212) );
  nand_x1_sg U69456 ( .A(n13032), .B(n40718), .X(n13031) );
  nand_x1_sg U69457 ( .A(n13851), .B(n40721), .X(n13850) );
  nand_x1_sg U69458 ( .A(n14670), .B(n40728), .X(n14669) );
  nand_x1_sg U69459 ( .A(n42160), .B(n40731), .X(n15488) );
  nand_x1_sg U69460 ( .A(n16308), .B(n40736), .X(n16307) );
  nand_x1_sg U69461 ( .A(n17125), .B(n40571), .X(n17124) );
  nand_x1_sg U69462 ( .A(n41670), .B(n42044), .X(n17945) );
  nand_x1_sg U69463 ( .A(n18767), .B(n40743), .X(n18766) );
  nor_x1_sg U69464 ( .A(n6171), .B(n46433), .X(n6170) );
  nor_x1_sg U69465 ( .A(n6173), .B(n6169), .X(n6171) );
  nand_x1_sg U69466 ( .A(n6169), .B(n6173), .X(n6172) );
  nand_x1_sg U69467 ( .A(n39677), .B(n40687), .X(n8419) );
  nand_x1_sg U69468 ( .A(n39676), .B(n40692), .X(n9237) );
  nand_x1_sg U69469 ( .A(n39674), .B(n40697), .X(n10057) );
  nand_x1_sg U69470 ( .A(n39675), .B(n40704), .X(n10876) );
  nand_x1_sg U69471 ( .A(n39673), .B(n40709), .X(n11695) );
  nand_x1_sg U69472 ( .A(n39672), .B(n40712), .X(n12514) );
  nand_x1_sg U69473 ( .A(n39670), .B(n40719), .X(n13333) );
  nand_x1_sg U69474 ( .A(n39671), .B(n40724), .X(n14152) );
  nand_x1_sg U69475 ( .A(n39669), .B(n40727), .X(n14971) );
  nand_x1_sg U69476 ( .A(n39668), .B(n40731), .X(n15790) );
  nand_x1_sg U69477 ( .A(n39666), .B(n40739), .X(n16609) );
  nand_x1_sg U69478 ( .A(n39667), .B(n40617), .X(n18247) );
  nand_x1_sg U69479 ( .A(n39665), .B(n40743), .X(n19068) );
  nand_x1_sg U69480 ( .A(n39798), .B(n40686), .X(n8261) );
  nand_x1_sg U69481 ( .A(n39800), .B(n40691), .X(n9079) );
  nand_x1_sg U69482 ( .A(n39794), .B(n40698), .X(n9899) );
  nand_x1_sg U69483 ( .A(n39796), .B(n40703), .X(n10718) );
  nand_x1_sg U69484 ( .A(n39790), .B(n40707), .X(n11537) );
  nand_x1_sg U69485 ( .A(n39792), .B(n40712), .X(n12356) );
  nand_x1_sg U69486 ( .A(n39786), .B(n40718), .X(n13175) );
  nand_x1_sg U69487 ( .A(n39788), .B(n40722), .X(n13994) );
  nand_x1_sg U69488 ( .A(n39782), .B(n40727), .X(n14813) );
  nand_x1_sg U69489 ( .A(n39784), .B(n40734), .X(n15632) );
  nand_x1_sg U69490 ( .A(n39778), .B(n40737), .X(n16451) );
  nand_x1_sg U69491 ( .A(n39780), .B(n40619), .X(n18089) );
  nand_x1_sg U69492 ( .A(n39776), .B(n40741), .X(n18910) );
  nand_x1_sg U69493 ( .A(n39563), .B(n40687), .X(n8004) );
  nand_x1_sg U69494 ( .A(n39566), .B(n40691), .X(n8822) );
  nand_x1_sg U69495 ( .A(n39569), .B(n40697), .X(n9642) );
  nand_x1_sg U69496 ( .A(n39572), .B(n40704), .X(n10461) );
  nand_x1_sg U69497 ( .A(n39575), .B(n40707), .X(n11280) );
  nand_x1_sg U69498 ( .A(n39578), .B(n40713), .X(n12099) );
  nand_x1_sg U69499 ( .A(n39581), .B(n40716), .X(n12918) );
  nand_x1_sg U69500 ( .A(n39584), .B(n40722), .X(n13737) );
  nand_x1_sg U69501 ( .A(n39587), .B(n40729), .X(n14556) );
  nand_x1_sg U69502 ( .A(n39590), .B(n40733), .X(n15375) );
  nand_x1_sg U69503 ( .A(n39593), .B(n40737), .X(n16194) );
  nand_x1_sg U69504 ( .A(n39599), .B(n40617), .X(n17832) );
  nand_x1_sg U69505 ( .A(n39596), .B(n40741), .X(n18653) );
  nand_x1_sg U69506 ( .A(n39560), .B(n40571), .X(n17010) );
  nor_x1_sg U69507 ( .A(n20309), .B(n20310), .X(n20308) );
  nor_x1_sg U69508 ( .A(n20142), .B(n20143), .X(n20141) );
  nor_x1_sg U69509 ( .A(n19944), .B(n46508), .X(n19943) );
  nor_x1_sg U69510 ( .A(n5978), .B(n46609), .X(n5976) );
  nor_x1_sg U69511 ( .A(n5980), .B(n38669), .X(n5978) );
  nand_x1_sg U69512 ( .A(n5974), .B(n5980), .X(n5979) );
  nor_x1_sg U69513 ( .A(n6079), .B(n46522), .X(n6078) );
  nor_x1_sg U69514 ( .A(n6081), .B(n38667), .X(n6079) );
  nand_x1_sg U69515 ( .A(n6077), .B(n6081), .X(n6080) );
  nor_x1_sg U69516 ( .A(n28135), .B(n28133), .X(n28249) );
  nor_x1_sg U69517 ( .A(n20501), .B(n20498), .X(n20653) );
  nor_x1_sg U69518 ( .A(n19844), .B(n19841), .X(n20013) );
  nor_x1_sg U69519 ( .A(n6715), .B(n6712), .X(n19209) );
  nor_x1_sg U69520 ( .A(n21270), .B(n21267), .X(n21423) );
  inv_x1_sg U69521 ( .A(n26035), .X(n50548) );
  inv_x1_sg U69522 ( .A(n21418), .X(n45959) );
  inv_x1_sg U69523 ( .A(n20648), .X(n45950) );
  inv_x1_sg U69524 ( .A(n20316), .X(n46400) );
  inv_x1_sg U69525 ( .A(n19790), .X(n46393) );
  inv_x1_sg U69526 ( .A(n20008), .X(n45941) );
  inv_x1_sg U69527 ( .A(n28244), .X(n45103) );
  inv_x1_sg U69528 ( .A(n19349), .X(n46437) );
  inv_x1_sg U69529 ( .A(n19204), .X(n45932) );
  nor_x1_sg U69530 ( .A(n6264), .B(n6265), .X(n6263) );
  nor_x1_sg U69531 ( .A(n46340), .B(n46297), .X(n6265) );
  nor_x1_sg U69532 ( .A(n6266), .B(n42282), .X(n6264) );
  inv_x1_sg U69533 ( .A(n6266), .X(n46297) );
  nor_x1_sg U69534 ( .A(n6309), .B(n6310), .X(n6308) );
  nor_x1_sg U69535 ( .A(n46294), .B(n46252), .X(n6310) );
  nor_x1_sg U69536 ( .A(n6311), .B(n42281), .X(n6309) );
  inv_x1_sg U69537 ( .A(n6311), .X(n46252) );
  nor_x1_sg U69538 ( .A(n6353), .B(n6354), .X(n6352) );
  nor_x1_sg U69539 ( .A(n46249), .B(n46206), .X(n6354) );
  nor_x1_sg U69540 ( .A(n6355), .B(n42280), .X(n6353) );
  inv_x1_sg U69541 ( .A(n6355), .X(n46206) );
  nor_x1_sg U69542 ( .A(n6398), .B(n6399), .X(n6397) );
  nor_x1_sg U69543 ( .A(n46203), .B(n46161), .X(n6399) );
  nor_x1_sg U69544 ( .A(n6400), .B(n42279), .X(n6398) );
  inv_x1_sg U69545 ( .A(n6400), .X(n46161) );
  nor_x1_sg U69546 ( .A(n6442), .B(n6443), .X(n6441) );
  nor_x1_sg U69547 ( .A(n46158), .B(n46115), .X(n6443) );
  nor_x1_sg U69548 ( .A(n6444), .B(n42268), .X(n6442) );
  inv_x1_sg U69549 ( .A(n6444), .X(n46115) );
  nor_x1_sg U69550 ( .A(n6487), .B(n6488), .X(n6486) );
  nor_x1_sg U69551 ( .A(n46112), .B(n46070), .X(n6488) );
  nor_x1_sg U69552 ( .A(n6489), .B(n42278), .X(n6487) );
  inv_x1_sg U69553 ( .A(n6489), .X(n46070) );
  nor_x1_sg U69554 ( .A(n6531), .B(n6532), .X(n6530) );
  nor_x1_sg U69555 ( .A(n46067), .B(n46024), .X(n6532) );
  nor_x1_sg U69556 ( .A(n6533), .B(n42277), .X(n6531) );
  inv_x1_sg U69557 ( .A(n6533), .X(n46024) );
  nor_x1_sg U69558 ( .A(n6576), .B(n6577), .X(n6575) );
  nor_x1_sg U69559 ( .A(n46021), .B(n45979), .X(n6577) );
  nor_x1_sg U69560 ( .A(n6578), .B(n42230), .X(n6576) );
  inv_x1_sg U69561 ( .A(n6578), .X(n45979) );
  nor_x1_sg U69562 ( .A(n6620), .B(n6621), .X(n6619) );
  nor_x1_sg U69563 ( .A(n45976), .B(n45934), .X(n6621) );
  nor_x1_sg U69564 ( .A(n6622), .B(n42276), .X(n6620) );
  inv_x1_sg U69565 ( .A(n6622), .X(n45934) );
  inv_x1_sg U69566 ( .A(n21402), .X(n46140) );
  inv_x1_sg U69567 ( .A(n21410), .X(n46049) );
  inv_x1_sg U69568 ( .A(n21394), .X(n46231) );
  inv_x1_sg U69569 ( .A(n21386), .X(n46322) );
  inv_x1_sg U69570 ( .A(n21378), .X(n46411) );
  inv_x1_sg U69571 ( .A(n21370), .X(n46497) );
  inv_x1_sg U69572 ( .A(n21406), .X(n46095) );
  inv_x1_sg U69573 ( .A(n21414), .X(n46004) );
  inv_x1_sg U69574 ( .A(n21398), .X(n46186) );
  inv_x1_sg U69575 ( .A(n21390), .X(n46277) );
  inv_x1_sg U69576 ( .A(n20612), .X(n46355) );
  inv_x1_sg U69577 ( .A(n20616), .X(n46313) );
  inv_x1_sg U69578 ( .A(n20620), .X(n46268) );
  inv_x1_sg U69579 ( .A(n20624), .X(n46222) );
  inv_x1_sg U69580 ( .A(n20628), .X(n46177) );
  inv_x1_sg U69581 ( .A(n20632), .X(n46131) );
  inv_x1_sg U69582 ( .A(n20636), .X(n46086) );
  inv_x1_sg U69583 ( .A(n20640), .X(n46040) );
  inv_x1_sg U69584 ( .A(n20644), .X(n45995) );
  inv_x1_sg U69585 ( .A(n21382), .X(n46364) );
  inv_x1_sg U69586 ( .A(n20608), .X(n46402) );
  inv_x1_sg U69587 ( .A(n21374), .X(n46459) );
  inv_x1_sg U69588 ( .A(n19976), .X(n46304) );
  inv_x1_sg U69589 ( .A(n19980), .X(n46259) );
  inv_x1_sg U69590 ( .A(n19984), .X(n46213) );
  inv_x1_sg U69591 ( .A(n19988), .X(n46168) );
  inv_x1_sg U69592 ( .A(n19992), .X(n46122) );
  inv_x1_sg U69593 ( .A(n19996), .X(n46077) );
  inv_x1_sg U69594 ( .A(n20000), .X(n46031) );
  inv_x1_sg U69595 ( .A(n20004), .X(n45986) );
  inv_x1_sg U69596 ( .A(n19172), .X(n46295) );
  inv_x1_sg U69597 ( .A(n19176), .X(n46250) );
  inv_x1_sg U69598 ( .A(n19180), .X(n46204) );
  inv_x1_sg U69599 ( .A(n19184), .X(n46159) );
  inv_x1_sg U69600 ( .A(n19188), .X(n46113) );
  inv_x1_sg U69601 ( .A(n19192), .X(n46068) );
  inv_x1_sg U69602 ( .A(n19196), .X(n46022) );
  inv_x1_sg U69603 ( .A(n19200), .X(n45977) );
  inv_x1_sg U69604 ( .A(n19786), .X(n46442) );
  inv_x1_sg U69605 ( .A(n28240), .X(n45149) );
  inv_x1_sg U69606 ( .A(n28236), .X(n45194) );
  inv_x1_sg U69607 ( .A(n28232), .X(n45240) );
  inv_x1_sg U69608 ( .A(n28228), .X(n45285) );
  inv_x1_sg U69609 ( .A(n28224), .X(n45330) );
  inv_x1_sg U69610 ( .A(n28220), .X(n45375) );
  inv_x1_sg U69611 ( .A(n28216), .X(n45421) );
  inv_x1_sg U69612 ( .A(n20604), .X(n46450) );
  nand_x1_sg U69613 ( .A(n42312), .B(n40314), .X(n7601) );
  nor_x1_sg U69614 ( .A(n6218), .B(n6219), .X(n6217) );
  nor_x1_sg U69615 ( .A(n46385), .B(n46342), .X(n6219) );
  nor_x1_sg U69616 ( .A(n6220), .B(n6216), .X(n6218) );
  inv_x1_sg U69617 ( .A(n6220), .X(n46342) );
  nand_x1_sg U69618 ( .A(n45127), .B(n45105), .X(n28144) );
  nand_x1_sg U69619 ( .A(n28145), .B(n22401), .X(n28143) );
  nand_x1_sg U69620 ( .A(n45172), .B(n45151), .X(n28149) );
  nand_x1_sg U69621 ( .A(n28150), .B(n22354), .X(n28148) );
  nand_x1_sg U69622 ( .A(n45218), .B(n45196), .X(n28154) );
  nand_x1_sg U69623 ( .A(n28155), .B(n22306), .X(n28153) );
  nand_x1_sg U69624 ( .A(n45263), .B(n45242), .X(n28159) );
  nand_x1_sg U69625 ( .A(n28160), .B(n22259), .X(n28158) );
  nand_x1_sg U69626 ( .A(n45308), .B(n45287), .X(n28164) );
  nand_x1_sg U69627 ( .A(n28165), .B(n22211), .X(n28163) );
  nand_x1_sg U69628 ( .A(n45353), .B(n45332), .X(n28169) );
  nand_x1_sg U69629 ( .A(n28170), .B(n22164), .X(n28168) );
  nand_x1_sg U69630 ( .A(n45399), .B(n45377), .X(n28174) );
  nand_x1_sg U69631 ( .A(n28175), .B(n22116), .X(n28173) );
  inv_x1_sg U69632 ( .A(n19779), .X(n46530) );
  inv_x1_sg U69633 ( .A(n20155), .X(n46447) );
  inv_x1_sg U69634 ( .A(n21201), .X(n46539) );
  inv_x1_sg U69635 ( .A(n28082), .X(n45465) );
  inv_x1_sg U69636 ( .A(n27920), .X(n45489) );
  inv_x1_sg U69637 ( .A(n27743), .X(n45533) );
  inv_x1_sg U69638 ( .A(n27549), .X(n45578) );
  inv_x1_sg U69639 ( .A(n21059), .X(n45908) );
  inv_x1_sg U69640 ( .A(n27336), .X(n45622) );
  inv_x1_sg U69641 ( .A(n27106), .X(n45666) );
  inv_x1_sg U69642 ( .A(n20350), .X(n45898) );
  inv_x1_sg U69643 ( .A(n19617), .X(n45888) );
  inv_x1_sg U69644 ( .A(n19963), .X(n46486) );
  inv_x1_sg U69645 ( .A(n21249), .X(n45911) );
  inv_x1_sg U69646 ( .A(n20481), .X(n45901) );
  inv_x1_sg U69647 ( .A(n19824), .X(n45891) );
  nand_x1_sg U69648 ( .A(n27988), .B(n27987), .X(n27985) );
  nor_x1_sg U69649 ( .A(n27987), .B(n27988), .X(n27986) );
  nand_x1_sg U69650 ( .A(n28998), .B(n28997), .X(n28995) );
  nor_x1_sg U69651 ( .A(n28997), .B(n28998), .X(n28996) );
  nand_x1_sg U69652 ( .A(n29011), .B(n29010), .X(n29008) );
  nor_x1_sg U69653 ( .A(n29010), .B(n29011), .X(n29009) );
  nand_x1_sg U69654 ( .A(n29024), .B(n29023), .X(n29021) );
  nor_x1_sg U69655 ( .A(n29023), .B(n29024), .X(n29022) );
  nand_x1_sg U69656 ( .A(n29037), .B(n29036), .X(n29034) );
  nor_x1_sg U69657 ( .A(n29036), .B(n29037), .X(n29035) );
  nand_x1_sg U69658 ( .A(n29050), .B(n29049), .X(n29047) );
  nor_x1_sg U69659 ( .A(n29049), .B(n29050), .X(n29048) );
  nand_x1_sg U69660 ( .A(n29063), .B(n29062), .X(n29060) );
  nor_x1_sg U69661 ( .A(n29062), .B(n29063), .X(n29061) );
  nand_x1_sg U69662 ( .A(n29076), .B(n29075), .X(n29073) );
  nor_x1_sg U69663 ( .A(n29075), .B(n29076), .X(n29074) );
  nand_x1_sg U69664 ( .A(n27981), .B(n27980), .X(n27978) );
  nor_x1_sg U69665 ( .A(n27980), .B(n27981), .X(n27979) );
  nand_x1_sg U69666 ( .A(n39807), .B(n40568), .X(n17426) );
  nand_x1_sg U69667 ( .A(n39774), .B(n40570), .X(n17268) );
  nand_x1_sg U69668 ( .A(n21597), .B(n21598), .X(n21595) );
  nor_x1_sg U69669 ( .A(n42187), .B(n21598), .X(n21596) );
  nand_x1_sg U69670 ( .A(n29148), .B(n29149), .X(n29146) );
  nor_x1_sg U69671 ( .A(n42194), .B(n29149), .X(n29147) );
  nand_x1_sg U69672 ( .A(n21609), .B(n21610), .X(n21607) );
  nor_x1_sg U69673 ( .A(n42188), .B(n21610), .X(n21608) );
  nand_x1_sg U69674 ( .A(n29160), .B(n29161), .X(n29158) );
  nor_x1_sg U69675 ( .A(n42195), .B(n29161), .X(n29159) );
  nand_x1_sg U69676 ( .A(n21621), .B(n21622), .X(n21619) );
  nor_x1_sg U69677 ( .A(n42189), .B(n21622), .X(n21620) );
  nand_x1_sg U69678 ( .A(n29172), .B(n29173), .X(n29170) );
  nor_x1_sg U69679 ( .A(n42196), .B(n29173), .X(n29171) );
  nand_x1_sg U69680 ( .A(n21633), .B(n21634), .X(n21631) );
  nor_x1_sg U69681 ( .A(n42190), .B(n21634), .X(n21632) );
  nand_x1_sg U69682 ( .A(n29184), .B(n29185), .X(n29182) );
  nor_x1_sg U69683 ( .A(n42197), .B(n29185), .X(n29183) );
  nand_x1_sg U69684 ( .A(n21645), .B(n21646), .X(n21643) );
  nor_x1_sg U69685 ( .A(n42191), .B(n21646), .X(n21644) );
  nand_x1_sg U69686 ( .A(n21657), .B(n21658), .X(n21655) );
  nor_x1_sg U69687 ( .A(n42192), .B(n21658), .X(n21656) );
  nand_x1_sg U69688 ( .A(n21352), .B(n21186), .X(n21350) );
  nor_x1_sg U69689 ( .A(n42193), .B(n21186), .X(n21351) );
  nand_x1_sg U69690 ( .A(n28916), .B(n28741), .X(n28914) );
  nor_x1_sg U69691 ( .A(n42198), .B(n28741), .X(n28915) );
  nand_x1_sg U69692 ( .A(n29196), .B(n29197), .X(n29194) );
  nor_x1_sg U69693 ( .A(n29196), .B(n29197), .X(n29195) );
  nand_x1_sg U69694 ( .A(n29208), .B(n29209), .X(n29206) );
  nor_x1_sg U69695 ( .A(n29208), .B(n29209), .X(n29207) );
  nand_x1_sg U69696 ( .A(n21669), .B(n21670), .X(n21667) );
  nor_x1_sg U69697 ( .A(n21669), .B(n21670), .X(n21668) );
  nand_x1_sg U69698 ( .A(n29220), .B(n29221), .X(n29218) );
  nor_x1_sg U69699 ( .A(n29220), .B(n29221), .X(n29219) );
  nand_x1_sg U69700 ( .A(n21534), .B(n21356), .X(n21532) );
  nor_x1_sg U69701 ( .A(n21534), .B(n21356), .X(n21533) );
  nand_x1_sg U69702 ( .A(n29085), .B(n28920), .X(n29083) );
  nor_x1_sg U69703 ( .A(n29085), .B(n28920), .X(n29084) );
  nor_x1_sg U69704 ( .A(n19133), .B(n46632), .X(n19132) );
  nor_x1_sg U69705 ( .A(n19135), .B(n19131), .X(n19133) );
  nand_x1_sg U69706 ( .A(n19131), .B(n19135), .X(n19134) );
  nand_x1_sg U69707 ( .A(n22514), .B(n22513), .X(n26945) );
  nand_x1_sg U69708 ( .A(n45020), .B(n45049), .X(n26947) );
  nand_x1_sg U69709 ( .A(n39802), .B(n6831), .X(n7443) );
  nand_x1_sg U69710 ( .A(n39850), .B(n40315), .X(n7185) );
  nand_x1_sg U69711 ( .A(n22503), .B(n28267), .X(n28360) );
  nand_x1_sg U69712 ( .A(n44994), .B(n45035), .X(n28362) );
  nand_x1_sg U69713 ( .A(n22457), .B(n28273), .X(n28357) );
  nand_x1_sg U69714 ( .A(n45060), .B(n45078), .X(n28359) );
  nand_x1_sg U69715 ( .A(n45037), .B(n27984), .X(n28115) );
  nand_x1_sg U69716 ( .A(n45001), .B(n27980), .X(n28117) );
  nand_x1_sg U69717 ( .A(n22411), .B(n28279), .X(n28354) );
  nand_x1_sg U69718 ( .A(n45106), .B(n45125), .X(n28356) );
  nand_x1_sg U69719 ( .A(n22483), .B(n27814), .X(n27962) );
  nand_x1_sg U69720 ( .A(n45004), .B(n45039), .X(n27964) );
  nand_x1_sg U69721 ( .A(n45081), .B(n27991), .X(n28112) );
  nand_x1_sg U69722 ( .A(n45057), .B(n27987), .X(n28114) );
  nand_x1_sg U69723 ( .A(n22363), .B(n28285), .X(n28351) );
  nand_x1_sg U69724 ( .A(n45152), .B(n45170), .X(n28353) );
  nand_x1_sg U69725 ( .A(n22492), .B(n27628), .X(n27794) );
  nand_x1_sg U69726 ( .A(n45007), .B(n45041), .X(n27796) );
  nand_x1_sg U69727 ( .A(n22437), .B(n27820), .X(n27959) );
  nand_x1_sg U69728 ( .A(n45056), .B(n45083), .X(n27961) );
  nand_x1_sg U69729 ( .A(n22394), .B(n27997), .X(n28109) );
  nand_x1_sg U69730 ( .A(n45101), .B(n45128), .X(n28111) );
  nand_x1_sg U69731 ( .A(n22316), .B(n28291), .X(n28348) );
  nand_x1_sg U69732 ( .A(n45197), .B(n45216), .X(n28350) );
  nand_x1_sg U69733 ( .A(n22502), .B(n28635), .X(n28803) );
  nand_x1_sg U69734 ( .A(n44985), .B(n45029), .X(n28805) );
  nand_x1_sg U69735 ( .A(n22487), .B(n27425), .X(n27609) );
  nand_x1_sg U69736 ( .A(n45010), .B(n45043), .X(n27611) );
  nand_x1_sg U69737 ( .A(n22446), .B(n27634), .X(n27791) );
  nand_x1_sg U69738 ( .A(n45055), .B(n45085), .X(n27793) );
  nand_x1_sg U69739 ( .A(n22389), .B(n27826), .X(n27956) );
  nand_x1_sg U69740 ( .A(n45100), .B(n45130), .X(n27958) );
  nand_x1_sg U69741 ( .A(n22347), .B(n28003), .X(n28106) );
  nand_x1_sg U69742 ( .A(n45148), .B(n45173), .X(n28108) );
  nand_x1_sg U69743 ( .A(n22268), .B(n28297), .X(n28345) );
  nand_x1_sg U69744 ( .A(n45243), .B(n45261), .X(n28347) );
  nand_x1_sg U69745 ( .A(n6723), .B(n21443), .X(n21582) );
  nand_x1_sg U69746 ( .A(n45815), .B(n45873), .X(n21584) );
  nand_x1_sg U69747 ( .A(n20870), .B(n20874), .X(n21050) );
  nand_x1_sg U69748 ( .A(n46000), .B(n46014), .X(n21052) );
  nand_x1_sg U69749 ( .A(n20684), .B(n20687), .X(n20829) );
  nand_x1_sg U69750 ( .A(n45953), .B(n42201), .X(n20831) );
  nand_x1_sg U69751 ( .A(n22496), .B(n28474), .X(n28615) );
  nand_x1_sg U69752 ( .A(n44988), .B(n45031), .X(n28617) );
  nand_x1_sg U69753 ( .A(n22456), .B(n28641), .X(n28800) );
  nand_x1_sg U69754 ( .A(n45063), .B(n45072), .X(n28802) );
  nand_x1_sg U69755 ( .A(n22497), .B(n28994), .X(n29133) );
  nand_x1_sg U69756 ( .A(n44979), .B(n45025), .X(n29135) );
  nand_x1_sg U69757 ( .A(n22484), .B(n27203), .X(n27405) );
  nand_x1_sg U69758 ( .A(n45013), .B(n45045), .X(n27407) );
  nand_x1_sg U69759 ( .A(n22441), .B(n27431), .X(n27606) );
  nand_x1_sg U69760 ( .A(n45054), .B(n45087), .X(n27608) );
  nand_x1_sg U69761 ( .A(n22399), .B(n27640), .X(n27788) );
  nand_x1_sg U69762 ( .A(n45099), .B(n45132), .X(n27790) );
  nand_x1_sg U69763 ( .A(n22342), .B(n27832), .X(n27953) );
  nand_x1_sg U69764 ( .A(n45147), .B(n45175), .X(n27955) );
  nand_x1_sg U69765 ( .A(n22299), .B(n28009), .X(n28103) );
  nand_x1_sg U69766 ( .A(n45193), .B(n45219), .X(n28105) );
  nand_x1_sg U69767 ( .A(n22221), .B(n28303), .X(n28342) );
  nand_x1_sg U69768 ( .A(n45288), .B(n45306), .X(n28344) );
  nand_x1_sg U69769 ( .A(n45919), .B(n21450), .X(n21579) );
  nand_x1_sg U69770 ( .A(n45916), .B(n21445), .X(n21581) );
  nand_x1_sg U69771 ( .A(n20877), .B(n20881), .X(n21047) );
  nand_x1_sg U69772 ( .A(n46045), .B(n46060), .X(n21049) );
  nand_x1_sg U69773 ( .A(n20691), .B(n20694), .X(n20826) );
  nand_x1_sg U69774 ( .A(n45998), .B(n42148), .X(n20828) );
  nand_x1_sg U69775 ( .A(n22517), .B(n28380), .X(n28455) );
  nand_x1_sg U69776 ( .A(n44991), .B(n45033), .X(n28457) );
  nand_x1_sg U69777 ( .A(n22451), .B(n28480), .X(n28612) );
  nand_x1_sg U69778 ( .A(n45062), .B(n45074), .X(n28614) );
  nand_x1_sg U69779 ( .A(n22410), .B(n28647), .X(n28797) );
  nand_x1_sg U69780 ( .A(n45109), .B(n45119), .X(n28799) );
  nand_x1_sg U69781 ( .A(n22518), .B(n28823), .X(n28973) );
  nand_x1_sg U69782 ( .A(n44982), .B(n45027), .X(n28975) );
  nand_x1_sg U69783 ( .A(n45068), .B(n29001), .X(n29130) );
  nand_x1_sg U69784 ( .A(n45065), .B(n28997), .X(n29132) );
  nand_x1_sg U69785 ( .A(n22493), .B(n26964), .X(n27184) );
  nand_x1_sg U69786 ( .A(n45016), .B(n45047), .X(n27186) );
  nand_x1_sg U69787 ( .A(n22438), .B(n27209), .X(n27402) );
  nand_x1_sg U69788 ( .A(n45053), .B(n45089), .X(n27404) );
  nand_x1_sg U69789 ( .A(n22393), .B(n27437), .X(n27603) );
  nand_x1_sg U69790 ( .A(n45098), .B(n45134), .X(n27605) );
  nand_x1_sg U69791 ( .A(n22352), .B(n27646), .X(n27785) );
  nand_x1_sg U69792 ( .A(n45146), .B(n45177), .X(n27787) );
  nand_x1_sg U69793 ( .A(n22294), .B(n27838), .X(n27950) );
  nand_x1_sg U69794 ( .A(n45192), .B(n45221), .X(n27952) );
  nand_x1_sg U69795 ( .A(n22252), .B(n28015), .X(n28100) );
  nand_x1_sg U69796 ( .A(n45239), .B(n45264), .X(n28102) );
  nand_x1_sg U69797 ( .A(n22173), .B(n28309), .X(n28339) );
  nand_x1_sg U69798 ( .A(n45333), .B(n45351), .X(n28341) );
  nand_x1_sg U69799 ( .A(n6631), .B(n21456), .X(n21576) );
  nand_x1_sg U69800 ( .A(n45962), .B(n45965), .X(n21578) );
  nand_x1_sg U69801 ( .A(n20884), .B(n20888), .X(n21044) );
  nand_x1_sg U69802 ( .A(n46091), .B(n46105), .X(n21046) );
  nand_x1_sg U69803 ( .A(n20698), .B(n20701), .X(n20823) );
  nand_x1_sg U69804 ( .A(n46043), .B(n42204), .X(n20825) );
  nand_x1_sg U69805 ( .A(n22471), .B(n28386), .X(n28452) );
  nand_x1_sg U69806 ( .A(n45061), .B(n45076), .X(n28454) );
  nand_x1_sg U69807 ( .A(n22404), .B(n28486), .X(n28609) );
  nand_x1_sg U69808 ( .A(n45108), .B(n45121), .X(n28611) );
  nand_x1_sg U69809 ( .A(n22362), .B(n28653), .X(n28794) );
  nand_x1_sg U69810 ( .A(n45155), .B(n45164), .X(n28796) );
  nand_x1_sg U69811 ( .A(n22472), .B(n28829), .X(n28970) );
  nand_x1_sg U69812 ( .A(n45064), .B(n45070), .X(n28972) );
  nand_x1_sg U69813 ( .A(n22405), .B(n29007), .X(n29127) );
  nand_x1_sg U69814 ( .A(n45111), .B(n45115), .X(n29129) );
  nand_x1_sg U69815 ( .A(n22468), .B(n22467), .X(n26942) );
  nand_x1_sg U69816 ( .A(n45051), .B(n45093), .X(n26944) );
  nand_x1_sg U69817 ( .A(n22447), .B(n26970), .X(n27181) );
  nand_x1_sg U69818 ( .A(n45052), .B(n45091), .X(n27183) );
  nand_x1_sg U69819 ( .A(n22390), .B(n27215), .X(n27399) );
  nand_x1_sg U69820 ( .A(n45097), .B(n45136), .X(n27401) );
  nand_x1_sg U69821 ( .A(n22346), .B(n27443), .X(n27600) );
  nand_x1_sg U69822 ( .A(n45145), .B(n45179), .X(n27602) );
  nand_x1_sg U69823 ( .A(n22304), .B(n27652), .X(n27782) );
  nand_x1_sg U69824 ( .A(n45191), .B(n45223), .X(n27784) );
  nand_x1_sg U69825 ( .A(n22247), .B(n27844), .X(n27947) );
  nand_x1_sg U69826 ( .A(n45238), .B(n45266), .X(n27949) );
  nand_x1_sg U69827 ( .A(n22204), .B(n28021), .X(n28097) );
  nand_x1_sg U69828 ( .A(n45284), .B(n45309), .X(n28099) );
  nand_x1_sg U69829 ( .A(n22126), .B(n28315), .X(n28336) );
  nand_x1_sg U69830 ( .A(n45378), .B(n45397), .X(n28338) );
  nand_x1_sg U69831 ( .A(n46010), .B(n21463), .X(n21573) );
  nand_x1_sg U69832 ( .A(n46007), .B(n21458), .X(n21575) );
  nand_x1_sg U69833 ( .A(n20891), .B(n20895), .X(n21041) );
  nand_x1_sg U69834 ( .A(n46136), .B(n46151), .X(n21043) );
  nand_x1_sg U69835 ( .A(n20705), .B(n20708), .X(n20820) );
  nand_x1_sg U69836 ( .A(n46089), .B(n42150), .X(n20822) );
  nand_x1_sg U69837 ( .A(n20227), .B(n20231), .X(n20341) );
  nand_x1_sg U69838 ( .A(n45991), .B(n46017), .X(n20343) );
  nand_x1_sg U69839 ( .A(n22425), .B(n28392), .X(n28449) );
  nand_x1_sg U69840 ( .A(n45107), .B(n45123), .X(n28451) );
  nand_x1_sg U69841 ( .A(n22357), .B(n28492), .X(n28606) );
  nand_x1_sg U69842 ( .A(n45154), .B(n45166), .X(n28608) );
  nand_x1_sg U69843 ( .A(n22315), .B(n28659), .X(n28791) );
  nand_x1_sg U69844 ( .A(n45200), .B(n45210), .X(n28793) );
  nand_x1_sg U69845 ( .A(n22426), .B(n28835), .X(n28967) );
  nand_x1_sg U69846 ( .A(n45110), .B(n45117), .X(n28969) );
  nand_x1_sg U69847 ( .A(n45160), .B(n29014), .X(n29124) );
  nand_x1_sg U69848 ( .A(n45157), .B(n29010), .X(n29126) );
  nand_x1_sg U69849 ( .A(n22422), .B(n22421), .X(n26939) );
  nand_x1_sg U69850 ( .A(n45095), .B(n45140), .X(n26941) );
  nand_x1_sg U69851 ( .A(n22400), .B(n26976), .X(n27178) );
  nand_x1_sg U69852 ( .A(n45096), .B(n45138), .X(n27180) );
  nand_x1_sg U69853 ( .A(n22343), .B(n27221), .X(n27396) );
  nand_x1_sg U69854 ( .A(n45144), .B(n45181), .X(n27398) );
  nand_x1_sg U69855 ( .A(n22298), .B(n27449), .X(n27597) );
  nand_x1_sg U69856 ( .A(n45190), .B(n45225), .X(n27599) );
  nand_x1_sg U69857 ( .A(n22257), .B(n27658), .X(n27779) );
  nand_x1_sg U69858 ( .A(n45237), .B(n45268), .X(n27781) );
  nand_x1_sg U69859 ( .A(n22199), .B(n27850), .X(n27944) );
  nand_x1_sg U69860 ( .A(n45283), .B(n45311), .X(n27946) );
  nand_x1_sg U69861 ( .A(n22157), .B(n28027), .X(n28094) );
  nand_x1_sg U69862 ( .A(n45329), .B(n45354), .X(n28096) );
  nand_x1_sg U69863 ( .A(n22078), .B(n28210), .X(n28207) );
  nand_x1_sg U69864 ( .A(n45424), .B(n45442), .X(n28209) );
  nand_x1_sg U69865 ( .A(n6542), .B(n21469), .X(n21570) );
  nand_x1_sg U69866 ( .A(n46052), .B(n46056), .X(n21572) );
  nand_x1_sg U69867 ( .A(n20898), .B(n20902), .X(n21038) );
  nand_x1_sg U69868 ( .A(n46182), .B(n46196), .X(n21040) );
  nand_x1_sg U69869 ( .A(n20712), .B(n20715), .X(n20817) );
  nand_x1_sg U69870 ( .A(n46134), .B(n42151), .X(n20819) );
  nand_x1_sg U69871 ( .A(n20044), .B(n20047), .X(n20186) );
  nand_x1_sg U69872 ( .A(n45944), .B(n42202), .X(n20188) );
  nand_x1_sg U69873 ( .A(n20234), .B(n20238), .X(n20338) );
  nand_x1_sg U69874 ( .A(n46036), .B(n46063), .X(n20340) );
  nand_x1_sg U69875 ( .A(n22377), .B(n28398), .X(n28446) );
  nand_x1_sg U69876 ( .A(n45153), .B(n45168), .X(n28448) );
  nand_x1_sg U69877 ( .A(n22309), .B(n28498), .X(n28603) );
  nand_x1_sg U69878 ( .A(n45199), .B(n45212), .X(n28605) );
  nand_x1_sg U69879 ( .A(n22267), .B(n28665), .X(n28788) );
  nand_x1_sg U69880 ( .A(n45246), .B(n45255), .X(n28790) );
  nand_x1_sg U69881 ( .A(n22378), .B(n28841), .X(n28964) );
  nand_x1_sg U69882 ( .A(n45156), .B(n45162), .X(n28966) );
  nand_x1_sg U69883 ( .A(n22310), .B(n29020), .X(n29121) );
  nand_x1_sg U69884 ( .A(n45202), .B(n45206), .X(n29123) );
  nand_x1_sg U69885 ( .A(n22374), .B(n22373), .X(n26936) );
  nand_x1_sg U69886 ( .A(n45142), .B(n45185), .X(n26938) );
  nand_x1_sg U69887 ( .A(n22353), .B(n26982), .X(n27175) );
  nand_x1_sg U69888 ( .A(n45143), .B(n45183), .X(n27177) );
  nand_x1_sg U69889 ( .A(n22295), .B(n27227), .X(n27393) );
  nand_x1_sg U69890 ( .A(n45189), .B(n45227), .X(n27395) );
  nand_x1_sg U69891 ( .A(n22251), .B(n27455), .X(n27594) );
  nand_x1_sg U69892 ( .A(n45236), .B(n45270), .X(n27596) );
  nand_x1_sg U69893 ( .A(n22209), .B(n27664), .X(n27776) );
  nand_x1_sg U69894 ( .A(n45282), .B(n45313), .X(n27778) );
  nand_x1_sg U69895 ( .A(n22152), .B(n27856), .X(n27941) );
  nand_x1_sg U69896 ( .A(n45328), .B(n45356), .X(n27943) );
  nand_x1_sg U69897 ( .A(n22109), .B(n28033), .X(n28091) );
  nand_x1_sg U69898 ( .A(n45374), .B(n45400), .X(n28093) );
  nand_x1_sg U69899 ( .A(n22032), .B(n28075), .X(n28072) );
  nand_x1_sg U69900 ( .A(n45468), .B(n45487), .X(n28074) );
  nand_x1_sg U69901 ( .A(n46101), .B(n21476), .X(n21567) );
  nand_x1_sg U69902 ( .A(n46098), .B(n21471), .X(n21569) );
  nand_x1_sg U69903 ( .A(n20905), .B(n20909), .X(n21035) );
  nand_x1_sg U69904 ( .A(n46227), .B(n46242), .X(n21037) );
  nand_x1_sg U69905 ( .A(n20719), .B(n20722), .X(n20814) );
  nand_x1_sg U69906 ( .A(n46180), .B(n42207), .X(n20816) );
  nand_x1_sg U69907 ( .A(n20051), .B(n20054), .X(n20183) );
  nand_x1_sg U69908 ( .A(n45989), .B(n42203), .X(n20185) );
  nand_x1_sg U69909 ( .A(n20241), .B(n20245), .X(n20335) );
  nand_x1_sg U69910 ( .A(n46082), .B(n46108), .X(n20337) );
  nand_x1_sg U69911 ( .A(n22330), .B(n28404), .X(n28443) );
  nand_x1_sg U69912 ( .A(n45198), .B(n45214), .X(n28445) );
  nand_x1_sg U69913 ( .A(n22262), .B(n28504), .X(n28600) );
  nand_x1_sg U69914 ( .A(n45245), .B(n45257), .X(n28602) );
  nand_x1_sg U69915 ( .A(n22220), .B(n28671), .X(n28785) );
  nand_x1_sg U69916 ( .A(n45291), .B(n45300), .X(n28787) );
  nand_x1_sg U69917 ( .A(n22331), .B(n28847), .X(n28961) );
  nand_x1_sg U69918 ( .A(n45201), .B(n45208), .X(n28963) );
  nand_x1_sg U69919 ( .A(n45251), .B(n29027), .X(n29118) );
  nand_x1_sg U69920 ( .A(n45248), .B(n29023), .X(n29120) );
  nand_x1_sg U69921 ( .A(n22327), .B(n22326), .X(n26933) );
  nand_x1_sg U69922 ( .A(n45187), .B(n45231), .X(n26935) );
  nand_x1_sg U69923 ( .A(n22305), .B(n26988), .X(n27172) );
  nand_x1_sg U69924 ( .A(n45188), .B(n45229), .X(n27174) );
  nand_x1_sg U69925 ( .A(n22248), .B(n27233), .X(n27390) );
  nand_x1_sg U69926 ( .A(n45235), .B(n45272), .X(n27392) );
  nand_x1_sg U69927 ( .A(n22203), .B(n27461), .X(n27591) );
  nand_x1_sg U69928 ( .A(n45281), .B(n45315), .X(n27593) );
  nand_x1_sg U69929 ( .A(n22162), .B(n27670), .X(n27773) );
  nand_x1_sg U69930 ( .A(n45327), .B(n45358), .X(n27775) );
  nand_x1_sg U69931 ( .A(n22104), .B(n27862), .X(n27938) );
  nand_x1_sg U69932 ( .A(n45373), .B(n45402), .X(n27940) );
  nand_x1_sg U69933 ( .A(n22063), .B(n28039), .X(n28088) );
  nand_x1_sg U69934 ( .A(n45420), .B(n45444), .X(n28090) );
  nand_x1_sg U69935 ( .A(n21985), .B(n27913), .X(n27910) );
  nand_x1_sg U69936 ( .A(n45513), .B(n45531), .X(n27912) );
  nand_x1_sg U69937 ( .A(n6453), .B(n21482), .X(n21564) );
  nand_x1_sg U69938 ( .A(n46143), .B(n46147), .X(n21566) );
  nand_x1_sg U69939 ( .A(n20912), .B(n20916), .X(n21032) );
  nand_x1_sg U69940 ( .A(n46273), .B(n46287), .X(n21034) );
  nand_x1_sg U69941 ( .A(n20726), .B(n20729), .X(n20811) );
  nand_x1_sg U69942 ( .A(n46225), .B(n42152), .X(n20813) );
  nand_x1_sg U69943 ( .A(n20058), .B(n20061), .X(n20180) );
  nand_x1_sg U69944 ( .A(n46034), .B(n42149), .X(n20182) );
  nand_x1_sg U69945 ( .A(n20248), .B(n20252), .X(n20332) );
  nand_x1_sg U69946 ( .A(n46127), .B(n46154), .X(n20334) );
  nand_x1_sg U69947 ( .A(n22282), .B(n28410), .X(n28440) );
  nand_x1_sg U69948 ( .A(n45244), .B(n45259), .X(n28442) );
  nand_x1_sg U69949 ( .A(n22214), .B(n28510), .X(n28597) );
  nand_x1_sg U69950 ( .A(n45290), .B(n45302), .X(n28599) );
  nand_x1_sg U69951 ( .A(n22172), .B(n28677), .X(n28782) );
  nand_x1_sg U69952 ( .A(n45336), .B(n45345), .X(n28784) );
  nand_x1_sg U69953 ( .A(n22283), .B(n28853), .X(n28958) );
  nand_x1_sg U69954 ( .A(n45247), .B(n45253), .X(n28960) );
  nand_x1_sg U69955 ( .A(n22215), .B(n29033), .X(n29115) );
  nand_x1_sg U69956 ( .A(n45293), .B(n45296), .X(n29117) );
  nand_x1_sg U69957 ( .A(n22279), .B(n22278), .X(n26930) );
  nand_x1_sg U69958 ( .A(n45233), .B(n45276), .X(n26932) );
  nand_x1_sg U69959 ( .A(n22258), .B(n26994), .X(n27169) );
  nand_x1_sg U69960 ( .A(n45234), .B(n45274), .X(n27171) );
  nand_x1_sg U69961 ( .A(n22200), .B(n27239), .X(n27387) );
  nand_x1_sg U69962 ( .A(n45280), .B(n45317), .X(n27389) );
  nand_x1_sg U69963 ( .A(n22156), .B(n27467), .X(n27588) );
  nand_x1_sg U69964 ( .A(n45326), .B(n45360), .X(n27590) );
  nand_x1_sg U69965 ( .A(n22114), .B(n27676), .X(n27770) );
  nand_x1_sg U69966 ( .A(n45372), .B(n45404), .X(n27772) );
  nand_x1_sg U69967 ( .A(n22058), .B(n27868), .X(n27935) );
  nand_x1_sg U69968 ( .A(n45419), .B(n45446), .X(n27937) );
  nand_x1_sg U69969 ( .A(n22016), .B(n28045), .X(n28085) );
  nand_x1_sg U69970 ( .A(n45464), .B(n45492), .X(n28087) );
  nand_x1_sg U69971 ( .A(n21939), .B(n27736), .X(n27733) );
  nand_x1_sg U69972 ( .A(n45557), .B(n45576), .X(n27735) );
  nand_x1_sg U69973 ( .A(n46192), .B(n21489), .X(n21561) );
  nand_x1_sg U69974 ( .A(n46189), .B(n21484), .X(n21563) );
  nand_x1_sg U69975 ( .A(n20919), .B(n20923), .X(n21029) );
  nand_x1_sg U69976 ( .A(n46318), .B(n46333), .X(n21031) );
  nand_x1_sg U69977 ( .A(n20733), .B(n20736), .X(n20808) );
  nand_x1_sg U69978 ( .A(n46271), .B(n42210), .X(n20810) );
  nand_x1_sg U69979 ( .A(n20065), .B(n20068), .X(n20177) );
  nand_x1_sg U69980 ( .A(n46080), .B(n42205), .X(n20179) );
  nand_x1_sg U69981 ( .A(n20255), .B(n20259), .X(n20329) );
  nand_x1_sg U69982 ( .A(n46173), .B(n46199), .X(n20331) );
  nand_x1_sg U69983 ( .A(n19240), .B(n19243), .X(n19380) );
  nand_x1_sg U69984 ( .A(n45935), .B(n42218), .X(n19382) );
  nand_x1_sg U69985 ( .A(n22235), .B(n28416), .X(n28437) );
  nand_x1_sg U69986 ( .A(n45289), .B(n45304), .X(n28439) );
  nand_x1_sg U69987 ( .A(n22167), .B(n28516), .X(n28594) );
  nand_x1_sg U69988 ( .A(n45335), .B(n45347), .X(n28596) );
  nand_x1_sg U69989 ( .A(n22125), .B(n28683), .X(n28779) );
  nand_x1_sg U69990 ( .A(n45381), .B(n45391), .X(n28781) );
  nand_x1_sg U69991 ( .A(n22236), .B(n28859), .X(n28955) );
  nand_x1_sg U69992 ( .A(n45292), .B(n45298), .X(n28957) );
  nand_x1_sg U69993 ( .A(n45341), .B(n29040), .X(n29112) );
  nand_x1_sg U69994 ( .A(n45338), .B(n29036), .X(n29114) );
  nand_x1_sg U69995 ( .A(n22232), .B(n22231), .X(n26927) );
  nand_x1_sg U69996 ( .A(n45278), .B(n45321), .X(n26929) );
  nand_x1_sg U69997 ( .A(n22210), .B(n27000), .X(n27166) );
  nand_x1_sg U69998 ( .A(n45279), .B(n45319), .X(n27168) );
  nand_x1_sg U69999 ( .A(n22153), .B(n27245), .X(n27384) );
  nand_x1_sg U70000 ( .A(n45325), .B(n45362), .X(n27386) );
  nand_x1_sg U70001 ( .A(n22108), .B(n27473), .X(n27585) );
  nand_x1_sg U70002 ( .A(n45371), .B(n45406), .X(n27587) );
  nand_x1_sg U70003 ( .A(n22068), .B(n27682), .X(n27767) );
  nand_x1_sg U70004 ( .A(n45418), .B(n45448), .X(n27769) );
  nand_x1_sg U70005 ( .A(n22011), .B(n27874), .X(n27932) );
  nand_x1_sg U70006 ( .A(n45463), .B(n45494), .X(n27934) );
  nand_x1_sg U70007 ( .A(n21970), .B(n27926), .X(n27923) );
  nand_x1_sg U70008 ( .A(n45512), .B(n45536), .X(n27925) );
  nand_x1_sg U70009 ( .A(n21892), .B(n27542), .X(n27539) );
  nand_x1_sg U70010 ( .A(n45602), .B(n45620), .X(n27541) );
  nand_x1_sg U70011 ( .A(n6364), .B(n21495), .X(n21558) );
  nand_x1_sg U70012 ( .A(n46234), .B(n46238), .X(n21560) );
  nand_x1_sg U70013 ( .A(n20926), .B(n20930), .X(n21026) );
  nand_x1_sg U70014 ( .A(n46360), .B(n46374), .X(n21028) );
  nand_x1_sg U70015 ( .A(n20740), .B(n20743), .X(n20805) );
  nand_x1_sg U70016 ( .A(n46316), .B(n42212), .X(n20807) );
  nand_x1_sg U70017 ( .A(n19421), .B(n19425), .X(n19608) );
  nand_x1_sg U70018 ( .A(n45982), .B(n46020), .X(n19610) );
  nand_x1_sg U70019 ( .A(n20072), .B(n20075), .X(n20174) );
  nand_x1_sg U70020 ( .A(n46125), .B(n42206), .X(n20176) );
  nand_x1_sg U70021 ( .A(n20262), .B(n20266), .X(n20326) );
  nand_x1_sg U70022 ( .A(n46218), .B(n46245), .X(n20328) );
  nand_x1_sg U70023 ( .A(n19247), .B(n19250), .X(n19377) );
  nand_x1_sg U70024 ( .A(n45980), .B(n42261), .X(n19379) );
  nand_x1_sg U70025 ( .A(n22187), .B(n28422), .X(n28434) );
  nand_x1_sg U70026 ( .A(n45334), .B(n45349), .X(n28436) );
  nand_x1_sg U70027 ( .A(n22119), .B(n28431), .X(n28591) );
  nand_x1_sg U70028 ( .A(n45380), .B(n45393), .X(n28593) );
  nand_x1_sg U70029 ( .A(n22077), .B(n28689), .X(n28776) );
  nand_x1_sg U70030 ( .A(n45427), .B(n45436), .X(n28778) );
  nand_x1_sg U70031 ( .A(n22188), .B(n28865), .X(n28952) );
  nand_x1_sg U70032 ( .A(n45337), .B(n45343), .X(n28954) );
  nand_x1_sg U70033 ( .A(n22120), .B(n29046), .X(n29109) );
  nand_x1_sg U70034 ( .A(n45383), .B(n45387), .X(n29111) );
  nand_x1_sg U70035 ( .A(n22184), .B(n22183), .X(n26924) );
  nand_x1_sg U70036 ( .A(n45323), .B(n45366), .X(n26926) );
  nand_x1_sg U70037 ( .A(n22163), .B(n27006), .X(n27163) );
  nand_x1_sg U70038 ( .A(n45324), .B(n45364), .X(n27165) );
  nand_x1_sg U70039 ( .A(n22105), .B(n27251), .X(n27381) );
  nand_x1_sg U70040 ( .A(n45370), .B(n45408), .X(n27383) );
  nand_x1_sg U70041 ( .A(n22062), .B(n27479), .X(n27582) );
  nand_x1_sg U70042 ( .A(n45417), .B(n45450), .X(n27584) );
  nand_x1_sg U70043 ( .A(n22021), .B(n27688), .X(n27764) );
  nand_x1_sg U70044 ( .A(n45462), .B(n45496), .X(n27766) );
  nand_x1_sg U70045 ( .A(n21965), .B(n27880), .X(n27929) );
  nand_x1_sg U70046 ( .A(n45511), .B(n45538), .X(n27931) );
  nand_x1_sg U70047 ( .A(n21923), .B(n27749), .X(n27746) );
  nand_x1_sg U70048 ( .A(n45556), .B(n45581), .X(n27748) );
  nand_x1_sg U70049 ( .A(n21846), .B(n27329), .X(n27326) );
  nand_x1_sg U70050 ( .A(n45664), .B(n45646), .X(n27328) );
  nand_x1_sg U70051 ( .A(n46283), .B(n21502), .X(n21555) );
  nand_x1_sg U70052 ( .A(n46280), .B(n21497), .X(n21557) );
  nand_x1_sg U70053 ( .A(n20933), .B(n20937), .X(n21023) );
  nand_x1_sg U70054 ( .A(n46407), .B(n46422), .X(n21025) );
  nand_x1_sg U70055 ( .A(n20747), .B(n20750), .X(n20802) );
  nand_x1_sg U70056 ( .A(n46358), .B(n42214), .X(n20804) );
  nand_x1_sg U70057 ( .A(n19428), .B(n19432), .X(n19605) );
  nand_x1_sg U70058 ( .A(n46027), .B(n46066), .X(n19607) );
  nand_x1_sg U70059 ( .A(n20079), .B(n20082), .X(n20171) );
  nand_x1_sg U70060 ( .A(n46171), .B(n42208), .X(n20173) );
  nand_x1_sg U70061 ( .A(n20269), .B(n20273), .X(n20323) );
  nand_x1_sg U70062 ( .A(n46264), .B(n46290), .X(n20325) );
  nand_x1_sg U70063 ( .A(n19254), .B(n19257), .X(n19374) );
  nand_x1_sg U70064 ( .A(n46025), .B(n42219), .X(n19376) );
  nand_x1_sg U70065 ( .A(n22140), .B(n28333), .X(n28330) );
  nand_x1_sg U70066 ( .A(n45379), .B(n45395), .X(n28332) );
  nand_x1_sg U70067 ( .A(n22072), .B(n28327), .X(n28588) );
  nand_x1_sg U70068 ( .A(n45426), .B(n45438), .X(n28590) );
  nand_x1_sg U70069 ( .A(n22031), .B(n28695), .X(n28773) );
  nand_x1_sg U70070 ( .A(n45471), .B(n45481), .X(n28775) );
  nand_x1_sg U70071 ( .A(n22141), .B(n28871), .X(n28949) );
  nand_x1_sg U70072 ( .A(n45382), .B(n45389), .X(n28951) );
  nand_x1_sg U70073 ( .A(n45432), .B(n29053), .X(n29106) );
  nand_x1_sg U70074 ( .A(n45429), .B(n29049), .X(n29108) );
  nand_x1_sg U70075 ( .A(n22137), .B(n22136), .X(n26921) );
  nand_x1_sg U70076 ( .A(n45368), .B(n45412), .X(n26923) );
  nand_x1_sg U70077 ( .A(n22115), .B(n27012), .X(n27160) );
  nand_x1_sg U70078 ( .A(n45369), .B(n45410), .X(n27162) );
  nand_x1_sg U70079 ( .A(n22059), .B(n27257), .X(n27378) );
  nand_x1_sg U70080 ( .A(n45416), .B(n45452), .X(n27380) );
  nand_x1_sg U70081 ( .A(n22015), .B(n27485), .X(n27579) );
  nand_x1_sg U70082 ( .A(n45461), .B(n45498), .X(n27581) );
  nand_x1_sg U70083 ( .A(n21975), .B(n27694), .X(n27761) );
  nand_x1_sg U70084 ( .A(n45510), .B(n45540), .X(n27763) );
  nand_x1_sg U70085 ( .A(n21918), .B(n27755), .X(n27752) );
  nand_x1_sg U70086 ( .A(n45555), .B(n45583), .X(n27754) );
  nand_x1_sg U70087 ( .A(n21877), .B(n27555), .X(n27552) );
  nand_x1_sg U70088 ( .A(n45601), .B(n45625), .X(n27554) );
  nand_x1_sg U70089 ( .A(n21799), .B(n27099), .X(n27096) );
  nand_x1_sg U70090 ( .A(n45690), .B(n45708), .X(n27098) );
  nand_x1_sg U70091 ( .A(n6275), .B(n21508), .X(n21552) );
  nand_x1_sg U70092 ( .A(n46325), .B(n46329), .X(n21554) );
  nand_x1_sg U70093 ( .A(n20940), .B(n20944), .X(n21020) );
  nand_x1_sg U70094 ( .A(n46455), .B(n46469), .X(n21022) );
  nand_x1_sg U70095 ( .A(n20754), .B(n20757), .X(n20799) );
  nand_x1_sg U70096 ( .A(n46405), .B(n42256), .X(n20801) );
  nand_x1_sg U70097 ( .A(n19435), .B(n19439), .X(n19602) );
  nand_x1_sg U70098 ( .A(n46073), .B(n46111), .X(n19604) );
  nand_x1_sg U70099 ( .A(n20086), .B(n20089), .X(n20168) );
  nand_x1_sg U70100 ( .A(n46216), .B(n42209), .X(n20170) );
  nand_x1_sg U70101 ( .A(n19261), .B(n19264), .X(n19371) );
  nand_x1_sg U70102 ( .A(n46071), .B(n42220), .X(n19373) );
  nand_x1_sg U70103 ( .A(n22092), .B(n28204), .X(n28201) );
  nand_x1_sg U70104 ( .A(n45425), .B(n45440), .X(n28203) );
  nand_x1_sg U70105 ( .A(n22025), .B(n28198), .X(n28585) );
  nand_x1_sg U70106 ( .A(n45470), .B(n45483), .X(n28587) );
  nand_x1_sg U70107 ( .A(n21984), .B(n28701), .X(n28770) );
  nand_x1_sg U70108 ( .A(n45516), .B(n45525), .X(n28772) );
  nand_x1_sg U70109 ( .A(n22093), .B(n28877), .X(n28946) );
  nand_x1_sg U70110 ( .A(n45428), .B(n45434), .X(n28948) );
  nand_x1_sg U70111 ( .A(n22026), .B(n29059), .X(n29103) );
  nand_x1_sg U70112 ( .A(n45473), .B(n45477), .X(n29105) );
  nand_x1_sg U70113 ( .A(n22089), .B(n22088), .X(n26918) );
  nand_x1_sg U70114 ( .A(n45414), .B(n45456), .X(n26920) );
  nand_x1_sg U70115 ( .A(n22069), .B(n27018), .X(n27157) );
  nand_x1_sg U70116 ( .A(n45415), .B(n45454), .X(n27159) );
  nand_x1_sg U70117 ( .A(n22012), .B(n27263), .X(n27375) );
  nand_x1_sg U70118 ( .A(n45460), .B(n45500), .X(n27377) );
  nand_x1_sg U70119 ( .A(n21969), .B(n27491), .X(n27576) );
  nand_x1_sg U70120 ( .A(n45509), .B(n45542), .X(n27578) );
  nand_x1_sg U70121 ( .A(n21928), .B(n27700), .X(n27758) );
  nand_x1_sg U70122 ( .A(n45554), .B(n45585), .X(n27760) );
  nand_x1_sg U70123 ( .A(n21872), .B(n27561), .X(n27558) );
  nand_x1_sg U70124 ( .A(n45600), .B(n45627), .X(n27560) );
  nand_x1_sg U70125 ( .A(n21830), .B(n27342), .X(n27339) );
  nand_x1_sg U70126 ( .A(n45669), .B(n45645), .X(n27341) );
  nand_x1_sg U70127 ( .A(n46370), .B(n21515), .X(n21549) );
  nand_x1_sg U70128 ( .A(n46367), .B(n21510), .X(n21551) );
  nand_x1_sg U70129 ( .A(n20761), .B(n20764), .X(n20796) );
  nand_x1_sg U70130 ( .A(n46453), .B(n42257), .X(n20798) );
  nand_x1_sg U70131 ( .A(n19442), .B(n19446), .X(n19599) );
  nand_x1_sg U70132 ( .A(n46118), .B(n46157), .X(n19601) );
  nand_x1_sg U70133 ( .A(n20093), .B(n20096), .X(n20165) );
  nand_x1_sg U70134 ( .A(n46262), .B(n42211), .X(n20167) );
  nand_x1_sg U70135 ( .A(n19268), .B(n19271), .X(n19368) );
  nand_x1_sg U70136 ( .A(n46116), .B(n42216), .X(n19370) );
  nand_x1_sg U70137 ( .A(n22046), .B(n28069), .X(n28066) );
  nand_x1_sg U70138 ( .A(n45469), .B(n45485), .X(n28068) );
  nand_x1_sg U70139 ( .A(n21979), .B(n28063), .X(n28582) );
  nand_x1_sg U70140 ( .A(n45515), .B(n45527), .X(n28584) );
  nand_x1_sg U70141 ( .A(n21938), .B(n28707), .X(n28767) );
  nand_x1_sg U70142 ( .A(n45560), .B(n45570), .X(n28769) );
  nand_x1_sg U70143 ( .A(n22047), .B(n28883), .X(n28943) );
  nand_x1_sg U70144 ( .A(n45472), .B(n45479), .X(n28945) );
  nand_x1_sg U70145 ( .A(n45521), .B(n29066), .X(n29100) );
  nand_x1_sg U70146 ( .A(n45518), .B(n29062), .X(n29102) );
  nand_x1_sg U70147 ( .A(n22043), .B(n22042), .X(n26915) );
  nand_x1_sg U70148 ( .A(n45458), .B(n45504), .X(n26917) );
  nand_x1_sg U70149 ( .A(n22022), .B(n27024), .X(n27154) );
  nand_x1_sg U70150 ( .A(n45459), .B(n45502), .X(n27156) );
  nand_x1_sg U70151 ( .A(n21966), .B(n27269), .X(n27372) );
  nand_x1_sg U70152 ( .A(n45508), .B(n45544), .X(n27374) );
  nand_x1_sg U70153 ( .A(n21922), .B(n27497), .X(n27573) );
  nand_x1_sg U70154 ( .A(n45553), .B(n45587), .X(n27575) );
  nand_x1_sg U70155 ( .A(n21882), .B(n27567), .X(n27564) );
  nand_x1_sg U70156 ( .A(n45599), .B(n45629), .X(n27566) );
  nand_x1_sg U70157 ( .A(n21825), .B(n27348), .X(n27345) );
  nand_x1_sg U70158 ( .A(n45671), .B(n45644), .X(n27347) );
  nand_x1_sg U70159 ( .A(n21783), .B(n27112), .X(n27109) );
  nand_x1_sg U70160 ( .A(n45689), .B(n45712), .X(n27111) );
  nand_x1_sg U70161 ( .A(n6184), .B(n21521), .X(n21546) );
  nand_x1_sg U70162 ( .A(n46414), .B(n46418), .X(n21548) );
  nand_x1_sg U70163 ( .A(n19449), .B(n19453), .X(n19596) );
  nand_x1_sg U70164 ( .A(n46164), .B(n46202), .X(n19598) );
  nand_x1_sg U70165 ( .A(n19275), .B(n19278), .X(n19365) );
  nand_x1_sg U70166 ( .A(n46162), .B(n42221), .X(n19367) );
  nand_x1_sg U70167 ( .A(n21999), .B(n27907), .X(n27904) );
  nand_x1_sg U70168 ( .A(n45514), .B(n45529), .X(n27906) );
  nand_x1_sg U70169 ( .A(n21932), .B(n27901), .X(n28579) );
  nand_x1_sg U70170 ( .A(n45559), .B(n45572), .X(n28581) );
  nand_x1_sg U70171 ( .A(n21891), .B(n28713), .X(n28764) );
  nand_x1_sg U70172 ( .A(n45605), .B(n45614), .X(n28766) );
  nand_x1_sg U70173 ( .A(n22000), .B(n28889), .X(n28940) );
  nand_x1_sg U70174 ( .A(n45517), .B(n45523), .X(n28942) );
  nand_x1_sg U70175 ( .A(n21933), .B(n29072), .X(n29097) );
  nand_x1_sg U70176 ( .A(n45562), .B(n45566), .X(n29099) );
  nand_x1_sg U70177 ( .A(n21996), .B(n21995), .X(n26912) );
  nand_x1_sg U70178 ( .A(n45506), .B(n45548), .X(n26914) );
  nand_x1_sg U70179 ( .A(n21976), .B(n27030), .X(n27151) );
  nand_x1_sg U70180 ( .A(n45507), .B(n45546), .X(n27153) );
  nand_x1_sg U70181 ( .A(n21919), .B(n27275), .X(n27369) );
  nand_x1_sg U70182 ( .A(n45552), .B(n45589), .X(n27371) );
  nand_x1_sg U70183 ( .A(n21876), .B(n27503), .X(n27570) );
  nand_x1_sg U70184 ( .A(n45598), .B(n45631), .X(n27572) );
  nand_x1_sg U70185 ( .A(n21835), .B(n27354), .X(n27351) );
  nand_x1_sg U70186 ( .A(n45673), .B(n45643), .X(n27353) );
  nand_x1_sg U70187 ( .A(n21778), .B(n27118), .X(n27115) );
  nand_x1_sg U70188 ( .A(n45688), .B(n45714), .X(n27117) );
  nand_x1_sg U70189 ( .A(n46465), .B(n21528), .X(n21543) );
  nand_x1_sg U70190 ( .A(n46462), .B(n21523), .X(n21545) );
  nand_x1_sg U70191 ( .A(n19456), .B(n19460), .X(n19593) );
  nand_x1_sg U70192 ( .A(n46209), .B(n46248), .X(n19595) );
  nand_x1_sg U70193 ( .A(n19282), .B(n19285), .X(n19362) );
  nand_x1_sg U70194 ( .A(n46207), .B(n42222), .X(n19364) );
  nand_x1_sg U70195 ( .A(n21953), .B(n27730), .X(n27727) );
  nand_x1_sg U70196 ( .A(n45558), .B(n45574), .X(n27729) );
  nand_x1_sg U70197 ( .A(n21886), .B(n27724), .X(n28576) );
  nand_x1_sg U70198 ( .A(n45604), .B(n45616), .X(n28578) );
  nand_x1_sg U70199 ( .A(n21845), .B(n28719), .X(n28761) );
  nand_x1_sg U70200 ( .A(n45658), .B(n45649), .X(n28763) );
  nand_x1_sg U70201 ( .A(n21954), .B(n28895), .X(n28937) );
  nand_x1_sg U70202 ( .A(n45561), .B(n45568), .X(n28939) );
  nand_x1_sg U70203 ( .A(n45610), .B(n29079), .X(n29094) );
  nand_x1_sg U70204 ( .A(n45607), .B(n29075), .X(n29096) );
  nand_x1_sg U70205 ( .A(n21950), .B(n21949), .X(n26909) );
  nand_x1_sg U70206 ( .A(n45550), .B(n45593), .X(n26911) );
  nand_x1_sg U70207 ( .A(n21929), .B(n27036), .X(n27148) );
  nand_x1_sg U70208 ( .A(n45551), .B(n45591), .X(n27150) );
  nand_x1_sg U70209 ( .A(n21873), .B(n27281), .X(n27366) );
  nand_x1_sg U70210 ( .A(n45597), .B(n45633), .X(n27368) );
  nand_x1_sg U70211 ( .A(n21829), .B(n27360), .X(n27357) );
  nand_x1_sg U70212 ( .A(n45675), .B(n45642), .X(n27359) );
  nand_x1_sg U70213 ( .A(n21788), .B(n27124), .X(n27121) );
  nand_x1_sg U70214 ( .A(n45687), .B(n45716), .X(n27123) );
  nand_x1_sg U70215 ( .A(n6093), .B(n21364), .X(n21361) );
  nand_x1_sg U70216 ( .A(n46500), .B(n46503), .X(n21363) );
  nand_x1_sg U70217 ( .A(n19463), .B(n19467), .X(n19590) );
  nand_x1_sg U70218 ( .A(n46255), .B(n46293), .X(n19592) );
  nand_x1_sg U70219 ( .A(n19289), .B(n19292), .X(n19359) );
  nand_x1_sg U70220 ( .A(n46253), .B(n42223), .X(n19361) );
  nand_x1_sg U70221 ( .A(n21906), .B(n27536), .X(n27533) );
  nand_x1_sg U70222 ( .A(n45603), .B(n45618), .X(n27535) );
  nand_x1_sg U70223 ( .A(n21839), .B(n27530), .X(n28573) );
  nand_x1_sg U70224 ( .A(n45660), .B(n45648), .X(n28575) );
  nand_x1_sg U70225 ( .A(n21798), .B(n28725), .X(n28758) );
  nand_x1_sg U70226 ( .A(n45693), .B(n45702), .X(n28760) );
  nand_x1_sg U70227 ( .A(n21907), .B(n28901), .X(n28934) );
  nand_x1_sg U70228 ( .A(n45606), .B(n45612), .X(n28936) );
  nand_x1_sg U70229 ( .A(n21840), .B(n28928), .X(n28925) );
  nand_x1_sg U70230 ( .A(n45654), .B(n45651), .X(n28927) );
  nand_x1_sg U70231 ( .A(n21903), .B(n21902), .X(n26906) );
  nand_x1_sg U70232 ( .A(n45595), .B(n45637), .X(n26908) );
  nand_x1_sg U70233 ( .A(n21883), .B(n27042), .X(n27145) );
  nand_x1_sg U70234 ( .A(n45596), .B(n45635), .X(n27147) );
  nand_x1_sg U70235 ( .A(n21826), .B(n27287), .X(n27363) );
  nand_x1_sg U70236 ( .A(n45677), .B(n45641), .X(n27365) );
  nand_x1_sg U70237 ( .A(n21782), .B(n27130), .X(n27127) );
  nand_x1_sg U70238 ( .A(n45686), .B(n45718), .X(n27129) );
  nand_x1_sg U70239 ( .A(n6043), .B(n21194), .X(n21191) );
  nand_x1_sg U70240 ( .A(n46542), .B(n46545), .X(n21193) );
  nand_x1_sg U70241 ( .A(n21860), .B(n27323), .X(n27320) );
  nand_x1_sg U70242 ( .A(n45662), .B(n45647), .X(n27322) );
  nand_x1_sg U70243 ( .A(n21792), .B(n27317), .X(n28570) );
  nand_x1_sg U70244 ( .A(n45692), .B(n45704), .X(n28572) );
  nand_x1_sg U70245 ( .A(n21861), .B(n28907), .X(n28931) );
  nand_x1_sg U70246 ( .A(n45656), .B(n45650), .X(n28933) );
  nand_x1_sg U70247 ( .A(n21793), .B(n28749), .X(n28746) );
  nand_x1_sg U70248 ( .A(n45695), .B(n45698), .X(n28748) );
  nand_x1_sg U70249 ( .A(n21857), .B(n21856), .X(n26903) );
  nand_x1_sg U70250 ( .A(n45681), .B(n45639), .X(n26905) );
  nand_x1_sg U70251 ( .A(n21836), .B(n27048), .X(n27142) );
  nand_x1_sg U70252 ( .A(n45679), .B(n45640), .X(n27144) );
  nand_x1_sg U70253 ( .A(n21779), .B(n27136), .X(n27133) );
  nand_x1_sg U70254 ( .A(n45685), .B(n45720), .X(n27135) );
  nand_x1_sg U70255 ( .A(n21813), .B(n27093), .X(n27090) );
  nand_x1_sg U70256 ( .A(n45691), .B(n45706), .X(n27092) );
  nand_x1_sg U70257 ( .A(n21814), .B(n28755), .X(n28752) );
  nand_x1_sg U70258 ( .A(n45694), .B(n45700), .X(n28754) );
  nand_x1_sg U70259 ( .A(n21810), .B(n21809), .X(n26900) );
  nand_x1_sg U70260 ( .A(n45683), .B(n45724), .X(n26902) );
  nand_x1_sg U70261 ( .A(n21789), .B(n27054), .X(n27139) );
  nand_x1_sg U70262 ( .A(n45684), .B(n45722), .X(n27141) );
  nand_x1_sg U70263 ( .A(n20677), .B(n45906), .X(n20832) );
  nand_x1_sg U70264 ( .A(n20680), .B(n42199), .X(n20834) );
  nand_x1_sg U70265 ( .A(n20037), .B(n45896), .X(n20189) );
  nand_x1_sg U70266 ( .A(n20040), .B(n42200), .X(n20191) );
  nand_x1_sg U70267 ( .A(n19233), .B(n45886), .X(n19383) );
  nand_x1_sg U70268 ( .A(n19236), .B(n42217), .X(n19385) );
  nand_x1_sg U70269 ( .A(n6127), .B(n46434), .X(n19160) );
  nand_x1_sg U70270 ( .A(n6131), .B(n42258), .X(n19162) );
  nand_x1_sg U70271 ( .A(n28181), .B(n42153), .X(n28178) );
  nand_x1_sg U70272 ( .A(n28180), .B(n45423), .X(n28179) );
  nand_x1_sg U70273 ( .A(n28186), .B(n42154), .X(n28184) );
  nand_x1_sg U70274 ( .A(n28081), .B(n45467), .X(n28185) );
  nand_x1_sg U70275 ( .A(n28051), .B(n42155), .X(n28049) );
  nand_x1_sg U70276 ( .A(n27919), .B(n45491), .X(n28050) );
  nand_x1_sg U70277 ( .A(n27889), .B(n42156), .X(n27887) );
  nand_x1_sg U70278 ( .A(n27742), .B(n45535), .X(n27888) );
  nand_x1_sg U70279 ( .A(n27712), .B(n42157), .X(n27710) );
  nand_x1_sg U70280 ( .A(n27548), .B(n45580), .X(n27711) );
  nand_x1_sg U70281 ( .A(n27518), .B(n42158), .X(n27516) );
  nand_x1_sg U70282 ( .A(n27335), .B(n45624), .X(n27517) );
  nand_x1_sg U70283 ( .A(n27305), .B(n42228), .X(n27303) );
  nand_x1_sg U70284 ( .A(n27105), .B(n45668), .X(n27304) );
  nand_x1_sg U70285 ( .A(n20863), .B(n45955), .X(n21053) );
  nand_x1_sg U70286 ( .A(n20867), .B(n45969), .X(n21055) );
  nand_x1_sg U70287 ( .A(n20220), .B(n45946), .X(n20344) );
  nand_x1_sg U70288 ( .A(n20224), .B(n45972), .X(n20346) );
  nand_x1_sg U70289 ( .A(n19414), .B(n45937), .X(n19611) );
  nand_x1_sg U70290 ( .A(n19418), .B(n45975), .X(n19613) );
  nand_x1_sg U70291 ( .A(n27811), .B(n45039), .X(n27809) );
  nor_x1_sg U70292 ( .A(n45039), .B(n27811), .X(n27810) );
  nand_x1_sg U70293 ( .A(n27817), .B(n45083), .X(n27815) );
  nor_x1_sg U70294 ( .A(n45083), .B(n27817), .X(n27816) );
  nand_x1_sg U70295 ( .A(n27994), .B(n45128), .X(n27992) );
  nor_x1_sg U70296 ( .A(n45128), .B(n27994), .X(n27993) );
  nand_x1_sg U70297 ( .A(n28000), .B(n45173), .X(n27998) );
  nor_x1_sg U70298 ( .A(n45173), .B(n28000), .X(n27999) );
  nand_x1_sg U70299 ( .A(n28006), .B(n45219), .X(n28004) );
  nor_x1_sg U70300 ( .A(n45219), .B(n28006), .X(n28005) );
  nand_x1_sg U70301 ( .A(n28012), .B(n45264), .X(n28010) );
  nor_x1_sg U70302 ( .A(n45264), .B(n28012), .X(n28011) );
  nand_x1_sg U70303 ( .A(n28018), .B(n45309), .X(n28016) );
  nor_x1_sg U70304 ( .A(n45309), .B(n28018), .X(n28017) );
  nand_x1_sg U70305 ( .A(n28024), .B(n45354), .X(n28022) );
  nor_x1_sg U70306 ( .A(n45354), .B(n28024), .X(n28023) );
  nand_x1_sg U70307 ( .A(n28030), .B(n45400), .X(n28028) );
  nor_x1_sg U70308 ( .A(n45400), .B(n28030), .X(n28029) );
  nand_x1_sg U70309 ( .A(n28898), .B(n45612), .X(n28896) );
  nor_x1_sg U70310 ( .A(n45612), .B(n28898), .X(n28897) );
  nand_x1_sg U70311 ( .A(n28886), .B(n45523), .X(n28884) );
  nor_x1_sg U70312 ( .A(n45523), .B(n28886), .X(n28885) );
  nand_x1_sg U70313 ( .A(n28874), .B(n45434), .X(n28872) );
  nor_x1_sg U70314 ( .A(n45434), .B(n28874), .X(n28873) );
  nand_x1_sg U70315 ( .A(n28862), .B(n45343), .X(n28860) );
  nor_x1_sg U70316 ( .A(n45343), .B(n28862), .X(n28861) );
  nand_x1_sg U70317 ( .A(n28850), .B(n45253), .X(n28848) );
  nor_x1_sg U70318 ( .A(n45253), .B(n28850), .X(n28849) );
  nand_x1_sg U70319 ( .A(n28838), .B(n45162), .X(n28836) );
  nor_x1_sg U70320 ( .A(n45162), .B(n28838), .X(n28837) );
  nand_x1_sg U70321 ( .A(n28826), .B(n45070), .X(n28824) );
  nor_x1_sg U70322 ( .A(n45070), .B(n28826), .X(n28825) );
  nand_x1_sg U70323 ( .A(n27625), .B(n45041), .X(n27623) );
  nor_x1_sg U70324 ( .A(n45041), .B(n27625), .X(n27624) );
  nand_x1_sg U70325 ( .A(n28632), .B(n45029), .X(n28630) );
  nor_x1_sg U70326 ( .A(n45029), .B(n28632), .X(n28631) );
  nand_x1_sg U70327 ( .A(n27422), .B(n45043), .X(n27420) );
  nor_x1_sg U70328 ( .A(n45043), .B(n27422), .X(n27421) );
  nand_x1_sg U70329 ( .A(n27631), .B(n45085), .X(n27629) );
  nor_x1_sg U70330 ( .A(n45085), .B(n27631), .X(n27630) );
  nand_x1_sg U70331 ( .A(n27823), .B(n45130), .X(n27821) );
  nor_x1_sg U70332 ( .A(n45130), .B(n27823), .X(n27822) );
  nand_x1_sg U70333 ( .A(n28471), .B(n45031), .X(n28469) );
  nor_x1_sg U70334 ( .A(n45031), .B(n28471), .X(n28470) );
  nand_x1_sg U70335 ( .A(n28638), .B(n45072), .X(n28636) );
  nor_x1_sg U70336 ( .A(n45072), .B(n28638), .X(n28637) );
  nand_x1_sg U70337 ( .A(n28991), .B(n45025), .X(n28989) );
  nor_x1_sg U70338 ( .A(n45025), .B(n28991), .X(n28990) );
  nand_x1_sg U70339 ( .A(n27200), .B(n45045), .X(n27198) );
  nor_x1_sg U70340 ( .A(n45045), .B(n27200), .X(n27199) );
  nand_x1_sg U70341 ( .A(n27428), .B(n45087), .X(n27426) );
  nor_x1_sg U70342 ( .A(n45087), .B(n27428), .X(n27427) );
  nand_x1_sg U70343 ( .A(n27637), .B(n45132), .X(n27635) );
  nor_x1_sg U70344 ( .A(n45132), .B(n27637), .X(n27636) );
  nand_x1_sg U70345 ( .A(n27829), .B(n45175), .X(n27827) );
  nor_x1_sg U70346 ( .A(n45175), .B(n27829), .X(n27828) );
  nand_x1_sg U70347 ( .A(n28477), .B(n45074), .X(n28475) );
  nor_x1_sg U70348 ( .A(n45074), .B(n28477), .X(n28476) );
  nand_x1_sg U70349 ( .A(n28644), .B(n45119), .X(n28642) );
  nor_x1_sg U70350 ( .A(n45119), .B(n28644), .X(n28643) );
  nand_x1_sg U70351 ( .A(n27206), .B(n45089), .X(n27204) );
  nor_x1_sg U70352 ( .A(n45089), .B(n27206), .X(n27205) );
  nand_x1_sg U70353 ( .A(n27434), .B(n45134), .X(n27432) );
  nor_x1_sg U70354 ( .A(n45134), .B(n27434), .X(n27433) );
  nand_x1_sg U70355 ( .A(n27643), .B(n45177), .X(n27641) );
  nor_x1_sg U70356 ( .A(n45177), .B(n27643), .X(n27642) );
  nand_x1_sg U70357 ( .A(n27835), .B(n45221), .X(n27833) );
  nor_x1_sg U70358 ( .A(n45221), .B(n27835), .X(n27834) );
  nand_x1_sg U70359 ( .A(n28483), .B(n45121), .X(n28481) );
  nor_x1_sg U70360 ( .A(n45121), .B(n28483), .X(n28482) );
  nand_x1_sg U70361 ( .A(n28650), .B(n45164), .X(n28648) );
  nor_x1_sg U70362 ( .A(n45164), .B(n28650), .X(n28649) );
  nand_x1_sg U70363 ( .A(n29004), .B(n45115), .X(n29002) );
  nor_x1_sg U70364 ( .A(n45115), .B(n29004), .X(n29003) );
  nand_x1_sg U70365 ( .A(n27212), .B(n45136), .X(n27210) );
  nor_x1_sg U70366 ( .A(n45136), .B(n27212), .X(n27211) );
  nand_x1_sg U70367 ( .A(n27440), .B(n45179), .X(n27438) );
  nor_x1_sg U70368 ( .A(n45179), .B(n27440), .X(n27439) );
  nand_x1_sg U70369 ( .A(n27649), .B(n45223), .X(n27647) );
  nor_x1_sg U70370 ( .A(n45223), .B(n27649), .X(n27648) );
  nand_x1_sg U70371 ( .A(n27841), .B(n45266), .X(n27839) );
  nor_x1_sg U70372 ( .A(n45266), .B(n27841), .X(n27840) );
  nand_x1_sg U70373 ( .A(n28489), .B(n45166), .X(n28487) );
  nor_x1_sg U70374 ( .A(n45166), .B(n28489), .X(n28488) );
  nand_x1_sg U70375 ( .A(n28656), .B(n45210), .X(n28654) );
  nor_x1_sg U70376 ( .A(n45210), .B(n28656), .X(n28655) );
  nand_x1_sg U70377 ( .A(n27218), .B(n45181), .X(n27216) );
  nor_x1_sg U70378 ( .A(n45181), .B(n27218), .X(n27217) );
  nand_x1_sg U70379 ( .A(n27446), .B(n45225), .X(n27444) );
  nor_x1_sg U70380 ( .A(n45225), .B(n27446), .X(n27445) );
  nand_x1_sg U70381 ( .A(n27655), .B(n45268), .X(n27653) );
  nor_x1_sg U70382 ( .A(n45268), .B(n27655), .X(n27654) );
  nand_x1_sg U70383 ( .A(n27847), .B(n45311), .X(n27845) );
  nor_x1_sg U70384 ( .A(n45311), .B(n27847), .X(n27846) );
  nand_x1_sg U70385 ( .A(n28495), .B(n45212), .X(n28493) );
  nor_x1_sg U70386 ( .A(n45212), .B(n28495), .X(n28494) );
  nand_x1_sg U70387 ( .A(n28662), .B(n45255), .X(n28660) );
  nor_x1_sg U70388 ( .A(n45255), .B(n28662), .X(n28661) );
  nand_x1_sg U70389 ( .A(n29017), .B(n45206), .X(n29015) );
  nor_x1_sg U70390 ( .A(n45206), .B(n29017), .X(n29016) );
  nand_x1_sg U70391 ( .A(n27224), .B(n45227), .X(n27222) );
  nor_x1_sg U70392 ( .A(n45227), .B(n27224), .X(n27223) );
  nand_x1_sg U70393 ( .A(n27452), .B(n45270), .X(n27450) );
  nor_x1_sg U70394 ( .A(n45270), .B(n27452), .X(n27451) );
  nand_x1_sg U70395 ( .A(n27661), .B(n45313), .X(n27659) );
  nor_x1_sg U70396 ( .A(n45313), .B(n27661), .X(n27660) );
  nand_x1_sg U70397 ( .A(n27853), .B(n45356), .X(n27851) );
  nor_x1_sg U70398 ( .A(n45356), .B(n27853), .X(n27852) );
  nand_x1_sg U70399 ( .A(n28501), .B(n45257), .X(n28499) );
  nor_x1_sg U70400 ( .A(n45257), .B(n28501), .X(n28500) );
  nand_x1_sg U70401 ( .A(n28668), .B(n45300), .X(n28666) );
  nor_x1_sg U70402 ( .A(n45300), .B(n28668), .X(n28667) );
  nand_x1_sg U70403 ( .A(n27230), .B(n45272), .X(n27228) );
  nor_x1_sg U70404 ( .A(n45272), .B(n27230), .X(n27229) );
  nand_x1_sg U70405 ( .A(n27458), .B(n45315), .X(n27456) );
  nor_x1_sg U70406 ( .A(n45315), .B(n27458), .X(n27457) );
  nand_x1_sg U70407 ( .A(n27667), .B(n45358), .X(n27665) );
  nor_x1_sg U70408 ( .A(n45358), .B(n27667), .X(n27666) );
  nand_x1_sg U70409 ( .A(n27859), .B(n45402), .X(n27857) );
  nor_x1_sg U70410 ( .A(n45402), .B(n27859), .X(n27858) );
  nand_x1_sg U70411 ( .A(n28036), .B(n45444), .X(n28034) );
  nor_x1_sg U70412 ( .A(n45444), .B(n28036), .X(n28035) );
  nand_x1_sg U70413 ( .A(n28507), .B(n45302), .X(n28505) );
  nor_x1_sg U70414 ( .A(n45302), .B(n28507), .X(n28506) );
  nand_x1_sg U70415 ( .A(n28674), .B(n45345), .X(n28672) );
  nor_x1_sg U70416 ( .A(n45345), .B(n28674), .X(n28673) );
  nand_x1_sg U70417 ( .A(n29030), .B(n45296), .X(n29028) );
  nor_x1_sg U70418 ( .A(n45296), .B(n29030), .X(n29029) );
  nand_x1_sg U70419 ( .A(n27236), .B(n45317), .X(n27234) );
  nor_x1_sg U70420 ( .A(n45317), .B(n27236), .X(n27235) );
  nand_x1_sg U70421 ( .A(n27464), .B(n45360), .X(n27462) );
  nor_x1_sg U70422 ( .A(n45360), .B(n27464), .X(n27463) );
  nand_x1_sg U70423 ( .A(n27673), .B(n45404), .X(n27671) );
  nor_x1_sg U70424 ( .A(n45404), .B(n27673), .X(n27672) );
  nand_x1_sg U70425 ( .A(n27865), .B(n45446), .X(n27863) );
  nor_x1_sg U70426 ( .A(n45446), .B(n27865), .X(n27864) );
  nand_x1_sg U70427 ( .A(n28042), .B(n45492), .X(n28040) );
  nor_x1_sg U70428 ( .A(n45492), .B(n28042), .X(n28041) );
  nand_x1_sg U70429 ( .A(n28513), .B(n45347), .X(n28511) );
  nor_x1_sg U70430 ( .A(n45347), .B(n28513), .X(n28512) );
  nand_x1_sg U70431 ( .A(n28680), .B(n45391), .X(n28678) );
  nor_x1_sg U70432 ( .A(n45391), .B(n28680), .X(n28679) );
  nand_x1_sg U70433 ( .A(n27242), .B(n45362), .X(n27240) );
  nor_x1_sg U70434 ( .A(n45362), .B(n27242), .X(n27241) );
  nand_x1_sg U70435 ( .A(n27470), .B(n45406), .X(n27468) );
  nor_x1_sg U70436 ( .A(n45406), .B(n27470), .X(n27469) );
  nand_x1_sg U70437 ( .A(n27679), .B(n45448), .X(n27677) );
  nor_x1_sg U70438 ( .A(n45448), .B(n27679), .X(n27678) );
  nand_x1_sg U70439 ( .A(n27871), .B(n45494), .X(n27869) );
  nor_x1_sg U70440 ( .A(n45494), .B(n27871), .X(n27870) );
  nand_x1_sg U70441 ( .A(n28048), .B(n45536), .X(n28046) );
  nor_x1_sg U70442 ( .A(n45536), .B(n28048), .X(n28047) );
  nand_x1_sg U70443 ( .A(n28428), .B(n45393), .X(n28426) );
  nor_x1_sg U70444 ( .A(n45393), .B(n28428), .X(n28427) );
  nand_x1_sg U70445 ( .A(n28686), .B(n45436), .X(n28684) );
  nor_x1_sg U70446 ( .A(n45436), .B(n28686), .X(n28685) );
  nand_x1_sg U70447 ( .A(n29043), .B(n45387), .X(n29041) );
  nor_x1_sg U70448 ( .A(n45387), .B(n29043), .X(n29042) );
  nand_x1_sg U70449 ( .A(n27248), .B(n45408), .X(n27246) );
  nor_x1_sg U70450 ( .A(n45408), .B(n27248), .X(n27247) );
  nand_x1_sg U70451 ( .A(n27476), .B(n45450), .X(n27474) );
  nor_x1_sg U70452 ( .A(n45450), .B(n27476), .X(n27475) );
  nand_x1_sg U70453 ( .A(n27685), .B(n45496), .X(n27683) );
  nor_x1_sg U70454 ( .A(n45496), .B(n27685), .X(n27684) );
  nand_x1_sg U70455 ( .A(n27877), .B(n45538), .X(n27875) );
  nor_x1_sg U70456 ( .A(n45538), .B(n27877), .X(n27876) );
  nand_x1_sg U70457 ( .A(n27886), .B(n45581), .X(n27884) );
  nor_x1_sg U70458 ( .A(n45581), .B(n27886), .X(n27885) );
  nand_x1_sg U70459 ( .A(n28324), .B(n45438), .X(n28322) );
  nor_x1_sg U70460 ( .A(n45438), .B(n28324), .X(n28323) );
  nand_x1_sg U70461 ( .A(n28692), .B(n45481), .X(n28690) );
  nor_x1_sg U70462 ( .A(n45481), .B(n28692), .X(n28691) );
  nand_x1_sg U70463 ( .A(n27254), .B(n45452), .X(n27252) );
  nor_x1_sg U70464 ( .A(n45452), .B(n27254), .X(n27253) );
  nand_x1_sg U70465 ( .A(n27482), .B(n45498), .X(n27480) );
  nor_x1_sg U70466 ( .A(n45498), .B(n27482), .X(n27481) );
  nand_x1_sg U70467 ( .A(n27691), .B(n45540), .X(n27689) );
  nor_x1_sg U70468 ( .A(n45540), .B(n27691), .X(n27690) );
  nand_x1_sg U70469 ( .A(n27883), .B(n45583), .X(n27881) );
  nor_x1_sg U70470 ( .A(n45583), .B(n27883), .X(n27882) );
  nand_x1_sg U70471 ( .A(n27709), .B(n45625), .X(n27707) );
  nor_x1_sg U70472 ( .A(n45625), .B(n27709), .X(n27708) );
  nand_x1_sg U70473 ( .A(n28195), .B(n45483), .X(n28193) );
  nor_x1_sg U70474 ( .A(n45483), .B(n28195), .X(n28194) );
  nand_x1_sg U70475 ( .A(n28698), .B(n45525), .X(n28696) );
  nor_x1_sg U70476 ( .A(n45525), .B(n28698), .X(n28697) );
  nand_x1_sg U70477 ( .A(n29056), .B(n45477), .X(n29054) );
  nor_x1_sg U70478 ( .A(n45477), .B(n29056), .X(n29055) );
  nand_x1_sg U70479 ( .A(n27260), .B(n45500), .X(n27258) );
  nor_x1_sg U70480 ( .A(n45500), .B(n27260), .X(n27259) );
  nand_x1_sg U70481 ( .A(n27488), .B(n45542), .X(n27486) );
  nor_x1_sg U70482 ( .A(n45542), .B(n27488), .X(n27487) );
  nand_x1_sg U70483 ( .A(n27697), .B(n45585), .X(n27695) );
  nor_x1_sg U70484 ( .A(n45585), .B(n27697), .X(n27696) );
  nand_x1_sg U70485 ( .A(n27706), .B(n45627), .X(n27704) );
  nor_x1_sg U70486 ( .A(n45627), .B(n27706), .X(n27705) );
  nand_x1_sg U70487 ( .A(n27515), .B(n45669), .X(n27513) );
  nor_x1_sg U70488 ( .A(n45669), .B(n27515), .X(n27514) );
  nand_x1_sg U70489 ( .A(n27078), .B(n45751), .X(n27076) );
  nor_x1_sg U70490 ( .A(n45751), .B(n27078), .X(n27077) );
  nand_x1_sg U70491 ( .A(n28060), .B(n45527), .X(n28058) );
  nor_x1_sg U70492 ( .A(n45527), .B(n28060), .X(n28059) );
  nand_x1_sg U70493 ( .A(n28704), .B(n45570), .X(n28702) );
  nor_x1_sg U70494 ( .A(n45570), .B(n28704), .X(n28703) );
  nand_x1_sg U70495 ( .A(n27266), .B(n45544), .X(n27264) );
  nor_x1_sg U70496 ( .A(n45544), .B(n27266), .X(n27265) );
  nand_x1_sg U70497 ( .A(n27494), .B(n45587), .X(n27492) );
  nor_x1_sg U70498 ( .A(n45587), .B(n27494), .X(n27493) );
  nand_x1_sg U70499 ( .A(n27703), .B(n45629), .X(n27701) );
  nor_x1_sg U70500 ( .A(n45629), .B(n27703), .X(n27702) );
  nand_x1_sg U70501 ( .A(n27512), .B(n45671), .X(n27510) );
  nor_x1_sg U70502 ( .A(n45671), .B(n27512), .X(n27511) );
  nand_x1_sg U70503 ( .A(n27302), .B(n45712), .X(n27300) );
  nor_x1_sg U70504 ( .A(n45712), .B(n27302), .X(n27301) );
  nand_x1_sg U70505 ( .A(n27075), .B(n45753), .X(n27073) );
  nand_x1_sg U70506 ( .A(n26851), .B(n45711), .X(n27074) );
  nand_x1_sg U70507 ( .A(n27898), .B(n45572), .X(n27896) );
  nor_x1_sg U70508 ( .A(n45572), .B(n27898), .X(n27897) );
  nand_x1_sg U70509 ( .A(n28710), .B(n45614), .X(n28708) );
  nor_x1_sg U70510 ( .A(n45614), .B(n28710), .X(n28709) );
  nand_x1_sg U70511 ( .A(n29069), .B(n45566), .X(n29067) );
  nor_x1_sg U70512 ( .A(n45566), .B(n29069), .X(n29068) );
  nand_x1_sg U70513 ( .A(n27272), .B(n45589), .X(n27270) );
  nor_x1_sg U70514 ( .A(n45589), .B(n27272), .X(n27271) );
  nand_x1_sg U70515 ( .A(n27500), .B(n45631), .X(n27498) );
  nor_x1_sg U70516 ( .A(n45631), .B(n27500), .X(n27499) );
  nand_x1_sg U70517 ( .A(n27509), .B(n45673), .X(n27507) );
  nor_x1_sg U70518 ( .A(n45673), .B(n27509), .X(n27508) );
  nand_x1_sg U70519 ( .A(n27299), .B(n45714), .X(n27297) );
  nor_x1_sg U70520 ( .A(n45714), .B(n27299), .X(n27298) );
  nand_x1_sg U70521 ( .A(n27072), .B(n45755), .X(n27070) );
  nor_x1_sg U70522 ( .A(n45755), .B(n27072), .X(n27071) );
  nand_x1_sg U70523 ( .A(n27721), .B(n45616), .X(n27719) );
  nor_x1_sg U70524 ( .A(n45616), .B(n27721), .X(n27720) );
  nand_x1_sg U70525 ( .A(n28716), .B(n45658), .X(n28714) );
  nor_x1_sg U70526 ( .A(n45658), .B(n28716), .X(n28715) );
  nand_x1_sg U70527 ( .A(n27278), .B(n45633), .X(n27276) );
  nor_x1_sg U70528 ( .A(n45633), .B(n27278), .X(n27277) );
  nand_x1_sg U70529 ( .A(n27506), .B(n45675), .X(n27504) );
  nor_x1_sg U70530 ( .A(n45675), .B(n27506), .X(n27505) );
  nand_x1_sg U70531 ( .A(n27296), .B(n45716), .X(n27294) );
  nor_x1_sg U70532 ( .A(n45716), .B(n27296), .X(n27295) );
  nand_x1_sg U70533 ( .A(n27069), .B(n45757), .X(n27067) );
  nor_x1_sg U70534 ( .A(n45757), .B(n27069), .X(n27068) );
  nand_x1_sg U70535 ( .A(n27527), .B(n45660), .X(n27525) );
  nor_x1_sg U70536 ( .A(n45660), .B(n27527), .X(n27526) );
  nand_x1_sg U70537 ( .A(n28722), .B(n45702), .X(n28720) );
  nor_x1_sg U70538 ( .A(n45702), .B(n28722), .X(n28721) );
  nand_x1_sg U70539 ( .A(n29082), .B(n45654), .X(n29080) );
  nor_x1_sg U70540 ( .A(n45654), .B(n29082), .X(n29081) );
  nand_x1_sg U70541 ( .A(n27284), .B(n45677), .X(n27282) );
  nor_x1_sg U70542 ( .A(n45677), .B(n27284), .X(n27283) );
  nand_x1_sg U70543 ( .A(n27293), .B(n45718), .X(n27291) );
  nor_x1_sg U70544 ( .A(n45718), .B(n27293), .X(n27292) );
  nand_x1_sg U70545 ( .A(n27066), .B(n45759), .X(n27064) );
  nor_x1_sg U70546 ( .A(n45759), .B(n27066), .X(n27065) );
  nand_x1_sg U70547 ( .A(n27314), .B(n45704), .X(n27312) );
  nor_x1_sg U70548 ( .A(n45704), .B(n27314), .X(n27313) );
  nand_x1_sg U70549 ( .A(n28728), .B(n45745), .X(n28726) );
  nor_x1_sg U70550 ( .A(n45745), .B(n28728), .X(n28727) );
  nand_x1_sg U70551 ( .A(n28913), .B(n45698), .X(n28911) );
  nor_x1_sg U70552 ( .A(n45698), .B(n28913), .X(n28912) );
  nand_x1_sg U70553 ( .A(n27290), .B(n45720), .X(n27288) );
  nor_x1_sg U70554 ( .A(n45720), .B(n27290), .X(n27289) );
  nand_x1_sg U70555 ( .A(n27063), .B(n45761), .X(n27061) );
  nor_x1_sg U70556 ( .A(n45761), .B(n27063), .X(n27062) );
  nand_x1_sg U70557 ( .A(n27084), .B(n45747), .X(n27082) );
  nor_x1_sg U70558 ( .A(n45747), .B(n27084), .X(n27083) );
  nand_x1_sg U70559 ( .A(n28734), .B(n45741), .X(n28732) );
  nor_x1_sg U70560 ( .A(n45741), .B(n28734), .X(n28733) );
  nand_x1_sg U70561 ( .A(n27060), .B(n45763), .X(n27058) );
  nor_x1_sg U70562 ( .A(n45763), .B(n27060), .X(n27059) );
  nand_x1_sg U70563 ( .A(n27081), .B(n45749), .X(n27079) );
  nor_x1_sg U70564 ( .A(n45749), .B(n27081), .X(n27080) );
  nand_x1_sg U70565 ( .A(n28731), .B(n45743), .X(n28729) );
  nor_x1_sg U70566 ( .A(n45743), .B(n28731), .X(n28730) );
  nand_x1_sg U70567 ( .A(n27057), .B(n45765), .X(n27055) );
  nor_x1_sg U70568 ( .A(n45765), .B(n27057), .X(n27056) );
  nand_x1_sg U70569 ( .A(n27311), .B(n45706), .X(n27309) );
  nor_x1_sg U70570 ( .A(n45706), .B(n27311), .X(n27310) );
  nand_x1_sg U70571 ( .A(n28910), .B(n45700), .X(n28908) );
  nor_x1_sg U70572 ( .A(n45700), .B(n28910), .X(n28909) );
  nand_x1_sg U70573 ( .A(n27051), .B(n45722), .X(n27049) );
  nor_x1_sg U70574 ( .A(n45722), .B(n27051), .X(n27050) );
  nand_x1_sg U70575 ( .A(n27524), .B(n45662), .X(n27522) );
  nor_x1_sg U70576 ( .A(n45662), .B(n27524), .X(n27523) );
  nand_x1_sg U70577 ( .A(n28904), .B(n45656), .X(n28902) );
  nor_x1_sg U70578 ( .A(n45656), .B(n28904), .X(n28903) );
  nand_x1_sg U70579 ( .A(n27045), .B(n45679), .X(n27043) );
  nor_x1_sg U70580 ( .A(n45679), .B(n27045), .X(n27044) );
  nand_x1_sg U70581 ( .A(n27718), .B(n45618), .X(n27716) );
  nor_x1_sg U70582 ( .A(n45618), .B(n27718), .X(n27717) );
  nand_x1_sg U70583 ( .A(n27039), .B(n45635), .X(n27037) );
  nor_x1_sg U70584 ( .A(n45635), .B(n27039), .X(n27038) );
  nand_x1_sg U70585 ( .A(n27895), .B(n45574), .X(n27893) );
  nor_x1_sg U70586 ( .A(n45574), .B(n27895), .X(n27894) );
  nand_x1_sg U70587 ( .A(n28892), .B(n45568), .X(n28890) );
  nor_x1_sg U70588 ( .A(n45568), .B(n28892), .X(n28891) );
  nand_x1_sg U70589 ( .A(n27033), .B(n45591), .X(n27031) );
  nor_x1_sg U70590 ( .A(n45591), .B(n27033), .X(n27032) );
  nand_x1_sg U70591 ( .A(n28057), .B(n45529), .X(n28055) );
  nor_x1_sg U70592 ( .A(n45529), .B(n28057), .X(n28056) );
  nand_x1_sg U70593 ( .A(n27027), .B(n45546), .X(n27025) );
  nor_x1_sg U70594 ( .A(n45546), .B(n27027), .X(n27026) );
  nand_x1_sg U70595 ( .A(n28192), .B(n45485), .X(n28190) );
  nor_x1_sg U70596 ( .A(n45485), .B(n28192), .X(n28191) );
  nand_x1_sg U70597 ( .A(n28880), .B(n45479), .X(n28878) );
  nor_x1_sg U70598 ( .A(n45479), .B(n28880), .X(n28879) );
  nand_x1_sg U70599 ( .A(n27021), .B(n45502), .X(n27019) );
  nor_x1_sg U70600 ( .A(n45502), .B(n27021), .X(n27020) );
  nand_x1_sg U70601 ( .A(n28321), .B(n45440), .X(n28319) );
  nor_x1_sg U70602 ( .A(n45440), .B(n28321), .X(n28320) );
  nand_x1_sg U70603 ( .A(n27015), .B(n45454), .X(n27013) );
  nor_x1_sg U70604 ( .A(n45454), .B(n27015), .X(n27014) );
  nand_x1_sg U70605 ( .A(n28425), .B(n45395), .X(n28423) );
  nor_x1_sg U70606 ( .A(n45395), .B(n28425), .X(n28424) );
  nand_x1_sg U70607 ( .A(n28868), .B(n45389), .X(n28866) );
  nor_x1_sg U70608 ( .A(n45389), .B(n28868), .X(n28867) );
  nand_x1_sg U70609 ( .A(n27009), .B(n45410), .X(n27007) );
  nor_x1_sg U70610 ( .A(n45410), .B(n27009), .X(n27008) );
  nand_x1_sg U70611 ( .A(n28419), .B(n45349), .X(n28417) );
  nor_x1_sg U70612 ( .A(n45349), .B(n28419), .X(n28418) );
  nand_x1_sg U70613 ( .A(n27003), .B(n45364), .X(n27001) );
  nor_x1_sg U70614 ( .A(n45364), .B(n27003), .X(n27002) );
  nand_x1_sg U70615 ( .A(n28413), .B(n45304), .X(n28411) );
  nor_x1_sg U70616 ( .A(n45304), .B(n28413), .X(n28412) );
  nand_x1_sg U70617 ( .A(n28856), .B(n45298), .X(n28854) );
  nor_x1_sg U70618 ( .A(n45298), .B(n28856), .X(n28855) );
  nand_x1_sg U70619 ( .A(n26997), .B(n45319), .X(n26995) );
  nor_x1_sg U70620 ( .A(n45319), .B(n26997), .X(n26996) );
  nand_x1_sg U70621 ( .A(n28407), .B(n45259), .X(n28405) );
  nor_x1_sg U70622 ( .A(n45259), .B(n28407), .X(n28406) );
  nand_x1_sg U70623 ( .A(n26991), .B(n45274), .X(n26989) );
  nor_x1_sg U70624 ( .A(n45274), .B(n26991), .X(n26990) );
  nand_x1_sg U70625 ( .A(n28401), .B(n45214), .X(n28399) );
  nor_x1_sg U70626 ( .A(n45214), .B(n28401), .X(n28400) );
  nand_x1_sg U70627 ( .A(n28844), .B(n45208), .X(n28842) );
  nor_x1_sg U70628 ( .A(n45208), .B(n28844), .X(n28843) );
  nand_x1_sg U70629 ( .A(n26985), .B(n45229), .X(n26983) );
  nor_x1_sg U70630 ( .A(n45229), .B(n26985), .X(n26984) );
  nand_x1_sg U70631 ( .A(n28395), .B(n45168), .X(n28393) );
  nor_x1_sg U70632 ( .A(n45168), .B(n28395), .X(n28394) );
  nand_x1_sg U70633 ( .A(n26979), .B(n45183), .X(n26977) );
  nor_x1_sg U70634 ( .A(n45183), .B(n26979), .X(n26978) );
  nand_x1_sg U70635 ( .A(n28389), .B(n45123), .X(n28387) );
  nor_x1_sg U70636 ( .A(n45123), .B(n28389), .X(n28388) );
  nand_x1_sg U70637 ( .A(n28832), .B(n45117), .X(n28830) );
  nor_x1_sg U70638 ( .A(n45117), .B(n28832), .X(n28831) );
  nand_x1_sg U70639 ( .A(n26973), .B(n45138), .X(n26971) );
  nor_x1_sg U70640 ( .A(n45138), .B(n26973), .X(n26972) );
  nand_x1_sg U70641 ( .A(n28383), .B(n45076), .X(n28381) );
  nor_x1_sg U70642 ( .A(n45076), .B(n28383), .X(n28382) );
  nand_x1_sg U70643 ( .A(n26967), .B(n45091), .X(n26965) );
  nor_x1_sg U70644 ( .A(n45091), .B(n26967), .X(n26966) );
  nand_x1_sg U70645 ( .A(n28377), .B(n45033), .X(n28375) );
  nor_x1_sg U70646 ( .A(n45033), .B(n28377), .X(n28376) );
  nand_x1_sg U70647 ( .A(n28820), .B(n45027), .X(n28818) );
  nor_x1_sg U70648 ( .A(n45027), .B(n28820), .X(n28819) );
  nand_x1_sg U70649 ( .A(n26961), .B(n45047), .X(n26959) );
  nor_x1_sg U70650 ( .A(n45047), .B(n26961), .X(n26960) );
  nand_x1_sg U70651 ( .A(n21181), .B(n46583), .X(n21180) );
  nor_x1_sg U70652 ( .A(n21181), .B(n46583), .X(n21182) );
  nand_x1_sg U70653 ( .A(n28736), .B(n45739), .X(n28735) );
  nor_x1_sg U70654 ( .A(n28736), .B(n45739), .X(n28737) );
  nand_x1_sg U70655 ( .A(n7474), .B(n40314), .X(n7472) );
  nor_x1_sg U70656 ( .A(n6030), .B(n46571), .X(n6029) );
  nor_x1_sg U70657 ( .A(n6032), .B(n46570), .X(n6030) );
  nand_x1_sg U70658 ( .A(n46570), .B(n6032), .X(n6031) );
  nor_x1_sg U70659 ( .A(n7829), .B(n22992), .X(n22995) );
  nor_x1_sg U70660 ( .A(n8647), .B(n23272), .X(n23275) );
  nor_x1_sg U70661 ( .A(n9467), .B(n23551), .X(n23554) );
  nor_x1_sg U70662 ( .A(n10286), .B(n23830), .X(n23833) );
  nor_x1_sg U70663 ( .A(n11105), .B(n24109), .X(n24112) );
  nor_x1_sg U70664 ( .A(n11924), .B(n24388), .X(n24391) );
  nor_x1_sg U70665 ( .A(n12743), .B(n24666), .X(n24669) );
  nor_x1_sg U70666 ( .A(n13562), .B(n24945), .X(n24948) );
  nor_x1_sg U70667 ( .A(n14381), .B(n25224), .X(n25227) );
  nor_x1_sg U70668 ( .A(n15200), .B(n25503), .X(n25506) );
  nor_x1_sg U70669 ( .A(n16019), .B(n25780), .X(n25783) );
  nor_x1_sg U70670 ( .A(n17657), .B(n26340), .X(n26343) );
  nor_x1_sg U70671 ( .A(n18478), .B(n26618), .X(n26621) );
  nor_x1_sg U70672 ( .A(n6709), .B(n41277), .X(n6707) );
  nor_x1_sg U70673 ( .A(n6710), .B(n6711), .X(n6709) );
  nor_x1_sg U70674 ( .A(n6713), .B(n41530), .X(n6710) );
  nor_x1_sg U70675 ( .A(n6712), .B(n45867), .X(n6711) );
  nand_x1_sg U70676 ( .A(n39352), .B(n40686), .X(n8346) );
  nand_x1_sg U70677 ( .A(n39351), .B(n40694), .X(n9164) );
  nand_x1_sg U70678 ( .A(n39353), .B(n40699), .X(n9984) );
  nand_x1_sg U70679 ( .A(n39355), .B(n40702), .X(n10803) );
  nand_x1_sg U70680 ( .A(n39354), .B(n40708), .X(n11622) );
  nand_x1_sg U70681 ( .A(n39356), .B(n40714), .X(n12441) );
  nand_x1_sg U70682 ( .A(n39358), .B(n40717), .X(n13260) );
  nand_x1_sg U70683 ( .A(n39357), .B(n40723), .X(n14079) );
  nand_x1_sg U70684 ( .A(n39359), .B(n40727), .X(n14898) );
  nand_x1_sg U70685 ( .A(n39361), .B(n40732), .X(n15717) );
  nand_x1_sg U70686 ( .A(n39360), .B(n40738), .X(n16536) );
  nand_x1_sg U70687 ( .A(n39363), .B(n38909), .X(n18174) );
  nand_x1_sg U70688 ( .A(n39362), .B(n40744), .X(n18995) );
  nand_x1_sg U70689 ( .A(n39506), .B(n40689), .X(n8290) );
  nand_x1_sg U70690 ( .A(n39505), .B(n40693), .X(n9108) );
  nand_x1_sg U70691 ( .A(n39507), .B(n40699), .X(n9928) );
  nand_x1_sg U70692 ( .A(n39509), .B(n40703), .X(n10747) );
  nand_x1_sg U70693 ( .A(n39508), .B(n40709), .X(n11566) );
  nand_x1_sg U70694 ( .A(n39511), .B(n40714), .X(n12385) );
  nand_x1_sg U70695 ( .A(n39510), .B(n40718), .X(n13204) );
  nand_x1_sg U70696 ( .A(n39513), .B(n40724), .X(n14023) );
  nand_x1_sg U70697 ( .A(n39512), .B(n40728), .X(n14842) );
  nand_x1_sg U70698 ( .A(n39515), .B(n40733), .X(n15661) );
  nand_x1_sg U70699 ( .A(n39514), .B(n40739), .X(n16480) );
  nand_x1_sg U70700 ( .A(n39516), .B(n40619), .X(n18118) );
  nand_x1_sg U70701 ( .A(n39517), .B(n40743), .X(n18939) );
  nand_x1_sg U70702 ( .A(n40648), .B(n40618), .X(n17775) );
  nand_x1_sg U70703 ( .A(n8451), .B(n40689), .X(n8450) );
  nand_x1_sg U70704 ( .A(n9269), .B(n40693), .X(n9268) );
  nand_x1_sg U70705 ( .A(n10089), .B(n40697), .X(n10088) );
  nand_x1_sg U70706 ( .A(n10908), .B(n40701), .X(n10907) );
  nand_x1_sg U70707 ( .A(n11727), .B(n40706), .X(n11726) );
  nand_x1_sg U70708 ( .A(n12546), .B(n40712), .X(n12545) );
  nand_x1_sg U70709 ( .A(n13365), .B(n40719), .X(n13364) );
  nand_x1_sg U70710 ( .A(n14184), .B(n40721), .X(n14183) );
  nand_x1_sg U70711 ( .A(n15003), .B(n40728), .X(n15002) );
  nand_x1_sg U70712 ( .A(n15822), .B(n40733), .X(n15821) );
  nand_x1_sg U70713 ( .A(n16641), .B(n40736), .X(n16640) );
  nand_x1_sg U70714 ( .A(n18279), .B(n40619), .X(n18278) );
  nand_x1_sg U70715 ( .A(n19100), .B(n40742), .X(n19099) );
  nand_x1_sg U70716 ( .A(n7648), .B(n40689), .X(n7646) );
  nand_x1_sg U70717 ( .A(n40242), .B(n40306), .X(n7649) );
  nand_x1_sg U70718 ( .A(n42105), .B(n40560), .X(n7650) );
  nand_x1_sg U70719 ( .A(n8466), .B(n40694), .X(n8464) );
  nand_x1_sg U70720 ( .A(n40248), .B(n41844), .X(n8467) );
  nand_x1_sg U70721 ( .A(n40361), .B(n40556), .X(n8468) );
  nand_x1_sg U70722 ( .A(n9286), .B(n40696), .X(n9284) );
  nand_x1_sg U70723 ( .A(n40255), .B(n41853), .X(n9287) );
  nand_x1_sg U70724 ( .A(n40356), .B(n40552), .X(n9288) );
  nand_x1_sg U70725 ( .A(n10105), .B(n40704), .X(n10103) );
  nand_x1_sg U70726 ( .A(n40257), .B(n41855), .X(n10106) );
  nand_x1_sg U70727 ( .A(n40352), .B(n40548), .X(n10107) );
  nand_x1_sg U70728 ( .A(n10924), .B(n40706), .X(n10922) );
  nand_x1_sg U70729 ( .A(n40265), .B(n41851), .X(n10925) );
  nand_x1_sg U70730 ( .A(n40348), .B(n40544), .X(n10926) );
  nand_x1_sg U70731 ( .A(n11743), .B(n40711), .X(n11741) );
  nand_x1_sg U70732 ( .A(n40268), .B(n41857), .X(n11744) );
  nand_x1_sg U70733 ( .A(n40328), .B(n40540), .X(n11745) );
  nand_x1_sg U70734 ( .A(n12562), .B(n40719), .X(n12560) );
  nand_x1_sg U70735 ( .A(n40272), .B(n41859), .X(n12563) );
  nand_x1_sg U70736 ( .A(n40340), .B(n40536), .X(n12564) );
  nand_x1_sg U70737 ( .A(n13381), .B(n40721), .X(n13379) );
  nand_x1_sg U70738 ( .A(n40279), .B(n41849), .X(n13382) );
  nand_x1_sg U70739 ( .A(n40336), .B(n40532), .X(n13383) );
  nand_x1_sg U70740 ( .A(n14200), .B(n40726), .X(n14198) );
  nand_x1_sg U70741 ( .A(n40283), .B(n41837), .X(n14201) );
  nand_x1_sg U70742 ( .A(n40344), .B(n40528), .X(n14202) );
  nand_x1_sg U70743 ( .A(n15019), .B(n40734), .X(n15017) );
  nand_x1_sg U70744 ( .A(n40287), .B(n41846), .X(n15020) );
  nand_x1_sg U70745 ( .A(n42095), .B(n40524), .X(n15021) );
  nand_x1_sg U70746 ( .A(n15838), .B(n40736), .X(n15836) );
  nand_x1_sg U70747 ( .A(n40295), .B(n41839), .X(n15839) );
  nand_x1_sg U70748 ( .A(n40324), .B(n40520), .X(n15840) );
  nand_x1_sg U70749 ( .A(n17476), .B(n40618), .X(n17474) );
  nand_x1_sg U70750 ( .A(n40237), .B(n40364), .X(n17477) );
  nand_x1_sg U70751 ( .A(n40068), .B(n40516), .X(n17478) );
  nand_x1_sg U70752 ( .A(n18297), .B(n40741), .X(n18295) );
  nand_x1_sg U70753 ( .A(n40298), .B(n41841), .X(n18298) );
  nand_x1_sg U70754 ( .A(n40332), .B(n40512), .X(n18299) );
  nand_x1_sg U70755 ( .A(n39662), .B(n40570), .X(n17297) );
  nor_x1_sg U70756 ( .A(n6125), .B(n6126), .X(n6124) );
  nor_x1_sg U70757 ( .A(n6128), .B(n42258), .X(n6125) );
  nor_x1_sg U70758 ( .A(n6127), .B(n46435), .X(n6126) );
  inv_x1_sg U70759 ( .A(n6128), .X(n46435) );
  nor_x1_sg U70760 ( .A(n47074), .B(n42016), .X(n7013) );
  nor_x1_sg U70761 ( .A(n47360), .B(n42017), .X(n7831) );
  nor_x1_sg U70762 ( .A(n47645), .B(n42011), .X(n8649) );
  nor_x1_sg U70763 ( .A(n47930), .B(n42012), .X(n9469) );
  nor_x1_sg U70764 ( .A(n48215), .B(n42013), .X(n10288) );
  nor_x1_sg U70765 ( .A(n48500), .B(n42014), .X(n11107) );
  nor_x1_sg U70766 ( .A(n48785), .B(n42007), .X(n11926) );
  nor_x1_sg U70767 ( .A(n49072), .B(n42008), .X(n12745) );
  nor_x1_sg U70768 ( .A(n49358), .B(n42009), .X(n13564) );
  nor_x1_sg U70769 ( .A(n49644), .B(n42010), .X(n14383) );
  nor_x1_sg U70770 ( .A(n49930), .B(n42003), .X(n15202) );
  nor_x1_sg U70771 ( .A(n50216), .B(n42004), .X(n16021) );
  nor_x1_sg U70772 ( .A(n50790), .B(n42006), .X(n17659) );
  nor_x1_sg U70773 ( .A(n51077), .B(n42001), .X(n18480) );
  nand_x1_sg U70774 ( .A(n39364), .B(n40568), .X(n17353) );
  nand_x1_sg U70775 ( .A(n40581), .B(n40571), .X(n16954) );
  nand_x1_sg U70776 ( .A(n17458), .B(n40569), .X(n17457) );
  nand_x1_sg U70777 ( .A(n16654), .B(n40570), .X(n16652) );
  nand_x1_sg U70778 ( .A(n40069), .B(n40302), .X(n16656) );
  nand_x1_sg U70779 ( .A(n40563), .B(n40310), .X(n16657) );
  nand_x1_sg U70780 ( .A(n26822), .B(n26781), .X(n26820) );
  nor_x1_sg U70781 ( .A(n26781), .B(n26822), .X(n26821) );
  nand_x1_sg U70782 ( .A(n39350), .B(n6831), .X(n7528) );
  nand_x1_sg U70783 ( .A(n40575), .B(n40314), .X(n7129) );
  nand_x1_sg U70784 ( .A(n7633), .B(n6831), .X(n7632) );
  nand_x1_sg U70785 ( .A(n6830), .B(n40316), .X(n6828) );
  nand_x1_sg U70786 ( .A(n40162), .B(n40368), .X(n6832) );
  nand_x1_sg U70787 ( .A(n39957), .B(n40615), .X(n6833) );
  nor_x1_sg U70788 ( .A(n20977), .B(n42237), .X(n20976) );
  nor_x1_sg U70789 ( .A(n28535), .B(n42238), .X(n28534) );
  nor_x1_sg U70790 ( .A(n45868), .B(n6755), .X(n6754) );
  nor_x1_sg U70791 ( .A(n6756), .B(n6757), .X(n6755) );
  nand_x1_sg U70792 ( .A(n6757), .B(n6756), .X(n6758) );
  nand_x1_sg U70793 ( .A(n26771), .B(n26818), .X(n26817) );
  nor_x1_sg U70794 ( .A(n26818), .B(n26771), .X(n26819) );
  nand_x1_sg U70795 ( .A(n26765), .B(n26815), .X(n26814) );
  nor_x1_sg U70796 ( .A(n26815), .B(n26765), .X(n26816) );
  nand_x1_sg U70797 ( .A(n26777), .B(n26812), .X(n26811) );
  nor_x1_sg U70798 ( .A(n26812), .B(n26777), .X(n26813) );
  nand_x1_sg U70799 ( .A(n26790), .B(n28525), .X(n28524) );
  nor_x1_sg U70800 ( .A(n28525), .B(n26790), .X(n28526) );
  nand_x1_sg U70801 ( .A(n26770), .B(n26809), .X(n26808) );
  nor_x1_sg U70802 ( .A(n26809), .B(n26770), .X(n26810) );
  nand_x1_sg U70803 ( .A(n26784), .B(n28522), .X(n28521) );
  nor_x1_sg U70804 ( .A(n28522), .B(n26784), .X(n28523) );
  nand_x1_sg U70805 ( .A(n26785), .B(n28531), .X(n28530) );
  nor_x1_sg U70806 ( .A(n28531), .B(n26785), .X(n28532) );
  nand_x1_sg U70807 ( .A(n26766), .B(n26806), .X(n26805) );
  nor_x1_sg U70808 ( .A(n26806), .B(n26766), .X(n26807) );
  nand_x1_sg U70809 ( .A(n26827), .B(n26828), .X(n26826) );
  nor_x1_sg U70810 ( .A(n26828), .B(n26827), .X(n26829) );
  nand_x1_sg U70811 ( .A(n28519), .B(n28528), .X(n28527) );
  nor_x1_sg U70812 ( .A(n28528), .B(n28519), .X(n28529) );
  nand_x1_sg U70813 ( .A(n26780), .B(n26803), .X(n26802) );
  nor_x1_sg U70814 ( .A(n26803), .B(n26780), .X(n26804) );
  nand_x1_sg U70815 ( .A(n26953), .B(n26954), .X(n26952) );
  nor_x1_sg U70816 ( .A(n26954), .B(n26953), .X(n26955) );
  inv_x1_sg U70817 ( .A(n20359), .X(n45804) );
  inv_x1_sg U70818 ( .A(n19626), .X(n45808) );
  inv_x1_sg U70819 ( .A(n19216), .X(n45810) );
  inv_x1_sg U70820 ( .A(n20020), .X(n45806) );
  inv_x1_sg U70821 ( .A(n20660), .X(n45802) );
  inv_x1_sg U70822 ( .A(n21068), .X(n45800) );
  nor_x1_sg U70823 ( .A(n40021), .B(n25917), .X(\L1_0/n3476 ) );
  nand_x1_sg U70824 ( .A(n40570), .B(n41114), .X(n25917) );
  inv_x1_sg U70825 ( .A(n19903), .X(n46348) );
  inv_x1_sg U70826 ( .A(n19755), .X(n46510) );
  nand_x1_sg U70827 ( .A(n19311), .B(n38675), .X(n19352) );
  nand_x1_sg U70828 ( .A(n38756), .B(n38134), .X(n28814) );
  nand_x1_sg U70829 ( .A(n22721), .B(n22719), .X(n22726) );
  nand_x1_sg U70830 ( .A(n22998), .B(n22996), .X(n23003) );
  nand_x1_sg U70831 ( .A(n23278), .B(n23276), .X(n23283) );
  nand_x1_sg U70832 ( .A(n23557), .B(n23555), .X(n23562) );
  nand_x1_sg U70833 ( .A(n23836), .B(n23834), .X(n23841) );
  nand_x1_sg U70834 ( .A(n24115), .B(n24113), .X(n24120) );
  nand_x1_sg U70835 ( .A(n24394), .B(n24392), .X(n24399) );
  nand_x1_sg U70836 ( .A(n24672), .B(n24670), .X(n24677) );
  nand_x1_sg U70837 ( .A(n24951), .B(n24949), .X(n24956) );
  nand_x1_sg U70838 ( .A(n25230), .B(n25228), .X(n25235) );
  nand_x1_sg U70839 ( .A(n25509), .B(n25507), .X(n25514) );
  nand_x1_sg U70840 ( .A(n25786), .B(n25784), .X(n25791) );
  nand_x1_sg U70841 ( .A(n26132), .B(n26133), .X(n26131) );
  nand_x1_sg U70842 ( .A(n26346), .B(n26344), .X(n26351) );
  nand_x1_sg U70843 ( .A(n26624), .B(n26622), .X(n26629) );
  nand_x1_sg U70844 ( .A(n28142), .B(n38714), .X(n28247) );
  nand_x1_sg U70845 ( .A(n20508), .B(n38701), .X(n20651) );
  nand_x1_sg U70846 ( .A(n21277), .B(n38720), .X(n21421) );
  nand_x1_sg U70847 ( .A(n19851), .B(n38673), .X(n20011) );
  nand_x1_sg U70848 ( .A(n6671), .B(n38606), .X(n19207) );
  nand_x1_sg U70849 ( .A(n22718), .B(n47096), .X(n22717) );
  nand_x1_sg U70850 ( .A(n6003), .B(n19536), .X(n19535) );
  nand_x1_sg U70851 ( .A(n5969), .B(n19550), .X(n19549) );
  nand_x1_sg U70852 ( .A(n5965), .B(n19564), .X(n19563) );
  nand_x1_sg U70853 ( .A(n5974), .B(n5983), .X(n19152) );
  nor_x1_sg U70854 ( .A(n22810), .B(n22811), .X(n7094) );
  nor_x1_sg U70855 ( .A(n46868), .B(n22807), .X(n22811) );
  nor_x1_sg U70856 ( .A(n23087), .B(n23088), .X(n7912) );
  nor_x1_sg U70857 ( .A(n47161), .B(n23084), .X(n23088) );
  nor_x1_sg U70858 ( .A(n23367), .B(n23368), .X(n8730) );
  nor_x1_sg U70859 ( .A(n47446), .B(n23364), .X(n23368) );
  nor_x1_sg U70860 ( .A(n23646), .B(n23647), .X(n9550) );
  nor_x1_sg U70861 ( .A(n47731), .B(n23643), .X(n23647) );
  nor_x1_sg U70862 ( .A(n23925), .B(n23926), .X(n10369) );
  nor_x1_sg U70863 ( .A(n48016), .B(n23922), .X(n23926) );
  nor_x1_sg U70864 ( .A(n24204), .B(n24205), .X(n11188) );
  nor_x1_sg U70865 ( .A(n48301), .B(n24201), .X(n24205) );
  nor_x1_sg U70866 ( .A(n24483), .B(n24484), .X(n12007) );
  nor_x1_sg U70867 ( .A(n48586), .B(n24480), .X(n24484) );
  nor_x1_sg U70868 ( .A(n24761), .B(n24762), .X(n12826) );
  nor_x1_sg U70869 ( .A(n48872), .B(n24758), .X(n24762) );
  nor_x1_sg U70870 ( .A(n25040), .B(n25041), .X(n13645) );
  nor_x1_sg U70871 ( .A(n49159), .B(n25037), .X(n25041) );
  nor_x1_sg U70872 ( .A(n25319), .B(n25320), .X(n14464) );
  nor_x1_sg U70873 ( .A(n49445), .B(n25316), .X(n25320) );
  nor_x1_sg U70874 ( .A(n25598), .B(n25599), .X(n15283) );
  nor_x1_sg U70875 ( .A(n49730), .B(n25595), .X(n25599) );
  nor_x1_sg U70876 ( .A(n25875), .B(n25876), .X(n16102) );
  nor_x1_sg U70877 ( .A(n50017), .B(n25872), .X(n25876) );
  nor_x1_sg U70878 ( .A(n26435), .B(n26436), .X(n17740) );
  nor_x1_sg U70879 ( .A(n50591), .B(n26432), .X(n26436) );
  nor_x1_sg U70880 ( .A(n26713), .B(n26714), .X(n18561) );
  nor_x1_sg U70881 ( .A(n50878), .B(n26710), .X(n26714) );
  nand_x1_sg U70882 ( .A(n19325), .B(n38608), .X(n19323) );
  nor_x1_sg U70883 ( .A(n6038), .B(n19325), .X(n19324) );
  nand_x1_sg U70884 ( .A(n26049), .B(n26050), .X(n26048) );
  nand_x1_sg U70885 ( .A(n50435), .B(n26055), .X(n26152) );
  nand_x1_sg U70886 ( .A(n22771), .B(n22769), .X(n22775) );
  nand_x1_sg U70887 ( .A(n46903), .B(n22778), .X(n22777) );
  nand_x1_sg U70888 ( .A(n26061), .B(n26062), .X(n26060) );
  nand_x1_sg U70889 ( .A(n50395), .B(n26067), .X(n26154) );
  nand_x1_sg U70890 ( .A(n23062), .B(n23060), .X(n23066) );
  nand_x1_sg U70891 ( .A(n23342), .B(n23340), .X(n23346) );
  nand_x1_sg U70892 ( .A(n23621), .B(n23619), .X(n23625) );
  nand_x1_sg U70893 ( .A(n23900), .B(n23898), .X(n23904) );
  nand_x1_sg U70894 ( .A(n24179), .B(n24177), .X(n24183) );
  nand_x1_sg U70895 ( .A(n24458), .B(n24456), .X(n24462) );
  nand_x1_sg U70896 ( .A(n24736), .B(n24734), .X(n24740) );
  nand_x1_sg U70897 ( .A(n25015), .B(n25013), .X(n25019) );
  nand_x1_sg U70898 ( .A(n25294), .B(n25292), .X(n25298) );
  nand_x1_sg U70899 ( .A(n25573), .B(n25571), .X(n25577) );
  nand_x1_sg U70900 ( .A(n25850), .B(n25848), .X(n25854) );
  nand_x1_sg U70901 ( .A(n26085), .B(n26086), .X(n26083) );
  nand_x1_sg U70902 ( .A(n26410), .B(n26408), .X(n26414) );
  nand_x1_sg U70903 ( .A(n26688), .B(n26686), .X(n26692) );
  nand_x1_sg U70904 ( .A(n26073), .B(n26074), .X(n26072) );
  nand_x1_sg U70905 ( .A(n50356), .B(n26079), .X(n26156) );
  nand_x1_sg U70906 ( .A(n22785), .B(n22786), .X(n22784) );
  nand_x1_sg U70907 ( .A(n22778), .B(n22776), .X(n22782) );
  nand_x1_sg U70908 ( .A(n46924), .B(n22771), .X(n22770) );
  nand_x1_sg U70909 ( .A(n22764), .B(n22762), .X(n22768) );
  nand_x1_sg U70910 ( .A(n22757), .B(n22755), .X(n22761) );
  nand_x1_sg U70911 ( .A(n46942), .B(n22764), .X(n22763) );
  nand_x1_sg U70912 ( .A(n46965), .B(n22757), .X(n22756) );
  nand_x1_sg U70913 ( .A(n22750), .B(n22748), .X(n22754) );
  nand_x1_sg U70914 ( .A(n22743), .B(n22741), .X(n22747) );
  nand_x1_sg U70915 ( .A(n46984), .B(n22750), .X(n22749) );
  nand_x1_sg U70916 ( .A(n47007), .B(n22743), .X(n22742) );
  nand_x1_sg U70917 ( .A(n22736), .B(n22734), .X(n22740) );
  nand_x1_sg U70918 ( .A(n23062), .B(n23063), .X(n23061) );
  nand_x1_sg U70919 ( .A(n23055), .B(n23053), .X(n23059) );
  nand_x1_sg U70920 ( .A(n23048), .B(n23046), .X(n23052) );
  nand_x1_sg U70921 ( .A(n47196), .B(n23055), .X(n23054) );
  nand_x1_sg U70922 ( .A(n47216), .B(n23048), .X(n23047) );
  nand_x1_sg U70923 ( .A(n23041), .B(n23039), .X(n23045) );
  nand_x1_sg U70924 ( .A(n23034), .B(n23032), .X(n23038) );
  nand_x1_sg U70925 ( .A(n47233), .B(n23041), .X(n23040) );
  nand_x1_sg U70926 ( .A(n47255), .B(n23034), .X(n23033) );
  nand_x1_sg U70927 ( .A(n23027), .B(n23025), .X(n23031) );
  nand_x1_sg U70928 ( .A(n23020), .B(n23018), .X(n23024) );
  nand_x1_sg U70929 ( .A(n47273), .B(n23027), .X(n23026) );
  nand_x1_sg U70930 ( .A(n47295), .B(n23020), .X(n23019) );
  nand_x1_sg U70931 ( .A(n23013), .B(n23011), .X(n23017) );
  nand_x1_sg U70932 ( .A(n23342), .B(n23343), .X(n23341) );
  nand_x1_sg U70933 ( .A(n23335), .B(n23333), .X(n23339) );
  nand_x1_sg U70934 ( .A(n23328), .B(n23326), .X(n23332) );
  nand_x1_sg U70935 ( .A(n47481), .B(n23335), .X(n23334) );
  nand_x1_sg U70936 ( .A(n47501), .B(n23328), .X(n23327) );
  nand_x1_sg U70937 ( .A(n23321), .B(n23319), .X(n23325) );
  nand_x1_sg U70938 ( .A(n23314), .B(n23312), .X(n23318) );
  nand_x1_sg U70939 ( .A(n47518), .B(n23321), .X(n23320) );
  nand_x1_sg U70940 ( .A(n47540), .B(n23314), .X(n23313) );
  nand_x1_sg U70941 ( .A(n23307), .B(n23305), .X(n23311) );
  nand_x1_sg U70942 ( .A(n23300), .B(n23298), .X(n23304) );
  nand_x1_sg U70943 ( .A(n47558), .B(n23307), .X(n23306) );
  nand_x1_sg U70944 ( .A(n47580), .B(n23300), .X(n23299) );
  nand_x1_sg U70945 ( .A(n23293), .B(n23291), .X(n23297) );
  nand_x1_sg U70946 ( .A(n23621), .B(n23622), .X(n23620) );
  nand_x1_sg U70947 ( .A(n23614), .B(n23612), .X(n23618) );
  nand_x1_sg U70948 ( .A(n23607), .B(n23605), .X(n23611) );
  nand_x1_sg U70949 ( .A(n47766), .B(n23614), .X(n23613) );
  nand_x1_sg U70950 ( .A(n47786), .B(n23607), .X(n23606) );
  nand_x1_sg U70951 ( .A(n23600), .B(n23598), .X(n23604) );
  nand_x1_sg U70952 ( .A(n23593), .B(n23591), .X(n23597) );
  nand_x1_sg U70953 ( .A(n47803), .B(n23600), .X(n23599) );
  nand_x1_sg U70954 ( .A(n47825), .B(n23593), .X(n23592) );
  nand_x1_sg U70955 ( .A(n23586), .B(n23584), .X(n23590) );
  nand_x1_sg U70956 ( .A(n23579), .B(n23577), .X(n23583) );
  nand_x1_sg U70957 ( .A(n47843), .B(n23586), .X(n23585) );
  nand_x1_sg U70958 ( .A(n47865), .B(n23579), .X(n23578) );
  nand_x1_sg U70959 ( .A(n23572), .B(n23570), .X(n23576) );
  nand_x1_sg U70960 ( .A(n23900), .B(n23901), .X(n23899) );
  nand_x1_sg U70961 ( .A(n23893), .B(n23891), .X(n23897) );
  nand_x1_sg U70962 ( .A(n23886), .B(n23884), .X(n23890) );
  nand_x1_sg U70963 ( .A(n48051), .B(n23893), .X(n23892) );
  nand_x1_sg U70964 ( .A(n48071), .B(n23886), .X(n23885) );
  nand_x1_sg U70965 ( .A(n23879), .B(n23877), .X(n23883) );
  nand_x1_sg U70966 ( .A(n23872), .B(n23870), .X(n23876) );
  nand_x1_sg U70967 ( .A(n48088), .B(n23879), .X(n23878) );
  nand_x1_sg U70968 ( .A(n48110), .B(n23872), .X(n23871) );
  nand_x1_sg U70969 ( .A(n23865), .B(n23863), .X(n23869) );
  nand_x1_sg U70970 ( .A(n23858), .B(n23856), .X(n23862) );
  nand_x1_sg U70971 ( .A(n48128), .B(n23865), .X(n23864) );
  nand_x1_sg U70972 ( .A(n48150), .B(n23858), .X(n23857) );
  nand_x1_sg U70973 ( .A(n23851), .B(n23849), .X(n23855) );
  nand_x1_sg U70974 ( .A(n24179), .B(n24180), .X(n24178) );
  nand_x1_sg U70975 ( .A(n24172), .B(n24170), .X(n24176) );
  nand_x1_sg U70976 ( .A(n24165), .B(n24163), .X(n24169) );
  nand_x1_sg U70977 ( .A(n48336), .B(n24172), .X(n24171) );
  nand_x1_sg U70978 ( .A(n48356), .B(n24165), .X(n24164) );
  nand_x1_sg U70979 ( .A(n24158), .B(n24156), .X(n24162) );
  nand_x1_sg U70980 ( .A(n24151), .B(n24149), .X(n24155) );
  nand_x1_sg U70981 ( .A(n48373), .B(n24158), .X(n24157) );
  nand_x1_sg U70982 ( .A(n48395), .B(n24151), .X(n24150) );
  nand_x1_sg U70983 ( .A(n24144), .B(n24142), .X(n24148) );
  nand_x1_sg U70984 ( .A(n24137), .B(n24135), .X(n24141) );
  nand_x1_sg U70985 ( .A(n48413), .B(n24144), .X(n24143) );
  nand_x1_sg U70986 ( .A(n48435), .B(n24137), .X(n24136) );
  nand_x1_sg U70987 ( .A(n24130), .B(n24128), .X(n24134) );
  nand_x1_sg U70988 ( .A(n24458), .B(n24459), .X(n24457) );
  nand_x1_sg U70989 ( .A(n24451), .B(n24449), .X(n24455) );
  nand_x1_sg U70990 ( .A(n24444), .B(n24442), .X(n24448) );
  nand_x1_sg U70991 ( .A(n48621), .B(n24451), .X(n24450) );
  nand_x1_sg U70992 ( .A(n48641), .B(n24444), .X(n24443) );
  nand_x1_sg U70993 ( .A(n24437), .B(n24435), .X(n24441) );
  nand_x1_sg U70994 ( .A(n24430), .B(n24428), .X(n24434) );
  nand_x1_sg U70995 ( .A(n48658), .B(n24437), .X(n24436) );
  nand_x1_sg U70996 ( .A(n48680), .B(n24430), .X(n24429) );
  nand_x1_sg U70997 ( .A(n24423), .B(n24421), .X(n24427) );
  nand_x1_sg U70998 ( .A(n24416), .B(n24414), .X(n24420) );
  nand_x1_sg U70999 ( .A(n48698), .B(n24423), .X(n24422) );
  nand_x1_sg U71000 ( .A(n48720), .B(n24416), .X(n24415) );
  nand_x1_sg U71001 ( .A(n24409), .B(n24407), .X(n24413) );
  nand_x1_sg U71002 ( .A(n24736), .B(n24737), .X(n24735) );
  nand_x1_sg U71003 ( .A(n24729), .B(n24727), .X(n24733) );
  nand_x1_sg U71004 ( .A(n24722), .B(n24720), .X(n24726) );
  nand_x1_sg U71005 ( .A(n48907), .B(n24729), .X(n24728) );
  nand_x1_sg U71006 ( .A(n48927), .B(n24722), .X(n24721) );
  nand_x1_sg U71007 ( .A(n24715), .B(n24713), .X(n24719) );
  nand_x1_sg U71008 ( .A(n24708), .B(n24706), .X(n24712) );
  nand_x1_sg U71009 ( .A(n48944), .B(n24715), .X(n24714) );
  nand_x1_sg U71010 ( .A(n48966), .B(n24708), .X(n24707) );
  nand_x1_sg U71011 ( .A(n24701), .B(n24699), .X(n24705) );
  nand_x1_sg U71012 ( .A(n24694), .B(n24692), .X(n24698) );
  nand_x1_sg U71013 ( .A(n48984), .B(n24701), .X(n24700) );
  nand_x1_sg U71014 ( .A(n49006), .B(n24694), .X(n24693) );
  nand_x1_sg U71015 ( .A(n24687), .B(n24685), .X(n24691) );
  nand_x1_sg U71016 ( .A(n25015), .B(n25016), .X(n25014) );
  nand_x1_sg U71017 ( .A(n25008), .B(n25006), .X(n25012) );
  nand_x1_sg U71018 ( .A(n25001), .B(n24999), .X(n25005) );
  nand_x1_sg U71019 ( .A(n49194), .B(n25008), .X(n25007) );
  nand_x1_sg U71020 ( .A(n49214), .B(n25001), .X(n25000) );
  nand_x1_sg U71021 ( .A(n24994), .B(n24992), .X(n24998) );
  nand_x1_sg U71022 ( .A(n24987), .B(n24985), .X(n24991) );
  nand_x1_sg U71023 ( .A(n49231), .B(n24994), .X(n24993) );
  nand_x1_sg U71024 ( .A(n49253), .B(n24987), .X(n24986) );
  nand_x1_sg U71025 ( .A(n24980), .B(n24978), .X(n24984) );
  nand_x1_sg U71026 ( .A(n24973), .B(n24971), .X(n24977) );
  nand_x1_sg U71027 ( .A(n49271), .B(n24980), .X(n24979) );
  nand_x1_sg U71028 ( .A(n49293), .B(n24973), .X(n24972) );
  nand_x1_sg U71029 ( .A(n24966), .B(n24964), .X(n24970) );
  nand_x1_sg U71030 ( .A(n25294), .B(n25295), .X(n25293) );
  nand_x1_sg U71031 ( .A(n25287), .B(n25285), .X(n25291) );
  nand_x1_sg U71032 ( .A(n25280), .B(n25278), .X(n25284) );
  nand_x1_sg U71033 ( .A(n49480), .B(n25287), .X(n25286) );
  nand_x1_sg U71034 ( .A(n49500), .B(n25280), .X(n25279) );
  nand_x1_sg U71035 ( .A(n25273), .B(n25271), .X(n25277) );
  nand_x1_sg U71036 ( .A(n25266), .B(n25264), .X(n25270) );
  nand_x1_sg U71037 ( .A(n49517), .B(n25273), .X(n25272) );
  nand_x1_sg U71038 ( .A(n49539), .B(n25266), .X(n25265) );
  nand_x1_sg U71039 ( .A(n25259), .B(n25257), .X(n25263) );
  nand_x1_sg U71040 ( .A(n25252), .B(n25250), .X(n25256) );
  nand_x1_sg U71041 ( .A(n49557), .B(n25259), .X(n25258) );
  nand_x1_sg U71042 ( .A(n49579), .B(n25252), .X(n25251) );
  nand_x1_sg U71043 ( .A(n25245), .B(n25243), .X(n25249) );
  nand_x1_sg U71044 ( .A(n25573), .B(n25574), .X(n25572) );
  nand_x1_sg U71045 ( .A(n25566), .B(n25564), .X(n25570) );
  nand_x1_sg U71046 ( .A(n25559), .B(n25557), .X(n25563) );
  nand_x1_sg U71047 ( .A(n49766), .B(n25566), .X(n25565) );
  nand_x1_sg U71048 ( .A(n49786), .B(n25559), .X(n25558) );
  nand_x1_sg U71049 ( .A(n25552), .B(n25550), .X(n25556) );
  nand_x1_sg U71050 ( .A(n25545), .B(n25543), .X(n25549) );
  nand_x1_sg U71051 ( .A(n49803), .B(n25552), .X(n25551) );
  nand_x1_sg U71052 ( .A(n49825), .B(n25545), .X(n25544) );
  nand_x1_sg U71053 ( .A(n25538), .B(n25536), .X(n25542) );
  nand_x1_sg U71054 ( .A(n25531), .B(n25529), .X(n25535) );
  nand_x1_sg U71055 ( .A(n49843), .B(n25538), .X(n25537) );
  nand_x1_sg U71056 ( .A(n49865), .B(n25531), .X(n25530) );
  nand_x1_sg U71057 ( .A(n25524), .B(n25522), .X(n25528) );
  nand_x1_sg U71058 ( .A(n25850), .B(n25851), .X(n25849) );
  nand_x1_sg U71059 ( .A(n25843), .B(n25841), .X(n25847) );
  nand_x1_sg U71060 ( .A(n25836), .B(n25834), .X(n25840) );
  nand_x1_sg U71061 ( .A(n50052), .B(n25843), .X(n25842) );
  nand_x1_sg U71062 ( .A(n50072), .B(n25836), .X(n25835) );
  nand_x1_sg U71063 ( .A(n25829), .B(n25827), .X(n25833) );
  nand_x1_sg U71064 ( .A(n25822), .B(n25820), .X(n25826) );
  nand_x1_sg U71065 ( .A(n50089), .B(n25829), .X(n25828) );
  nand_x1_sg U71066 ( .A(n50111), .B(n25822), .X(n25821) );
  nand_x1_sg U71067 ( .A(n25815), .B(n25813), .X(n25819) );
  nand_x1_sg U71068 ( .A(n25808), .B(n25806), .X(n25812) );
  nand_x1_sg U71069 ( .A(n50129), .B(n25815), .X(n25814) );
  nand_x1_sg U71070 ( .A(n50151), .B(n25808), .X(n25807) );
  nand_x1_sg U71071 ( .A(n25801), .B(n25799), .X(n25805) );
  nand_x1_sg U71072 ( .A(n26085), .B(n26084), .X(n26157) );
  nand_x1_sg U71073 ( .A(n26079), .B(n26080), .X(n26077) );
  nand_x1_sg U71074 ( .A(n50373), .B(n26073), .X(n26155) );
  nand_x1_sg U71075 ( .A(n26067), .B(n26068), .X(n26065) );
  nand_x1_sg U71076 ( .A(n50413), .B(n26061), .X(n26153) );
  nand_x1_sg U71077 ( .A(n26055), .B(n26056), .X(n26053) );
  nand_x1_sg U71078 ( .A(n50453), .B(n26049), .X(n26151) );
  nand_x1_sg U71079 ( .A(n26043), .B(n26044), .X(n26041) );
  nand_x1_sg U71080 ( .A(n26410), .B(n26411), .X(n26409) );
  nand_x1_sg U71081 ( .A(n26403), .B(n26401), .X(n26407) );
  nand_x1_sg U71082 ( .A(n26396), .B(n26394), .X(n26400) );
  nand_x1_sg U71083 ( .A(n50626), .B(n26403), .X(n26402) );
  nand_x1_sg U71084 ( .A(n50646), .B(n26396), .X(n26395) );
  nand_x1_sg U71085 ( .A(n26389), .B(n26387), .X(n26393) );
  nand_x1_sg U71086 ( .A(n26382), .B(n26380), .X(n26386) );
  nand_x1_sg U71087 ( .A(n50663), .B(n26389), .X(n26388) );
  nand_x1_sg U71088 ( .A(n50685), .B(n26382), .X(n26381) );
  nand_x1_sg U71089 ( .A(n26375), .B(n26373), .X(n26379) );
  nand_x1_sg U71090 ( .A(n26368), .B(n26366), .X(n26372) );
  nand_x1_sg U71091 ( .A(n50703), .B(n26375), .X(n26374) );
  nand_x1_sg U71092 ( .A(n50725), .B(n26368), .X(n26367) );
  nand_x1_sg U71093 ( .A(n26361), .B(n26359), .X(n26365) );
  nand_x1_sg U71094 ( .A(n26688), .B(n26689), .X(n26687) );
  nand_x1_sg U71095 ( .A(n26681), .B(n26679), .X(n26685) );
  nand_x1_sg U71096 ( .A(n26674), .B(n26672), .X(n26678) );
  nand_x1_sg U71097 ( .A(n50913), .B(n26681), .X(n26680) );
  nand_x1_sg U71098 ( .A(n50933), .B(n26674), .X(n26673) );
  nand_x1_sg U71099 ( .A(n26667), .B(n26665), .X(n26671) );
  nand_x1_sg U71100 ( .A(n26660), .B(n26658), .X(n26664) );
  nand_x1_sg U71101 ( .A(n50950), .B(n26667), .X(n26666) );
  nand_x1_sg U71102 ( .A(n50972), .B(n26660), .X(n26659) );
  nand_x1_sg U71103 ( .A(n26653), .B(n26651), .X(n26657) );
  nand_x1_sg U71104 ( .A(n26646), .B(n26644), .X(n26650) );
  nand_x1_sg U71105 ( .A(n50990), .B(n26653), .X(n26652) );
  nand_x1_sg U71106 ( .A(n51012), .B(n26646), .X(n26645) );
  nand_x1_sg U71107 ( .A(n26639), .B(n26637), .X(n26643) );
  nand_x1_sg U71108 ( .A(n22785), .B(n22783), .X(n22789) );
  nand_x1_sg U71109 ( .A(n22729), .B(n22727), .X(n22733) );
  nand_x1_sg U71110 ( .A(n47026), .B(n22736), .X(n22735) );
  nand_x1_sg U71111 ( .A(n23006), .B(n23004), .X(n23010) );
  nand_x1_sg U71112 ( .A(n47313), .B(n23013), .X(n23012) );
  nand_x1_sg U71113 ( .A(n23286), .B(n23284), .X(n23290) );
  nand_x1_sg U71114 ( .A(n47598), .B(n23293), .X(n23292) );
  nand_x1_sg U71115 ( .A(n23565), .B(n23563), .X(n23569) );
  nand_x1_sg U71116 ( .A(n47883), .B(n23572), .X(n23571) );
  nand_x1_sg U71117 ( .A(n23844), .B(n23842), .X(n23848) );
  nand_x1_sg U71118 ( .A(n48168), .B(n23851), .X(n23850) );
  nand_x1_sg U71119 ( .A(n24123), .B(n24121), .X(n24127) );
  nand_x1_sg U71120 ( .A(n48453), .B(n24130), .X(n24129) );
  nand_x1_sg U71121 ( .A(n24402), .B(n24400), .X(n24406) );
  nand_x1_sg U71122 ( .A(n48738), .B(n24409), .X(n24408) );
  nand_x1_sg U71123 ( .A(n24680), .B(n24678), .X(n24684) );
  nand_x1_sg U71124 ( .A(n49024), .B(n24687), .X(n24686) );
  nand_x1_sg U71125 ( .A(n24959), .B(n24957), .X(n24963) );
  nand_x1_sg U71126 ( .A(n49311), .B(n24966), .X(n24965) );
  nand_x1_sg U71127 ( .A(n25238), .B(n25236), .X(n25242) );
  nand_x1_sg U71128 ( .A(n49597), .B(n25245), .X(n25244) );
  nand_x1_sg U71129 ( .A(n25517), .B(n25515), .X(n25521) );
  nand_x1_sg U71130 ( .A(n49883), .B(n25524), .X(n25523) );
  nand_x1_sg U71131 ( .A(n25794), .B(n25792), .X(n25798) );
  nand_x1_sg U71132 ( .A(n50169), .B(n25801), .X(n25800) );
  nand_x1_sg U71133 ( .A(n26138), .B(n26139), .X(n26137) );
  nand_x1_sg U71134 ( .A(n50482), .B(n26043), .X(n26150) );
  nand_x1_sg U71135 ( .A(n26354), .B(n26352), .X(n26358) );
  nand_x1_sg U71136 ( .A(n50743), .B(n26361), .X(n26360) );
  nand_x1_sg U71137 ( .A(n26632), .B(n26630), .X(n26636) );
  nand_x1_sg U71138 ( .A(n51030), .B(n26639), .X(n26638) );
  nand_x1_sg U71139 ( .A(n38634), .B(n21005), .X(n21004) );
  nand_x1_sg U71140 ( .A(n38695), .B(n19337), .X(n19569) );
  nand_x1_sg U71141 ( .A(n38718), .B(n19145), .X(n19144) );
  nand_x1_sg U71142 ( .A(n20567), .B(n38756), .X(n22592) );
  nand_x1_sg U71143 ( .A(n22594), .B(n41093), .X(n22593) );
  nand_x1_sg U71144 ( .A(n21258), .B(n38140), .X(n21262) );
  nand_x1_sg U71145 ( .A(n42159), .B(n38133), .X(n27974) );
  inv_x1_sg U71146 ( .A(n20116), .X(n46397) );
  inv_x1_sg U71147 ( .A(n19328), .X(n46526) );
  inv_x1_sg U71148 ( .A(n19322), .X(n46481) );
  inv_x1_sg U71149 ( .A(n19722), .X(n46484) );
  inv_x1_sg U71150 ( .A(n23077), .X(n47170) );
  inv_x1_sg U71151 ( .A(n23357), .X(n47455) );
  inv_x1_sg U71152 ( .A(n23636), .X(n47740) );
  inv_x1_sg U71153 ( .A(n23915), .X(n48025) );
  inv_x1_sg U71154 ( .A(n24194), .X(n48310) );
  inv_x1_sg U71155 ( .A(n24473), .X(n48595) );
  inv_x1_sg U71156 ( .A(n24751), .X(n48881) );
  inv_x1_sg U71157 ( .A(n25030), .X(n49168) );
  inv_x1_sg U71158 ( .A(n25309), .X(n49454) );
  inv_x1_sg U71159 ( .A(n25588), .X(n49739) );
  inv_x1_sg U71160 ( .A(n25865), .X(n50026) );
  inv_x1_sg U71161 ( .A(n26425), .X(n50600) );
  inv_x1_sg U71162 ( .A(n26703), .X(n50887) );
  inv_x1_sg U71163 ( .A(n22800), .X(n46877) );
  nand_x1_sg U71164 ( .A(n19328), .B(n38608), .X(n19342) );
  nand_x1_sg U71165 ( .A(n19322), .B(n38716), .X(n19345) );
  nand_x1_sg U71166 ( .A(n44964), .B(n38196), .X(n28985) );
  nand_x1_sg U71167 ( .A(n45798), .B(n38197), .X(n21434) );
  nand_x1_sg U71168 ( .A(n45803), .B(n38136), .X(n20493) );
  nand_x1_sg U71169 ( .A(n45807), .B(n38138), .X(n19836) );
  nand_x1_sg U71170 ( .A(n45809), .B(n38139), .X(n19397) );
  nand_x1_sg U71171 ( .A(n45805), .B(n38137), .X(n20203) );
  nand_x1_sg U71172 ( .A(n45801), .B(n38135), .X(n20846) );
  nor_x1_sg U71173 ( .A(n41057), .B(n7010), .X(n7008) );
  nor_x1_sg U71174 ( .A(n7011), .B(n47120), .X(n7010) );
  nor_x1_sg U71175 ( .A(n7012), .B(n7013), .X(n7011) );
  nand_x1_sg U71176 ( .A(n23070), .B(n23067), .X(n23072) );
  nand_x1_sg U71177 ( .A(n23350), .B(n23347), .X(n23352) );
  nand_x1_sg U71178 ( .A(n23629), .B(n23626), .X(n23631) );
  nand_x1_sg U71179 ( .A(n23908), .B(n23905), .X(n23910) );
  nand_x1_sg U71180 ( .A(n24187), .B(n24184), .X(n24189) );
  nand_x1_sg U71181 ( .A(n24466), .B(n24463), .X(n24468) );
  nand_x1_sg U71182 ( .A(n24744), .B(n24741), .X(n24746) );
  nand_x1_sg U71183 ( .A(n25023), .B(n25020), .X(n25025) );
  nand_x1_sg U71184 ( .A(n25302), .B(n25299), .X(n25304) );
  nand_x1_sg U71185 ( .A(n25581), .B(n25578), .X(n25583) );
  nand_x1_sg U71186 ( .A(n25858), .B(n25855), .X(n25860) );
  nand_x1_sg U71187 ( .A(n26418), .B(n26415), .X(n26420) );
  nand_x1_sg U71188 ( .A(n26696), .B(n26693), .X(n26698) );
  nand_x1_sg U71189 ( .A(n22793), .B(n22790), .X(n22796) );
  nand_x1_sg U71190 ( .A(n26091), .B(n26092), .X(n26090) );
  nor_x1_sg U71191 ( .A(n41929), .B(n7827), .X(n7825) );
  nor_x1_sg U71192 ( .A(n7828), .B(n7829), .X(n7827) );
  nor_x1_sg U71193 ( .A(n7830), .B(n7831), .X(n7828) );
  nor_x1_sg U71194 ( .A(n39969), .B(n8645), .X(n8643) );
  nor_x1_sg U71195 ( .A(n8646), .B(n8647), .X(n8645) );
  nor_x1_sg U71196 ( .A(n8648), .B(n8649), .X(n8646) );
  nor_x1_sg U71197 ( .A(n39971), .B(n9465), .X(n9463) );
  nor_x1_sg U71198 ( .A(n9466), .B(n9467), .X(n9465) );
  nor_x1_sg U71199 ( .A(n9468), .B(n9469), .X(n9466) );
  nor_x1_sg U71200 ( .A(n41926), .B(n10284), .X(n10282) );
  nor_x1_sg U71201 ( .A(n10285), .B(n10286), .X(n10284) );
  nor_x1_sg U71202 ( .A(n10287), .B(n10288), .X(n10285) );
  nor_x1_sg U71203 ( .A(n39981), .B(n11103), .X(n11101) );
  nor_x1_sg U71204 ( .A(n11104), .B(n11105), .X(n11103) );
  nor_x1_sg U71205 ( .A(n11106), .B(n11107), .X(n11104) );
  nor_x1_sg U71206 ( .A(n41943), .B(n11922), .X(n11920) );
  nor_x1_sg U71207 ( .A(n11923), .B(n11924), .X(n11922) );
  nor_x1_sg U71208 ( .A(n11925), .B(n11926), .X(n11923) );
  nor_x1_sg U71209 ( .A(n41923), .B(n12741), .X(n12739) );
  nor_x1_sg U71210 ( .A(n12742), .B(n12743), .X(n12741) );
  nor_x1_sg U71211 ( .A(n12744), .B(n12745), .X(n12742) );
  nor_x1_sg U71212 ( .A(n40720), .B(n13560), .X(n13558) );
  nor_x1_sg U71213 ( .A(n13561), .B(n13562), .X(n13560) );
  nor_x1_sg U71214 ( .A(n13563), .B(n13564), .X(n13561) );
  nor_x1_sg U71215 ( .A(n41921), .B(n14379), .X(n14377) );
  nor_x1_sg U71216 ( .A(n14380), .B(n14381), .X(n14379) );
  nor_x1_sg U71217 ( .A(n14382), .B(n14383), .X(n14380) );
  nor_x1_sg U71218 ( .A(n41920), .B(n15198), .X(n15196) );
  nor_x1_sg U71219 ( .A(n15199), .B(n15200), .X(n15198) );
  nor_x1_sg U71220 ( .A(n15201), .B(n15202), .X(n15199) );
  nor_x1_sg U71221 ( .A(n40005), .B(n16017), .X(n16015) );
  nor_x1_sg U71222 ( .A(n16018), .B(n16019), .X(n16017) );
  nor_x1_sg U71223 ( .A(n16020), .B(n16021), .X(n16018) );
  nor_x1_sg U71224 ( .A(n40999), .B(n17655), .X(n17653) );
  nor_x1_sg U71225 ( .A(n17656), .B(n17657), .X(n17655) );
  nor_x1_sg U71226 ( .A(n17658), .B(n17659), .X(n17656) );
  nor_x1_sg U71227 ( .A(n40007), .B(n18476), .X(n18474) );
  nor_x1_sg U71228 ( .A(n18477), .B(n18478), .X(n18476) );
  nor_x1_sg U71229 ( .A(n18479), .B(n18480), .X(n18477) );
  nand_x1_sg U71230 ( .A(n50548), .B(n16834), .X(n16833) );
  nor_x1_sg U71231 ( .A(n40994), .B(n16835), .X(n16832) );
  nor_x1_sg U71232 ( .A(n16836), .B(n50548), .X(n16835) );
  nand_x1_sg U71233 ( .A(n44964), .B(n41395), .X(n22576) );
  nand_x1_sg U71234 ( .A(n39266), .B(n22578), .X(n22577) );
  nand_x1_sg U71235 ( .A(n21173), .B(n38634), .X(n21171) );
  nor_x1_sg U71236 ( .A(n5998), .B(n21173), .X(n21172) );
  nand_x1_sg U71237 ( .A(n46430), .B(n46395), .X(n19706) );
  nand_x1_sg U71238 ( .A(n19707), .B(n6162), .X(n19705) );
  nand_x1_sg U71239 ( .A(n19761), .B(n38626), .X(n19760) );
  nand_x1_sg U71240 ( .A(n20276), .B(n20280), .X(n20320) );
  nand_x1_sg U71241 ( .A(n46309), .B(n46336), .X(n20322) );
  nand_x1_sg U71242 ( .A(n20947), .B(n20951), .X(n21017) );
  nand_x1_sg U71243 ( .A(n46493), .B(n46506), .X(n21019) );
  nand_x1_sg U71244 ( .A(n19296), .B(n19299), .X(n19356) );
  nand_x1_sg U71245 ( .A(n46298), .B(n42224), .X(n19358) );
  inv_x1_sg U71246 ( .A(n6802), .X(n45811) );
  nand_x1_sg U71247 ( .A(n21092), .B(n38642), .X(n21245) );
  nand_x1_sg U71248 ( .A(n20383), .B(n38722), .X(n20477) );
  nand_x1_sg U71249 ( .A(n19650), .B(n38689), .X(n19820) );
  nand_x1_sg U71250 ( .A(n19773), .B(n38636), .X(n19772) );
  nand_x1_sg U71251 ( .A(n19956), .B(n38640), .X(n19955) );
  nand_x1_sg U71252 ( .A(n20148), .B(n38699), .X(n20147) );
  nand_x1_sg U71253 ( .A(n19795), .B(n38583), .X(n19794) );
  nor_x1_sg U71254 ( .A(n6255), .B(n19698), .X(n19796) );
  inv_x1_sg U71255 ( .A(n19550), .X(n46562) );
  inv_x1_sg U71256 ( .A(n6131), .X(n46434) );
  inv_x1_sg U71257 ( .A(n20786), .X(n46580) );
  inv_x1_sg U71258 ( .A(n19536), .X(n46558) );
  inv_x1_sg U71259 ( .A(n6223), .X(n46341) );
  inv_x1_sg U71260 ( .A(n20867), .X(n45955) );
  inv_x1_sg U71261 ( .A(n20224), .X(n45946) );
  inv_x1_sg U71262 ( .A(n19418), .X(n45937) );
  inv_x1_sg U71263 ( .A(n20136), .X(n46489) );
  inv_x1_sg U71264 ( .A(n19909), .X(n46396) );
  inv_x1_sg U71265 ( .A(n19564), .X(n46576) );
  inv_x1_sg U71266 ( .A(n26850), .X(n45710) );
  inv_x1_sg U71267 ( .A(n20998), .X(n46547) );
  inv_x1_sg U71268 ( .A(n5983), .X(n46572) );
  inv_x1_sg U71269 ( .A(n20680), .X(n45906) );
  inv_x1_sg U71270 ( .A(n20040), .X(n45896) );
  inv_x1_sg U71271 ( .A(n19236), .X(n45886) );
  inv_x1_sg U71272 ( .A(n19500), .X(n46483) );
  inv_x1_sg U71273 ( .A(n22816), .X(n46850) );
  nand_x1_sg U71274 ( .A(n7829), .B(n22992), .X(n7826) );
  nand_x1_sg U71275 ( .A(n8647), .B(n23272), .X(n8644) );
  nand_x1_sg U71276 ( .A(n9467), .B(n23551), .X(n9464) );
  nand_x1_sg U71277 ( .A(n10286), .B(n23830), .X(n10283) );
  nand_x1_sg U71278 ( .A(n11105), .B(n24109), .X(n11102) );
  nand_x1_sg U71279 ( .A(n11924), .B(n24388), .X(n11921) );
  nand_x1_sg U71280 ( .A(n12743), .B(n24666), .X(n12740) );
  nand_x1_sg U71281 ( .A(n13562), .B(n24945), .X(n13559) );
  nand_x1_sg U71282 ( .A(n14381), .B(n25224), .X(n14378) );
  nand_x1_sg U71283 ( .A(n15200), .B(n25503), .X(n15197) );
  nand_x1_sg U71284 ( .A(n16019), .B(n25780), .X(n16016) );
  nand_x1_sg U71285 ( .A(n17657), .B(n26340), .X(n17654) );
  nand_x1_sg U71286 ( .A(n18478), .B(n26618), .X(n18475) );
  inv_x1_sg U71287 ( .A(n21258), .X(n45799) );
  nand_x1_sg U71288 ( .A(n21146), .B(n38563), .X(n21144) );
  nor_x1_sg U71289 ( .A(n38563), .B(n21146), .X(n21145) );
  nand_x1_sg U71290 ( .A(n21140), .B(n38564), .X(n21138) );
  nor_x1_sg U71291 ( .A(n38564), .B(n21140), .X(n21139) );
  nand_x1_sg U71292 ( .A(n21134), .B(n38565), .X(n21132) );
  nor_x1_sg U71293 ( .A(n38565), .B(n21134), .X(n21133) );
  nand_x1_sg U71294 ( .A(n21128), .B(n38566), .X(n21126) );
  nor_x1_sg U71295 ( .A(n38566), .B(n21128), .X(n21127) );
  nand_x1_sg U71296 ( .A(n21122), .B(n38567), .X(n21120) );
  nor_x1_sg U71297 ( .A(n38567), .B(n21122), .X(n21121) );
  nand_x1_sg U71298 ( .A(n21116), .B(n38568), .X(n21114) );
  nor_x1_sg U71299 ( .A(n38568), .B(n21116), .X(n21115) );
  nand_x1_sg U71300 ( .A(n21110), .B(n38569), .X(n21108) );
  nor_x1_sg U71301 ( .A(n38569), .B(n21110), .X(n21109) );
  nand_x1_sg U71302 ( .A(n21104), .B(n38570), .X(n21102) );
  nor_x1_sg U71303 ( .A(n38570), .B(n21104), .X(n21103) );
  nand_x1_sg U71304 ( .A(n21098), .B(n38571), .X(n21096) );
  nor_x1_sg U71305 ( .A(n38571), .B(n21098), .X(n21097) );
  nand_x1_sg U71306 ( .A(n21152), .B(n38572), .X(n21150) );
  nor_x1_sg U71307 ( .A(n38572), .B(n21152), .X(n21151) );
  nand_x1_sg U71308 ( .A(n21158), .B(n38573), .X(n21156) );
  nor_x1_sg U71309 ( .A(n38573), .B(n21158), .X(n21157) );
  nand_x1_sg U71310 ( .A(n21164), .B(n38574), .X(n21162) );
  nor_x1_sg U71311 ( .A(n38574), .B(n21164), .X(n21163) );
  nand_x1_sg U71312 ( .A(n20431), .B(n38575), .X(n20429) );
  nor_x1_sg U71313 ( .A(n38575), .B(n20431), .X(n20430) );
  nand_x1_sg U71314 ( .A(n20425), .B(n38576), .X(n20423) );
  nor_x1_sg U71315 ( .A(n38576), .B(n20425), .X(n20424) );
  nand_x1_sg U71316 ( .A(n20419), .B(n38577), .X(n20417) );
  nor_x1_sg U71317 ( .A(n38577), .B(n20419), .X(n20418) );
  nand_x1_sg U71318 ( .A(n20413), .B(n38578), .X(n20411) );
  nor_x1_sg U71319 ( .A(n38578), .B(n20413), .X(n20412) );
  nand_x1_sg U71320 ( .A(n20407), .B(n38579), .X(n20405) );
  nor_x1_sg U71321 ( .A(n38579), .B(n20407), .X(n20406) );
  nand_x1_sg U71322 ( .A(n20401), .B(n38580), .X(n20399) );
  nor_x1_sg U71323 ( .A(n38580), .B(n20401), .X(n20400) );
  nand_x1_sg U71324 ( .A(n20395), .B(n38581), .X(n20393) );
  nor_x1_sg U71325 ( .A(n38581), .B(n20395), .X(n20394) );
  nand_x1_sg U71326 ( .A(n20389), .B(n38582), .X(n20387) );
  nor_x1_sg U71327 ( .A(n38582), .B(n20389), .X(n20388) );
  nand_x1_sg U71328 ( .A(n19698), .B(n38583), .X(n19696) );
  nor_x1_sg U71329 ( .A(n38583), .B(n19698), .X(n19697) );
  nand_x1_sg U71330 ( .A(n19692), .B(n38584), .X(n19690) );
  nor_x1_sg U71331 ( .A(n38584), .B(n19692), .X(n19691) );
  nand_x1_sg U71332 ( .A(n19686), .B(n38585), .X(n19684) );
  nor_x1_sg U71333 ( .A(n38585), .B(n19686), .X(n19685) );
  nand_x1_sg U71334 ( .A(n19680), .B(n38586), .X(n19678) );
  nor_x1_sg U71335 ( .A(n38586), .B(n19680), .X(n19679) );
  nand_x1_sg U71336 ( .A(n19674), .B(n38587), .X(n19672) );
  nor_x1_sg U71337 ( .A(n38587), .B(n19674), .X(n19673) );
  nand_x1_sg U71338 ( .A(n19668), .B(n38588), .X(n19666) );
  nor_x1_sg U71339 ( .A(n38588), .B(n19668), .X(n19667) );
  nand_x1_sg U71340 ( .A(n19662), .B(n38589), .X(n19660) );
  nor_x1_sg U71341 ( .A(n38589), .B(n19662), .X(n19661) );
  nand_x1_sg U71342 ( .A(n19656), .B(n38590), .X(n19654) );
  nor_x1_sg U71343 ( .A(n38590), .B(n19656), .X(n19655) );
  nand_x1_sg U71344 ( .A(n21092), .B(n38591), .X(n21090) );
  nor_x1_sg U71345 ( .A(n38591), .B(n21092), .X(n21091) );
  nand_x1_sg U71346 ( .A(n20383), .B(n38592), .X(n20381) );
  nor_x1_sg U71347 ( .A(n38592), .B(n20383), .X(n20382) );
  nand_x1_sg U71348 ( .A(n19650), .B(n38593), .X(n19648) );
  nor_x1_sg U71349 ( .A(n38593), .B(n19650), .X(n19649) );
  nand_x1_sg U71350 ( .A(n19956), .B(n38594), .X(n20150) );
  nor_x1_sg U71351 ( .A(n38594), .B(n19956), .X(n20151) );
  nand_x1_sg U71352 ( .A(n19773), .B(n38595), .X(n19958) );
  nor_x1_sg U71353 ( .A(n38595), .B(n19773), .X(n19959) );
  nand_x1_sg U71354 ( .A(n20148), .B(n38596), .X(n20311) );
  nor_x1_sg U71355 ( .A(n38596), .B(n20148), .X(n20312) );
  nand_x1_sg U71356 ( .A(n28142), .B(n38128), .X(n28140) );
  nor_x1_sg U71357 ( .A(n38128), .B(n28142), .X(n28141) );
  nand_x1_sg U71358 ( .A(n20508), .B(n38129), .X(n20506) );
  nor_x1_sg U71359 ( .A(n38129), .B(n20508), .X(n20507) );
  nand_x1_sg U71360 ( .A(n19851), .B(n38130), .X(n19849) );
  nor_x1_sg U71361 ( .A(n38130), .B(n19851), .X(n19850) );
  nand_x1_sg U71362 ( .A(n6671), .B(n38131), .X(n6669) );
  nor_x1_sg U71363 ( .A(n38131), .B(n6671), .X(n6670) );
  nand_x1_sg U71364 ( .A(n21277), .B(n38132), .X(n21275) );
  nor_x1_sg U71365 ( .A(n38132), .B(n21277), .X(n21276) );
  nand_x1_sg U71366 ( .A(n40157), .B(n40686), .X(n22861) );
  nand_x1_sg U71367 ( .A(n40360), .B(n40694), .X(n23138) );
  nand_x1_sg U71368 ( .A(n42103), .B(n40696), .X(n23418) );
  nand_x1_sg U71369 ( .A(n42102), .B(n40702), .X(n23697) );
  nand_x1_sg U71370 ( .A(n42101), .B(n40709), .X(n23976) );
  nand_x1_sg U71371 ( .A(n42100), .B(n40711), .X(n24255) );
  nand_x1_sg U71372 ( .A(n42099), .B(n40717), .X(n24534) );
  nand_x1_sg U71373 ( .A(n42098), .B(n40724), .X(n24812) );
  nand_x1_sg U71374 ( .A(n42097), .B(n40726), .X(n25091) );
  nand_x1_sg U71375 ( .A(n40318), .B(n40731), .X(n25370) );
  nand_x1_sg U71376 ( .A(n42094), .B(n40739), .X(n25649) );
  nand_x1_sg U71377 ( .A(n42093), .B(n40744), .X(n26486) );
  nand_x1_sg U71378 ( .A(n21752), .B(n26843), .X(n26840) );
  nand_x1_sg U71379 ( .A(n45751), .B(n45733), .X(n26842) );
  nand_x1_sg U71380 ( .A(n21736), .B(n26858), .X(n26855) );
  nand_x1_sg U71381 ( .A(n45755), .B(n45732), .X(n26857) );
  nand_x1_sg U71382 ( .A(n21731), .B(n26865), .X(n26862) );
  nand_x1_sg U71383 ( .A(n45757), .B(n45731), .X(n26864) );
  nand_x1_sg U71384 ( .A(n21741), .B(n26872), .X(n26869) );
  nand_x1_sg U71385 ( .A(n45759), .B(n45730), .X(n26871) );
  nand_x1_sg U71386 ( .A(n21751), .B(n28563), .X(n28560) );
  nand_x1_sg U71387 ( .A(n45745), .B(n45736), .X(n28562) );
  nand_x1_sg U71388 ( .A(n21735), .B(n26879), .X(n26876) );
  nand_x1_sg U71389 ( .A(n45761), .B(n45729), .X(n26878) );
  nand_x1_sg U71390 ( .A(n5995), .B(n20991), .X(n20988) );
  nand_x1_sg U71391 ( .A(n46585), .B(n46582), .X(n20990) );
  nand_x1_sg U71392 ( .A(n21745), .B(n27087), .X(n28567) );
  nand_x1_sg U71393 ( .A(n45747), .B(n45735), .X(n28569) );
  nand_x1_sg U71394 ( .A(n21746), .B(n28549), .X(n28546) );
  nand_x1_sg U71395 ( .A(n45741), .B(n45738), .X(n28548) );
  nand_x1_sg U71396 ( .A(n21732), .B(n26886), .X(n26883) );
  nand_x1_sg U71397 ( .A(n45763), .B(n45728), .X(n26885) );
  nand_x1_sg U71398 ( .A(n21766), .B(n26836), .X(n26833) );
  nand_x1_sg U71399 ( .A(n45749), .B(n45734), .X(n26835) );
  nand_x1_sg U71400 ( .A(n21767), .B(n28556), .X(n28553) );
  nand_x1_sg U71401 ( .A(n45743), .B(n45737), .X(n28555) );
  nand_x1_sg U71402 ( .A(n21763), .B(n21762), .X(n26897) );
  nand_x1_sg U71403 ( .A(n45767), .B(n45726), .X(n26899) );
  nand_x1_sg U71404 ( .A(n21742), .B(n26893), .X(n26890) );
  nand_x1_sg U71405 ( .A(n45765), .B(n45727), .X(n26892) );
  nand_x1_sg U71406 ( .A(n20999), .B(n46547), .X(n20995) );
  nand_x1_sg U71407 ( .A(n42260), .B(n20998), .X(n20997) );
  nand_x1_sg U71408 ( .A(n26851), .B(n45710), .X(n26847) );
  nand_x1_sg U71409 ( .A(n45753), .B(n26850), .X(n26849) );
  nand_x1_sg U71410 ( .A(n21013), .B(n46580), .X(n21010) );
  nand_x1_sg U71411 ( .A(n42023), .B(n20786), .X(n21012) );
  nand_x1_sg U71412 ( .A(n40070), .B(n40569), .X(n25923) );
  nand_x1_sg U71413 ( .A(n40067), .B(n40618), .X(n26190) );
  nor_x1_sg U71414 ( .A(n42335), .B(n46578), .X(n20588) );
  nor_x1_sg U71415 ( .A(n42334), .B(n19337), .X(n19570) );
  nor_x1_sg U71416 ( .A(n42342), .B(n19145), .X(n19146) );
  nor_x1_sg U71417 ( .A(n5998), .B(n21005), .X(n21006) );
  nand_x1_sg U71418 ( .A(n41099), .B(n22565), .X(n22564) );
  nand_x1_sg U71419 ( .A(n39664), .B(n40316), .X(n7369) );
  nand_x1_sg U71420 ( .A(n39532), .B(n40687), .X(n8187) );
  nand_x1_sg U71421 ( .A(n39533), .B(n40692), .X(n9005) );
  nand_x1_sg U71422 ( .A(n39534), .B(n40699), .X(n9825) );
  nand_x1_sg U71423 ( .A(n39535), .B(n40702), .X(n10644) );
  nand_x1_sg U71424 ( .A(n39536), .B(n40708), .X(n11463) );
  nand_x1_sg U71425 ( .A(n39537), .B(n40711), .X(n12282) );
  nand_x1_sg U71426 ( .A(n39538), .B(n40717), .X(n13101) );
  nand_x1_sg U71427 ( .A(n39539), .B(n40723), .X(n13920) );
  nand_x1_sg U71428 ( .A(n39540), .B(n40726), .X(n14739) );
  nand_x1_sg U71429 ( .A(n39541), .B(n40732), .X(n15558) );
  nand_x1_sg U71430 ( .A(n39542), .B(n40738), .X(n16377) );
  nand_x1_sg U71431 ( .A(n39543), .B(n42044), .X(n18015) );
  nand_x1_sg U71432 ( .A(n39544), .B(n40744), .X(n18836) );
  nand_x1_sg U71433 ( .A(n40081), .B(n40315), .X(n7154) );
  nand_x1_sg U71434 ( .A(n40077), .B(n40568), .X(n16979) );
  nand_x1_sg U71435 ( .A(n39661), .B(n40569), .X(n17194) );
  nand_x1_sg U71436 ( .A(n19909), .B(n6161), .X(n19969) );
  nand_x1_sg U71437 ( .A(n22987), .B(n22988), .X(n22986) );
  nand_x1_sg U71438 ( .A(n23267), .B(n23268), .X(n23266) );
  nand_x1_sg U71439 ( .A(n23546), .B(n23547), .X(n23545) );
  nand_x1_sg U71440 ( .A(n23825), .B(n23826), .X(n23824) );
  nand_x1_sg U71441 ( .A(n24104), .B(n24105), .X(n24103) );
  nand_x1_sg U71442 ( .A(n24383), .B(n24384), .X(n24382) );
  nand_x1_sg U71443 ( .A(n24661), .B(n24662), .X(n24660) );
  nand_x1_sg U71444 ( .A(n24940), .B(n24941), .X(n24939) );
  nand_x1_sg U71445 ( .A(n25219), .B(n25220), .X(n25218) );
  nand_x1_sg U71446 ( .A(n25498), .B(n25499), .X(n25497) );
  nand_x1_sg U71447 ( .A(n25775), .B(n25776), .X(n25774) );
  nand_x1_sg U71448 ( .A(n26335), .B(n26336), .X(n26334) );
  nand_x1_sg U71449 ( .A(n26613), .B(n26614), .X(n26612) );
  nand_x1_sg U71450 ( .A(n19500), .B(n6087), .X(n19576) );
  nand_x1_sg U71451 ( .A(n41306), .B(n40315), .X(n22600) );
  nand_x1_sg U71452 ( .A(n46659), .B(n22992), .X(n22991) );
  nand_x1_sg U71453 ( .A(n46673), .B(n23272), .X(n23271) );
  nand_x1_sg U71454 ( .A(n46687), .B(n23551), .X(n23550) );
  nand_x1_sg U71455 ( .A(n46701), .B(n23830), .X(n23829) );
  nand_x1_sg U71456 ( .A(n46715), .B(n24109), .X(n24108) );
  nand_x1_sg U71457 ( .A(n46729), .B(n24388), .X(n24387) );
  nand_x1_sg U71458 ( .A(n46743), .B(n24666), .X(n24665) );
  nand_x1_sg U71459 ( .A(n46757), .B(n24945), .X(n24944) );
  nand_x1_sg U71460 ( .A(n46771), .B(n25224), .X(n25223) );
  nand_x1_sg U71461 ( .A(n46785), .B(n25503), .X(n25502) );
  nand_x1_sg U71462 ( .A(n46799), .B(n25780), .X(n25779) );
  nand_x1_sg U71463 ( .A(n46826), .B(n26340), .X(n26339) );
  nand_x1_sg U71464 ( .A(n46840), .B(n26618), .X(n26617) );
  nand_x1_sg U71465 ( .A(n40988), .B(n22566), .X(n22563) );
  inv_x1_sg U71466 ( .A(n29154), .X(n45022) );
  inv_x1_sg U71467 ( .A(n21603), .X(n45870) );
  inv_x1_sg U71468 ( .A(n29166), .X(n45112) );
  inv_x1_sg U71469 ( .A(n29178), .X(n45203) );
  inv_x1_sg U71470 ( .A(n29190), .X(n45294) );
  inv_x1_sg U71471 ( .A(n21663), .X(n46326) );
  inv_x1_sg U71472 ( .A(n21651), .X(n46235) );
  inv_x1_sg U71473 ( .A(n21639), .X(n46144) );
  inv_x1_sg U71474 ( .A(n21627), .X(n46053) );
  inv_x1_sg U71475 ( .A(n21615), .X(n45963) );
  inv_x1_sg U71476 ( .A(n29202), .X(n45384) );
  inv_x1_sg U71477 ( .A(n29214), .X(n45474) );
  inv_x1_sg U71478 ( .A(n29089), .X(n45563) );
  inv_x1_sg U71479 ( .A(n21538), .X(n46415) );
  inv_x1_sg U71480 ( .A(n20855), .X(n45826) );
  inv_x1_sg U71481 ( .A(n20212), .X(n45842) );
  inv_x1_sg U71482 ( .A(n19406), .X(n45858) );
  nor_x1_sg U71483 ( .A(n41376), .B(n23130), .X(\L1_0/n4276 ) );
  nand_x1_sg U71484 ( .A(n41316), .B(n40692), .X(n23130) );
  nor_x1_sg U71485 ( .A(n39458), .B(n23410), .X(\L1_0/n4196 ) );
  nand_x1_sg U71486 ( .A(n39475), .B(n40698), .X(n23410) );
  nor_x1_sg U71487 ( .A(n41341), .B(n23689), .X(\L1_0/n4116 ) );
  nand_x1_sg U71488 ( .A(n39928), .B(n40701), .X(n23689) );
  nor_x1_sg U71489 ( .A(n38969), .B(n23968), .X(\L1_0/n4036 ) );
  nand_x1_sg U71490 ( .A(n39277), .B(n40707), .X(n23968) );
  nor_x1_sg U71491 ( .A(n39452), .B(n24247), .X(\L1_0/n3956 ) );
  nand_x1_sg U71492 ( .A(n41315), .B(n40713), .X(n24247) );
  nor_x1_sg U71493 ( .A(n38955), .B(n24526), .X(\L1_0/n3876 ) );
  nand_x1_sg U71494 ( .A(n39279), .B(n40716), .X(n24526) );
  nor_x1_sg U71495 ( .A(n38951), .B(n24804), .X(\L1_0/n3796 ) );
  nand_x1_sg U71496 ( .A(n38943), .B(n40722), .X(n24804) );
  nor_x1_sg U71497 ( .A(n41327), .B(n25083), .X(\L1_0/n3716 ) );
  nand_x1_sg U71498 ( .A(n41462), .B(n40729), .X(n25083) );
  nor_x1_sg U71499 ( .A(n39905), .B(n25362), .X(\L1_0/n3636 ) );
  nand_x1_sg U71500 ( .A(n39276), .B(n40732), .X(n25362) );
  nor_x1_sg U71501 ( .A(n39901), .B(n25641), .X(\L1_0/n3556 ) );
  nand_x1_sg U71502 ( .A(n39929), .B(n40737), .X(n25641) );
  nor_x1_sg U71503 ( .A(n39455), .B(n26478), .X(\L1_0/n3316 ) );
  nand_x1_sg U71504 ( .A(n41316), .B(n40742), .X(n26478) );
  inv_x2_sg U71505 ( .A(n22589), .X(n44975) );
  nor_x1_sg U71506 ( .A(n39962), .B(n7642), .X(\L2_0/n3444 ) );
  nand_x1_sg U71507 ( .A(n41554), .B(n42105), .X(n7642) );
  nor_x1_sg U71508 ( .A(n39966), .B(n8460), .X(\L2_0/n3364 ) );
  nand_x1_sg U71509 ( .A(n41565), .B(n40359), .X(n8460) );
  nor_x1_sg U71510 ( .A(n39970), .B(n9280), .X(\L2_0/n3284 ) );
  nand_x1_sg U71511 ( .A(n41555), .B(n40356), .X(n9280) );
  nor_x1_sg U71512 ( .A(n40703), .B(n10099), .X(\L2_0/n3204 ) );
  nand_x1_sg U71513 ( .A(n41556), .B(n40352), .X(n10099) );
  nor_x1_sg U71514 ( .A(n40708), .B(n10918), .X(\L2_0/n3124 ) );
  nand_x1_sg U71515 ( .A(n41564), .B(n40348), .X(n10918) );
  nor_x1_sg U71516 ( .A(n39982), .B(n11737), .X(\L2_0/n3044 ) );
  nand_x1_sg U71517 ( .A(n41563), .B(n40328), .X(n11737) );
  nor_x1_sg U71518 ( .A(n40718), .B(n12556), .X(\L2_0/n2964 ) );
  nand_x1_sg U71519 ( .A(n41562), .B(n40340), .X(n12556) );
  nor_x1_sg U71520 ( .A(n40723), .B(n13375), .X(\L2_0/n2884 ) );
  nand_x1_sg U71521 ( .A(n41561), .B(n40336), .X(n13375) );
  nor_x1_sg U71522 ( .A(n39994), .B(n14194), .X(\L2_0/n2804 ) );
  nand_x1_sg U71523 ( .A(n41560), .B(n40344), .X(n14194) );
  nor_x1_sg U71524 ( .A(n40733), .B(n15013), .X(\L2_0/n2724 ) );
  nand_x1_sg U71525 ( .A(n41559), .B(n40319), .X(n15013) );
  nor_x1_sg U71526 ( .A(n40738), .B(n15832), .X(\L2_0/n2644 ) );
  nand_x1_sg U71527 ( .A(n41558), .B(n40324), .X(n15832) );
  nor_x1_sg U71528 ( .A(n40617), .B(n51421), .X(\L2_0/n2484 ) );
  nor_x1_sg U71529 ( .A(n17466), .B(n40364), .X(n17470) );
  nor_x1_sg U71530 ( .A(n40743), .B(n18291), .X(\L2_0/n2404 ) );
  nand_x1_sg U71531 ( .A(n41557), .B(n40332), .X(n18291) );
  nand_x1_sg U71532 ( .A(n42185), .B(n40688), .X(n7973) );
  nand_x1_sg U71533 ( .A(n40135), .B(n40693), .X(n8791) );
  nand_x1_sg U71534 ( .A(n40137), .B(n40698), .X(n9611) );
  nand_x1_sg U71535 ( .A(n40139), .B(n40701), .X(n10430) );
  nand_x1_sg U71536 ( .A(n40141), .B(n40708), .X(n11249) );
  nand_x1_sg U71537 ( .A(n40143), .B(n40713), .X(n12068) );
  nand_x1_sg U71538 ( .A(n40145), .B(n40716), .X(n12887) );
  nand_x1_sg U71539 ( .A(n40147), .B(n40723), .X(n13706) );
  nand_x1_sg U71540 ( .A(n40149), .B(n40729), .X(n14525) );
  nand_x1_sg U71541 ( .A(n40151), .B(n40734), .X(n15344) );
  nand_x1_sg U71542 ( .A(n40153), .B(n40738), .X(n16163) );
  nand_x1_sg U71543 ( .A(n40160), .B(n42044), .X(n17801) );
  nand_x1_sg U71544 ( .A(n40156), .B(n40742), .X(n18622) );
  nand_x1_sg U71545 ( .A(n26112), .B(n26113), .X(n26114) );
  nand_x1_sg U71546 ( .A(n23115), .B(n23111), .X(n23116) );
  nand_x1_sg U71547 ( .A(n23395), .B(n23391), .X(n23396) );
  nand_x1_sg U71548 ( .A(n23674), .B(n23670), .X(n23675) );
  nand_x1_sg U71549 ( .A(n23953), .B(n23949), .X(n23954) );
  nand_x1_sg U71550 ( .A(n24232), .B(n24228), .X(n24233) );
  nand_x1_sg U71551 ( .A(n24511), .B(n24507), .X(n24512) );
  nand_x1_sg U71552 ( .A(n24789), .B(n24785), .X(n24790) );
  nand_x1_sg U71553 ( .A(n25068), .B(n25064), .X(n25069) );
  nand_x1_sg U71554 ( .A(n25347), .B(n25343), .X(n25348) );
  nand_x1_sg U71555 ( .A(n25626), .B(n25622), .X(n25627) );
  nand_x1_sg U71556 ( .A(n25903), .B(n25899), .X(n25904) );
  nand_x1_sg U71557 ( .A(n26463), .B(n26459), .X(n26464) );
  nand_x1_sg U71558 ( .A(n26741), .B(n26737), .X(n26742) );
  nand_x1_sg U71559 ( .A(n22838), .B(n22834), .X(n22839) );
  inv_x1_sg U71560 ( .A(n23093), .X(n47143) );
  inv_x1_sg U71561 ( .A(n23373), .X(n47428) );
  inv_x1_sg U71562 ( .A(n23652), .X(n47713) );
  inv_x1_sg U71563 ( .A(n23931), .X(n47998) );
  inv_x1_sg U71564 ( .A(n24210), .X(n48283) );
  inv_x1_sg U71565 ( .A(n24489), .X(n48568) );
  inv_x1_sg U71566 ( .A(n24767), .X(n48853) );
  inv_x1_sg U71567 ( .A(n25046), .X(n49140) );
  inv_x1_sg U71568 ( .A(n25325), .X(n49426) );
  inv_x1_sg U71569 ( .A(n25604), .X(n49712) );
  inv_x1_sg U71570 ( .A(n25881), .X(n49998) );
  inv_x1_sg U71571 ( .A(n26441), .X(n50573) );
  inv_x1_sg U71572 ( .A(n26719), .X(n50859) );
  inv_x1_sg U71573 ( .A(n22513), .X(n45020) );
  inv_x1_sg U71574 ( .A(n42087), .X(n46391) );
  inv_x1_sg U71575 ( .A(n28267), .X(n44994) );
  inv_x1_sg U71576 ( .A(n27984), .X(n45001) );
  inv_x1_sg U71577 ( .A(n27814), .X(n45004) );
  inv_x1_sg U71578 ( .A(n27628), .X(n45007) );
  inv_x1_sg U71579 ( .A(n28635), .X(n44985) );
  inv_x1_sg U71580 ( .A(n27425), .X(n45010) );
  inv_x1_sg U71581 ( .A(n21443), .X(n45815) );
  inv_x1_sg U71582 ( .A(n28474), .X(n44988) );
  inv_x1_sg U71583 ( .A(n28994), .X(n44979) );
  inv_x1_sg U71584 ( .A(n27203), .X(n45013) );
  inv_x1_sg U71585 ( .A(n28380), .X(n44991) );
  inv_x1_sg U71586 ( .A(n28823), .X(n44982) );
  inv_x1_sg U71587 ( .A(n26964), .X(n45016) );
  nand_x1_sg U71588 ( .A(n46802), .B(n26102), .X(n26164) );
  inv_x1_sg U71589 ( .A(n26107), .X(n50283) );
  nor_x1_sg U71590 ( .A(n6800), .B(n6801), .X(n6799) );
  nor_x1_sg U71591 ( .A(n6805), .B(n6806), .X(n6798) );
  nor_x1_sg U71592 ( .A(n39123), .B(n6803), .X(n6800) );
  nor_x1_sg U71593 ( .A(n39249), .B(n26180), .X(\L1_0/n3396 ) );
  nand_x1_sg U71594 ( .A(n39477), .B(n40617), .X(n26180) );
  nand_x1_sg U71595 ( .A(n41111), .B(n22583), .X(n22582) );
  nand_x1_sg U71596 ( .A(n39261), .B(n22584), .X(n22581) );
  inv_x1_sg U71597 ( .A(n22812), .X(n46868) );
  inv_x1_sg U71598 ( .A(n23089), .X(n47161) );
  inv_x1_sg U71599 ( .A(n23369), .X(n47446) );
  inv_x1_sg U71600 ( .A(n23648), .X(n47731) );
  inv_x1_sg U71601 ( .A(n23927), .X(n48016) );
  inv_x1_sg U71602 ( .A(n24206), .X(n48301) );
  inv_x1_sg U71603 ( .A(n24485), .X(n48586) );
  inv_x1_sg U71604 ( .A(n24763), .X(n48872) );
  inv_x1_sg U71605 ( .A(n25042), .X(n49159) );
  inv_x1_sg U71606 ( .A(n25321), .X(n49445) );
  inv_x1_sg U71607 ( .A(n25600), .X(n49730) );
  inv_x1_sg U71608 ( .A(n25877), .X(n50017) );
  inv_x1_sg U71609 ( .A(n26437), .X(n50591) );
  inv_x1_sg U71610 ( .A(n26715), .X(n50878) );
  nand_x1_sg U71611 ( .A(n22588), .B(n44975), .X(n22587) );
  nand_x1_sg U71612 ( .A(n22589), .B(n22590), .X(n22586) );
  nand_x1_sg U71613 ( .A(n40990), .B(n22575), .X(n22572) );
  nand_x1_sg U71614 ( .A(n19118), .B(n22574), .X(n22573) );
  nor_x1_sg U71615 ( .A(n41388), .B(n22853), .X(\L1_0/n4356 ) );
  nand_x1_sg U71616 ( .A(n39927), .B(n40688), .X(n22853) );
  inv_x1_sg U71617 ( .A(n26113), .X(n50279) );
  nand_x1_sg U71618 ( .A(n22549), .B(n22548), .X(n22546) );
  nor_x1_sg U71619 ( .A(n22548), .B(n22549), .X(n22547) );
  nor_x1_sg U71620 ( .A(n26327), .B(n26328), .X(\L1_0/n3320 ) );
  nand_x1_sg U71621 ( .A(n50843), .B(n41051), .X(n26328) );
  nand_x1_sg U71622 ( .A(n21759), .B(n45767), .X(n21757) );
  nor_x1_sg U71623 ( .A(n45767), .B(n21759), .X(n21758) );
  nand_x1_sg U71624 ( .A(n21806), .B(n45724), .X(n21804) );
  nor_x1_sg U71625 ( .A(n45724), .B(n21806), .X(n21805) );
  nand_x1_sg U71626 ( .A(n21853), .B(n45681), .X(n21851) );
  nor_x1_sg U71627 ( .A(n45681), .B(n21853), .X(n21852) );
  nand_x1_sg U71628 ( .A(n21899), .B(n45637), .X(n21897) );
  nor_x1_sg U71629 ( .A(n45637), .B(n21899), .X(n21898) );
  nand_x1_sg U71630 ( .A(n21946), .B(n45593), .X(n21944) );
  nor_x1_sg U71631 ( .A(n45593), .B(n21946), .X(n21945) );
  nand_x1_sg U71632 ( .A(n21992), .B(n45548), .X(n21990) );
  nor_x1_sg U71633 ( .A(n45548), .B(n21992), .X(n21991) );
  nand_x1_sg U71634 ( .A(n22039), .B(n45504), .X(n22037) );
  nor_x1_sg U71635 ( .A(n45504), .B(n22039), .X(n22038) );
  nand_x1_sg U71636 ( .A(n22085), .B(n45456), .X(n22083) );
  nor_x1_sg U71637 ( .A(n45456), .B(n22085), .X(n22084) );
  nand_x1_sg U71638 ( .A(n22133), .B(n45412), .X(n22131) );
  nor_x1_sg U71639 ( .A(n45412), .B(n22133), .X(n22132) );
  nand_x1_sg U71640 ( .A(n22180), .B(n45366), .X(n22178) );
  nor_x1_sg U71641 ( .A(n45366), .B(n22180), .X(n22179) );
  nand_x1_sg U71642 ( .A(n22228), .B(n45321), .X(n22226) );
  nor_x1_sg U71643 ( .A(n45321), .B(n22228), .X(n22227) );
  nand_x1_sg U71644 ( .A(n22275), .B(n45276), .X(n22273) );
  nor_x1_sg U71645 ( .A(n45276), .B(n22275), .X(n22274) );
  nand_x1_sg U71646 ( .A(n22323), .B(n45231), .X(n22321) );
  nor_x1_sg U71647 ( .A(n45231), .B(n22323), .X(n22322) );
  nand_x1_sg U71648 ( .A(n22370), .B(n45185), .X(n22368) );
  nor_x1_sg U71649 ( .A(n45185), .B(n22370), .X(n22369) );
  nand_x1_sg U71650 ( .A(n22418), .B(n45140), .X(n22416) );
  nor_x1_sg U71651 ( .A(n45140), .B(n22418), .X(n22417) );
  nand_x1_sg U71652 ( .A(n22464), .B(n45093), .X(n22462) );
  nor_x1_sg U71653 ( .A(n45093), .B(n22464), .X(n22463) );
  nand_x1_sg U71654 ( .A(n22510), .B(n45049), .X(n22508) );
  nor_x1_sg U71655 ( .A(n45049), .B(n22510), .X(n22509) );
  nand_x1_sg U71656 ( .A(n26796), .B(n26800), .X(n26799) );
  nor_x1_sg U71657 ( .A(n26800), .B(n26796), .X(n26801) );
  inv_x1_sg U71658 ( .A(n29149), .X(n45021) );
  inv_x1_sg U71659 ( .A(n21598), .X(n45869) );
  inv_x1_sg U71660 ( .A(n21186), .X(n46543) );
  inv_x1_sg U71661 ( .A(n28741), .X(n45696) );
  inv_x1_sg U71662 ( .A(n29161), .X(n45066) );
  inv_x1_sg U71663 ( .A(n29173), .X(n45158) );
  inv_x1_sg U71664 ( .A(n29185), .X(n45249) );
  inv_x1_sg U71665 ( .A(n21658), .X(n46281) );
  inv_x1_sg U71666 ( .A(n21646), .X(n46190) );
  inv_x1_sg U71667 ( .A(n21634), .X(n46099) );
  inv_x1_sg U71668 ( .A(n21622), .X(n46008) );
  inv_x1_sg U71669 ( .A(n21610), .X(n45917) );
  inv_x1_sg U71670 ( .A(n6713), .X(n45867) );
  nand_x1_sg U71671 ( .A(n26182), .B(n41050), .X(n26183) );
  nand_x1_sg U71672 ( .A(n26192), .B(n38912), .X(n26193) );
  nand_x1_sg U71673 ( .A(n26200), .B(n38912), .X(n26201) );
  nand_x1_sg U71674 ( .A(n26208), .B(n41050), .X(n26209) );
  nand_x1_sg U71675 ( .A(n26216), .B(n41050), .X(n26217) );
  nand_x1_sg U71676 ( .A(n26224), .B(n41049), .X(n26225) );
  nand_x1_sg U71677 ( .A(n26248), .B(n38912), .X(n26249) );
  nand_x1_sg U71678 ( .A(n26264), .B(n41048), .X(n26265) );
  nand_x1_sg U71679 ( .A(n26280), .B(n41050), .X(n26281) );
  nand_x1_sg U71680 ( .A(n26296), .B(n41049), .X(n26297) );
  nand_x1_sg U71681 ( .A(n26304), .B(n41049), .X(n26305) );
  nand_x1_sg U71682 ( .A(n26310), .B(n41048), .X(n26311) );
  nand_x1_sg U71683 ( .A(n26318), .B(n41048), .X(n26319) );
  nand_x1_sg U71684 ( .A(n38912), .B(n26233), .X(n26232) );
  nand_x1_sg U71685 ( .A(n41051), .B(n26241), .X(n26240) );
  nand_x1_sg U71686 ( .A(n41048), .B(n26257), .X(n26256) );
  nand_x1_sg U71687 ( .A(n41049), .B(n26273), .X(n26272) );
  nand_x1_sg U71688 ( .A(n41051), .B(n26289), .X(n26288) );
  nor_x1_sg U71689 ( .A(n42022), .B(n29275), .X(n29274) );
  nand_x1_sg U71690 ( .A(num[3]), .B(n38834), .X(n38118) );
  nand_x1_sg U71691 ( .A(reg_num[3]), .B(n40395), .X(n38119) );
  nand_x1_sg U71692 ( .A(\yHat[0][6] ), .B(n40834), .X(n36924) );
  nand_x1_sg U71693 ( .A(n40092), .B(\reg_yHat[0][6] ), .X(n36925) );
  nand_x1_sg U71694 ( .A(\yHat[0][18] ), .B(n41494), .X(n36948) );
  nand_x1_sg U71695 ( .A(n40413), .B(\reg_yHat[0][18] ), .X(n36949) );
  nand_x1_sg U71696 ( .A(\yHat[12][6] ), .B(n40833), .X(n37404) );
  nand_x1_sg U71697 ( .A(n40593), .B(\reg_yHat[12][6] ), .X(n37405) );
  nand_x1_sg U71698 ( .A(\yHat[12][18] ), .B(n40834), .X(n37428) );
  nand_x1_sg U71699 ( .A(n40588), .B(\reg_yHat[12][18] ), .X(n37429) );
  nand_x1_sg U71700 ( .A(\y[0][18] ), .B(n40840), .X(n37548) );
  nand_x1_sg U71701 ( .A(n40598), .B(\reg_y[0][18] ), .X(n37549) );
  nand_x1_sg U71702 ( .A(\y[12][18] ), .B(n40828), .X(n38028) );
  nand_x1_sg U71703 ( .A(n40603), .B(\reg_y[12][18] ), .X(n38029) );
  nand_x1_sg U71704 ( .A(\yHat[0][17] ), .B(n41516), .X(n36946) );
  nand_x1_sg U71705 ( .A(\reg_yHat[0][17] ), .B(n40399), .X(n36947) );
  nand_x1_sg U71706 ( .A(\yHat[12][2] ), .B(n38847), .X(n37396) );
  nand_x1_sg U71707 ( .A(\reg_yHat[12][2] ), .B(n41448), .X(n37397) );
  nand_x1_sg U71708 ( .A(\yHat[12][3] ), .B(n40768), .X(n37398) );
  nand_x1_sg U71709 ( .A(\reg_yHat[12][3] ), .B(n39192), .X(n37399) );
  nand_x1_sg U71710 ( .A(\yHat[12][17] ), .B(n41044), .X(n37426) );
  nand_x1_sg U71711 ( .A(\reg_yHat[12][17] ), .B(n40377), .X(n37427) );
  nand_x1_sg U71712 ( .A(\y[0][17] ), .B(n40780), .X(n37546) );
  nand_x1_sg U71713 ( .A(\reg_y[0][17] ), .B(n40382), .X(n37547) );
  nand_x1_sg U71714 ( .A(\y[12][3] ), .B(n40809), .X(n37998) );
  nand_x1_sg U71715 ( .A(\reg_y[12][3] ), .B(n39649), .X(n37999) );
  nand_x1_sg U71716 ( .A(\y[12][17] ), .B(n38843), .X(n38026) );
  nand_x1_sg U71717 ( .A(\reg_y[12][17] ), .B(n40450), .X(n38027) );
  nand_x1_sg U71718 ( .A(num[0]), .B(n41496), .X(n38112) );
  nand_x1_sg U71719 ( .A(reg_num[0]), .B(n40440), .X(n38113) );
  nand_x1_sg U71720 ( .A(\yHat[0][1] ), .B(n39406), .X(n36914) );
  nand_x1_sg U71721 ( .A(\reg_yHat[0][1] ), .B(n40603), .X(n36915) );
  nand_x1_sg U71722 ( .A(\yHat[12][1] ), .B(n40815), .X(n37394) );
  nand_x1_sg U71723 ( .A(\reg_yHat[12][1] ), .B(n40599), .X(n37395) );
  nand_x1_sg U71724 ( .A(\y[0][4] ), .B(n40761), .X(n37520) );
  nand_x1_sg U71725 ( .A(\reg_y[0][4] ), .B(n40405), .X(n37521) );
  nand_x1_sg U71726 ( .A(\y[12][2] ), .B(n38854), .X(n37996) );
  nand_x1_sg U71727 ( .A(\reg_y[12][2] ), .B(n40410), .X(n37997) );
  nand_x1_sg U71728 ( .A(\y[12][4] ), .B(n40811), .X(n38000) );
  nand_x1_sg U71729 ( .A(\reg_y[12][4] ), .B(n38985), .X(n38001) );
  nand_x1_sg U71730 ( .A(\y[0][5] ), .B(n41518), .X(n37522) );
  nand_x1_sg U71731 ( .A(\reg_y[0][5] ), .B(n41474), .X(n37523) );
  nand_x1_sg U71732 ( .A(model), .B(n41503), .X(n36909) );
  nand_x1_sg U71733 ( .A(n41267), .B(n40402), .X(n36910) );
  nand_x1_sg U71734 ( .A(\yHat[0][0] ), .B(n38848), .X(n36912) );
  nand_x1_sg U71735 ( .A(\reg_yHat[0][0] ), .B(n41443), .X(n36913) );
  nand_x1_sg U71736 ( .A(\yHat[0][4] ), .B(n40816), .X(n36920) );
  nand_x1_sg U71737 ( .A(\reg_yHat[0][4] ), .B(n40594), .X(n36921) );
  nand_x1_sg U71738 ( .A(\yHat[0][5] ), .B(n41519), .X(n36922) );
  nand_x1_sg U71739 ( .A(\reg_yHat[0][5] ), .B(n40425), .X(n36923) );
  nand_x1_sg U71740 ( .A(\yHat[0][7] ), .B(n40809), .X(n36926) );
  nand_x1_sg U71741 ( .A(\reg_yHat[0][7] ), .B(n40591), .X(n36927) );
  nand_x1_sg U71742 ( .A(\yHat[0][8] ), .B(n40791), .X(n36928) );
  nand_x1_sg U71743 ( .A(\reg_yHat[0][8] ), .B(n40377), .X(n36929) );
  nand_x1_sg U71744 ( .A(\yHat[0][9] ), .B(n40798), .X(n36930) );
  nand_x1_sg U71745 ( .A(\reg_yHat[0][9] ), .B(n41478), .X(n36931) );
  nand_x1_sg U71746 ( .A(\yHat[0][10] ), .B(n41517), .X(n36932) );
  nand_x1_sg U71747 ( .A(\reg_yHat[0][10] ), .B(n41427), .X(n36933) );
  nand_x1_sg U71748 ( .A(\yHat[0][11] ), .B(n39411), .X(n36934) );
  nand_x1_sg U71749 ( .A(\reg_yHat[0][11] ), .B(n40429), .X(n36935) );
  nand_x1_sg U71750 ( .A(\yHat[0][12] ), .B(n40760), .X(n36936) );
  nand_x1_sg U71751 ( .A(\reg_yHat[0][12] ), .B(n40417), .X(n36937) );
  nand_x1_sg U71752 ( .A(\yHat[0][13] ), .B(n40784), .X(n36938) );
  nand_x1_sg U71753 ( .A(\reg_yHat[0][13] ), .B(n39898), .X(n36939) );
  nand_x1_sg U71754 ( .A(\yHat[0][14] ), .B(n40795), .X(n36940) );
  nand_x1_sg U71755 ( .A(\reg_yHat[0][14] ), .B(n40442), .X(n36941) );
  nand_x1_sg U71756 ( .A(\yHat[0][15] ), .B(n40790), .X(n36942) );
  nand_x1_sg U71757 ( .A(\reg_yHat[0][15] ), .B(n41429), .X(n36943) );
  nand_x1_sg U71758 ( .A(\yHat[0][16] ), .B(n39415), .X(n36944) );
  nand_x1_sg U71759 ( .A(\reg_yHat[0][16] ), .B(n41435), .X(n36945) );
  nand_x1_sg U71760 ( .A(\yHat[0][19] ), .B(n40755), .X(n36950) );
  nand_x1_sg U71761 ( .A(\reg_yHat[0][19] ), .B(n41450), .X(n36951) );
  nand_x1_sg U71762 ( .A(\yHat[12][0] ), .B(n40803), .X(n37392) );
  nand_x1_sg U71763 ( .A(\reg_yHat[12][0] ), .B(n40385), .X(n37393) );
  nand_x1_sg U71764 ( .A(\yHat[12][4] ), .B(n41516), .X(n37400) );
  nand_x1_sg U71765 ( .A(\reg_yHat[12][4] ), .B(n40414), .X(n37401) );
  nand_x1_sg U71766 ( .A(\yHat[12][5] ), .B(n40803), .X(n37402) );
  nand_x1_sg U71767 ( .A(\reg_yHat[12][5] ), .B(n39178), .X(n37403) );
  nand_x1_sg U71768 ( .A(\yHat[12][7] ), .B(n41490), .X(n37406) );
  nand_x1_sg U71769 ( .A(\reg_yHat[12][7] ), .B(n41475), .X(n37407) );
  nand_x1_sg U71770 ( .A(\yHat[12][8] ), .B(n40795), .X(n37408) );
  nand_x1_sg U71771 ( .A(\reg_yHat[12][8] ), .B(n40403), .X(n37409) );
  nand_x1_sg U71772 ( .A(\yHat[12][9] ), .B(n39392), .X(n37410) );
  nand_x1_sg U71773 ( .A(\reg_yHat[12][9] ), .B(n40394), .X(n37411) );
  nand_x1_sg U71774 ( .A(\yHat[12][10] ), .B(n41491), .X(n37412) );
  nand_x1_sg U71775 ( .A(\reg_yHat[12][10] ), .B(n40387), .X(n37413) );
  nand_x1_sg U71776 ( .A(\yHat[12][11] ), .B(n40834), .X(n37414) );
  nand_x1_sg U71777 ( .A(\reg_yHat[12][11] ), .B(n41476), .X(n37415) );
  nand_x1_sg U71778 ( .A(\yHat[12][12] ), .B(n40783), .X(n37416) );
  nand_x1_sg U71779 ( .A(\reg_yHat[12][12] ), .B(n40398), .X(n37417) );
  nand_x1_sg U71780 ( .A(\yHat[12][13] ), .B(n41512), .X(n37418) );
  nand_x1_sg U71781 ( .A(\reg_yHat[12][13] ), .B(n41450), .X(n37419) );
  nand_x1_sg U71782 ( .A(\yHat[12][14] ), .B(n40827), .X(n37420) );
  nand_x1_sg U71783 ( .A(\reg_yHat[12][14] ), .B(n40384), .X(n37421) );
  nand_x1_sg U71784 ( .A(\yHat[12][15] ), .B(n39393), .X(n37422) );
  nand_x1_sg U71785 ( .A(\reg_yHat[12][15] ), .B(n40383), .X(n37423) );
  nand_x1_sg U71786 ( .A(\yHat[12][16] ), .B(n39426), .X(n37424) );
  nand_x1_sg U71787 ( .A(\reg_yHat[12][16] ), .B(n41459), .X(n37425) );
  nand_x1_sg U71788 ( .A(\yHat[12][19] ), .B(n40818), .X(n37430) );
  nand_x1_sg U71789 ( .A(\reg_yHat[12][19] ), .B(n41474), .X(n37431) );
  nand_x1_sg U71790 ( .A(\y[0][0] ), .B(n40780), .X(n37512) );
  nand_x1_sg U71791 ( .A(\reg_y[0][0] ), .B(n39172), .X(n37513) );
  nand_x1_sg U71792 ( .A(\y[0][1] ), .B(n40813), .X(n37514) );
  nand_x1_sg U71793 ( .A(\reg_y[0][1] ), .B(n38987), .X(n37515) );
  nand_x1_sg U71794 ( .A(\y[0][2] ), .B(n39415), .X(n37516) );
  nand_x1_sg U71795 ( .A(\reg_y[0][2] ), .B(n39898), .X(n37517) );
  nand_x1_sg U71796 ( .A(\y[0][3] ), .B(n40768), .X(n37518) );
  nand_x1_sg U71797 ( .A(\reg_y[0][3] ), .B(n41482), .X(n37519) );
  nand_x1_sg U71798 ( .A(\y[0][6] ), .B(n40826), .X(n37524) );
  nand_x1_sg U71799 ( .A(\reg_y[0][6] ), .B(n40446), .X(n37525) );
  nand_x1_sg U71800 ( .A(\y[0][7] ), .B(n39425), .X(n37526) );
  nand_x1_sg U71801 ( .A(\reg_y[0][7] ), .B(n40451), .X(n37527) );
  nand_x1_sg U71802 ( .A(\y[0][8] ), .B(n40803), .X(n37528) );
  nand_x1_sg U71803 ( .A(\reg_y[0][8] ), .B(n40440), .X(n37529) );
  nand_x1_sg U71804 ( .A(\y[0][9] ), .B(n40830), .X(n37530) );
  nand_x1_sg U71805 ( .A(\reg_y[0][9] ), .B(n40425), .X(n37531) );
  nand_x1_sg U71806 ( .A(\y[0][10] ), .B(n39412), .X(n37532) );
  nand_x1_sg U71807 ( .A(\reg_y[0][10] ), .B(n39431), .X(n37533) );
  nand_x1_sg U71808 ( .A(\y[0][11] ), .B(n40835), .X(n37534) );
  nand_x1_sg U71809 ( .A(\reg_y[0][11] ), .B(n40446), .X(n37535) );
  nand_x1_sg U71810 ( .A(\y[0][12] ), .B(n40774), .X(n37536) );
  nand_x1_sg U71811 ( .A(\reg_y[0][12] ), .B(n40435), .X(n37537) );
  nand_x1_sg U71812 ( .A(\y[0][13] ), .B(n39268), .X(n37538) );
  nand_x1_sg U71813 ( .A(\reg_y[0][13] ), .B(n40421), .X(n37539) );
  nand_x1_sg U71814 ( .A(\y[0][14] ), .B(n41511), .X(n37540) );
  nand_x1_sg U71815 ( .A(\reg_y[0][14] ), .B(n40409), .X(n37541) );
  nand_x1_sg U71816 ( .A(\y[0][15] ), .B(n40772), .X(n37542) );
  nand_x1_sg U71817 ( .A(\reg_y[0][15] ), .B(n40406), .X(n37543) );
  nand_x1_sg U71818 ( .A(\y[0][16] ), .B(n41492), .X(n37544) );
  nand_x1_sg U71819 ( .A(\reg_y[0][16] ), .B(n41412), .X(n37545) );
  nand_x1_sg U71820 ( .A(\y[0][19] ), .B(n41521), .X(n37550) );
  nand_x1_sg U71821 ( .A(\reg_y[0][19] ), .B(n41425), .X(n37551) );
  nand_x1_sg U71822 ( .A(\y[12][0] ), .B(n38848), .X(n37992) );
  nand_x1_sg U71823 ( .A(\reg_y[12][0] ), .B(n39167), .X(n37993) );
  nand_x1_sg U71824 ( .A(\y[12][1] ), .B(n40838), .X(n37994) );
  nand_x1_sg U71825 ( .A(\reg_y[12][1] ), .B(n40398), .X(n37995) );
  nand_x1_sg U71826 ( .A(\y[12][5] ), .B(n40794), .X(n38002) );
  nand_x1_sg U71827 ( .A(\reg_y[12][5] ), .B(n41448), .X(n38003) );
  nand_x1_sg U71828 ( .A(\y[12][6] ), .B(n40787), .X(n38004) );
  nand_x1_sg U71829 ( .A(\reg_y[12][6] ), .B(n40434), .X(n38005) );
  nand_x1_sg U71830 ( .A(\y[12][7] ), .B(n40813), .X(n38006) );
  nand_x1_sg U71831 ( .A(\reg_y[12][7] ), .B(n39192), .X(n38007) );
  nand_x1_sg U71832 ( .A(\y[12][8] ), .B(n40778), .X(n38008) );
  nand_x1_sg U71833 ( .A(\reg_y[12][8] ), .B(n40094), .X(n38009) );
  nand_x1_sg U71834 ( .A(\y[12][9] ), .B(n41499), .X(n38010) );
  nand_x1_sg U71835 ( .A(\reg_y[12][9] ), .B(n40606), .X(n38011) );
  nand_x1_sg U71836 ( .A(\y[12][10] ), .B(n41516), .X(n38012) );
  nand_x1_sg U71837 ( .A(\reg_y[12][10] ), .B(n40598), .X(n38013) );
  nand_x1_sg U71838 ( .A(\y[12][11] ), .B(n39410), .X(n38014) );
  nand_x1_sg U71839 ( .A(\reg_y[12][11] ), .B(n40593), .X(n38015) );
  nand_x1_sg U71840 ( .A(\y[12][12] ), .B(n40838), .X(n38016) );
  nand_x1_sg U71841 ( .A(\reg_y[12][12] ), .B(n40378), .X(n38017) );
  nand_x1_sg U71842 ( .A(\y[12][13] ), .B(n39430), .X(n38018) );
  nand_x1_sg U71843 ( .A(\reg_y[12][13] ), .B(n40590), .X(n38019) );
  nand_x1_sg U71844 ( .A(\y[12][14] ), .B(n41509), .X(n38020) );
  nand_x1_sg U71845 ( .A(\reg_y[12][14] ), .B(n41422), .X(n38021) );
  nand_x1_sg U71846 ( .A(\y[12][15] ), .B(n40798), .X(n38022) );
  nand_x1_sg U71847 ( .A(\reg_y[12][15] ), .B(n41425), .X(n38023) );
  nand_x1_sg U71848 ( .A(\y[12][16] ), .B(n39425), .X(n38024) );
  nand_x1_sg U71849 ( .A(\reg_y[12][16] ), .B(n39168), .X(n38025) );
  nand_x1_sg U71850 ( .A(\y[12][19] ), .B(n40768), .X(n38030) );
  nand_x1_sg U71851 ( .A(\reg_y[12][19] ), .B(n40418), .X(n38031) );
  nand_x1_sg U71852 ( .A(num[2]), .B(n41523), .X(n38116) );
  nand_x1_sg U71853 ( .A(reg_num[2]), .B(n40422), .X(n38117) );
  nand_x1_sg U71854 ( .A(\yHat[0][2] ), .B(n38840), .X(n36916) );
  nand_x1_sg U71855 ( .A(\reg_yHat[0][2] ), .B(n40387), .X(n36917) );
  nand_x1_sg U71856 ( .A(\yHat[0][3] ), .B(n40751), .X(n36918) );
  nand_x1_sg U71857 ( .A(\reg_yHat[0][3] ), .B(n39157), .X(n36919) );
  nand_x1_sg U71858 ( .A(num[1]), .B(n41518), .X(n38114) );
  nand_x1_sg U71859 ( .A(reg_num[1]), .B(n40414), .X(n38115) );
  nand_x1_sg U71860 ( .A(\yHat[1][0] ), .B(n40810), .X(n36952) );
  nand_x1_sg U71861 ( .A(\reg_yHat[1][0] ), .B(n40389), .X(n36953) );
  nand_x1_sg U71862 ( .A(\yHat[1][19] ), .B(n40784), .X(n36990) );
  nand_x1_sg U71863 ( .A(\reg_yHat[1][19] ), .B(n41480), .X(n36991) );
  nand_x1_sg U71864 ( .A(\yHat[2][0] ), .B(n40782), .X(n36992) );
  nand_x1_sg U71865 ( .A(\reg_yHat[2][0] ), .B(n41429), .X(n36993) );
  nand_x1_sg U71866 ( .A(\yHat[3][19] ), .B(n39392), .X(n37070) );
  nand_x1_sg U71867 ( .A(\reg_yHat[3][19] ), .B(n40390), .X(n37071) );
  nand_x1_sg U71868 ( .A(\yHat[4][0] ), .B(n40832), .X(n37072) );
  nand_x1_sg U71869 ( .A(\reg_yHat[4][0] ), .B(n40392), .X(n37073) );
  nand_x1_sg U71870 ( .A(\yHat[4][19] ), .B(n39412), .X(n37110) );
  nand_x1_sg U71871 ( .A(\reg_yHat[4][19] ), .B(n41454), .X(n37111) );
  nand_x1_sg U71872 ( .A(\yHat[5][0] ), .B(n40806), .X(n37112) );
  nand_x1_sg U71873 ( .A(\reg_yHat[5][0] ), .B(n41413), .X(n37113) );
  nand_x1_sg U71874 ( .A(\yHat[5][19] ), .B(n40796), .X(n37150) );
  nand_x1_sg U71875 ( .A(\reg_yHat[5][19] ), .B(n41481), .X(n37151) );
  nand_x1_sg U71876 ( .A(\yHat[6][0] ), .B(n39429), .X(n37152) );
  nand_x1_sg U71877 ( .A(\reg_yHat[6][0] ), .B(n39649), .X(n37153) );
  nand_x1_sg U71878 ( .A(\yHat[6][19] ), .B(n40820), .X(n37190) );
  nand_x1_sg U71879 ( .A(\reg_yHat[6][19] ), .B(n40438), .X(n37191) );
  nand_x1_sg U71880 ( .A(\yHat[7][0] ), .B(n40779), .X(n37192) );
  nand_x1_sg U71881 ( .A(\reg_yHat[7][0] ), .B(n41433), .X(n37193) );
  nand_x1_sg U71882 ( .A(\yHat[7][19] ), .B(n41515), .X(n37230) );
  nand_x1_sg U71883 ( .A(\reg_yHat[7][19] ), .B(n41480), .X(n37231) );
  nand_x1_sg U71884 ( .A(\yHat[8][0] ), .B(n40758), .X(n37232) );
  nand_x1_sg U71885 ( .A(\reg_yHat[8][0] ), .B(n40589), .X(n37233) );
  nand_x1_sg U71886 ( .A(\yHat[8][19] ), .B(n40756), .X(n37270) );
  nand_x1_sg U71887 ( .A(\reg_yHat[8][19] ), .B(n40444), .X(n37271) );
  nand_x1_sg U71888 ( .A(\yHat[9][0] ), .B(n40827), .X(n37272) );
  nand_x1_sg U71889 ( .A(\reg_yHat[9][0] ), .B(n40426), .X(n37273) );
  nand_x1_sg U71890 ( .A(\yHat[9][19] ), .B(n41045), .X(n37310) );
  nand_x1_sg U71891 ( .A(\reg_yHat[9][19] ), .B(n40414), .X(n37311) );
  nand_x1_sg U71892 ( .A(\yHat[10][0] ), .B(n40795), .X(n37312) );
  nand_x1_sg U71893 ( .A(\reg_yHat[10][0] ), .B(n41426), .X(n37313) );
  nand_x1_sg U71894 ( .A(\yHat[11][19] ), .B(n40775), .X(n37390) );
  nand_x1_sg U71895 ( .A(\reg_yHat[11][19] ), .B(n41479), .X(n37391) );
  nand_x1_sg U71896 ( .A(\yHat[13][0] ), .B(n41492), .X(n37432) );
  nand_x1_sg U71897 ( .A(\reg_yHat[13][0] ), .B(n41414), .X(n37433) );
  nand_x1_sg U71898 ( .A(\yHat[13][19] ), .B(n40799), .X(n37470) );
  nand_x1_sg U71899 ( .A(\reg_yHat[13][19] ), .B(n40604), .X(n37471) );
  nand_x1_sg U71900 ( .A(\yHat[14][0] ), .B(n40772), .X(n37472) );
  nand_x1_sg U71901 ( .A(\reg_yHat[14][0] ), .B(n40606), .X(n37473) );
  nand_x1_sg U71902 ( .A(\yHat[14][19] ), .B(n40823), .X(n37510) );
  nand_x1_sg U71903 ( .A(\reg_yHat[14][19] ), .B(n40392), .X(n37511) );
  nand_x1_sg U71904 ( .A(\yHat[1][4] ), .B(n41508), .X(n36960) );
  nand_x1_sg U71905 ( .A(\reg_yHat[1][4] ), .B(n41479), .X(n36961) );
  nand_x1_sg U71906 ( .A(\yHat[1][7] ), .B(n41522), .X(n36966) );
  nand_x1_sg U71907 ( .A(\reg_yHat[1][7] ), .B(n40433), .X(n36967) );
  nand_x1_sg U71908 ( .A(\yHat[1][8] ), .B(n40750), .X(n36968) );
  nand_x1_sg U71909 ( .A(\reg_yHat[1][8] ), .B(n40010), .X(n36969) );
  nand_x1_sg U71910 ( .A(\yHat[1][9] ), .B(n40787), .X(n36970) );
  nand_x1_sg U71911 ( .A(\reg_yHat[1][9] ), .B(n41431), .X(n36971) );
  nand_x1_sg U71912 ( .A(\yHat[1][10] ), .B(n39418), .X(n36972) );
  nand_x1_sg U71913 ( .A(\reg_yHat[1][10] ), .B(n40411), .X(n36973) );
  nand_x1_sg U71914 ( .A(\yHat[1][11] ), .B(n40770), .X(n36974) );
  nand_x1_sg U71915 ( .A(\reg_yHat[1][11] ), .B(n41457), .X(n36975) );
  nand_x1_sg U71916 ( .A(\yHat[1][12] ), .B(n40765), .X(n36976) );
  nand_x1_sg U71917 ( .A(\reg_yHat[1][12] ), .B(n41459), .X(n36977) );
  nand_x1_sg U71918 ( .A(\yHat[1][13] ), .B(n40754), .X(n36978) );
  nand_x1_sg U71919 ( .A(\reg_yHat[1][13] ), .B(n41449), .X(n36979) );
  nand_x1_sg U71920 ( .A(\yHat[1][14] ), .B(n40810), .X(n36980) );
  nand_x1_sg U71921 ( .A(\reg_yHat[1][14] ), .B(n40381), .X(n36981) );
  nand_x1_sg U71922 ( .A(\yHat[1][15] ), .B(n40832), .X(n36982) );
  nand_x1_sg U71923 ( .A(\reg_yHat[1][15] ), .B(n40606), .X(n36983) );
  nand_x1_sg U71924 ( .A(\yHat[1][16] ), .B(n40766), .X(n36984) );
  nand_x1_sg U71925 ( .A(\reg_yHat[1][16] ), .B(n41422), .X(n36985) );
  nand_x1_sg U71926 ( .A(\yHat[2][4] ), .B(n40814), .X(n37000) );
  nand_x1_sg U71927 ( .A(\reg_yHat[2][4] ), .B(n39650), .X(n37001) );
  nand_x1_sg U71928 ( .A(\yHat[2][7] ), .B(n40801), .X(n37006) );
  nand_x1_sg U71929 ( .A(\reg_yHat[2][7] ), .B(n40415), .X(n37007) );
  nand_x1_sg U71930 ( .A(\yHat[2][8] ), .B(n39407), .X(n37008) );
  nand_x1_sg U71931 ( .A(\reg_yHat[2][8] ), .B(n39193), .X(n37009) );
  nand_x1_sg U71932 ( .A(\yHat[2][9] ), .B(n41495), .X(n37010) );
  nand_x1_sg U71933 ( .A(\reg_yHat[2][9] ), .B(n40601), .X(n37011) );
  nand_x1_sg U71934 ( .A(\yHat[2][10] ), .B(n40767), .X(n37012) );
  nand_x1_sg U71935 ( .A(\reg_yHat[2][10] ), .B(n40422), .X(n37013) );
  nand_x1_sg U71936 ( .A(\yHat[2][11] ), .B(n40753), .X(n37014) );
  nand_x1_sg U71937 ( .A(\reg_yHat[2][11] ), .B(n39192), .X(n37015) );
  nand_x1_sg U71938 ( .A(\yHat[2][12] ), .B(n40765), .X(n37016) );
  nand_x1_sg U71939 ( .A(\reg_yHat[2][12] ), .B(n40415), .X(n37017) );
  nand_x1_sg U71940 ( .A(\yHat[2][13] ), .B(n40838), .X(n37018) );
  nand_x1_sg U71941 ( .A(\reg_yHat[2][13] ), .B(n40595), .X(n37019) );
  nand_x1_sg U71942 ( .A(\yHat[2][14] ), .B(n41497), .X(n37020) );
  nand_x1_sg U71943 ( .A(\reg_yHat[2][14] ), .B(n40380), .X(n37021) );
  nand_x1_sg U71944 ( .A(\yHat[2][15] ), .B(n40814), .X(n37022) );
  nand_x1_sg U71945 ( .A(\reg_yHat[2][15] ), .B(n38987), .X(n37023) );
  nand_x1_sg U71946 ( .A(\yHat[2][16] ), .B(n40816), .X(n37024) );
  nand_x1_sg U71947 ( .A(\reg_yHat[2][16] ), .B(n41478), .X(n37025) );
  nand_x1_sg U71948 ( .A(\yHat[4][4] ), .B(n40831), .X(n37080) );
  nand_x1_sg U71949 ( .A(\reg_yHat[4][4] ), .B(n39157), .X(n37081) );
  nand_x1_sg U71950 ( .A(\yHat[4][7] ), .B(n41488), .X(n37086) );
  nand_x1_sg U71951 ( .A(\reg_yHat[4][7] ), .B(n40377), .X(n37087) );
  nand_x1_sg U71952 ( .A(\yHat[4][8] ), .B(n41501), .X(n37088) );
  nand_x1_sg U71953 ( .A(\reg_yHat[4][8] ), .B(n40435), .X(n37089) );
  nand_x1_sg U71954 ( .A(\yHat[4][9] ), .B(n40775), .X(n37090) );
  nand_x1_sg U71955 ( .A(\reg_yHat[4][9] ), .B(n40402), .X(n37091) );
  nand_x1_sg U71956 ( .A(\yHat[4][10] ), .B(n41493), .X(n37092) );
  nand_x1_sg U71957 ( .A(\reg_yHat[4][10] ), .B(n40389), .X(n37093) );
  nand_x1_sg U71958 ( .A(\yHat[4][11] ), .B(n40799), .X(n37094) );
  nand_x1_sg U71959 ( .A(\reg_yHat[4][11] ), .B(n40423), .X(n37095) );
  nand_x1_sg U71960 ( .A(\yHat[4][12] ), .B(n40826), .X(n37096) );
  nand_x1_sg U71961 ( .A(\reg_yHat[4][12] ), .B(n41442), .X(n37097) );
  nand_x1_sg U71962 ( .A(\yHat[4][13] ), .B(n40765), .X(n37098) );
  nand_x1_sg U71963 ( .A(\reg_yHat[4][13] ), .B(n41456), .X(n37099) );
  nand_x1_sg U71964 ( .A(\yHat[4][14] ), .B(n40771), .X(n37100) );
  nand_x1_sg U71965 ( .A(\reg_yHat[4][14] ), .B(n40011), .X(n37101) );
  nand_x1_sg U71966 ( .A(\yHat[4][15] ), .B(n39420), .X(n37102) );
  nand_x1_sg U71967 ( .A(\reg_yHat[4][15] ), .B(n41453), .X(n37103) );
  nand_x1_sg U71968 ( .A(\yHat[4][16] ), .B(n39407), .X(n37104) );
  nand_x1_sg U71969 ( .A(\reg_yHat[4][16] ), .B(n41481), .X(n37105) );
  nand_x1_sg U71970 ( .A(\yHat[5][9] ), .B(n39268), .X(n37130) );
  nand_x1_sg U71971 ( .A(\reg_yHat[5][9] ), .B(n39193), .X(n37131) );
  nand_x1_sg U71972 ( .A(\yHat[5][10] ), .B(n39394), .X(n37132) );
  nand_x1_sg U71973 ( .A(\reg_yHat[5][10] ), .B(n41440), .X(n37133) );
  nand_x1_sg U71974 ( .A(\yHat[5][11] ), .B(n40831), .X(n37134) );
  nand_x1_sg U71975 ( .A(\reg_yHat[5][11] ), .B(n40396), .X(n37135) );
  nand_x1_sg U71976 ( .A(\yHat[5][12] ), .B(n41043), .X(n37136) );
  nand_x1_sg U71977 ( .A(\reg_yHat[5][12] ), .B(n40439), .X(n37137) );
  nand_x1_sg U71978 ( .A(\yHat[5][13] ), .B(n40807), .X(n37138) );
  nand_x1_sg U71979 ( .A(\reg_yHat[5][13] ), .B(n41430), .X(n37139) );
  nand_x1_sg U71980 ( .A(\yHat[5][14] ), .B(n40802), .X(n37140) );
  nand_x1_sg U71981 ( .A(\reg_yHat[5][14] ), .B(n39188), .X(n37141) );
  nand_x1_sg U71982 ( .A(\yHat[5][15] ), .B(n39393), .X(n37142) );
  nand_x1_sg U71983 ( .A(\reg_yHat[5][15] ), .B(n41447), .X(n37143) );
  nand_x1_sg U71984 ( .A(\yHat[5][16] ), .B(n39403), .X(n37144) );
  nand_x1_sg U71985 ( .A(\reg_yHat[5][16] ), .B(n40605), .X(n37145) );
  nand_x1_sg U71986 ( .A(\yHat[6][4] ), .B(n41511), .X(n37160) );
  nand_x1_sg U71987 ( .A(\reg_yHat[6][4] ), .B(n40405), .X(n37161) );
  nand_x1_sg U71988 ( .A(\yHat[6][7] ), .B(n39421), .X(n37166) );
  nand_x1_sg U71989 ( .A(\reg_yHat[6][7] ), .B(n39187), .X(n37167) );
  nand_x1_sg U71990 ( .A(\yHat[6][8] ), .B(n41498), .X(n37168) );
  nand_x1_sg U71991 ( .A(\reg_yHat[6][8] ), .B(n40426), .X(n37169) );
  nand_x1_sg U71992 ( .A(\yHat[6][9] ), .B(n40760), .X(n37170) );
  nand_x1_sg U71993 ( .A(\reg_yHat[6][9] ), .B(n41413), .X(n37171) );
  nand_x1_sg U71994 ( .A(\yHat[6][10] ), .B(n40798), .X(n37172) );
  nand_x1_sg U71995 ( .A(\reg_yHat[6][10] ), .B(n40598), .X(n37173) );
  nand_x1_sg U71996 ( .A(\yHat[6][11] ), .B(n40783), .X(n37174) );
  nand_x1_sg U71997 ( .A(\reg_yHat[6][11] ), .B(n40432), .X(n37175) );
  nand_x1_sg U71998 ( .A(\yHat[6][12] ), .B(n40782), .X(n37176) );
  nand_x1_sg U71999 ( .A(\reg_yHat[6][12] ), .B(n39188), .X(n37177) );
  nand_x1_sg U72000 ( .A(\yHat[6][13] ), .B(n40832), .X(n37178) );
  nand_x1_sg U72001 ( .A(\reg_yHat[6][13] ), .B(n41443), .X(n37179) );
  nand_x1_sg U72002 ( .A(\yHat[6][14] ), .B(n40789), .X(n37180) );
  nand_x1_sg U72003 ( .A(\reg_yHat[6][14] ), .B(n41451), .X(n37181) );
  nand_x1_sg U72004 ( .A(\yHat[6][15] ), .B(n39419), .X(n37182) );
  nand_x1_sg U72005 ( .A(\reg_yHat[6][15] ), .B(n39484), .X(n37183) );
  nand_x1_sg U72006 ( .A(\yHat[6][16] ), .B(n41497), .X(n37184) );
  nand_x1_sg U72007 ( .A(\reg_yHat[6][16] ), .B(n40427), .X(n37185) );
  nand_x1_sg U72008 ( .A(\yHat[7][4] ), .B(n40814), .X(n37200) );
  nand_x1_sg U72009 ( .A(\reg_yHat[7][4] ), .B(n41427), .X(n37201) );
  nand_x1_sg U72010 ( .A(\yHat[7][7] ), .B(n41515), .X(n37206) );
  nand_x1_sg U72011 ( .A(\reg_yHat[7][7] ), .B(n40428), .X(n37207) );
  nand_x1_sg U72012 ( .A(\yHat[7][8] ), .B(n40839), .X(n37208) );
  nand_x1_sg U72013 ( .A(\reg_yHat[7][8] ), .B(n40596), .X(n37209) );
  nand_x1_sg U72014 ( .A(\yHat[7][9] ), .B(n40808), .X(n37210) );
  nand_x1_sg U72015 ( .A(\reg_yHat[7][9] ), .B(n40416), .X(n37211) );
  nand_x1_sg U72016 ( .A(\yHat[7][10] ), .B(n40755), .X(n37212) );
  nand_x1_sg U72017 ( .A(\reg_yHat[7][10] ), .B(n40410), .X(n37213) );
  nand_x1_sg U72018 ( .A(\yHat[7][11] ), .B(n41511), .X(n37214) );
  nand_x1_sg U72019 ( .A(\reg_yHat[7][11] ), .B(n39198), .X(n37215) );
  nand_x1_sg U72020 ( .A(\yHat[7][12] ), .B(n40826), .X(n37216) );
  nand_x1_sg U72021 ( .A(\reg_yHat[7][12] ), .B(n40410), .X(n37217) );
  nand_x1_sg U72022 ( .A(\yHat[7][13] ), .B(n40796), .X(n37218) );
  nand_x1_sg U72023 ( .A(\reg_yHat[7][13] ), .B(n40450), .X(n37219) );
  nand_x1_sg U72024 ( .A(\yHat[7][14] ), .B(n40797), .X(n37220) );
  nand_x1_sg U72025 ( .A(\reg_yHat[7][14] ), .B(n40391), .X(n37221) );
  nand_x1_sg U72026 ( .A(\yHat[7][15] ), .B(n40774), .X(n37222) );
  nand_x1_sg U72027 ( .A(\reg_yHat[7][15] ), .B(n40385), .X(n37223) );
  nand_x1_sg U72028 ( .A(\yHat[7][16] ), .B(n39413), .X(n37224) );
  nand_x1_sg U72029 ( .A(\reg_yHat[7][16] ), .B(n40452), .X(n37225) );
  nand_x1_sg U72030 ( .A(\yHat[8][4] ), .B(n38990), .X(n37240) );
  nand_x1_sg U72031 ( .A(\reg_yHat[8][4] ), .B(n40399), .X(n37241) );
  nand_x1_sg U72032 ( .A(\yHat[8][7] ), .B(n40771), .X(n37246) );
  nand_x1_sg U72033 ( .A(\reg_yHat[8][7] ), .B(n40432), .X(n37247) );
  nand_x1_sg U72034 ( .A(\yHat[8][8] ), .B(n40779), .X(n37248) );
  nand_x1_sg U72035 ( .A(\reg_yHat[8][8] ), .B(n40430), .X(n37249) );
  nand_x1_sg U72036 ( .A(\yHat[8][9] ), .B(n40821), .X(n37250) );
  nand_x1_sg U72037 ( .A(\reg_yHat[8][9] ), .B(n40404), .X(n37251) );
  nand_x1_sg U72038 ( .A(\yHat[8][10] ), .B(n41043), .X(n37252) );
  nand_x1_sg U72039 ( .A(\reg_yHat[8][10] ), .B(n40409), .X(n37253) );
  nand_x1_sg U72040 ( .A(\yHat[8][11] ), .B(n41509), .X(n37254) );
  nand_x1_sg U72041 ( .A(\reg_yHat[8][11] ), .B(n41459), .X(n37255) );
  nand_x1_sg U72042 ( .A(\yHat[8][12] ), .B(n38858), .X(n37256) );
  nand_x1_sg U72043 ( .A(\reg_yHat[8][12] ), .B(n41426), .X(n37257) );
  nand_x1_sg U72044 ( .A(\yHat[8][13] ), .B(n41495), .X(n37258) );
  nand_x1_sg U72045 ( .A(\reg_yHat[8][13] ), .B(n40439), .X(n37259) );
  nand_x1_sg U72046 ( .A(\yHat[8][14] ), .B(n40773), .X(n37260) );
  nand_x1_sg U72047 ( .A(\reg_yHat[8][14] ), .B(n41422), .X(n37261) );
  nand_x1_sg U72048 ( .A(\yHat[8][15] ), .B(n40777), .X(n37262) );
  nand_x1_sg U72049 ( .A(\reg_yHat[8][15] ), .B(n38985), .X(n37263) );
  nand_x1_sg U72050 ( .A(\yHat[8][16] ), .B(n40806), .X(n37264) );
  nand_x1_sg U72051 ( .A(\reg_yHat[8][16] ), .B(n39182), .X(n37265) );
  nand_x1_sg U72052 ( .A(\yHat[9][4] ), .B(n40820), .X(n37280) );
  nand_x1_sg U72053 ( .A(\reg_yHat[9][4] ), .B(n39173), .X(n37281) );
  nand_x1_sg U72054 ( .A(\yHat[9][7] ), .B(n41520), .X(n37286) );
  nand_x1_sg U72055 ( .A(\reg_yHat[9][7] ), .B(n41431), .X(n37287) );
  nand_x1_sg U72056 ( .A(\yHat[9][8] ), .B(n38911), .X(n37288) );
  nand_x1_sg U72057 ( .A(\reg_yHat[9][8] ), .B(n41473), .X(n37289) );
  nand_x1_sg U72058 ( .A(\yHat[9][9] ), .B(n41514), .X(n37290) );
  nand_x1_sg U72059 ( .A(\reg_yHat[9][9] ), .B(n39167), .X(n37291) );
  nand_x1_sg U72060 ( .A(\yHat[9][10] ), .B(n40813), .X(n37292) );
  nand_x1_sg U72061 ( .A(\reg_yHat[9][10] ), .B(n40600), .X(n37293) );
  nand_x1_sg U72062 ( .A(\yHat[9][11] ), .B(n39416), .X(n37294) );
  nand_x1_sg U72063 ( .A(\reg_yHat[9][11] ), .B(n40446), .X(n37295) );
  nand_x1_sg U72064 ( .A(\yHat[9][12] ), .B(n41519), .X(n37296) );
  nand_x1_sg U72065 ( .A(\reg_yHat[9][12] ), .B(n40441), .X(n37297) );
  nand_x1_sg U72066 ( .A(\yHat[9][13] ), .B(n39411), .X(n37298) );
  nand_x1_sg U72067 ( .A(\reg_yHat[9][13] ), .B(n40439), .X(n37299) );
  nand_x1_sg U72068 ( .A(\yHat[9][14] ), .B(n40771), .X(n37300) );
  nand_x1_sg U72069 ( .A(\reg_yHat[9][14] ), .B(n40390), .X(n37301) );
  nand_x1_sg U72070 ( .A(\yHat[9][15] ), .B(n40770), .X(n37302) );
  nand_x1_sg U72071 ( .A(\reg_yHat[9][15] ), .B(n39198), .X(n37303) );
  nand_x1_sg U72072 ( .A(\yHat[9][16] ), .B(n38858), .X(n37304) );
  nand_x1_sg U72073 ( .A(\reg_yHat[9][16] ), .B(n40426), .X(n37305) );
  nand_x1_sg U72074 ( .A(\yHat[10][4] ), .B(n41508), .X(n37320) );
  nand_x1_sg U72075 ( .A(\reg_yHat[10][4] ), .B(n41434), .X(n37321) );
  nand_x1_sg U72076 ( .A(\yHat[10][7] ), .B(n39414), .X(n37326) );
  nand_x1_sg U72077 ( .A(\reg_yHat[10][7] ), .B(n41458), .X(n37327) );
  nand_x1_sg U72078 ( .A(\yHat[10][8] ), .B(n40827), .X(n37328) );
  nand_x1_sg U72079 ( .A(\reg_yHat[10][8] ), .B(n40447), .X(n37329) );
  nand_x1_sg U72080 ( .A(\yHat[10][9] ), .B(n41494), .X(n37330) );
  nand_x1_sg U72081 ( .A(\reg_yHat[10][9] ), .B(n41439), .X(n37331) );
  nand_x1_sg U72082 ( .A(\yHat[10][10] ), .B(n39420), .X(n37332) );
  nand_x1_sg U72083 ( .A(\reg_yHat[10][10] ), .B(n41445), .X(n37333) );
  nand_x1_sg U72084 ( .A(\yHat[10][11] ), .B(n40814), .X(n37334) );
  nand_x1_sg U72085 ( .A(\reg_yHat[10][11] ), .B(n40416), .X(n37335) );
  nand_x1_sg U72086 ( .A(\yHat[10][12] ), .B(n41495), .X(n37336) );
  nand_x1_sg U72087 ( .A(\reg_yHat[10][12] ), .B(n40604), .X(n37337) );
  nand_x1_sg U72088 ( .A(\yHat[10][13] ), .B(n40762), .X(n37338) );
  nand_x1_sg U72089 ( .A(\reg_yHat[10][13] ), .B(n39899), .X(n37339) );
  nand_x1_sg U72090 ( .A(\yHat[13][4] ), .B(n40753), .X(n37440) );
  nand_x1_sg U72091 ( .A(\reg_yHat[13][4] ), .B(n41429), .X(n37441) );
  nand_x1_sg U72092 ( .A(\yHat[13][7] ), .B(n40779), .X(n37446) );
  nand_x1_sg U72093 ( .A(\reg_yHat[13][7] ), .B(n41412), .X(n37447) );
  nand_x1_sg U72094 ( .A(\yHat[13][8] ), .B(n39407), .X(n37448) );
  nand_x1_sg U72095 ( .A(\reg_yHat[13][8] ), .B(n40406), .X(n37449) );
  nand_x1_sg U72096 ( .A(\yHat[13][9] ), .B(n40840), .X(n37450) );
  nand_x1_sg U72097 ( .A(\reg_yHat[13][9] ), .B(n40417), .X(n37451) );
  nand_x1_sg U72098 ( .A(\yHat[13][10] ), .B(n38860), .X(n37452) );
  nand_x1_sg U72099 ( .A(\reg_yHat[13][10] ), .B(n39182), .X(n37453) );
  nand_x1_sg U72100 ( .A(\yHat[13][11] ), .B(n40813), .X(n37454) );
  nand_x1_sg U72101 ( .A(\reg_yHat[13][11] ), .B(n40593), .X(n37455) );
  nand_x1_sg U72102 ( .A(\yHat[13][12] ), .B(n39396), .X(n37456) );
  nand_x1_sg U72103 ( .A(\reg_yHat[13][12] ), .B(n41481), .X(n37457) );
  nand_x1_sg U72104 ( .A(\yHat[13][13] ), .B(n40810), .X(n37458) );
  nand_x1_sg U72105 ( .A(\reg_yHat[13][13] ), .B(n41445), .X(n37459) );
  nand_x1_sg U72106 ( .A(\yHat[13][14] ), .B(n41502), .X(n37460) );
  nand_x1_sg U72107 ( .A(\reg_yHat[13][14] ), .B(n41438), .X(n37461) );
  nand_x1_sg U72108 ( .A(\yHat[13][15] ), .B(n40766), .X(n37462) );
  nand_x1_sg U72109 ( .A(\reg_yHat[13][15] ), .B(n41445), .X(n37463) );
  nand_x1_sg U72110 ( .A(\yHat[13][16] ), .B(n40762), .X(n37464) );
  nand_x1_sg U72111 ( .A(\reg_yHat[13][16] ), .B(n41453), .X(n37465) );
  nand_x1_sg U72112 ( .A(\yHat[14][4] ), .B(n40770), .X(n37480) );
  nand_x1_sg U72113 ( .A(\reg_yHat[14][4] ), .B(n40600), .X(n37481) );
  nand_x1_sg U72114 ( .A(\yHat[14][7] ), .B(n39203), .X(n37486) );
  nand_x1_sg U72115 ( .A(\reg_yHat[14][7] ), .B(n39650), .X(n37487) );
  nand_x1_sg U72116 ( .A(\yHat[14][8] ), .B(n39203), .X(n37488) );
  nand_x1_sg U72117 ( .A(\reg_yHat[14][8] ), .B(n40603), .X(n37489) );
  nand_x1_sg U72118 ( .A(\yHat[14][9] ), .B(n39415), .X(n37490) );
  nand_x1_sg U72119 ( .A(\reg_yHat[14][9] ), .B(n40449), .X(n37491) );
  nand_x1_sg U72120 ( .A(\yHat[14][10] ), .B(n40773), .X(n37492) );
  nand_x1_sg U72121 ( .A(\reg_yHat[14][10] ), .B(n41430), .X(n37493) );
  nand_x1_sg U72122 ( .A(\yHat[14][11] ), .B(n41521), .X(n37494) );
  nand_x1_sg U72123 ( .A(\reg_yHat[14][11] ), .B(n40388), .X(n37495) );
  nand_x1_sg U72124 ( .A(\yHat[14][12] ), .B(n40811), .X(n37496) );
  nand_x1_sg U72125 ( .A(\reg_yHat[14][12] ), .B(n41435), .X(n37497) );
  nand_x1_sg U72126 ( .A(\yHat[14][13] ), .B(n40777), .X(n37498) );
  nand_x1_sg U72127 ( .A(\reg_yHat[14][13] ), .B(n41452), .X(n37499) );
  nand_x1_sg U72128 ( .A(\yHat[14][14] ), .B(n40753), .X(n37500) );
  nand_x1_sg U72129 ( .A(\reg_yHat[14][14] ), .B(n40404), .X(n37501) );
  nand_x1_sg U72130 ( .A(\yHat[14][15] ), .B(n40786), .X(n37502) );
  nand_x1_sg U72131 ( .A(\reg_yHat[14][15] ), .B(n40429), .X(n37503) );
  nand_x1_sg U72132 ( .A(\yHat[14][16] ), .B(n40802), .X(n37504) );
  nand_x1_sg U72133 ( .A(\reg_yHat[14][16] ), .B(n41480), .X(n37505) );
  nand_x1_sg U72134 ( .A(\y[1][1] ), .B(n40771), .X(n37554) );
  nand_x1_sg U72135 ( .A(\reg_y[1][1] ), .B(n40595), .X(n37555) );
  nand_x1_sg U72136 ( .A(\y[1][2] ), .B(n39414), .X(n37556) );
  nand_x1_sg U72137 ( .A(\reg_y[1][2] ), .B(n40399), .X(n37557) );
  nand_x1_sg U72138 ( .A(\y[1][7] ), .B(n40755), .X(n37566) );
  nand_x1_sg U72139 ( .A(\reg_y[1][7] ), .B(n40591), .X(n37567) );
  nand_x1_sg U72140 ( .A(\y[1][8] ), .B(n39405), .X(n37568) );
  nand_x1_sg U72141 ( .A(\reg_y[1][8] ), .B(n40427), .X(n37569) );
  nand_x1_sg U72142 ( .A(\y[1][9] ), .B(n40831), .X(n37570) );
  nand_x1_sg U72143 ( .A(\reg_y[1][9] ), .B(n40409), .X(n37571) );
  nand_x1_sg U72144 ( .A(\y[1][10] ), .B(n40751), .X(n37572) );
  nand_x1_sg U72145 ( .A(\reg_y[1][10] ), .B(n40420), .X(n37573) );
  nand_x1_sg U72146 ( .A(\y[1][11] ), .B(n38993), .X(n37574) );
  nand_x1_sg U72147 ( .A(\reg_y[1][11] ), .B(n39162), .X(n37575) );
  nand_x1_sg U72148 ( .A(\y[1][12] ), .B(n40775), .X(n37576) );
  nand_x1_sg U72149 ( .A(\reg_y[1][12] ), .B(n40430), .X(n37577) );
  nand_x1_sg U72150 ( .A(\y[1][13] ), .B(n40785), .X(n37578) );
  nand_x1_sg U72151 ( .A(\reg_y[1][13] ), .B(n39168), .X(n37579) );
  nand_x1_sg U72152 ( .A(\y[1][14] ), .B(n40822), .X(n37580) );
  nand_x1_sg U72153 ( .A(\reg_y[1][14] ), .B(n41474), .X(n37581) );
  nand_x1_sg U72154 ( .A(\y[1][15] ), .B(n41513), .X(n37582) );
  nand_x1_sg U72155 ( .A(\reg_y[1][15] ), .B(n40596), .X(n37583) );
  nand_x1_sg U72156 ( .A(\y[1][16] ), .B(n39402), .X(n37584) );
  nand_x1_sg U72157 ( .A(\reg_y[1][16] ), .B(n40403), .X(n37585) );
  nand_x1_sg U72158 ( .A(\y[2][1] ), .B(n40775), .X(n37594) );
  nand_x1_sg U72159 ( .A(\reg_y[2][1] ), .B(n39158), .X(n37595) );
  nand_x1_sg U72160 ( .A(\y[2][2] ), .B(n40834), .X(n37596) );
  nand_x1_sg U72161 ( .A(\reg_y[2][2] ), .B(n40440), .X(n37597) );
  nand_x1_sg U72162 ( .A(\y[3][9] ), .B(n39394), .X(n37650) );
  nand_x1_sg U72163 ( .A(\reg_y[3][9] ), .B(n41413), .X(n37651) );
  nand_x1_sg U72164 ( .A(\y[3][10] ), .B(n39392), .X(n37652) );
  nand_x1_sg U72165 ( .A(\reg_y[3][10] ), .B(n39483), .X(n37653) );
  nand_x1_sg U72166 ( .A(\y[3][11] ), .B(n38848), .X(n37654) );
  nand_x1_sg U72167 ( .A(\reg_y[3][11] ), .B(n41456), .X(n37655) );
  nand_x1_sg U72168 ( .A(\y[3][12] ), .B(n39404), .X(n37656) );
  nand_x1_sg U72169 ( .A(\reg_y[3][12] ), .B(n39182), .X(n37657) );
  nand_x1_sg U72170 ( .A(\y[3][13] ), .B(n39203), .X(n37658) );
  nand_x1_sg U72171 ( .A(\reg_y[3][13] ), .B(n40414), .X(n37659) );
  nand_x1_sg U72172 ( .A(\y[3][14] ), .B(n41500), .X(n37660) );
  nand_x1_sg U72173 ( .A(\reg_y[3][14] ), .B(n40450), .X(n37661) );
  nand_x1_sg U72174 ( .A(\y[3][15] ), .B(n40802), .X(n37662) );
  nand_x1_sg U72175 ( .A(\reg_y[3][15] ), .B(n41458), .X(n37663) );
  nand_x1_sg U72176 ( .A(\y[3][16] ), .B(n40808), .X(n37664) );
  nand_x1_sg U72177 ( .A(\reg_y[3][16] ), .B(n40092), .X(n37665) );
  nand_x1_sg U72178 ( .A(\y[4][1] ), .B(n40778), .X(n37674) );
  nand_x1_sg U72179 ( .A(\reg_y[4][1] ), .B(n41454), .X(n37675) );
  nand_x1_sg U72180 ( .A(\y[4][2] ), .B(n41510), .X(n37676) );
  nand_x1_sg U72181 ( .A(\reg_y[4][2] ), .B(n41427), .X(n37677) );
  nand_x1_sg U72182 ( .A(\y[4][7] ), .B(n39411), .X(n37686) );
  nand_x1_sg U72183 ( .A(\reg_y[4][7] ), .B(n40387), .X(n37687) );
  nand_x1_sg U72184 ( .A(\y[4][8] ), .B(n40786), .X(n37688) );
  nand_x1_sg U72185 ( .A(\reg_y[4][8] ), .B(n41431), .X(n37689) );
  nand_x1_sg U72186 ( .A(\y[4][9] ), .B(n40760), .X(n37690) );
  nand_x1_sg U72187 ( .A(\reg_y[4][9] ), .B(n40418), .X(n37691) );
  nand_x1_sg U72188 ( .A(\y[4][10] ), .B(n40779), .X(n37692) );
  nand_x1_sg U72189 ( .A(\reg_y[4][10] ), .B(n40421), .X(n37693) );
  nand_x1_sg U72190 ( .A(\y[4][11] ), .B(n38855), .X(n37694) );
  nand_x1_sg U72191 ( .A(\reg_y[4][11] ), .B(n40384), .X(n37695) );
  nand_x1_sg U72192 ( .A(\y[4][12] ), .B(n40766), .X(n37696) );
  nand_x1_sg U72193 ( .A(\reg_y[4][12] ), .B(n39649), .X(n37697) );
  nand_x1_sg U72194 ( .A(\y[4][13] ), .B(n40751), .X(n37698) );
  nand_x1_sg U72195 ( .A(\reg_y[4][13] ), .B(n40395), .X(n37699) );
  nand_x1_sg U72196 ( .A(\y[4][14] ), .B(n41500), .X(n37700) );
  nand_x1_sg U72197 ( .A(\reg_y[4][14] ), .B(n41449), .X(n37701) );
  nand_x1_sg U72198 ( .A(\y[4][15] ), .B(n40803), .X(n37702) );
  nand_x1_sg U72199 ( .A(\reg_y[4][15] ), .B(n40447), .X(n37703) );
  nand_x1_sg U72200 ( .A(\y[4][16] ), .B(n38994), .X(n37704) );
  nand_x1_sg U72201 ( .A(\reg_y[4][16] ), .B(n40601), .X(n37705) );
  nand_x1_sg U72202 ( .A(\y[6][1] ), .B(n40819), .X(n37754) );
  nand_x1_sg U72203 ( .A(\reg_y[6][1] ), .B(n41414), .X(n37755) );
  nand_x1_sg U72204 ( .A(\y[6][2] ), .B(n39416), .X(n37756) );
  nand_x1_sg U72205 ( .A(\reg_y[6][2] ), .B(n40442), .X(n37757) );
  nand_x1_sg U72206 ( .A(\y[6][7] ), .B(n40755), .X(n37766) );
  nand_x1_sg U72207 ( .A(\reg_y[6][7] ), .B(n41435), .X(n37767) );
  nand_x1_sg U72208 ( .A(\y[6][8] ), .B(n40767), .X(n37768) );
  nand_x1_sg U72209 ( .A(\reg_y[6][8] ), .B(n40433), .X(n37769) );
  nand_x1_sg U72210 ( .A(\y[6][9] ), .B(n39395), .X(n37770) );
  nand_x1_sg U72211 ( .A(\reg_y[6][9] ), .B(n40438), .X(n37771) );
  nand_x1_sg U72212 ( .A(\y[6][10] ), .B(n41046), .X(n37772) );
  nand_x1_sg U72213 ( .A(\reg_y[6][10] ), .B(n41454), .X(n37773) );
  nand_x1_sg U72214 ( .A(\y[6][11] ), .B(n39403), .X(n37774) );
  nand_x1_sg U72215 ( .A(\reg_y[6][11] ), .B(n39484), .X(n37775) );
  nand_x1_sg U72216 ( .A(\y[6][12] ), .B(n40811), .X(n37776) );
  nand_x1_sg U72217 ( .A(\reg_y[6][12] ), .B(n40010), .X(n37777) );
  nand_x1_sg U72218 ( .A(\y[6][13] ), .B(n41512), .X(n37778) );
  nand_x1_sg U72219 ( .A(\reg_y[6][13] ), .B(n40418), .X(n37779) );
  nand_x1_sg U72220 ( .A(\y[6][14] ), .B(n40782), .X(n37780) );
  nand_x1_sg U72221 ( .A(\reg_y[6][14] ), .B(n40435), .X(n37781) );
  nand_x1_sg U72222 ( .A(\y[6][15] ), .B(n40833), .X(n37782) );
  nand_x1_sg U72223 ( .A(\reg_y[6][15] ), .B(n40605), .X(n37783) );
  nand_x1_sg U72224 ( .A(\y[6][16] ), .B(n39396), .X(n37784) );
  nand_x1_sg U72225 ( .A(\reg_y[6][16] ), .B(n40378), .X(n37785) );
  nand_x1_sg U72226 ( .A(\y[7][1] ), .B(n39285), .X(n37794) );
  nand_x1_sg U72227 ( .A(\reg_y[7][1] ), .B(n40595), .X(n37795) );
  nand_x1_sg U72228 ( .A(\y[7][2] ), .B(n40839), .X(n37796) );
  nand_x1_sg U72229 ( .A(\reg_y[7][2] ), .B(n40588), .X(n37797) );
  nand_x1_sg U72230 ( .A(\y[7][7] ), .B(n40838), .X(n37806) );
  nand_x1_sg U72231 ( .A(\reg_y[7][7] ), .B(n40438), .X(n37807) );
  nand_x1_sg U72232 ( .A(\y[7][8] ), .B(n40754), .X(n37808) );
  nand_x1_sg U72233 ( .A(\reg_y[7][8] ), .B(n41439), .X(n37809) );
  nand_x1_sg U72234 ( .A(\y[7][9] ), .B(n41513), .X(n37810) );
  nand_x1_sg U72235 ( .A(\reg_y[7][9] ), .B(n39163), .X(n37811) );
  nand_x1_sg U72236 ( .A(\y[7][10] ), .B(n39404), .X(n37812) );
  nand_x1_sg U72237 ( .A(\reg_y[7][10] ), .B(n39172), .X(n37813) );
  nand_x1_sg U72238 ( .A(\y[7][11] ), .B(n40782), .X(n37814) );
  nand_x1_sg U72239 ( .A(\reg_y[7][11] ), .B(n39483), .X(n37815) );
  nand_x1_sg U72240 ( .A(\y[7][12] ), .B(n40767), .X(n37816) );
  nand_x1_sg U72241 ( .A(\reg_y[7][12] ), .B(n40449), .X(n37817) );
  nand_x1_sg U72242 ( .A(\y[7][13] ), .B(n40832), .X(n37818) );
  nand_x1_sg U72243 ( .A(\reg_y[7][13] ), .B(n41457), .X(n37819) );
  nand_x1_sg U72244 ( .A(\y[7][14] ), .B(n40753), .X(n37820) );
  nand_x1_sg U72245 ( .A(\reg_y[7][14] ), .B(n41442), .X(n37821) );
  nand_x1_sg U72246 ( .A(\y[7][15] ), .B(n41498), .X(n37822) );
  nand_x1_sg U72247 ( .A(\reg_y[7][15] ), .B(n40441), .X(n37823) );
  nand_x1_sg U72248 ( .A(\y[7][16] ), .B(n41515), .X(n37824) );
  nand_x1_sg U72249 ( .A(\reg_y[7][16] ), .B(n40413), .X(n37825) );
  nand_x1_sg U72250 ( .A(\y[8][1] ), .B(n40796), .X(n37834) );
  nand_x1_sg U72251 ( .A(\reg_y[8][1] ), .B(n39178), .X(n37835) );
  nand_x1_sg U72252 ( .A(\y[8][2] ), .B(n41523), .X(n37836) );
  nand_x1_sg U72253 ( .A(\reg_y[8][2] ), .B(n39431), .X(n37837) );
  nand_x1_sg U72254 ( .A(\y[8][7] ), .B(n40785), .X(n37846) );
  nand_x1_sg U72255 ( .A(\reg_y[8][7] ), .B(n40411), .X(n37847) );
  nand_x1_sg U72256 ( .A(\y[8][8] ), .B(n39393), .X(n37848) );
  nand_x1_sg U72257 ( .A(\reg_y[8][8] ), .B(n40401), .X(n37849) );
  nand_x1_sg U72258 ( .A(\y[8][9] ), .B(n39272), .X(n37850) );
  nand_x1_sg U72259 ( .A(\reg_y[8][9] ), .B(n40589), .X(n37851) );
  nand_x1_sg U72260 ( .A(\y[8][10] ), .B(n40791), .X(n37852) );
  nand_x1_sg U72261 ( .A(\reg_y[8][10] ), .B(n41473), .X(n37853) );
  nand_x1_sg U72262 ( .A(\y[8][11] ), .B(n39426), .X(n37854) );
  nand_x1_sg U72263 ( .A(\reg_y[8][11] ), .B(n40445), .X(n37855) );
  nand_x1_sg U72264 ( .A(\y[8][12] ), .B(n40759), .X(n37856) );
  nand_x1_sg U72265 ( .A(\reg_y[8][12] ), .B(n39431), .X(n37857) );
  nand_x1_sg U72266 ( .A(\y[8][13] ), .B(n40815), .X(n37858) );
  nand_x1_sg U72267 ( .A(\reg_y[8][13] ), .B(n41479), .X(n37859) );
  nand_x1_sg U72268 ( .A(\y[10][7] ), .B(n41520), .X(n37926) );
  nand_x1_sg U72269 ( .A(\reg_y[10][7] ), .B(n41472), .X(n37927) );
  nand_x1_sg U72270 ( .A(\y[10][8] ), .B(n41511), .X(n37928) );
  nand_x1_sg U72271 ( .A(\reg_y[10][8] ), .B(n41414), .X(n37929) );
  nand_x1_sg U72272 ( .A(\y[10][9] ), .B(n40754), .X(n37930) );
  nand_x1_sg U72273 ( .A(\reg_y[10][9] ), .B(n40593), .X(n37931) );
  nand_x1_sg U72274 ( .A(\y[10][10] ), .B(n41490), .X(n37932) );
  nand_x1_sg U72275 ( .A(\reg_y[10][10] ), .B(n41436), .X(n37933) );
  nand_x1_sg U72276 ( .A(\y[10][11] ), .B(n40754), .X(n37934) );
  nand_x1_sg U72277 ( .A(\reg_y[10][11] ), .B(n40401), .X(n37935) );
  nand_x1_sg U72278 ( .A(\y[10][12] ), .B(n39395), .X(n37936) );
  nand_x1_sg U72279 ( .A(\reg_y[10][12] ), .B(n40387), .X(n37937) );
  nand_x1_sg U72280 ( .A(\y[10][13] ), .B(n40839), .X(n37938) );
  nand_x1_sg U72281 ( .A(\reg_y[10][13] ), .B(n40397), .X(n37939) );
  nand_x1_sg U72282 ( .A(\y[10][14] ), .B(n41490), .X(n37940) );
  nand_x1_sg U72283 ( .A(\reg_y[10][14] ), .B(n40432), .X(n37941) );
  nand_x1_sg U72284 ( .A(\y[10][15] ), .B(n40801), .X(n37942) );
  nand_x1_sg U72285 ( .A(\reg_y[10][15] ), .B(n41438), .X(n37943) );
  nand_x1_sg U72286 ( .A(\y[10][16] ), .B(n40790), .X(n37944) );
  nand_x1_sg U72287 ( .A(\reg_y[10][16] ), .B(n40094), .X(n37945) );
  nand_x1_sg U72288 ( .A(\y[11][1] ), .B(n40808), .X(n37954) );
  nand_x1_sg U72289 ( .A(\reg_y[11][1] ), .B(n39157), .X(n37955) );
  nand_x1_sg U72290 ( .A(\y[11][2] ), .B(n41499), .X(n37956) );
  nand_x1_sg U72291 ( .A(\reg_y[11][2] ), .B(n41444), .X(n37957) );
  nand_x1_sg U72292 ( .A(\y[11][7] ), .B(n40839), .X(n37966) );
  nand_x1_sg U72293 ( .A(\reg_y[11][7] ), .B(n41421), .X(n37967) );
  nand_x1_sg U72294 ( .A(\y[11][8] ), .B(n39417), .X(n37968) );
  nand_x1_sg U72295 ( .A(\reg_y[11][8] ), .B(n40590), .X(n37969) );
  nand_x1_sg U72296 ( .A(\y[11][9] ), .B(n41503), .X(n37970) );
  nand_x1_sg U72297 ( .A(\reg_y[11][9] ), .B(n40437), .X(n37971) );
  nand_x1_sg U72298 ( .A(\y[11][10] ), .B(n40837), .X(n37972) );
  nand_x1_sg U72299 ( .A(\reg_y[11][10] ), .B(n40389), .X(n37973) );
  nand_x1_sg U72300 ( .A(\y[11][11] ), .B(n40806), .X(n37974) );
  nand_x1_sg U72301 ( .A(\reg_y[11][11] ), .B(n41424), .X(n37975) );
  nand_x1_sg U72302 ( .A(\y[11][12] ), .B(n39396), .X(n37976) );
  nand_x1_sg U72303 ( .A(\reg_y[11][12] ), .B(n40391), .X(n37977) );
  nand_x1_sg U72304 ( .A(\y[11][13] ), .B(n41500), .X(n37978) );
  nand_x1_sg U72305 ( .A(\reg_y[11][13] ), .B(n40381), .X(n37979) );
  nand_x1_sg U72306 ( .A(\y[11][14] ), .B(n39419), .X(n37980) );
  nand_x1_sg U72307 ( .A(\reg_y[11][14] ), .B(n40441), .X(n37981) );
  nand_x1_sg U72308 ( .A(\y[11][15] ), .B(n41520), .X(n37982) );
  nand_x1_sg U72309 ( .A(\reg_y[11][15] ), .B(n40392), .X(n37983) );
  nand_x1_sg U72310 ( .A(\y[11][16] ), .B(n40837), .X(n37984) );
  nand_x1_sg U72311 ( .A(\reg_y[11][16] ), .B(n39172), .X(n37985) );
  nand_x1_sg U72312 ( .A(\y[13][1] ), .B(n39410), .X(n38034) );
  nand_x1_sg U72313 ( .A(\reg_y[13][1] ), .B(n41482), .X(n38035) );
  nand_x1_sg U72314 ( .A(\y[13][2] ), .B(n39271), .X(n38036) );
  nand_x1_sg U72315 ( .A(\reg_y[13][2] ), .B(n40011), .X(n38037) );
  nand_x1_sg U72316 ( .A(\y[13][7] ), .B(n39413), .X(n38046) );
  nand_x1_sg U72317 ( .A(\reg_y[13][7] ), .B(n39193), .X(n38047) );
  nand_x1_sg U72318 ( .A(\y[13][8] ), .B(n39404), .X(n38048) );
  nand_x1_sg U72319 ( .A(\reg_y[13][8] ), .B(n40388), .X(n38049) );
  nand_x1_sg U72320 ( .A(\y[13][9] ), .B(n39402), .X(n38050) );
  nand_x1_sg U72321 ( .A(\reg_y[13][9] ), .B(n40011), .X(n38051) );
  nand_x1_sg U72322 ( .A(\y[13][10] ), .B(n39417), .X(n38052) );
  nand_x1_sg U72323 ( .A(\reg_y[13][10] ), .B(n40434), .X(n38053) );
  nand_x1_sg U72324 ( .A(\y[13][11] ), .B(n40789), .X(n38054) );
  nand_x1_sg U72325 ( .A(\reg_y[13][11] ), .B(n40385), .X(n38055) );
  nand_x1_sg U72326 ( .A(\y[13][12] ), .B(n39429), .X(n38056) );
  nand_x1_sg U72327 ( .A(\reg_y[13][12] ), .B(n41440), .X(n38057) );
  nand_x1_sg U72328 ( .A(\y[13][13] ), .B(n39418), .X(n38058) );
  nand_x1_sg U72329 ( .A(\reg_y[13][13] ), .B(n40402), .X(n38059) );
  nand_x1_sg U72330 ( .A(\y[13][14] ), .B(n39271), .X(n38060) );
  nand_x1_sg U72331 ( .A(\reg_y[13][14] ), .B(n41433), .X(n38061) );
  nand_x1_sg U72332 ( .A(\y[13][15] ), .B(n40770), .X(n38062) );
  nand_x1_sg U72333 ( .A(\reg_y[13][15] ), .B(n41425), .X(n38063) );
  nand_x1_sg U72334 ( .A(\y[13][16] ), .B(n40799), .X(n38064) );
  nand_x1_sg U72335 ( .A(\reg_y[13][16] ), .B(n40601), .X(n38065) );
  nand_x1_sg U72336 ( .A(\y[14][1] ), .B(n41502), .X(n38074) );
  nand_x1_sg U72337 ( .A(\reg_y[14][1] ), .B(n40442), .X(n38075) );
  nand_x1_sg U72338 ( .A(\y[14][2] ), .B(n39285), .X(n38076) );
  nand_x1_sg U72339 ( .A(\reg_y[14][2] ), .B(n41415), .X(n38077) );
  nand_x1_sg U72340 ( .A(\y[14][7] ), .B(n40790), .X(n38086) );
  nand_x1_sg U72341 ( .A(\reg_y[14][7] ), .B(n39197), .X(n38087) );
  nand_x1_sg U72342 ( .A(\y[14][8] ), .B(n39414), .X(n38088) );
  nand_x1_sg U72343 ( .A(\reg_y[14][8] ), .B(n41421), .X(n38089) );
  nand_x1_sg U72344 ( .A(\y[14][9] ), .B(n40773), .X(n38090) );
  nand_x1_sg U72345 ( .A(\reg_y[14][9] ), .B(n41415), .X(n38091) );
  nand_x1_sg U72346 ( .A(\y[14][10] ), .B(n38990), .X(n38092) );
  nand_x1_sg U72347 ( .A(\reg_y[14][10] ), .B(n40382), .X(n38093) );
  nand_x1_sg U72348 ( .A(\y[14][11] ), .B(n40801), .X(n38094) );
  nand_x1_sg U72349 ( .A(\reg_y[14][11] ), .B(n40452), .X(n38095) );
  nand_x1_sg U72350 ( .A(\y[14][12] ), .B(n41495), .X(n38096) );
  nand_x1_sg U72351 ( .A(\reg_y[14][12] ), .B(n39192), .X(n38097) );
  nand_x1_sg U72352 ( .A(\y[14][13] ), .B(n39405), .X(n38098) );
  nand_x1_sg U72353 ( .A(\reg_y[14][13] ), .B(n40420), .X(n38099) );
  nand_x1_sg U72354 ( .A(\y[14][14] ), .B(n40802), .X(n38100) );
  nand_x1_sg U72355 ( .A(\reg_y[14][14] ), .B(n41433), .X(n38101) );
  nand_x1_sg U72356 ( .A(\y[14][15] ), .B(n40794), .X(n38102) );
  nand_x1_sg U72357 ( .A(\reg_y[14][15] ), .B(n41426), .X(n38103) );
  nand_x1_sg U72358 ( .A(\y[14][16] ), .B(n41503), .X(n38104) );
  nand_x1_sg U72359 ( .A(\reg_y[14][16] ), .B(n40433), .X(n38105) );
  nand_x1_sg U72360 ( .A(\yHat[1][2] ), .B(n38847), .X(n36956) );
  nand_x1_sg U72361 ( .A(\reg_yHat[1][2] ), .B(n40403), .X(n36957) );
  nand_x1_sg U72362 ( .A(\yHat[1][3] ), .B(n39411), .X(n36958) );
  nand_x1_sg U72363 ( .A(\reg_yHat[1][3] ), .B(n41458), .X(n36959) );
  nand_x1_sg U72364 ( .A(\yHat[2][2] ), .B(n39394), .X(n36996) );
  nand_x1_sg U72365 ( .A(\reg_yHat[2][2] ), .B(n41475), .X(n36997) );
  nand_x1_sg U72366 ( .A(\yHat[2][3] ), .B(n39429), .X(n36998) );
  nand_x1_sg U72367 ( .A(\reg_yHat[2][3] ), .B(n40402), .X(n36999) );
  nand_x1_sg U72368 ( .A(\yHat[4][2] ), .B(n40809), .X(n37076) );
  nand_x1_sg U72369 ( .A(\reg_yHat[4][2] ), .B(n39158), .X(n37077) );
  nand_x1_sg U72370 ( .A(\yHat[4][3] ), .B(n38834), .X(n37078) );
  nand_x1_sg U72371 ( .A(\reg_yHat[4][3] ), .B(n40385), .X(n37079) );
  nand_x1_sg U72372 ( .A(\yHat[5][2] ), .B(n40763), .X(n37116) );
  nand_x1_sg U72373 ( .A(\reg_yHat[5][2] ), .B(n40444), .X(n37117) );
  nand_x1_sg U72374 ( .A(\yHat[5][3] ), .B(n38846), .X(n37118) );
  nand_x1_sg U72375 ( .A(\reg_yHat[5][3] ), .B(n39197), .X(n37119) );
  nand_x1_sg U72376 ( .A(\yHat[6][2] ), .B(n38831), .X(n37156) );
  nand_x1_sg U72377 ( .A(\reg_yHat[6][2] ), .B(n40388), .X(n37157) );
  nand_x1_sg U72378 ( .A(\yHat[6][3] ), .B(n40780), .X(n37158) );
  nand_x1_sg U72379 ( .A(\reg_yHat[6][3] ), .B(n40094), .X(n37159) );
  nand_x1_sg U72380 ( .A(\yHat[7][2] ), .B(n41498), .X(n37196) );
  nand_x1_sg U72381 ( .A(\reg_yHat[7][2] ), .B(n39177), .X(n37197) );
  nand_x1_sg U72382 ( .A(\yHat[7][3] ), .B(n41045), .X(n37198) );
  nand_x1_sg U72383 ( .A(\reg_yHat[7][3] ), .B(n41427), .X(n37199) );
  nand_x1_sg U72384 ( .A(\yHat[8][2] ), .B(n41497), .X(n37236) );
  nand_x1_sg U72385 ( .A(\reg_yHat[8][2] ), .B(n40392), .X(n37237) );
  nand_x1_sg U72386 ( .A(\yHat[8][3] ), .B(n40797), .X(n37238) );
  nand_x1_sg U72387 ( .A(\reg_yHat[8][3] ), .B(n40415), .X(n37239) );
  nand_x1_sg U72388 ( .A(\yHat[9][2] ), .B(n40825), .X(n37276) );
  nand_x1_sg U72389 ( .A(\reg_yHat[9][2] ), .B(n40432), .X(n37277) );
  nand_x1_sg U72390 ( .A(\yHat[9][3] ), .B(n40804), .X(n37278) );
  nand_x1_sg U72391 ( .A(\reg_yHat[9][3] ), .B(n40378), .X(n37279) );
  nand_x1_sg U72392 ( .A(\yHat[10][2] ), .B(n41518), .X(n37316) );
  nand_x1_sg U72393 ( .A(\reg_yHat[10][2] ), .B(n40605), .X(n37317) );
  nand_x1_sg U72394 ( .A(\yHat[10][3] ), .B(n39203), .X(n37318) );
  nand_x1_sg U72395 ( .A(\reg_yHat[10][3] ), .B(n40590), .X(n37319) );
  nand_x1_sg U72396 ( .A(\yHat[13][2] ), .B(n40791), .X(n37436) );
  nand_x1_sg U72397 ( .A(\reg_yHat[13][2] ), .B(n41436), .X(n37437) );
  nand_x1_sg U72398 ( .A(\yHat[13][3] ), .B(n38831), .X(n37438) );
  nand_x1_sg U72399 ( .A(\reg_yHat[13][3] ), .B(n40394), .X(n37439) );
  nand_x1_sg U72400 ( .A(\yHat[14][2] ), .B(n40774), .X(n37476) );
  nand_x1_sg U72401 ( .A(\reg_yHat[14][2] ), .B(n40093), .X(n37477) );
  nand_x1_sg U72402 ( .A(\yHat[14][3] ), .B(n39406), .X(n37478) );
  nand_x1_sg U72403 ( .A(\reg_yHat[14][3] ), .B(n40408), .X(n37479) );
  nand_x1_sg U72404 ( .A(\yHat[1][17] ), .B(n40837), .X(n36986) );
  nand_x1_sg U72405 ( .A(\reg_yHat[1][17] ), .B(n41453), .X(n36987) );
  nand_x1_sg U72406 ( .A(\yHat[2][17] ), .B(n38851), .X(n37026) );
  nand_x1_sg U72407 ( .A(\reg_yHat[2][17] ), .B(n40600), .X(n37027) );
  nand_x1_sg U72408 ( .A(\yHat[4][17] ), .B(n41501), .X(n37106) );
  nand_x1_sg U72409 ( .A(\reg_yHat[4][17] ), .B(n40426), .X(n37107) );
  nand_x1_sg U72410 ( .A(\yHat[5][17] ), .B(n40750), .X(n37146) );
  nand_x1_sg U72411 ( .A(\reg_yHat[5][17] ), .B(n40427), .X(n37147) );
  nand_x1_sg U72412 ( .A(\yHat[6][17] ), .B(n40792), .X(n37186) );
  nand_x1_sg U72413 ( .A(\reg_yHat[6][17] ), .B(n40092), .X(n37187) );
  nand_x1_sg U72414 ( .A(\yHat[7][17] ), .B(n41502), .X(n37226) );
  nand_x1_sg U72415 ( .A(\reg_yHat[7][17] ), .B(n41481), .X(n37227) );
  nand_x1_sg U72416 ( .A(\yHat[8][17] ), .B(n39415), .X(n37266) );
  nand_x1_sg U72417 ( .A(\reg_yHat[8][17] ), .B(n39188), .X(n37267) );
  nand_x1_sg U72418 ( .A(\yHat[9][17] ), .B(n40786), .X(n37306) );
  nand_x1_sg U72419 ( .A(\reg_yHat[9][17] ), .B(n41447), .X(n37307) );
  nand_x1_sg U72420 ( .A(\yHat[13][17] ), .B(n39396), .X(n37466) );
  nand_x1_sg U72421 ( .A(\reg_yHat[13][17] ), .B(n40445), .X(n37467) );
  nand_x1_sg U72422 ( .A(\yHat[14][17] ), .B(n40833), .X(n37506) );
  nand_x1_sg U72423 ( .A(\reg_yHat[14][17] ), .B(n40391), .X(n37507) );
  nand_x1_sg U72424 ( .A(\y[1][17] ), .B(n41488), .X(n37586) );
  nand_x1_sg U72425 ( .A(\reg_y[1][17] ), .B(n39193), .X(n37587) );
  nand_x1_sg U72426 ( .A(\y[3][17] ), .B(n40815), .X(n37666) );
  nand_x1_sg U72427 ( .A(\reg_y[3][17] ), .B(n41473), .X(n37667) );
  nand_x1_sg U72428 ( .A(\y[4][17] ), .B(n39418), .X(n37706) );
  nand_x1_sg U72429 ( .A(\reg_y[4][17] ), .B(n39162), .X(n37707) );
  nand_x1_sg U72430 ( .A(\y[6][17] ), .B(n40758), .X(n37786) );
  nand_x1_sg U72431 ( .A(\reg_y[6][17] ), .B(n40413), .X(n37787) );
  nand_x1_sg U72432 ( .A(\y[7][17] ), .B(n39270), .X(n37826) );
  nand_x1_sg U72433 ( .A(\reg_y[7][17] ), .B(n40433), .X(n37827) );
  nand_x1_sg U72434 ( .A(\y[10][17] ), .B(n40837), .X(n37946) );
  nand_x1_sg U72435 ( .A(\reg_y[10][17] ), .B(n40383), .X(n37947) );
  nand_x1_sg U72436 ( .A(\y[11][17] ), .B(n38846), .X(n37986) );
  nand_x1_sg U72437 ( .A(\reg_y[11][17] ), .B(n40442), .X(n37987) );
  nand_x1_sg U72438 ( .A(\y[13][17] ), .B(n39404), .X(n38066) );
  nand_x1_sg U72439 ( .A(\reg_y[13][17] ), .B(n40394), .X(n38067) );
  nand_x1_sg U72440 ( .A(\y[14][17] ), .B(n41508), .X(n38106) );
  nand_x1_sg U72441 ( .A(\reg_y[14][17] ), .B(n38987), .X(n38107) );
  nand_x1_sg U72442 ( .A(\yHat[1][5] ), .B(n40761), .X(n36962) );
  nand_x1_sg U72443 ( .A(\reg_yHat[1][5] ), .B(n41457), .X(n36963) );
  nand_x1_sg U72444 ( .A(\yHat[2][5] ), .B(n40840), .X(n37002) );
  nand_x1_sg U72445 ( .A(\reg_yHat[2][5] ), .B(n41439), .X(n37003) );
  nand_x1_sg U72446 ( .A(\yHat[4][5] ), .B(n40819), .X(n37082) );
  nand_x1_sg U72447 ( .A(\reg_yHat[4][5] ), .B(n41472), .X(n37083) );
  nand_x1_sg U72448 ( .A(\yHat[6][5] ), .B(n39421), .X(n37162) );
  nand_x1_sg U72449 ( .A(\reg_yHat[6][5] ), .B(n40429), .X(n37163) );
  nand_x1_sg U72450 ( .A(\yHat[7][5] ), .B(n39405), .X(n37202) );
  nand_x1_sg U72451 ( .A(\reg_yHat[7][5] ), .B(n41454), .X(n37203) );
  nand_x1_sg U72452 ( .A(\yHat[8][5] ), .B(n38855), .X(n37242) );
  nand_x1_sg U72453 ( .A(\reg_yHat[8][5] ), .B(n39432), .X(n37243) );
  nand_x1_sg U72454 ( .A(\yHat[9][5] ), .B(n39413), .X(n37282) );
  nand_x1_sg U72455 ( .A(\reg_yHat[9][5] ), .B(n40601), .X(n37283) );
  nand_x1_sg U72456 ( .A(\yHat[10][5] ), .B(n38991), .X(n37322) );
  nand_x1_sg U72457 ( .A(\reg_yHat[10][5] ), .B(n40589), .X(n37323) );
  nand_x1_sg U72458 ( .A(\yHat[13][5] ), .B(n38854), .X(n37442) );
  nand_x1_sg U72459 ( .A(\reg_yHat[13][5] ), .B(n41438), .X(n37443) );
  nand_x1_sg U72460 ( .A(\yHat[14][5] ), .B(n39268), .X(n37482) );
  nand_x1_sg U72461 ( .A(\reg_yHat[14][5] ), .B(n40423), .X(n37483) );
  nand_x1_sg U72462 ( .A(\y[1][3] ), .B(n40791), .X(n37558) );
  nand_x1_sg U72463 ( .A(\reg_y[1][3] ), .B(n40391), .X(n37559) );
  nand_x1_sg U72464 ( .A(\y[1][6] ), .B(n40798), .X(n37564) );
  nand_x1_sg U72465 ( .A(\reg_y[1][6] ), .B(n41452), .X(n37565) );
  nand_x1_sg U72466 ( .A(\y[2][3] ), .B(n41046), .X(n37598) );
  nand_x1_sg U72467 ( .A(\reg_y[2][3] ), .B(n40428), .X(n37599) );
  nand_x1_sg U72468 ( .A(\y[4][3] ), .B(n41514), .X(n37678) );
  nand_x1_sg U72469 ( .A(\reg_y[4][3] ), .B(n40451), .X(n37679) );
  nand_x1_sg U72470 ( .A(\y[4][6] ), .B(n40822), .X(n37684) );
  nand_x1_sg U72471 ( .A(\reg_y[4][6] ), .B(n39163), .X(n37685) );
  nand_x1_sg U72472 ( .A(\y[6][3] ), .B(n40816), .X(n37758) );
  nand_x1_sg U72473 ( .A(\reg_y[6][3] ), .B(n41449), .X(n37759) );
  nand_x1_sg U72474 ( .A(\y[6][6] ), .B(n40807), .X(n37764) );
  nand_x1_sg U72475 ( .A(\reg_y[6][6] ), .B(n41430), .X(n37765) );
  nand_x1_sg U72476 ( .A(\y[7][3] ), .B(n39407), .X(n37798) );
  nand_x1_sg U72477 ( .A(\reg_y[7][3] ), .B(n39649), .X(n37799) );
  nand_x1_sg U72478 ( .A(\y[7][6] ), .B(n40762), .X(n37804) );
  nand_x1_sg U72479 ( .A(\reg_y[7][6] ), .B(n39484), .X(n37805) );
  nand_x1_sg U72480 ( .A(\y[8][3] ), .B(n38846), .X(n37838) );
  nand_x1_sg U72481 ( .A(\reg_y[8][3] ), .B(n40447), .X(n37839) );
  nand_x1_sg U72482 ( .A(\y[8][6] ), .B(n40811), .X(n37844) );
  nand_x1_sg U72483 ( .A(\reg_y[8][6] ), .B(n41435), .X(n37845) );
  nand_x1_sg U72484 ( .A(\y[10][6] ), .B(n40761), .X(n37924) );
  nand_x1_sg U72485 ( .A(\reg_y[10][6] ), .B(n40381), .X(n37925) );
  nand_x1_sg U72486 ( .A(\y[11][3] ), .B(n40804), .X(n37958) );
  nand_x1_sg U72487 ( .A(\reg_y[11][3] ), .B(n39173), .X(n37959) );
  nand_x1_sg U72488 ( .A(\y[11][6] ), .B(n41515), .X(n37964) );
  nand_x1_sg U72489 ( .A(\reg_y[11][6] ), .B(n41450), .X(n37965) );
  nand_x1_sg U72490 ( .A(\y[13][3] ), .B(n40818), .X(n38038) );
  nand_x1_sg U72491 ( .A(\reg_y[13][3] ), .B(n41456), .X(n38039) );
  nand_x1_sg U72492 ( .A(\y[13][6] ), .B(n38858), .X(n38044) );
  nand_x1_sg U72493 ( .A(\reg_y[13][6] ), .B(n40380), .X(n38045) );
  nand_x1_sg U72494 ( .A(\y[14][3] ), .B(n39406), .X(n38078) );
  nand_x1_sg U72495 ( .A(\reg_y[14][3] ), .B(n40417), .X(n38079) );
  nand_x1_sg U72496 ( .A(\y[14][6] ), .B(n40809), .X(n38084) );
  nand_x1_sg U72497 ( .A(\reg_y[14][6] ), .B(n41451), .X(n38085) );
  nand_x1_sg U72498 ( .A(\y[1][4] ), .B(n40823), .X(n37560) );
  nand_x1_sg U72499 ( .A(\reg_y[1][4] ), .B(n40398), .X(n37561) );
  nand_x1_sg U72500 ( .A(\y[4][4] ), .B(n39410), .X(n37680) );
  nand_x1_sg U72501 ( .A(\reg_y[4][4] ), .B(n40408), .X(n37681) );
  nand_x1_sg U72502 ( .A(\y[6][4] ), .B(n39417), .X(n37760) );
  nand_x1_sg U72503 ( .A(\reg_y[6][4] ), .B(n40093), .X(n37761) );
  nand_x1_sg U72504 ( .A(\y[7][4] ), .B(n41491), .X(n37800) );
  nand_x1_sg U72505 ( .A(\reg_y[7][4] ), .B(n41478), .X(n37801) );
  nand_x1_sg U72506 ( .A(\y[8][4] ), .B(n40822), .X(n37840) );
  nand_x1_sg U72507 ( .A(\reg_y[8][4] ), .B(n41415), .X(n37841) );
  nand_x1_sg U72508 ( .A(\y[10][4] ), .B(n40785), .X(n37920) );
  nand_x1_sg U72509 ( .A(\reg_y[10][4] ), .B(n40604), .X(n37921) );
  nand_x1_sg U72510 ( .A(\y[11][4] ), .B(n40756), .X(n37960) );
  nand_x1_sg U72511 ( .A(\reg_y[11][4] ), .B(n40596), .X(n37961) );
  nand_x1_sg U72512 ( .A(\y[13][4] ), .B(n40785), .X(n38040) );
  nand_x1_sg U72513 ( .A(\reg_y[13][4] ), .B(n41453), .X(n38041) );
  nand_x1_sg U72514 ( .A(\y[14][4] ), .B(n40756), .X(n38080) );
  nand_x1_sg U72515 ( .A(\reg_y[14][4] ), .B(n41441), .X(n38081) );
  nand_x1_sg U72516 ( .A(\yHat[1][18] ), .B(n38849), .X(n36988) );
  nand_x1_sg U72517 ( .A(\reg_yHat[1][18] ), .B(n40596), .X(n36989) );
  nand_x1_sg U72518 ( .A(\yHat[2][18] ), .B(n40833), .X(n37028) );
  nand_x1_sg U72519 ( .A(\reg_yHat[2][18] ), .B(n40398), .X(n37029) );
  nand_x1_sg U72520 ( .A(\yHat[4][18] ), .B(n41512), .X(n37108) );
  nand_x1_sg U72521 ( .A(\reg_yHat[4][18] ), .B(n39168), .X(n37109) );
  nand_x1_sg U72522 ( .A(\yHat[5][18] ), .B(n39394), .X(n37148) );
  nand_x1_sg U72523 ( .A(\reg_yHat[5][18] ), .B(n39898), .X(n37149) );
  nand_x1_sg U72524 ( .A(\yHat[6][18] ), .B(n40787), .X(n37188) );
  nand_x1_sg U72525 ( .A(\reg_yHat[6][18] ), .B(n39432), .X(n37189) );
  nand_x1_sg U72526 ( .A(\yHat[7][18] ), .B(n39403), .X(n37228) );
  nand_x1_sg U72527 ( .A(\reg_yHat[7][18] ), .B(n40417), .X(n37229) );
  nand_x1_sg U72528 ( .A(\yHat[8][18] ), .B(n40828), .X(n37268) );
  nand_x1_sg U72529 ( .A(\reg_yHat[8][18] ), .B(n39178), .X(n37269) );
  nand_x1_sg U72530 ( .A(\yHat[9][18] ), .B(n38837), .X(n37308) );
  nand_x1_sg U72531 ( .A(\reg_yHat[9][18] ), .B(n39484), .X(n37309) );
  nand_x1_sg U72532 ( .A(\yHat[13][18] ), .B(n41521), .X(n37468) );
  nand_x1_sg U72533 ( .A(\reg_yHat[13][18] ), .B(n40588), .X(n37469) );
  nand_x1_sg U72534 ( .A(\yHat[14][18] ), .B(n41044), .X(n37508) );
  nand_x1_sg U72535 ( .A(\reg_yHat[14][18] ), .B(n40427), .X(n37509) );
  nand_x1_sg U72536 ( .A(\y[1][0] ), .B(n40821), .X(n37552) );
  nand_x1_sg U72537 ( .A(\reg_y[1][0] ), .B(n40383), .X(n37553) );
  nand_x1_sg U72538 ( .A(\y[1][19] ), .B(n38855), .X(n37590) );
  nand_x1_sg U72539 ( .A(\reg_y[1][19] ), .B(n39183), .X(n37591) );
  nand_x1_sg U72540 ( .A(\y[2][0] ), .B(n41045), .X(n37592) );
  nand_x1_sg U72541 ( .A(\reg_y[2][0] ), .B(n40591), .X(n37593) );
  nand_x1_sg U72542 ( .A(\y[3][19] ), .B(n38911), .X(n37670) );
  nand_x1_sg U72543 ( .A(\reg_y[3][19] ), .B(n40389), .X(n37671) );
  nand_x1_sg U72544 ( .A(\y[4][0] ), .B(n40840), .X(n37672) );
  nand_x1_sg U72545 ( .A(\reg_y[4][0] ), .B(n40406), .X(n37673) );
  nand_x1_sg U72546 ( .A(\y[5][19] ), .B(n41510), .X(n37750) );
  nand_x1_sg U72547 ( .A(\reg_y[5][19] ), .B(n39158), .X(n37751) );
  nand_x1_sg U72548 ( .A(\y[6][0] ), .B(n39403), .X(n37752) );
  nand_x1_sg U72549 ( .A(\reg_y[6][0] ), .B(n40422), .X(n37753) );
  nand_x1_sg U72550 ( .A(\y[6][19] ), .B(n38837), .X(n37790) );
  nand_x1_sg U72551 ( .A(\reg_y[6][19] ), .B(n41441), .X(n37791) );
  nand_x1_sg U72552 ( .A(\y[7][0] ), .B(n38911), .X(n37792) );
  nand_x1_sg U72553 ( .A(\reg_y[7][0] ), .B(n41424), .X(n37793) );
  nand_x1_sg U72554 ( .A(\y[7][19] ), .B(n40761), .X(n37830) );
  nand_x1_sg U72555 ( .A(\reg_y[7][19] ), .B(n39188), .X(n37831) );
  nand_x1_sg U72556 ( .A(\y[8][0] ), .B(n38847), .X(n37832) );
  nand_x1_sg U72557 ( .A(\reg_y[8][0] ), .B(n41482), .X(n37833) );
  nand_x1_sg U72558 ( .A(\y[10][19] ), .B(n39430), .X(n37950) );
  nand_x1_sg U72559 ( .A(\reg_y[10][19] ), .B(n39197), .X(n37951) );
  nand_x1_sg U72560 ( .A(\y[11][0] ), .B(n38993), .X(n37952) );
  nand_x1_sg U72561 ( .A(\reg_y[11][0] ), .B(n41436), .X(n37953) );
  nand_x1_sg U72562 ( .A(\y[11][19] ), .B(n41522), .X(n37990) );
  nand_x1_sg U72563 ( .A(\reg_y[11][19] ), .B(n40382), .X(n37991) );
  nand_x1_sg U72564 ( .A(\y[13][0] ), .B(n41488), .X(n38032) );
  nand_x1_sg U72565 ( .A(\reg_y[13][0] ), .B(n39157), .X(n38033) );
  nand_x1_sg U72566 ( .A(\y[13][19] ), .B(n41502), .X(n38070) );
  nand_x1_sg U72567 ( .A(\reg_y[13][19] ), .B(n41421), .X(n38071) );
  nand_x1_sg U72568 ( .A(\y[14][0] ), .B(n41513), .X(n38072) );
  nand_x1_sg U72569 ( .A(\reg_y[14][0] ), .B(n40434), .X(n38073) );
  nand_x1_sg U72570 ( .A(\y[14][19] ), .B(n39270), .X(n38110) );
  nand_x1_sg U72571 ( .A(\reg_y[14][19] ), .B(n39162), .X(n38111) );
  nand_x1_sg U72572 ( .A(\yHat[1][1] ), .B(n40772), .X(n36954) );
  nand_x1_sg U72573 ( .A(\reg_yHat[1][1] ), .B(n40594), .X(n36955) );
  nand_x1_sg U72574 ( .A(\yHat[2][1] ), .B(n38854), .X(n36994) );
  nand_x1_sg U72575 ( .A(\reg_yHat[2][1] ), .B(n41436), .X(n36995) );
  nand_x1_sg U72576 ( .A(\yHat[4][1] ), .B(n39402), .X(n37074) );
  nand_x1_sg U72577 ( .A(\reg_yHat[4][1] ), .B(n41444), .X(n37075) );
  nand_x1_sg U72578 ( .A(\yHat[5][1] ), .B(n41491), .X(n37114) );
  nand_x1_sg U72579 ( .A(\reg_yHat[5][1] ), .B(n39187), .X(n37115) );
  nand_x1_sg U72580 ( .A(\yHat[6][1] ), .B(n40767), .X(n37154) );
  nand_x1_sg U72581 ( .A(\reg_yHat[6][1] ), .B(n40378), .X(n37155) );
  nand_x1_sg U72582 ( .A(\yHat[7][1] ), .B(n38859), .X(n37194) );
  nand_x1_sg U72583 ( .A(\reg_yHat[7][1] ), .B(n40408), .X(n37195) );
  nand_x1_sg U72584 ( .A(\yHat[8][1] ), .B(n38859), .X(n37234) );
  nand_x1_sg U72585 ( .A(\reg_yHat[8][1] ), .B(n41441), .X(n37235) );
  nand_x1_sg U72586 ( .A(\yHat[9][1] ), .B(n39420), .X(n37274) );
  nand_x1_sg U72587 ( .A(\reg_yHat[9][1] ), .B(n39899), .X(n37275) );
  nand_x1_sg U72588 ( .A(\yHat[10][1] ), .B(n40818), .X(n37314) );
  nand_x1_sg U72589 ( .A(\reg_yHat[10][1] ), .B(n40445), .X(n37315) );
  nand_x1_sg U72590 ( .A(\yHat[13][1] ), .B(n41519), .X(n37434) );
  nand_x1_sg U72591 ( .A(\reg_yHat[13][1] ), .B(n40428), .X(n37435) );
  nand_x1_sg U72592 ( .A(\yHat[14][1] ), .B(n39412), .X(n37474) );
  nand_x1_sg U72593 ( .A(\reg_yHat[14][1] ), .B(n41458), .X(n37475) );
  nand_x1_sg U72594 ( .A(\y[1][5] ), .B(n40825), .X(n37562) );
  nand_x1_sg U72595 ( .A(\reg_y[1][5] ), .B(n40396), .X(n37563) );
  nand_x1_sg U72596 ( .A(\y[1][18] ), .B(n40830), .X(n37588) );
  nand_x1_sg U72597 ( .A(\reg_y[1][18] ), .B(n40416), .X(n37589) );
  nand_x1_sg U72598 ( .A(\y[3][18] ), .B(n38831), .X(n37668) );
  nand_x1_sg U72599 ( .A(\reg_y[3][18] ), .B(n40595), .X(n37669) );
  nand_x1_sg U72600 ( .A(\y[4][5] ), .B(n39271), .X(n37682) );
  nand_x1_sg U72601 ( .A(\reg_y[4][5] ), .B(n39431), .X(n37683) );
  nand_x1_sg U72602 ( .A(\y[4][18] ), .B(n40816), .X(n37708) );
  nand_x1_sg U72603 ( .A(\reg_y[4][18] ), .B(n39167), .X(n37709) );
  nand_x1_sg U72604 ( .A(\y[6][5] ), .B(n40826), .X(n37762) );
  nand_x1_sg U72605 ( .A(\reg_y[6][5] ), .B(n40397), .X(n37763) );
  nand_x1_sg U72606 ( .A(\y[6][18] ), .B(n41043), .X(n37788) );
  nand_x1_sg U72607 ( .A(\reg_y[6][18] ), .B(n40093), .X(n37789) );
  nand_x1_sg U72608 ( .A(\y[7][5] ), .B(n39402), .X(n37802) );
  nand_x1_sg U72609 ( .A(\reg_y[7][5] ), .B(n41440), .X(n37803) );
  nand_x1_sg U72610 ( .A(\y[7][18] ), .B(n41493), .X(n37828) );
  nand_x1_sg U72611 ( .A(\reg_y[7][18] ), .B(n40606), .X(n37829) );
  nand_x1_sg U72612 ( .A(\y[8][5] ), .B(n40797), .X(n37842) );
  nand_x1_sg U72613 ( .A(\reg_y[8][5] ), .B(n40381), .X(n37843) );
  nand_x1_sg U72614 ( .A(\y[10][5] ), .B(n40792), .X(n37922) );
  nand_x1_sg U72615 ( .A(\reg_y[10][5] ), .B(n39172), .X(n37923) );
  nand_x1_sg U72616 ( .A(\y[10][18] ), .B(n41519), .X(n37948) );
  nand_x1_sg U72617 ( .A(\reg_y[10][18] ), .B(n39198), .X(n37949) );
  nand_x1_sg U72618 ( .A(\y[11][5] ), .B(n39405), .X(n37962) );
  nand_x1_sg U72619 ( .A(\reg_y[11][5] ), .B(n40603), .X(n37963) );
  nand_x1_sg U72620 ( .A(\y[11][18] ), .B(n40821), .X(n37988) );
  nand_x1_sg U72621 ( .A(\reg_y[11][18] ), .B(n40380), .X(n37989) );
  nand_x1_sg U72622 ( .A(\y[13][5] ), .B(n40825), .X(n38042) );
  nand_x1_sg U72623 ( .A(\reg_y[13][5] ), .B(n40384), .X(n38043) );
  nand_x1_sg U72624 ( .A(\y[13][18] ), .B(n40756), .X(n38068) );
  nand_x1_sg U72625 ( .A(\reg_y[13][18] ), .B(n41479), .X(n38069) );
  nand_x1_sg U72626 ( .A(\y[14][5] ), .B(n38837), .X(n38082) );
  nand_x1_sg U72627 ( .A(\reg_y[14][5] ), .B(n40418), .X(n38083) );
  nand_x1_sg U72628 ( .A(\y[14][18] ), .B(n39418), .X(n38108) );
  nand_x1_sg U72629 ( .A(\reg_y[14][18] ), .B(n40594), .X(n38109) );
  nand_x1_sg U72630 ( .A(\yHat[1][6] ), .B(n38849), .X(n36964) );
  nand_x1_sg U72631 ( .A(\reg_yHat[1][6] ), .B(n41450), .X(n36965) );
  nand_x1_sg U72632 ( .A(\yHat[2][6] ), .B(n38991), .X(n37004) );
  nand_x1_sg U72633 ( .A(\reg_yHat[2][6] ), .B(n41441), .X(n37005) );
  nand_x1_sg U72634 ( .A(\yHat[4][6] ), .B(n41496), .X(n37084) );
  nand_x1_sg U72635 ( .A(\reg_yHat[4][6] ), .B(n40401), .X(n37085) );
  nand_x1_sg U72636 ( .A(\yHat[6][6] ), .B(n40835), .X(n37164) );
  nand_x1_sg U72637 ( .A(\reg_yHat[6][6] ), .B(n41431), .X(n37165) );
  nand_x1_sg U72638 ( .A(\yHat[7][6] ), .B(n41523), .X(n37204) );
  nand_x1_sg U72639 ( .A(\reg_yHat[7][6] ), .B(n40604), .X(n37205) );
  nand_x1_sg U72640 ( .A(\yHat[8][6] ), .B(n40768), .X(n37244) );
  nand_x1_sg U72641 ( .A(\reg_yHat[8][6] ), .B(n40437), .X(n37245) );
  nand_x1_sg U72642 ( .A(\yHat[9][6] ), .B(n40823), .X(n37284) );
  nand_x1_sg U72643 ( .A(\reg_yHat[9][6] ), .B(n40438), .X(n37285) );
  nand_x1_sg U72644 ( .A(\yHat[10][6] ), .B(n38851), .X(n37324) );
  nand_x1_sg U72645 ( .A(\reg_yHat[10][6] ), .B(n40589), .X(n37325) );
  nand_x1_sg U72646 ( .A(\yHat[13][6] ), .B(n40825), .X(n37444) );
  nand_x1_sg U72647 ( .A(\reg_yHat[13][6] ), .B(n40420), .X(n37445) );
  nand_x1_sg U72648 ( .A(\yHat[14][6] ), .B(n40763), .X(n37484) );
  nand_x1_sg U72649 ( .A(\reg_yHat[14][6] ), .B(n41476), .X(n37485) );
  nand_x1_sg U72650 ( .A(\yHat[3][2] ), .B(n40830), .X(n37036) );
  nand_x1_sg U72651 ( .A(\reg_yHat[3][2] ), .B(n40449), .X(n37037) );
  nand_x1_sg U72652 ( .A(\yHat[3][3] ), .B(n41488), .X(n37038) );
  nand_x1_sg U72653 ( .A(\reg_yHat[3][3] ), .B(n39187), .X(n37039) );
  nand_x1_sg U72654 ( .A(\yHat[11][2] ), .B(n41489), .X(n37356) );
  nand_x1_sg U72655 ( .A(\reg_yHat[11][2] ), .B(n40406), .X(n37357) );
  nand_x1_sg U72656 ( .A(\yHat[11][3] ), .B(n40797), .X(n37358) );
  nand_x1_sg U72657 ( .A(\reg_yHat[11][3] ), .B(n40092), .X(n37359) );
  nand_x1_sg U72658 ( .A(\yHat[3][17] ), .B(n40821), .X(n37066) );
  nand_x1_sg U72659 ( .A(\reg_yHat[3][17] ), .B(n40405), .X(n37067) );
  nand_x1_sg U72660 ( .A(\yHat[10][17] ), .B(n41503), .X(n37346) );
  nand_x1_sg U72661 ( .A(\reg_yHat[10][17] ), .B(n40094), .X(n37347) );
  nand_x1_sg U72662 ( .A(\yHat[11][17] ), .B(n41509), .X(n37386) );
  nand_x1_sg U72663 ( .A(\reg_yHat[11][17] ), .B(n39182), .X(n37387) );
  nand_x1_sg U72664 ( .A(\y[2][17] ), .B(n40786), .X(n37626) );
  nand_x1_sg U72665 ( .A(\reg_y[2][17] ), .B(n41412), .X(n37627) );
  nand_x1_sg U72666 ( .A(\y[5][17] ), .B(n40792), .X(n37746) );
  nand_x1_sg U72667 ( .A(\reg_y[5][17] ), .B(n41412), .X(n37747) );
  nand_x1_sg U72668 ( .A(\y[8][17] ), .B(n39410), .X(n37866) );
  nand_x1_sg U72669 ( .A(\reg_y[8][17] ), .B(n39899), .X(n37867) );
  nand_x1_sg U72670 ( .A(\y[9][17] ), .B(n41494), .X(n37906) );
  nand_x1_sg U72671 ( .A(\reg_y[9][17] ), .B(n41449), .X(n37907) );
  nand_x1_sg U72672 ( .A(\yHat[3][5] ), .B(n41489), .X(n37042) );
  nand_x1_sg U72673 ( .A(\reg_yHat[3][5] ), .B(n40409), .X(n37043) );
  nand_x1_sg U72674 ( .A(\yHat[5][5] ), .B(n38843), .X(n37122) );
  nand_x1_sg U72675 ( .A(\reg_yHat[5][5] ), .B(n41444), .X(n37123) );
  nand_x1_sg U72676 ( .A(\yHat[11][5] ), .B(n40777), .X(n37362) );
  nand_x1_sg U72677 ( .A(\reg_yHat[11][5] ), .B(n40437), .X(n37363) );
  nand_x1_sg U72678 ( .A(\y[2][6] ), .B(n40789), .X(n37604) );
  nand_x1_sg U72679 ( .A(\reg_y[2][6] ), .B(n40588), .X(n37605) );
  nand_x1_sg U72680 ( .A(\y[3][3] ), .B(n38840), .X(n37638) );
  nand_x1_sg U72681 ( .A(\reg_y[3][3] ), .B(n41421), .X(n37639) );
  nand_x1_sg U72682 ( .A(\y[3][6] ), .B(n39425), .X(n37644) );
  nand_x1_sg U72683 ( .A(\reg_y[3][6] ), .B(n39898), .X(n37645) );
  nand_x1_sg U72684 ( .A(\y[5][3] ), .B(n40828), .X(n37718) );
  nand_x1_sg U72685 ( .A(\reg_y[5][3] ), .B(n41434), .X(n37719) );
  nand_x1_sg U72686 ( .A(\y[5][6] ), .B(n38840), .X(n37724) );
  nand_x1_sg U72687 ( .A(\reg_y[5][6] ), .B(n39183), .X(n37725) );
  nand_x1_sg U72688 ( .A(\y[9][3] ), .B(n41514), .X(n37878) );
  nand_x1_sg U72689 ( .A(\reg_y[9][3] ), .B(n41459), .X(n37879) );
  nand_x1_sg U72690 ( .A(\y[9][6] ), .B(n40763), .X(n37884) );
  nand_x1_sg U72691 ( .A(\reg_y[9][6] ), .B(n39168), .X(n37885) );
  nand_x1_sg U72692 ( .A(\y[10][3] ), .B(n40804), .X(n37918) );
  nand_x1_sg U72693 ( .A(\reg_y[10][3] ), .B(n41415), .X(n37919) );
  nand_x1_sg U72694 ( .A(\yHat[2][19] ), .B(n40784), .X(n37030) );
  nand_x1_sg U72695 ( .A(\reg_yHat[2][19] ), .B(n40445), .X(n37031) );
  nand_x1_sg U72696 ( .A(\yHat[3][0] ), .B(n40835), .X(n37032) );
  nand_x1_sg U72697 ( .A(\reg_yHat[3][0] ), .B(n41428), .X(n37033) );
  nand_x1_sg U72698 ( .A(\yHat[10][19] ), .B(n41491), .X(n37350) );
  nand_x1_sg U72699 ( .A(\reg_yHat[10][19] ), .B(n41442), .X(n37351) );
  nand_x1_sg U72700 ( .A(\yHat[11][0] ), .B(n40807), .X(n37352) );
  nand_x1_sg U72701 ( .A(\reg_yHat[11][0] ), .B(n40404), .X(n37353) );
  nand_x1_sg U72702 ( .A(\yHat[3][4] ), .B(n40799), .X(n37040) );
  nand_x1_sg U72703 ( .A(\reg_yHat[3][4] ), .B(n40377), .X(n37041) );
  nand_x1_sg U72704 ( .A(\yHat[3][7] ), .B(n39430), .X(n37046) );
  nand_x1_sg U72705 ( .A(\reg_yHat[3][7] ), .B(n40010), .X(n37047) );
  nand_x1_sg U72706 ( .A(\yHat[3][8] ), .B(n39419), .X(n37048) );
  nand_x1_sg U72707 ( .A(\reg_yHat[3][8] ), .B(n40599), .X(n37049) );
  nand_x1_sg U72708 ( .A(\yHat[3][9] ), .B(n41523), .X(n37050) );
  nand_x1_sg U72709 ( .A(\reg_yHat[3][9] ), .B(n41447), .X(n37051) );
  nand_x1_sg U72710 ( .A(\yHat[3][10] ), .B(n39393), .X(n37052) );
  nand_x1_sg U72711 ( .A(\reg_yHat[3][10] ), .B(n40396), .X(n37053) );
  nand_x1_sg U72712 ( .A(\yHat[3][11] ), .B(n40794), .X(n37054) );
  nand_x1_sg U72713 ( .A(\reg_yHat[3][11] ), .B(n40403), .X(n37055) );
  nand_x1_sg U72714 ( .A(\yHat[3][12] ), .B(n40827), .X(n37056) );
  nand_x1_sg U72715 ( .A(\reg_yHat[3][12] ), .B(n40422), .X(n37057) );
  nand_x1_sg U72716 ( .A(\yHat[3][13] ), .B(n40759), .X(n37058) );
  nand_x1_sg U72717 ( .A(\reg_yHat[3][13] ), .B(n40093), .X(n37059) );
  nand_x1_sg U72718 ( .A(\yHat[3][14] ), .B(n40783), .X(n37060) );
  nand_x1_sg U72719 ( .A(\reg_yHat[3][14] ), .B(n41451), .X(n37061) );
  nand_x1_sg U72720 ( .A(\yHat[3][15] ), .B(n40815), .X(n37062) );
  nand_x1_sg U72721 ( .A(\reg_yHat[3][15] ), .B(n41482), .X(n37063) );
  nand_x1_sg U72722 ( .A(\yHat[3][16] ), .B(n41522), .X(n37064) );
  nand_x1_sg U72723 ( .A(\reg_yHat[3][16] ), .B(n40450), .X(n37065) );
  nand_x1_sg U72724 ( .A(\yHat[5][4] ), .B(n40750), .X(n37120) );
  nand_x1_sg U72725 ( .A(\reg_yHat[5][4] ), .B(n40395), .X(n37121) );
  nand_x1_sg U72726 ( .A(\yHat[5][7] ), .B(n40801), .X(n37126) );
  nand_x1_sg U72727 ( .A(\reg_yHat[5][7] ), .B(n40444), .X(n37127) );
  nand_x1_sg U72728 ( .A(\yHat[5][8] ), .B(n39395), .X(n37128) );
  nand_x1_sg U72729 ( .A(\reg_yHat[5][8] ), .B(n40405), .X(n37129) );
  nand_x1_sg U72730 ( .A(\yHat[10][14] ), .B(n40774), .X(n37340) );
  nand_x1_sg U72731 ( .A(\reg_yHat[10][14] ), .B(n39432), .X(n37341) );
  nand_x1_sg U72732 ( .A(\yHat[10][15] ), .B(n40784), .X(n37342) );
  nand_x1_sg U72733 ( .A(\reg_yHat[10][15] ), .B(n39483), .X(n37343) );
  nand_x1_sg U72734 ( .A(\yHat[10][16] ), .B(n40783), .X(n37344) );
  nand_x1_sg U72735 ( .A(\reg_yHat[10][16] ), .B(n40420), .X(n37345) );
  nand_x1_sg U72736 ( .A(\yHat[11][4] ), .B(n40789), .X(n37360) );
  nand_x1_sg U72737 ( .A(\reg_yHat[11][4] ), .B(n40423), .X(n37361) );
  nand_x1_sg U72738 ( .A(\yHat[11][7] ), .B(n39421), .X(n37366) );
  nand_x1_sg U72739 ( .A(\reg_yHat[11][7] ), .B(n40388), .X(n37367) );
  nand_x1_sg U72740 ( .A(\yHat[11][8] ), .B(n40759), .X(n37368) );
  nand_x1_sg U72741 ( .A(\reg_yHat[11][8] ), .B(n40408), .X(n37369) );
  nand_x1_sg U72742 ( .A(\yHat[11][9] ), .B(n41518), .X(n37370) );
  nand_x1_sg U72743 ( .A(\reg_yHat[11][9] ), .B(n39167), .X(n37371) );
  nand_x1_sg U72744 ( .A(\yHat[11][10] ), .B(n40778), .X(n37372) );
  nand_x1_sg U72745 ( .A(\reg_yHat[11][10] ), .B(n40434), .X(n37373) );
  nand_x1_sg U72746 ( .A(\yHat[11][11] ), .B(n40766), .X(n37374) );
  nand_x1_sg U72747 ( .A(\reg_yHat[11][11] ), .B(n41452), .X(n37375) );
  nand_x1_sg U72748 ( .A(\yHat[11][12] ), .B(n38860), .X(n37376) );
  nand_x1_sg U72749 ( .A(\reg_yHat[11][12] ), .B(n40401), .X(n37377) );
  nand_x1_sg U72750 ( .A(\yHat[11][13] ), .B(n39429), .X(n37378) );
  nand_x1_sg U72751 ( .A(\reg_yHat[11][13] ), .B(n41430), .X(n37379) );
  nand_x1_sg U72752 ( .A(\yHat[11][14] ), .B(n41045), .X(n37380) );
  nand_x1_sg U72753 ( .A(\reg_yHat[11][14] ), .B(n39899), .X(n37381) );
  nand_x1_sg U72754 ( .A(\yHat[11][15] ), .B(n40758), .X(n37382) );
  nand_x1_sg U72755 ( .A(\reg_yHat[11][15] ), .B(n41413), .X(n37383) );
  nand_x1_sg U72756 ( .A(\yHat[11][16] ), .B(n40790), .X(n37384) );
  nand_x1_sg U72757 ( .A(\reg_yHat[11][16] ), .B(n40600), .X(n37385) );
  nand_x1_sg U72758 ( .A(\y[2][7] ), .B(n40762), .X(n37606) );
  nand_x1_sg U72759 ( .A(\reg_y[2][7] ), .B(n40437), .X(n37607) );
  nand_x1_sg U72760 ( .A(\y[2][8] ), .B(n40820), .X(n37608) );
  nand_x1_sg U72761 ( .A(\reg_y[2][8] ), .B(n40380), .X(n37609) );
  nand_x1_sg U72762 ( .A(\y[2][9] ), .B(n40760), .X(n37610) );
  nand_x1_sg U72763 ( .A(\reg_y[2][9] ), .B(n40415), .X(n37611) );
  nand_x1_sg U72764 ( .A(\y[2][10] ), .B(n39417), .X(n37612) );
  nand_x1_sg U72765 ( .A(\reg_y[2][10] ), .B(n39650), .X(n37613) );
  nand_x1_sg U72766 ( .A(\y[2][11] ), .B(n39406), .X(n37614) );
  nand_x1_sg U72767 ( .A(\reg_y[2][11] ), .B(n41434), .X(n37615) );
  nand_x1_sg U72768 ( .A(\y[2][12] ), .B(n40831), .X(n37616) );
  nand_x1_sg U72769 ( .A(\reg_y[2][12] ), .B(n40425), .X(n37617) );
  nand_x1_sg U72770 ( .A(\y[2][13] ), .B(n40792), .X(n37618) );
  nand_x1_sg U72771 ( .A(\reg_y[2][13] ), .B(n39432), .X(n37619) );
  nand_x1_sg U72772 ( .A(\y[2][14] ), .B(n41490), .X(n37620) );
  nand_x1_sg U72773 ( .A(\reg_y[2][14] ), .B(n39163), .X(n37621) );
  nand_x1_sg U72774 ( .A(\y[2][15] ), .B(n40823), .X(n37622) );
  nand_x1_sg U72775 ( .A(\reg_y[2][15] ), .B(n40605), .X(n37623) );
  nand_x1_sg U72776 ( .A(\y[2][16] ), .B(n40835), .X(n37624) );
  nand_x1_sg U72777 ( .A(\reg_y[2][16] ), .B(n40410), .X(n37625) );
  nand_x1_sg U72778 ( .A(\y[3][1] ), .B(n41517), .X(n37634) );
  nand_x1_sg U72779 ( .A(\reg_y[3][1] ), .B(n40010), .X(n37635) );
  nand_x1_sg U72780 ( .A(\y[3][2] ), .B(n39425), .X(n37636) );
  nand_x1_sg U72781 ( .A(\reg_y[3][2] ), .B(n40011), .X(n37637) );
  nand_x1_sg U72782 ( .A(\y[3][7] ), .B(n39419), .X(n37646) );
  nand_x1_sg U72783 ( .A(\reg_y[3][7] ), .B(n40413), .X(n37647) );
  nand_x1_sg U72784 ( .A(\y[3][8] ), .B(n41044), .X(n37648) );
  nand_x1_sg U72785 ( .A(\reg_y[3][8] ), .B(n40452), .X(n37649) );
  nand_x1_sg U72786 ( .A(\y[5][1] ), .B(n40777), .X(n37714) );
  nand_x1_sg U72787 ( .A(\reg_y[5][1] ), .B(n40451), .X(n37715) );
  nand_x1_sg U72788 ( .A(\y[5][2] ), .B(n40822), .X(n37716) );
  nand_x1_sg U72789 ( .A(\reg_y[5][2] ), .B(n40598), .X(n37717) );
  nand_x1_sg U72790 ( .A(\y[5][7] ), .B(n40807), .X(n37726) );
  nand_x1_sg U72791 ( .A(\reg_y[5][7] ), .B(n40399), .X(n37727) );
  nand_x1_sg U72792 ( .A(\y[5][8] ), .B(n41493), .X(n37728) );
  nand_x1_sg U72793 ( .A(\reg_y[5][8] ), .B(n41448), .X(n37729) );
  nand_x1_sg U72794 ( .A(\y[5][9] ), .B(n40806), .X(n37730) );
  nand_x1_sg U72795 ( .A(\reg_y[5][9] ), .B(n41424), .X(n37731) );
  nand_x1_sg U72796 ( .A(\y[5][10] ), .B(n40830), .X(n37732) );
  nand_x1_sg U72797 ( .A(\reg_y[5][10] ), .B(n40451), .X(n37733) );
  nand_x1_sg U72798 ( .A(\y[5][11] ), .B(n40758), .X(n37734) );
  nand_x1_sg U72799 ( .A(\reg_y[5][11] ), .B(n40397), .X(n37735) );
  nand_x1_sg U72800 ( .A(\y[5][12] ), .B(n38911), .X(n37736) );
  nand_x1_sg U72801 ( .A(\reg_y[5][12] ), .B(n40590), .X(n37737) );
  nand_x1_sg U72802 ( .A(\y[5][13] ), .B(n40794), .X(n37738) );
  nand_x1_sg U72803 ( .A(\reg_y[5][13] ), .B(n39158), .X(n37739) );
  nand_x1_sg U72804 ( .A(\y[5][14] ), .B(n40795), .X(n37740) );
  nand_x1_sg U72805 ( .A(\reg_y[5][14] ), .B(n40446), .X(n37741) );
  nand_x1_sg U72806 ( .A(\y[5][15] ), .B(n40772), .X(n37742) );
  nand_x1_sg U72807 ( .A(\reg_y[5][15] ), .B(n39183), .X(n37743) );
  nand_x1_sg U72808 ( .A(\y[5][16] ), .B(n40763), .X(n37744) );
  nand_x1_sg U72809 ( .A(\reg_y[5][16] ), .B(n39177), .X(n37745) );
  nand_x1_sg U72810 ( .A(\y[8][14] ), .B(n39272), .X(n37860) );
  nand_x1_sg U72811 ( .A(\reg_y[8][14] ), .B(n40449), .X(n37861) );
  nand_x1_sg U72812 ( .A(\y[8][15] ), .B(n39426), .X(n37862) );
  nand_x1_sg U72813 ( .A(\reg_y[8][15] ), .B(n40384), .X(n37863) );
  nand_x1_sg U72814 ( .A(\y[8][16] ), .B(n40773), .X(n37864) );
  nand_x1_sg U72815 ( .A(\reg_y[8][16] ), .B(n40395), .X(n37865) );
  nand_x1_sg U72816 ( .A(\y[9][1] ), .B(n39285), .X(n37874) );
  nand_x1_sg U72817 ( .A(\reg_y[9][1] ), .B(n41444), .X(n37875) );
  nand_x1_sg U72818 ( .A(\y[9][2] ), .B(n40818), .X(n37876) );
  nand_x1_sg U72819 ( .A(\reg_y[9][2] ), .B(n39162), .X(n37877) );
  nand_x1_sg U72820 ( .A(\y[9][7] ), .B(n40820), .X(n37886) );
  nand_x1_sg U72821 ( .A(\reg_y[9][7] ), .B(n39177), .X(n37887) );
  nand_x1_sg U72822 ( .A(\y[9][8] ), .B(n41510), .X(n37888) );
  nand_x1_sg U72823 ( .A(\reg_y[9][8] ), .B(n39173), .X(n37889) );
  nand_x1_sg U72824 ( .A(\y[9][9] ), .B(n39421), .X(n37890) );
  nand_x1_sg U72825 ( .A(\reg_y[9][9] ), .B(n41443), .X(n37891) );
  nand_x1_sg U72826 ( .A(\y[9][10] ), .B(n40808), .X(n37892) );
  nand_x1_sg U72827 ( .A(\reg_y[9][10] ), .B(n41414), .X(n37893) );
  nand_x1_sg U72828 ( .A(\y[9][11] ), .B(n40787), .X(n37894) );
  nand_x1_sg U72829 ( .A(\reg_y[9][11] ), .B(n40394), .X(n37895) );
  nand_x1_sg U72830 ( .A(\y[9][12] ), .B(n41501), .X(n37896) );
  nand_x1_sg U72831 ( .A(\reg_y[9][12] ), .B(n39183), .X(n37897) );
  nand_x1_sg U72832 ( .A(\y[9][13] ), .B(n40796), .X(n37898) );
  nand_x1_sg U72833 ( .A(\reg_y[9][13] ), .B(n40396), .X(n37899) );
  nand_x1_sg U72834 ( .A(\y[9][14] ), .B(n41514), .X(n37900) );
  nand_x1_sg U72835 ( .A(\reg_y[9][14] ), .B(n39197), .X(n37901) );
  nand_x1_sg U72836 ( .A(\y[9][15] ), .B(n40804), .X(n37902) );
  nand_x1_sg U72837 ( .A(\reg_y[9][15] ), .B(n41428), .X(n37903) );
  nand_x1_sg U72838 ( .A(\y[9][16] ), .B(n41046), .X(n37904) );
  nand_x1_sg U72839 ( .A(\reg_y[9][16] ), .B(n40429), .X(n37905) );
  nand_x1_sg U72840 ( .A(\y[10][1] ), .B(n39416), .X(n37914) );
  nand_x1_sg U72841 ( .A(\reg_y[10][1] ), .B(n40444), .X(n37915) );
  nand_x1_sg U72842 ( .A(\y[10][2] ), .B(n40765), .X(n37916) );
  nand_x1_sg U72843 ( .A(\reg_y[10][2] ), .B(n41428), .X(n37917) );
  nand_x1_sg U72844 ( .A(\y[2][4] ), .B(n41046), .X(n37600) );
  nand_x1_sg U72845 ( .A(\reg_y[2][4] ), .B(n41440), .X(n37601) );
  nand_x1_sg U72846 ( .A(\y[3][4] ), .B(n40819), .X(n37640) );
  nand_x1_sg U72847 ( .A(\reg_y[3][4] ), .B(n41475), .X(n37641) );
  nand_x1_sg U72848 ( .A(\y[5][4] ), .B(n40780), .X(n37720) );
  nand_x1_sg U72849 ( .A(\reg_y[5][4] ), .B(n40411), .X(n37721) );
  nand_x1_sg U72850 ( .A(\y[9][4] ), .B(n41499), .X(n37880) );
  nand_x1_sg U72851 ( .A(\reg_y[9][4] ), .B(n41476), .X(n37881) );
  nand_x1_sg U72852 ( .A(\yHat[3][18] ), .B(n39270), .X(n37068) );
  nand_x1_sg U72853 ( .A(\reg_yHat[3][18] ), .B(n39163), .X(n37069) );
  nand_x1_sg U72854 ( .A(\yHat[10][18] ), .B(n41498), .X(n37348) );
  nand_x1_sg U72855 ( .A(\reg_yHat[10][18] ), .B(n40441), .X(n37349) );
  nand_x1_sg U72856 ( .A(\yHat[11][18] ), .B(n38851), .X(n37388) );
  nand_x1_sg U72857 ( .A(\reg_yHat[11][18] ), .B(n40382), .X(n37389) );
  nand_x1_sg U72858 ( .A(\y[2][19] ), .B(n41494), .X(n37630) );
  nand_x1_sg U72859 ( .A(\reg_y[2][19] ), .B(n39187), .X(n37631) );
  nand_x1_sg U72860 ( .A(\y[3][0] ), .B(n39271), .X(n37632) );
  nand_x1_sg U72861 ( .A(\reg_y[3][0] ), .B(n41426), .X(n37633) );
  nand_x1_sg U72862 ( .A(\y[4][19] ), .B(n40759), .X(n37710) );
  nand_x1_sg U72863 ( .A(\reg_y[4][19] ), .B(n39198), .X(n37711) );
  nand_x1_sg U72864 ( .A(\y[5][0] ), .B(n41499), .X(n37712) );
  nand_x1_sg U72865 ( .A(\reg_y[5][0] ), .B(n40421), .X(n37713) );
  nand_x1_sg U72866 ( .A(\y[8][19] ), .B(n40828), .X(n37870) );
  nand_x1_sg U72867 ( .A(\reg_y[8][19] ), .B(n40599), .X(n37871) );
  nand_x1_sg U72868 ( .A(\y[9][0] ), .B(n38849), .X(n37872) );
  nand_x1_sg U72869 ( .A(\reg_y[9][0] ), .B(n39173), .X(n37873) );
  nand_x1_sg U72870 ( .A(\y[9][19] ), .B(n38843), .X(n37910) );
  nand_x1_sg U72871 ( .A(\reg_y[9][19] ), .B(n40430), .X(n37911) );
  nand_x1_sg U72872 ( .A(\y[10][0] ), .B(n40819), .X(n37912) );
  nand_x1_sg U72873 ( .A(\reg_y[10][0] ), .B(n39177), .X(n37913) );
  nand_x1_sg U72874 ( .A(\yHat[3][1] ), .B(n39272), .X(n37034) );
  nand_x1_sg U72875 ( .A(\reg_yHat[3][1] ), .B(n40390), .X(n37035) );
  nand_x1_sg U72876 ( .A(\yHat[11][1] ), .B(n39414), .X(n37354) );
  nand_x1_sg U72877 ( .A(\reg_yHat[11][1] ), .B(n40594), .X(n37355) );
  nand_x1_sg U72878 ( .A(\y[2][5] ), .B(n38834), .X(n37602) );
  nand_x1_sg U72879 ( .A(\reg_y[2][5] ), .B(n41445), .X(n37603) );
  nand_x1_sg U72880 ( .A(\y[2][18] ), .B(n40750), .X(n37628) );
  nand_x1_sg U72881 ( .A(\reg_y[2][18] ), .B(n39650), .X(n37629) );
  nand_x1_sg U72882 ( .A(\y[3][5] ), .B(n39426), .X(n37642) );
  nand_x1_sg U72883 ( .A(\reg_y[3][5] ), .B(n40430), .X(n37643) );
  nand_x1_sg U72884 ( .A(\y[5][5] ), .B(n40778), .X(n37722) );
  nand_x1_sg U72885 ( .A(\reg_y[5][5] ), .B(n39178), .X(n37723) );
  nand_x1_sg U72886 ( .A(\y[5][18] ), .B(n38859), .X(n37748) );
  nand_x1_sg U72887 ( .A(\reg_y[5][18] ), .B(n40591), .X(n37749) );
  nand_x1_sg U72888 ( .A(\y[8][18] ), .B(n41510), .X(n37868) );
  nand_x1_sg U72889 ( .A(\reg_y[8][18] ), .B(n40439), .X(n37869) );
  nand_x1_sg U72890 ( .A(\y[9][5] ), .B(n40751), .X(n37882) );
  nand_x1_sg U72891 ( .A(\reg_y[9][5] ), .B(n40425), .X(n37883) );
  nand_x1_sg U72892 ( .A(\y[9][18] ), .B(n38860), .X(n37908) );
  nand_x1_sg U72893 ( .A(\reg_y[9][18] ), .B(n39483), .X(n37909) );
  nand_x1_sg U72894 ( .A(\yHat[3][6] ), .B(n41517), .X(n37044) );
  nand_x1_sg U72895 ( .A(\reg_yHat[3][6] ), .B(n40421), .X(n37045) );
  nand_x1_sg U72896 ( .A(\yHat[5][6] ), .B(n39420), .X(n37124) );
  nand_x1_sg U72897 ( .A(\reg_yHat[5][6] ), .B(n40599), .X(n37125) );
  nand_x1_sg U72898 ( .A(\yHat[11][6] ), .B(n41508), .X(n37364) );
  nand_x1_sg U72899 ( .A(\reg_yHat[11][6] ), .B(n41480), .X(n37365) );
  inv_x1_sg U72900 ( .A(state[0]), .X(n51530) );
  nand_x1_sg U72901 ( .A(output_taken), .B(n51530), .X(n29275) );
  nor_x1_sg U72902 ( .A(state[1]), .B(state[0]), .X(n38120) );
  nor_x1_sg U72903 ( .A(n36903), .B(n39728), .X(n1999) );
  nor_x1_sg U72904 ( .A(state[1]), .B(n36904), .X(n36903) );
  nor_x1_sg U72905 ( .A(n36908), .B(n51530), .X(n36904) );
  nand_x1_sg U72906 ( .A(n42022), .B(done), .X(n36908) );
  nand_x1_sg U72907 ( .A(out_L2[2]), .B(n39267), .X(n36876) );
  nand_x1_sg U72908 ( .A(out_L1[2]), .B(n41267), .X(n36877) );
  nand_x1_sg U72909 ( .A(out_L2[9]), .B(n41054), .X(n36862) );
  nand_x1_sg U72910 ( .A(n41269), .B(out_L1[9]), .X(n36863) );
  nand_x1_sg U72911 ( .A(out_L2[0]), .B(n39267), .X(n36900) );
  nand_x1_sg U72912 ( .A(out_L1[0]), .B(n41269), .X(n36901) );
  nand_x1_sg U72913 ( .A(out_L2[10]), .B(n41053), .X(n36898) );
  nand_x1_sg U72914 ( .A(out_L1[10]), .B(n41270), .X(n36899) );
  nand_x1_sg U72915 ( .A(out_L2[11]), .B(n41054), .X(n36896) );
  nand_x1_sg U72916 ( .A(out_L1[11]), .B(n41268), .X(n36897) );
  nand_x1_sg U72917 ( .A(out_L2[12]), .B(n41054), .X(n36894) );
  nand_x1_sg U72918 ( .A(out_L1[12]), .B(n41269), .X(n36895) );
  nand_x1_sg U72919 ( .A(out_L2[13]), .B(n41053), .X(n36892) );
  nand_x1_sg U72920 ( .A(out_L1[13]), .B(n41273), .X(n36893) );
  nand_x1_sg U72921 ( .A(out_L2[14]), .B(n41053), .X(n36890) );
  nand_x1_sg U72922 ( .A(out_L1[14]), .B(n41274), .X(n36891) );
  nand_x1_sg U72923 ( .A(out_L2[15]), .B(n41055), .X(n36888) );
  nand_x1_sg U72924 ( .A(out_L1[15]), .B(n41271), .X(n36889) );
  nand_x1_sg U72925 ( .A(out_L2[17]), .B(n41052), .X(n36884) );
  nand_x1_sg U72926 ( .A(out_L1[17]), .B(n41269), .X(n36885) );
  nand_x1_sg U72927 ( .A(out_L2[18]), .B(n41055), .X(n36882) );
  nand_x1_sg U72928 ( .A(out_L1[18]), .B(n41270), .X(n36883) );
  nand_x1_sg U72929 ( .A(out_L2[19]), .B(n39267), .X(n36880) );
  nand_x1_sg U72930 ( .A(out_L1[19]), .B(n41274), .X(n36881) );
  nand_x1_sg U72931 ( .A(out_L2[3]), .B(n39267), .X(n36874) );
  nand_x1_sg U72932 ( .A(out_L1[3]), .B(n41268), .X(n36875) );
  nand_x1_sg U72933 ( .A(out_L2[4]), .B(n41052), .X(n36872) );
  nand_x1_sg U72934 ( .A(out_L1[4]), .B(n41271), .X(n36873) );
  nand_x1_sg U72935 ( .A(out_L2[5]), .B(n41052), .X(n36870) );
  nand_x1_sg U72936 ( .A(out_L1[5]), .B(n41270), .X(n36871) );
  nand_x1_sg U72937 ( .A(out_L2[6]), .B(n41055), .X(n36868) );
  nand_x1_sg U72938 ( .A(out_L1[6]), .B(n41272), .X(n36869) );
  nand_x1_sg U72939 ( .A(out_L2[7]), .B(n41055), .X(n36866) );
  nand_x1_sg U72940 ( .A(out_L1[7]), .B(n41272), .X(n36867) );
  nand_x1_sg U72941 ( .A(out_L2[8]), .B(n41945), .X(n36864) );
  nand_x1_sg U72942 ( .A(out_L1[8]), .B(n41273), .X(n36865) );
  nand_x1_sg U72943 ( .A(out_L2[1]), .B(n41054), .X(n36878) );
  nand_x1_sg U72944 ( .A(out_L2[16]), .B(n41053), .X(n36886) );
  nand_x1_sg U72945 ( .A(n39288), .B(n26772), .X(n24937) );
  nand_x1_sg U72946 ( .A(n26767), .B(n42021), .X(n26772) );
  nand_x1_sg U72947 ( .A(n39288), .B(n26779), .X(n25216) );
  nand_x1_sg U72948 ( .A(n41660), .B(n42021), .X(n26779) );
  nor_x1_sg U72949 ( .A(reg_num[2]), .B(reg_num[3]), .X(n23543) );
  nor_x1_sg U72950 ( .A(reg_num[0]), .B(n39486), .X(n26767) );
  nor_x1_sg U72951 ( .A(n39139), .B(n26331), .X(n26184) );
  nor_x1_sg U72952 ( .A(n39727), .B(reg_num[1]), .X(n26331) );
  nor_x1_sg U72953 ( .A(n38133), .B(n42159), .X(n27969) );
  nor_x1_sg U72954 ( .A(n27970), .B(n5726), .X(n27968) );
  nor_x1_sg U72955 ( .A(n41524), .B(n5720), .X(n28809) );
  nor_x1_sg U72956 ( .A(n38134), .B(n22595), .X(n28810) );
  nor_x1_sg U72957 ( .A(n6071), .B(n46474), .X(n19948) );
  nor_x1_sg U72958 ( .A(n19951), .B(n41552), .X(n19950) );
  nor_x1_sg U72959 ( .A(n46573), .B(n5438), .X(n19341) );
  nor_x1_sg U72960 ( .A(n6038), .B(n19328), .X(n19340) );
  nor_x1_sg U72961 ( .A(n46388), .B(n5442), .X(n19354) );
  nor_x1_sg U72962 ( .A(n6226), .B(n46343), .X(n19353) );
  nor_x1_sg U72963 ( .A(n42295), .B(n21170), .X(n21204) );
  nor_x1_sg U72964 ( .A(n46537), .B(n46549), .X(n21206) );
  nor_x1_sg U72965 ( .A(n38135), .B(n45801), .X(n20842) );
  nor_x1_sg U72966 ( .A(n6821), .B(n5707), .X(n20841) );
  nor_x1_sg U72967 ( .A(n38136), .B(n45803), .X(n20489) );
  nor_x1_sg U72968 ( .A(n6818), .B(n5709), .X(n20488) );
  nor_x1_sg U72969 ( .A(n38137), .B(n45805), .X(n20199) );
  nor_x1_sg U72970 ( .A(n6797), .B(n5711), .X(n20198) );
  nor_x1_sg U72971 ( .A(n38138), .B(n45807), .X(n19832) );
  nor_x1_sg U72972 ( .A(n6794), .B(n5713), .X(n19831) );
  nor_x1_sg U72973 ( .A(n38139), .B(n45809), .X(n19393) );
  nor_x1_sg U72974 ( .A(n6807), .B(n5715), .X(n19392) );
  nor_x1_sg U72975 ( .A(n26113), .B(n42015), .X(n26168) );
  nor_x1_sg U72976 ( .A(n26170), .B(\reg_y[12][3] ), .X(n26169) );
  nor_x1_sg U72977 ( .A(\reg_yHat[12][3] ), .B(n50279), .X(n26170) );
  nor_x1_sg U72978 ( .A(n41971), .B(n46528), .X(n19571) );
  nor_x1_sg U72979 ( .A(n19507), .B(n19504), .X(n19573) );
  nor_x1_sg U72980 ( .A(n38140), .B(n21258), .X(n21257) );
  nor_x1_sg U72981 ( .A(n45799), .B(n5705), .X(n21256) );
  nor_x1_sg U72982 ( .A(n42215), .B(n46843), .X(n22832) );
  nor_x1_sg U72983 ( .A(n22834), .B(\reg_yHat[0][2] ), .X(n22831) );
  inv_x1_sg U72984 ( .A(n22833), .X(n46843) );
  nor_x1_sg U72985 ( .A(n23111), .B(\reg_yHat[1][2] ), .X(n23108) );
  nand_x1_sg U72986 ( .A(\reg_y[1][2] ), .B(n23110), .X(n23109) );
  nor_x1_sg U72987 ( .A(n23391), .B(\reg_yHat[2][2] ), .X(n23388) );
  nand_x1_sg U72988 ( .A(\reg_y[2][2] ), .B(n23390), .X(n23389) );
  nor_x1_sg U72989 ( .A(n23670), .B(\reg_yHat[3][2] ), .X(n23667) );
  nand_x1_sg U72990 ( .A(\reg_y[3][2] ), .B(n23669), .X(n23668) );
  nor_x1_sg U72991 ( .A(n23949), .B(\reg_yHat[4][2] ), .X(n23946) );
  nand_x1_sg U72992 ( .A(\reg_y[4][2] ), .B(n23948), .X(n23947) );
  nor_x1_sg U72993 ( .A(n24228), .B(\reg_yHat[5][2] ), .X(n24225) );
  nand_x1_sg U72994 ( .A(\reg_y[5][2] ), .B(n24227), .X(n24226) );
  nor_x1_sg U72995 ( .A(n24507), .B(\reg_yHat[6][2] ), .X(n24504) );
  nand_x1_sg U72996 ( .A(\reg_y[6][2] ), .B(n24506), .X(n24505) );
  nor_x1_sg U72997 ( .A(n24785), .B(\reg_yHat[7][2] ), .X(n24782) );
  nand_x1_sg U72998 ( .A(\reg_y[7][2] ), .B(n24784), .X(n24783) );
  nor_x1_sg U72999 ( .A(n25064), .B(\reg_yHat[8][2] ), .X(n25061) );
  nand_x1_sg U73000 ( .A(\reg_y[8][2] ), .B(n25063), .X(n25062) );
  nor_x1_sg U73001 ( .A(n25343), .B(\reg_yHat[9][2] ), .X(n25340) );
  nand_x1_sg U73002 ( .A(\reg_y[9][2] ), .B(n25342), .X(n25341) );
  nor_x1_sg U73003 ( .A(n25622), .B(\reg_yHat[10][2] ), .X(n25619) );
  nand_x1_sg U73004 ( .A(\reg_y[10][2] ), .B(n25621), .X(n25620) );
  nor_x1_sg U73005 ( .A(n25899), .B(\reg_yHat[11][2] ), .X(n25896) );
  nand_x1_sg U73006 ( .A(\reg_y[11][2] ), .B(n25898), .X(n25897) );
  nor_x1_sg U73007 ( .A(n26459), .B(\reg_yHat[13][2] ), .X(n26456) );
  nand_x1_sg U73008 ( .A(\reg_y[13][2] ), .B(n26458), .X(n26457) );
  nor_x1_sg U73009 ( .A(n26737), .B(\reg_yHat[14][2] ), .X(n26734) );
  nand_x1_sg U73010 ( .A(\reg_y[14][2] ), .B(n26736), .X(n26735) );
  nand_x1_sg U73011 ( .A(\reg_yHat[1][0] ), .B(n47133), .X(n23123) );
  nand_x1_sg U73012 ( .A(\reg_yHat[2][0] ), .B(n47419), .X(n23403) );
  nand_x1_sg U73013 ( .A(\reg_yHat[3][0] ), .B(n47704), .X(n23682) );
  nand_x1_sg U73014 ( .A(\reg_yHat[4][0] ), .B(n47989), .X(n23961) );
  nand_x1_sg U73015 ( .A(\reg_yHat[5][0] ), .B(n48274), .X(n24240) );
  nand_x1_sg U73016 ( .A(\reg_yHat[6][0] ), .B(n48559), .X(n24519) );
  nand_x1_sg U73017 ( .A(\reg_yHat[7][0] ), .B(n48844), .X(n24797) );
  nand_x1_sg U73018 ( .A(\reg_yHat[8][0] ), .B(n49131), .X(n25076) );
  nand_x1_sg U73019 ( .A(\reg_yHat[9][0] ), .B(n49417), .X(n25355) );
  nand_x1_sg U73020 ( .A(\reg_yHat[10][0] ), .B(n49703), .X(n25634) );
  nand_x1_sg U73021 ( .A(\reg_yHat[11][0] ), .B(n49989), .X(n25911) );
  nand_x1_sg U73022 ( .A(\reg_yHat[13][0] ), .B(n50562), .X(n26471) );
  nand_x1_sg U73023 ( .A(\reg_yHat[14][0] ), .B(n50849), .X(n26749) );
  nor_x1_sg U73024 ( .A(n42302), .B(n21249), .X(n21246) );
  nor_x1_sg U73025 ( .A(n45911), .B(n45922), .X(n21248) );
  nor_x1_sg U73026 ( .A(n42298), .B(n20481), .X(n20478) );
  nor_x1_sg U73027 ( .A(n45901), .B(n45925), .X(n20480) );
  nor_x1_sg U73028 ( .A(n42285), .B(n19824), .X(n19821) );
  nor_x1_sg U73029 ( .A(n45891), .B(n45928), .X(n19823) );
  nor_x1_sg U73030 ( .A(n6119), .B(n20155), .X(n20152) );
  nor_x1_sg U73031 ( .A(n46447), .B(n46476), .X(n20154) );
  nor_x1_sg U73032 ( .A(n6068), .B(n19963), .X(n19960) );
  nor_x1_sg U73033 ( .A(n46486), .B(n46518), .X(n19962) );
  nor_x1_sg U73034 ( .A(n41537), .B(n20316), .X(n20313) );
  nor_x1_sg U73035 ( .A(n46400), .B(n20288), .X(n20315) );
  nand_x1_sg U73036 ( .A(n28133), .B(n28135), .X(n28250) );
  nand_x1_sg U73037 ( .A(n20498), .B(n20501), .X(n20654) );
  nand_x1_sg U73038 ( .A(n19841), .B(n19844), .X(n20014) );
  nand_x1_sg U73039 ( .A(n6712), .B(n6715), .X(n19210) );
  nand_x1_sg U73040 ( .A(n21267), .B(n21270), .X(n21424) );
  nand_x1_sg U73041 ( .A(\reg_yHat[12][0] ), .B(n50275), .X(n26128) );
  nand_x1_sg U73042 ( .A(\reg_yHat[0][0] ), .B(n46841), .X(n22851) );
  nand_x1_sg U73043 ( .A(n41419), .B(n39288), .X(n13370) );
  nor_x1_sg U73044 ( .A(n42294), .B(n19976), .X(n19973) );
  nor_x1_sg U73045 ( .A(n46304), .B(n46337), .X(n19975) );
  nor_x1_sg U73046 ( .A(n38141), .B(n45802), .X(n20659) );
  nor_x1_sg U73047 ( .A(n20660), .B(n5708), .X(n20658) );
  nor_x1_sg U73048 ( .A(n38142), .B(n45804), .X(n20358) );
  nor_x1_sg U73049 ( .A(n20359), .B(n5710), .X(n20357) );
  nor_x1_sg U73050 ( .A(n38143), .B(n45806), .X(n20019) );
  nor_x1_sg U73051 ( .A(n20020), .B(n5712), .X(n20018) );
  nor_x1_sg U73052 ( .A(n38144), .B(n45808), .X(n19625) );
  nor_x1_sg U73053 ( .A(n19626), .B(n5714), .X(n19624) );
  nor_x1_sg U73054 ( .A(n38145), .B(n45800), .X(n21067) );
  nor_x1_sg U73055 ( .A(n21068), .B(n5706), .X(n21066) );
  nand_x1_sg U73056 ( .A(n46508), .B(n19944), .X(n19945) );
  nor_x1_sg U73057 ( .A(n6211), .B(n46349), .X(n20159) );
  nor_x1_sg U73058 ( .A(n20108), .B(n41551), .X(n20161) );
  nor_x1_sg U73059 ( .A(n46525), .B(n5439), .X(n19344) );
  nor_x1_sg U73060 ( .A(n42341), .B(n19322), .X(n19343) );
  nor_x1_sg U73061 ( .A(n6134), .B(n19349), .X(n19346) );
  nor_x1_sg U73062 ( .A(n46437), .B(n46479), .X(n19348) );
  nor_x1_sg U73063 ( .A(n38146), .B(n45810), .X(n19215) );
  nor_x1_sg U73064 ( .A(n19216), .B(n5716), .X(n19214) );
  nor_x1_sg U73065 ( .A(n42262), .B(n19786), .X(n19783) );
  nor_x1_sg U73066 ( .A(n46442), .B(n19712), .X(n19785) );
  nor_x1_sg U73067 ( .A(n23084), .B(n46648), .X(n23081) );
  nor_x1_sg U73068 ( .A(n23083), .B(\reg_y[1][5] ), .X(n23082) );
  nor_x1_sg U73069 ( .A(\reg_yHat[1][5] ), .B(n42145), .X(n23083) );
  nor_x1_sg U73070 ( .A(n23364), .B(n46662), .X(n23361) );
  nor_x1_sg U73071 ( .A(n23363), .B(\reg_y[2][5] ), .X(n23362) );
  nor_x1_sg U73072 ( .A(\reg_yHat[2][5] ), .B(n42144), .X(n23363) );
  nor_x1_sg U73073 ( .A(n23643), .B(n46676), .X(n23640) );
  nor_x1_sg U73074 ( .A(n23642), .B(\reg_y[3][5] ), .X(n23641) );
  nor_x1_sg U73075 ( .A(\reg_yHat[3][5] ), .B(n42143), .X(n23642) );
  nor_x1_sg U73076 ( .A(n23922), .B(n46690), .X(n23919) );
  nor_x1_sg U73077 ( .A(n23921), .B(\reg_y[4][5] ), .X(n23920) );
  nor_x1_sg U73078 ( .A(\reg_yHat[4][5] ), .B(n42142), .X(n23921) );
  nor_x1_sg U73079 ( .A(n24201), .B(n46704), .X(n24198) );
  nor_x1_sg U73080 ( .A(n24200), .B(\reg_y[5][5] ), .X(n24199) );
  nor_x1_sg U73081 ( .A(\reg_yHat[5][5] ), .B(n42141), .X(n24200) );
  nor_x1_sg U73082 ( .A(n24480), .B(n46718), .X(n24477) );
  nor_x1_sg U73083 ( .A(n24479), .B(\reg_y[6][5] ), .X(n24478) );
  nor_x1_sg U73084 ( .A(\reg_yHat[6][5] ), .B(n42140), .X(n24479) );
  nor_x1_sg U73085 ( .A(n24758), .B(n46732), .X(n24755) );
  nor_x1_sg U73086 ( .A(n24757), .B(\reg_y[7][5] ), .X(n24756) );
  nor_x1_sg U73087 ( .A(\reg_yHat[7][5] ), .B(n42139), .X(n24757) );
  nor_x1_sg U73088 ( .A(n25037), .B(n46746), .X(n25034) );
  nor_x1_sg U73089 ( .A(n25036), .B(\reg_y[8][5] ), .X(n25035) );
  nor_x1_sg U73090 ( .A(\reg_yHat[8][5] ), .B(n42138), .X(n25036) );
  nor_x1_sg U73091 ( .A(n25316), .B(n46760), .X(n25313) );
  nor_x1_sg U73092 ( .A(n25315), .B(\reg_y[9][5] ), .X(n25314) );
  nor_x1_sg U73093 ( .A(\reg_yHat[9][5] ), .B(n42137), .X(n25315) );
  nor_x1_sg U73094 ( .A(n25595), .B(n46774), .X(n25592) );
  nor_x1_sg U73095 ( .A(n25594), .B(\reg_y[10][5] ), .X(n25593) );
  nor_x1_sg U73096 ( .A(\reg_yHat[10][5] ), .B(n42060), .X(n25594) );
  nor_x1_sg U73097 ( .A(n25872), .B(n46788), .X(n25869) );
  nor_x1_sg U73098 ( .A(n25871), .B(\reg_y[11][5] ), .X(n25870) );
  nor_x1_sg U73099 ( .A(\reg_yHat[11][5] ), .B(n42136), .X(n25871) );
  nor_x1_sg U73100 ( .A(n26432), .B(n46815), .X(n26429) );
  nor_x1_sg U73101 ( .A(n26431), .B(\reg_y[13][5] ), .X(n26430) );
  nor_x1_sg U73102 ( .A(\reg_yHat[13][5] ), .B(n42135), .X(n26431) );
  nor_x1_sg U73103 ( .A(n26710), .B(n46829), .X(n26707) );
  nor_x1_sg U73104 ( .A(n26709), .B(\reg_y[14][5] ), .X(n26708) );
  nor_x1_sg U73105 ( .A(\reg_yHat[14][5] ), .B(n42134), .X(n26709) );
  nor_x1_sg U73106 ( .A(n46635), .B(n22807), .X(n22804) );
  nor_x1_sg U73107 ( .A(n22806), .B(\reg_y[0][5] ), .X(n22805) );
  nor_x1_sg U73108 ( .A(\reg_yHat[0][5] ), .B(n42146), .X(n22806) );
  nor_x1_sg U73109 ( .A(n6024), .B(n46516), .X(n19764) );
  nor_x1_sg U73110 ( .A(n19767), .B(n41550), .X(n19766) );
  nor_x1_sg U73111 ( .A(n6169), .B(n46386), .X(n19163) );
  nor_x1_sg U73112 ( .A(n6175), .B(n41553), .X(n19165) );
  nor_x1_sg U73113 ( .A(n46579), .B(n5609), .X(n21015) );
  nor_x1_sg U73114 ( .A(n6055), .B(n46535), .X(n21014) );
  nor_x1_sg U73115 ( .A(n42283), .B(n19755), .X(n19752) );
  nor_x1_sg U73116 ( .A(n46510), .B(n46557), .X(n19754) );
  nor_x1_sg U73117 ( .A(n42282), .B(n19172), .X(n19169) );
  nor_x1_sg U73118 ( .A(n46295), .B(n46340), .X(n19171) );
  nor_x1_sg U73119 ( .A(n6691), .B(n21059), .X(n21056) );
  nor_x1_sg U73120 ( .A(n45908), .B(n45923), .X(n21058) );
  nor_x1_sg U73121 ( .A(n6659), .B(n20350), .X(n20347) );
  nor_x1_sg U73122 ( .A(n45898), .B(n45926), .X(n20349) );
  nor_x1_sg U73123 ( .A(n6674), .B(n19617), .X(n19614) );
  nor_x1_sg U73124 ( .A(n45888), .B(n45929), .X(n19616) );
  nor_x1_sg U73125 ( .A(n6147), .B(n20604), .X(n20601) );
  nor_x1_sg U73126 ( .A(n46450), .B(n46470), .X(n20603) );
  nor_x1_sg U73127 ( .A(n41538), .B(n19903), .X(n19970) );
  nor_x1_sg U73128 ( .A(n46348), .B(n19899), .X(n19972) );
  nor_x1_sg U73129 ( .A(n6020), .B(n19779), .X(n19776) );
  nor_x1_sg U73130 ( .A(n46530), .B(n46567), .X(n19778) );
  nor_x1_sg U73131 ( .A(n42228), .B(n27106), .X(n27102) );
  nor_x1_sg U73132 ( .A(n45666), .B(n27105), .X(n27104) );
  nor_x1_sg U73133 ( .A(n41968), .B(n21201), .X(n21197) );
  nor_x1_sg U73134 ( .A(n46539), .B(n21200), .X(n21199) );
  nor_x1_sg U73135 ( .A(n46570), .B(n46523), .X(n19153) );
  nor_x1_sg U73136 ( .A(n6034), .B(n19156), .X(n19155) );
  nor_x1_sg U73137 ( .A(n41529), .B(n45830), .X(n20835) );
  inv_x1_sg U73138 ( .A(n20673), .X(n45830) );
  nor_x1_sg U73139 ( .A(n41528), .B(n45846), .X(n20192) );
  inv_x1_sg U73140 ( .A(n20033), .X(n45846) );
  nor_x1_sg U73141 ( .A(n41527), .B(n45862), .X(n19386) );
  inv_x1_sg U73142 ( .A(n19229), .X(n45862) );
  nor_x1_sg U73143 ( .A(n41533), .B(n46440), .X(n19577) );
  inv_x1_sg U73144 ( .A(n19494), .X(n46440) );
  nor_x1_sg U73145 ( .A(n22823), .B(\reg_y[0][3] ), .X(n22822) );
  nand_x1_sg U73146 ( .A(n38760), .B(n22824), .X(n22825) );
  nor_x1_sg U73147 ( .A(n47171), .B(n23076), .X(n23075) );
  nor_x1_sg U73148 ( .A(n47170), .B(\reg_yHat[1][6] ), .X(n23074) );
  nor_x1_sg U73149 ( .A(n42041), .B(n23077), .X(n23076) );
  nor_x1_sg U73150 ( .A(n47456), .B(n23356), .X(n23355) );
  nor_x1_sg U73151 ( .A(n47455), .B(\reg_yHat[2][6] ), .X(n23354) );
  nor_x1_sg U73152 ( .A(n42035), .B(n23357), .X(n23356) );
  nor_x1_sg U73153 ( .A(n47741), .B(n23635), .X(n23634) );
  nor_x1_sg U73154 ( .A(n47740), .B(\reg_yHat[3][6] ), .X(n23633) );
  nor_x1_sg U73155 ( .A(n42036), .B(n23636), .X(n23635) );
  nor_x1_sg U73156 ( .A(n48026), .B(n23914), .X(n23913) );
  nor_x1_sg U73157 ( .A(n48025), .B(\reg_yHat[4][6] ), .X(n23912) );
  nor_x1_sg U73158 ( .A(n42037), .B(n23915), .X(n23914) );
  nor_x1_sg U73159 ( .A(n48311), .B(n24193), .X(n24192) );
  nor_x1_sg U73160 ( .A(n48310), .B(\reg_yHat[5][6] ), .X(n24191) );
  nor_x1_sg U73161 ( .A(n42038), .B(n24194), .X(n24193) );
  nor_x1_sg U73162 ( .A(n48596), .B(n24472), .X(n24471) );
  nor_x1_sg U73163 ( .A(n48595), .B(\reg_yHat[6][6] ), .X(n24470) );
  nor_x1_sg U73164 ( .A(n42031), .B(n24473), .X(n24472) );
  nor_x1_sg U73165 ( .A(n48882), .B(n24750), .X(n24749) );
  nor_x1_sg U73166 ( .A(n48881), .B(\reg_yHat[7][6] ), .X(n24748) );
  nor_x1_sg U73167 ( .A(n42032), .B(n24751), .X(n24750) );
  nor_x1_sg U73168 ( .A(n49169), .B(n25029), .X(n25028) );
  nor_x1_sg U73169 ( .A(n49168), .B(\reg_yHat[8][6] ), .X(n25027) );
  nor_x1_sg U73170 ( .A(n42033), .B(n25030), .X(n25029) );
  nor_x1_sg U73171 ( .A(n49455), .B(n25308), .X(n25307) );
  nor_x1_sg U73172 ( .A(n49454), .B(\reg_yHat[9][6] ), .X(n25306) );
  nor_x1_sg U73173 ( .A(n42034), .B(n25309), .X(n25308) );
  nor_x1_sg U73174 ( .A(n49740), .B(n25587), .X(n25586) );
  nor_x1_sg U73175 ( .A(n49739), .B(\reg_yHat[10][6] ), .X(n25585) );
  nor_x1_sg U73176 ( .A(n42027), .B(n25588), .X(n25587) );
  nor_x1_sg U73177 ( .A(n50027), .B(n25864), .X(n25863) );
  nor_x1_sg U73178 ( .A(n50026), .B(\reg_yHat[11][6] ), .X(n25862) );
  nor_x1_sg U73179 ( .A(n42028), .B(n25865), .X(n25864) );
  nor_x1_sg U73180 ( .A(n50601), .B(n26424), .X(n26423) );
  nor_x1_sg U73181 ( .A(n50600), .B(\reg_yHat[13][6] ), .X(n26422) );
  nor_x1_sg U73182 ( .A(n42025), .B(n26425), .X(n26424) );
  nor_x1_sg U73183 ( .A(n50888), .B(n26702), .X(n26701) );
  nor_x1_sg U73184 ( .A(n50887), .B(\reg_yHat[14][6] ), .X(n26700) );
  nor_x1_sg U73185 ( .A(n42026), .B(n26703), .X(n26702) );
  nor_x1_sg U73186 ( .A(n46878), .B(n22799), .X(n22798) );
  nor_x1_sg U73187 ( .A(n46877), .B(\reg_yHat[0][6] ), .X(n22797) );
  nor_x1_sg U73188 ( .A(n42039), .B(n22800), .X(n22799) );
  nor_x1_sg U73189 ( .A(n50312), .B(n26161), .X(n26160) );
  nor_x1_sg U73190 ( .A(n50311), .B(\reg_yHat[12][6] ), .X(n26159) );
  nor_x1_sg U73191 ( .A(n42029), .B(n26096), .X(n26161) );
  inv_x1_sg U73192 ( .A(reg_num[0]), .X(n51136) );
  nor_x1_sg U73193 ( .A(n46841), .B(\reg_yHat[0][0] ), .X(n22843) );
  nor_x1_sg U73194 ( .A(n47133), .B(\reg_yHat[1][0] ), .X(n23120) );
  nor_x1_sg U73195 ( .A(n47419), .B(\reg_yHat[2][0] ), .X(n23400) );
  nor_x1_sg U73196 ( .A(n47704), .B(\reg_yHat[3][0] ), .X(n23679) );
  nor_x1_sg U73197 ( .A(n47989), .B(\reg_yHat[4][0] ), .X(n23958) );
  nor_x1_sg U73198 ( .A(n48274), .B(\reg_yHat[5][0] ), .X(n24237) );
  nor_x1_sg U73199 ( .A(n48559), .B(\reg_yHat[6][0] ), .X(n24516) );
  nor_x1_sg U73200 ( .A(n48844), .B(\reg_yHat[7][0] ), .X(n24794) );
  nor_x1_sg U73201 ( .A(n49131), .B(\reg_yHat[8][0] ), .X(n25073) );
  nor_x1_sg U73202 ( .A(n49417), .B(\reg_yHat[9][0] ), .X(n25352) );
  nor_x1_sg U73203 ( .A(n49703), .B(\reg_yHat[10][0] ), .X(n25631) );
  nor_x1_sg U73204 ( .A(n49989), .B(\reg_yHat[11][0] ), .X(n25908) );
  nor_x1_sg U73205 ( .A(n50562), .B(\reg_yHat[13][0] ), .X(n26468) );
  nor_x1_sg U73206 ( .A(n50849), .B(\reg_yHat[14][0] ), .X(n26746) );
  nor_x1_sg U73207 ( .A(n50275), .B(\reg_yHat[12][0] ), .X(n26177) );
  nor_x1_sg U73208 ( .A(n42030), .B(\reg_y[12][18] ), .X(n26036) );
  nor_x1_sg U73209 ( .A(n50547), .B(\reg_yHat[12][18] ), .X(n26037) );
  inv_x1_sg U73210 ( .A(\reg_y[12][18] ), .X(n50547) );
  nor_x1_sg U73211 ( .A(n22817), .B(n46867), .X(n22812) );
  nor_x1_sg U73212 ( .A(n46635), .B(\reg_y[0][5] ), .X(n22817) );
  nand_x1_sg U73213 ( .A(\reg_y[0][5] ), .B(n46635), .X(n22818) );
  nor_x1_sg U73214 ( .A(n23094), .B(n47160), .X(n23089) );
  nor_x1_sg U73215 ( .A(n46648), .B(\reg_y[1][5] ), .X(n23094) );
  nand_x1_sg U73216 ( .A(\reg_y[1][5] ), .B(n46648), .X(n23095) );
  nor_x1_sg U73217 ( .A(n23374), .B(n47445), .X(n23369) );
  nor_x1_sg U73218 ( .A(n46662), .B(\reg_y[2][5] ), .X(n23374) );
  nand_x1_sg U73219 ( .A(\reg_y[2][5] ), .B(n46662), .X(n23375) );
  nor_x1_sg U73220 ( .A(n23653), .B(n47730), .X(n23648) );
  nor_x1_sg U73221 ( .A(n46676), .B(\reg_y[3][5] ), .X(n23653) );
  nand_x1_sg U73222 ( .A(\reg_y[3][5] ), .B(n46676), .X(n23654) );
  nor_x1_sg U73223 ( .A(n23932), .B(n48015), .X(n23927) );
  nor_x1_sg U73224 ( .A(n46690), .B(\reg_y[4][5] ), .X(n23932) );
  nand_x1_sg U73225 ( .A(\reg_y[4][5] ), .B(n46690), .X(n23933) );
  nor_x1_sg U73226 ( .A(n24211), .B(n48300), .X(n24206) );
  nor_x1_sg U73227 ( .A(n46704), .B(\reg_y[5][5] ), .X(n24211) );
  nand_x1_sg U73228 ( .A(\reg_y[5][5] ), .B(n46704), .X(n24212) );
  nor_x1_sg U73229 ( .A(n24490), .B(n48585), .X(n24485) );
  nor_x1_sg U73230 ( .A(n46718), .B(\reg_y[6][5] ), .X(n24490) );
  nand_x1_sg U73231 ( .A(\reg_y[6][5] ), .B(n46718), .X(n24491) );
  nor_x1_sg U73232 ( .A(n24768), .B(n48871), .X(n24763) );
  nor_x1_sg U73233 ( .A(n46732), .B(\reg_y[7][5] ), .X(n24768) );
  nand_x1_sg U73234 ( .A(\reg_y[7][5] ), .B(n46732), .X(n24769) );
  nor_x1_sg U73235 ( .A(n25047), .B(n49158), .X(n25042) );
  nor_x1_sg U73236 ( .A(n46746), .B(\reg_y[8][5] ), .X(n25047) );
  nand_x1_sg U73237 ( .A(\reg_y[8][5] ), .B(n46746), .X(n25048) );
  nor_x1_sg U73238 ( .A(n25326), .B(n49444), .X(n25321) );
  nor_x1_sg U73239 ( .A(n46760), .B(\reg_y[9][5] ), .X(n25326) );
  nand_x1_sg U73240 ( .A(\reg_y[9][5] ), .B(n46760), .X(n25327) );
  nor_x1_sg U73241 ( .A(n25605), .B(n49729), .X(n25600) );
  nor_x1_sg U73242 ( .A(n46774), .B(\reg_y[10][5] ), .X(n25605) );
  nand_x1_sg U73243 ( .A(\reg_y[10][5] ), .B(n46774), .X(n25606) );
  nor_x1_sg U73244 ( .A(n25882), .B(n50016), .X(n25877) );
  nor_x1_sg U73245 ( .A(n46788), .B(\reg_y[11][5] ), .X(n25882) );
  nand_x1_sg U73246 ( .A(\reg_y[11][5] ), .B(n46788), .X(n25883) );
  nor_x1_sg U73247 ( .A(n26442), .B(n50590), .X(n26437) );
  nor_x1_sg U73248 ( .A(n46815), .B(\reg_y[13][5] ), .X(n26442) );
  nand_x1_sg U73249 ( .A(\reg_y[13][5] ), .B(n46815), .X(n26443) );
  nor_x1_sg U73250 ( .A(n26720), .B(n50877), .X(n26715) );
  nor_x1_sg U73251 ( .A(n46829), .B(\reg_y[14][5] ), .X(n26720) );
  nand_x1_sg U73252 ( .A(\reg_y[14][5] ), .B(n46829), .X(n26721) );
  nor_x1_sg U73253 ( .A(n46399), .B(n5537), .X(n20318) );
  nor_x1_sg U73254 ( .A(n6210), .B(n46351), .X(n20317) );
  nor_x1_sg U73255 ( .A(n46392), .B(n5480), .X(n19792) );
  nor_x1_sg U73256 ( .A(n6207), .B(n46347), .X(n19791) );
  nor_x1_sg U73257 ( .A(n45102), .B(n5281), .X(n28246) );
  nor_x1_sg U73258 ( .A(n42340), .B(n28142), .X(n28245) );
  nor_x1_sg U73259 ( .A(n45949), .B(n5585), .X(n20650) );
  nor_x1_sg U73260 ( .A(n6687), .B(n20508), .X(n20649) );
  nor_x1_sg U73261 ( .A(n45958), .B(n5661), .X(n21420) );
  nor_x1_sg U73262 ( .A(n42343), .B(n21277), .X(n21419) );
  nor_x1_sg U73263 ( .A(n45940), .B(n5509), .X(n20010) );
  nor_x1_sg U73264 ( .A(n6655), .B(n19851), .X(n20009) );
  nor_x1_sg U73265 ( .A(n45931), .B(n5433), .X(n19206) );
  nor_x1_sg U73266 ( .A(n6664), .B(n6671), .X(n19205) );
  nor_x1_sg U73267 ( .A(n46436), .B(n5441), .X(n19351) );
  nor_x1_sg U73268 ( .A(n42333), .B(n19311), .X(n19350) );
  nor_x1_sg U73269 ( .A(n42300), .B(n20648), .X(n20645) );
  nor_x1_sg U73270 ( .A(n45950), .B(n45970), .X(n20647) );
  nor_x1_sg U73271 ( .A(n42233), .B(n20644), .X(n20641) );
  nor_x1_sg U73272 ( .A(n45995), .B(n46015), .X(n20643) );
  nor_x1_sg U73273 ( .A(n42301), .B(n20640), .X(n20637) );
  nor_x1_sg U73274 ( .A(n46040), .B(n46061), .X(n20639) );
  nor_x1_sg U73275 ( .A(n42234), .B(n20636), .X(n20633) );
  nor_x1_sg U73276 ( .A(n46086), .B(n46106), .X(n20635) );
  nor_x1_sg U73277 ( .A(n42287), .B(n20008), .X(n20005) );
  nor_x1_sg U73278 ( .A(n45941), .B(n45973), .X(n20007) );
  nor_x1_sg U73279 ( .A(n42232), .B(n20632), .X(n20629) );
  nor_x1_sg U73280 ( .A(n46131), .B(n46152), .X(n20631) );
  nor_x1_sg U73281 ( .A(n42288), .B(n20004), .X(n20001) );
  nor_x1_sg U73282 ( .A(n45986), .B(n46018), .X(n20003) );
  nor_x1_sg U73283 ( .A(n42299), .B(n20628), .X(n20625) );
  nor_x1_sg U73284 ( .A(n46177), .B(n46197), .X(n20627) );
  nor_x1_sg U73285 ( .A(n42289), .B(n20000), .X(n19997) );
  nor_x1_sg U73286 ( .A(n46031), .B(n46064), .X(n19999) );
  nor_x1_sg U73287 ( .A(n42276), .B(n19204), .X(n19201) );
  nor_x1_sg U73288 ( .A(n45932), .B(n45976), .X(n19203) );
  nor_x1_sg U73289 ( .A(n42231), .B(n20624), .X(n20621) );
  nor_x1_sg U73290 ( .A(n46222), .B(n46243), .X(n20623) );
  nor_x1_sg U73291 ( .A(n42290), .B(n19996), .X(n19993) );
  nor_x1_sg U73292 ( .A(n46077), .B(n46109), .X(n19995) );
  nor_x1_sg U73293 ( .A(n42230), .B(n19200), .X(n19197) );
  nor_x1_sg U73294 ( .A(n45977), .B(n46021), .X(n19199) );
  nor_x1_sg U73295 ( .A(n42297), .B(n20620), .X(n20617) );
  nor_x1_sg U73296 ( .A(n46268), .B(n46288), .X(n20619) );
  nor_x1_sg U73297 ( .A(n42286), .B(n19992), .X(n19989) );
  nor_x1_sg U73298 ( .A(n46122), .B(n46155), .X(n19991) );
  nor_x1_sg U73299 ( .A(n42296), .B(n20616), .X(n20613) );
  nor_x1_sg U73300 ( .A(n46313), .B(n46334), .X(n20615) );
  nor_x1_sg U73301 ( .A(n42277), .B(n19196), .X(n19193) );
  nor_x1_sg U73302 ( .A(n46022), .B(n46067), .X(n19195) );
  nor_x1_sg U73303 ( .A(n42291), .B(n19988), .X(n19985) );
  nor_x1_sg U73304 ( .A(n46168), .B(n46200), .X(n19987) );
  nor_x1_sg U73305 ( .A(n42284), .B(n20612), .X(n20609) );
  nor_x1_sg U73306 ( .A(n46355), .B(n46375), .X(n20611) );
  nor_x1_sg U73307 ( .A(n42278), .B(n19192), .X(n19189) );
  nor_x1_sg U73308 ( .A(n46068), .B(n46112), .X(n19191) );
  nor_x1_sg U73309 ( .A(n42292), .B(n19984), .X(n19981) );
  nor_x1_sg U73310 ( .A(n46213), .B(n46246), .X(n19983) );
  nor_x1_sg U73311 ( .A(n42268), .B(n19188), .X(n19185) );
  nor_x1_sg U73312 ( .A(n46113), .B(n46158), .X(n19187) );
  nor_x1_sg U73313 ( .A(n42293), .B(n19980), .X(n19977) );
  nor_x1_sg U73314 ( .A(n46259), .B(n46291), .X(n19979) );
  nor_x1_sg U73315 ( .A(n42279), .B(n19184), .X(n19181) );
  nor_x1_sg U73316 ( .A(n46159), .B(n46203), .X(n19183) );
  nor_x1_sg U73317 ( .A(n42280), .B(n19180), .X(n19177) );
  nor_x1_sg U73318 ( .A(n46204), .B(n46249), .X(n19179) );
  nor_x1_sg U73319 ( .A(n42281), .B(n19176), .X(n19173) );
  nor_x1_sg U73320 ( .A(n46250), .B(n46294), .X(n19175) );
  nor_x1_sg U73321 ( .A(n42263), .B(n21418), .X(n21415) );
  nor_x1_sg U73322 ( .A(n45959), .B(n45967), .X(n21417) );
  nor_x1_sg U73323 ( .A(n42264), .B(n21414), .X(n21411) );
  nor_x1_sg U73324 ( .A(n46004), .B(n46012), .X(n21413) );
  nor_x1_sg U73325 ( .A(n42265), .B(n21410), .X(n21407) );
  nor_x1_sg U73326 ( .A(n46049), .B(n46058), .X(n21409) );
  nor_x1_sg U73327 ( .A(n42266), .B(n21406), .X(n21403) );
  nor_x1_sg U73328 ( .A(n46095), .B(n46103), .X(n21405) );
  nor_x1_sg U73329 ( .A(n42267), .B(n21402), .X(n21399) );
  nor_x1_sg U73330 ( .A(n46140), .B(n46149), .X(n21401) );
  nor_x1_sg U73331 ( .A(n42269), .B(n21398), .X(n21395) );
  nor_x1_sg U73332 ( .A(n46186), .B(n46194), .X(n21397) );
  nor_x1_sg U73333 ( .A(n42270), .B(n21394), .X(n21391) );
  nor_x1_sg U73334 ( .A(n46231), .B(n46240), .X(n21393) );
  nor_x1_sg U73335 ( .A(n42271), .B(n21390), .X(n21387) );
  nor_x1_sg U73336 ( .A(n46277), .B(n46285), .X(n21389) );
  nor_x1_sg U73337 ( .A(n42272), .B(n21386), .X(n21383) );
  nor_x1_sg U73338 ( .A(n46322), .B(n46331), .X(n21385) );
  nor_x1_sg U73339 ( .A(n42273), .B(n21382), .X(n21379) );
  nor_x1_sg U73340 ( .A(n46364), .B(n46372), .X(n21381) );
  nor_x1_sg U73341 ( .A(n42274), .B(n21378), .X(n21375) );
  nor_x1_sg U73342 ( .A(n46411), .B(n46420), .X(n21377) );
  nor_x1_sg U73343 ( .A(n42275), .B(n21374), .X(n21371) );
  nor_x1_sg U73344 ( .A(n46459), .B(n46467), .X(n21373) );
  nor_x1_sg U73345 ( .A(n6193), .B(n20608), .X(n20605) );
  nor_x1_sg U73346 ( .A(n46402), .B(n46423), .X(n20607) );
  nor_x1_sg U73347 ( .A(n22401), .B(n28244), .X(n28241) );
  nor_x1_sg U73348 ( .A(n45103), .B(n45127), .X(n28243) );
  nor_x1_sg U73349 ( .A(n22354), .B(n28240), .X(n28237) );
  nor_x1_sg U73350 ( .A(n45149), .B(n45172), .X(n28239) );
  nor_x1_sg U73351 ( .A(n22306), .B(n28236), .X(n28233) );
  nor_x1_sg U73352 ( .A(n45194), .B(n45218), .X(n28235) );
  nor_x1_sg U73353 ( .A(n22259), .B(n28232), .X(n28229) );
  nor_x1_sg U73354 ( .A(n45240), .B(n45263), .X(n28231) );
  nor_x1_sg U73355 ( .A(n22211), .B(n28228), .X(n28225) );
  nor_x1_sg U73356 ( .A(n45285), .B(n45308), .X(n28227) );
  nor_x1_sg U73357 ( .A(n22164), .B(n28224), .X(n28221) );
  nor_x1_sg U73358 ( .A(n45330), .B(n45353), .X(n28223) );
  nor_x1_sg U73359 ( .A(n22116), .B(n28220), .X(n28217) );
  nor_x1_sg U73360 ( .A(n45375), .B(n45399), .X(n28219) );
  nor_x1_sg U73361 ( .A(n6162), .B(n19790), .X(n19787) );
  nor_x1_sg U73362 ( .A(n46393), .B(n46430), .X(n19789) );
  nor_x1_sg U73363 ( .A(n38147), .B(n44969), .X(n28122) );
  nor_x1_sg U73364 ( .A(n28123), .B(n5725), .X(n28121) );
  nor_x1_sg U73365 ( .A(n41970), .B(n20116), .X(n20156) );
  nor_x1_sg U73366 ( .A(n46397), .B(n20113), .X(n20158) );
  nor_x1_sg U73367 ( .A(n41953), .B(n19722), .X(n19780) );
  nor_x1_sg U73368 ( .A(n46484), .B(n19719), .X(n19782) );
  nor_x1_sg U73369 ( .A(n42153), .B(n28216), .X(n28213) );
  nor_x1_sg U73370 ( .A(n45421), .B(n28180), .X(n28215) );
  nor_x1_sg U73371 ( .A(n41969), .B(n21370), .X(n21367) );
  nor_x1_sg U73372 ( .A(n46497), .B(n21341), .X(n21369) );
  nor_x1_sg U73373 ( .A(n42154), .B(n28082), .X(n28078) );
  nor_x1_sg U73374 ( .A(n45465), .B(n28081), .X(n28080) );
  nor_x1_sg U73375 ( .A(n42155), .B(n27920), .X(n27916) );
  nor_x1_sg U73376 ( .A(n45489), .B(n27919), .X(n27918) );
  nor_x1_sg U73377 ( .A(n42156), .B(n27743), .X(n27739) );
  nor_x1_sg U73378 ( .A(n45533), .B(n27742), .X(n27741) );
  nor_x1_sg U73379 ( .A(n42157), .B(n27549), .X(n27545) );
  nor_x1_sg U73380 ( .A(n45578), .B(n27548), .X(n27547) );
  nor_x1_sg U73381 ( .A(n42158), .B(n27336), .X(n27332) );
  nor_x1_sg U73382 ( .A(n27335), .B(n45622), .X(n27334) );
  nor_x1_sg U73383 ( .A(n20435), .B(n46353), .X(n20434) );
  nor_x1_sg U73384 ( .A(n20437), .B(n5556), .X(n20435) );
  nand_x1_sg U73385 ( .A(n5556), .B(n20437), .X(n20436) );
  nor_x1_sg U73386 ( .A(n42229), .B(n45826), .X(n21060) );
  nor_x1_sg U73387 ( .A(n20855), .B(n20851), .X(n21062) );
  nor_x1_sg U73388 ( .A(n42227), .B(n45842), .X(n20351) );
  nor_x1_sg U73389 ( .A(n20212), .B(n20208), .X(n20353) );
  nor_x1_sg U73390 ( .A(n42225), .B(n45858), .X(n19618) );
  nor_x1_sg U73391 ( .A(n19406), .B(n19402), .X(n19620) );
  nor_x1_sg U73392 ( .A(n42226), .B(n46445), .X(n19964) );
  nor_x1_sg U73393 ( .A(n19916), .B(n19912), .X(n19966) );
  nor_x1_sg U73394 ( .A(n46537), .B(n5628), .X(n21168) );
  nor_x1_sg U73395 ( .A(n38539), .B(n21170), .X(n21169) );
  nor_x1_sg U73396 ( .A(n46510), .B(n5552), .X(n19940) );
  nor_x1_sg U73397 ( .A(n38540), .B(n19755), .X(n19941) );
  nor_x1_sg U73398 ( .A(n41536), .B(n45822), .X(n21250) );
  inv_x1_sg U73399 ( .A(n21081), .X(n45822) );
  nor_x1_sg U73400 ( .A(n41535), .B(n45838), .X(n20482) );
  inv_x1_sg U73401 ( .A(n20372), .X(n45838) );
  nor_x1_sg U73402 ( .A(n41534), .B(n45854), .X(n19825) );
  inv_x1_sg U73403 ( .A(n19639), .X(n45854) );
  nor_x1_sg U73404 ( .A(n38541), .B(n5414), .X(n29157) );
  nor_x1_sg U73405 ( .A(n38154), .B(out_L1[3]), .X(n29156) );
  nor_x1_sg U73406 ( .A(n38542), .B(n5412), .X(n29169) );
  nor_x1_sg U73407 ( .A(n38155), .B(out_L1[5]), .X(n29168) );
  nor_x1_sg U73408 ( .A(n38543), .B(n5410), .X(n29181) );
  nor_x1_sg U73409 ( .A(n38156), .B(out_L1[7]), .X(n29180) );
  nor_x1_sg U73410 ( .A(n38544), .B(n5408), .X(n29193) );
  nor_x1_sg U73411 ( .A(n38162), .B(out_L1[9]), .X(n29192) );
  nor_x1_sg U73412 ( .A(n38545), .B(n5406), .X(n29205) );
  nor_x1_sg U73413 ( .A(n38163), .B(out_L1[11]), .X(n29204) );
  nor_x1_sg U73414 ( .A(n38546), .B(n5404), .X(n29217) );
  nor_x1_sg U73415 ( .A(n38164), .B(out_L1[13]), .X(n29216) );
  nor_x1_sg U73416 ( .A(n38547), .B(n5402), .X(n29269) );
  nor_x1_sg U73417 ( .A(n38166), .B(out_L1[15]), .X(n29268) );
  nor_x1_sg U73418 ( .A(n38548), .B(n5699), .X(n21606) );
  nor_x1_sg U73419 ( .A(n38161), .B(out_L2[3]), .X(n21605) );
  nor_x1_sg U73420 ( .A(n38549), .B(n5687), .X(n21718) );
  nor_x1_sg U73421 ( .A(n38165), .B(out_L2[15]), .X(n21717) );
  nor_x1_sg U73422 ( .A(n38550), .B(n5689), .X(n21666) );
  nor_x1_sg U73423 ( .A(n38167), .B(out_L2[13]), .X(n21665) );
  nor_x1_sg U73424 ( .A(n38551), .B(n5691), .X(n21654) );
  nor_x1_sg U73425 ( .A(n38157), .B(out_L2[11]), .X(n21653) );
  nor_x1_sg U73426 ( .A(n38552), .B(n5693), .X(n21642) );
  nor_x1_sg U73427 ( .A(n38158), .B(out_L2[9]), .X(n21641) );
  nor_x1_sg U73428 ( .A(n38553), .B(n5695), .X(n21630) );
  nor_x1_sg U73429 ( .A(n38159), .B(out_L2[7]), .X(n21629) );
  nor_x1_sg U73430 ( .A(n38554), .B(n5697), .X(n21618) );
  nor_x1_sg U73431 ( .A(n38160), .B(out_L2[5]), .X(n21617) );
  nand_x1_sg U73432 ( .A(n39929), .B(reg_num[0]), .X(n29272) );
  nor_x1_sg U73433 ( .A(\reg_yHat[1][3] ), .B(n23102), .X(n23101) );
  nor_x1_sg U73434 ( .A(\reg_yHat[2][3] ), .B(n23382), .X(n23381) );
  nor_x1_sg U73435 ( .A(\reg_yHat[3][3] ), .B(n23661), .X(n23660) );
  nor_x1_sg U73436 ( .A(\reg_yHat[4][3] ), .B(n23940), .X(n23939) );
  nor_x1_sg U73437 ( .A(\reg_yHat[5][3] ), .B(n24219), .X(n24218) );
  nor_x1_sg U73438 ( .A(\reg_yHat[6][3] ), .B(n24498), .X(n24497) );
  nor_x1_sg U73439 ( .A(\reg_yHat[7][3] ), .B(n24776), .X(n24775) );
  nor_x1_sg U73440 ( .A(\reg_yHat[8][3] ), .B(n25055), .X(n25054) );
  nor_x1_sg U73441 ( .A(\reg_yHat[9][3] ), .B(n25334), .X(n25333) );
  nor_x1_sg U73442 ( .A(\reg_yHat[10][3] ), .B(n25613), .X(n25612) );
  nor_x1_sg U73443 ( .A(\reg_yHat[11][3] ), .B(n25890), .X(n25889) );
  nor_x1_sg U73444 ( .A(\reg_yHat[13][3] ), .B(n26450), .X(n26449) );
  nor_x1_sg U73445 ( .A(\reg_yHat[14][3] ), .B(n26728), .X(n26727) );
  nor_x1_sg U73446 ( .A(\reg_yHat[0][3] ), .B(n22824), .X(n22823) );
  nor_x1_sg U73447 ( .A(n42040), .B(\reg_y[0][18] ), .X(n22722) );
  nor_x1_sg U73448 ( .A(n47119), .B(\reg_yHat[0][18] ), .X(n22723) );
  inv_x1_sg U73449 ( .A(\reg_y[0][18] ), .X(n47119) );
  nor_x1_sg U73450 ( .A(n23103), .B(n47150), .X(n23098) );
  nor_x1_sg U73451 ( .A(n46647), .B(\reg_y[1][4] ), .X(n23103) );
  nand_x1_sg U73452 ( .A(\reg_y[1][4] ), .B(n46647), .X(n23104) );
  nor_x1_sg U73453 ( .A(n23383), .B(n47435), .X(n23378) );
  nor_x1_sg U73454 ( .A(n46661), .B(\reg_y[2][4] ), .X(n23383) );
  nand_x1_sg U73455 ( .A(\reg_y[2][4] ), .B(n46661), .X(n23384) );
  nor_x1_sg U73456 ( .A(n23662), .B(n47720), .X(n23657) );
  nor_x1_sg U73457 ( .A(n46675), .B(\reg_y[3][4] ), .X(n23662) );
  nand_x1_sg U73458 ( .A(\reg_y[3][4] ), .B(n46675), .X(n23663) );
  nor_x1_sg U73459 ( .A(n23941), .B(n48005), .X(n23936) );
  nor_x1_sg U73460 ( .A(n46689), .B(\reg_y[4][4] ), .X(n23941) );
  nand_x1_sg U73461 ( .A(\reg_y[4][4] ), .B(n46689), .X(n23942) );
  nor_x1_sg U73462 ( .A(n24220), .B(n48290), .X(n24215) );
  nor_x1_sg U73463 ( .A(n46703), .B(\reg_y[5][4] ), .X(n24220) );
  nand_x1_sg U73464 ( .A(\reg_y[5][4] ), .B(n46703), .X(n24221) );
  nor_x1_sg U73465 ( .A(n24499), .B(n48575), .X(n24494) );
  nor_x1_sg U73466 ( .A(n46717), .B(\reg_y[6][4] ), .X(n24499) );
  nand_x1_sg U73467 ( .A(\reg_y[6][4] ), .B(n46717), .X(n24500) );
  nor_x1_sg U73468 ( .A(n24777), .B(n48861), .X(n24772) );
  nor_x1_sg U73469 ( .A(n46731), .B(\reg_y[7][4] ), .X(n24777) );
  nand_x1_sg U73470 ( .A(\reg_y[7][4] ), .B(n46731), .X(n24778) );
  nor_x1_sg U73471 ( .A(n25056), .B(n49148), .X(n25051) );
  nor_x1_sg U73472 ( .A(n46745), .B(\reg_y[8][4] ), .X(n25056) );
  nand_x1_sg U73473 ( .A(\reg_y[8][4] ), .B(n46745), .X(n25057) );
  nor_x1_sg U73474 ( .A(n25335), .B(n49434), .X(n25330) );
  nor_x1_sg U73475 ( .A(n46759), .B(\reg_y[9][4] ), .X(n25335) );
  nand_x1_sg U73476 ( .A(\reg_y[9][4] ), .B(n46759), .X(n25336) );
  nor_x1_sg U73477 ( .A(n25614), .B(n49719), .X(n25609) );
  nor_x1_sg U73478 ( .A(n46773), .B(\reg_y[10][4] ), .X(n25614) );
  nand_x1_sg U73479 ( .A(\reg_y[10][4] ), .B(n46773), .X(n25615) );
  nor_x1_sg U73480 ( .A(n25891), .B(n50006), .X(n25886) );
  nor_x1_sg U73481 ( .A(n46787), .B(\reg_y[11][4] ), .X(n25891) );
  nand_x1_sg U73482 ( .A(\reg_y[11][4] ), .B(n46787), .X(n25892) );
  nor_x1_sg U73483 ( .A(n26451), .B(n50580), .X(n26446) );
  nor_x1_sg U73484 ( .A(n46814), .B(\reg_y[13][4] ), .X(n26451) );
  nand_x1_sg U73485 ( .A(\reg_y[13][4] ), .B(n46814), .X(n26452) );
  nor_x1_sg U73486 ( .A(n26729), .B(n50867), .X(n26724) );
  nor_x1_sg U73487 ( .A(n46828), .B(\reg_y[14][4] ), .X(n26729) );
  nand_x1_sg U73488 ( .A(\reg_y[14][4] ), .B(n46828), .X(n26730) );
  nor_x1_sg U73489 ( .A(n22826), .B(n46857), .X(n22821) );
  nor_x1_sg U73490 ( .A(n46634), .B(\reg_y[0][4] ), .X(n22826) );
  nand_x1_sg U73491 ( .A(\reg_y[0][4] ), .B(n46634), .X(n22827) );
  nor_x1_sg U73492 ( .A(n42041), .B(\reg_y[1][6] ), .X(n23085) );
  nor_x1_sg U73493 ( .A(n47171), .B(\reg_yHat[1][6] ), .X(n23086) );
  nor_x1_sg U73494 ( .A(n42035), .B(\reg_y[2][6] ), .X(n23365) );
  nor_x1_sg U73495 ( .A(n47456), .B(\reg_yHat[2][6] ), .X(n23366) );
  nor_x1_sg U73496 ( .A(n42036), .B(\reg_y[3][6] ), .X(n23644) );
  nor_x1_sg U73497 ( .A(n47741), .B(\reg_yHat[3][6] ), .X(n23645) );
  nor_x1_sg U73498 ( .A(n42037), .B(\reg_y[4][6] ), .X(n23923) );
  nor_x1_sg U73499 ( .A(n48026), .B(\reg_yHat[4][6] ), .X(n23924) );
  nor_x1_sg U73500 ( .A(n42038), .B(\reg_y[5][6] ), .X(n24202) );
  nor_x1_sg U73501 ( .A(n48311), .B(\reg_yHat[5][6] ), .X(n24203) );
  nor_x1_sg U73502 ( .A(n42031), .B(\reg_y[6][6] ), .X(n24481) );
  nor_x1_sg U73503 ( .A(n48596), .B(\reg_yHat[6][6] ), .X(n24482) );
  nor_x1_sg U73504 ( .A(n42032), .B(\reg_y[7][6] ), .X(n24759) );
  nor_x1_sg U73505 ( .A(n48882), .B(\reg_yHat[7][6] ), .X(n24760) );
  nor_x1_sg U73506 ( .A(n42033), .B(\reg_y[8][6] ), .X(n25038) );
  nor_x1_sg U73507 ( .A(n49169), .B(\reg_yHat[8][6] ), .X(n25039) );
  nor_x1_sg U73508 ( .A(n42034), .B(\reg_y[9][6] ), .X(n25317) );
  nor_x1_sg U73509 ( .A(n49455), .B(\reg_yHat[9][6] ), .X(n25318) );
  nor_x1_sg U73510 ( .A(n42027), .B(\reg_y[10][6] ), .X(n25596) );
  nor_x1_sg U73511 ( .A(n49740), .B(\reg_yHat[10][6] ), .X(n25597) );
  nor_x1_sg U73512 ( .A(n42028), .B(\reg_y[11][6] ), .X(n25873) );
  nor_x1_sg U73513 ( .A(n50027), .B(\reg_yHat[11][6] ), .X(n25874) );
  nor_x1_sg U73514 ( .A(n42025), .B(\reg_y[13][6] ), .X(n26433) );
  nor_x1_sg U73515 ( .A(n50601), .B(\reg_yHat[13][6] ), .X(n26434) );
  nor_x1_sg U73516 ( .A(n42026), .B(\reg_y[14][6] ), .X(n26711) );
  nor_x1_sg U73517 ( .A(n50888), .B(\reg_yHat[14][6] ), .X(n26712) );
  nor_x1_sg U73518 ( .A(n42039), .B(\reg_y[0][6] ), .X(n22808) );
  nor_x1_sg U73519 ( .A(n46878), .B(\reg_yHat[0][6] ), .X(n22809) );
  nor_x1_sg U73520 ( .A(n42029), .B(\reg_y[12][6] ), .X(n26097) );
  nor_x1_sg U73521 ( .A(n50312), .B(\reg_yHat[12][6] ), .X(n26098) );
  nor_x1_sg U73522 ( .A(n38555), .B(out_L1[1]), .X(n29144) );
  nor_x1_sg U73523 ( .A(n19315), .B(n46438), .X(n19314) );
  nor_x1_sg U73524 ( .A(n46437), .B(n5440), .X(n19315) );
  nand_x1_sg U73525 ( .A(n5440), .B(n46437), .X(n19316) );
  nor_x1_sg U73526 ( .A(n26109), .B(n50290), .X(n26106) );
  nor_x1_sg U73527 ( .A(n46801), .B(\reg_y[12][4] ), .X(n26109) );
  nand_x1_sg U73528 ( .A(\reg_y[12][4] ), .B(n46801), .X(n26110) );
  nor_x1_sg U73529 ( .A(\reg_y[0][17] ), .B(n7014), .X(n7012) );
  nor_x1_sg U73530 ( .A(\reg_yHat[0][17] ), .B(n7015), .X(n7014) );
  nor_x1_sg U73531 ( .A(\reg_y[1][17] ), .B(n7832), .X(n7830) );
  nor_x1_sg U73532 ( .A(\reg_yHat[1][17] ), .B(n7833), .X(n7832) );
  nor_x1_sg U73533 ( .A(\reg_y[2][17] ), .B(n8650), .X(n8648) );
  nor_x1_sg U73534 ( .A(\reg_yHat[2][17] ), .B(n8651), .X(n8650) );
  nor_x1_sg U73535 ( .A(\reg_y[3][17] ), .B(n9470), .X(n9468) );
  nor_x1_sg U73536 ( .A(\reg_yHat[3][17] ), .B(n9471), .X(n9470) );
  nor_x1_sg U73537 ( .A(\reg_y[4][17] ), .B(n10289), .X(n10287) );
  nor_x1_sg U73538 ( .A(\reg_yHat[4][17] ), .B(n10290), .X(n10289) );
  nor_x1_sg U73539 ( .A(\reg_y[5][17] ), .B(n11108), .X(n11106) );
  nor_x1_sg U73540 ( .A(\reg_yHat[5][17] ), .B(n11109), .X(n11108) );
  nor_x1_sg U73541 ( .A(\reg_y[6][17] ), .B(n11927), .X(n11925) );
  nor_x1_sg U73542 ( .A(\reg_yHat[6][17] ), .B(n11928), .X(n11927) );
  nor_x1_sg U73543 ( .A(\reg_y[7][17] ), .B(n12746), .X(n12744) );
  nor_x1_sg U73544 ( .A(\reg_yHat[7][17] ), .B(n12747), .X(n12746) );
  nor_x1_sg U73545 ( .A(\reg_y[8][17] ), .B(n13565), .X(n13563) );
  nor_x1_sg U73546 ( .A(\reg_yHat[8][17] ), .B(n13566), .X(n13565) );
  nor_x1_sg U73547 ( .A(\reg_y[9][17] ), .B(n14384), .X(n14382) );
  nor_x1_sg U73548 ( .A(\reg_yHat[9][17] ), .B(n14385), .X(n14384) );
  nor_x1_sg U73549 ( .A(\reg_y[10][17] ), .B(n15203), .X(n15201) );
  nor_x1_sg U73550 ( .A(\reg_yHat[10][17] ), .B(n15204), .X(n15203) );
  nor_x1_sg U73551 ( .A(\reg_y[11][17] ), .B(n16022), .X(n16020) );
  nor_x1_sg U73552 ( .A(\reg_yHat[11][17] ), .B(n16023), .X(n16022) );
  nor_x1_sg U73553 ( .A(\reg_y[13][17] ), .B(n17660), .X(n17658) );
  nor_x1_sg U73554 ( .A(\reg_yHat[13][17] ), .B(n17661), .X(n17660) );
  nor_x1_sg U73555 ( .A(\reg_y[14][17] ), .B(n18481), .X(n18479) );
  nor_x1_sg U73556 ( .A(\reg_yHat[14][17] ), .B(n18482), .X(n18481) );
  nor_x1_sg U73557 ( .A(n28986), .B(n28987), .X(n28984) );
  nor_x1_sg U73558 ( .A(n28988), .B(n5397), .X(n28987) );
  nor_x1_sg U73559 ( .A(n28815), .B(n28816), .X(n28813) );
  nor_x1_sg U73560 ( .A(n28817), .B(n5378), .X(n28816) );
  nor_x1_sg U73561 ( .A(n28627), .B(n28628), .X(n28625) );
  nor_x1_sg U73562 ( .A(n28629), .B(n5359), .X(n28628) );
  nor_x1_sg U73563 ( .A(n28466), .B(n28467), .X(n28465) );
  nor_x1_sg U73564 ( .A(n28468), .B(n5340), .X(n28467) );
  nor_x1_sg U73565 ( .A(n28372), .B(n28373), .X(n28370) );
  nor_x1_sg U73566 ( .A(n28374), .B(n5321), .X(n28373) );
  nor_x1_sg U73567 ( .A(n28259), .B(n28260), .X(n28258) );
  nor_x1_sg U73568 ( .A(n28261), .B(n5302), .X(n28260) );
  nor_x1_sg U73569 ( .A(n27975), .B(n27976), .X(n27973) );
  nor_x1_sg U73570 ( .A(n27977), .B(n5264), .X(n27976) );
  nor_x1_sg U73571 ( .A(n27806), .B(n27807), .X(n27804) );
  nor_x1_sg U73572 ( .A(n27808), .B(n5245), .X(n27807) );
  nor_x1_sg U73573 ( .A(n27620), .B(n27621), .X(n27619) );
  nor_x1_sg U73574 ( .A(n27622), .B(n5226), .X(n27621) );
  nor_x1_sg U73575 ( .A(n27417), .B(n27418), .X(n27415) );
  nor_x1_sg U73576 ( .A(n27419), .B(n5207), .X(n27418) );
  nor_x1_sg U73577 ( .A(n27195), .B(n27196), .X(n27194) );
  nor_x1_sg U73578 ( .A(n27197), .B(n5188), .X(n27196) );
  nor_x1_sg U73579 ( .A(n21435), .B(n21436), .X(n21433) );
  nor_x1_sg U73580 ( .A(n21437), .B(n5682), .X(n21436) );
  nor_x1_sg U73581 ( .A(n26956), .B(n26957), .X(n26953) );
  nor_x1_sg U73582 ( .A(n26958), .B(n5169), .X(n26957) );
  nor_x1_sg U73583 ( .A(n28128), .B(n28129), .X(n28126) );
  nor_x1_sg U73584 ( .A(n22535), .B(n5283), .X(n28129) );
  nor_x1_sg U73585 ( .A(n21073), .B(n21074), .X(n21071) );
  nor_x1_sg U73586 ( .A(n6772), .B(n5644), .X(n21074) );
  nor_x1_sg U73587 ( .A(n20665), .B(n20666), .X(n20663) );
  nor_x1_sg U73588 ( .A(n6782), .B(n5606), .X(n20666) );
  nor_x1_sg U73589 ( .A(n20494), .B(n20495), .X(n20492) );
  nor_x1_sg U73590 ( .A(n6777), .B(n5587), .X(n20495) );
  nor_x1_sg U73591 ( .A(n20025), .B(n20026), .X(n20023) );
  nor_x1_sg U73592 ( .A(n6748), .B(n5530), .X(n20026) );
  nor_x1_sg U73593 ( .A(n20364), .B(n20365), .X(n20362) );
  nor_x1_sg U73594 ( .A(n6778), .B(n5568), .X(n20365) );
  nor_x1_sg U73595 ( .A(n19837), .B(n19838), .X(n19835) );
  nor_x1_sg U73596 ( .A(n6743), .B(n5511), .X(n19838) );
  nor_x1_sg U73597 ( .A(n19631), .B(n19632), .X(n19629) );
  nor_x1_sg U73598 ( .A(n6744), .B(n5492), .X(n19632) );
  nor_x1_sg U73599 ( .A(n19398), .B(n19399), .X(n19396) );
  nor_x1_sg U73600 ( .A(n6763), .B(n5473), .X(n19399) );
  nor_x1_sg U73601 ( .A(n19221), .B(n19222), .X(n19219) );
  nor_x1_sg U73602 ( .A(n6764), .B(n5454), .X(n19222) );
  nor_x1_sg U73603 ( .A(n6759), .B(n6760), .X(n6756) );
  nor_x1_sg U73604 ( .A(n6753), .B(n5435), .X(n6760) );
  nor_x1_sg U73605 ( .A(n20204), .B(n20205), .X(n20202) );
  nor_x1_sg U73606 ( .A(n6747), .B(n5549), .X(n20205) );
  nor_x1_sg U73607 ( .A(n21263), .B(n21264), .X(n21261) );
  nor_x1_sg U73608 ( .A(n6771), .B(n5663), .X(n21264) );
  nor_x1_sg U73609 ( .A(n20847), .B(n20848), .X(n20845) );
  nor_x1_sg U73610 ( .A(n6781), .B(n5625), .X(n20848) );
  nand_x1_sg U73611 ( .A(n28981), .B(n38196), .X(n28979) );
  nor_x1_sg U73612 ( .A(n22992), .B(n46659), .X(n22989) );
  nor_x1_sg U73613 ( .A(n47382), .B(\reg_y[1][18] ), .X(n22990) );
  nor_x1_sg U73614 ( .A(n23272), .B(n46673), .X(n23269) );
  nor_x1_sg U73615 ( .A(n47667), .B(\reg_y[2][18] ), .X(n23270) );
  nor_x1_sg U73616 ( .A(n23551), .B(n46687), .X(n23548) );
  nor_x1_sg U73617 ( .A(n47952), .B(\reg_y[3][18] ), .X(n23549) );
  nor_x1_sg U73618 ( .A(n23830), .B(n46701), .X(n23827) );
  nor_x1_sg U73619 ( .A(n48237), .B(\reg_y[4][18] ), .X(n23828) );
  nor_x1_sg U73620 ( .A(n24109), .B(n46715), .X(n24106) );
  nor_x1_sg U73621 ( .A(n48522), .B(\reg_y[5][18] ), .X(n24107) );
  nor_x1_sg U73622 ( .A(n24388), .B(n46729), .X(n24385) );
  nor_x1_sg U73623 ( .A(n48807), .B(\reg_y[6][18] ), .X(n24386) );
  nor_x1_sg U73624 ( .A(n24666), .B(n46743), .X(n24663) );
  nor_x1_sg U73625 ( .A(n49094), .B(\reg_y[7][18] ), .X(n24664) );
  nor_x1_sg U73626 ( .A(n24945), .B(n46757), .X(n24942) );
  nor_x1_sg U73627 ( .A(n49380), .B(\reg_y[8][18] ), .X(n24943) );
  nor_x1_sg U73628 ( .A(n25224), .B(n46771), .X(n25221) );
  nor_x1_sg U73629 ( .A(n49666), .B(\reg_y[9][18] ), .X(n25222) );
  nor_x1_sg U73630 ( .A(n25503), .B(n46785), .X(n25500) );
  nor_x1_sg U73631 ( .A(n49952), .B(\reg_y[10][18] ), .X(n25501) );
  nor_x1_sg U73632 ( .A(n25780), .B(n46799), .X(n25777) );
  nor_x1_sg U73633 ( .A(n50238), .B(\reg_y[11][18] ), .X(n25778) );
  nor_x1_sg U73634 ( .A(n26340), .B(n46826), .X(n26337) );
  nor_x1_sg U73635 ( .A(n50812), .B(\reg_y[13][18] ), .X(n26338) );
  nor_x1_sg U73636 ( .A(n26618), .B(n46840), .X(n26615) );
  nor_x1_sg U73637 ( .A(n51099), .B(\reg_y[14][18] ), .X(n26616) );
  nor_x1_sg U73638 ( .A(n42030), .B(n16834), .X(n26145) );
  nor_x1_sg U73639 ( .A(n26147), .B(\reg_y[12][18] ), .X(n26146) );
  nor_x1_sg U73640 ( .A(\reg_yHat[12][18] ), .B(n41526), .X(n26147) );
  nor_x1_sg U73641 ( .A(n42040), .B(n22714), .X(n22711) );
  nor_x1_sg U73642 ( .A(n22713), .B(\reg_y[0][18] ), .X(n22712) );
  nor_x1_sg U73643 ( .A(\reg_yHat[0][18] ), .B(n47096), .X(n22713) );
  nor_x1_sg U73644 ( .A(n21079), .B(n45823), .X(n21077) );
  nor_x1_sg U73645 ( .A(n21081), .B(n5643), .X(n21079) );
  nor_x1_sg U73646 ( .A(n20671), .B(n45831), .X(n20669) );
  nor_x1_sg U73647 ( .A(n20673), .B(n5605), .X(n20671) );
  nor_x1_sg U73648 ( .A(n20370), .B(n45839), .X(n20368) );
  nor_x1_sg U73649 ( .A(n20372), .B(n5567), .X(n20370) );
  nor_x1_sg U73650 ( .A(n20031), .B(n45847), .X(n20029) );
  nor_x1_sg U73651 ( .A(n20033), .B(n5529), .X(n20031) );
  nor_x1_sg U73652 ( .A(n19637), .B(n45855), .X(n19635) );
  nor_x1_sg U73653 ( .A(n19639), .B(n5491), .X(n19637) );
  nor_x1_sg U73654 ( .A(n19492), .B(n46441), .X(n19491) );
  nor_x1_sg U73655 ( .A(n19494), .B(n5459), .X(n19492) );
  nor_x1_sg U73656 ( .A(n19227), .B(n45863), .X(n19225) );
  nor_x1_sg U73657 ( .A(n19229), .B(n5453), .X(n19227) );
  nor_x1_sg U73658 ( .A(n20775), .B(n46534), .X(n20774) );
  nor_x1_sg U73659 ( .A(n20777), .B(n5590), .X(n20775) );
  nand_x1_sg U73660 ( .A(n5590), .B(n20777), .X(n20776) );
  nor_x1_sg U73661 ( .A(n20291), .B(n46401), .X(n20289) );
  nor_x1_sg U73662 ( .A(n46400), .B(n5536), .X(n20291) );
  nand_x1_sg U73663 ( .A(n5536), .B(n46400), .X(n20292) );
  nor_x1_sg U73664 ( .A(n19726), .B(n46531), .X(n19724) );
  nor_x1_sg U73665 ( .A(n46530), .B(n5476), .X(n19726) );
  nand_x1_sg U73666 ( .A(n5476), .B(n46530), .X(n19727) );
  nor_x1_sg U73667 ( .A(n20120), .B(n46448), .X(n20118) );
  nor_x1_sg U73668 ( .A(n46447), .B(n5516), .X(n20120) );
  nand_x1_sg U73669 ( .A(n5516), .B(n46447), .X(n20121) );
  nor_x1_sg U73670 ( .A(n19920), .B(n46487), .X(n19918) );
  nor_x1_sg U73671 ( .A(n46486), .B(n5496), .X(n19920) );
  nand_x1_sg U73672 ( .A(n5496), .B(n46486), .X(n19921) );
  nor_x1_sg U73673 ( .A(n46348), .B(n5499), .X(n19901) );
  nor_x1_sg U73674 ( .A(n38556), .B(n19903), .X(n19902) );
  nor_x1_sg U73675 ( .A(n26837), .B(n45776), .X(n26825) );
  nor_x1_sg U73676 ( .A(n26839), .B(n5284), .X(n26837) );
  nor_x1_sg U73677 ( .A(n26852), .B(n45775), .X(n26818) );
  nor_x1_sg U73678 ( .A(n26854), .B(n5246), .X(n26852) );
  nor_x1_sg U73679 ( .A(n26859), .B(n45774), .X(n26815) );
  nor_x1_sg U73680 ( .A(n26861), .B(n5227), .X(n26859) );
  nor_x1_sg U73681 ( .A(n26866), .B(n45773), .X(n26812) );
  nor_x1_sg U73682 ( .A(n26868), .B(n5208), .X(n26866) );
  nor_x1_sg U73683 ( .A(n28557), .B(n45779), .X(n28525) );
  nor_x1_sg U73684 ( .A(n28559), .B(n5341), .X(n28557) );
  nor_x1_sg U73685 ( .A(n26873), .B(n45772), .X(n26809) );
  nor_x1_sg U73686 ( .A(n26875), .B(n5189), .X(n26873) );
  nor_x1_sg U73687 ( .A(n20985), .B(n46616), .X(n20974) );
  nor_x1_sg U73688 ( .A(n20987), .B(n5664), .X(n20985) );
  nor_x1_sg U73689 ( .A(n28564), .B(n45778), .X(n28522) );
  nor_x1_sg U73690 ( .A(n28566), .B(n5322), .X(n28564) );
  nor_x1_sg U73691 ( .A(n28543), .B(n45781), .X(n28531) );
  nor_x1_sg U73692 ( .A(n28545), .B(n5379), .X(n28543) );
  nor_x1_sg U73693 ( .A(n26880), .B(n45771), .X(n26806) );
  nor_x1_sg U73694 ( .A(n26882), .B(n5170), .X(n26880) );
  nor_x1_sg U73695 ( .A(n26830), .B(n45777), .X(n26828) );
  nor_x1_sg U73696 ( .A(n26832), .B(n5303), .X(n26830) );
  nor_x1_sg U73697 ( .A(n28550), .B(n45780), .X(n28528) );
  nor_x1_sg U73698 ( .A(n28552), .B(n5360), .X(n28550) );
  nor_x1_sg U73699 ( .A(n26894), .B(n45769), .X(n26800) );
  nor_x1_sg U73700 ( .A(n26896), .B(n5132), .X(n26894) );
  nor_x1_sg U73701 ( .A(n26887), .B(n45770), .X(n26803) );
  nor_x1_sg U73702 ( .A(n26889), .B(n5151), .X(n26887) );
  nor_x1_sg U73703 ( .A(n38557), .B(n5684), .X(n21188) );
  nor_x1_sg U73704 ( .A(n38189), .B(out_L2[18]), .X(n21187) );
  nor_x1_sg U73705 ( .A(n38558), .B(n5399), .X(n28743) );
  nor_x1_sg U73706 ( .A(n38190), .B(out_L1[18]), .X(n28742) );
  nor_x1_sg U73707 ( .A(n44975), .B(n5717), .X(n22549) );
  nor_x1_sg U73708 ( .A(n46852), .B(n22835), .X(n22829) );
  nor_x1_sg U73709 ( .A(n46851), .B(\reg_yHat[0][3] ), .X(n22835) );
  nand_x1_sg U73710 ( .A(n38760), .B(n46851), .X(n22836) );
  nor_x1_sg U73711 ( .A(n47145), .B(n23112), .X(n23106) );
  nor_x1_sg U73712 ( .A(n47144), .B(\reg_yHat[1][3] ), .X(n23112) );
  nand_x1_sg U73713 ( .A(n38764), .B(n47144), .X(n23113) );
  nor_x1_sg U73714 ( .A(n47430), .B(n23392), .X(n23386) );
  nor_x1_sg U73715 ( .A(n47429), .B(\reg_yHat[2][3] ), .X(n23392) );
  nand_x1_sg U73716 ( .A(n38768), .B(n47429), .X(n23393) );
  nor_x1_sg U73717 ( .A(n47715), .B(n23671), .X(n23665) );
  nor_x1_sg U73718 ( .A(n47714), .B(\reg_yHat[3][3] ), .X(n23671) );
  nand_x1_sg U73719 ( .A(n38772), .B(n47714), .X(n23672) );
  nor_x1_sg U73720 ( .A(n48000), .B(n23950), .X(n23944) );
  nor_x1_sg U73721 ( .A(n47999), .B(\reg_yHat[4][3] ), .X(n23950) );
  nand_x1_sg U73722 ( .A(n38776), .B(n47999), .X(n23951) );
  nor_x1_sg U73723 ( .A(n48285), .B(n24229), .X(n24223) );
  nor_x1_sg U73724 ( .A(n48284), .B(\reg_yHat[5][3] ), .X(n24229) );
  nand_x1_sg U73725 ( .A(n38780), .B(n48284), .X(n24230) );
  nor_x1_sg U73726 ( .A(n48570), .B(n24508), .X(n24502) );
  nor_x1_sg U73727 ( .A(n48569), .B(\reg_yHat[6][3] ), .X(n24508) );
  nand_x1_sg U73728 ( .A(n38784), .B(n48569), .X(n24509) );
  nor_x1_sg U73729 ( .A(n48855), .B(n24786), .X(n24780) );
  nor_x1_sg U73730 ( .A(n48854), .B(\reg_yHat[7][3] ), .X(n24786) );
  nand_x1_sg U73731 ( .A(n38788), .B(n48854), .X(n24787) );
  nor_x1_sg U73732 ( .A(n49142), .B(n25065), .X(n25059) );
  nor_x1_sg U73733 ( .A(n49141), .B(\reg_yHat[8][3] ), .X(n25065) );
  nand_x1_sg U73734 ( .A(n38792), .B(n49141), .X(n25066) );
  nor_x1_sg U73735 ( .A(n49428), .B(n25344), .X(n25338) );
  nor_x1_sg U73736 ( .A(n49427), .B(\reg_yHat[9][3] ), .X(n25344) );
  nand_x1_sg U73737 ( .A(n38796), .B(n49427), .X(n25345) );
  nor_x1_sg U73738 ( .A(n49714), .B(n25623), .X(n25617) );
  nor_x1_sg U73739 ( .A(n49713), .B(\reg_yHat[10][3] ), .X(n25623) );
  nand_x1_sg U73740 ( .A(n38800), .B(n49713), .X(n25624) );
  nor_x1_sg U73741 ( .A(n50000), .B(n25900), .X(n25894) );
  nor_x1_sg U73742 ( .A(n49999), .B(\reg_yHat[11][3] ), .X(n25900) );
  nand_x1_sg U73743 ( .A(n38804), .B(n49999), .X(n25901) );
  nor_x1_sg U73744 ( .A(n50575), .B(n26460), .X(n26454) );
  nor_x1_sg U73745 ( .A(n50574), .B(\reg_yHat[13][3] ), .X(n26460) );
  nand_x1_sg U73746 ( .A(n38808), .B(n50574), .X(n26461) );
  nor_x1_sg U73747 ( .A(n50861), .B(n26738), .X(n26732) );
  nor_x1_sg U73748 ( .A(n50860), .B(\reg_yHat[14][3] ), .X(n26738) );
  nand_x1_sg U73749 ( .A(n38812), .B(n50860), .X(n26739) );
  nor_x1_sg U73750 ( .A(n47414), .B(n22993), .X(n22988) );
  nor_x1_sg U73751 ( .A(n47413), .B(\reg_yHat[1][19] ), .X(n22993) );
  nand_x1_sg U73752 ( .A(\reg_yHat[1][19] ), .B(n47413), .X(n22994) );
  nor_x1_sg U73753 ( .A(n47699), .B(n23273), .X(n23268) );
  nor_x1_sg U73754 ( .A(n47698), .B(\reg_yHat[2][19] ), .X(n23273) );
  nand_x1_sg U73755 ( .A(\reg_yHat[2][19] ), .B(n47698), .X(n23274) );
  nor_x1_sg U73756 ( .A(n47984), .B(n23552), .X(n23547) );
  nor_x1_sg U73757 ( .A(n47983), .B(\reg_yHat[3][19] ), .X(n23552) );
  nand_x1_sg U73758 ( .A(\reg_yHat[3][19] ), .B(n47983), .X(n23553) );
  nor_x1_sg U73759 ( .A(n48269), .B(n23831), .X(n23826) );
  nor_x1_sg U73760 ( .A(n48268), .B(\reg_yHat[4][19] ), .X(n23831) );
  nand_x1_sg U73761 ( .A(\reg_yHat[4][19] ), .B(n48268), .X(n23832) );
  nor_x1_sg U73762 ( .A(n48554), .B(n24110), .X(n24105) );
  nor_x1_sg U73763 ( .A(n48553), .B(\reg_yHat[5][19] ), .X(n24110) );
  nand_x1_sg U73764 ( .A(\reg_yHat[5][19] ), .B(n48553), .X(n24111) );
  nor_x1_sg U73765 ( .A(n48839), .B(n24389), .X(n24384) );
  nor_x1_sg U73766 ( .A(n48838), .B(\reg_yHat[6][19] ), .X(n24389) );
  nand_x1_sg U73767 ( .A(\reg_yHat[6][19] ), .B(n48838), .X(n24390) );
  nor_x1_sg U73768 ( .A(n49126), .B(n24667), .X(n24662) );
  nor_x1_sg U73769 ( .A(n49125), .B(\reg_yHat[7][19] ), .X(n24667) );
  nand_x1_sg U73770 ( .A(\reg_yHat[7][19] ), .B(n49125), .X(n24668) );
  nor_x1_sg U73771 ( .A(n49412), .B(n24946), .X(n24941) );
  nor_x1_sg U73772 ( .A(n49411), .B(\reg_yHat[8][19] ), .X(n24946) );
  nand_x1_sg U73773 ( .A(\reg_yHat[8][19] ), .B(n49411), .X(n24947) );
  nor_x1_sg U73774 ( .A(n49698), .B(n25225), .X(n25220) );
  nor_x1_sg U73775 ( .A(n49697), .B(\reg_yHat[9][19] ), .X(n25225) );
  nand_x1_sg U73776 ( .A(\reg_yHat[9][19] ), .B(n49697), .X(n25226) );
  nor_x1_sg U73777 ( .A(n49984), .B(n25504), .X(n25499) );
  nor_x1_sg U73778 ( .A(n49983), .B(\reg_yHat[10][19] ), .X(n25504) );
  nand_x1_sg U73779 ( .A(\reg_yHat[10][19] ), .B(n49983), .X(n25505) );
  nor_x1_sg U73780 ( .A(n50270), .B(n25781), .X(n25776) );
  nor_x1_sg U73781 ( .A(n50269), .B(\reg_yHat[11][19] ), .X(n25781) );
  nand_x1_sg U73782 ( .A(\reg_yHat[11][19] ), .B(n50269), .X(n25782) );
  nor_x1_sg U73783 ( .A(n50845), .B(n26341), .X(n26336) );
  nor_x1_sg U73784 ( .A(n50844), .B(\reg_yHat[13][19] ), .X(n26341) );
  nand_x1_sg U73785 ( .A(\reg_yHat[13][19] ), .B(n50844), .X(n26342) );
  nor_x1_sg U73786 ( .A(n51131), .B(n26619), .X(n26614) );
  nor_x1_sg U73787 ( .A(n51130), .B(\reg_yHat[14][19] ), .X(n26619) );
  nand_x1_sg U73788 ( .A(\reg_yHat[14][19] ), .B(n51130), .X(n26620) );
  nor_x1_sg U73789 ( .A(n47129), .B(n22715), .X(n22710) );
  nor_x1_sg U73790 ( .A(n47128), .B(\reg_yHat[0][19] ), .X(n22715) );
  nand_x1_sg U73791 ( .A(\reg_yHat[0][19] ), .B(n47128), .X(n22716) );
  nor_x1_sg U73792 ( .A(n50558), .B(n26178), .X(n26144) );
  nor_x1_sg U73793 ( .A(n50557), .B(\reg_yHat[12][19] ), .X(n26178) );
  nand_x1_sg U73794 ( .A(\reg_yHat[12][19] ), .B(n50557), .X(n26179) );
  inv_x1_sg U73795 ( .A(\reg_yHat[1][18] ), .X(n46659) );
  inv_x1_sg U73796 ( .A(\reg_yHat[2][18] ), .X(n46673) );
  inv_x1_sg U73797 ( .A(\reg_yHat[3][18] ), .X(n46687) );
  inv_x1_sg U73798 ( .A(\reg_yHat[4][18] ), .X(n46701) );
  inv_x1_sg U73799 ( .A(\reg_yHat[5][18] ), .X(n46715) );
  inv_x1_sg U73800 ( .A(\reg_yHat[6][18] ), .X(n46729) );
  inv_x1_sg U73801 ( .A(\reg_yHat[7][18] ), .X(n46743) );
  inv_x1_sg U73802 ( .A(\reg_yHat[8][18] ), .X(n46757) );
  inv_x1_sg U73803 ( .A(\reg_yHat[9][18] ), .X(n46771) );
  inv_x1_sg U73804 ( .A(\reg_yHat[10][18] ), .X(n46785) );
  inv_x1_sg U73805 ( .A(\reg_yHat[11][18] ), .X(n46799) );
  inv_x1_sg U73806 ( .A(\reg_yHat[13][18] ), .X(n46826) );
  inv_x1_sg U73807 ( .A(\reg_yHat[14][18] ), .X(n46840) );
  inv_x1_sg U73808 ( .A(\reg_yHat[0][5] ), .X(n46635) );
  inv_x1_sg U73809 ( .A(\reg_yHat[1][5] ), .X(n46648) );
  inv_x1_sg U73810 ( .A(\reg_yHat[2][5] ), .X(n46662) );
  inv_x1_sg U73811 ( .A(\reg_yHat[3][5] ), .X(n46676) );
  inv_x1_sg U73812 ( .A(\reg_yHat[4][5] ), .X(n46690) );
  inv_x1_sg U73813 ( .A(\reg_yHat[5][5] ), .X(n46704) );
  inv_x1_sg U73814 ( .A(\reg_yHat[6][5] ), .X(n46718) );
  inv_x1_sg U73815 ( .A(\reg_yHat[7][5] ), .X(n46732) );
  inv_x1_sg U73816 ( .A(\reg_yHat[8][5] ), .X(n46746) );
  inv_x1_sg U73817 ( .A(\reg_yHat[9][5] ), .X(n46760) );
  inv_x1_sg U73818 ( .A(\reg_yHat[10][5] ), .X(n46774) );
  inv_x1_sg U73819 ( .A(\reg_yHat[11][5] ), .X(n46788) );
  inv_x1_sg U73820 ( .A(\reg_yHat[13][5] ), .X(n46815) );
  inv_x1_sg U73821 ( .A(\reg_yHat[14][5] ), .X(n46829) );
  nand_x1_sg U73822 ( .A(\reg_yHat[0][17] ), .B(n47095), .X(n22721) );
  inv_x1_sg U73823 ( .A(\reg_y[0][17] ), .X(n47095) );
  nand_x1_sg U73824 ( .A(\reg_yHat[1][17] ), .B(n47381), .X(n22998) );
  inv_x1_sg U73825 ( .A(\reg_y[1][17] ), .X(n47381) );
  nand_x1_sg U73826 ( .A(\reg_yHat[2][17] ), .B(n47666), .X(n23278) );
  inv_x1_sg U73827 ( .A(\reg_y[2][17] ), .X(n47666) );
  nand_x1_sg U73828 ( .A(\reg_yHat[3][17] ), .B(n47951), .X(n23557) );
  inv_x1_sg U73829 ( .A(\reg_y[3][17] ), .X(n47951) );
  nand_x1_sg U73830 ( .A(\reg_yHat[4][17] ), .B(n48236), .X(n23836) );
  inv_x1_sg U73831 ( .A(\reg_y[4][17] ), .X(n48236) );
  nand_x1_sg U73832 ( .A(\reg_yHat[5][17] ), .B(n48521), .X(n24115) );
  inv_x1_sg U73833 ( .A(\reg_y[5][17] ), .X(n48521) );
  nand_x1_sg U73834 ( .A(\reg_yHat[6][17] ), .B(n48806), .X(n24394) );
  inv_x1_sg U73835 ( .A(\reg_y[6][17] ), .X(n48806) );
  nand_x1_sg U73836 ( .A(\reg_yHat[7][17] ), .B(n49093), .X(n24672) );
  inv_x1_sg U73837 ( .A(\reg_y[7][17] ), .X(n49093) );
  nand_x1_sg U73838 ( .A(\reg_yHat[8][17] ), .B(n49379), .X(n24951) );
  inv_x1_sg U73839 ( .A(\reg_y[8][17] ), .X(n49379) );
  nand_x1_sg U73840 ( .A(\reg_yHat[9][17] ), .B(n49665), .X(n25230) );
  inv_x1_sg U73841 ( .A(\reg_y[9][17] ), .X(n49665) );
  nand_x1_sg U73842 ( .A(\reg_yHat[10][17] ), .B(n49951), .X(n25509) );
  inv_x1_sg U73843 ( .A(\reg_y[10][17] ), .X(n49951) );
  nand_x1_sg U73844 ( .A(\reg_yHat[11][17] ), .B(n50237), .X(n25786) );
  inv_x1_sg U73845 ( .A(\reg_y[11][17] ), .X(n50237) );
  nand_x1_sg U73846 ( .A(\reg_yHat[13][17] ), .B(n50811), .X(n26346) );
  inv_x1_sg U73847 ( .A(\reg_y[13][17] ), .X(n50811) );
  nand_x1_sg U73848 ( .A(\reg_yHat[14][17] ), .B(n51098), .X(n26624) );
  inv_x1_sg U73849 ( .A(\reg_y[14][17] ), .X(n51098) );
  nand_x1_sg U73850 ( .A(\reg_y[0][17] ), .B(n42016), .X(n22719) );
  nand_x1_sg U73851 ( .A(\reg_y[1][17] ), .B(n42017), .X(n22996) );
  nand_x1_sg U73852 ( .A(\reg_y[2][17] ), .B(n42011), .X(n23276) );
  nand_x1_sg U73853 ( .A(\reg_y[3][17] ), .B(n42012), .X(n23555) );
  nand_x1_sg U73854 ( .A(\reg_y[4][17] ), .B(n42013), .X(n23834) );
  nand_x1_sg U73855 ( .A(\reg_y[5][17] ), .B(n42014), .X(n24113) );
  nand_x1_sg U73856 ( .A(\reg_y[6][17] ), .B(n42007), .X(n24392) );
  nand_x1_sg U73857 ( .A(\reg_y[7][17] ), .B(n42008), .X(n24670) );
  nand_x1_sg U73858 ( .A(\reg_y[8][17] ), .B(n42009), .X(n24949) );
  nand_x1_sg U73859 ( .A(\reg_y[9][17] ), .B(n42010), .X(n25228) );
  nand_x1_sg U73860 ( .A(\reg_y[10][17] ), .B(n42003), .X(n25507) );
  nand_x1_sg U73861 ( .A(\reg_y[11][17] ), .B(n42004), .X(n25784) );
  nand_x1_sg U73862 ( .A(\reg_y[13][17] ), .B(n42006), .X(n26344) );
  nand_x1_sg U73863 ( .A(\reg_y[14][17] ), .B(n42001), .X(n26622) );
  nand_x1_sg U73864 ( .A(\reg_yHat[12][17] ), .B(n50523), .X(n26132) );
  inv_x1_sg U73865 ( .A(\reg_y[12][17] ), .X(n50523) );
  nand_x1_sg U73866 ( .A(\reg_y[12][17] ), .B(n42005), .X(n26133) );
  nand_x1_sg U73867 ( .A(n38758), .B(n22834), .X(n22833) );
  nand_x1_sg U73868 ( .A(n45821), .B(n38148), .X(n21253) );
  nand_x1_sg U73869 ( .A(n21255), .B(n21068), .X(n21254) );
  nor_x1_sg U73870 ( .A(n5706), .B(n21073), .X(n21255) );
  nand_x1_sg U73871 ( .A(n45829), .B(n38149), .X(n20838) );
  nand_x1_sg U73872 ( .A(n20840), .B(n20660), .X(n20839) );
  nor_x1_sg U73873 ( .A(n5708), .B(n20665), .X(n20840) );
  nand_x1_sg U73874 ( .A(n45837), .B(n38150), .X(n20485) );
  nand_x1_sg U73875 ( .A(n20487), .B(n20359), .X(n20486) );
  nor_x1_sg U73876 ( .A(n5710), .B(n20364), .X(n20487) );
  nand_x1_sg U73877 ( .A(n45845), .B(n38151), .X(n20195) );
  nand_x1_sg U73878 ( .A(n20197), .B(n20020), .X(n20196) );
  nor_x1_sg U73879 ( .A(n5712), .B(n20025), .X(n20197) );
  nand_x1_sg U73880 ( .A(n45853), .B(n38152), .X(n19828) );
  nand_x1_sg U73881 ( .A(n19830), .B(n19626), .X(n19829) );
  nor_x1_sg U73882 ( .A(n5714), .B(n19631), .X(n19830) );
  nand_x1_sg U73883 ( .A(n45861), .B(n38153), .X(n19389) );
  nand_x1_sg U73884 ( .A(n19391), .B(n19216), .X(n19390) );
  nor_x1_sg U73885 ( .A(n5716), .B(n19221), .X(n19391) );
  nand_x1_sg U73886 ( .A(\reg_y[12][2] ), .B(n26172), .X(n26171) );
  nor_x1_sg U73887 ( .A(n26120), .B(\reg_yHat[12][2] ), .X(n26173) );
  inv_x1_sg U73888 ( .A(\reg_yHat[1][4] ), .X(n46647) );
  inv_x1_sg U73889 ( .A(\reg_yHat[2][4] ), .X(n46661) );
  inv_x1_sg U73890 ( .A(\reg_yHat[3][4] ), .X(n46675) );
  inv_x1_sg U73891 ( .A(\reg_yHat[4][4] ), .X(n46689) );
  inv_x1_sg U73892 ( .A(\reg_yHat[5][4] ), .X(n46703) );
  inv_x1_sg U73893 ( .A(\reg_yHat[6][4] ), .X(n46717) );
  inv_x1_sg U73894 ( .A(\reg_yHat[7][4] ), .X(n46731) );
  inv_x1_sg U73895 ( .A(\reg_yHat[8][4] ), .X(n46745) );
  inv_x1_sg U73896 ( .A(\reg_yHat[9][4] ), .X(n46759) );
  inv_x1_sg U73897 ( .A(\reg_yHat[10][4] ), .X(n46773) );
  inv_x1_sg U73898 ( .A(\reg_yHat[11][4] ), .X(n46787) );
  inv_x1_sg U73899 ( .A(\reg_yHat[13][4] ), .X(n46814) );
  inv_x1_sg U73900 ( .A(\reg_yHat[14][4] ), .X(n46828) );
  inv_x1_sg U73901 ( .A(\reg_yHat[0][4] ), .X(n46634) );
  inv_x1_sg U73902 ( .A(\reg_yHat[12][4] ), .X(n46801) );
  inv_x1_sg U73903 ( .A(\reg_yHat[12][5] ), .X(n46802) );
  nor_x1_sg U73904 ( .A(n5718), .B(n29144), .X(n29267) );
  nor_x1_sg U73905 ( .A(n5703), .B(n21593), .X(n21716) );
  nand_x1_sg U73906 ( .A(n21356), .B(n38125), .X(n21353) );
  nand_x1_sg U73907 ( .A(n28920), .B(n38126), .X(n28917) );
  nand_x1_sg U73908 ( .A(n29154), .B(n38154), .X(n29260) );
  nand_x1_sg U73909 ( .A(n5414), .B(n45022), .X(n29262) );
  nand_x1_sg U73910 ( .A(n29166), .B(n38155), .X(n29254) );
  nand_x1_sg U73911 ( .A(n5412), .B(n45112), .X(n29256) );
  nand_x1_sg U73912 ( .A(n29178), .B(n38156), .X(n29248) );
  nand_x1_sg U73913 ( .A(n5410), .B(n45203), .X(n29250) );
  nand_x1_sg U73914 ( .A(n21651), .B(n38157), .X(n21685) );
  nand_x1_sg U73915 ( .A(n5691), .B(n46235), .X(n21687) );
  nand_x1_sg U73916 ( .A(n21639), .B(n38158), .X(n21691) );
  nand_x1_sg U73917 ( .A(n5693), .B(n46144), .X(n21693) );
  nand_x1_sg U73918 ( .A(n21627), .B(n38159), .X(n21697) );
  nand_x1_sg U73919 ( .A(n5695), .B(n46053), .X(n21699) );
  nand_x1_sg U73920 ( .A(n21615), .B(n38160), .X(n21703) );
  nand_x1_sg U73921 ( .A(n5697), .B(n45963), .X(n21705) );
  nand_x1_sg U73922 ( .A(n21603), .B(n38161), .X(n21709) );
  nand_x1_sg U73923 ( .A(n5699), .B(n45870), .X(n21711) );
  nand_x1_sg U73924 ( .A(n21430), .B(n38197), .X(n21428) );
  nand_x1_sg U73925 ( .A(n22842), .B(n46842), .X(n22841) );
  nand_x1_sg U73926 ( .A(\reg_yHat[0][1] ), .B(n42046), .X(n22840) );
  nand_x1_sg U73927 ( .A(n22843), .B(n46633), .X(n22842) );
  nand_x1_sg U73928 ( .A(n23119), .B(n47135), .X(n23118) );
  nand_x1_sg U73929 ( .A(\reg_yHat[1][1] ), .B(n47134), .X(n23117) );
  nand_x1_sg U73930 ( .A(n23120), .B(n46646), .X(n23119) );
  nand_x1_sg U73931 ( .A(n23399), .B(n47420), .X(n23398) );
  nand_x1_sg U73932 ( .A(\reg_yHat[2][1] ), .B(n42057), .X(n23397) );
  nand_x1_sg U73933 ( .A(n23400), .B(n46660), .X(n23399) );
  nand_x1_sg U73934 ( .A(n23678), .B(n47705), .X(n23677) );
  nand_x1_sg U73935 ( .A(\reg_yHat[3][1] ), .B(n42056), .X(n23676) );
  nand_x1_sg U73936 ( .A(n23679), .B(n46674), .X(n23678) );
  nand_x1_sg U73937 ( .A(n23957), .B(n47990), .X(n23956) );
  nand_x1_sg U73938 ( .A(\reg_yHat[4][1] ), .B(n42055), .X(n23955) );
  nand_x1_sg U73939 ( .A(n23958), .B(n46688), .X(n23957) );
  nand_x1_sg U73940 ( .A(n24236), .B(n48275), .X(n24235) );
  nand_x1_sg U73941 ( .A(\reg_yHat[5][1] ), .B(n42054), .X(n24234) );
  nand_x1_sg U73942 ( .A(n24237), .B(n46702), .X(n24236) );
  nand_x1_sg U73943 ( .A(n24515), .B(n48560), .X(n24514) );
  nand_x1_sg U73944 ( .A(\reg_yHat[6][1] ), .B(n42053), .X(n24513) );
  nand_x1_sg U73945 ( .A(n24516), .B(n46716), .X(n24515) );
  nand_x1_sg U73946 ( .A(n24793), .B(n48845), .X(n24792) );
  nand_x1_sg U73947 ( .A(\reg_yHat[7][1] ), .B(n42052), .X(n24791) );
  nand_x1_sg U73948 ( .A(n24794), .B(n46730), .X(n24793) );
  nand_x1_sg U73949 ( .A(n25072), .B(n49132), .X(n25071) );
  nand_x1_sg U73950 ( .A(\reg_yHat[8][1] ), .B(n42051), .X(n25070) );
  nand_x1_sg U73951 ( .A(n25073), .B(n46744), .X(n25072) );
  nand_x1_sg U73952 ( .A(n25351), .B(n49418), .X(n25350) );
  nand_x1_sg U73953 ( .A(\reg_yHat[9][1] ), .B(n42050), .X(n25349) );
  nand_x1_sg U73954 ( .A(n25352), .B(n46758), .X(n25351) );
  nand_x1_sg U73955 ( .A(n25630), .B(n49704), .X(n25629) );
  nand_x1_sg U73956 ( .A(\reg_yHat[10][1] ), .B(n42049), .X(n25628) );
  nand_x1_sg U73957 ( .A(n25631), .B(n46772), .X(n25630) );
  nand_x1_sg U73958 ( .A(n25907), .B(n49990), .X(n25906) );
  nand_x1_sg U73959 ( .A(\reg_yHat[11][1] ), .B(n42048), .X(n25905) );
  nand_x1_sg U73960 ( .A(n25908), .B(n46786), .X(n25907) );
  nand_x1_sg U73961 ( .A(n26467), .B(n50563), .X(n26466) );
  nand_x1_sg U73962 ( .A(\reg_yHat[13][1] ), .B(n42047), .X(n26465) );
  nand_x1_sg U73963 ( .A(n26468), .B(n46813), .X(n26467) );
  nand_x1_sg U73964 ( .A(n26745), .B(n50851), .X(n26744) );
  nand_x1_sg U73965 ( .A(\reg_yHat[14][1] ), .B(n50850), .X(n26743) );
  nand_x1_sg U73966 ( .A(n26746), .B(n46827), .X(n26745) );
  nand_x1_sg U73967 ( .A(n26176), .B(n50276), .X(n26175) );
  nand_x1_sg U73968 ( .A(\reg_yHat[12][1] ), .B(n42043), .X(n26174) );
  nand_x1_sg U73969 ( .A(n26177), .B(n46800), .X(n26176) );
  nand_x1_sg U73970 ( .A(n26107), .B(n46801), .X(n26165) );
  nand_x1_sg U73971 ( .A(\reg_y[12][4] ), .B(n26167), .X(n26166) );
  nand_x1_sg U73972 ( .A(\reg_yHat[12][4] ), .B(n50283), .X(n26167) );
  nand_x1_sg U73973 ( .A(n20310), .B(n20309), .X(n20306) );
  nor_x1_sg U73974 ( .A(n20308), .B(n5555), .X(n20307) );
  nand_x1_sg U73975 ( .A(n20143), .B(n20142), .X(n20139) );
  nor_x1_sg U73976 ( .A(n20141), .B(n5554), .X(n20140) );
  nand_x1_sg U73977 ( .A(n46552), .B(n19938), .X(n20595) );
  nor_x1_sg U73978 ( .A(n20597), .B(n5571), .X(n20596) );
  nand_x1_sg U73979 ( .A(n46376), .B(n20437), .X(n20448) );
  nor_x1_sg U73980 ( .A(n20450), .B(n5556), .X(n20449) );
  nand_x1_sg U73981 ( .A(n29190), .B(n38162), .X(n29242) );
  nand_x1_sg U73982 ( .A(n5408), .B(n45294), .X(n29244) );
  nand_x1_sg U73983 ( .A(n29202), .B(n38163), .X(n29236) );
  nand_x1_sg U73984 ( .A(n5406), .B(n45384), .X(n29238) );
  nand_x1_sg U73985 ( .A(n29214), .B(n38164), .X(n29230) );
  nand_x1_sg U73986 ( .A(n5404), .B(n45474), .X(n29232) );
  nand_x1_sg U73987 ( .A(n21538), .B(n38165), .X(n21535) );
  nand_x1_sg U73988 ( .A(n5687), .B(n46415), .X(n21537) );
  nand_x1_sg U73989 ( .A(n29089), .B(n38166), .X(n29086) );
  nand_x1_sg U73990 ( .A(n5402), .B(n45563), .X(n29088) );
  nand_x1_sg U73991 ( .A(n21663), .B(n38167), .X(n21679) );
  nand_x1_sg U73992 ( .A(n5689), .B(n46326), .X(n21681) );
  nand_x1_sg U73993 ( .A(n44996), .B(n38168), .X(n28251) );
  nand_x1_sg U73994 ( .A(n28253), .B(n28123), .X(n28252) );
  nor_x1_sg U73995 ( .A(n5725), .B(n28128), .X(n28253) );
  nand_x1_sg U73996 ( .A(n45833), .B(n38169), .X(n20655) );
  nand_x1_sg U73997 ( .A(n20657), .B(n45803), .X(n20656) );
  nor_x1_sg U73998 ( .A(n5709), .B(n20494), .X(n20657) );
  nand_x1_sg U73999 ( .A(n45849), .B(n38170), .X(n20015) );
  nand_x1_sg U74000 ( .A(n20017), .B(n45807), .X(n20016) );
  nor_x1_sg U74001 ( .A(n5713), .B(n19837), .X(n20017) );
  nand_x1_sg U74002 ( .A(n45817), .B(n38171), .X(n21425) );
  nand_x1_sg U74003 ( .A(n21427), .B(n21258), .X(n21426) );
  nor_x1_sg U74004 ( .A(n5705), .B(n21263), .X(n21427) );
  nand_x1_sg U74005 ( .A(n45865), .B(n38172), .X(n19211) );
  nand_x1_sg U74006 ( .A(n19213), .B(n45811), .X(n19212) );
  nor_x1_sg U74007 ( .A(n5702), .B(n6759), .X(n19213) );
  nor_x1_sg U74008 ( .A(n51137), .B(reg_num[1]), .X(n5994) );
  nand_x1_sg U74009 ( .A(n38762), .B(n23111), .X(n23110) );
  nand_x1_sg U74010 ( .A(n38766), .B(n23391), .X(n23390) );
  nand_x1_sg U74011 ( .A(n38770), .B(n23670), .X(n23669) );
  nand_x1_sg U74012 ( .A(n38774), .B(n23949), .X(n23948) );
  nand_x1_sg U74013 ( .A(n38778), .B(n24228), .X(n24227) );
  nand_x1_sg U74014 ( .A(n38782), .B(n24507), .X(n24506) );
  nand_x1_sg U74015 ( .A(n38786), .B(n24785), .X(n24784) );
  nand_x1_sg U74016 ( .A(n38790), .B(n25064), .X(n25063) );
  nand_x1_sg U74017 ( .A(n38794), .B(n25343), .X(n25342) );
  nand_x1_sg U74018 ( .A(n38798), .B(n25622), .X(n25621) );
  nand_x1_sg U74019 ( .A(n38802), .B(n25899), .X(n25898) );
  nand_x1_sg U74020 ( .A(n38806), .B(n26459), .X(n26458) );
  nand_x1_sg U74021 ( .A(n38810), .B(n26737), .X(n26736) );
  nand_x1_sg U74022 ( .A(\reg_yHat[12][13] ), .B(n50436), .X(n26055) );
  inv_x1_sg U74023 ( .A(\reg_y[12][13] ), .X(n50436) );
  nand_x1_sg U74024 ( .A(\reg_yHat[12][14] ), .B(n50454), .X(n26050) );
  inv_x1_sg U74025 ( .A(\reg_y[12][14] ), .X(n50454) );
  nand_x1_sg U74026 ( .A(\reg_y[12][14] ), .B(n46810), .X(n26049) );
  inv_x1_sg U74027 ( .A(\reg_yHat[12][14] ), .X(n46810) );
  nand_x1_sg U74028 ( .A(\reg_y[12][13] ), .B(n46809), .X(n26056) );
  inv_x1_sg U74029 ( .A(\reg_yHat[12][13] ), .X(n46809) );
  nand_x1_sg U74030 ( .A(\reg_yHat[0][9] ), .B(n46923), .X(n22778) );
  inv_x1_sg U74031 ( .A(\reg_y[0][9] ), .X(n46923) );
  nand_x1_sg U74032 ( .A(\reg_yHat[0][10] ), .B(n46941), .X(n22769) );
  inv_x1_sg U74033 ( .A(\reg_y[0][10] ), .X(n46941) );
  nand_x1_sg U74034 ( .A(\reg_y[0][10] ), .B(n46639), .X(n22771) );
  inv_x1_sg U74035 ( .A(\reg_yHat[0][10] ), .X(n46639) );
  nand_x1_sg U74036 ( .A(\reg_y[0][9] ), .B(n46638), .X(n22776) );
  inv_x1_sg U74037 ( .A(\reg_yHat[0][9] ), .X(n46638) );
  nand_x1_sg U74038 ( .A(\reg_yHat[1][7] ), .B(n47183), .X(n23067) );
  inv_x1_sg U74039 ( .A(\reg_y[1][7] ), .X(n47183) );
  nand_x1_sg U74040 ( .A(\reg_y[1][7] ), .B(n46649), .X(n23070) );
  inv_x1_sg U74041 ( .A(\reg_yHat[1][7] ), .X(n46649) );
  nand_x1_sg U74042 ( .A(\reg_yHat[2][7] ), .B(n47468), .X(n23347) );
  inv_x1_sg U74043 ( .A(\reg_y[2][7] ), .X(n47468) );
  nand_x1_sg U74044 ( .A(\reg_y[2][7] ), .B(n46663), .X(n23350) );
  inv_x1_sg U74045 ( .A(\reg_yHat[2][7] ), .X(n46663) );
  nand_x1_sg U74046 ( .A(\reg_yHat[3][7] ), .B(n47753), .X(n23626) );
  inv_x1_sg U74047 ( .A(\reg_y[3][7] ), .X(n47753) );
  nand_x1_sg U74048 ( .A(\reg_y[3][7] ), .B(n46677), .X(n23629) );
  inv_x1_sg U74049 ( .A(\reg_yHat[3][7] ), .X(n46677) );
  nand_x1_sg U74050 ( .A(\reg_yHat[4][7] ), .B(n48038), .X(n23905) );
  inv_x1_sg U74051 ( .A(\reg_y[4][7] ), .X(n48038) );
  nand_x1_sg U74052 ( .A(\reg_y[4][7] ), .B(n46691), .X(n23908) );
  inv_x1_sg U74053 ( .A(\reg_yHat[4][7] ), .X(n46691) );
  nand_x1_sg U74054 ( .A(\reg_yHat[5][7] ), .B(n48323), .X(n24184) );
  inv_x1_sg U74055 ( .A(\reg_y[5][7] ), .X(n48323) );
  nand_x1_sg U74056 ( .A(\reg_y[5][7] ), .B(n46705), .X(n24187) );
  inv_x1_sg U74057 ( .A(\reg_yHat[5][7] ), .X(n46705) );
  nand_x1_sg U74058 ( .A(\reg_yHat[6][7] ), .B(n48608), .X(n24463) );
  inv_x1_sg U74059 ( .A(\reg_y[6][7] ), .X(n48608) );
  nand_x1_sg U74060 ( .A(\reg_y[6][7] ), .B(n46719), .X(n24466) );
  inv_x1_sg U74061 ( .A(\reg_yHat[6][7] ), .X(n46719) );
  nand_x1_sg U74062 ( .A(\reg_yHat[7][7] ), .B(n48894), .X(n24741) );
  inv_x1_sg U74063 ( .A(\reg_y[7][7] ), .X(n48894) );
  nand_x1_sg U74064 ( .A(\reg_y[7][7] ), .B(n46733), .X(n24744) );
  inv_x1_sg U74065 ( .A(\reg_yHat[7][7] ), .X(n46733) );
  nand_x1_sg U74066 ( .A(\reg_yHat[8][7] ), .B(n49181), .X(n25020) );
  inv_x1_sg U74067 ( .A(\reg_y[8][7] ), .X(n49181) );
  nand_x1_sg U74068 ( .A(\reg_y[8][7] ), .B(n46747), .X(n25023) );
  inv_x1_sg U74069 ( .A(\reg_yHat[8][7] ), .X(n46747) );
  nand_x1_sg U74070 ( .A(\reg_yHat[9][7] ), .B(n49467), .X(n25299) );
  inv_x1_sg U74071 ( .A(\reg_y[9][7] ), .X(n49467) );
  nand_x1_sg U74072 ( .A(\reg_y[9][7] ), .B(n46761), .X(n25302) );
  inv_x1_sg U74073 ( .A(\reg_yHat[9][7] ), .X(n46761) );
  nand_x1_sg U74074 ( .A(\reg_yHat[10][7] ), .B(n49752), .X(n25578) );
  inv_x1_sg U74075 ( .A(\reg_y[10][7] ), .X(n49752) );
  nand_x1_sg U74076 ( .A(\reg_y[10][7] ), .B(n46775), .X(n25581) );
  inv_x1_sg U74077 ( .A(\reg_yHat[10][7] ), .X(n46775) );
  nand_x1_sg U74078 ( .A(\reg_yHat[11][7] ), .B(n50039), .X(n25855) );
  inv_x1_sg U74079 ( .A(\reg_y[11][7] ), .X(n50039) );
  nand_x1_sg U74080 ( .A(\reg_y[11][7] ), .B(n46789), .X(n25858) );
  inv_x1_sg U74081 ( .A(\reg_yHat[11][7] ), .X(n46789) );
  nand_x1_sg U74082 ( .A(\reg_yHat[13][7] ), .B(n50613), .X(n26415) );
  inv_x1_sg U74083 ( .A(\reg_y[13][7] ), .X(n50613) );
  nand_x1_sg U74084 ( .A(\reg_y[13][7] ), .B(n46816), .X(n26418) );
  inv_x1_sg U74085 ( .A(\reg_yHat[13][7] ), .X(n46816) );
  nand_x1_sg U74086 ( .A(\reg_yHat[14][7] ), .B(n50900), .X(n26693) );
  inv_x1_sg U74087 ( .A(\reg_y[14][7] ), .X(n50900) );
  nand_x1_sg U74088 ( .A(\reg_y[14][7] ), .B(n46830), .X(n26696) );
  inv_x1_sg U74089 ( .A(\reg_yHat[14][7] ), .X(n46830) );
  nand_x1_sg U74090 ( .A(\reg_yHat[12][11] ), .B(n50396), .X(n26067) );
  inv_x1_sg U74091 ( .A(\reg_y[12][11] ), .X(n50396) );
  nand_x1_sg U74092 ( .A(\reg_yHat[12][12] ), .B(n50414), .X(n26062) );
  inv_x1_sg U74093 ( .A(\reg_y[12][12] ), .X(n50414) );
  nand_x1_sg U74094 ( .A(\reg_y[12][12] ), .B(n46808), .X(n26061) );
  inv_x1_sg U74095 ( .A(\reg_yHat[12][12] ), .X(n46808) );
  nand_x1_sg U74096 ( .A(\reg_y[12][11] ), .B(n46807), .X(n26068) );
  inv_x1_sg U74097 ( .A(\reg_yHat[12][11] ), .X(n46807) );
  nand_x1_sg U74098 ( .A(\reg_y[12][7] ), .B(n46803), .X(n26091) );
  inv_x1_sg U74099 ( .A(\reg_yHat[12][7] ), .X(n46803) );
  nand_x1_sg U74100 ( .A(\reg_yHat[1][8] ), .B(n47195), .X(n23060) );
  inv_x1_sg U74101 ( .A(\reg_y[1][8] ), .X(n47195) );
  nand_x1_sg U74102 ( .A(\reg_y[1][8] ), .B(n46650), .X(n23062) );
  inv_x1_sg U74103 ( .A(\reg_yHat[1][8] ), .X(n46650) );
  nand_x1_sg U74104 ( .A(\reg_yHat[2][8] ), .B(n47480), .X(n23340) );
  inv_x1_sg U74105 ( .A(\reg_y[2][8] ), .X(n47480) );
  nand_x1_sg U74106 ( .A(\reg_y[2][8] ), .B(n46664), .X(n23342) );
  inv_x1_sg U74107 ( .A(\reg_yHat[2][8] ), .X(n46664) );
  nand_x1_sg U74108 ( .A(\reg_yHat[3][8] ), .B(n47765), .X(n23619) );
  inv_x1_sg U74109 ( .A(\reg_y[3][8] ), .X(n47765) );
  nand_x1_sg U74110 ( .A(\reg_y[3][8] ), .B(n46678), .X(n23621) );
  inv_x1_sg U74111 ( .A(\reg_yHat[3][8] ), .X(n46678) );
  nand_x1_sg U74112 ( .A(\reg_yHat[4][8] ), .B(n48050), .X(n23898) );
  inv_x1_sg U74113 ( .A(\reg_y[4][8] ), .X(n48050) );
  nand_x1_sg U74114 ( .A(\reg_y[4][8] ), .B(n46692), .X(n23900) );
  inv_x1_sg U74115 ( .A(\reg_yHat[4][8] ), .X(n46692) );
  nand_x1_sg U74116 ( .A(\reg_yHat[5][8] ), .B(n48335), .X(n24177) );
  inv_x1_sg U74117 ( .A(\reg_y[5][8] ), .X(n48335) );
  nand_x1_sg U74118 ( .A(\reg_y[5][8] ), .B(n46706), .X(n24179) );
  inv_x1_sg U74119 ( .A(\reg_yHat[5][8] ), .X(n46706) );
  nand_x1_sg U74120 ( .A(\reg_yHat[6][8] ), .B(n48620), .X(n24456) );
  inv_x1_sg U74121 ( .A(\reg_y[6][8] ), .X(n48620) );
  nand_x1_sg U74122 ( .A(\reg_y[6][8] ), .B(n46720), .X(n24458) );
  inv_x1_sg U74123 ( .A(\reg_yHat[6][8] ), .X(n46720) );
  nand_x1_sg U74124 ( .A(\reg_yHat[7][8] ), .B(n48906), .X(n24734) );
  inv_x1_sg U74125 ( .A(\reg_y[7][8] ), .X(n48906) );
  nand_x1_sg U74126 ( .A(\reg_y[7][8] ), .B(n46734), .X(n24736) );
  inv_x1_sg U74127 ( .A(\reg_yHat[7][8] ), .X(n46734) );
  nand_x1_sg U74128 ( .A(\reg_yHat[8][8] ), .B(n49193), .X(n25013) );
  inv_x1_sg U74129 ( .A(\reg_y[8][8] ), .X(n49193) );
  nand_x1_sg U74130 ( .A(\reg_y[8][8] ), .B(n46748), .X(n25015) );
  inv_x1_sg U74131 ( .A(\reg_yHat[8][8] ), .X(n46748) );
  nand_x1_sg U74132 ( .A(\reg_yHat[9][8] ), .B(n49479), .X(n25292) );
  inv_x1_sg U74133 ( .A(\reg_y[9][8] ), .X(n49479) );
  nand_x1_sg U74134 ( .A(\reg_y[9][8] ), .B(n46762), .X(n25294) );
  inv_x1_sg U74135 ( .A(\reg_yHat[9][8] ), .X(n46762) );
  nand_x1_sg U74136 ( .A(\reg_yHat[10][8] ), .B(n49765), .X(n25571) );
  inv_x1_sg U74137 ( .A(\reg_y[10][8] ), .X(n49765) );
  nand_x1_sg U74138 ( .A(\reg_y[10][8] ), .B(n46776), .X(n25573) );
  inv_x1_sg U74139 ( .A(\reg_yHat[10][8] ), .X(n46776) );
  nand_x1_sg U74140 ( .A(\reg_yHat[11][8] ), .B(n50051), .X(n25848) );
  inv_x1_sg U74141 ( .A(\reg_y[11][8] ), .X(n50051) );
  nand_x1_sg U74142 ( .A(\reg_y[11][8] ), .B(n46790), .X(n25850) );
  inv_x1_sg U74143 ( .A(\reg_yHat[11][8] ), .X(n46790) );
  nand_x1_sg U74144 ( .A(\reg_yHat[12][7] ), .B(n50324), .X(n26092) );
  inv_x1_sg U74145 ( .A(\reg_y[12][7] ), .X(n50324) );
  nand_x1_sg U74146 ( .A(\reg_yHat[12][8] ), .B(n50337), .X(n26086) );
  inv_x1_sg U74147 ( .A(\reg_y[12][8] ), .X(n50337) );
  nand_x1_sg U74148 ( .A(\reg_y[12][8] ), .B(n46804), .X(n26085) );
  inv_x1_sg U74149 ( .A(\reg_yHat[12][8] ), .X(n46804) );
  nand_x1_sg U74150 ( .A(\reg_yHat[13][8] ), .B(n50625), .X(n26408) );
  inv_x1_sg U74151 ( .A(\reg_y[13][8] ), .X(n50625) );
  nand_x1_sg U74152 ( .A(\reg_y[13][8] ), .B(n46817), .X(n26410) );
  inv_x1_sg U74153 ( .A(\reg_yHat[13][8] ), .X(n46817) );
  nand_x1_sg U74154 ( .A(\reg_yHat[14][8] ), .B(n50912), .X(n26686) );
  inv_x1_sg U74155 ( .A(\reg_y[14][8] ), .X(n50912) );
  nand_x1_sg U74156 ( .A(\reg_y[14][8] ), .B(n46831), .X(n26688) );
  inv_x1_sg U74157 ( .A(\reg_yHat[14][8] ), .X(n46831) );
  nand_x1_sg U74158 ( .A(\reg_yHat[12][9] ), .B(n50357), .X(n26079) );
  inv_x1_sg U74159 ( .A(\reg_y[12][9] ), .X(n50357) );
  nand_x1_sg U74160 ( .A(\reg_yHat[0][7] ), .B(n46890), .X(n22790) );
  inv_x1_sg U74161 ( .A(\reg_y[0][7] ), .X(n46890) );
  nand_x1_sg U74162 ( .A(\reg_y[0][7] ), .B(n46636), .X(n22793) );
  inv_x1_sg U74163 ( .A(\reg_yHat[0][7] ), .X(n46636) );
  nand_x1_sg U74164 ( .A(\reg_y[0][8] ), .B(n46637), .X(n22785) );
  inv_x1_sg U74165 ( .A(\reg_yHat[0][8] ), .X(n46637) );
  nand_x1_sg U74166 ( .A(\reg_yHat[12][10] ), .B(n50374), .X(n26074) );
  inv_x1_sg U74167 ( .A(\reg_y[12][10] ), .X(n50374) );
  nand_x1_sg U74168 ( .A(\reg_y[12][9] ), .B(n46805), .X(n26080) );
  inv_x1_sg U74169 ( .A(\reg_yHat[12][9] ), .X(n46805) );
  nand_x1_sg U74170 ( .A(\reg_y[12][10] ), .B(n46806), .X(n26073) );
  inv_x1_sg U74171 ( .A(\reg_yHat[12][10] ), .X(n46806) );
  nand_x1_sg U74172 ( .A(\reg_yHat[0][8] ), .B(n46902), .X(n22783) );
  inv_x1_sg U74173 ( .A(\reg_y[0][8] ), .X(n46902) );
  nand_x1_sg U74174 ( .A(\reg_yHat[0][11] ), .B(n46964), .X(n22764) );
  inv_x1_sg U74175 ( .A(\reg_y[0][11] ), .X(n46964) );
  nand_x1_sg U74176 ( .A(\reg_y[0][12] ), .B(n46641), .X(n22757) );
  inv_x1_sg U74177 ( .A(\reg_yHat[0][12] ), .X(n46641) );
  nand_x1_sg U74178 ( .A(\reg_y[0][11] ), .B(n46640), .X(n22762) );
  inv_x1_sg U74179 ( .A(\reg_yHat[0][11] ), .X(n46640) );
  nand_x1_sg U74180 ( .A(\reg_yHat[0][12] ), .B(n46983), .X(n22755) );
  inv_x1_sg U74181 ( .A(\reg_y[0][12] ), .X(n46983) );
  nand_x1_sg U74182 ( .A(\reg_yHat[0][13] ), .B(n47006), .X(n22750) );
  inv_x1_sg U74183 ( .A(\reg_y[0][13] ), .X(n47006) );
  nand_x1_sg U74184 ( .A(\reg_y[0][14] ), .B(n46643), .X(n22743) );
  inv_x1_sg U74185 ( .A(\reg_yHat[0][14] ), .X(n46643) );
  nand_x1_sg U74186 ( .A(\reg_y[0][13] ), .B(n46642), .X(n22748) );
  inv_x1_sg U74187 ( .A(\reg_yHat[0][13] ), .X(n46642) );
  nand_x1_sg U74188 ( .A(\reg_yHat[0][14] ), .B(n47025), .X(n22741) );
  inv_x1_sg U74189 ( .A(\reg_y[0][14] ), .X(n47025) );
  nand_x1_sg U74190 ( .A(\reg_y[0][15] ), .B(n46644), .X(n22734) );
  inv_x1_sg U74191 ( .A(\reg_yHat[0][15] ), .X(n46644) );
  nand_x1_sg U74192 ( .A(\reg_yHat[0][15] ), .B(n47055), .X(n22736) );
  inv_x1_sg U74193 ( .A(\reg_y[0][15] ), .X(n47055) );
  nand_x1_sg U74194 ( .A(\reg_yHat[1][9] ), .B(n47215), .X(n23055) );
  inv_x1_sg U74195 ( .A(\reg_y[1][9] ), .X(n47215) );
  nand_x1_sg U74196 ( .A(\reg_y[1][10] ), .B(n46652), .X(n23048) );
  inv_x1_sg U74197 ( .A(\reg_yHat[1][10] ), .X(n46652) );
  nand_x1_sg U74198 ( .A(\reg_y[1][9] ), .B(n46651), .X(n23053) );
  inv_x1_sg U74199 ( .A(\reg_yHat[1][9] ), .X(n46651) );
  nand_x1_sg U74200 ( .A(\reg_yHat[1][10] ), .B(n47232), .X(n23046) );
  inv_x1_sg U74201 ( .A(\reg_y[1][10] ), .X(n47232) );
  nand_x1_sg U74202 ( .A(\reg_yHat[1][11] ), .B(n47254), .X(n23041) );
  inv_x1_sg U74203 ( .A(\reg_y[1][11] ), .X(n47254) );
  nand_x1_sg U74204 ( .A(\reg_y[1][12] ), .B(n46654), .X(n23034) );
  inv_x1_sg U74205 ( .A(\reg_yHat[1][12] ), .X(n46654) );
  nand_x1_sg U74206 ( .A(\reg_y[1][11] ), .B(n46653), .X(n23039) );
  inv_x1_sg U74207 ( .A(\reg_yHat[1][11] ), .X(n46653) );
  nand_x1_sg U74208 ( .A(\reg_yHat[1][12] ), .B(n47272), .X(n23032) );
  inv_x1_sg U74209 ( .A(\reg_y[1][12] ), .X(n47272) );
  nand_x1_sg U74210 ( .A(\reg_yHat[1][13] ), .B(n47294), .X(n23027) );
  inv_x1_sg U74211 ( .A(\reg_y[1][13] ), .X(n47294) );
  nand_x1_sg U74212 ( .A(\reg_y[1][14] ), .B(n46656), .X(n23020) );
  inv_x1_sg U74213 ( .A(\reg_yHat[1][14] ), .X(n46656) );
  nand_x1_sg U74214 ( .A(\reg_y[1][13] ), .B(n46655), .X(n23025) );
  inv_x1_sg U74215 ( .A(\reg_yHat[1][13] ), .X(n46655) );
  nand_x1_sg U74216 ( .A(\reg_yHat[1][14] ), .B(n47312), .X(n23018) );
  inv_x1_sg U74217 ( .A(\reg_y[1][14] ), .X(n47312) );
  nand_x1_sg U74218 ( .A(\reg_y[1][15] ), .B(n46657), .X(n23011) );
  inv_x1_sg U74219 ( .A(\reg_yHat[1][15] ), .X(n46657) );
  nand_x1_sg U74220 ( .A(\reg_yHat[1][15] ), .B(n47341), .X(n23013) );
  inv_x1_sg U74221 ( .A(\reg_y[1][15] ), .X(n47341) );
  nand_x1_sg U74222 ( .A(\reg_yHat[2][9] ), .B(n47500), .X(n23335) );
  inv_x1_sg U74223 ( .A(\reg_y[2][9] ), .X(n47500) );
  nand_x1_sg U74224 ( .A(\reg_y[2][10] ), .B(n46666), .X(n23328) );
  inv_x1_sg U74225 ( .A(\reg_yHat[2][10] ), .X(n46666) );
  nand_x1_sg U74226 ( .A(\reg_y[2][9] ), .B(n46665), .X(n23333) );
  inv_x1_sg U74227 ( .A(\reg_yHat[2][9] ), .X(n46665) );
  nand_x1_sg U74228 ( .A(\reg_yHat[2][10] ), .B(n47517), .X(n23326) );
  inv_x1_sg U74229 ( .A(\reg_y[2][10] ), .X(n47517) );
  nand_x1_sg U74230 ( .A(\reg_yHat[2][11] ), .B(n47539), .X(n23321) );
  inv_x1_sg U74231 ( .A(\reg_y[2][11] ), .X(n47539) );
  nand_x1_sg U74232 ( .A(\reg_y[2][12] ), .B(n46668), .X(n23314) );
  inv_x1_sg U74233 ( .A(\reg_yHat[2][12] ), .X(n46668) );
  nand_x1_sg U74234 ( .A(\reg_y[2][11] ), .B(n46667), .X(n23319) );
  inv_x1_sg U74235 ( .A(\reg_yHat[2][11] ), .X(n46667) );
  nand_x1_sg U74236 ( .A(\reg_yHat[2][12] ), .B(n47557), .X(n23312) );
  inv_x1_sg U74237 ( .A(\reg_y[2][12] ), .X(n47557) );
  nand_x1_sg U74238 ( .A(\reg_yHat[2][13] ), .B(n47579), .X(n23307) );
  inv_x1_sg U74239 ( .A(\reg_y[2][13] ), .X(n47579) );
  nand_x1_sg U74240 ( .A(\reg_y[2][14] ), .B(n46670), .X(n23300) );
  inv_x1_sg U74241 ( .A(\reg_yHat[2][14] ), .X(n46670) );
  nand_x1_sg U74242 ( .A(\reg_y[2][13] ), .B(n46669), .X(n23305) );
  inv_x1_sg U74243 ( .A(\reg_yHat[2][13] ), .X(n46669) );
  nand_x1_sg U74244 ( .A(\reg_yHat[2][14] ), .B(n47597), .X(n23298) );
  inv_x1_sg U74245 ( .A(\reg_y[2][14] ), .X(n47597) );
  nand_x1_sg U74246 ( .A(\reg_y[2][15] ), .B(n46671), .X(n23291) );
  inv_x1_sg U74247 ( .A(\reg_yHat[2][15] ), .X(n46671) );
  nand_x1_sg U74248 ( .A(\reg_yHat[2][15] ), .B(n47626), .X(n23293) );
  inv_x1_sg U74249 ( .A(\reg_y[2][15] ), .X(n47626) );
  nand_x1_sg U74250 ( .A(\reg_yHat[3][9] ), .B(n47785), .X(n23614) );
  inv_x1_sg U74251 ( .A(\reg_y[3][9] ), .X(n47785) );
  nand_x1_sg U74252 ( .A(\reg_y[3][10] ), .B(n46680), .X(n23607) );
  inv_x1_sg U74253 ( .A(\reg_yHat[3][10] ), .X(n46680) );
  nand_x1_sg U74254 ( .A(\reg_y[3][9] ), .B(n46679), .X(n23612) );
  inv_x1_sg U74255 ( .A(\reg_yHat[3][9] ), .X(n46679) );
  nand_x1_sg U74256 ( .A(\reg_yHat[3][10] ), .B(n47802), .X(n23605) );
  inv_x1_sg U74257 ( .A(\reg_y[3][10] ), .X(n47802) );
  nand_x1_sg U74258 ( .A(\reg_yHat[3][11] ), .B(n47824), .X(n23600) );
  inv_x1_sg U74259 ( .A(\reg_y[3][11] ), .X(n47824) );
  nand_x1_sg U74260 ( .A(\reg_y[3][12] ), .B(n46682), .X(n23593) );
  inv_x1_sg U74261 ( .A(\reg_yHat[3][12] ), .X(n46682) );
  nand_x1_sg U74262 ( .A(\reg_y[3][11] ), .B(n46681), .X(n23598) );
  inv_x1_sg U74263 ( .A(\reg_yHat[3][11] ), .X(n46681) );
  nand_x1_sg U74264 ( .A(\reg_yHat[3][12] ), .B(n47842), .X(n23591) );
  inv_x1_sg U74265 ( .A(\reg_y[3][12] ), .X(n47842) );
  nand_x1_sg U74266 ( .A(\reg_yHat[3][13] ), .B(n47864), .X(n23586) );
  inv_x1_sg U74267 ( .A(\reg_y[3][13] ), .X(n47864) );
  nand_x1_sg U74268 ( .A(\reg_y[3][14] ), .B(n46684), .X(n23579) );
  inv_x1_sg U74269 ( .A(\reg_yHat[3][14] ), .X(n46684) );
  nand_x1_sg U74270 ( .A(\reg_y[3][13] ), .B(n46683), .X(n23584) );
  inv_x1_sg U74271 ( .A(\reg_yHat[3][13] ), .X(n46683) );
  nand_x1_sg U74272 ( .A(\reg_yHat[3][14] ), .B(n47882), .X(n23577) );
  inv_x1_sg U74273 ( .A(\reg_y[3][14] ), .X(n47882) );
  nand_x1_sg U74274 ( .A(\reg_y[3][15] ), .B(n46685), .X(n23570) );
  inv_x1_sg U74275 ( .A(\reg_yHat[3][15] ), .X(n46685) );
  nand_x1_sg U74276 ( .A(\reg_yHat[3][15] ), .B(n47911), .X(n23572) );
  inv_x1_sg U74277 ( .A(\reg_y[3][15] ), .X(n47911) );
  nand_x1_sg U74278 ( .A(\reg_yHat[4][9] ), .B(n48070), .X(n23893) );
  inv_x1_sg U74279 ( .A(\reg_y[4][9] ), .X(n48070) );
  nand_x1_sg U74280 ( .A(\reg_y[4][10] ), .B(n46694), .X(n23886) );
  inv_x1_sg U74281 ( .A(\reg_yHat[4][10] ), .X(n46694) );
  nand_x1_sg U74282 ( .A(\reg_y[4][9] ), .B(n46693), .X(n23891) );
  inv_x1_sg U74283 ( .A(\reg_yHat[4][9] ), .X(n46693) );
  nand_x1_sg U74284 ( .A(\reg_yHat[4][10] ), .B(n48087), .X(n23884) );
  inv_x1_sg U74285 ( .A(\reg_y[4][10] ), .X(n48087) );
  nand_x1_sg U74286 ( .A(\reg_yHat[4][11] ), .B(n48109), .X(n23879) );
  inv_x1_sg U74287 ( .A(\reg_y[4][11] ), .X(n48109) );
  nand_x1_sg U74288 ( .A(\reg_y[4][12] ), .B(n46696), .X(n23872) );
  inv_x1_sg U74289 ( .A(\reg_yHat[4][12] ), .X(n46696) );
  nand_x1_sg U74290 ( .A(\reg_y[4][11] ), .B(n46695), .X(n23877) );
  inv_x1_sg U74291 ( .A(\reg_yHat[4][11] ), .X(n46695) );
  nand_x1_sg U74292 ( .A(\reg_yHat[4][12] ), .B(n48127), .X(n23870) );
  inv_x1_sg U74293 ( .A(\reg_y[4][12] ), .X(n48127) );
  nand_x1_sg U74294 ( .A(\reg_yHat[4][13] ), .B(n48149), .X(n23865) );
  inv_x1_sg U74295 ( .A(\reg_y[4][13] ), .X(n48149) );
  nand_x1_sg U74296 ( .A(\reg_y[4][14] ), .B(n46698), .X(n23858) );
  inv_x1_sg U74297 ( .A(\reg_yHat[4][14] ), .X(n46698) );
  nand_x1_sg U74298 ( .A(\reg_y[4][13] ), .B(n46697), .X(n23863) );
  inv_x1_sg U74299 ( .A(\reg_yHat[4][13] ), .X(n46697) );
  nand_x1_sg U74300 ( .A(\reg_yHat[4][14] ), .B(n48167), .X(n23856) );
  inv_x1_sg U74301 ( .A(\reg_y[4][14] ), .X(n48167) );
  nand_x1_sg U74302 ( .A(\reg_y[4][15] ), .B(n46699), .X(n23849) );
  inv_x1_sg U74303 ( .A(\reg_yHat[4][15] ), .X(n46699) );
  nand_x1_sg U74304 ( .A(\reg_yHat[4][15] ), .B(n48196), .X(n23851) );
  inv_x1_sg U74305 ( .A(\reg_y[4][15] ), .X(n48196) );
  nand_x1_sg U74306 ( .A(\reg_yHat[5][9] ), .B(n48355), .X(n24172) );
  inv_x1_sg U74307 ( .A(\reg_y[5][9] ), .X(n48355) );
  nand_x1_sg U74308 ( .A(\reg_y[5][10] ), .B(n46708), .X(n24165) );
  inv_x1_sg U74309 ( .A(\reg_yHat[5][10] ), .X(n46708) );
  nand_x1_sg U74310 ( .A(\reg_y[5][9] ), .B(n46707), .X(n24170) );
  inv_x1_sg U74311 ( .A(\reg_yHat[5][9] ), .X(n46707) );
  nand_x1_sg U74312 ( .A(\reg_yHat[5][10] ), .B(n48372), .X(n24163) );
  inv_x1_sg U74313 ( .A(\reg_y[5][10] ), .X(n48372) );
  nand_x1_sg U74314 ( .A(\reg_yHat[5][11] ), .B(n48394), .X(n24158) );
  inv_x1_sg U74315 ( .A(\reg_y[5][11] ), .X(n48394) );
  nand_x1_sg U74316 ( .A(\reg_y[5][12] ), .B(n46710), .X(n24151) );
  inv_x1_sg U74317 ( .A(\reg_yHat[5][12] ), .X(n46710) );
  nand_x1_sg U74318 ( .A(\reg_y[5][11] ), .B(n46709), .X(n24156) );
  inv_x1_sg U74319 ( .A(\reg_yHat[5][11] ), .X(n46709) );
  nand_x1_sg U74320 ( .A(\reg_yHat[5][12] ), .B(n48412), .X(n24149) );
  inv_x1_sg U74321 ( .A(\reg_y[5][12] ), .X(n48412) );
  nand_x1_sg U74322 ( .A(\reg_yHat[5][13] ), .B(n48434), .X(n24144) );
  inv_x1_sg U74323 ( .A(\reg_y[5][13] ), .X(n48434) );
  nand_x1_sg U74324 ( .A(\reg_y[5][14] ), .B(n46712), .X(n24137) );
  inv_x1_sg U74325 ( .A(\reg_yHat[5][14] ), .X(n46712) );
  nand_x1_sg U74326 ( .A(\reg_y[5][13] ), .B(n46711), .X(n24142) );
  inv_x1_sg U74327 ( .A(\reg_yHat[5][13] ), .X(n46711) );
  nand_x1_sg U74328 ( .A(\reg_yHat[5][14] ), .B(n48452), .X(n24135) );
  inv_x1_sg U74329 ( .A(\reg_y[5][14] ), .X(n48452) );
  nand_x1_sg U74330 ( .A(\reg_y[5][15] ), .B(n46713), .X(n24128) );
  inv_x1_sg U74331 ( .A(\reg_yHat[5][15] ), .X(n46713) );
  nand_x1_sg U74332 ( .A(\reg_yHat[5][15] ), .B(n48481), .X(n24130) );
  inv_x1_sg U74333 ( .A(\reg_y[5][15] ), .X(n48481) );
  nand_x1_sg U74334 ( .A(\reg_yHat[6][9] ), .B(n48640), .X(n24451) );
  inv_x1_sg U74335 ( .A(\reg_y[6][9] ), .X(n48640) );
  nand_x1_sg U74336 ( .A(\reg_y[6][10] ), .B(n46722), .X(n24444) );
  inv_x1_sg U74337 ( .A(\reg_yHat[6][10] ), .X(n46722) );
  nand_x1_sg U74338 ( .A(\reg_y[6][9] ), .B(n46721), .X(n24449) );
  inv_x1_sg U74339 ( .A(\reg_yHat[6][9] ), .X(n46721) );
  nand_x1_sg U74340 ( .A(\reg_yHat[6][10] ), .B(n48657), .X(n24442) );
  inv_x1_sg U74341 ( .A(\reg_y[6][10] ), .X(n48657) );
  nand_x1_sg U74342 ( .A(\reg_yHat[6][11] ), .B(n48679), .X(n24437) );
  inv_x1_sg U74343 ( .A(\reg_y[6][11] ), .X(n48679) );
  nand_x1_sg U74344 ( .A(\reg_y[6][12] ), .B(n46724), .X(n24430) );
  inv_x1_sg U74345 ( .A(\reg_yHat[6][12] ), .X(n46724) );
  nand_x1_sg U74346 ( .A(\reg_y[6][11] ), .B(n46723), .X(n24435) );
  inv_x1_sg U74347 ( .A(\reg_yHat[6][11] ), .X(n46723) );
  nand_x1_sg U74348 ( .A(\reg_yHat[6][12] ), .B(n48697), .X(n24428) );
  inv_x1_sg U74349 ( .A(\reg_y[6][12] ), .X(n48697) );
  nand_x1_sg U74350 ( .A(\reg_yHat[6][13] ), .B(n48719), .X(n24423) );
  inv_x1_sg U74351 ( .A(\reg_y[6][13] ), .X(n48719) );
  nand_x1_sg U74352 ( .A(\reg_y[6][14] ), .B(n46726), .X(n24416) );
  inv_x1_sg U74353 ( .A(\reg_yHat[6][14] ), .X(n46726) );
  nand_x1_sg U74354 ( .A(\reg_y[6][13] ), .B(n46725), .X(n24421) );
  inv_x1_sg U74355 ( .A(\reg_yHat[6][13] ), .X(n46725) );
  nand_x1_sg U74356 ( .A(\reg_yHat[6][14] ), .B(n48737), .X(n24414) );
  inv_x1_sg U74357 ( .A(\reg_y[6][14] ), .X(n48737) );
  nand_x1_sg U74358 ( .A(\reg_y[6][15] ), .B(n46727), .X(n24407) );
  inv_x1_sg U74359 ( .A(\reg_yHat[6][15] ), .X(n46727) );
  nand_x1_sg U74360 ( .A(\reg_yHat[6][15] ), .B(n48766), .X(n24409) );
  inv_x1_sg U74361 ( .A(\reg_y[6][15] ), .X(n48766) );
  nand_x1_sg U74362 ( .A(\reg_yHat[7][9] ), .B(n48926), .X(n24729) );
  inv_x1_sg U74363 ( .A(\reg_y[7][9] ), .X(n48926) );
  nand_x1_sg U74364 ( .A(\reg_y[7][10] ), .B(n46736), .X(n24722) );
  inv_x1_sg U74365 ( .A(\reg_yHat[7][10] ), .X(n46736) );
  nand_x1_sg U74366 ( .A(\reg_y[7][9] ), .B(n46735), .X(n24727) );
  inv_x1_sg U74367 ( .A(\reg_yHat[7][9] ), .X(n46735) );
  nand_x1_sg U74368 ( .A(\reg_yHat[7][10] ), .B(n48943), .X(n24720) );
  inv_x1_sg U74369 ( .A(\reg_y[7][10] ), .X(n48943) );
  nand_x1_sg U74370 ( .A(\reg_yHat[7][11] ), .B(n48965), .X(n24715) );
  inv_x1_sg U74371 ( .A(\reg_y[7][11] ), .X(n48965) );
  nand_x1_sg U74372 ( .A(\reg_y[7][12] ), .B(n46738), .X(n24708) );
  inv_x1_sg U74373 ( .A(\reg_yHat[7][12] ), .X(n46738) );
  nand_x1_sg U74374 ( .A(\reg_y[7][11] ), .B(n46737), .X(n24713) );
  inv_x1_sg U74375 ( .A(\reg_yHat[7][11] ), .X(n46737) );
  nand_x1_sg U74376 ( .A(\reg_yHat[7][12] ), .B(n48983), .X(n24706) );
  inv_x1_sg U74377 ( .A(\reg_y[7][12] ), .X(n48983) );
  nand_x1_sg U74378 ( .A(\reg_yHat[7][13] ), .B(n49005), .X(n24701) );
  inv_x1_sg U74379 ( .A(\reg_y[7][13] ), .X(n49005) );
  nand_x1_sg U74380 ( .A(\reg_y[7][14] ), .B(n46740), .X(n24694) );
  inv_x1_sg U74381 ( .A(\reg_yHat[7][14] ), .X(n46740) );
  nand_x1_sg U74382 ( .A(\reg_y[7][13] ), .B(n46739), .X(n24699) );
  inv_x1_sg U74383 ( .A(\reg_yHat[7][13] ), .X(n46739) );
  nand_x1_sg U74384 ( .A(\reg_yHat[7][14] ), .B(n49023), .X(n24692) );
  inv_x1_sg U74385 ( .A(\reg_y[7][14] ), .X(n49023) );
  nand_x1_sg U74386 ( .A(\reg_y[7][15] ), .B(n46741), .X(n24685) );
  inv_x1_sg U74387 ( .A(\reg_yHat[7][15] ), .X(n46741) );
  nand_x1_sg U74388 ( .A(\reg_yHat[7][15] ), .B(n49052), .X(n24687) );
  inv_x1_sg U74389 ( .A(\reg_y[7][15] ), .X(n49052) );
  nand_x1_sg U74390 ( .A(\reg_yHat[8][9] ), .B(n49213), .X(n25008) );
  inv_x1_sg U74391 ( .A(\reg_y[8][9] ), .X(n49213) );
  nand_x1_sg U74392 ( .A(\reg_y[8][10] ), .B(n46750), .X(n25001) );
  inv_x1_sg U74393 ( .A(\reg_yHat[8][10] ), .X(n46750) );
  nand_x1_sg U74394 ( .A(\reg_y[8][9] ), .B(n46749), .X(n25006) );
  inv_x1_sg U74395 ( .A(\reg_yHat[8][9] ), .X(n46749) );
  nand_x1_sg U74396 ( .A(\reg_yHat[8][10] ), .B(n49230), .X(n24999) );
  inv_x1_sg U74397 ( .A(\reg_y[8][10] ), .X(n49230) );
  nand_x1_sg U74398 ( .A(\reg_yHat[8][11] ), .B(n49252), .X(n24994) );
  inv_x1_sg U74399 ( .A(\reg_y[8][11] ), .X(n49252) );
  nand_x1_sg U74400 ( .A(\reg_y[8][12] ), .B(n46752), .X(n24987) );
  inv_x1_sg U74401 ( .A(\reg_yHat[8][12] ), .X(n46752) );
  nand_x1_sg U74402 ( .A(\reg_y[8][11] ), .B(n46751), .X(n24992) );
  inv_x1_sg U74403 ( .A(\reg_yHat[8][11] ), .X(n46751) );
  nand_x1_sg U74404 ( .A(\reg_yHat[8][12] ), .B(n49270), .X(n24985) );
  inv_x1_sg U74405 ( .A(\reg_y[8][12] ), .X(n49270) );
  nand_x1_sg U74406 ( .A(\reg_yHat[8][13] ), .B(n49292), .X(n24980) );
  inv_x1_sg U74407 ( .A(\reg_y[8][13] ), .X(n49292) );
  nand_x1_sg U74408 ( .A(\reg_y[8][14] ), .B(n46754), .X(n24973) );
  inv_x1_sg U74409 ( .A(\reg_yHat[8][14] ), .X(n46754) );
  nand_x1_sg U74410 ( .A(\reg_y[8][13] ), .B(n46753), .X(n24978) );
  inv_x1_sg U74411 ( .A(\reg_yHat[8][13] ), .X(n46753) );
  nand_x1_sg U74412 ( .A(\reg_yHat[8][14] ), .B(n49310), .X(n24971) );
  inv_x1_sg U74413 ( .A(\reg_y[8][14] ), .X(n49310) );
  nand_x1_sg U74414 ( .A(\reg_y[8][15] ), .B(n46755), .X(n24964) );
  inv_x1_sg U74415 ( .A(\reg_yHat[8][15] ), .X(n46755) );
  nand_x1_sg U74416 ( .A(\reg_yHat[8][15] ), .B(n49339), .X(n24966) );
  inv_x1_sg U74417 ( .A(\reg_y[8][15] ), .X(n49339) );
  nand_x1_sg U74418 ( .A(\reg_yHat[9][9] ), .B(n49499), .X(n25287) );
  inv_x1_sg U74419 ( .A(\reg_y[9][9] ), .X(n49499) );
  nand_x1_sg U74420 ( .A(\reg_y[9][10] ), .B(n46764), .X(n25280) );
  inv_x1_sg U74421 ( .A(\reg_yHat[9][10] ), .X(n46764) );
  nand_x1_sg U74422 ( .A(\reg_y[9][9] ), .B(n46763), .X(n25285) );
  inv_x1_sg U74423 ( .A(\reg_yHat[9][9] ), .X(n46763) );
  nand_x1_sg U74424 ( .A(\reg_yHat[9][10] ), .B(n49516), .X(n25278) );
  inv_x1_sg U74425 ( .A(\reg_y[9][10] ), .X(n49516) );
  nand_x1_sg U74426 ( .A(\reg_yHat[9][11] ), .B(n49538), .X(n25273) );
  inv_x1_sg U74427 ( .A(\reg_y[9][11] ), .X(n49538) );
  nand_x1_sg U74428 ( .A(\reg_y[9][12] ), .B(n46766), .X(n25266) );
  inv_x1_sg U74429 ( .A(\reg_yHat[9][12] ), .X(n46766) );
  nand_x1_sg U74430 ( .A(\reg_y[9][11] ), .B(n46765), .X(n25271) );
  inv_x1_sg U74431 ( .A(\reg_yHat[9][11] ), .X(n46765) );
  nand_x1_sg U74432 ( .A(\reg_yHat[9][12] ), .B(n49556), .X(n25264) );
  inv_x1_sg U74433 ( .A(\reg_y[9][12] ), .X(n49556) );
  nand_x1_sg U74434 ( .A(\reg_yHat[9][13] ), .B(n49578), .X(n25259) );
  inv_x1_sg U74435 ( .A(\reg_y[9][13] ), .X(n49578) );
  nand_x1_sg U74436 ( .A(\reg_y[9][14] ), .B(n46768), .X(n25252) );
  inv_x1_sg U74437 ( .A(\reg_yHat[9][14] ), .X(n46768) );
  nand_x1_sg U74438 ( .A(\reg_y[9][13] ), .B(n46767), .X(n25257) );
  inv_x1_sg U74439 ( .A(\reg_yHat[9][13] ), .X(n46767) );
  nand_x1_sg U74440 ( .A(\reg_yHat[9][14] ), .B(n49596), .X(n25250) );
  inv_x1_sg U74441 ( .A(\reg_y[9][14] ), .X(n49596) );
  nand_x1_sg U74442 ( .A(\reg_y[9][15] ), .B(n46769), .X(n25243) );
  inv_x1_sg U74443 ( .A(\reg_yHat[9][15] ), .X(n46769) );
  nand_x1_sg U74444 ( .A(\reg_yHat[9][15] ), .B(n49625), .X(n25245) );
  inv_x1_sg U74445 ( .A(\reg_y[9][15] ), .X(n49625) );
  nand_x1_sg U74446 ( .A(\reg_yHat[10][9] ), .B(n49785), .X(n25566) );
  inv_x1_sg U74447 ( .A(\reg_y[10][9] ), .X(n49785) );
  nand_x1_sg U74448 ( .A(\reg_y[10][10] ), .B(n46778), .X(n25559) );
  inv_x1_sg U74449 ( .A(\reg_yHat[10][10] ), .X(n46778) );
  nand_x1_sg U74450 ( .A(\reg_y[10][9] ), .B(n46777), .X(n25564) );
  inv_x1_sg U74451 ( .A(\reg_yHat[10][9] ), .X(n46777) );
  nand_x1_sg U74452 ( .A(\reg_yHat[10][10] ), .B(n49802), .X(n25557) );
  inv_x1_sg U74453 ( .A(\reg_y[10][10] ), .X(n49802) );
  nand_x1_sg U74454 ( .A(\reg_yHat[10][11] ), .B(n49824), .X(n25552) );
  inv_x1_sg U74455 ( .A(\reg_y[10][11] ), .X(n49824) );
  nand_x1_sg U74456 ( .A(\reg_y[10][12] ), .B(n46780), .X(n25545) );
  inv_x1_sg U74457 ( .A(\reg_yHat[10][12] ), .X(n46780) );
  nand_x1_sg U74458 ( .A(\reg_y[10][11] ), .B(n46779), .X(n25550) );
  inv_x1_sg U74459 ( .A(\reg_yHat[10][11] ), .X(n46779) );
  nand_x1_sg U74460 ( .A(\reg_yHat[10][12] ), .B(n49842), .X(n25543) );
  inv_x1_sg U74461 ( .A(\reg_y[10][12] ), .X(n49842) );
  nand_x1_sg U74462 ( .A(\reg_yHat[10][13] ), .B(n49864), .X(n25538) );
  inv_x1_sg U74463 ( .A(\reg_y[10][13] ), .X(n49864) );
  nand_x1_sg U74464 ( .A(\reg_y[10][14] ), .B(n46782), .X(n25531) );
  inv_x1_sg U74465 ( .A(\reg_yHat[10][14] ), .X(n46782) );
  nand_x1_sg U74466 ( .A(\reg_y[10][13] ), .B(n46781), .X(n25536) );
  inv_x1_sg U74467 ( .A(\reg_yHat[10][13] ), .X(n46781) );
  nand_x1_sg U74468 ( .A(\reg_yHat[10][14] ), .B(n49882), .X(n25529) );
  inv_x1_sg U74469 ( .A(\reg_y[10][14] ), .X(n49882) );
  nand_x1_sg U74470 ( .A(\reg_y[10][15] ), .B(n46783), .X(n25522) );
  inv_x1_sg U74471 ( .A(\reg_yHat[10][15] ), .X(n46783) );
  nand_x1_sg U74472 ( .A(\reg_yHat[10][15] ), .B(n49911), .X(n25524) );
  inv_x1_sg U74473 ( .A(\reg_y[10][15] ), .X(n49911) );
  nand_x1_sg U74474 ( .A(\reg_yHat[11][9] ), .B(n50071), .X(n25843) );
  inv_x1_sg U74475 ( .A(\reg_y[11][9] ), .X(n50071) );
  nand_x1_sg U74476 ( .A(\reg_y[11][10] ), .B(n46792), .X(n25836) );
  inv_x1_sg U74477 ( .A(\reg_yHat[11][10] ), .X(n46792) );
  nand_x1_sg U74478 ( .A(\reg_y[11][9] ), .B(n46791), .X(n25841) );
  inv_x1_sg U74479 ( .A(\reg_yHat[11][9] ), .X(n46791) );
  nand_x1_sg U74480 ( .A(\reg_yHat[11][10] ), .B(n50088), .X(n25834) );
  inv_x1_sg U74481 ( .A(\reg_y[11][10] ), .X(n50088) );
  nand_x1_sg U74482 ( .A(\reg_yHat[11][11] ), .B(n50110), .X(n25829) );
  inv_x1_sg U74483 ( .A(\reg_y[11][11] ), .X(n50110) );
  nand_x1_sg U74484 ( .A(\reg_y[11][12] ), .B(n46794), .X(n25822) );
  inv_x1_sg U74485 ( .A(\reg_yHat[11][12] ), .X(n46794) );
  nand_x1_sg U74486 ( .A(\reg_y[11][11] ), .B(n46793), .X(n25827) );
  inv_x1_sg U74487 ( .A(\reg_yHat[11][11] ), .X(n46793) );
  nand_x1_sg U74488 ( .A(\reg_yHat[11][12] ), .B(n50128), .X(n25820) );
  inv_x1_sg U74489 ( .A(\reg_y[11][12] ), .X(n50128) );
  nand_x1_sg U74490 ( .A(\reg_yHat[11][13] ), .B(n50150), .X(n25815) );
  inv_x1_sg U74491 ( .A(\reg_y[11][13] ), .X(n50150) );
  nand_x1_sg U74492 ( .A(\reg_y[11][14] ), .B(n46796), .X(n25808) );
  inv_x1_sg U74493 ( .A(\reg_yHat[11][14] ), .X(n46796) );
  nand_x1_sg U74494 ( .A(\reg_y[11][13] ), .B(n46795), .X(n25813) );
  inv_x1_sg U74495 ( .A(\reg_yHat[11][13] ), .X(n46795) );
  nand_x1_sg U74496 ( .A(\reg_yHat[11][14] ), .B(n50168), .X(n25806) );
  inv_x1_sg U74497 ( .A(\reg_y[11][14] ), .X(n50168) );
  nand_x1_sg U74498 ( .A(\reg_y[11][15] ), .B(n46797), .X(n25799) );
  inv_x1_sg U74499 ( .A(\reg_yHat[11][15] ), .X(n46797) );
  nand_x1_sg U74500 ( .A(\reg_yHat[11][15] ), .B(n50197), .X(n25801) );
  inv_x1_sg U74501 ( .A(\reg_y[11][15] ), .X(n50197) );
  nand_x1_sg U74502 ( .A(\reg_y[12][15] ), .B(n46811), .X(n26044) );
  inv_x1_sg U74503 ( .A(\reg_yHat[12][15] ), .X(n46811) );
  nand_x1_sg U74504 ( .A(\reg_yHat[12][15] ), .B(n50483), .X(n26043) );
  inv_x1_sg U74505 ( .A(\reg_y[12][15] ), .X(n50483) );
  nand_x1_sg U74506 ( .A(\reg_yHat[13][9] ), .B(n50645), .X(n26403) );
  inv_x1_sg U74507 ( .A(\reg_y[13][9] ), .X(n50645) );
  nand_x1_sg U74508 ( .A(\reg_y[13][10] ), .B(n46819), .X(n26396) );
  inv_x1_sg U74509 ( .A(\reg_yHat[13][10] ), .X(n46819) );
  nand_x1_sg U74510 ( .A(\reg_y[13][9] ), .B(n46818), .X(n26401) );
  inv_x1_sg U74511 ( .A(\reg_yHat[13][9] ), .X(n46818) );
  nand_x1_sg U74512 ( .A(\reg_yHat[13][10] ), .B(n50662), .X(n26394) );
  inv_x1_sg U74513 ( .A(\reg_y[13][10] ), .X(n50662) );
  nand_x1_sg U74514 ( .A(\reg_yHat[13][11] ), .B(n50684), .X(n26389) );
  inv_x1_sg U74515 ( .A(\reg_y[13][11] ), .X(n50684) );
  nand_x1_sg U74516 ( .A(\reg_y[13][12] ), .B(n46821), .X(n26382) );
  inv_x1_sg U74517 ( .A(\reg_yHat[13][12] ), .X(n46821) );
  nand_x1_sg U74518 ( .A(\reg_y[13][11] ), .B(n46820), .X(n26387) );
  inv_x1_sg U74519 ( .A(\reg_yHat[13][11] ), .X(n46820) );
  nand_x1_sg U74520 ( .A(\reg_yHat[13][12] ), .B(n50702), .X(n26380) );
  inv_x1_sg U74521 ( .A(\reg_y[13][12] ), .X(n50702) );
  nand_x1_sg U74522 ( .A(\reg_yHat[13][13] ), .B(n50724), .X(n26375) );
  inv_x1_sg U74523 ( .A(\reg_y[13][13] ), .X(n50724) );
  nand_x1_sg U74524 ( .A(\reg_y[13][14] ), .B(n46823), .X(n26368) );
  inv_x1_sg U74525 ( .A(\reg_yHat[13][14] ), .X(n46823) );
  nand_x1_sg U74526 ( .A(\reg_y[13][13] ), .B(n46822), .X(n26373) );
  inv_x1_sg U74527 ( .A(\reg_yHat[13][13] ), .X(n46822) );
  nand_x1_sg U74528 ( .A(\reg_yHat[13][14] ), .B(n50742), .X(n26366) );
  inv_x1_sg U74529 ( .A(\reg_y[13][14] ), .X(n50742) );
  nand_x1_sg U74530 ( .A(\reg_y[13][15] ), .B(n46824), .X(n26359) );
  inv_x1_sg U74531 ( .A(\reg_yHat[13][15] ), .X(n46824) );
  nand_x1_sg U74532 ( .A(\reg_yHat[13][15] ), .B(n50771), .X(n26361) );
  inv_x1_sg U74533 ( .A(\reg_y[13][15] ), .X(n50771) );
  nand_x1_sg U74534 ( .A(\reg_yHat[14][9] ), .B(n50932), .X(n26681) );
  inv_x1_sg U74535 ( .A(\reg_y[14][9] ), .X(n50932) );
  nand_x1_sg U74536 ( .A(\reg_y[14][10] ), .B(n46833), .X(n26674) );
  inv_x1_sg U74537 ( .A(\reg_yHat[14][10] ), .X(n46833) );
  nand_x1_sg U74538 ( .A(\reg_y[14][9] ), .B(n46832), .X(n26679) );
  inv_x1_sg U74539 ( .A(\reg_yHat[14][9] ), .X(n46832) );
  nand_x1_sg U74540 ( .A(\reg_yHat[14][10] ), .B(n50949), .X(n26672) );
  inv_x1_sg U74541 ( .A(\reg_y[14][10] ), .X(n50949) );
  nand_x1_sg U74542 ( .A(\reg_yHat[14][11] ), .B(n50971), .X(n26667) );
  inv_x1_sg U74543 ( .A(\reg_y[14][11] ), .X(n50971) );
  nand_x1_sg U74544 ( .A(\reg_y[14][12] ), .B(n46835), .X(n26660) );
  inv_x1_sg U74545 ( .A(\reg_yHat[14][12] ), .X(n46835) );
  nand_x1_sg U74546 ( .A(\reg_y[14][11] ), .B(n46834), .X(n26665) );
  inv_x1_sg U74547 ( .A(\reg_yHat[14][11] ), .X(n46834) );
  nand_x1_sg U74548 ( .A(\reg_yHat[14][12] ), .B(n50989), .X(n26658) );
  inv_x1_sg U74549 ( .A(\reg_y[14][12] ), .X(n50989) );
  nand_x1_sg U74550 ( .A(\reg_yHat[14][13] ), .B(n51011), .X(n26653) );
  inv_x1_sg U74551 ( .A(\reg_y[14][13] ), .X(n51011) );
  nand_x1_sg U74552 ( .A(\reg_y[14][14] ), .B(n46837), .X(n26646) );
  inv_x1_sg U74553 ( .A(\reg_yHat[14][14] ), .X(n46837) );
  nand_x1_sg U74554 ( .A(\reg_y[14][13] ), .B(n46836), .X(n26651) );
  inv_x1_sg U74555 ( .A(\reg_yHat[14][13] ), .X(n46836) );
  nand_x1_sg U74556 ( .A(\reg_yHat[14][14] ), .B(n51029), .X(n26644) );
  inv_x1_sg U74557 ( .A(\reg_y[14][14] ), .X(n51029) );
  nand_x1_sg U74558 ( .A(\reg_y[14][15] ), .B(n46838), .X(n26637) );
  inv_x1_sg U74559 ( .A(\reg_yHat[14][15] ), .X(n46838) );
  nand_x1_sg U74560 ( .A(\reg_yHat[14][15] ), .B(n51058), .X(n26639) );
  inv_x1_sg U74561 ( .A(\reg_y[14][15] ), .X(n51058) );
  nand_x1_sg U74562 ( .A(\reg_y[0][16] ), .B(n46645), .X(n22729) );
  inv_x1_sg U74563 ( .A(\reg_yHat[0][16] ), .X(n46645) );
  nand_x1_sg U74564 ( .A(\reg_yHat[0][16] ), .B(n47073), .X(n22727) );
  inv_x1_sg U74565 ( .A(\reg_y[0][16] ), .X(n47073) );
  nand_x1_sg U74566 ( .A(\reg_y[1][16] ), .B(n46658), .X(n23006) );
  inv_x1_sg U74567 ( .A(\reg_yHat[1][16] ), .X(n46658) );
  nand_x1_sg U74568 ( .A(\reg_yHat[1][16] ), .B(n47359), .X(n23004) );
  inv_x1_sg U74569 ( .A(\reg_y[1][16] ), .X(n47359) );
  nand_x1_sg U74570 ( .A(\reg_y[2][16] ), .B(n46672), .X(n23286) );
  inv_x1_sg U74571 ( .A(\reg_yHat[2][16] ), .X(n46672) );
  nand_x1_sg U74572 ( .A(\reg_yHat[2][16] ), .B(n47644), .X(n23284) );
  inv_x1_sg U74573 ( .A(\reg_y[2][16] ), .X(n47644) );
  nand_x1_sg U74574 ( .A(\reg_y[3][16] ), .B(n46686), .X(n23565) );
  inv_x1_sg U74575 ( .A(\reg_yHat[3][16] ), .X(n46686) );
  nand_x1_sg U74576 ( .A(\reg_yHat[3][16] ), .B(n47929), .X(n23563) );
  inv_x1_sg U74577 ( .A(\reg_y[3][16] ), .X(n47929) );
  nand_x1_sg U74578 ( .A(\reg_y[4][16] ), .B(n46700), .X(n23844) );
  inv_x1_sg U74579 ( .A(\reg_yHat[4][16] ), .X(n46700) );
  nand_x1_sg U74580 ( .A(\reg_yHat[4][16] ), .B(n48214), .X(n23842) );
  inv_x1_sg U74581 ( .A(\reg_y[4][16] ), .X(n48214) );
  nand_x1_sg U74582 ( .A(\reg_y[5][16] ), .B(n46714), .X(n24123) );
  inv_x1_sg U74583 ( .A(\reg_yHat[5][16] ), .X(n46714) );
  nand_x1_sg U74584 ( .A(\reg_yHat[5][16] ), .B(n48499), .X(n24121) );
  inv_x1_sg U74585 ( .A(\reg_y[5][16] ), .X(n48499) );
  nand_x1_sg U74586 ( .A(\reg_y[6][16] ), .B(n46728), .X(n24402) );
  inv_x1_sg U74587 ( .A(\reg_yHat[6][16] ), .X(n46728) );
  nand_x1_sg U74588 ( .A(\reg_yHat[6][16] ), .B(n48784), .X(n24400) );
  inv_x1_sg U74589 ( .A(\reg_y[6][16] ), .X(n48784) );
  nand_x1_sg U74590 ( .A(\reg_y[7][16] ), .B(n46742), .X(n24680) );
  inv_x1_sg U74591 ( .A(\reg_yHat[7][16] ), .X(n46742) );
  nand_x1_sg U74592 ( .A(\reg_yHat[7][16] ), .B(n49071), .X(n24678) );
  inv_x1_sg U74593 ( .A(\reg_y[7][16] ), .X(n49071) );
  nand_x1_sg U74594 ( .A(\reg_y[8][16] ), .B(n46756), .X(n24959) );
  inv_x1_sg U74595 ( .A(\reg_yHat[8][16] ), .X(n46756) );
  nand_x1_sg U74596 ( .A(\reg_yHat[8][16] ), .B(n49357), .X(n24957) );
  inv_x1_sg U74597 ( .A(\reg_y[8][16] ), .X(n49357) );
  nand_x1_sg U74598 ( .A(\reg_y[9][16] ), .B(n46770), .X(n25238) );
  inv_x1_sg U74599 ( .A(\reg_yHat[9][16] ), .X(n46770) );
  nand_x1_sg U74600 ( .A(\reg_yHat[9][16] ), .B(n49643), .X(n25236) );
  inv_x1_sg U74601 ( .A(\reg_y[9][16] ), .X(n49643) );
  nand_x1_sg U74602 ( .A(\reg_y[10][16] ), .B(n46784), .X(n25517) );
  inv_x1_sg U74603 ( .A(\reg_yHat[10][16] ), .X(n46784) );
  nand_x1_sg U74604 ( .A(\reg_yHat[10][16] ), .B(n49929), .X(n25515) );
  inv_x1_sg U74605 ( .A(\reg_y[10][16] ), .X(n49929) );
  nand_x1_sg U74606 ( .A(\reg_y[11][16] ), .B(n46798), .X(n25794) );
  inv_x1_sg U74607 ( .A(\reg_yHat[11][16] ), .X(n46798) );
  nand_x1_sg U74608 ( .A(\reg_yHat[11][16] ), .B(n50215), .X(n25792) );
  inv_x1_sg U74609 ( .A(\reg_y[11][16] ), .X(n50215) );
  nand_x1_sg U74610 ( .A(\reg_y[12][16] ), .B(n46812), .X(n26138) );
  inv_x1_sg U74611 ( .A(\reg_yHat[12][16] ), .X(n46812) );
  nand_x1_sg U74612 ( .A(\reg_yHat[12][16] ), .B(n50501), .X(n26139) );
  inv_x1_sg U74613 ( .A(\reg_y[12][16] ), .X(n50501) );
  nand_x1_sg U74614 ( .A(\reg_y[13][16] ), .B(n46825), .X(n26354) );
  inv_x1_sg U74615 ( .A(\reg_yHat[13][16] ), .X(n46825) );
  nand_x1_sg U74616 ( .A(\reg_yHat[13][16] ), .B(n50789), .X(n26352) );
  inv_x1_sg U74617 ( .A(\reg_y[13][16] ), .X(n50789) );
  nand_x1_sg U74618 ( .A(\reg_y[14][16] ), .B(n46839), .X(n26632) );
  inv_x1_sg U74619 ( .A(\reg_yHat[14][16] ), .X(n46839) );
  nand_x1_sg U74620 ( .A(\reg_yHat[14][16] ), .B(n51076), .X(n26630) );
  inv_x1_sg U74621 ( .A(\reg_y[14][16] ), .X(n51076) );
  nand_x1_sg U74622 ( .A(n5727), .B(n22565), .X(n27800) );
  nor_x1_sg U74623 ( .A(n22565), .B(n5727), .X(n27801) );
  nand_x1_sg U74624 ( .A(n5721), .B(n22583), .X(n28621) );
  nor_x1_sg U74625 ( .A(n22583), .B(n5721), .X(n28622) );
  nand_x1_sg U74626 ( .A(n5729), .B(n22569), .X(n27411) );
  nor_x1_sg U74627 ( .A(n22569), .B(n5729), .X(n27412) );
  nor_x1_sg U74628 ( .A(n22594), .B(n5723), .X(n28367) );
  inv_x1_sg U74629 ( .A(\reg_y[1][6] ), .X(n47171) );
  inv_x1_sg U74630 ( .A(\reg_y[2][6] ), .X(n47456) );
  inv_x1_sg U74631 ( .A(\reg_y[3][6] ), .X(n47741) );
  inv_x1_sg U74632 ( .A(\reg_y[4][6] ), .X(n48026) );
  inv_x1_sg U74633 ( .A(\reg_y[5][6] ), .X(n48311) );
  inv_x1_sg U74634 ( .A(\reg_y[6][6] ), .X(n48596) );
  inv_x1_sg U74635 ( .A(\reg_y[7][6] ), .X(n48882) );
  inv_x1_sg U74636 ( .A(\reg_y[8][6] ), .X(n49169) );
  inv_x1_sg U74637 ( .A(\reg_y[9][6] ), .X(n49455) );
  inv_x1_sg U74638 ( .A(\reg_y[10][6] ), .X(n49740) );
  inv_x1_sg U74639 ( .A(\reg_y[11][6] ), .X(n50027) );
  inv_x1_sg U74640 ( .A(\reg_y[13][6] ), .X(n50601) );
  inv_x1_sg U74641 ( .A(\reg_y[14][6] ), .X(n50888) );
  inv_x1_sg U74642 ( .A(\reg_y[0][6] ), .X(n46878) );
  inv_x1_sg U74643 ( .A(\reg_y[12][6] ), .X(n50312) );
  inv_x1_sg U74644 ( .A(\reg_yHat[0][1] ), .X(n46633) );
  inv_x1_sg U74645 ( .A(\reg_yHat[1][1] ), .X(n46646) );
  inv_x1_sg U74646 ( .A(\reg_yHat[2][1] ), .X(n46660) );
  inv_x1_sg U74647 ( .A(\reg_yHat[3][1] ), .X(n46674) );
  inv_x1_sg U74648 ( .A(\reg_yHat[4][1] ), .X(n46688) );
  inv_x1_sg U74649 ( .A(\reg_yHat[5][1] ), .X(n46702) );
  inv_x1_sg U74650 ( .A(\reg_yHat[6][1] ), .X(n46716) );
  inv_x1_sg U74651 ( .A(\reg_yHat[7][1] ), .X(n46730) );
  inv_x1_sg U74652 ( .A(\reg_yHat[8][1] ), .X(n46744) );
  inv_x1_sg U74653 ( .A(\reg_yHat[9][1] ), .X(n46758) );
  inv_x1_sg U74654 ( .A(\reg_yHat[10][1] ), .X(n46772) );
  inv_x1_sg U74655 ( .A(\reg_yHat[11][1] ), .X(n46786) );
  inv_x1_sg U74656 ( .A(\reg_yHat[13][1] ), .X(n46813) );
  inv_x1_sg U74657 ( .A(\reg_yHat[14][1] ), .X(n46827) );
  inv_x1_sg U74658 ( .A(\reg_yHat[12][1] ), .X(n46800) );
  nand_x1_sg U74659 ( .A(n22816), .B(n46634), .X(n22813) );
  nand_x1_sg U74660 ( .A(\reg_y[0][4] ), .B(n22815), .X(n22814) );
  nand_x1_sg U74661 ( .A(\reg_yHat[0][4] ), .B(n46850), .X(n22815) );
  nand_x1_sg U74662 ( .A(n47143), .B(n46647), .X(n23090) );
  nand_x1_sg U74663 ( .A(\reg_y[1][4] ), .B(n23092), .X(n23091) );
  nand_x1_sg U74664 ( .A(\reg_yHat[1][4] ), .B(n23093), .X(n23092) );
  nand_x1_sg U74665 ( .A(n47428), .B(n46661), .X(n23370) );
  nand_x1_sg U74666 ( .A(\reg_y[2][4] ), .B(n23372), .X(n23371) );
  nand_x1_sg U74667 ( .A(\reg_yHat[2][4] ), .B(n23373), .X(n23372) );
  nand_x1_sg U74668 ( .A(n47713), .B(n46675), .X(n23649) );
  nand_x1_sg U74669 ( .A(\reg_y[3][4] ), .B(n23651), .X(n23650) );
  nand_x1_sg U74670 ( .A(\reg_yHat[3][4] ), .B(n23652), .X(n23651) );
  nand_x1_sg U74671 ( .A(n47998), .B(n46689), .X(n23928) );
  nand_x1_sg U74672 ( .A(\reg_y[4][4] ), .B(n23930), .X(n23929) );
  nand_x1_sg U74673 ( .A(\reg_yHat[4][4] ), .B(n23931), .X(n23930) );
  nand_x1_sg U74674 ( .A(n48283), .B(n46703), .X(n24207) );
  nand_x1_sg U74675 ( .A(\reg_y[5][4] ), .B(n24209), .X(n24208) );
  nand_x1_sg U74676 ( .A(\reg_yHat[5][4] ), .B(n24210), .X(n24209) );
  nand_x1_sg U74677 ( .A(n48568), .B(n46717), .X(n24486) );
  nand_x1_sg U74678 ( .A(\reg_y[6][4] ), .B(n24488), .X(n24487) );
  nand_x1_sg U74679 ( .A(\reg_yHat[6][4] ), .B(n24489), .X(n24488) );
  nand_x1_sg U74680 ( .A(n48853), .B(n46731), .X(n24764) );
  nand_x1_sg U74681 ( .A(\reg_y[7][4] ), .B(n24766), .X(n24765) );
  nand_x1_sg U74682 ( .A(\reg_yHat[7][4] ), .B(n24767), .X(n24766) );
  nand_x1_sg U74683 ( .A(n49140), .B(n46745), .X(n25043) );
  nand_x1_sg U74684 ( .A(\reg_y[8][4] ), .B(n25045), .X(n25044) );
  nand_x1_sg U74685 ( .A(\reg_yHat[8][4] ), .B(n25046), .X(n25045) );
  nand_x1_sg U74686 ( .A(n49426), .B(n46759), .X(n25322) );
  nand_x1_sg U74687 ( .A(\reg_y[9][4] ), .B(n25324), .X(n25323) );
  nand_x1_sg U74688 ( .A(\reg_yHat[9][4] ), .B(n25325), .X(n25324) );
  nand_x1_sg U74689 ( .A(n49712), .B(n46773), .X(n25601) );
  nand_x1_sg U74690 ( .A(\reg_y[10][4] ), .B(n25603), .X(n25602) );
  nand_x1_sg U74691 ( .A(\reg_yHat[10][4] ), .B(n25604), .X(n25603) );
  nand_x1_sg U74692 ( .A(n49998), .B(n46787), .X(n25878) );
  nand_x1_sg U74693 ( .A(\reg_y[11][4] ), .B(n25880), .X(n25879) );
  nand_x1_sg U74694 ( .A(\reg_yHat[11][4] ), .B(n25881), .X(n25880) );
  nand_x1_sg U74695 ( .A(n50573), .B(n46814), .X(n26438) );
  nand_x1_sg U74696 ( .A(\reg_y[13][4] ), .B(n26440), .X(n26439) );
  nand_x1_sg U74697 ( .A(\reg_yHat[13][4] ), .B(n26441), .X(n26440) );
  nand_x1_sg U74698 ( .A(n50859), .B(n46828), .X(n26716) );
  nand_x1_sg U74699 ( .A(\reg_y[14][4] ), .B(n26718), .X(n26717) );
  nand_x1_sg U74700 ( .A(\reg_yHat[14][4] ), .B(n26719), .X(n26718) );
  nand_x1_sg U74701 ( .A(\reg_yHat[12][2] ), .B(n26120), .X(n26172) );
  nand_x1_sg U74702 ( .A(n38623), .B(n38520), .X(n27805) );
  nand_x1_sg U74703 ( .A(n38602), .B(n38521), .X(n28626) );
  nand_x1_sg U74704 ( .A(n38621), .B(n38522), .X(n28371) );
  nand_x1_sg U74705 ( .A(n38628), .B(n38523), .X(n27416) );
  nand_x1_sg U74706 ( .A(n38619), .B(n38524), .X(n26954) );
  inv_x1_sg U74707 ( .A(\reg_y[0][3] ), .X(n46851) );
  inv_x1_sg U74708 ( .A(\reg_y[1][3] ), .X(n47144) );
  inv_x1_sg U74709 ( .A(\reg_y[2][3] ), .X(n47429) );
  inv_x1_sg U74710 ( .A(\reg_y[3][3] ), .X(n47714) );
  inv_x1_sg U74711 ( .A(\reg_y[4][3] ), .X(n47999) );
  inv_x1_sg U74712 ( .A(\reg_y[5][3] ), .X(n48284) );
  inv_x1_sg U74713 ( .A(\reg_y[6][3] ), .X(n48569) );
  inv_x1_sg U74714 ( .A(\reg_y[7][3] ), .X(n48854) );
  inv_x1_sg U74715 ( .A(\reg_y[8][3] ), .X(n49141) );
  inv_x1_sg U74716 ( .A(\reg_y[9][3] ), .X(n49427) );
  inv_x1_sg U74717 ( .A(\reg_y[10][3] ), .X(n49713) );
  inv_x1_sg U74718 ( .A(\reg_y[11][3] ), .X(n49999) );
  inv_x1_sg U74719 ( .A(\reg_y[13][3] ), .X(n50574) );
  inv_x1_sg U74720 ( .A(\reg_y[14][3] ), .X(n50860) );
  nand_x1_sg U74721 ( .A(n39486), .B(n17465), .X(n5977) );
  inv_x1_sg U74722 ( .A(\reg_y[1][2] ), .X(n47138) );
  inv_x1_sg U74723 ( .A(\reg_y[2][2] ), .X(n47423) );
  inv_x1_sg U74724 ( .A(\reg_y[3][2] ), .X(n47708) );
  inv_x1_sg U74725 ( .A(\reg_y[4][2] ), .X(n47993) );
  inv_x1_sg U74726 ( .A(\reg_y[5][2] ), .X(n48278) );
  inv_x1_sg U74727 ( .A(\reg_y[6][2] ), .X(n48563) );
  inv_x1_sg U74728 ( .A(\reg_y[7][2] ), .X(n48848) );
  inv_x1_sg U74729 ( .A(\reg_y[8][2] ), .X(n49135) );
  inv_x1_sg U74730 ( .A(\reg_y[9][2] ), .X(n49421) );
  inv_x1_sg U74731 ( .A(\reg_y[10][2] ), .X(n49707) );
  inv_x1_sg U74732 ( .A(\reg_y[11][2] ), .X(n49993) );
  inv_x1_sg U74733 ( .A(\reg_y[13][2] ), .X(n50568) );
  inv_x1_sg U74734 ( .A(\reg_y[14][2] ), .X(n50854) );
  nand_x1_sg U74735 ( .A(n29149), .B(n42114), .X(n29263) );
  nand_x1_sg U74736 ( .A(n29161), .B(n42115), .X(n29257) );
  nand_x1_sg U74737 ( .A(n29173), .B(n42116), .X(n29251) );
  nand_x1_sg U74738 ( .A(n29185), .B(n42117), .X(n29245) );
  nand_x1_sg U74739 ( .A(n21658), .B(n42112), .X(n21682) );
  nand_x1_sg U74740 ( .A(n21646), .B(n42111), .X(n21688) );
  nand_x1_sg U74741 ( .A(n21634), .B(n42110), .X(n21694) );
  nand_x1_sg U74742 ( .A(n21622), .B(n42109), .X(n21700) );
  nand_x1_sg U74743 ( .A(n29197), .B(n38121), .X(n29239) );
  nand_x1_sg U74744 ( .A(n29209), .B(n38122), .X(n29233) );
  nand_x1_sg U74745 ( .A(n29221), .B(n38124), .X(n29227) );
  nand_x1_sg U74746 ( .A(n21670), .B(n38123), .X(n21676) );
  nand_x1_sg U74747 ( .A(n23102), .B(n38764), .X(n23099) );
  nor_x1_sg U74748 ( .A(n23101), .B(\reg_y[1][3] ), .X(n23100) );
  nand_x1_sg U74749 ( .A(n23382), .B(n38768), .X(n23379) );
  nor_x1_sg U74750 ( .A(n23381), .B(\reg_y[2][3] ), .X(n23380) );
  nand_x1_sg U74751 ( .A(n23661), .B(n38772), .X(n23658) );
  nor_x1_sg U74752 ( .A(n23660), .B(\reg_y[3][3] ), .X(n23659) );
  nand_x1_sg U74753 ( .A(n23940), .B(n38776), .X(n23937) );
  nor_x1_sg U74754 ( .A(n23939), .B(\reg_y[4][3] ), .X(n23938) );
  nand_x1_sg U74755 ( .A(n24219), .B(n38780), .X(n24216) );
  nor_x1_sg U74756 ( .A(n24218), .B(\reg_y[5][3] ), .X(n24217) );
  nand_x1_sg U74757 ( .A(n24498), .B(n38784), .X(n24495) );
  nor_x1_sg U74758 ( .A(n24497), .B(\reg_y[6][3] ), .X(n24496) );
  nand_x1_sg U74759 ( .A(n24776), .B(n38788), .X(n24773) );
  nor_x1_sg U74760 ( .A(n24775), .B(\reg_y[7][3] ), .X(n24774) );
  nand_x1_sg U74761 ( .A(n25055), .B(n38792), .X(n25052) );
  nor_x1_sg U74762 ( .A(n25054), .B(\reg_y[8][3] ), .X(n25053) );
  nand_x1_sg U74763 ( .A(n25334), .B(n38796), .X(n25331) );
  nor_x1_sg U74764 ( .A(n25333), .B(\reg_y[9][3] ), .X(n25332) );
  nand_x1_sg U74765 ( .A(n25613), .B(n38800), .X(n25610) );
  nor_x1_sg U74766 ( .A(n25612), .B(\reg_y[10][3] ), .X(n25611) );
  nand_x1_sg U74767 ( .A(n25890), .B(n38804), .X(n25887) );
  nor_x1_sg U74768 ( .A(n25889), .B(\reg_y[11][3] ), .X(n25888) );
  nand_x1_sg U74769 ( .A(n26450), .B(n38808), .X(n26447) );
  nor_x1_sg U74770 ( .A(n26449), .B(\reg_y[13][3] ), .X(n26448) );
  nand_x1_sg U74771 ( .A(n26728), .B(n38812), .X(n26725) );
  nor_x1_sg U74772 ( .A(n26727), .B(\reg_y[14][3] ), .X(n26726) );
  nor_x1_sg U74773 ( .A(n16837), .B(n16838), .X(n16836) );
  nor_x1_sg U74774 ( .A(n50522), .B(n42005), .X(n16838) );
  nor_x1_sg U74775 ( .A(\reg_y[12][17] ), .B(n16839), .X(n16837) );
  nor_x1_sg U74776 ( .A(\reg_yHat[12][17] ), .B(n16840), .X(n16839) );
  nand_x1_sg U74777 ( .A(n45825), .B(n38173), .X(n21063) );
  nand_x1_sg U74778 ( .A(n21065), .B(n45801), .X(n21064) );
  nor_x1_sg U74779 ( .A(n5707), .B(n20847), .X(n21065) );
  nand_x1_sg U74780 ( .A(n45841), .B(n38174), .X(n20354) );
  nand_x1_sg U74781 ( .A(n20356), .B(n45805), .X(n20355) );
  nor_x1_sg U74782 ( .A(n5711), .B(n20204), .X(n20356) );
  nand_x1_sg U74783 ( .A(n45857), .B(n38175), .X(n19621) );
  nand_x1_sg U74784 ( .A(n19623), .B(n45809), .X(n19622) );
  nor_x1_sg U74785 ( .A(n5715), .B(n19398), .X(n19623) );
  nor_x1_sg U74786 ( .A(n41122), .B(n42162), .X(n26797) );
  nand_x1_sg U74787 ( .A(\reg_y[1][18] ), .B(n46659), .X(n22999) );
  nor_x1_sg U74788 ( .A(n46659), .B(\reg_y[1][18] ), .X(n23000) );
  nand_x1_sg U74789 ( .A(\reg_y[2][18] ), .B(n46673), .X(n23279) );
  nor_x1_sg U74790 ( .A(n46673), .B(\reg_y[2][18] ), .X(n23280) );
  nand_x1_sg U74791 ( .A(\reg_y[3][18] ), .B(n46687), .X(n23558) );
  nor_x1_sg U74792 ( .A(n46687), .B(\reg_y[3][18] ), .X(n23559) );
  nand_x1_sg U74793 ( .A(\reg_y[4][18] ), .B(n46701), .X(n23837) );
  nor_x1_sg U74794 ( .A(n46701), .B(\reg_y[4][18] ), .X(n23838) );
  nand_x1_sg U74795 ( .A(\reg_y[5][18] ), .B(n46715), .X(n24116) );
  nor_x1_sg U74796 ( .A(n46715), .B(\reg_y[5][18] ), .X(n24117) );
  nand_x1_sg U74797 ( .A(\reg_y[6][18] ), .B(n46729), .X(n24395) );
  nor_x1_sg U74798 ( .A(n46729), .B(\reg_y[6][18] ), .X(n24396) );
  nand_x1_sg U74799 ( .A(\reg_y[7][18] ), .B(n46743), .X(n24673) );
  nor_x1_sg U74800 ( .A(n46743), .B(\reg_y[7][18] ), .X(n24674) );
  nand_x1_sg U74801 ( .A(\reg_y[8][18] ), .B(n46757), .X(n24952) );
  nor_x1_sg U74802 ( .A(n46757), .B(\reg_y[8][18] ), .X(n24953) );
  nand_x1_sg U74803 ( .A(\reg_y[9][18] ), .B(n46771), .X(n25231) );
  nor_x1_sg U74804 ( .A(n46771), .B(\reg_y[9][18] ), .X(n25232) );
  nand_x1_sg U74805 ( .A(\reg_y[10][18] ), .B(n46785), .X(n25510) );
  nor_x1_sg U74806 ( .A(n46785), .B(\reg_y[10][18] ), .X(n25511) );
  nand_x1_sg U74807 ( .A(\reg_y[11][18] ), .B(n46799), .X(n25787) );
  nor_x1_sg U74808 ( .A(n46799), .B(\reg_y[11][18] ), .X(n25788) );
  nand_x1_sg U74809 ( .A(\reg_y[13][18] ), .B(n46826), .X(n26347) );
  nor_x1_sg U74810 ( .A(n46826), .B(\reg_y[13][18] ), .X(n26348) );
  nand_x1_sg U74811 ( .A(\reg_y[14][18] ), .B(n46840), .X(n26625) );
  nor_x1_sg U74812 ( .A(n46840), .B(\reg_y[14][18] ), .X(n26626) );
  nor_x1_sg U74813 ( .A(n5717), .B(n22551), .X(n26949) );
  inv_x1_sg U74814 ( .A(\reg_y[0][1] ), .X(n46842) );
  inv_x1_sg U74815 ( .A(\reg_y[1][1] ), .X(n47135) );
  inv_x1_sg U74816 ( .A(\reg_y[2][1] ), .X(n47420) );
  inv_x1_sg U74817 ( .A(\reg_y[3][1] ), .X(n47705) );
  inv_x1_sg U74818 ( .A(\reg_y[4][1] ), .X(n47990) );
  inv_x1_sg U74819 ( .A(\reg_y[5][1] ), .X(n48275) );
  inv_x1_sg U74820 ( .A(\reg_y[6][1] ), .X(n48560) );
  inv_x1_sg U74821 ( .A(\reg_y[7][1] ), .X(n48845) );
  inv_x1_sg U74822 ( .A(\reg_y[8][1] ), .X(n49132) );
  inv_x1_sg U74823 ( .A(\reg_y[9][1] ), .X(n49418) );
  inv_x1_sg U74824 ( .A(\reg_y[10][1] ), .X(n49704) );
  inv_x1_sg U74825 ( .A(\reg_y[11][1] ), .X(n49990) );
  inv_x1_sg U74826 ( .A(\reg_y[12][5] ), .X(n50300) );
  inv_x1_sg U74827 ( .A(\reg_y[13][1] ), .X(n50563) );
  inv_x1_sg U74828 ( .A(\reg_y[14][1] ), .X(n50851) );
  inv_x1_sg U74829 ( .A(\reg_y[12][1] ), .X(n50276) );
  nand_x1_sg U74830 ( .A(n19478), .B(n19480), .X(n19584) );
  nor_x1_sg U74831 ( .A(n19586), .B(n5461), .X(n19585) );
  nand_x1_sg U74832 ( .A(n28365), .B(n22584), .X(n28364) );
  nand_x1_sg U74833 ( .A(n44993), .B(n38176), .X(n28363) );
  nor_x1_sg U74834 ( .A(n5724), .B(n28259), .X(n28365) );
  nand_x1_sg U74835 ( .A(n28120), .B(n42159), .X(n28119) );
  nand_x1_sg U74836 ( .A(n45000), .B(n38177), .X(n28118) );
  nor_x1_sg U74837 ( .A(n5726), .B(n27975), .X(n28120) );
  nand_x1_sg U74838 ( .A(n45003), .B(n38178), .X(n27965) );
  nand_x1_sg U74839 ( .A(n27967), .B(n38623), .X(n27966) );
  nor_x1_sg U74840 ( .A(n5727), .B(n27806), .X(n27967) );
  nand_x1_sg U74841 ( .A(n27799), .B(n22574), .X(n27798) );
  nand_x1_sg U74842 ( .A(n45006), .B(n38179), .X(n27797) );
  nor_x1_sg U74843 ( .A(n5728), .B(n27620), .X(n27799) );
  nand_x1_sg U74844 ( .A(n44984), .B(n38180), .X(n28806) );
  nand_x1_sg U74845 ( .A(n28808), .B(n38602), .X(n28807) );
  nor_x1_sg U74846 ( .A(n5721), .B(n28627), .X(n28808) );
  nand_x1_sg U74847 ( .A(n45009), .B(n38181), .X(n27612) );
  nand_x1_sg U74848 ( .A(n27614), .B(n22569), .X(n27613) );
  nor_x1_sg U74849 ( .A(n5729), .B(n27417), .X(n27614) );
  nand_x1_sg U74850 ( .A(n21587), .B(n45798), .X(n21586) );
  nand_x1_sg U74851 ( .A(n45814), .B(n38182), .X(n21585) );
  nor_x1_sg U74852 ( .A(n5704), .B(n21435), .X(n21587) );
  nand_x1_sg U74853 ( .A(n28620), .B(n22578), .X(n28619) );
  nand_x1_sg U74854 ( .A(n44987), .B(n38183), .X(n28618) );
  nor_x1_sg U74855 ( .A(n5722), .B(n28466), .X(n28620) );
  nand_x1_sg U74856 ( .A(n29138), .B(n44964), .X(n29137) );
  nand_x1_sg U74857 ( .A(n44978), .B(n38184), .X(n29136) );
  nor_x1_sg U74858 ( .A(n5719), .B(n28986), .X(n29138) );
  nand_x1_sg U74859 ( .A(n27410), .B(n22566), .X(n27409) );
  nand_x1_sg U74860 ( .A(n45012), .B(n38185), .X(n27408) );
  nor_x1_sg U74861 ( .A(n5730), .B(n27195), .X(n27410) );
  nand_x1_sg U74862 ( .A(n44990), .B(n38186), .X(n28458) );
  nand_x1_sg U74863 ( .A(n28460), .B(n38621), .X(n28459) );
  nor_x1_sg U74864 ( .A(n5723), .B(n28372), .X(n28460) );
  nand_x1_sg U74865 ( .A(n44981), .B(n38187), .X(n28976) );
  nand_x1_sg U74866 ( .A(n28978), .B(n38756), .X(n28977) );
  nor_x1_sg U74867 ( .A(n5720), .B(n28815), .X(n28978) );
  nand_x1_sg U74868 ( .A(n45015), .B(n38188), .X(n27187) );
  nand_x1_sg U74869 ( .A(n27189), .B(n38619), .X(n27188) );
  nor_x1_sg U74870 ( .A(n5731), .B(n26956), .X(n27189) );
  nor_x1_sg U74871 ( .A(n22575), .B(n5731), .X(n26951) );
  inv_x1_sg U74872 ( .A(\reg_y[0][0] ), .X(n46841) );
  inv_x1_sg U74873 ( .A(\reg_y[1][0] ), .X(n47133) );
  inv_x1_sg U74874 ( .A(\reg_y[2][0] ), .X(n47419) );
  inv_x1_sg U74875 ( .A(\reg_y[3][0] ), .X(n47704) );
  inv_x1_sg U74876 ( .A(\reg_y[4][0] ), .X(n47989) );
  inv_x1_sg U74877 ( .A(\reg_y[5][0] ), .X(n48274) );
  inv_x1_sg U74878 ( .A(\reg_y[6][0] ), .X(n48559) );
  inv_x1_sg U74879 ( .A(\reg_y[7][0] ), .X(n48844) );
  inv_x1_sg U74880 ( .A(\reg_y[8][0] ), .X(n49131) );
  inv_x1_sg U74881 ( .A(\reg_y[9][0] ), .X(n49417) );
  inv_x1_sg U74882 ( .A(\reg_y[10][0] ), .X(n49703) );
  inv_x1_sg U74883 ( .A(\reg_y[11][0] ), .X(n49989) );
  inv_x1_sg U74884 ( .A(\reg_y[13][0] ), .X(n50562) );
  inv_x1_sg U74885 ( .A(\reg_y[14][0] ), .X(n50849) );
  inv_x1_sg U74886 ( .A(\reg_y[1][19] ), .X(n47413) );
  inv_x1_sg U74887 ( .A(\reg_y[2][19] ), .X(n47698) );
  inv_x1_sg U74888 ( .A(\reg_y[3][19] ), .X(n47983) );
  inv_x1_sg U74889 ( .A(\reg_y[4][19] ), .X(n48268) );
  inv_x1_sg U74890 ( .A(\reg_y[5][19] ), .X(n48553) );
  inv_x1_sg U74891 ( .A(\reg_y[6][19] ), .X(n48838) );
  inv_x1_sg U74892 ( .A(\reg_y[7][19] ), .X(n49125) );
  inv_x1_sg U74893 ( .A(\reg_y[8][19] ), .X(n49411) );
  inv_x1_sg U74894 ( .A(\reg_y[9][19] ), .X(n49697) );
  inv_x1_sg U74895 ( .A(\reg_y[10][19] ), .X(n49983) );
  inv_x1_sg U74896 ( .A(\reg_y[11][19] ), .X(n50269) );
  inv_x1_sg U74897 ( .A(\reg_y[13][19] ), .X(n50844) );
  inv_x1_sg U74898 ( .A(\reg_y[14][19] ), .X(n51130) );
  inv_x1_sg U74899 ( .A(\reg_y[12][0] ), .X(n50275) );
  inv_x1_sg U74900 ( .A(\reg_y[0][19] ), .X(n47128) );
  inv_x1_sg U74901 ( .A(\reg_y[12][19] ), .X(n50557) );
  nand_x1_sg U74902 ( .A(n5517), .B(n46397), .X(n20115) );
  nand_x1_sg U74903 ( .A(n20116), .B(n38525), .X(n20114) );
  nand_x1_sg U74904 ( .A(n5477), .B(n46484), .X(n19721) );
  nand_x1_sg U74905 ( .A(n19722), .B(n38526), .X(n19720) );
  nand_x1_sg U74906 ( .A(n5421), .B(n46434), .X(n6130) );
  nand_x1_sg U74907 ( .A(n6131), .B(n38198), .X(n6129) );
  nand_x1_sg U74908 ( .A(n5572), .B(n46489), .X(n20135) );
  nand_x1_sg U74909 ( .A(n20136), .B(n38199), .X(n20134) );
  nand_x1_sg U74910 ( .A(n5423), .B(n46341), .X(n6222) );
  nand_x1_sg U74911 ( .A(n6223), .B(n38200), .X(n6221) );
  nand_x1_sg U74912 ( .A(n5646), .B(n46547), .X(n21196) );
  nand_x1_sg U74913 ( .A(n20998), .B(n38201), .X(n21195) );
  nand_x1_sg U74914 ( .A(n5604), .B(n45906), .X(n20679) );
  nand_x1_sg U74915 ( .A(n20680), .B(n38202), .X(n20678) );
  nand_x1_sg U74916 ( .A(n5528), .B(n45896), .X(n20039) );
  nand_x1_sg U74917 ( .A(n20040), .B(n38203), .X(n20038) );
  nand_x1_sg U74918 ( .A(n5452), .B(n45886), .X(n19235) );
  nand_x1_sg U74919 ( .A(n19236), .B(n38204), .X(n19234) );
  nor_x1_sg U74920 ( .A(n5717), .B(n41276), .X(n22588) );
  nand_x1_sg U74921 ( .A(n46528), .B(n38527), .X(n19505) );
  nand_x1_sg U74922 ( .A(n5457), .B(n19507), .X(n19506) );
  nand_x1_sg U74923 ( .A(n46358), .B(n38205), .X(n20748) );
  nand_x1_sg U74924 ( .A(n46316), .B(n38206), .X(n20741) );
  nand_x1_sg U74925 ( .A(n46271), .B(n38207), .X(n20734) );
  nand_x1_sg U74926 ( .A(n46225), .B(n38208), .X(n20727) );
  nand_x1_sg U74927 ( .A(n46180), .B(n38209), .X(n20720) );
  nand_x1_sg U74928 ( .A(n46134), .B(n38210), .X(n20713) );
  nand_x1_sg U74929 ( .A(n46089), .B(n38211), .X(n20706) );
  nand_x1_sg U74930 ( .A(n46043), .B(n38212), .X(n20699) );
  nand_x1_sg U74931 ( .A(n45998), .B(n38213), .X(n20692) );
  nand_x1_sg U74932 ( .A(n45953), .B(n38214), .X(n20685) );
  nand_x1_sg U74933 ( .A(n46405), .B(n38215), .X(n20755) );
  nand_x1_sg U74934 ( .A(n46453), .B(n38216), .X(n20762) );
  nand_x1_sg U74935 ( .A(n46491), .B(n38217), .X(n20769) );
  nand_x1_sg U74936 ( .A(n46307), .B(n38218), .X(n20101) );
  nand_x1_sg U74937 ( .A(n46262), .B(n38219), .X(n20094) );
  nand_x1_sg U74938 ( .A(n46216), .B(n38220), .X(n20087) );
  nand_x1_sg U74939 ( .A(n46171), .B(n38221), .X(n20080) );
  nand_x1_sg U74940 ( .A(n46125), .B(n38222), .X(n20073) );
  nand_x1_sg U74941 ( .A(n46080), .B(n38223), .X(n20066) );
  nand_x1_sg U74942 ( .A(n46034), .B(n38224), .X(n20059) );
  nand_x1_sg U74943 ( .A(n45989), .B(n38225), .X(n20052) );
  nand_x1_sg U74944 ( .A(n45944), .B(n38226), .X(n20045) );
  nand_x1_sg U74945 ( .A(n46298), .B(n38227), .X(n19297) );
  nand_x1_sg U74946 ( .A(n46253), .B(n38228), .X(n19290) );
  nand_x1_sg U74947 ( .A(n46207), .B(n38229), .X(n19283) );
  nand_x1_sg U74948 ( .A(n46162), .B(n38230), .X(n19276) );
  nand_x1_sg U74949 ( .A(n46116), .B(n38231), .X(n19269) );
  nand_x1_sg U74950 ( .A(n46071), .B(n38232), .X(n19262) );
  nand_x1_sg U74951 ( .A(n46025), .B(n38233), .X(n19255) );
  nand_x1_sg U74952 ( .A(n45980), .B(n38234), .X(n19248) );
  nand_x1_sg U74953 ( .A(n45935), .B(n38235), .X(n19241) );
  nand_x1_sg U74954 ( .A(n5282), .B(n28135), .X(n28134) );
  nor_x1_sg U74955 ( .A(n28135), .B(n5282), .X(n28136) );
  nand_x1_sg U74956 ( .A(n5654), .B(n46231), .X(n21311) );
  nor_x1_sg U74957 ( .A(n46231), .B(n5654), .X(n21312) );
  nand_x1_sg U74958 ( .A(n5655), .B(n46186), .X(n21306) );
  nor_x1_sg U74959 ( .A(n46186), .B(n5655), .X(n21307) );
  nand_x1_sg U74960 ( .A(n5656), .B(n46140), .X(n21301) );
  nor_x1_sg U74961 ( .A(n46140), .B(n5656), .X(n21302) );
  nand_x1_sg U74962 ( .A(n5657), .B(n46095), .X(n21296) );
  nor_x1_sg U74963 ( .A(n46095), .B(n5657), .X(n21297) );
  nand_x1_sg U74964 ( .A(n5658), .B(n46049), .X(n21291) );
  nor_x1_sg U74965 ( .A(n46049), .B(n5658), .X(n21292) );
  nand_x1_sg U74966 ( .A(n5659), .B(n46004), .X(n21286) );
  nor_x1_sg U74967 ( .A(n46004), .B(n5659), .X(n21287) );
  nand_x1_sg U74968 ( .A(n5660), .B(n45959), .X(n21281) );
  nor_x1_sg U74969 ( .A(n45959), .B(n5660), .X(n21282) );
  nand_x1_sg U74970 ( .A(n5653), .B(n46277), .X(n21316) );
  nor_x1_sg U74971 ( .A(n46277), .B(n5653), .X(n21317) );
  nand_x1_sg U74972 ( .A(n5642), .B(n45911), .X(n21085) );
  nor_x1_sg U74973 ( .A(n45911), .B(n5642), .X(n21086) );
  nand_x1_sg U74974 ( .A(n5652), .B(n46322), .X(n21321) );
  nor_x1_sg U74975 ( .A(n46322), .B(n5652), .X(n21322) );
  nand_x1_sg U74976 ( .A(n5651), .B(n46364), .X(n21326) );
  nor_x1_sg U74977 ( .A(n46364), .B(n5651), .X(n21327) );
  nand_x1_sg U74978 ( .A(n5650), .B(n46411), .X(n21331) );
  nor_x1_sg U74979 ( .A(n46411), .B(n5650), .X(n21332) );
  nand_x1_sg U74980 ( .A(n5575), .B(n46355), .X(n20557) );
  nor_x1_sg U74981 ( .A(n46355), .B(n5575), .X(n20558) );
  nand_x1_sg U74982 ( .A(n5576), .B(n46313), .X(n20552) );
  nor_x1_sg U74983 ( .A(n46313), .B(n5576), .X(n20553) );
  nand_x1_sg U74984 ( .A(n5577), .B(n46268), .X(n20547) );
  nor_x1_sg U74985 ( .A(n46268), .B(n5577), .X(n20548) );
  nand_x1_sg U74986 ( .A(n5578), .B(n46222), .X(n20542) );
  nor_x1_sg U74987 ( .A(n46222), .B(n5578), .X(n20543) );
  nand_x1_sg U74988 ( .A(n5579), .B(n46177), .X(n20537) );
  nor_x1_sg U74989 ( .A(n46177), .B(n5579), .X(n20538) );
  nand_x1_sg U74990 ( .A(n5580), .B(n46131), .X(n20532) );
  nor_x1_sg U74991 ( .A(n46131), .B(n5580), .X(n20533) );
  nand_x1_sg U74992 ( .A(n5581), .B(n46086), .X(n20527) );
  nor_x1_sg U74993 ( .A(n46086), .B(n5581), .X(n20528) );
  nand_x1_sg U74994 ( .A(n5582), .B(n46040), .X(n20522) );
  nor_x1_sg U74995 ( .A(n46040), .B(n5582), .X(n20523) );
  nand_x1_sg U74996 ( .A(n5583), .B(n45995), .X(n20517) );
  nor_x1_sg U74997 ( .A(n45995), .B(n5583), .X(n20518) );
  nand_x1_sg U74998 ( .A(n5584), .B(n45950), .X(n20512) );
  nor_x1_sg U74999 ( .A(n45950), .B(n5584), .X(n20513) );
  nand_x1_sg U75000 ( .A(n5649), .B(n46459), .X(n21336) );
  nor_x1_sg U75001 ( .A(n46459), .B(n5649), .X(n21337) );
  nand_x1_sg U75002 ( .A(n5566), .B(n45901), .X(n20376) );
  nor_x1_sg U75003 ( .A(n45901), .B(n5566), .X(n20377) );
  nand_x1_sg U75004 ( .A(n5648), .B(n46497), .X(n21342) );
  nor_x1_sg U75005 ( .A(n46497), .B(n5648), .X(n21343) );
  nand_x1_sg U75006 ( .A(n5554), .B(n20142), .X(n20304) );
  nor_x1_sg U75007 ( .A(n20142), .B(n5554), .X(n20305) );
  nand_x1_sg U75008 ( .A(n5647), .B(n46539), .X(n21365) );
  nor_x1_sg U75009 ( .A(n46539), .B(n5647), .X(n21366) );
  nand_x1_sg U75010 ( .A(n5500), .B(n46304), .X(n19895) );
  nor_x1_sg U75011 ( .A(n46304), .B(n5500), .X(n19896) );
  nand_x1_sg U75012 ( .A(n5501), .B(n46259), .X(n19890) );
  nor_x1_sg U75013 ( .A(n46259), .B(n5501), .X(n19891) );
  nand_x1_sg U75014 ( .A(n5502), .B(n46213), .X(n19885) );
  nor_x1_sg U75015 ( .A(n46213), .B(n5502), .X(n19886) );
  nand_x1_sg U75016 ( .A(n5503), .B(n46168), .X(n19880) );
  nor_x1_sg U75017 ( .A(n46168), .B(n5503), .X(n19881) );
  nand_x1_sg U75018 ( .A(n5504), .B(n46122), .X(n19875) );
  nor_x1_sg U75019 ( .A(n46122), .B(n5504), .X(n19876) );
  nand_x1_sg U75020 ( .A(n5505), .B(n46077), .X(n19870) );
  nor_x1_sg U75021 ( .A(n46077), .B(n5505), .X(n19871) );
  nand_x1_sg U75022 ( .A(n5506), .B(n46031), .X(n19865) );
  nor_x1_sg U75023 ( .A(n46031), .B(n5506), .X(n19866) );
  nand_x1_sg U75024 ( .A(n5507), .B(n45986), .X(n19860) );
  nor_x1_sg U75025 ( .A(n45986), .B(n5507), .X(n19861) );
  nand_x1_sg U75026 ( .A(n5508), .B(n45941), .X(n19855) );
  nor_x1_sg U75027 ( .A(n45941), .B(n5508), .X(n19856) );
  nand_x1_sg U75028 ( .A(n5490), .B(n45891), .X(n19643) );
  nor_x1_sg U75029 ( .A(n45891), .B(n5490), .X(n19644) );
  nand_x1_sg U75030 ( .A(n5570), .B(n19748), .X(n19747) );
  nor_x1_sg U75031 ( .A(n19748), .B(n5570), .X(n19749) );
  nand_x1_sg U75032 ( .A(n5461), .B(n19480), .X(n19479) );
  nor_x1_sg U75033 ( .A(n19480), .B(n5461), .X(n19481) );
  nand_x1_sg U75034 ( .A(n5424), .B(n46295), .X(n6267) );
  nor_x1_sg U75035 ( .A(n46295), .B(n5424), .X(n6268) );
  nand_x1_sg U75036 ( .A(n5425), .B(n46250), .X(n6312) );
  nor_x1_sg U75037 ( .A(n46250), .B(n5425), .X(n6313) );
  nand_x1_sg U75038 ( .A(n5426), .B(n46204), .X(n6356) );
  nor_x1_sg U75039 ( .A(n46204), .B(n5426), .X(n6357) );
  nand_x1_sg U75040 ( .A(n5427), .B(n46159), .X(n6401) );
  nor_x1_sg U75041 ( .A(n46159), .B(n5427), .X(n6402) );
  nand_x1_sg U75042 ( .A(n5428), .B(n46113), .X(n6445) );
  nor_x1_sg U75043 ( .A(n46113), .B(n5428), .X(n6446) );
  nand_x1_sg U75044 ( .A(n5429), .B(n46068), .X(n6490) );
  nor_x1_sg U75045 ( .A(n46068), .B(n5429), .X(n6491) );
  nand_x1_sg U75046 ( .A(n5430), .B(n46022), .X(n6534) );
  nor_x1_sg U75047 ( .A(n46022), .B(n5430), .X(n6535) );
  nand_x1_sg U75048 ( .A(n5431), .B(n45977), .X(n6579) );
  nor_x1_sg U75049 ( .A(n45977), .B(n5431), .X(n6580) );
  nand_x1_sg U75050 ( .A(n5432), .B(n45932), .X(n6623) );
  nor_x1_sg U75051 ( .A(n45932), .B(n5432), .X(n6624) );
  nand_x1_sg U75052 ( .A(n5434), .B(n6715), .X(n6714) );
  nor_x1_sg U75053 ( .A(n6715), .B(n5434), .X(n6716) );
  nand_x1_sg U75054 ( .A(n38762), .B(n47138), .X(n23121) );
  nor_x1_sg U75055 ( .A(n47138), .B(\reg_yHat[1][2] ), .X(n23122) );
  nand_x1_sg U75056 ( .A(n38766), .B(n47423), .X(n23401) );
  nor_x1_sg U75057 ( .A(n47423), .B(\reg_yHat[2][2] ), .X(n23402) );
  nand_x1_sg U75058 ( .A(n38770), .B(n47708), .X(n23680) );
  nor_x1_sg U75059 ( .A(n47708), .B(\reg_yHat[3][2] ), .X(n23681) );
  nand_x1_sg U75060 ( .A(n38774), .B(n47993), .X(n23959) );
  nor_x1_sg U75061 ( .A(n47993), .B(\reg_yHat[4][2] ), .X(n23960) );
  nand_x1_sg U75062 ( .A(n38778), .B(n48278), .X(n24238) );
  nor_x1_sg U75063 ( .A(n48278), .B(\reg_yHat[5][2] ), .X(n24239) );
  nand_x1_sg U75064 ( .A(n38782), .B(n48563), .X(n24517) );
  nor_x1_sg U75065 ( .A(n48563), .B(\reg_yHat[6][2] ), .X(n24518) );
  nand_x1_sg U75066 ( .A(n38786), .B(n48848), .X(n24795) );
  nor_x1_sg U75067 ( .A(n48848), .B(\reg_yHat[7][2] ), .X(n24796) );
  nand_x1_sg U75068 ( .A(n38790), .B(n49135), .X(n25074) );
  nor_x1_sg U75069 ( .A(n49135), .B(\reg_yHat[8][2] ), .X(n25075) );
  nand_x1_sg U75070 ( .A(n38794), .B(n49421), .X(n25353) );
  nor_x1_sg U75071 ( .A(n49421), .B(\reg_yHat[9][2] ), .X(n25354) );
  nand_x1_sg U75072 ( .A(n38798), .B(n49707), .X(n25632) );
  nor_x1_sg U75073 ( .A(n49707), .B(\reg_yHat[10][2] ), .X(n25633) );
  nand_x1_sg U75074 ( .A(n38802), .B(n49993), .X(n25909) );
  nor_x1_sg U75075 ( .A(n49993), .B(\reg_yHat[11][2] ), .X(n25910) );
  nand_x1_sg U75076 ( .A(n38806), .B(n50568), .X(n26469) );
  nor_x1_sg U75077 ( .A(n50568), .B(\reg_yHat[13][2] ), .X(n26470) );
  nand_x1_sg U75078 ( .A(n38810), .B(n50854), .X(n26747) );
  nor_x1_sg U75079 ( .A(n50854), .B(\reg_yHat[14][2] ), .X(n26748) );
  nand_x1_sg U75080 ( .A(n38758), .B(n42215), .X(n22844) );
  nor_x1_sg U75081 ( .A(n42215), .B(\reg_yHat[0][2] ), .X(n22845) );
  nand_x1_sg U75082 ( .A(\reg_yHat[12][3] ), .B(n50284), .X(n26115) );
  nand_x1_sg U75083 ( .A(\reg_y[12][3] ), .B(n42015), .X(n26116) );
  inv_x1_sg U75084 ( .A(\reg_y[12][3] ), .X(n50284) );
  nand_x1_sg U75085 ( .A(\reg_y[0][1] ), .B(n46633), .X(n22850) );
  nand_x1_sg U75086 ( .A(\reg_yHat[0][1] ), .B(n46842), .X(n22849) );
  nand_x1_sg U75087 ( .A(\reg_y[1][1] ), .B(n46646), .X(n23128) );
  nand_x1_sg U75088 ( .A(\reg_yHat[1][1] ), .B(n47135), .X(n23127) );
  nand_x1_sg U75089 ( .A(\reg_y[2][1] ), .B(n46660), .X(n23408) );
  nand_x1_sg U75090 ( .A(\reg_yHat[2][1] ), .B(n47420), .X(n23407) );
  nand_x1_sg U75091 ( .A(\reg_y[3][1] ), .B(n46674), .X(n23687) );
  nand_x1_sg U75092 ( .A(\reg_yHat[3][1] ), .B(n47705), .X(n23686) );
  nand_x1_sg U75093 ( .A(\reg_y[4][1] ), .B(n46688), .X(n23966) );
  nand_x1_sg U75094 ( .A(\reg_yHat[4][1] ), .B(n47990), .X(n23965) );
  nand_x1_sg U75095 ( .A(\reg_y[5][1] ), .B(n46702), .X(n24245) );
  nand_x1_sg U75096 ( .A(\reg_yHat[5][1] ), .B(n48275), .X(n24244) );
  nand_x1_sg U75097 ( .A(\reg_y[6][1] ), .B(n46716), .X(n24524) );
  nand_x1_sg U75098 ( .A(\reg_yHat[6][1] ), .B(n48560), .X(n24523) );
  nand_x1_sg U75099 ( .A(\reg_y[7][1] ), .B(n46730), .X(n24802) );
  nand_x1_sg U75100 ( .A(\reg_yHat[7][1] ), .B(n48845), .X(n24801) );
  nand_x1_sg U75101 ( .A(\reg_y[8][1] ), .B(n46744), .X(n25081) );
  nand_x1_sg U75102 ( .A(\reg_yHat[8][1] ), .B(n49132), .X(n25080) );
  nand_x1_sg U75103 ( .A(\reg_y[9][1] ), .B(n46758), .X(n25360) );
  nand_x1_sg U75104 ( .A(\reg_yHat[9][1] ), .B(n49418), .X(n25359) );
  nand_x1_sg U75105 ( .A(\reg_y[10][1] ), .B(n46772), .X(n25639) );
  nand_x1_sg U75106 ( .A(\reg_yHat[10][1] ), .B(n49704), .X(n25638) );
  nand_x1_sg U75107 ( .A(\reg_y[11][1] ), .B(n46786), .X(n25916) );
  nand_x1_sg U75108 ( .A(\reg_yHat[11][1] ), .B(n49990), .X(n25915) );
  nand_x1_sg U75109 ( .A(\reg_y[12][1] ), .B(n46800), .X(n26127) );
  nand_x1_sg U75110 ( .A(\reg_yHat[12][1] ), .B(n50276), .X(n26126) );
  nand_x1_sg U75111 ( .A(\reg_y[14][1] ), .B(n46827), .X(n26754) );
  nand_x1_sg U75112 ( .A(\reg_yHat[14][1] ), .B(n50851), .X(n26753) );
  nand_x1_sg U75113 ( .A(\reg_y[13][1] ), .B(n46813), .X(n26476) );
  nand_x1_sg U75114 ( .A(\reg_yHat[13][1] ), .B(n50563), .X(n26475) );
  nand_x1_sg U75115 ( .A(n5622), .B(n45955), .X(n20866) );
  nand_x1_sg U75116 ( .A(n20867), .B(n38236), .X(n20865) );
  nand_x1_sg U75117 ( .A(n5546), .B(n45946), .X(n20223) );
  nand_x1_sg U75118 ( .A(n20224), .B(n38237), .X(n20222) );
  nand_x1_sg U75119 ( .A(n5470), .B(n45937), .X(n19417) );
  nand_x1_sg U75120 ( .A(n19418), .B(n38238), .X(n19416) );
  nand_x1_sg U75121 ( .A(n5266), .B(n45710), .X(n27101) );
  nand_x1_sg U75122 ( .A(n26850), .B(n38239), .X(n27100) );
  nand_x1_sg U75123 ( .A(n42339), .B(n20777), .X(n20790) );
  nor_x1_sg U75124 ( .A(n20792), .B(n5590), .X(n20791) );
  nand_x1_sg U75125 ( .A(n21186), .B(n42113), .X(n21183) );
  nand_x1_sg U75126 ( .A(n28741), .B(n42118), .X(n28738) );
  nand_x2_sg U75127 ( .A(n5703), .B(n38561), .X(n21588) );
  nand_x2_sg U75128 ( .A(n5718), .B(n38562), .X(n29139) );
  nand_x1_sg U75129 ( .A(n45826), .B(n38528), .X(n20853) );
  nand_x1_sg U75130 ( .A(n5624), .B(n20855), .X(n20854) );
  nand_x1_sg U75131 ( .A(n45842), .B(n38529), .X(n20210) );
  nand_x1_sg U75132 ( .A(n5548), .B(n20212), .X(n20211) );
  nand_x1_sg U75133 ( .A(n46445), .B(n38530), .X(n19914) );
  nand_x1_sg U75134 ( .A(n5497), .B(n19916), .X(n19915) );
  nand_x1_sg U75135 ( .A(n45858), .B(n38531), .X(n19404) );
  nand_x1_sg U75136 ( .A(n5472), .B(n19406), .X(n19405) );
  nand_x1_sg U75137 ( .A(\reg_yHat[12][5] ), .B(n50300), .X(n26103) );
  nand_x1_sg U75138 ( .A(\reg_y[12][5] ), .B(n46802), .X(n26104) );
  nand_x1_sg U75139 ( .A(n46360), .B(n38240), .X(n20928) );
  nand_x1_sg U75140 ( .A(n46318), .B(n38241), .X(n20921) );
  nand_x1_sg U75141 ( .A(n46273), .B(n38242), .X(n20914) );
  nand_x1_sg U75142 ( .A(n46227), .B(n38243), .X(n20907) );
  nand_x1_sg U75143 ( .A(n46182), .B(n38244), .X(n20900) );
  nand_x1_sg U75144 ( .A(n46136), .B(n38245), .X(n20893) );
  nand_x1_sg U75145 ( .A(n46091), .B(n38246), .X(n20886) );
  nand_x1_sg U75146 ( .A(n46045), .B(n38247), .X(n20879) );
  nand_x1_sg U75147 ( .A(n46000), .B(n38248), .X(n20872) );
  nand_x1_sg U75148 ( .A(n46407), .B(n38249), .X(n20935) );
  nand_x1_sg U75149 ( .A(n46455), .B(n38250), .X(n20942) );
  nand_x1_sg U75150 ( .A(n46493), .B(n38251), .X(n20949) );
  nand_x1_sg U75151 ( .A(n46309), .B(n38252), .X(n20278) );
  nand_x1_sg U75152 ( .A(n46264), .B(n38253), .X(n20271) );
  nand_x1_sg U75153 ( .A(n46218), .B(n38254), .X(n20264) );
  nand_x1_sg U75154 ( .A(n46173), .B(n38255), .X(n20257) );
  nand_x1_sg U75155 ( .A(n46127), .B(n38256), .X(n20250) );
  nand_x1_sg U75156 ( .A(n46082), .B(n38257), .X(n20243) );
  nand_x1_sg U75157 ( .A(n46036), .B(n38258), .X(n20236) );
  nand_x1_sg U75158 ( .A(n45991), .B(n38259), .X(n20229) );
  nand_x1_sg U75159 ( .A(n46300), .B(n38260), .X(n19472) );
  nand_x1_sg U75160 ( .A(n46255), .B(n38261), .X(n19465) );
  nand_x1_sg U75161 ( .A(n46209), .B(n38262), .X(n19458) );
  nand_x1_sg U75162 ( .A(n46164), .B(n38263), .X(n19451) );
  nand_x1_sg U75163 ( .A(n46118), .B(n38264), .X(n19444) );
  nand_x1_sg U75164 ( .A(n46073), .B(n38265), .X(n19437) );
  nand_x1_sg U75165 ( .A(n46027), .B(n38266), .X(n19430) );
  nand_x1_sg U75166 ( .A(n45982), .B(n38267), .X(n19423) );
  nand_x1_sg U75167 ( .A(n5662), .B(n21270), .X(n21269) );
  nor_x1_sg U75168 ( .A(n21270), .B(n5662), .X(n21271) );
  nand_x1_sg U75169 ( .A(n5555), .B(n20309), .X(n20446) );
  nor_x1_sg U75170 ( .A(n20309), .B(n5555), .X(n20447) );
  nand_x1_sg U75171 ( .A(n5586), .B(n20501), .X(n20500) );
  nor_x1_sg U75172 ( .A(n20501), .B(n5586), .X(n20502) );
  nand_x1_sg U75173 ( .A(n5510), .B(n19844), .X(n19843) );
  nor_x1_sg U75174 ( .A(n19844), .B(n5510), .X(n19845) );
  nand_x1_sg U75175 ( .A(n5280), .B(n45103), .X(n28146) );
  nor_x1_sg U75176 ( .A(n45103), .B(n5280), .X(n28147) );
  nand_x1_sg U75177 ( .A(n5279), .B(n45149), .X(n28151) );
  nor_x1_sg U75178 ( .A(n45149), .B(n5279), .X(n28152) );
  nand_x1_sg U75179 ( .A(n5278), .B(n45194), .X(n28156) );
  nor_x1_sg U75180 ( .A(n45194), .B(n5278), .X(n28157) );
  nand_x1_sg U75181 ( .A(n5277), .B(n45240), .X(n28161) );
  nor_x1_sg U75182 ( .A(n45240), .B(n5277), .X(n28162) );
  nand_x1_sg U75183 ( .A(n5276), .B(n45285), .X(n28166) );
  nor_x1_sg U75184 ( .A(n45285), .B(n5276), .X(n28167) );
  nand_x1_sg U75185 ( .A(n5275), .B(n45330), .X(n28171) );
  nor_x1_sg U75186 ( .A(n45330), .B(n5275), .X(n28172) );
  nand_x1_sg U75187 ( .A(n5274), .B(n45375), .X(n28176) );
  nor_x1_sg U75188 ( .A(n45375), .B(n5274), .X(n28177) );
  nand_x1_sg U75189 ( .A(n5273), .B(n45421), .X(n28182) );
  nor_x1_sg U75190 ( .A(n45421), .B(n5273), .X(n28183) );
  nand_x1_sg U75191 ( .A(n5272), .B(n45465), .X(n28211) );
  nor_x1_sg U75192 ( .A(n45465), .B(n5272), .X(n28212) );
  nand_x1_sg U75193 ( .A(n5271), .B(n45489), .X(n28076) );
  nor_x1_sg U75194 ( .A(n45489), .B(n5271), .X(n28077) );
  nand_x1_sg U75195 ( .A(n5270), .B(n45533), .X(n27914) );
  nor_x1_sg U75196 ( .A(n45533), .B(n5270), .X(n27915) );
  nand_x1_sg U75197 ( .A(n5269), .B(n45578), .X(n27737) );
  nor_x1_sg U75198 ( .A(n45578), .B(n5269), .X(n27738) );
  nand_x1_sg U75199 ( .A(n5623), .B(n45908), .X(n20859) );
  nor_x1_sg U75200 ( .A(n45908), .B(n5623), .X(n20860) );
  nand_x1_sg U75201 ( .A(n5268), .B(n45622), .X(n27543) );
  nor_x1_sg U75202 ( .A(n45622), .B(n5268), .X(n27544) );
  nand_x1_sg U75203 ( .A(n5574), .B(n46402), .X(n20444) );
  nor_x1_sg U75204 ( .A(n46402), .B(n5574), .X(n20445) );
  nand_x1_sg U75205 ( .A(n5267), .B(n45666), .X(n27330) );
  nor_x1_sg U75206 ( .A(n45666), .B(n5267), .X(n27331) );
  nand_x1_sg U75207 ( .A(n5573), .B(n46450), .X(n20302) );
  nor_x1_sg U75208 ( .A(n46450), .B(n5573), .X(n20303) );
  nand_x1_sg U75209 ( .A(n5547), .B(n45898), .X(n20216) );
  nor_x1_sg U75210 ( .A(n45898), .B(n5547), .X(n20217) );
  nand_x1_sg U75211 ( .A(n5479), .B(n46393), .X(n19708) );
  nor_x1_sg U75212 ( .A(n46393), .B(n5479), .X(n19709) );
  nand_x1_sg U75213 ( .A(n5478), .B(n46442), .X(n19714) );
  nor_x1_sg U75214 ( .A(n46442), .B(n5478), .X(n19715) );
  nand_x1_sg U75215 ( .A(n5471), .B(n45888), .X(n19410) );
  nor_x1_sg U75216 ( .A(n45888), .B(n5471), .X(n19411) );
  nand_x1_sg U75217 ( .A(\reg_y[12][2] ), .B(n42002), .X(n26121) );
  nor_x1_sg U75218 ( .A(n42002), .B(\reg_y[12][2] ), .X(n26122) );
  nand_x1_sg U75219 ( .A(n19761), .B(n38268), .X(n19946) );
  inv_x1_sg U75220 ( .A(n19761), .X(n46513) );
  nand_x1_sg U75221 ( .A(n19145), .B(n38269), .X(n19338) );
  inv_x1_sg U75222 ( .A(n19145), .X(n46574) );
  nand_x1_sg U75223 ( .A(n19311), .B(n38532), .X(n19309) );
  inv_x1_sg U75224 ( .A(n19311), .X(n46389) );
  nand_x1_sg U75225 ( .A(n21005), .B(n38270), .X(n21202) );
  inv_x1_sg U75226 ( .A(n21005), .X(n46581) );
  nand_x1_sg U75227 ( .A(n19337), .B(n38271), .X(n19335) );
  inv_x1_sg U75228 ( .A(n19337), .X(n46575) );
  nand_x1_sg U75229 ( .A(n5513), .B(n46562), .X(n19763) );
  nand_x1_sg U75230 ( .A(n19550), .B(n38272), .X(n19762) );
  nand_x1_sg U75231 ( .A(n5494), .B(n46565), .X(n19769) );
  nand_x1_sg U75232 ( .A(n19557), .B(n38273), .X(n19768) );
  nand_x1_sg U75233 ( .A(n5608), .B(n46580), .X(n20785) );
  nand_x1_sg U75234 ( .A(n20786), .B(n38274), .X(n20784) );
  nand_x1_sg U75235 ( .A(n5532), .B(n46560), .X(n19757) );
  nand_x1_sg U75236 ( .A(n19543), .B(n38275), .X(n19756) );
  nand_x1_sg U75237 ( .A(n5551), .B(n46558), .X(n19751) );
  nand_x1_sg U75238 ( .A(n19536), .B(n38276), .X(n19750) );
  nand_x1_sg U75239 ( .A(n5475), .B(n46576), .X(n19775) );
  nand_x1_sg U75240 ( .A(n19564), .B(n38277), .X(n19774) );
  nand_x1_sg U75241 ( .A(n5418), .B(n46572), .X(n5982) );
  nand_x1_sg U75242 ( .A(n5983), .B(n38278), .X(n5981) );
  nand_x1_sg U75243 ( .A(n5498), .B(n46396), .X(n19908) );
  nand_x1_sg U75244 ( .A(n5458), .B(n46483), .X(n19499) );
  nand_x1_sg U75245 ( .A(n19746), .B(n19748), .X(n20592) );
  nor_x1_sg U75246 ( .A(n20594), .B(n5570), .X(n20593) );
  nand_x1_sg U75247 ( .A(n46535), .B(n38533), .X(n20955) );
  nand_x1_sg U75248 ( .A(n46351), .B(n38534), .X(n20284) );
  nand_x1_sg U75249 ( .A(n46578), .B(n38279), .X(n20787) );
  nand_x1_sg U75250 ( .A(n46343), .B(n38535), .X(n19303) );
  nand_x1_sg U75251 ( .A(n46347), .B(n38536), .X(n19702) );
  nand_x1_sg U75252 ( .A(n20982), .B(n38189), .X(n20979) );
  nand_x1_sg U75253 ( .A(n28540), .B(n38190), .X(n28537) );
  nand_x1_sg U75254 ( .A(n46474), .B(n38537), .X(n20144) );
  nand_x1_sg U75255 ( .A(n5534), .B(n19951), .X(n20145) );
  nand_x1_sg U75256 ( .A(n46516), .B(n38538), .X(n19952) );
  nand_x1_sg U75257 ( .A(n5514), .B(n19767), .X(n19953) );
  nand_x1_sg U75258 ( .A(n45020), .B(n38280), .X(n22511) );
  nand_x1_sg U75259 ( .A(n44994), .B(n38281), .X(n28265) );
  nand_x1_sg U75260 ( .A(n45060), .B(n38282), .X(n28271) );
  nand_x1_sg U75261 ( .A(n45001), .B(n38283), .X(n27982) );
  nand_x1_sg U75262 ( .A(n45106), .B(n38284), .X(n28277) );
  nand_x1_sg U75263 ( .A(n45004), .B(n38285), .X(n27812) );
  nand_x1_sg U75264 ( .A(n45152), .B(n38286), .X(n28283) );
  nand_x1_sg U75265 ( .A(n45007), .B(n38287), .X(n27626) );
  nand_x1_sg U75266 ( .A(n45056), .B(n38288), .X(n27818) );
  nand_x1_sg U75267 ( .A(n44985), .B(n38289), .X(n28633) );
  nand_x1_sg U75268 ( .A(n45010), .B(n38290), .X(n27423) );
  nand_x1_sg U75269 ( .A(n45057), .B(n38291), .X(n27989) );
  nand_x1_sg U75270 ( .A(n45101), .B(n38292), .X(n27995) );
  nand_x1_sg U75271 ( .A(n45197), .B(n38293), .X(n28289) );
  nand_x1_sg U75272 ( .A(n45055), .B(n38294), .X(n27632) );
  nand_x1_sg U75273 ( .A(n45100), .B(n38295), .X(n27824) );
  nand_x1_sg U75274 ( .A(n45148), .B(n38296), .X(n28001) );
  nand_x1_sg U75275 ( .A(n45243), .B(n38297), .X(n28295) );
  nand_x1_sg U75276 ( .A(n44988), .B(n38298), .X(n28472) );
  nand_x1_sg U75277 ( .A(n45063), .B(n38299), .X(n28639) );
  nand_x1_sg U75278 ( .A(n44979), .B(n38300), .X(n28992) );
  nand_x1_sg U75279 ( .A(n45013), .B(n38301), .X(n27201) );
  nand_x1_sg U75280 ( .A(n45054), .B(n38302), .X(n27429) );
  nand_x1_sg U75281 ( .A(n45099), .B(n38303), .X(n27638) );
  nand_x1_sg U75282 ( .A(n45147), .B(n38304), .X(n27830) );
  nand_x1_sg U75283 ( .A(n45193), .B(n38305), .X(n28007) );
  nand_x1_sg U75284 ( .A(n45288), .B(n38306), .X(n28301) );
  nand_x1_sg U75285 ( .A(n45062), .B(n38307), .X(n28478) );
  nand_x1_sg U75286 ( .A(n45109), .B(n38308), .X(n28645) );
  nand_x1_sg U75287 ( .A(n45065), .B(n38309), .X(n28999) );
  nand_x1_sg U75288 ( .A(n45053), .B(n38310), .X(n27207) );
  nand_x1_sg U75289 ( .A(n45098), .B(n38311), .X(n27435) );
  nand_x1_sg U75290 ( .A(n45146), .B(n38312), .X(n27644) );
  nand_x1_sg U75291 ( .A(n45192), .B(n38313), .X(n27836) );
  nand_x1_sg U75292 ( .A(n45239), .B(n38314), .X(n28013) );
  nand_x1_sg U75293 ( .A(n45333), .B(n38315), .X(n28307) );
  nand_x1_sg U75294 ( .A(n45108), .B(n38316), .X(n28484) );
  nand_x1_sg U75295 ( .A(n45155), .B(n38317), .X(n28651) );
  nand_x1_sg U75296 ( .A(n45111), .B(n38318), .X(n29005) );
  nand_x1_sg U75297 ( .A(n45097), .B(n38319), .X(n27213) );
  nand_x1_sg U75298 ( .A(n45145), .B(n38320), .X(n27441) );
  nand_x1_sg U75299 ( .A(n45191), .B(n38321), .X(n27650) );
  nand_x1_sg U75300 ( .A(n45238), .B(n38322), .X(n27842) );
  nand_x1_sg U75301 ( .A(n45284), .B(n38323), .X(n28019) );
  nand_x1_sg U75302 ( .A(n45378), .B(n38324), .X(n28313) );
  nand_x1_sg U75303 ( .A(n45154), .B(n38325), .X(n28490) );
  nand_x1_sg U75304 ( .A(n45200), .B(n38326), .X(n28657) );
  nand_x1_sg U75305 ( .A(n45157), .B(n38327), .X(n29012) );
  nand_x1_sg U75306 ( .A(n45144), .B(n38328), .X(n27219) );
  nand_x1_sg U75307 ( .A(n45190), .B(n38329), .X(n27447) );
  nand_x1_sg U75308 ( .A(n45237), .B(n38330), .X(n27656) );
  nand_x1_sg U75309 ( .A(n45283), .B(n38331), .X(n27848) );
  nand_x1_sg U75310 ( .A(n45329), .B(n38332), .X(n28025) );
  nand_x1_sg U75311 ( .A(n45424), .B(n38333), .X(n28334) );
  nand_x1_sg U75312 ( .A(n45199), .B(n38334), .X(n28496) );
  nand_x1_sg U75313 ( .A(n45246), .B(n38335), .X(n28663) );
  nand_x1_sg U75314 ( .A(n45202), .B(n38336), .X(n29018) );
  nand_x1_sg U75315 ( .A(n45189), .B(n38337), .X(n27225) );
  nand_x1_sg U75316 ( .A(n45236), .B(n38338), .X(n27453) );
  nand_x1_sg U75317 ( .A(n45282), .B(n38339), .X(n27662) );
  nand_x1_sg U75318 ( .A(n45328), .B(n38340), .X(n27854) );
  nand_x1_sg U75319 ( .A(n45374), .B(n38341), .X(n28031) );
  nand_x1_sg U75320 ( .A(n45468), .B(n38342), .X(n28205) );
  nand_x1_sg U75321 ( .A(n45245), .B(n38343), .X(n28502) );
  nand_x1_sg U75322 ( .A(n45291), .B(n38344), .X(n28669) );
  nand_x1_sg U75323 ( .A(n45248), .B(n38345), .X(n29025) );
  nand_x1_sg U75324 ( .A(n45235), .B(n38346), .X(n27231) );
  nand_x1_sg U75325 ( .A(n45281), .B(n38347), .X(n27459) );
  nand_x1_sg U75326 ( .A(n45327), .B(n38348), .X(n27668) );
  nand_x1_sg U75327 ( .A(n45373), .B(n38349), .X(n27860) );
  nand_x1_sg U75328 ( .A(n45420), .B(n38350), .X(n28037) );
  nand_x1_sg U75329 ( .A(n45513), .B(n38351), .X(n28070) );
  nand_x1_sg U75330 ( .A(n45290), .B(n38352), .X(n28508) );
  nand_x1_sg U75331 ( .A(n45336), .B(n38353), .X(n28675) );
  nand_x1_sg U75332 ( .A(n45293), .B(n38354), .X(n29031) );
  nand_x1_sg U75333 ( .A(n45280), .B(n38355), .X(n27237) );
  nand_x1_sg U75334 ( .A(n45326), .B(n38356), .X(n27465) );
  nand_x1_sg U75335 ( .A(n45372), .B(n38357), .X(n27674) );
  nand_x1_sg U75336 ( .A(n45419), .B(n38358), .X(n27866) );
  nand_x1_sg U75337 ( .A(n45464), .B(n38359), .X(n28043) );
  nand_x1_sg U75338 ( .A(n45557), .B(n38360), .X(n27908) );
  nand_x1_sg U75339 ( .A(n45335), .B(n38361), .X(n28514) );
  nand_x1_sg U75340 ( .A(n45381), .B(n38362), .X(n28681) );
  nand_x1_sg U75341 ( .A(n45338), .B(n38363), .X(n29038) );
  nand_x1_sg U75342 ( .A(n45325), .B(n38364), .X(n27243) );
  nand_x1_sg U75343 ( .A(n45371), .B(n38365), .X(n27471) );
  nand_x1_sg U75344 ( .A(n45418), .B(n38366), .X(n27680) );
  nand_x1_sg U75345 ( .A(n45463), .B(n38367), .X(n27872) );
  nand_x1_sg U75346 ( .A(n45512), .B(n38368), .X(n28083) );
  nand_x1_sg U75347 ( .A(n45602), .B(n38369), .X(n27731) );
  nand_x1_sg U75348 ( .A(n45380), .B(n38370), .X(n28429) );
  nand_x1_sg U75349 ( .A(n45427), .B(n38371), .X(n28687) );
  nand_x1_sg U75350 ( .A(n45383), .B(n38372), .X(n29044) );
  nand_x1_sg U75351 ( .A(n45370), .B(n38373), .X(n27249) );
  nand_x1_sg U75352 ( .A(n45417), .B(n38374), .X(n27477) );
  nand_x1_sg U75353 ( .A(n45462), .B(n38375), .X(n27686) );
  nand_x1_sg U75354 ( .A(n45511), .B(n38376), .X(n27878) );
  nand_x1_sg U75355 ( .A(n45556), .B(n38377), .X(n27921) );
  nand_x1_sg U75356 ( .A(n45646), .B(n38378), .X(n27537) );
  nand_x1_sg U75357 ( .A(n45426), .B(n38379), .X(n28325) );
  nand_x1_sg U75358 ( .A(n45471), .B(n38380), .X(n28693) );
  nand_x1_sg U75359 ( .A(n45429), .B(n38381), .X(n29051) );
  nand_x1_sg U75360 ( .A(n45416), .B(n38382), .X(n27255) );
  nand_x1_sg U75361 ( .A(n45461), .B(n38383), .X(n27483) );
  nand_x1_sg U75362 ( .A(n45510), .B(n38384), .X(n27692) );
  nand_x1_sg U75363 ( .A(n45555), .B(n38385), .X(n27927) );
  nand_x1_sg U75364 ( .A(n45601), .B(n38386), .X(n27744) );
  nand_x1_sg U75365 ( .A(n45690), .B(n38387), .X(n27324) );
  nand_x1_sg U75366 ( .A(n45470), .B(n38388), .X(n28196) );
  nand_x1_sg U75367 ( .A(n45516), .B(n38389), .X(n28699) );
  nand_x1_sg U75368 ( .A(n45473), .B(n38390), .X(n29057) );
  nand_x1_sg U75369 ( .A(n45460), .B(n38391), .X(n27261) );
  nand_x1_sg U75370 ( .A(n45509), .B(n38392), .X(n27489) );
  nand_x1_sg U75371 ( .A(n45554), .B(n38393), .X(n27698) );
  nand_x1_sg U75372 ( .A(n45600), .B(n38394), .X(n27750) );
  nand_x1_sg U75373 ( .A(n45645), .B(n38395), .X(n27550) );
  nand_x1_sg U75374 ( .A(n45733), .B(n38396), .X(n27094) );
  nand_x1_sg U75375 ( .A(n45515), .B(n38397), .X(n28061) );
  nand_x1_sg U75376 ( .A(n45560), .B(n38398), .X(n28705) );
  nand_x1_sg U75377 ( .A(n45518), .B(n38399), .X(n29064) );
  nand_x1_sg U75378 ( .A(n45508), .B(n38400), .X(n27267) );
  nand_x1_sg U75379 ( .A(n45553), .B(n38401), .X(n27495) );
  nand_x1_sg U75380 ( .A(n45599), .B(n38402), .X(n27756) );
  nand_x1_sg U75381 ( .A(n45644), .B(n38403), .X(n27556) );
  nand_x1_sg U75382 ( .A(n45689), .B(n38404), .X(n27337) );
  nand_x1_sg U75383 ( .A(n45559), .B(n38405), .X(n27899) );
  nand_x1_sg U75384 ( .A(n45605), .B(n38406), .X(n28711) );
  nand_x1_sg U75385 ( .A(n45562), .B(n38407), .X(n29070) );
  nand_x1_sg U75386 ( .A(n45552), .B(n38408), .X(n27273) );
  nand_x1_sg U75387 ( .A(n45598), .B(n38409), .X(n27501) );
  nand_x1_sg U75388 ( .A(n45643), .B(n38410), .X(n27562) );
  nand_x1_sg U75389 ( .A(n45688), .B(n38411), .X(n27343) );
  nand_x1_sg U75390 ( .A(n45732), .B(n38412), .X(n27107) );
  nand_x1_sg U75391 ( .A(n46500), .B(n38413), .X(n21541) );
  nand_x1_sg U75392 ( .A(n45604), .B(n38414), .X(n27722) );
  nand_x1_sg U75393 ( .A(n45649), .B(n38415), .X(n28717) );
  nand_x1_sg U75394 ( .A(n45607), .B(n38416), .X(n29077) );
  nand_x1_sg U75395 ( .A(n45597), .B(n38417), .X(n27279) );
  nand_x1_sg U75396 ( .A(n45642), .B(n38418), .X(n27568) );
  nand_x1_sg U75397 ( .A(n45687), .B(n38419), .X(n27349) );
  nand_x1_sg U75398 ( .A(n45731), .B(n38420), .X(n27113) );
  nand_x1_sg U75399 ( .A(n46542), .B(n38421), .X(n21359) );
  nand_x1_sg U75400 ( .A(n45648), .B(n38422), .X(n27528) );
  nand_x1_sg U75401 ( .A(n45693), .B(n38423), .X(n28723) );
  nand_x1_sg U75402 ( .A(n45651), .B(n38424), .X(n29092) );
  nand_x1_sg U75403 ( .A(n45641), .B(n38425), .X(n27285) );
  nand_x1_sg U75404 ( .A(n45686), .B(n38426), .X(n27355) );
  nand_x1_sg U75405 ( .A(n45730), .B(n38427), .X(n27119) );
  nand_x1_sg U75406 ( .A(n45815), .B(n38428), .X(n21441) );
  nand_x1_sg U75407 ( .A(n45692), .B(n38429), .X(n27315) );
  nand_x1_sg U75408 ( .A(n45736), .B(n38430), .X(n28756) );
  nand_x1_sg U75409 ( .A(n45695), .B(n38431), .X(n28923) );
  nand_x1_sg U75410 ( .A(n45685), .B(n38432), .X(n27361) );
  nand_x1_sg U75411 ( .A(n45729), .B(n38433), .X(n27125) );
  nand_x1_sg U75412 ( .A(n46582), .B(n38434), .X(n21189) );
  nand_x1_sg U75413 ( .A(n45735), .B(n38435), .X(n27085) );
  nand_x1_sg U75414 ( .A(n45738), .B(n38436), .X(n28744) );
  nand_x1_sg U75415 ( .A(n45728), .B(n38437), .X(n27131) );
  nand_x1_sg U75416 ( .A(n46391), .B(n38438), .X(n19485) );
  nand_x1_sg U75417 ( .A(n45916), .B(n38439), .X(n21448) );
  nand_x1_sg U75418 ( .A(n46480), .B(n38440), .X(n6082) );
  nand_x1_sg U75419 ( .A(n46462), .B(n38441), .X(n21526) );
  nand_x1_sg U75420 ( .A(n46414), .B(n38442), .X(n21519) );
  nand_x1_sg U75421 ( .A(n46367), .B(n38443), .X(n21513) );
  nand_x1_sg U75422 ( .A(n46325), .B(n38444), .X(n21506) );
  nand_x1_sg U75423 ( .A(n46280), .B(n38445), .X(n21500) );
  nand_x1_sg U75424 ( .A(n46234), .B(n38446), .X(n21493) );
  nand_x1_sg U75425 ( .A(n46189), .B(n38447), .X(n21487) );
  nand_x1_sg U75426 ( .A(n46143), .B(n38448), .X(n21480) );
  nand_x1_sg U75427 ( .A(n46098), .B(n38449), .X(n21474) );
  nand_x1_sg U75428 ( .A(n46052), .B(n38450), .X(n21467) );
  nand_x1_sg U75429 ( .A(n46007), .B(n38451), .X(n21461) );
  nand_x1_sg U75430 ( .A(n45962), .B(n38452), .X(n21454) );
  nand_x1_sg U75431 ( .A(n45734), .B(n38453), .X(n27088) );
  nand_x1_sg U75432 ( .A(n45737), .B(n38454), .X(n28750) );
  nand_x1_sg U75433 ( .A(n45726), .B(n38455), .X(n21760) );
  nand_x1_sg U75434 ( .A(n45727), .B(n38456), .X(n27137) );
  nand_x1_sg U75435 ( .A(n45691), .B(n38457), .X(n27318) );
  nand_x1_sg U75436 ( .A(n45694), .B(n38458), .X(n28929) );
  nand_x1_sg U75437 ( .A(n45683), .B(n38459), .X(n21807) );
  nand_x1_sg U75438 ( .A(n45684), .B(n38460), .X(n27052) );
  nand_x1_sg U75439 ( .A(n45647), .B(n38461), .X(n27531) );
  nand_x1_sg U75440 ( .A(n45650), .B(n38462), .X(n28905) );
  nand_x1_sg U75441 ( .A(n45639), .B(n38463), .X(n21854) );
  nand_x1_sg U75442 ( .A(n45640), .B(n38464), .X(n27046) );
  nand_x1_sg U75443 ( .A(n45603), .B(n38465), .X(n27725) );
  nand_x1_sg U75444 ( .A(n45606), .B(n38466), .X(n28899) );
  nand_x1_sg U75445 ( .A(n45595), .B(n38467), .X(n21900) );
  nand_x1_sg U75446 ( .A(n45596), .B(n38468), .X(n27040) );
  nand_x1_sg U75447 ( .A(n45558), .B(n38469), .X(n27902) );
  nand_x1_sg U75448 ( .A(n45561), .B(n38470), .X(n28893) );
  nand_x1_sg U75449 ( .A(n45550), .B(n38471), .X(n21947) );
  nand_x1_sg U75450 ( .A(n45551), .B(n38472), .X(n27034) );
  nand_x1_sg U75451 ( .A(n45514), .B(n38473), .X(n28064) );
  nand_x1_sg U75452 ( .A(n45517), .B(n38474), .X(n28887) );
  nand_x1_sg U75453 ( .A(n45506), .B(n38475), .X(n21993) );
  nand_x1_sg U75454 ( .A(n45507), .B(n38476), .X(n27028) );
  nand_x1_sg U75455 ( .A(n45469), .B(n38477), .X(n28199) );
  nand_x1_sg U75456 ( .A(n45472), .B(n38478), .X(n28881) );
  nand_x1_sg U75457 ( .A(n45458), .B(n38479), .X(n22040) );
  nand_x1_sg U75458 ( .A(n45459), .B(n38480), .X(n27022) );
  nand_x1_sg U75459 ( .A(n45425), .B(n38481), .X(n28328) );
  nand_x1_sg U75460 ( .A(n45428), .B(n38482), .X(n28875) );
  nand_x1_sg U75461 ( .A(n45414), .B(n38483), .X(n22086) );
  nand_x1_sg U75462 ( .A(n45415), .B(n38484), .X(n27016) );
  nand_x1_sg U75463 ( .A(n45379), .B(n38485), .X(n28432) );
  nand_x1_sg U75464 ( .A(n45382), .B(n38486), .X(n28869) );
  nand_x1_sg U75465 ( .A(n45368), .B(n38487), .X(n22134) );
  nand_x1_sg U75466 ( .A(n45369), .B(n38488), .X(n27010) );
  nand_x1_sg U75467 ( .A(n45334), .B(n38489), .X(n28420) );
  nand_x1_sg U75468 ( .A(n45337), .B(n38490), .X(n28863) );
  nand_x1_sg U75469 ( .A(n45323), .B(n38491), .X(n22181) );
  nand_x1_sg U75470 ( .A(n45324), .B(n38492), .X(n27004) );
  nand_x1_sg U75471 ( .A(n45289), .B(n38493), .X(n28414) );
  nand_x1_sg U75472 ( .A(n45292), .B(n38494), .X(n28857) );
  nand_x1_sg U75473 ( .A(n45278), .B(n38495), .X(n22229) );
  nand_x1_sg U75474 ( .A(n45279), .B(n38496), .X(n26998) );
  nand_x1_sg U75475 ( .A(n45244), .B(n38497), .X(n28408) );
  nand_x1_sg U75476 ( .A(n45247), .B(n38498), .X(n28851) );
  nand_x1_sg U75477 ( .A(n45233), .B(n38499), .X(n22276) );
  nand_x1_sg U75478 ( .A(n45234), .B(n38500), .X(n26992) );
  nand_x1_sg U75479 ( .A(n45198), .B(n38501), .X(n28402) );
  nand_x1_sg U75480 ( .A(n45201), .B(n38502), .X(n28845) );
  nand_x1_sg U75481 ( .A(n45187), .B(n38503), .X(n22324) );
  nand_x1_sg U75482 ( .A(n45188), .B(n38504), .X(n26986) );
  nand_x1_sg U75483 ( .A(n45153), .B(n38505), .X(n28396) );
  nand_x1_sg U75484 ( .A(n45156), .B(n38506), .X(n28839) );
  nand_x1_sg U75485 ( .A(n45142), .B(n38507), .X(n22371) );
  nand_x1_sg U75486 ( .A(n45143), .B(n38508), .X(n26980) );
  nand_x1_sg U75487 ( .A(n45107), .B(n38509), .X(n28390) );
  nand_x1_sg U75488 ( .A(n45110), .B(n38510), .X(n28833) );
  nand_x1_sg U75489 ( .A(n45095), .B(n38511), .X(n22419) );
  nand_x1_sg U75490 ( .A(n45096), .B(n38512), .X(n26974) );
  nand_x1_sg U75491 ( .A(n45061), .B(n38513), .X(n28384) );
  nand_x1_sg U75492 ( .A(n45064), .B(n38514), .X(n28827) );
  nand_x1_sg U75493 ( .A(n45051), .B(n38515), .X(n22465) );
  nand_x1_sg U75494 ( .A(n45052), .B(n38516), .X(n26968) );
  nand_x1_sg U75495 ( .A(n44991), .B(n38517), .X(n28378) );
  nand_x1_sg U75496 ( .A(n44982), .B(n38518), .X(n28821) );
  nand_x1_sg U75497 ( .A(n45016), .B(n38519), .X(n26962) );
  nor_x1_sg U75498 ( .A(n20108), .B(n5518), .X(n20109) );
  nor_x1_sg U75499 ( .A(n6034), .B(n5419), .X(n6035) );
  nor_x1_sg U75500 ( .A(n6175), .B(n5422), .X(n6176) );
  nor_x1_sg U75501 ( .A(n38121), .B(out_L1[10]), .X(n29199) );
  nor_x1_sg U75502 ( .A(n38122), .B(out_L1[12]), .X(n29211) );
  nor_x1_sg U75503 ( .A(n38123), .B(out_L2[14]), .X(n21672) );
  nor_x1_sg U75504 ( .A(n38124), .B(out_L1[14]), .X(n29223) );
  nor_x1_sg U75505 ( .A(n38125), .B(out_L2[16]), .X(n21540) );
  nor_x1_sg U75506 ( .A(n38126), .B(out_L1[16]), .X(n29091) );
  nand_x1_sg U75507 ( .A(n5553), .B(n19944), .X(n20137) );
  nor_x1_sg U75508 ( .A(n19944), .B(n5553), .X(n20138) );
  nand_x1_sg U75509 ( .A(n5571), .B(n19938), .X(n19937) );
  nor_x1_sg U75510 ( .A(n19938), .B(n5571), .X(n19939) );
  nand_x1_sg U75511 ( .A(n5438), .B(n46526), .X(n19326) );
  nor_x1_sg U75512 ( .A(n46526), .B(n5438), .X(n19327) );
  nand_x1_sg U75513 ( .A(n5439), .B(n46481), .X(n19320) );
  nor_x1_sg U75514 ( .A(n46481), .B(n5439), .X(n19321) );
  nor_x1_sg U75515 ( .A(n26845), .B(n5265), .X(n26846) );
  nor_x1_sg U75516 ( .A(n19545), .B(n5512), .X(n19546) );
  nor_x1_sg U75517 ( .A(n19552), .B(n5493), .X(n19553) );
  nor_x1_sg U75518 ( .A(n19559), .B(n5474), .X(n19560) );
  nand_x1_sg U75519 ( .A(n5588), .B(n20584), .X(n20583) );
  nor_x1_sg U75520 ( .A(n20584), .B(n5588), .X(n20585) );
  nand_x1_sg U75521 ( .A(n5455), .B(n19566), .X(n19565) );
  nor_x1_sg U75522 ( .A(n19566), .B(n5455), .X(n19567) );
  nand_x1_sg U75523 ( .A(n5569), .B(n20590), .X(n20589) );
  nor_x1_sg U75524 ( .A(n20590), .B(n5569), .X(n20591) );
  nand_x1_sg U75525 ( .A(n5436), .B(n19141), .X(n19140) );
  nor_x1_sg U75526 ( .A(n19141), .B(n5436), .X(n19142) );
  nor_x1_sg U75527 ( .A(n19531), .B(n5550), .X(n19532) );
  nand_x1_sg U75528 ( .A(n5626), .B(n21001), .X(n21000) );
  nor_x1_sg U75529 ( .A(n21001), .B(n5626), .X(n21002) );
  nor_x1_sg U75530 ( .A(n19148), .B(n5417), .X(n19149) );
  nor_x1_sg U75531 ( .A(n19538), .B(n5531), .X(n19539) );
  nor_x1_sg U75532 ( .A(n20993), .B(n5645), .X(n20994) );
  nor_x1_sg U75533 ( .A(n21008), .B(n5607), .X(n21009) );
  nand_x1_sg U75534 ( .A(n5702), .B(n6802), .X(n6804) );
  nand_x1_sg U75535 ( .A(n41251), .B(n22591), .X(n22590) );
  nand_x1_sg U75536 ( .A(n5717), .B(n41124), .X(n22591) );
endmodule

