
module post_sparsity ( clk, reset, .i_im({\i_im[15][19] , \i_im[15][18] , 
        \i_im[15][17] , \i_im[15][16] , \i_im[15][15] , \i_im[15][14] , 
        \i_im[15][13] , \i_im[15][12] , \i_im[15][11] , \i_im[15][10] , 
        \i_im[15][9] , \i_im[15][8] , \i_im[15][7] , \i_im[15][6] , 
        \i_im[15][5] , \i_im[15][4] , \i_im[15][3] , \i_im[15][2] , 
        \i_im[15][1] , \i_im[15][0] , \i_im[14][19] , \i_im[14][18] , 
        \i_im[14][17] , \i_im[14][16] , \i_im[14][15] , \i_im[14][14] , 
        \i_im[14][13] , \i_im[14][12] , \i_im[14][11] , \i_im[14][10] , 
        \i_im[14][9] , \i_im[14][8] , \i_im[14][7] , \i_im[14][6] , 
        \i_im[14][5] , \i_im[14][4] , \i_im[14][3] , \i_im[14][2] , 
        \i_im[14][1] , \i_im[14][0] , \i_im[13][19] , \i_im[13][18] , 
        \i_im[13][17] , \i_im[13][16] , \i_im[13][15] , \i_im[13][14] , 
        \i_im[13][13] , \i_im[13][12] , \i_im[13][11] , \i_im[13][10] , 
        \i_im[13][9] , \i_im[13][8] , \i_im[13][7] , \i_im[13][6] , 
        \i_im[13][5] , \i_im[13][4] , \i_im[13][3] , \i_im[13][2] , 
        \i_im[13][1] , \i_im[13][0] , \i_im[12][19] , \i_im[12][18] , 
        \i_im[12][17] , \i_im[12][16] , \i_im[12][15] , \i_im[12][14] , 
        \i_im[12][13] , \i_im[12][12] , \i_im[12][11] , \i_im[12][10] , 
        \i_im[12][9] , \i_im[12][8] , \i_im[12][7] , \i_im[12][6] , 
        \i_im[12][5] , \i_im[12][4] , \i_im[12][3] , \i_im[12][2] , 
        \i_im[12][1] , \i_im[12][0] , \i_im[11][19] , \i_im[11][18] , 
        \i_im[11][17] , \i_im[11][16] , \i_im[11][15] , \i_im[11][14] , 
        \i_im[11][13] , \i_im[11][12] , \i_im[11][11] , \i_im[11][10] , 
        \i_im[11][9] , \i_im[11][8] , \i_im[11][7] , \i_im[11][6] , 
        \i_im[11][5] , \i_im[11][4] , \i_im[11][3] , \i_im[11][2] , 
        \i_im[11][1] , \i_im[11][0] , \i_im[10][19] , \i_im[10][18] , 
        \i_im[10][17] , \i_im[10][16] , \i_im[10][15] , \i_im[10][14] , 
        \i_im[10][13] , \i_im[10][12] , \i_im[10][11] , \i_im[10][10] , 
        \i_im[10][9] , \i_im[10][8] , \i_im[10][7] , \i_im[10][6] , 
        \i_im[10][5] , \i_im[10][4] , \i_im[10][3] , \i_im[10][2] , 
        \i_im[10][1] , \i_im[10][0] , \i_im[9][19] , \i_im[9][18] , 
        \i_im[9][17] , \i_im[9][16] , \i_im[9][15] , \i_im[9][14] , 
        \i_im[9][13] , \i_im[9][12] , \i_im[9][11] , \i_im[9][10] , 
        \i_im[9][9] , \i_im[9][8] , \i_im[9][7] , \i_im[9][6] , \i_im[9][5] , 
        \i_im[9][4] , \i_im[9][3] , \i_im[9][2] , \i_im[9][1] , \i_im[9][0] , 
        \i_im[8][19] , \i_im[8][18] , \i_im[8][17] , \i_im[8][16] , 
        \i_im[8][15] , \i_im[8][14] , \i_im[8][13] , \i_im[8][12] , 
        \i_im[8][11] , \i_im[8][10] , \i_im[8][9] , \i_im[8][8] , \i_im[8][7] , 
        \i_im[8][6] , \i_im[8][5] , \i_im[8][4] , \i_im[8][3] , \i_im[8][2] , 
        \i_im[8][1] , \i_im[8][0] , \i_im[7][19] , \i_im[7][18] , 
        \i_im[7][17] , \i_im[7][16] , \i_im[7][15] , \i_im[7][14] , 
        \i_im[7][13] , \i_im[7][12] , \i_im[7][11] , \i_im[7][10] , 
        \i_im[7][9] , \i_im[7][8] , \i_im[7][7] , \i_im[7][6] , \i_im[7][5] , 
        \i_im[7][4] , \i_im[7][3] , \i_im[7][2] , \i_im[7][1] , \i_im[7][0] , 
        \i_im[6][19] , \i_im[6][18] , \i_im[6][17] , \i_im[6][16] , 
        \i_im[6][15] , \i_im[6][14] , \i_im[6][13] , \i_im[6][12] , 
        \i_im[6][11] , \i_im[6][10] , \i_im[6][9] , \i_im[6][8] , \i_im[6][7] , 
        \i_im[6][6] , \i_im[6][5] , \i_im[6][4] , \i_im[6][3] , \i_im[6][2] , 
        \i_im[6][1] , \i_im[6][0] , \i_im[5][19] , \i_im[5][18] , 
        \i_im[5][17] , \i_im[5][16] , \i_im[5][15] , \i_im[5][14] , 
        \i_im[5][13] , \i_im[5][12] , \i_im[5][11] , \i_im[5][10] , 
        \i_im[5][9] , \i_im[5][8] , \i_im[5][7] , \i_im[5][6] , \i_im[5][5] , 
        \i_im[5][4] , \i_im[5][3] , \i_im[5][2] , \i_im[5][1] , \i_im[5][0] , 
        \i_im[4][19] , \i_im[4][18] , \i_im[4][17] , \i_im[4][16] , 
        \i_im[4][15] , \i_im[4][14] , \i_im[4][13] , \i_im[4][12] , 
        \i_im[4][11] , \i_im[4][10] , \i_im[4][9] , \i_im[4][8] , \i_im[4][7] , 
        \i_im[4][6] , \i_im[4][5] , \i_im[4][4] , \i_im[4][3] , \i_im[4][2] , 
        \i_im[4][1] , \i_im[4][0] , \i_im[3][19] , \i_im[3][18] , 
        \i_im[3][17] , \i_im[3][16] , \i_im[3][15] , \i_im[3][14] , 
        \i_im[3][13] , \i_im[3][12] , \i_im[3][11] , \i_im[3][10] , 
        \i_im[3][9] , \i_im[3][8] , \i_im[3][7] , \i_im[3][6] , \i_im[3][5] , 
        \i_im[3][4] , \i_im[3][3] , \i_im[3][2] , \i_im[3][1] , \i_im[3][0] , 
        \i_im[2][19] , \i_im[2][18] , \i_im[2][17] , \i_im[2][16] , 
        \i_im[2][15] , \i_im[2][14] , \i_im[2][13] , \i_im[2][12] , 
        \i_im[2][11] , \i_im[2][10] , \i_im[2][9] , \i_im[2][8] , \i_im[2][7] , 
        \i_im[2][6] , \i_im[2][5] , \i_im[2][4] , \i_im[2][3] , \i_im[2][2] , 
        \i_im[2][1] , \i_im[2][0] , \i_im[1][19] , \i_im[1][18] , 
        \i_im[1][17] , \i_im[1][16] , \i_im[1][15] , \i_im[1][14] , 
        \i_im[1][13] , \i_im[1][12] , \i_im[1][11] , \i_im[1][10] , 
        \i_im[1][9] , \i_im[1][8] , \i_im[1][7] , \i_im[1][6] , \i_im[1][5] , 
        \i_im[1][4] , \i_im[1][3] , \i_im[1][2] , \i_im[1][1] , \i_im[1][0] , 
        \i_im[0][19] , \i_im[0][18] , \i_im[0][17] , \i_im[0][16] , 
        \i_im[0][15] , \i_im[0][14] , \i_im[0][13] , \i_im[0][12] , 
        \i_im[0][11] , \i_im[0][10] , \i_im[0][9] , \i_im[0][8] , \i_im[0][7] , 
        \i_im[0][6] , \i_im[0][5] , \i_im[0][4] , \i_im[0][3] , \i_im[0][2] , 
        \i_im[0][1] , \i_im[0][0] }), i_mask, input_ready, output_taken, 
    .o_im({\o_im[15][19] , \o_im[15][18] , \o_im[15][17] , \o_im[15][16] , 
        \o_im[15][15] , \o_im[15][14] , \o_im[15][13] , \o_im[15][12] , 
        \o_im[15][11] , \o_im[15][10] , \o_im[15][9] , \o_im[15][8] , 
        \o_im[15][7] , \o_im[15][6] , \o_im[15][5] , \o_im[15][4] , 
        \o_im[15][3] , \o_im[15][2] , \o_im[15][1] , \o_im[15][0] , 
        \o_im[14][19] , \o_im[14][18] , \o_im[14][17] , \o_im[14][16] , 
        \o_im[14][15] , \o_im[14][14] , \o_im[14][13] , \o_im[14][12] , 
        \o_im[14][11] , \o_im[14][10] , \o_im[14][9] , \o_im[14][8] , 
        \o_im[14][7] , \o_im[14][6] , \o_im[14][5] , \o_im[14][4] , 
        \o_im[14][3] , \o_im[14][2] , \o_im[14][1] , \o_im[14][0] , 
        \o_im[13][19] , \o_im[13][18] , \o_im[13][17] , \o_im[13][16] , 
        \o_im[13][15] , \o_im[13][14] , \o_im[13][13] , \o_im[13][12] , 
        \o_im[13][11] , \o_im[13][10] , \o_im[13][9] , \o_im[13][8] , 
        \o_im[13][7] , \o_im[13][6] , \o_im[13][5] , \o_im[13][4] , 
        \o_im[13][3] , \o_im[13][2] , \o_im[13][1] , \o_im[13][0] , 
        \o_im[12][19] , \o_im[12][18] , \o_im[12][17] , \o_im[12][16] , 
        \o_im[12][15] , \o_im[12][14] , \o_im[12][13] , \o_im[12][12] , 
        \o_im[12][11] , \o_im[12][10] , \o_im[12][9] , \o_im[12][8] , 
        \o_im[12][7] , \o_im[12][6] , \o_im[12][5] , \o_im[12][4] , 
        \o_im[12][3] , \o_im[12][2] , \o_im[12][1] , \o_im[12][0] , 
        \o_im[11][19] , \o_im[11][18] , \o_im[11][17] , \o_im[11][16] , 
        \o_im[11][15] , \o_im[11][14] , \o_im[11][13] , \o_im[11][12] , 
        \o_im[11][11] , \o_im[11][10] , \o_im[11][9] , \o_im[11][8] , 
        \o_im[11][7] , \o_im[11][6] , \o_im[11][5] , \o_im[11][4] , 
        \o_im[11][3] , \o_im[11][2] , \o_im[11][1] , \o_im[11][0] , 
        \o_im[10][19] , \o_im[10][18] , \o_im[10][17] , \o_im[10][16] , 
        \o_im[10][15] , \o_im[10][14] , \o_im[10][13] , \o_im[10][12] , 
        \o_im[10][11] , \o_im[10][10] , \o_im[10][9] , \o_im[10][8] , 
        \o_im[10][7] , \o_im[10][6] , \o_im[10][5] , \o_im[10][4] , 
        \o_im[10][3] , \o_im[10][2] , \o_im[10][1] , \o_im[10][0] , 
        \o_im[9][19] , \o_im[9][18] , \o_im[9][17] , \o_im[9][16] , 
        \o_im[9][15] , \o_im[9][14] , \o_im[9][13] , \o_im[9][12] , 
        \o_im[9][11] , \o_im[9][10] , \o_im[9][9] , \o_im[9][8] , \o_im[9][7] , 
        \o_im[9][6] , \o_im[9][5] , \o_im[9][4] , \o_im[9][3] , \o_im[9][2] , 
        \o_im[9][1] , \o_im[9][0] , \o_im[8][19] , \o_im[8][18] , 
        \o_im[8][17] , \o_im[8][16] , \o_im[8][15] , \o_im[8][14] , 
        \o_im[8][13] , \o_im[8][12] , \o_im[8][11] , \o_im[8][10] , 
        \o_im[8][9] , \o_im[8][8] , \o_im[8][7] , \o_im[8][6] , \o_im[8][5] , 
        \o_im[8][4] , \o_im[8][3] , \o_im[8][2] , \o_im[8][1] , \o_im[8][0] , 
        \o_im[7][19] , \o_im[7][18] , \o_im[7][17] , \o_im[7][16] , 
        \o_im[7][15] , \o_im[7][14] , \o_im[7][13] , \o_im[7][12] , 
        \o_im[7][11] , \o_im[7][10] , \o_im[7][9] , \o_im[7][8] , \o_im[7][7] , 
        \o_im[7][6] , \o_im[7][5] , \o_im[7][4] , \o_im[7][3] , \o_im[7][2] , 
        \o_im[7][1] , \o_im[7][0] , \o_im[6][19] , \o_im[6][18] , 
        \o_im[6][17] , \o_im[6][16] , \o_im[6][15] , \o_im[6][14] , 
        \o_im[6][13] , \o_im[6][12] , \o_im[6][11] , \o_im[6][10] , 
        \o_im[6][9] , \o_im[6][8] , \o_im[6][7] , \o_im[6][6] , \o_im[6][5] , 
        \o_im[6][4] , \o_im[6][3] , \o_im[6][2] , \o_im[6][1] , \o_im[6][0] , 
        \o_im[5][19] , \o_im[5][18] , \o_im[5][17] , \o_im[5][16] , 
        \o_im[5][15] , \o_im[5][14] , \o_im[5][13] , \o_im[5][12] , 
        \o_im[5][11] , \o_im[5][10] , \o_im[5][9] , \o_im[5][8] , \o_im[5][7] , 
        \o_im[5][6] , \o_im[5][5] , \o_im[5][4] , \o_im[5][3] , \o_im[5][2] , 
        \o_im[5][1] , \o_im[5][0] , \o_im[4][19] , \o_im[4][18] , 
        \o_im[4][17] , \o_im[4][16] , \o_im[4][15] , \o_im[4][14] , 
        \o_im[4][13] , \o_im[4][12] , \o_im[4][11] , \o_im[4][10] , 
        \o_im[4][9] , \o_im[4][8] , \o_im[4][7] , \o_im[4][6] , \o_im[4][5] , 
        \o_im[4][4] , \o_im[4][3] , \o_im[4][2] , \o_im[4][1] , \o_im[4][0] , 
        \o_im[3][19] , \o_im[3][18] , \o_im[3][17] , \o_im[3][16] , 
        \o_im[3][15] , \o_im[3][14] , \o_im[3][13] , \o_im[3][12] , 
        \o_im[3][11] , \o_im[3][10] , \o_im[3][9] , \o_im[3][8] , \o_im[3][7] , 
        \o_im[3][6] , \o_im[3][5] , \o_im[3][4] , \o_im[3][3] , \o_im[3][2] , 
        \o_im[3][1] , \o_im[3][0] , \o_im[2][19] , \o_im[2][18] , 
        \o_im[2][17] , \o_im[2][16] , \o_im[2][15] , \o_im[2][14] , 
        \o_im[2][13] , \o_im[2][12] , \o_im[2][11] , \o_im[2][10] , 
        \o_im[2][9] , \o_im[2][8] , \o_im[2][7] , \o_im[2][6] , \o_im[2][5] , 
        \o_im[2][4] , \o_im[2][3] , \o_im[2][2] , \o_im[2][1] , \o_im[2][0] , 
        \o_im[1][19] , \o_im[1][18] , \o_im[1][17] , \o_im[1][16] , 
        \o_im[1][15] , \o_im[1][14] , \o_im[1][13] , \o_im[1][12] , 
        \o_im[1][11] , \o_im[1][10] , \o_im[1][9] , \o_im[1][8] , \o_im[1][7] , 
        \o_im[1][6] , \o_im[1][5] , \o_im[1][4] , \o_im[1][3] , \o_im[1][2] , 
        \o_im[1][1] , \o_im[1][0] , \o_im[0][19] , \o_im[0][18] , 
        \o_im[0][17] , \o_im[0][16] , \o_im[0][15] , \o_im[0][14] , 
        \o_im[0][13] , \o_im[0][12] , \o_im[0][11] , \o_im[0][10] , 
        \o_im[0][9] , \o_im[0][8] , \o_im[0][7] , \o_im[0][6] , \o_im[0][5] , 
        \o_im[0][4] , \o_im[0][3] , \o_im[0][2] , \o_im[0][1] , \o_im[0][0] }), 
        o_mask, state );
  input [31:0] i_mask;
  output [31:0] o_mask;
  output [1:0] state;
  input clk, reset, \i_im[15][19] , \i_im[15][18] , \i_im[15][17] ,
         \i_im[15][16] , \i_im[15][15] , \i_im[15][14] , \i_im[15][13] ,
         \i_im[15][12] , \i_im[15][11] , \i_im[15][10] , \i_im[15][9] ,
         \i_im[15][8] , \i_im[15][7] , \i_im[15][6] , \i_im[15][5] ,
         \i_im[15][4] , \i_im[15][3] , \i_im[15][2] , \i_im[15][1] ,
         \i_im[15][0] , \i_im[14][19] , \i_im[14][18] , \i_im[14][17] ,
         \i_im[14][16] , \i_im[14][15] , \i_im[14][14] , \i_im[14][13] ,
         \i_im[14][12] , \i_im[14][11] , \i_im[14][10] , \i_im[14][9] ,
         \i_im[14][8] , \i_im[14][7] , \i_im[14][6] , \i_im[14][5] ,
         \i_im[14][4] , \i_im[14][3] , \i_im[14][2] , \i_im[14][1] ,
         \i_im[14][0] , \i_im[13][19] , \i_im[13][18] , \i_im[13][17] ,
         \i_im[13][16] , \i_im[13][15] , \i_im[13][14] , \i_im[13][13] ,
         \i_im[13][12] , \i_im[13][11] , \i_im[13][10] , \i_im[13][9] ,
         \i_im[13][8] , \i_im[13][7] , \i_im[13][6] , \i_im[13][5] ,
         \i_im[13][4] , \i_im[13][3] , \i_im[13][2] , \i_im[13][1] ,
         \i_im[13][0] , \i_im[12][19] , \i_im[12][18] , \i_im[12][17] ,
         \i_im[12][16] , \i_im[12][15] , \i_im[12][14] , \i_im[12][13] ,
         \i_im[12][12] , \i_im[12][11] , \i_im[12][10] , \i_im[12][9] ,
         \i_im[12][8] , \i_im[12][7] , \i_im[12][6] , \i_im[12][5] ,
         \i_im[12][4] , \i_im[12][3] , \i_im[12][2] , \i_im[12][1] ,
         \i_im[12][0] , \i_im[11][19] , \i_im[11][18] , \i_im[11][17] ,
         \i_im[11][16] , \i_im[11][15] , \i_im[11][14] , \i_im[11][13] ,
         \i_im[11][12] , \i_im[11][11] , \i_im[11][10] , \i_im[11][9] ,
         \i_im[11][8] , \i_im[11][7] , \i_im[11][6] , \i_im[11][5] ,
         \i_im[11][4] , \i_im[11][3] , \i_im[11][2] , \i_im[11][1] ,
         \i_im[11][0] , \i_im[10][19] , \i_im[10][18] , \i_im[10][17] ,
         \i_im[10][16] , \i_im[10][15] , \i_im[10][14] , \i_im[10][13] ,
         \i_im[10][12] , \i_im[10][11] , \i_im[10][10] , \i_im[10][9] ,
         \i_im[10][8] , \i_im[10][7] , \i_im[10][6] , \i_im[10][5] ,
         \i_im[10][4] , \i_im[10][3] , \i_im[10][2] , \i_im[10][1] ,
         \i_im[10][0] , \i_im[9][19] , \i_im[9][18] , \i_im[9][17] ,
         \i_im[9][16] , \i_im[9][15] , \i_im[9][14] , \i_im[9][13] ,
         \i_im[9][12] , \i_im[9][11] , \i_im[9][10] , \i_im[9][9] ,
         \i_im[9][8] , \i_im[9][7] , \i_im[9][6] , \i_im[9][5] , \i_im[9][4] ,
         \i_im[9][3] , \i_im[9][2] , \i_im[9][1] , \i_im[9][0] , \i_im[8][19] ,
         \i_im[8][18] , \i_im[8][17] , \i_im[8][16] , \i_im[8][15] ,
         \i_im[8][14] , \i_im[8][13] , \i_im[8][12] , \i_im[8][11] ,
         \i_im[8][10] , \i_im[8][9] , \i_im[8][8] , \i_im[8][7] , \i_im[8][6] ,
         \i_im[8][5] , \i_im[8][4] , \i_im[8][3] , \i_im[8][2] , \i_im[8][1] ,
         \i_im[8][0] , \i_im[7][19] , \i_im[7][18] , \i_im[7][17] ,
         \i_im[7][16] , \i_im[7][15] , \i_im[7][14] , \i_im[7][13] ,
         \i_im[7][12] , \i_im[7][11] , \i_im[7][10] , \i_im[7][9] ,
         \i_im[7][8] , \i_im[7][7] , \i_im[7][6] , \i_im[7][5] , \i_im[7][4] ,
         \i_im[7][3] , \i_im[7][2] , \i_im[7][1] , \i_im[7][0] , \i_im[6][19] ,
         \i_im[6][18] , \i_im[6][17] , \i_im[6][16] , \i_im[6][15] ,
         \i_im[6][14] , \i_im[6][13] , \i_im[6][12] , \i_im[6][11] ,
         \i_im[6][10] , \i_im[6][9] , \i_im[6][8] , \i_im[6][7] , \i_im[6][6] ,
         \i_im[6][5] , \i_im[6][4] , \i_im[6][3] , \i_im[6][2] , \i_im[6][1] ,
         \i_im[6][0] , \i_im[5][19] , \i_im[5][18] , \i_im[5][17] ,
         \i_im[5][16] , \i_im[5][15] , \i_im[5][14] , \i_im[5][13] ,
         \i_im[5][12] , \i_im[5][11] , \i_im[5][10] , \i_im[5][9] ,
         \i_im[5][8] , \i_im[5][7] , \i_im[5][6] , \i_im[5][5] , \i_im[5][4] ,
         \i_im[5][3] , \i_im[5][2] , \i_im[5][1] , \i_im[5][0] , \i_im[4][19] ,
         \i_im[4][18] , \i_im[4][17] , \i_im[4][16] , \i_im[4][15] ,
         \i_im[4][14] , \i_im[4][13] , \i_im[4][12] , \i_im[4][11] ,
         \i_im[4][10] , \i_im[4][9] , \i_im[4][8] , \i_im[4][7] , \i_im[4][6] ,
         \i_im[4][5] , \i_im[4][4] , \i_im[4][3] , \i_im[4][2] , \i_im[4][1] ,
         \i_im[4][0] , \i_im[3][19] , \i_im[3][18] , \i_im[3][17] ,
         \i_im[3][16] , \i_im[3][15] , \i_im[3][14] , \i_im[3][13] ,
         \i_im[3][12] , \i_im[3][11] , \i_im[3][10] , \i_im[3][9] ,
         \i_im[3][8] , \i_im[3][7] , \i_im[3][6] , \i_im[3][5] , \i_im[3][4] ,
         \i_im[3][3] , \i_im[3][2] , \i_im[3][1] , \i_im[3][0] , \i_im[2][19] ,
         \i_im[2][18] , \i_im[2][17] , \i_im[2][16] , \i_im[2][15] ,
         \i_im[2][14] , \i_im[2][13] , \i_im[2][12] , \i_im[2][11] ,
         \i_im[2][10] , \i_im[2][9] , \i_im[2][8] , \i_im[2][7] , \i_im[2][6] ,
         \i_im[2][5] , \i_im[2][4] , \i_im[2][3] , \i_im[2][2] , \i_im[2][1] ,
         \i_im[2][0] , \i_im[1][19] , \i_im[1][18] , \i_im[1][17] ,
         \i_im[1][16] , \i_im[1][15] , \i_im[1][14] , \i_im[1][13] ,
         \i_im[1][12] , \i_im[1][11] , \i_im[1][10] , \i_im[1][9] ,
         \i_im[1][8] , \i_im[1][7] , \i_im[1][6] , \i_im[1][5] , \i_im[1][4] ,
         \i_im[1][3] , \i_im[1][2] , \i_im[1][1] , \i_im[1][0] , \i_im[0][19] ,
         \i_im[0][18] , \i_im[0][17] , \i_im[0][16] , \i_im[0][15] ,
         \i_im[0][14] , \i_im[0][13] , \i_im[0][12] , \i_im[0][11] ,
         \i_im[0][10] , \i_im[0][9] , \i_im[0][8] , \i_im[0][7] , \i_im[0][6] ,
         \i_im[0][5] , \i_im[0][4] , \i_im[0][3] , \i_im[0][2] , \i_im[0][1] ,
         \i_im[0][0] , input_ready, output_taken;
  output \o_im[15][19] , \o_im[15][18] , \o_im[15][17] , \o_im[15][16] ,
         \o_im[15][15] , \o_im[15][14] , \o_im[15][13] , \o_im[15][12] ,
         \o_im[15][11] , \o_im[15][10] , \o_im[15][9] , \o_im[15][8] ,
         \o_im[15][7] , \o_im[15][6] , \o_im[15][5] , \o_im[15][4] ,
         \o_im[15][3] , \o_im[15][2] , \o_im[15][1] , \o_im[15][0] ,
         \o_im[14][19] , \o_im[14][18] , \o_im[14][17] , \o_im[14][16] ,
         \o_im[14][15] , \o_im[14][14] , \o_im[14][13] , \o_im[14][12] ,
         \o_im[14][11] , \o_im[14][10] , \o_im[14][9] , \o_im[14][8] ,
         \o_im[14][7] , \o_im[14][6] , \o_im[14][5] , \o_im[14][4] ,
         \o_im[14][3] , \o_im[14][2] , \o_im[14][1] , \o_im[14][0] ,
         \o_im[13][19] , \o_im[13][18] , \o_im[13][17] , \o_im[13][16] ,
         \o_im[13][15] , \o_im[13][14] , \o_im[13][13] , \o_im[13][12] ,
         \o_im[13][11] , \o_im[13][10] , \o_im[13][9] , \o_im[13][8] ,
         \o_im[13][7] , \o_im[13][6] , \o_im[13][5] , \o_im[13][4] ,
         \o_im[13][3] , \o_im[13][2] , \o_im[13][1] , \o_im[13][0] ,
         \o_im[12][19] , \o_im[12][18] , \o_im[12][17] , \o_im[12][16] ,
         \o_im[12][15] , \o_im[12][14] , \o_im[12][13] , \o_im[12][12] ,
         \o_im[12][11] , \o_im[12][10] , \o_im[12][9] , \o_im[12][8] ,
         \o_im[12][7] , \o_im[12][6] , \o_im[12][5] , \o_im[12][4] ,
         \o_im[12][3] , \o_im[12][2] , \o_im[12][1] , \o_im[12][0] ,
         \o_im[11][19] , \o_im[11][18] , \o_im[11][17] , \o_im[11][16] ,
         \o_im[11][15] , \o_im[11][14] , \o_im[11][13] , \o_im[11][12] ,
         \o_im[11][11] , \o_im[11][10] , \o_im[11][9] , \o_im[11][8] ,
         \o_im[11][7] , \o_im[11][6] , \o_im[11][5] , \o_im[11][4] ,
         \o_im[11][3] , \o_im[11][2] , \o_im[11][1] , \o_im[11][0] ,
         \o_im[10][19] , \o_im[10][18] , \o_im[10][17] , \o_im[10][16] ,
         \o_im[10][15] , \o_im[10][14] , \o_im[10][13] , \o_im[10][12] ,
         \o_im[10][11] , \o_im[10][10] , \o_im[10][9] , \o_im[10][8] ,
         \o_im[10][7] , \o_im[10][6] , \o_im[10][5] , \o_im[10][4] ,
         \o_im[10][3] , \o_im[10][2] , \o_im[10][1] , \o_im[10][0] ,
         \o_im[9][19] , \o_im[9][18] , \o_im[9][17] , \o_im[9][16] ,
         \o_im[9][15] , \o_im[9][14] , \o_im[9][13] , \o_im[9][12] ,
         \o_im[9][11] , \o_im[9][10] , \o_im[9][9] , \o_im[9][8] ,
         \o_im[9][7] , \o_im[9][6] , \o_im[9][5] , \o_im[9][4] , \o_im[9][3] ,
         \o_im[9][2] , \o_im[9][1] , \o_im[9][0] , \o_im[8][19] ,
         \o_im[8][18] , \o_im[8][17] , \o_im[8][16] , \o_im[8][15] ,
         \o_im[8][14] , \o_im[8][13] , \o_im[8][12] , \o_im[8][11] ,
         \o_im[8][10] , \o_im[8][9] , \o_im[8][8] , \o_im[8][7] , \o_im[8][6] ,
         \o_im[8][5] , \o_im[8][4] , \o_im[8][3] , \o_im[8][2] , \o_im[8][1] ,
         \o_im[8][0] , \o_im[7][19] , \o_im[7][18] , \o_im[7][17] ,
         \o_im[7][16] , \o_im[7][15] , \o_im[7][14] , \o_im[7][13] ,
         \o_im[7][12] , \o_im[7][11] , \o_im[7][10] , \o_im[7][9] ,
         \o_im[7][8] , \o_im[7][7] , \o_im[7][6] , \o_im[7][5] , \o_im[7][4] ,
         \o_im[7][3] , \o_im[7][2] , \o_im[7][1] , \o_im[7][0] , \o_im[6][19] ,
         \o_im[6][18] , \o_im[6][17] , \o_im[6][16] , \o_im[6][15] ,
         \o_im[6][14] , \o_im[6][13] , \o_im[6][12] , \o_im[6][11] ,
         \o_im[6][10] , \o_im[6][9] , \o_im[6][8] , \o_im[6][7] , \o_im[6][6] ,
         \o_im[6][5] , \o_im[6][4] , \o_im[6][3] , \o_im[6][2] , \o_im[6][1] ,
         \o_im[6][0] , \o_im[5][19] , \o_im[5][18] , \o_im[5][17] ,
         \o_im[5][16] , \o_im[5][15] , \o_im[5][14] , \o_im[5][13] ,
         \o_im[5][12] , \o_im[5][11] , \o_im[5][10] , \o_im[5][9] ,
         \o_im[5][8] , \o_im[5][7] , \o_im[5][6] , \o_im[5][5] , \o_im[5][4] ,
         \o_im[5][3] , \o_im[5][2] , \o_im[5][1] , \o_im[5][0] , \o_im[4][19] ,
         \o_im[4][18] , \o_im[4][17] , \o_im[4][16] , \o_im[4][15] ,
         \o_im[4][14] , \o_im[4][13] , \o_im[4][12] , \o_im[4][11] ,
         \o_im[4][10] , \o_im[4][9] , \o_im[4][8] , \o_im[4][7] , \o_im[4][6] ,
         \o_im[4][5] , \o_im[4][4] , \o_im[4][3] , \o_im[4][2] , \o_im[4][1] ,
         \o_im[4][0] , \o_im[3][19] , \o_im[3][18] , \o_im[3][17] ,
         \o_im[3][16] , \o_im[3][15] , \o_im[3][14] , \o_im[3][13] ,
         \o_im[3][12] , \o_im[3][11] , \o_im[3][10] , \o_im[3][9] ,
         \o_im[3][8] , \o_im[3][7] , \o_im[3][6] , \o_im[3][5] , \o_im[3][4] ,
         \o_im[3][3] , \o_im[3][2] , \o_im[3][1] , \o_im[3][0] , \o_im[2][19] ,
         \o_im[2][18] , \o_im[2][17] , \o_im[2][16] , \o_im[2][15] ,
         \o_im[2][14] , \o_im[2][13] , \o_im[2][12] , \o_im[2][11] ,
         \o_im[2][10] , \o_im[2][9] , \o_im[2][8] , \o_im[2][7] , \o_im[2][6] ,
         \o_im[2][5] , \o_im[2][4] , \o_im[2][3] , \o_im[2][2] , \o_im[2][1] ,
         \o_im[2][0] , \o_im[1][19] , \o_im[1][18] , \o_im[1][17] ,
         \o_im[1][16] , \o_im[1][15] , \o_im[1][14] , \o_im[1][13] ,
         \o_im[1][12] , \o_im[1][11] , \o_im[1][10] , \o_im[1][9] ,
         \o_im[1][8] , \o_im[1][7] , \o_im[1][6] , \o_im[1][5] , \o_im[1][4] ,
         \o_im[1][3] , \o_im[1][2] , \o_im[1][1] , \o_im[1][0] , \o_im[0][19] ,
         \o_im[0][18] , \o_im[0][17] , \o_im[0][16] , \o_im[0][15] ,
         \o_im[0][14] , \o_im[0][13] , \o_im[0][12] , \o_im[0][11] ,
         \o_im[0][10] , \o_im[0][9] , \o_im[0][8] , \o_im[0][7] , \o_im[0][6] ,
         \o_im[0][5] , \o_im[0][4] , \o_im[0][3] , \o_im[0][2] , \o_im[0][1] ,
         \o_im[0][0] ;
  wire   n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257,
         n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267,
         n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277,
         n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287,
         n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297,
         n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307,
         n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317,
         n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327,
         n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337,
         n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347,
         n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357,
         n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367,
         n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377,
         n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387,
         n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397,
         n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407,
         n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417,
         n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427,
         n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437,
         n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447,
         n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457,
         n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467,
         n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477,
         n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487,
         n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497,
         n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507,
         n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517,
         n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527,
         n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537,
         n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547,
         n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557,
         n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567,
         n19, n20, n9568, n9569, \update_mask_0/n1480 , \update_mask_0/n1479 ,
         \update_mask_0/n1478 , \update_mask_0/n1477 , \update_mask_0/n1476 ,
         \update_mask_0/n1475 , \update_mask_0/n1474 , \update_mask_0/n1473 ,
         \update_mask_0/n1472 , \update_mask_0/n1471 , \update_mask_0/n1470 ,
         \update_mask_0/n1469 , \update_mask_0/n1468 , \update_mask_0/n1467 ,
         \update_mask_0/n1466 , \update_mask_0/n1465 , \update_mask_0/n1464 ,
         \update_mask_0/n1463 , \update_mask_0/n1462 , \update_mask_0/n1461 ,
         \update_mask_0/n1460 , \update_mask_0/n1459 , \update_mask_0/n1458 ,
         \update_mask_0/n1457 , \update_mask_0/n1456 , \update_mask_0/n1455 ,
         \update_mask_0/n1454 , \update_mask_0/n1453 , \update_mask_0/n1452 ,
         \update_mask_0/n1451 , \update_mask_0/n1450 , \update_mask_0/n1449 ,
         \update_mask_0/n1448 , \update_mask_0/n1447 , \update_mask_0/n1446 ,
         \update_mask_0/n1445 , \update_mask_0/n1444 , \update_mask_0/n1443 ,
         \update_mask_0/n1442 , \update_mask_0/n1441 , \update_mask_0/n1440 ,
         \update_mask_0/n1439 , \update_mask_0/n1438 , \update_mask_0/n1437 ,
         \update_mask_0/n1436 , \update_mask_0/n1435 , \update_mask_0/n1434 ,
         \update_mask_0/n1433 , \update_mask_0/n1432 , \update_mask_0/n1431 ,
         \update_mask_0/n1430 , \update_mask_0/n1429 , \update_mask_0/n1428 ,
         \update_mask_0/n1427 , \update_mask_0/n1426 , \update_mask_0/n1425 ,
         \update_mask_0/n1424 , \update_mask_0/n1423 , \update_mask_0/n1422 ,
         \update_mask_0/n1421 , \update_mask_0/n1420 , \update_mask_0/n1419 ,
         \update_mask_0/n1418 , \update_mask_0/n1417 , \update_mask_0/n1416 ,
         \update_mask_0/n1415 , \update_mask_0/n1414 , \update_mask_0/n1413 ,
         \update_mask_0/n1412 , \update_mask_0/n1411 , \update_mask_0/n1410 ,
         \update_mask_0/n1409 , \update_mask_0/n1408 , \update_mask_0/n1407 ,
         \update_mask_0/n1406 , \update_mask_0/n1405 , \update_mask_0/n1404 ,
         \update_mask_0/n1403 , \update_mask_0/n1402 , \update_mask_0/n1401 ,
         \update_mask_0/n1400 , \update_mask_0/n1399 , \update_mask_0/n1398 ,
         \update_mask_0/n1397 , \update_mask_0/n1396 , \update_mask_0/n1395 ,
         \update_mask_0/n1394 , \update_mask_0/n1393 , \update_mask_0/n1392 ,
         \update_mask_0/n1391 , \update_mask_0/n1390 , \update_mask_0/n1389 ,
         \update_mask_0/n1388 , \update_mask_0/n1387 , \update_mask_0/n1386 ,
         \update_mask_0/n1385 , \update_mask_0/n1384 , \update_mask_0/n1383 ,
         \update_mask_0/n1382 , \update_mask_0/n1381 , \update_mask_0/n1380 ,
         \update_mask_0/n1379 , \update_mask_0/n1378 , \update_mask_0/n1377 ,
         \update_mask_0/n1376 , \update_mask_0/n1375 , \update_mask_0/n1374 ,
         \update_mask_0/n1373 , \update_mask_0/n1372 , \update_mask_0/n1371 ,
         \update_mask_0/n1370 , \update_mask_0/n1369 , \update_mask_0/n1368 ,
         \update_mask_0/n1367 , \update_mask_0/n1366 , \update_mask_0/n1365 ,
         \update_mask_0/n1364 , \update_mask_0/n1363 , \update_mask_0/n1362 ,
         \update_mask_0/n1361 , \update_mask_0/n1360 , \update_mask_0/n1359 ,
         \update_mask_0/n1358 , \update_mask_0/n1357 , \update_mask_0/n1356 ,
         \update_mask_0/n1355 , \update_mask_0/n1354 , \update_mask_0/n1353 ,
         \update_mask_0/n1352 , \update_mask_0/n1351 , \update_mask_0/n1350 ,
         \update_mask_0/n1349 , \update_mask_0/n1348 , \update_mask_0/n1347 ,
         \update_mask_0/n1346 , \update_mask_0/n1345 , \update_mask_0/n1344 ,
         \update_mask_0/n1343 , \update_mask_0/n1342 , \update_mask_0/n1341 ,
         \update_mask_0/n1340 , \update_mask_0/n1339 , \update_mask_0/n1338 ,
         \update_mask_0/n1337 , \update_mask_0/n1336 , \update_mask_0/n1335 ,
         \update_mask_0/n1334 , \update_mask_0/n1333 , \update_mask_0/n1332 ,
         \update_mask_0/n1331 , \update_mask_0/n1330 , \update_mask_0/n1329 ,
         \update_mask_0/n1328 , \update_mask_0/n1327 , \update_mask_0/n1326 ,
         \update_mask_0/n1325 , \update_mask_0/n1324 , \update_mask_0/n1323 ,
         \update_mask_0/n1322 , \update_mask_0/n1321 , \update_mask_0/n1320 ,
         \update_mask_0/n1319 , \update_mask_0/n1318 , \update_mask_0/n1317 ,
         \update_mask_0/n1316 , \update_mask_0/n1315 , \update_mask_0/n1314 ,
         \update_mask_0/n1313 , \update_mask_0/n1312 , \update_mask_0/n1311 ,
         \update_mask_0/n1310 , \update_mask_0/n1309 , \update_mask_0/n1308 ,
         \update_mask_0/n1307 , \update_mask_0/n1306 , \update_mask_0/n1305 ,
         \update_mask_0/n1304 , \update_mask_0/n1303 , \update_mask_0/n1302 ,
         \update_mask_0/n1301 , \update_mask_0/n1300 , \update_mask_0/n1299 ,
         \update_mask_0/n1298 , \update_mask_0/n1297 , \update_mask_0/n1296 ,
         \update_mask_0/n1295 , \update_mask_0/n1294 , \update_mask_0/n1293 ,
         \update_mask_0/n1292 , \update_mask_0/n1291 , \update_mask_0/n1290 ,
         \update_mask_0/n1289 , \update_mask_0/n1288 , \update_mask_0/n1287 ,
         \update_mask_0/n1286 , \update_mask_0/n1285 , \update_mask_0/n1284 ,
         \update_mask_0/n1283 , \update_mask_0/n1282 , \update_mask_0/n1281 ,
         \update_mask_0/n1280 , \update_mask_0/n1279 , \update_mask_0/n1278 ,
         \update_mask_0/n1277 , \update_mask_0/n1276 , \update_mask_0/n1275 ,
         \update_mask_0/n1274 , \update_mask_0/n1273 , \update_mask_0/n1272 ,
         \update_mask_0/n1271 , \update_mask_0/n1270 , \update_mask_0/n1269 ,
         \update_mask_0/n1268 , \update_mask_0/n1267 , \update_mask_0/n1266 ,
         \update_mask_0/n1265 , \update_mask_0/n1264 , \update_mask_0/n1263 ,
         \update_mask_0/n1262 , \update_mask_0/n1261 , \update_mask_0/n1260 ,
         \update_mask_0/n1259 , \update_mask_0/n1258 , \update_mask_0/n1257 ,
         \update_mask_0/n1256 , \update_mask_0/n1255 , \update_mask_0/n1254 ,
         \update_mask_0/n1253 , \update_mask_0/n1252 , \update_mask_0/n1251 ,
         \update_mask_0/n1250 , \update_mask_0/n1249 , \update_mask_0/n1248 ,
         \update_mask_0/n1247 , \update_mask_0/n1246 , \update_mask_0/n1245 ,
         \update_mask_0/n1244 , \update_mask_0/n1243 , \update_mask_0/n1242 ,
         \update_mask_0/n1241 , \update_mask_0/n1240 , \update_mask_0/n1239 ,
         \update_mask_0/n1238 , \update_mask_0/n1237 , \update_mask_0/n1236 ,
         \update_mask_0/n1235 , \update_mask_0/n1234 , \update_mask_0/n1233 ,
         \update_mask_0/n1232 , \update_mask_0/n1231 , \update_mask_0/n1230 ,
         \update_mask_0/n1229 , \update_mask_0/n1228 , \update_mask_0/n1227 ,
         \update_mask_0/n1226 , \update_mask_0/n1225 , \update_mask_0/n1224 ,
         \update_mask_0/n1223 , \update_mask_0/n1222 , \update_mask_0/n1221 ,
         \update_mask_0/n1220 , \update_mask_0/n1219 , \update_mask_0/n1218 ,
         \update_mask_0/n1217 , \update_mask_0/n1216 , \update_mask_0/n1215 ,
         \update_mask_0/n1214 , \update_mask_0/n1213 , \update_mask_0/n1212 ,
         \update_mask_0/n1211 , \update_mask_0/n1210 , \update_mask_0/n1209 ,
         \update_mask_0/n1208 , \update_mask_0/n1207 , \update_mask_0/n1206 ,
         \update_mask_0/n1205 , \update_mask_0/n1204 , \update_mask_0/n1203 ,
         \update_mask_0/n1202 , \update_mask_0/n1201 , \update_mask_0/n1200 ,
         \update_mask_0/n1199 , \update_mask_0/n1198 , \update_mask_0/n1197 ,
         \update_mask_0/n1196 , \update_mask_0/n1195 , \update_mask_0/n1194 ,
         \update_mask_0/n1193 , \update_mask_0/n1192 , \update_mask_0/n1191 ,
         \update_mask_0/n1190 , \update_mask_0/n1189 , \update_mask_0/n1188 ,
         \update_mask_0/n1187 , \update_mask_0/n1186 , \update_mask_0/n1185 ,
         \update_mask_0/n1184 , \update_mask_0/n1183 , \update_mask_0/n1182 ,
         \update_mask_0/n1181 , \update_mask_0/n1180 , \update_mask_0/n1179 ,
         \update_mask_0/n1178 , \update_mask_0/n1177 , \update_mask_0/n1176 ,
         \update_mask_0/n1175 , \update_mask_0/n1174 , \update_mask_0/n1173 ,
         \update_mask_0/n1172 , \update_mask_0/n1171 , \update_mask_0/n1170 ,
         \update_mask_0/n1169 , \update_mask_0/n1168 , \update_mask_0/n1167 ,
         \update_mask_0/n1166 , \update_mask_0/n1165 , \update_mask_0/n1164 ,
         \update_mask_0/n1163 , \update_mask_0/n1162 , \update_mask_0/n1161 ,
         \update_mask_0/n1160 , \update_mask_0/n1159 , \update_mask_0/n1158 ,
         \update_mask_0/n1157 , \update_mask_0/n1156 , \update_mask_0/n1155 ,
         \update_mask_0/n1154 , \update_mask_0/n1153 , \update_mask_0/n1152 ,
         \update_mask_0/n1151 , \update_mask_0/n1150 , \update_mask_0/n1149 ,
         \update_mask_0/n1148 , \update_mask_0/n1147 , \update_mask_0/n1146 ,
         \update_mask_0/n1145 , \update_mask_0/n1144 , \update_mask_0/n1143 ,
         \update_mask_0/n1142 , \update_mask_0/n1141 , \update_mask_0/n1140 ,
         \update_mask_0/n1139 , \update_mask_0/n1138 , \update_mask_0/n1137 ,
         \update_mask_0/n1136 , \update_mask_0/n1135 , \update_mask_0/n1134 ,
         \update_mask_0/n1133 , \update_mask_0/n1132 , \update_mask_0/n1131 ,
         \update_mask_0/n1130 , \update_mask_0/n1129 , \update_mask_0/n1128 ,
         \update_mask_0/n1127 , \update_mask_0/n919 ,
         \update_mask_0/reg_out[15][19] , \update_mask_0/reg_out[15][18] ,
         \update_mask_0/reg_out[15][17] , \update_mask_0/reg_out[15][16] ,
         \update_mask_0/reg_out[15][15] , \update_mask_0/reg_out[15][14] ,
         \update_mask_0/reg_out[15][13] , \update_mask_0/reg_out[15][12] ,
         \update_mask_0/reg_out[15][11] , \update_mask_0/reg_out[15][10] ,
         \update_mask_0/reg_out[15][9] , \update_mask_0/reg_out[15][8] ,
         \update_mask_0/reg_out[15][7] , \update_mask_0/reg_out[15][6] ,
         \update_mask_0/reg_out[15][5] , \update_mask_0/reg_out[15][4] ,
         \update_mask_0/reg_out[15][3] , \update_mask_0/reg_out[15][2] ,
         \update_mask_0/reg_out[15][1] , \update_mask_0/reg_out[15][0] ,
         \update_mask_0/reg_out[14][19] , \update_mask_0/reg_out[14][18] ,
         \update_mask_0/reg_out[14][17] , \update_mask_0/reg_out[14][16] ,
         \update_mask_0/reg_out[14][15] , \update_mask_0/reg_out[14][14] ,
         \update_mask_0/reg_out[14][13] , \update_mask_0/reg_out[14][12] ,
         \update_mask_0/reg_out[14][11] , \update_mask_0/reg_out[14][10] ,
         \update_mask_0/reg_out[14][9] , \update_mask_0/reg_out[14][8] ,
         \update_mask_0/reg_out[14][7] , \update_mask_0/reg_out[14][6] ,
         \update_mask_0/reg_out[14][5] , \update_mask_0/reg_out[14][4] ,
         \update_mask_0/reg_out[14][3] , \update_mask_0/reg_out[14][2] ,
         \update_mask_0/reg_out[14][1] , \update_mask_0/reg_out[14][0] ,
         \update_mask_0/reg_out[13][19] , \update_mask_0/reg_out[13][18] ,
         \update_mask_0/reg_out[13][17] , \update_mask_0/reg_out[13][16] ,
         \update_mask_0/reg_out[13][15] , \update_mask_0/reg_out[13][14] ,
         \update_mask_0/reg_out[13][13] , \update_mask_0/reg_out[13][12] ,
         \update_mask_0/reg_out[13][11] , \update_mask_0/reg_out[13][10] ,
         \update_mask_0/reg_out[13][9] , \update_mask_0/reg_out[13][8] ,
         \update_mask_0/reg_out[13][7] , \update_mask_0/reg_out[13][6] ,
         \update_mask_0/reg_out[13][5] , \update_mask_0/reg_out[13][4] ,
         \update_mask_0/reg_out[13][3] , \update_mask_0/reg_out[13][2] ,
         \update_mask_0/reg_out[13][1] , \update_mask_0/reg_out[13][0] ,
         \update_mask_0/reg_out[12][19] , \update_mask_0/reg_out[12][18] ,
         \update_mask_0/reg_out[12][17] , \update_mask_0/reg_out[12][16] ,
         \update_mask_0/reg_out[12][15] , \update_mask_0/reg_out[12][14] ,
         \update_mask_0/reg_out[12][13] , \update_mask_0/reg_out[12][12] ,
         \update_mask_0/reg_out[12][11] , \update_mask_0/reg_out[12][10] ,
         \update_mask_0/reg_out[12][9] , \update_mask_0/reg_out[12][8] ,
         \update_mask_0/reg_out[12][7] , \update_mask_0/reg_out[12][6] ,
         \update_mask_0/reg_out[12][5] , \update_mask_0/reg_out[12][4] ,
         \update_mask_0/reg_out[12][3] , \update_mask_0/reg_out[12][2] ,
         \update_mask_0/reg_out[12][1] , \update_mask_0/reg_out[12][0] ,
         \update_mask_0/reg_out[11][19] , \update_mask_0/reg_out[11][18] ,
         \update_mask_0/reg_out[11][17] , \update_mask_0/reg_out[11][16] ,
         \update_mask_0/reg_out[11][15] , \update_mask_0/reg_out[11][14] ,
         \update_mask_0/reg_out[11][13] , \update_mask_0/reg_out[11][12] ,
         \update_mask_0/reg_out[11][11] , \update_mask_0/reg_out[11][10] ,
         \update_mask_0/reg_out[11][9] , \update_mask_0/reg_out[11][8] ,
         \update_mask_0/reg_out[11][7] , \update_mask_0/reg_out[11][6] ,
         \update_mask_0/reg_out[11][5] , \update_mask_0/reg_out[11][4] ,
         \update_mask_0/reg_out[11][3] , \update_mask_0/reg_out[11][2] ,
         \update_mask_0/reg_out[11][1] , \update_mask_0/reg_out[11][0] ,
         \update_mask_0/reg_out[10][19] , \update_mask_0/reg_out[10][18] ,
         \update_mask_0/reg_out[10][17] , \update_mask_0/reg_out[10][16] ,
         \update_mask_0/reg_out[10][15] , \update_mask_0/reg_out[10][14] ,
         \update_mask_0/reg_out[10][13] , \update_mask_0/reg_out[10][12] ,
         \update_mask_0/reg_out[10][11] , \update_mask_0/reg_out[10][10] ,
         \update_mask_0/reg_out[10][9] , \update_mask_0/reg_out[10][8] ,
         \update_mask_0/reg_out[10][7] , \update_mask_0/reg_out[10][6] ,
         \update_mask_0/reg_out[10][5] , \update_mask_0/reg_out[10][4] ,
         \update_mask_0/reg_out[10][3] , \update_mask_0/reg_out[10][2] ,
         \update_mask_0/reg_out[10][1] , \update_mask_0/reg_out[10][0] ,
         \update_mask_0/reg_out[9][19] , \update_mask_0/reg_out[9][18] ,
         \update_mask_0/reg_out[9][17] , \update_mask_0/reg_out[9][16] ,
         \update_mask_0/reg_out[9][15] , \update_mask_0/reg_out[9][14] ,
         \update_mask_0/reg_out[9][13] , \update_mask_0/reg_out[9][12] ,
         \update_mask_0/reg_out[9][11] , \update_mask_0/reg_out[9][10] ,
         \update_mask_0/reg_out[9][9] , \update_mask_0/reg_out[9][8] ,
         \update_mask_0/reg_out[9][7] , \update_mask_0/reg_out[9][6] ,
         \update_mask_0/reg_out[9][5] , \update_mask_0/reg_out[9][4] ,
         \update_mask_0/reg_out[9][3] , \update_mask_0/reg_out[9][2] ,
         \update_mask_0/reg_out[9][1] , \update_mask_0/reg_out[9][0] ,
         \update_mask_0/reg_out[8][19] , \update_mask_0/reg_out[8][18] ,
         \update_mask_0/reg_out[8][17] , \update_mask_0/reg_out[8][16] ,
         \update_mask_0/reg_out[8][15] , \update_mask_0/reg_out[8][14] ,
         \update_mask_0/reg_out[8][13] , \update_mask_0/reg_out[8][12] ,
         \update_mask_0/reg_out[8][11] , \update_mask_0/reg_out[8][10] ,
         \update_mask_0/reg_out[8][9] , \update_mask_0/reg_out[8][8] ,
         \update_mask_0/reg_out[8][7] , \update_mask_0/reg_out[8][6] ,
         \update_mask_0/reg_out[8][5] , \update_mask_0/reg_out[8][4] ,
         \update_mask_0/reg_out[8][3] , \update_mask_0/reg_out[8][2] ,
         \update_mask_0/reg_out[8][1] , \update_mask_0/reg_out[8][0] ,
         \update_mask_0/reg_out[7][19] , \update_mask_0/reg_out[7][18] ,
         \update_mask_0/reg_out[7][17] , \update_mask_0/reg_out[7][16] ,
         \update_mask_0/reg_out[7][15] , \update_mask_0/reg_out[7][14] ,
         \update_mask_0/reg_out[7][13] , \update_mask_0/reg_out[7][12] ,
         \update_mask_0/reg_out[7][11] , \update_mask_0/reg_out[7][10] ,
         \update_mask_0/reg_out[7][9] , \update_mask_0/reg_out[7][8] ,
         \update_mask_0/reg_out[7][7] , \update_mask_0/reg_out[7][6] ,
         \update_mask_0/reg_out[7][5] , \update_mask_0/reg_out[7][4] ,
         \update_mask_0/reg_out[7][3] , \update_mask_0/reg_out[7][2] ,
         \update_mask_0/reg_out[7][1] , \update_mask_0/reg_out[7][0] ,
         \update_mask_0/reg_out[6][19] , \update_mask_0/reg_out[6][18] ,
         \update_mask_0/reg_out[6][17] , \update_mask_0/reg_out[6][16] ,
         \update_mask_0/reg_out[6][15] , \update_mask_0/reg_out[6][14] ,
         \update_mask_0/reg_out[6][13] , \update_mask_0/reg_out[6][12] ,
         \update_mask_0/reg_out[6][11] , \update_mask_0/reg_out[6][10] ,
         \update_mask_0/reg_out[6][9] , \update_mask_0/reg_out[6][8] ,
         \update_mask_0/reg_out[6][7] , \update_mask_0/reg_out[6][6] ,
         \update_mask_0/reg_out[6][5] , \update_mask_0/reg_out[6][4] ,
         \update_mask_0/reg_out[6][3] , \update_mask_0/reg_out[6][2] ,
         \update_mask_0/reg_out[6][1] , \update_mask_0/reg_out[6][0] ,
         \update_mask_0/reg_out[5][19] , \update_mask_0/reg_out[5][18] ,
         \update_mask_0/reg_out[5][17] , \update_mask_0/reg_out[5][16] ,
         \update_mask_0/reg_out[5][15] , \update_mask_0/reg_out[5][14] ,
         \update_mask_0/reg_out[5][13] , \update_mask_0/reg_out[5][12] ,
         \update_mask_0/reg_out[5][11] , \update_mask_0/reg_out[5][10] ,
         \update_mask_0/reg_out[5][9] , \update_mask_0/reg_out[5][8] ,
         \update_mask_0/reg_out[5][7] , \update_mask_0/reg_out[5][6] ,
         \update_mask_0/reg_out[5][5] , \update_mask_0/reg_out[5][4] ,
         \update_mask_0/reg_out[5][3] , \update_mask_0/reg_out[5][2] ,
         \update_mask_0/reg_out[5][1] , \update_mask_0/reg_out[5][0] ,
         \update_mask_0/reg_out[4][19] , \update_mask_0/reg_out[4][18] ,
         \update_mask_0/reg_out[4][17] , \update_mask_0/reg_out[4][16] ,
         \update_mask_0/reg_out[4][15] , \update_mask_0/reg_out[4][14] ,
         \update_mask_0/reg_out[4][13] , \update_mask_0/reg_out[4][12] ,
         \update_mask_0/reg_out[4][11] , \update_mask_0/reg_out[4][10] ,
         \update_mask_0/reg_out[4][9] , \update_mask_0/reg_out[4][8] ,
         \update_mask_0/reg_out[4][7] , \update_mask_0/reg_out[4][6] ,
         \update_mask_0/reg_out[4][5] , \update_mask_0/reg_out[4][4] ,
         \update_mask_0/reg_out[4][3] , \update_mask_0/reg_out[4][2] ,
         \update_mask_0/reg_out[4][1] , \update_mask_0/reg_out[4][0] ,
         \update_mask_0/reg_out[3][19] , \update_mask_0/reg_out[3][18] ,
         \update_mask_0/reg_out[3][17] , \update_mask_0/reg_out[3][16] ,
         \update_mask_0/reg_out[3][15] , \update_mask_0/reg_out[3][14] ,
         \update_mask_0/reg_out[3][13] , \update_mask_0/reg_out[3][12] ,
         \update_mask_0/reg_out[3][11] , \update_mask_0/reg_out[3][10] ,
         \update_mask_0/reg_out[3][9] , \update_mask_0/reg_out[3][8] ,
         \update_mask_0/reg_out[3][7] , \update_mask_0/reg_out[3][6] ,
         \update_mask_0/reg_out[3][5] , \update_mask_0/reg_out[3][4] ,
         \update_mask_0/reg_out[3][3] , \update_mask_0/reg_out[3][2] ,
         \update_mask_0/reg_out[3][1] , \update_mask_0/reg_out[3][0] ,
         \update_mask_0/reg_out[2][19] , \update_mask_0/reg_out[2][18] ,
         \update_mask_0/reg_out[2][17] , \update_mask_0/reg_out[2][16] ,
         \update_mask_0/reg_out[2][15] , \update_mask_0/reg_out[2][14] ,
         \update_mask_0/reg_out[2][13] , \update_mask_0/reg_out[2][12] ,
         \update_mask_0/reg_out[2][11] , \update_mask_0/reg_out[2][10] ,
         \update_mask_0/reg_out[2][9] , \update_mask_0/reg_out[2][8] ,
         \update_mask_0/reg_out[2][7] , \update_mask_0/reg_out[2][6] ,
         \update_mask_0/reg_out[2][5] , \update_mask_0/reg_out[2][4] ,
         \update_mask_0/reg_out[2][3] , \update_mask_0/reg_out[2][2] ,
         \update_mask_0/reg_out[2][1] , \update_mask_0/reg_out[2][0] ,
         \update_mask_0/reg_out[1][19] , \update_mask_0/reg_out[1][18] ,
         \update_mask_0/reg_out[1][17] , \update_mask_0/reg_out[1][16] ,
         \update_mask_0/reg_out[1][15] , \update_mask_0/reg_out[1][14] ,
         \update_mask_0/reg_out[1][13] , \update_mask_0/reg_out[1][12] ,
         \update_mask_0/reg_out[1][11] , \update_mask_0/reg_out[1][10] ,
         \update_mask_0/reg_out[1][9] , \update_mask_0/reg_out[1][8] ,
         \update_mask_0/reg_out[1][7] , \update_mask_0/reg_out[1][6] ,
         \update_mask_0/reg_out[1][5] , \update_mask_0/reg_out[1][4] ,
         \update_mask_0/reg_out[1][3] , \update_mask_0/reg_out[1][2] ,
         \update_mask_0/reg_out[1][1] , \update_mask_0/reg_out[1][0] ,
         \update_mask_0/reg_out[0][19] , \update_mask_0/reg_out[0][18] ,
         \update_mask_0/reg_out[0][17] , \update_mask_0/reg_out[0][16] ,
         \update_mask_0/reg_out[0][15] , \update_mask_0/reg_out[0][14] ,
         \update_mask_0/reg_out[0][13] , \update_mask_0/reg_out[0][12] ,
         \update_mask_0/reg_out[0][11] , \update_mask_0/reg_out[0][10] ,
         \update_mask_0/reg_out[0][9] , \update_mask_0/reg_out[0][8] ,
         \update_mask_0/reg_out[0][7] , \update_mask_0/reg_out[0][6] ,
         \update_mask_0/reg_out[0][5] , \update_mask_0/reg_out[0][4] ,
         \update_mask_0/reg_out[0][3] , \update_mask_0/reg_out[0][2] ,
         \update_mask_0/reg_out[0][1] , \update_mask_0/reg_out[0][0] ,
         \update_mask_0/n4206 , \update_mask_0/n4205 , \update_mask_0/N31 ,
         \update_mask_0/N30 , \update_mask_0/N29 , \update_mask_0/N28 ,
         \update_mask_0/N27 , \update_mask_0/N26 , \update_mask_0/N25 ,
         \update_mask_0/N24 , \update_mask_0/N23 , \update_output_0/n6703 ,
         \update_output_0/n6702 , \update_output_0/n6701 ,
         \update_output_0/n6700 , \update_output_0/n6699 ,
         \update_output_0/n6698 , \update_output_0/n6697 ,
         \update_output_0/n6696 , \update_output_0/n6695 ,
         \update_output_0/n6694 , \update_output_0/n6693 ,
         \update_output_0/n6692 , \update_output_0/n6691 ,
         \update_output_0/n6690 , \update_output_0/n6689 ,
         \update_output_0/n6688 , \update_output_0/n6687 ,
         \update_output_0/n6686 , \update_output_0/n6685 ,
         \update_output_0/n6684 , \update_output_0/n6683 ,
         \update_output_0/n6682 , \update_output_0/n6681 ,
         \update_output_0/n6680 , \update_output_0/n6679 ,
         \update_output_0/n6678 , \update_output_0/n6677 ,
         \update_output_0/n6676 , \update_output_0/n6675 ,
         \update_output_0/n6674 , \update_output_0/n6673 ,
         \update_output_0/n6672 , \update_output_0/n6671 ,
         \update_output_0/n6670 , \update_output_0/n6669 ,
         \update_output_0/n6668 , \update_output_0/n6667 ,
         \update_output_0/n6666 , \update_output_0/n6665 ,
         \update_output_0/n6664 , \update_output_0/n6583 ,
         \update_output_0/n6582 , \update_output_0/n6581 ,
         \update_output_0/n6580 , \update_output_0/n6579 ,
         \update_output_0/n6578 , \update_output_0/n6577 ,
         \update_output_0/n6576 , \update_output_0/n6575 ,
         \update_output_0/n6574 , \update_output_0/n6573 ,
         \update_output_0/n6572 , \update_output_0/n6571 ,
         \update_output_0/n6570 , \update_output_0/n6569 ,
         \update_output_0/n6568 , \update_output_0/n6567 ,
         \update_output_0/n6566 , \update_output_0/n6565 ,
         \update_output_0/n6564 , \update_output_0/n6563 ,
         \update_output_0/n6562 , \update_output_0/n6561 ,
         \update_output_0/n6560 , \update_output_0/n6559 ,
         \update_output_0/n6558 , \update_output_0/n6557 ,
         \update_output_0/n6556 , \update_output_0/n6555 ,
         \update_output_0/n6554 , \update_output_0/n6553 ,
         \update_output_0/n6552 , \update_output_0/n6551 ,
         \update_output_0/n6550 , \update_output_0/n6549 ,
         \update_output_0/n6548 , \update_output_0/n6547 ,
         \update_output_0/n6546 , \update_output_0/n6545 ,
         \update_output_0/n6544 , \update_output_0/n6443 ,
         \update_output_0/n6442 , \update_output_0/n6441 ,
         \update_output_0/n6440 , \update_output_0/n6439 ,
         \update_output_0/n6438 , \update_output_0/n6437 ,
         \update_output_0/n6436 , \update_output_0/n6435 ,
         \update_output_0/n6434 , \update_output_0/n6433 ,
         \update_output_0/n6432 , \update_output_0/n6431 ,
         \update_output_0/n6430 , \update_output_0/n6429 ,
         \update_output_0/n6428 , \update_output_0/n6427 ,
         \update_output_0/n6426 , \update_output_0/n6425 ,
         \update_output_0/n6424 , \update_output_0/n3549 ,
         \update_output_0/n1535 , \update_output_0/n9020 ,
         \update_output_0/n9019 , \update_output_0/N34 , \update_output_0/N33 ,
         \update_output_0/N32 , \update_output_0/N31 , \update_output_0/N30 ,
         \update_output_0/N29 , \update_output_0/N28 , \update_output_0/N27 ,
         n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099,
         n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109,
         n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119,
         n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129,
         n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139,
         n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149,
         n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159,
         n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169,
         n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179,
         n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189,
         n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199,
         n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209,
         n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219,
         n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229,
         n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239,
         n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249,
         n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259,
         n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269,
         n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279,
         n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289,
         n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299,
         n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309,
         n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319,
         n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329,
         n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339,
         n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349,
         n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359,
         n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369,
         n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379,
         n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389,
         n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399,
         n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409,
         n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419,
         n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429,
         n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439,
         n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449,
         n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459,
         n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469,
         n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479,
         n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489,
         n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499,
         n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509,
         n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519,
         n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529,
         n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539,
         n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549,
         n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559,
         n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569,
         n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579,
         n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589,
         n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599,
         n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609,
         n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619,
         n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629,
         n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639,
         n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649,
         n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659,
         n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669,
         n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679,
         n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689,
         n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699,
         n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709,
         n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719,
         n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729,
         n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739,
         n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749,
         n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759,
         n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769,
         n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779,
         n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789,
         n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799,
         n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809,
         n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819,
         n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829,
         n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839,
         n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849,
         n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859,
         n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869,
         n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879,
         n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889,
         n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899,
         n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909,
         n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919,
         n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929,
         n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939,
         n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949,
         n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959,
         n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969,
         n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979,
         n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989,
         n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999,
         n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009,
         n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019,
         n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029,
         n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039,
         n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049,
         n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059,
         n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069,
         n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079,
         n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089,
         n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099,
         n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109,
         n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119,
         n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129,
         n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139,
         n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149,
         n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159,
         n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169,
         n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179,
         n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189,
         n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199,
         n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209,
         n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219,
         n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229,
         n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239,
         n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249,
         n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259,
         n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269,
         n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279,
         n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289,
         n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299,
         n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309,
         n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319,
         n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329,
         n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339,
         n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349,
         n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359,
         n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369,
         n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379,
         n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389,
         n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399,
         n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409,
         n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419,
         n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429,
         n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439,
         n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449,
         n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459,
         n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469,
         n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479,
         n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489,
         n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499,
         n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509,
         n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519,
         n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529,
         n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539,
         n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549,
         n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559,
         n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569,
         n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579,
         n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589,
         n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599,
         n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609,
         n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619,
         n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629,
         n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639,
         n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649,
         n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659,
         n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669,
         n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679,
         n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689,
         n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699,
         n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709,
         n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719,
         n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729,
         n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739,
         n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749,
         n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759,
         n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769,
         n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779,
         n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789,
         n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799,
         n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809,
         n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819,
         n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829,
         n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839,
         n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849,
         n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859,
         n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869,
         n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879,
         n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889,
         n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899,
         n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909,
         n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919,
         n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929,
         n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939,
         n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949,
         n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959,
         n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969,
         n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979,
         n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989,
         n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999,
         n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009,
         n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019,
         n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029,
         n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039,
         n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049,
         n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059,
         n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069,
         n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079,
         n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089,
         n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099,
         n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109,
         n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119,
         n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129,
         n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139,
         n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149,
         n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159,
         n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169,
         n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179,
         n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189,
         n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199,
         n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209,
         n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219,
         n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229,
         n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239,
         n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249,
         n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259,
         n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269,
         n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279,
         n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289,
         n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299,
         n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309,
         n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319,
         n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329,
         n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339,
         n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349,
         n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359,
         n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369,
         n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379,
         n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389,
         n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399,
         n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409,
         n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419,
         n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429,
         n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439,
         n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449,
         n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459,
         n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469,
         n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479,
         n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489,
         n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499,
         n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509,
         n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519,
         n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529,
         n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539,
         n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549,
         n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559,
         n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569,
         n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579,
         n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589,
         n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599,
         n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609,
         n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619,
         n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629,
         n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639,
         n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649,
         n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659,
         n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669,
         n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679,
         n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689,
         n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699,
         n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709,
         n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719,
         n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729,
         n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739,
         n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749,
         n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759,
         n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769,
         n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779,
         n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789,
         n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799,
         n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809,
         n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819,
         n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829,
         n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839,
         n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849,
         n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859,
         n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869,
         n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879,
         n5880, n5881, n5882, n5883, n5884, n5885, \update_output_0/n3460 ,
         \update_output_0/n3459 , \update_output_0/n3456 ,
         \update_output_0/n3455 , \update_output_0/n3452 ,
         \update_output_0/n3451 , \update_output_0/n3448 ,
         \update_output_0/n3447 , \update_output_0/n3444 ,
         \update_output_0/n3443 , \update_output_0/n3440 ,
         \update_output_0/n3439 , \update_output_0/n3436 ,
         \update_output_0/n3435 , \update_output_0/n3432 ,
         \update_output_0/n3431 , \update_output_0/n3428 ,
         \update_output_0/n3427 , \update_output_0/n3424 ,
         \update_output_0/n3423 , \update_output_0/n3420 ,
         \update_output_0/n3419 , \update_output_0/n3416 ,
         \update_output_0/n3415 , \update_output_0/n3412 ,
         \update_output_0/n3411 , \update_output_0/n3408 ,
         \update_output_0/n3407 , \update_output_0/n3404 ,
         \update_output_0/n3403 , \update_output_0/n3400 ,
         \update_output_0/n3399 , \update_output_0/n3396 ,
         \update_output_0/n3395 , \update_output_0/n3392 ,
         \update_output_0/n3391 , \update_output_0/n3388 ,
         \update_output_0/n3387 , \update_output_0/n3384 ,
         \update_output_0/n3383 , \update_output_0/n3380 ,
         \update_output_0/n3379 , \update_output_0/n3376 ,
         \update_output_0/n3375 , \update_output_0/n3372 ,
         \update_output_0/n3371 , \update_output_0/n3368 ,
         \update_output_0/n3367 , \update_output_0/n3364 ,
         \update_output_0/n3363 , \update_output_0/n3360 ,
         \update_output_0/n3359 , \update_output_0/n3356 ,
         \update_output_0/n3355 , \update_output_0/n3352 ,
         \update_output_0/n3351 , \update_output_0/n3348 ,
         \update_output_0/n3347 , \update_output_0/n3344 ,
         \update_output_0/n3343 , \update_output_0/n3340 ,
         \update_output_0/n3339 , \update_output_0/n3336 ,
         \update_output_0/n3335 , \update_output_0/n3332 ,
         \update_output_0/n3331 , \update_output_0/n3328 ,
         \update_output_0/n3327 , \update_output_0/n3324 ,
         \update_output_0/n3323 , \update_output_0/n3320 ,
         \update_output_0/n3319 , \update_output_0/n3316 ,
         \update_output_0/n3315 , \update_output_0/n3312 ,
         \update_output_0/n3311 , \update_output_0/n3308 ,
         \update_output_0/n3307 , \update_output_0/n3304 ,
         \update_output_0/n3303 , \update_output_0/n3300 ,
         \update_output_0/n3299 , \update_output_0/n3296 ,
         \update_output_0/n3295 , \update_output_0/n3292 ,
         \update_output_0/n3291 , \update_output_0/n3288 ,
         \update_output_0/n3287 , \update_output_0/n3284 ,
         \update_output_0/n3283 , \update_output_0/n3280 ,
         \update_output_0/n3279 , \update_output_0/n3276 ,
         \update_output_0/n3275 , \update_output_0/n3272 ,
         \update_output_0/n3271 , \update_output_0/n3268 ,
         \update_output_0/n3267 , \update_output_0/n3264 ,
         \update_output_0/n3263 , \update_output_0/n3260 ,
         \update_output_0/n3259 , \update_output_0/n3256 ,
         \update_output_0/n3255 , \update_output_0/n3252 ,
         \update_output_0/n3251 , \update_output_0/n3248 ,
         \update_output_0/n3247 , \update_output_0/n3244 ,
         \update_output_0/n3243 , \update_output_0/n3240 ,
         \update_output_0/n3239 , \update_output_0/n3236 ,
         \update_output_0/n3235 , \update_output_0/n3232 ,
         \update_output_0/n3231 , \update_output_0/n3228 ,
         \update_output_0/n3227 , \update_output_0/n3224 ,
         \update_output_0/n3223 , \update_output_0/n3220 ,
         \update_output_0/n3219 , \update_output_0/n3216 ,
         \update_output_0/n3215 , \update_output_0/n3212 ,
         \update_output_0/n3211 , \update_output_0/n3208 ,
         \update_output_0/n3207 , \update_output_0/n3204 ,
         \update_output_0/n3203 , \update_output_0/n3200 ,
         \update_output_0/n3199 , \update_output_0/n3196 ,
         \update_output_0/n3195 , \update_output_0/n3192 ,
         \update_output_0/n3191 , \update_output_0/n3188 ,
         \update_output_0/n3187 , \update_output_0/n3184 ,
         \update_output_0/n3183 , \update_output_0/n3180 ,
         \update_output_0/n3179 , \update_output_0/n3176 ,
         \update_output_0/n3175 , \update_output_0/n3172 ,
         \update_output_0/n3171 , \update_output_0/n3168 ,
         \update_output_0/n3167 , \update_output_0/n3164 ,
         \update_output_0/n3163 , \update_output_0/n3160 ,
         \update_output_0/n3159 , \update_output_0/n3156 ,
         \update_output_0/n3155 , \update_output_0/n3152 ,
         \update_output_0/n3151 , \update_output_0/n3148 ,
         \update_output_0/n3147 , \update_output_0/n3144 ,
         \update_output_0/n3143 , \update_output_0/n3140 ,
         \update_output_0/n3139 , \update_output_0/n3136 ,
         \update_output_0/n3135 , \update_output_0/n3132 ,
         \update_output_0/n3131 , \update_output_0/n3128 ,
         \update_output_0/n3127 , \update_output_0/n3124 ,
         \update_output_0/n3123 , \update_output_0/n3120 ,
         \update_output_0/n3119 , \update_output_0/n3116 ,
         \update_output_0/n3115 , \update_output_0/n3112 ,
         \update_output_0/n3111 , \update_output_0/n3108 ,
         \update_output_0/n3107 , \update_output_0/n3104 ,
         \update_output_0/n3103 , \update_output_0/n3100 ,
         \update_output_0/n3099 , \update_output_0/n3096 ,
         \update_output_0/n3095 , \update_output_0/n3092 ,
         \update_output_0/n3091 , \update_output_0/n3088 ,
         \update_output_0/n3087 , \update_output_0/n3084 ,
         \update_output_0/n3083 , \update_output_0/n3080 ,
         \update_output_0/n3079 , \update_output_0/n3076 ,
         \update_output_0/n3075 , \update_output_0/n3072 ,
         \update_output_0/n3071 , \update_output_0/n3068 ,
         \update_output_0/n3067 , \update_output_0/n3064 ,
         \update_output_0/n3063 , \update_output_0/n3060 ,
         \update_output_0/n3059 , \update_output_0/n3056 ,
         \update_output_0/n3055 , \update_output_0/n3052 ,
         \update_output_0/n3051 , \update_output_0/n3048 ,
         \update_output_0/n3047 , \update_output_0/n3044 ,
         \update_output_0/n3043 , \update_output_0/n3040 ,
         \update_output_0/n3039 , \update_output_0/n3036 ,
         \update_output_0/n3035 , \update_output_0/n3032 ,
         \update_output_0/n3031 , \update_output_0/n3028 ,
         \update_output_0/n3027 , \update_output_0/n3024 ,
         \update_output_0/n3023 , \update_output_0/n3020 ,
         \update_output_0/n3019 , \update_output_0/n3016 ,
         \update_output_0/n3015 , \update_output_0/n3012 ,
         \update_output_0/n3011 , \update_output_0/n3008 ,
         \update_output_0/n3007 , \update_output_0/n3004 ,
         \update_output_0/n3003 , \update_output_0/n3000 ,
         \update_output_0/n2999 , \update_output_0/n2996 ,
         \update_output_0/n2995 , \update_output_0/n2992 ,
         \update_output_0/n2991 , \update_output_0/n2988 ,
         \update_output_0/n2987 , \update_output_0/n2984 ,
         \update_output_0/n2983 , \update_output_0/n2980 ,
         \update_output_0/n2979 , \update_output_0/n2976 ,
         \update_output_0/n2975 , \update_output_0/n2972 ,
         \update_output_0/n2971 , \update_output_0/n2968 ,
         \update_output_0/n2967 , \update_output_0/n2964 ,
         \update_output_0/n2963 , \update_output_0/n2960 ,
         \update_output_0/n2959 , \update_output_0/n2956 ,
         \update_output_0/n2955 , \update_output_0/n2952 ,
         \update_output_0/n2951 , \update_output_0/n2948 ,
         \update_output_0/n2947 , \update_output_0/n2944 ,
         \update_output_0/n2943 , \update_output_0/n2940 ,
         \update_output_0/n2939 , \update_output_0/n2936 ,
         \update_output_0/n2935 , \update_output_0/n2932 ,
         \update_output_0/n2931 , \update_output_0/n2928 ,
         \update_output_0/n2927 , \update_output_0/n2924 ,
         \update_output_0/n2923 , \update_output_0/n2920 ,
         \update_output_0/n2919 , \update_output_0/n2916 ,
         \update_output_0/n2915 , \update_output_0/n2912 ,
         \update_output_0/n2911 , \update_output_0/n2908 ,
         \update_output_0/n2907 , \update_output_0/n2904 ,
         \update_output_0/n2903 , \update_output_0/n2900 ,
         \update_output_0/n2899 , \update_output_0/n2896 ,
         \update_output_0/n2895 , \update_output_0/n2892 ,
         \update_output_0/n2891 , \update_output_0/n2888 ,
         \update_output_0/n2887 , \update_output_0/n2884 ,
         \update_output_0/n2883 , \update_output_0/n2880 ,
         \update_output_0/n2879 , \update_output_0/n2876 ,
         \update_output_0/n2875 , \update_output_0/n2872 ,
         \update_output_0/n2871 , \update_output_0/n2868 ,
         \update_output_0/n2867 , \update_output_0/n2864 ,
         \update_output_0/n2863 , \update_output_0/n2860 ,
         \update_output_0/n2859 , \update_output_0/n2856 ,
         \update_output_0/n2855 , \update_output_0/n2852 ,
         \update_output_0/n2851 , \update_output_0/n2848 ,
         \update_output_0/n2847 , \update_output_0/n2844 ,
         \update_output_0/n2843 , \update_output_0/n2840 ,
         \update_output_0/n2839 , \update_output_0/n2836 ,
         \update_output_0/n2835 , \update_output_0/n2832 ,
         \update_output_0/n2831 , \update_output_0/n2828 ,
         \update_output_0/n2827 , \update_output_0/n2824 ,
         \update_output_0/n2823 , \update_output_0/n2820 ,
         \update_output_0/n2819 , \update_output_0/n2816 ,
         \update_output_0/n2815 , \update_output_0/n2812 ,
         \update_output_0/n2811 , \update_output_0/n2808 ,
         \update_output_0/n2807 , \update_output_0/n2804 ,
         \update_output_0/n2803 , \update_output_0/n2800 ,
         \update_output_0/n2799 , \update_output_0/n2796 ,
         \update_output_0/n2795 , \update_output_0/n2792 ,
         \update_output_0/n2791 , \update_output_0/n2788 ,
         \update_output_0/n2787 , \update_output_0/n2784 ,
         \update_output_0/n2783 , \update_output_0/n2780 ,
         \update_output_0/n2779 , \update_output_0/n2776 ,
         \update_output_0/n2775 , \update_output_0/n2772 ,
         \update_output_0/n2771 , \update_output_0/n2768 ,
         \update_output_0/n2767 , \update_output_0/n2764 ,
         \update_output_0/n2763 , \update_output_0/n2760 ,
         \update_output_0/n2759 , \update_output_0/n2756 ,
         \update_output_0/n2755 , \update_output_0/n2752 ,
         \update_output_0/n2751 , \update_output_0/n2748 ,
         \update_output_0/n2747 , \update_output_0/n2744 ,
         \update_output_0/n2743 , \update_output_0/n2740 ,
         \update_output_0/n2739 , \update_output_0/n2736 ,
         \update_output_0/n2735 , \update_output_0/n2732 ,
         \update_output_0/n2731 , \update_output_0/n2728 ,
         \update_output_0/n2727 , \update_output_0/n2724 ,
         \update_output_0/n2723 , \update_output_0/n2720 ,
         \update_output_0/n2719 , \update_output_0/n2716 ,
         \update_output_0/n2715 , \update_output_0/n2712 ,
         \update_output_0/n2711 , \update_output_0/n2708 ,
         \update_output_0/n2707 , \update_output_0/n2704 ,
         \update_output_0/n2703 , \update_output_0/n2700 ,
         \update_output_0/n2699 , \update_output_0/n2696 ,
         \update_output_0/n2695 , \update_output_0/n2692 ,
         \update_output_0/n2691 , \update_output_0/n2688 ,
         \update_output_0/n2687 , \update_output_0/n2684 ,
         \update_output_0/n2683 , \update_output_0/n2680 ,
         \update_output_0/n2679 , \update_output_0/n2676 ,
         \update_output_0/n2675 , \update_output_0/n2672 ,
         \update_output_0/n2671 , \update_output_0/n2668 ,
         \update_output_0/n2667 , \update_output_0/n2664 ,
         \update_output_0/n2663 , \update_output_0/n2660 ,
         \update_output_0/n2659 , \update_output_0/n2656 ,
         \update_output_0/n2655 , \update_output_0/n2652 ,
         \update_output_0/n2651 , \update_output_0/n2648 ,
         \update_output_0/n2647 , \update_output_0/n2644 ,
         \update_output_0/n2643 , \update_output_0/n2640 ,
         \update_output_0/n2639 , \update_output_0/n2636 ,
         \update_output_0/n2635 , \update_output_0/n2632 ,
         \update_output_0/n2631 , \update_output_0/n2628 ,
         \update_output_0/n2627 , \update_output_0/n2624 ,
         \update_output_0/n2623 , \update_output_0/n2620 ,
         \update_output_0/n2619 , \update_output_0/n2616 ,
         \update_output_0/n2615 , \update_output_0/n2612 ,
         \update_output_0/n2611 , \update_output_0/n2608 ,
         \update_output_0/n2607 , \update_output_0/n2604 ,
         \update_output_0/n2603 , \update_output_0/n2600 ,
         \update_output_0/n2599 , \update_output_0/n2596 ,
         \update_output_0/n2595 , \update_output_0/n2592 ,
         \update_output_0/n2591 , \update_output_0/n2588 ,
         \update_output_0/n2587 , \update_output_0/n2584 ,
         \update_output_0/n2583 , \update_output_0/n2580 ,
         \update_output_0/n2579 , \update_output_0/n2576 ,
         \update_output_0/n2575 , \update_output_0/n2572 ,
         \update_output_0/n2571 , \update_output_0/n2568 ,
         \update_output_0/n2567 , \update_output_0/n2564 ,
         \update_output_0/n2563 , \update_output_0/n2560 ,
         \update_output_0/n2559 , \update_output_0/n2556 ,
         \update_output_0/n2555 , \update_output_0/n2552 ,
         \update_output_0/n2551 , \update_output_0/n2548 ,
         \update_output_0/n2547 , \update_output_0/n2544 ,
         \update_output_0/n2543 , \update_output_0/n2540 ,
         \update_output_0/n2539 , \update_output_0/n2536 ,
         \update_output_0/n2535 , \update_output_0/n2532 ,
         \update_output_0/n2531 , \update_output_0/n2528 ,
         \update_output_0/n2527 , \update_output_0/n2524 ,
         \update_output_0/n2523 , \update_output_0/n2520 ,
         \update_output_0/n2519 , \update_output_0/n2516 ,
         \update_output_0/n2515 , \update_output_0/n2512 ,
         \update_output_0/n2511 , \update_output_0/n2508 ,
         \update_output_0/n2507 , \update_output_0/n2504 ,
         \update_output_0/n2503 , \update_output_0/n2500 ,
         \update_output_0/n2499 , \update_output_0/n2496 ,
         \update_output_0/n2495 , \update_output_0/n2492 ,
         \update_output_0/n2491 , \update_output_0/n2488 ,
         \update_output_0/n2487 , \update_output_0/n2484 ,
         \update_output_0/n2483 , \update_output_0/n2480 ,
         \update_output_0/n2479 , \update_output_0/n2476 ,
         \update_output_0/n2475 , \update_output_0/n2472 ,
         \update_output_0/n2471 , \update_output_0/n2468 ,
         \update_output_0/n2467 , \update_output_0/n2464 ,
         \update_output_0/n2463 , \update_output_0/n2460 ,
         \update_output_0/n2459 , \update_output_0/n2456 ,
         \update_output_0/n2455 , \update_output_0/n2452 ,
         \update_output_0/n2451 , \update_output_0/n2448 ,
         \update_output_0/n2447 , \update_output_0/n2444 ,
         \update_output_0/n2443 , \update_output_0/n2440 ,
         \update_output_0/n2439 , \update_output_0/n2436 ,
         \update_output_0/n2435 , \update_output_0/n2432 ,
         \update_output_0/n2431 , \update_output_0/n2428 ,
         \update_output_0/n2427 , \update_output_0/n2424 ,
         \update_output_0/n2423 , \update_output_0/n2420 ,
         \update_output_0/n2419 , \update_output_0/n2416 ,
         \update_output_0/n2415 , \update_output_0/n2412 ,
         \update_output_0/n2411 , \update_output_0/n2408 ,
         \update_output_0/n2407 , \update_output_0/n2404 ,
         \update_output_0/n2403 , \update_output_0/n2400 ,
         \update_output_0/n2399 , \update_output_0/n2396 ,
         \update_output_0/n2395 , \update_output_0/n2392 ,
         \update_output_0/n2391 , \update_output_0/n2388 ,
         \update_output_0/n2387 , \update_output_0/n2384 ,
         \update_output_0/n2383 , \update_output_0/n2380 ,
         \update_output_0/n2379 , \update_output_0/n2376 ,
         \update_output_0/n2375 , \update_output_0/n2372 ,
         \update_output_0/n2371 , \update_output_0/n2368 ,
         \update_output_0/n2367 , \update_output_0/n2364 ,
         \update_output_0/n2363 , \update_output_0/n2360 ,
         \update_output_0/n2359 , \update_output_0/n2356 ,
         \update_output_0/n2355 , \update_output_0/n2352 ,
         \update_output_0/n2351 , \update_output_0/n2348 ,
         \update_output_0/n2347 , \update_output_0/n2344 ,
         \update_output_0/n2343 , \update_output_0/n2340 ,
         \update_output_0/n2339 , \update_output_0/n2336 ,
         \update_output_0/n2335 , \update_output_0/n2332 ,
         \update_output_0/n2331 , \update_output_0/n2328 ,
         \update_output_0/n2327 , \update_output_0/n2324 ,
         \update_output_0/n2323 , \update_output_0/n2320 ,
         \update_output_0/n2319 , \update_output_0/n2316 ,
         \update_output_0/n2315 , \update_output_0/n2312 ,
         \update_output_0/n2311 , \update_output_0/n2308 ,
         \update_output_0/n2307 , \update_output_0/n2304 ,
         \update_output_0/n2303 , \update_output_0/n2300 ,
         \update_output_0/n2299 , \update_output_0/n2296 ,
         \update_output_0/n2295 , \update_output_0/n2292 ,
         \update_output_0/n2291 , \update_output_0/n2288 ,
         \update_output_0/n2287 , \update_output_0/n2284 ,
         \update_output_0/n2283 , \update_output_0/n2280 ,
         \update_output_0/n2279 , \update_output_0/n2276 ,
         \update_output_0/n2275 , \update_output_0/n2272 ,
         \update_output_0/n2271 , \update_output_0/n2268 ,
         \update_output_0/n2267 , \update_output_0/n2264 ,
         \update_output_0/n2263 , \update_output_0/n2260 ,
         \update_output_0/n2259 , \update_output_0/n2256 ,
         \update_output_0/n2255 , \update_output_0/n2252 ,
         \update_output_0/n2251 , \update_output_0/n2248 ,
         \update_output_0/n2247 , \update_output_0/n2244 ,
         \update_output_0/n2243 , \update_output_0/n2240 ,
         \update_output_0/n2239 , \update_output_0/n2236 ,
         \update_output_0/n2235 , \update_output_0/n2232 ,
         \update_output_0/n2231 , \update_output_0/n2228 ,
         \update_output_0/n2227 , \update_output_0/n2224 ,
         \update_output_0/n2223 , \update_output_0/n2220 ,
         \update_output_0/n2219 , \update_output_0/n2216 ,
         \update_output_0/n2215 , \update_output_0/n2212 ,
         \update_output_0/n2211 , \update_output_0/n2208 ,
         \update_output_0/n2207 , \update_output_0/n2204 ,
         \update_output_0/n2203 , \update_output_0/n2200 ,
         \update_output_0/n2199 , \update_output_0/n2196 ,
         \update_output_0/n2195 , \update_output_0/n2192 ,
         \update_output_0/n2191 , \update_output_0/n2188 ,
         \update_output_0/n2187 , \update_output_0/n2183 ,
         \update_output_0/n2180 , \update_output_0/n2179 ,
         \update_mask_0/n996 , \update_mask_0/n991 , \update_mask_0/n988 ,
         \update_mask_0/n1116 , \update_mask_0/n1112 , \update_mask_0/n1108 ,
         \update_mask_0/n1104 , \update_mask_0/n1100 , \update_mask_0/n1096 ,
         \update_mask_0/n1092 , \update_mask_0/n1088 , \update_mask_0/n1084 ,
         \update_mask_0/n1080 , \update_mask_0/n1076 , \update_mask_0/n1072 ,
         \update_mask_0/n1068 , \update_mask_0/n1064 , \update_mask_0/n1060 ,
         \update_mask_0/n1056 , \update_mask_0/n1052 , \update_mask_0/n1048 ,
         \update_mask_0/n1044 , \update_mask_0/n1040 , \update_mask_0/n1036 ,
         \update_mask_0/n1032 , \update_mask_0/n1028 , \update_mask_0/n1024 ,
         \update_mask_0/n1020 , \update_mask_0/n1016 , \update_mask_0/n1012 ,
         \update_mask_0/n1008 , \update_mask_0/n1004 , \update_mask_0/n1000 ,
         n999, n998, n997, n996, n995, n994, n993, n992, n991, n990, n989,
         n988, n987, n986, n985, n984, n983, n982, n981, n980, n979, n978,
         n977, n976, n975, n974, n973, n972, n971, n970, n969, n968, n967,
         n966, n965, n964, n963, n962, n961, n960, n959, n958, n957, n956,
         n955, n954, n953, n952, n951, n950, n949, n948, n947, n946, n945,
         n944, n943, n942, n941, n940, n939, n938, n937, n936, n935, n934,
         n933, n932, n931, n930, n929, n928, n927, n926, n925, n924, n923,
         n922, n921, n920, n919, n918, n917, n916, n915, n914, n913, n912,
         n911, n910, n909, n908, n907, n906, n905, n904, n903, n902, n901,
         n900, n899, n898, n897, n896, n895, n894, n893, n892, n891, n890,
         n889, n888, n887, n886, n885, n884, n883, n882, n881, n880, n879,
         n878, n877, n876, n875, n874, n873, n872, n871, n870, n869, n868,
         n867, n866, n865, n864, n863, n862, n861, n860, n859, n858, n857,
         n856, n855, n854, n853, n852, n851, n850, n849, n848, n847, n846,
         n845, n844, n843, n842, n841, n840, n839, n838, n837, n836, n835,
         n834, n833, n832, n831, n830, n829, n828, n827, n826, n825, n824,
         n823, n822, n821, n820, n819, n818, n817, n816, n815, n814, n813,
         n812, n811, n810, n809, n808, n807, n806, n805, n804, n803, n802,
         n801, n800, n799, n798, n797, n796, n795, n794, n793, n792, n791,
         n790, n789, n788, n787, n786, n785, n784, n783, n782, n781, n780,
         n779, n778, n777, n776, n775, n774, n773, n772, n771, n770, n769,
         n768, n767, n766, n765, n764, n763, n762, n761, n760, n759, n758,
         n757, n756, n755, n754, n753, n752, n751, n750, n749, n748, n747,
         n746, n745, n744, n743, n742, n741, n740, n2070, n2069, n2068, n2067,
         n2066, n2065, n2064, n2063, n2062, n2061, n2060, n2059, n2058, n2057,
         n2056, n2055, n2054, n2053, n2052, n2051, n2050, n2049, n2048, n2047,
         n2046, n2045, n2044, n2043, n2042, n2041, n2040, n2039, n2038, n2037,
         n2036, n2035, n2034, n2033, n2032, n2031, n2030, n2029, n2028, n2027,
         n2026, n2025, n2024, n2023, n2022, n2021, n2020, n2019, n2018, n2017,
         n2016, n2015, n2014, n2013, n2012, n2011, n2010, n2009, n2008, n2007,
         n2006, n2005, n2004, n2003, n2002, n2001, n2000, n1999, n1998, n1997,
         n1996, n1995, n1994, n1993, n1992, n1991, n1990, n1989, n1988, n1987,
         n1986, n1985, n1984, n1983, n1982, n1981, n1980, n1979, n1978, n1977,
         n1976, n1975, n1974, n1973, n1972, n1971, n1970, n1969, n1968, n1967,
         n1966, n1965, n1964, n1963, n1962, n1961, n1960, n1959, n1958, n1957,
         n1956, n1955, n1954, n1953, n1952, n1951, n1950, n1949, n1948, n1947,
         n1946, n1945, n1944, n1943, n1942, n1941, n1940, n1939, n1938, n1937,
         n1936, n1935, n1934, n1933, n1932, n1931, n1930, n1929, n1928, n1927,
         n1926, n1925, n1924, n1923, n1922, n1921, n1920, n1919, n1918, n1917,
         n1916, n1915, n1914, n1913, n1912, n1911, n1910, n1909, n1908, n1907,
         n1906, n1905, n1904, n1903, n1902, n1901, n1900, n1899, n1898, n1897,
         n1896, n1895, n1894, n1893, n1892, n1891, n1890, n1889, n1888, n1887,
         n1886, n1885, n1884, n1883, n1882, n1881, n1880, n1879, n1878, n1877,
         n1876, n1875, n1874, n1873, n1872, n1871, n1870, n1869, n1868, n1867,
         n1866, n1865, n1864, n1863, n1862, n1861, n1860, n1859, n1858, n1857,
         n1856, n1855, n1854, n1853, n1852, n1851, n1850, n1849, n1848, n1847,
         n1846, n1845, n1844, n1843, n1842, n1841, n1840, n1839, n1838, n1837,
         n1836, n1835, n1834, n1833, n1832, n1831, n1830, n1829, n1828, n1827,
         n1826, n1825, n1824, n1823, n1822, n1821, n1820, n1819, n1818, n1817,
         n1816, n1815, n1814, n1813, n1812, n1811, n1810, n1809, n1808, n1807,
         n1806, n1805, n1804, n1803, n1802, n1801, n1800, n1799, n1798, n1797,
         n1796, n1795, n1794, n1793, n1792, n1791, n1790, n1789, n1788, n1787,
         n1786, n1785, n1784, n1783, n1782, n1781, n1780, n1779, n1778, n1777,
         n1776, n1775, n1774, n1773, n1772, n1771, n1770, n1769, n1768, n1767,
         n1766, n1765, n1764, n1763, n1762, n1761, n1760, n1759, n1758, n1757,
         n1756, n1755, n1754, n1753, n1752, n1751, n1750, n1749, n1748, n1747,
         n1746, n1745, n1744, n1743, n1742, n1741, n1740, n1739, n1738, n1737,
         n1736, n1735, n1734, n1733, n1732, n1731, n1730, n1729, n1728, n1727,
         n1726, n1725, n1724, n1723, n1722, n1721, n1720, n1719, n1718, n1717,
         n1716, n1715, n1714, n1713, n1712, n1711, n1710, n1709, n1708, n1707,
         n1706, n1705, n1704, n1703, n1702, n1701, n1700, n1699, n1698, n1697,
         n1696, n1695, n1694, n1693, n1692, n1691, n1690, n1689, n1688, n1687,
         n1686, n1685, n1684, n1683, n1682, n1681, n1680, n1679, n1678, n1677,
         n1676, n1675, n1674, n1673, n1672, n1671, n1670, n1669, n1668, n1667,
         n1666, n1665, n1664, n1663, n1662, n1661, n1660, n1659, n1658, n1657,
         n1656, n1655, n1654, n1653, n1652, n1651, n1650, n1649, n1648, n1647,
         n1646, n1645, n1644, n1643, n1642, n1641, n1640, n1639, n1638, n1637,
         n1636, n1635, n1634, n1633, n1632, n1631, n1630, n1629, n1628, n1627,
         n1626, n1625, n1624, n1623, n1622, n1621, n1620, n1619, n1618, n1617,
         n1616, n1615, n1614, n1613, n1612, n1611, n1610, n1609, n1608, n1607,
         n1606, n1605, n1604, n1603, n1602, n1601, n1600, n1599, n1598, n1597,
         n1596, n1595, n1594, n1593, n1592, n1591, n1590, n1589, n1588, n1587,
         n1586, n1585, n1584, n1583, n1582, n1581, n1580, n1579, n1578, n1577,
         n1576, n1575, n1574, n1573, n1572, n1571, n1570, n1569, n1568, n1567,
         n1566, n1565, n1564, n1563, n1562, n1561, n1560, n1559, n1558, n1557,
         n1556, n1555, n1554, n1553, n1552, n1551, n1550, n1549, n1548, n1547,
         n1546, n1545, n1544, n1543, n1542, n1541, n1540, n1539, n1538, n1537,
         n1536, n1535, n1534, n1533, n1532, n1531, n1530, n1529, n1528, n1527,
         n1526, n1525, n1524, n1523, n1522, n1521, n1520, n1519, n1518, n1517,
         n1516, n1515, n1514, n1513, n1512, n1511, n1510, n1509, n1508, n1507,
         n1506, n1505, n1504, n1503, n1502, n1501, n1500, n1499, n1498, n1497,
         n1496, n1495, n1494, n1493, n1492, n1491, n1490, n1489, n1488, n1487,
         n1486, n1485, n1484, n1483, n1482, n1481, n1480, n1479, n1478, n1477,
         n1476, n1475, n1474, n1473, n1472, n1471, n1470, n1469, n1468, n1467,
         n1466, n1465, n1464, n1463, n1462, n1461, n1460, n1459, n1458, n1457,
         n1456, n1455, n1454, n1453, n1452, n1451, n1450, n1449, n1448, n1447,
         n1446, n1445, n1444, n1443, n1442, n1441, n1440, n1439, n1438, n1437,
         n1436, n1435, n1434, n1433, n1432, n1431, n1430, n1429, n1428, n1427,
         n1426, n1425, n1424, n1423, n1422, n1421, n1420, n1419, n1418, n1417,
         n1416, n1415, n1414, n1413, n1412, n1411, n1410, n1409, n1408, n1407,
         n1406, n1405, n1404, n1403, n1402, n1401, n1400, n1399, n1398, n1397,
         n1396, n1395, n1394, n1393, n1392, n1391, n1390, n1389, n1388, n1387,
         n1386, n1385, n1384, n1383, n1382, n1381, n1380, n1379, n1378, n1377,
         n1376, n1375, n1374, n1373, n1372, n1371, n1370, n1369, n1368, n1367,
         n1366, n1365, n1364, n1363, n1362, n1361, n1360, n1359, n1358, n1357,
         n1356, n1355, n1354, n1353, n1352, n1351, n1350, n1349, n1348, n1347,
         n1346, n1345, n1344, n1343, n1342, n1341, n1340, n1339, n1338, n1337,
         n1336, n1335, n1334, n1333, n1332, n1331, n1330, n1329, n1328, n1327,
         n1326, n1325, n1324, n1323, n1322, n1321, n1320, n1319, n1318, n1317,
         n1316, n1315, n1314, n1313, n1312, n1311, n1310, n1309, n1308, n1307,
         n1306, n1305, n1304, n1303, n1302, n1301, n1300, n1299, n1298, n1297,
         n1296, n1295, n1294, n1293, n1292, n1291, n1290, n1289, n1288, n1287,
         n1286, n1285, n1284, n1283, n1282, n1281, n1280, n1279, n1278, n1277,
         n1276, n1275, n1274, n1273, n1272, n1271, n1270, n1269, n1268, n1267,
         n1266, n1265, n1264, n1263, n1262, n1261, n1260, n1259, n1258, n1257,
         n1256, n1255, n1254, n1253, n1252, n1251, n1250, n1249, n1248, n1247,
         n1246, n1245, n1244, n1243, n1242, n1241, n1240, n1239, n1238, n1237,
         n1236, n1235, n1234, n1233, n1232, n1231, n1230, n1229, n1228, n1227,
         n1226, n1225, n1224, n1223, n1222, n1221, n1220, n1219, n1218, n1217,
         n1216, n1215, n1214, n1213, n1212, n1211, n1210, n1209, n1208, n1207,
         n1206, n1205, n1204, n1203, n1202, n1201, n1200, n1199, n1198, n1197,
         n1196, n1195, n1194, n1193, n1192, n1191, n1190, n1189, n1188, n1187,
         n1186, n1185, n1184, n1183, n1182, n1181, n1180, n1179, n1178, n1177,
         n1176, n1175, n1174, n1173, n1172, n1171, n1170, n1169, n1168, n1167,
         n1166, n1165, n1164, n1163, n1162, n1161, n1160, n1159, n1158, n1157,
         n1156, n1155, n1154, n1153, n1152, n1151, n1150, n1149, n1148, n1147,
         n1146, n1145, n1144, n1143, n1142, n1141, n1140, n1139, n1138, n1137,
         n1136, n1135, n1134, n1133, n1132, n1131, n1130, n1129, n1128, n1127,
         n1126, n1125, n1124, n1123, n1122, n1121, n1120, n1119, n1118, n1117,
         n1116, n1115, n1114, n1113, n1112, n1111, n1110, n1109, n1108, n1107,
         n1106, n1105, n1104, n1103, n1102, n1101, n1100, n1099, n1098, n1097,
         n1096, n1095, n1094, n1093, n1092, n1091, n1090, n1089, n1088, n1087,
         n1086, n1085, n1084, n1083, n1082, n1081, n1080, n1079, n1078, n1077,
         n1076, n1075, n1074, n1073, n1072, n1071, n1070, n1069, n1068, n1067,
         n1066, n1065, n1064, n1063, n1062, n1061, n1060, n1059, n1058, n1057,
         n1056, n1055, n1054, n1053, n1052, n1051, n1050, n1049, n1048, n1047,
         n1046, n1045, n1044, n1043, n1042, n1041, n1040, n1039, n1038, n1037,
         n1036, n1035, n1034, n1033, n1032, n1031, n1030, n1029, n1028, n1027,
         n1026, n1025, n1024, n1023, n1022, n1021, n1020, n1019, n1018, n1017,
         n1016, n1015, n1014, n1013, n1012, n1011, n1010, n1009, n1008, n1007,
         n1006, n1005, n1004, n1003, n1002, n1001, n1000, n5886, n5887, n5888,
         n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898,
         n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908,
         n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918,
         n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928,
         n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938,
         n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948,
         n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958,
         n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968,
         n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978,
         n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988,
         n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998,
         n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008,
         n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018,
         n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028,
         n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038,
         n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048,
         n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058,
         n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068,
         n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078,
         n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088,
         n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098,
         n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108,
         n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118,
         n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128,
         n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138,
         n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148,
         n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158,
         n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168,
         n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178,
         n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188,
         n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198,
         n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208,
         n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218,
         n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228,
         n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238,
         n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248,
         n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258,
         n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268,
         n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278,
         n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288,
         n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298,
         n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308,
         n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318,
         n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328,
         n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338,
         n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348,
         n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358,
         n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368,
         n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378,
         n6379, n6380, n6381, n6382, n6383, n6384, n6386, n6388, n6390, n6392,
         n6394, n6396, n6398, n6400, n6402, n6404, n6406, n6408, n6410, n6412,
         n6414, n6416, n6418, n6420, n6422, n6424, n6426, n6428, n6430, n6432,
         n6434, n6436, n6438, n6440, n6442, n6444, n6446, n6448, n6450, n6452,
         n6454, n6456, n6458, n6460, n6462, n6464, n6466, n6468, n6470, n6472,
         n6474, n6476, n6478, n6480, n6482, n6484, n6486, n6488, n6490, n6492,
         n6494, n6496, n6498, n6500, n6502, n6504, n6506, n6508, n6510, n6512,
         n6514, n6516, n6518, n6520, n6522, n6524, n6526, n6528, n6530, n6532,
         n6534, n6536, n6538, n6540, n6542, n6544, n6546, n6548, n6550, n6552,
         n6554, n6556, n6558, n6560, n6562, n6564, n6566, n6568, n6570, n6572,
         n6574, n6576, n6578, n6580, n6582, n6584, n6586, n6588, n6590, n6592,
         n6594, n6596, n6598, n6600, n6602, n6604, n6606, n6608, n6610, n6612,
         n6614, n6616, n6618, n6620, n6622, n6624, n6626, n6628, n6630, n6632,
         n6634, n6636, n6638, n6640, n6642, n6644, n6646, n6648, n6650, n6652,
         n6654, n6656, n6658, n6660, n6662, n6664, n6666, n6668, n6670, n6672,
         n6674, n6676, n6678, n6680, n6682, n6684, n6686, n6688, n6690, n6692,
         n6694, n6696, n6698, n6700, n6702, n6704, n6706, n6708, n6710, n6712,
         n6714, n6716, n6718, n6720, n6722, n6724, n6726, n6728, n6730, n6732,
         n6734, n6736, n6738, n6740, n6742, n6744, n6746, n6748, n6750, n6752,
         n6754, n6756, n6758, n6760, n6762, n6764, n6766, n6768, n6770, n6772,
         n6774, n6776, n6778, n6780, n6782, n6784, n6786, n6788, n6790, n6792,
         n6794, n6796, n6798, n6800, n6802, n6804, n6806, n6808, n6810, n6812,
         n6814, n6816, n6818, n6820, n6822, n6824, n6826, n6828, n6830, n6832,
         n6834, n6836, n6838, n6840, n6842, n6844, n6846, n6848, n6850, n6852,
         n6854, n6856, n6858, n6860, n6862, n6864, n6866, n6868, n6870, n6872,
         n6874, n6876, n6878, n6880, n6882, n6884, n6886, n6888, n6890, n6892,
         n6894, n6896, n6898, n6900, n6902, n6904, n6906, n6908, n6910, n6912,
         n6914, n6916, n6918, n6920, n6922, n6924, n6926, n6928, n6930, n6932,
         n6934, n6936, n6938, n6940, n6942, n6944, n6946, n6948, n6950, n6952,
         n6954, n6956, n6958, n6960, n6962, n6964, n6966, n6968, n6970, n6972,
         n6974, n6976, n6978, n6980, n6982, n6984, n6986, n6988, n6990, n6992,
         n6994, n6996, n6998, n7000, n7002, n7004, n7006, n7008, n7010, n7012,
         n7014, n7016, n7018, n7020, n7022, n7024, n7025, n7026, n7027, n7028,
         n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038,
         n7039, n7040, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049,
         n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059,
         n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069,
         n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079,
         n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089,
         n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099,
         n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109,
         n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119,
         n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129,
         n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139,
         n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149,
         n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159,
         n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169,
         n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179,
         n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189,
         n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199,
         n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209,
         n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219,
         n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229,
         n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239,
         n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249,
         n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259,
         n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269,
         n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279,
         n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289,
         n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299,
         n7300, n7301, n7302, n7303, n7304, n7305, n7307, n7308, n7309, n7310,
         n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320,
         n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330,
         n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340,
         n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350,
         n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360,
         n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370,
         n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380,
         n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390,
         n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400,
         n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410,
         n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420,
         n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430,
         n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440,
         n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450,
         n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460,
         n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470,
         n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480,
         n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490,
         n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500,
         n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510,
         n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520,
         n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530,
         n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540,
         n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550,
         n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560,
         n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570,
         n7571, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996,
         n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006,
         n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016,
         n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026,
         n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036,
         n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046,
         n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056,
         n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066,
         n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076,
         n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086,
         n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096,
         n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106,
         n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116,
         n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126,
         n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136,
         n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146,
         n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156,
         n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166,
         n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176,
         n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186,
         n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196,
         n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206,
         n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216,
         n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226,
         n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236,
         n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246,
         n9247;
  wire   [31:0] \update_mask_0/reg_i_mask ;

  dff_sg \state_reg[0]  ( .D(n20), .CP(clk), .Q(n9569) );
  dff_sg \state_reg[1]  ( .D(n19), .CP(clk), .Q(n9568) );
  dff_sg \update_mask_0/o_pointer_reg[3]  ( .D(\update_mask_0/n1128 ), .CP(clk), .Q(\update_mask_0/N31 ) );
  dff_sg \update_mask_0/o_pointer_reg[2]  ( .D(n5879), .CP(clk), .Q(
        \update_mask_0/N30 ) );
  dff_sg \update_mask_0/o_pointer_reg[1]  ( .D(n5878), .CP(clk), .Q(
        \update_mask_0/N29 ) );
  dff_sg \update_mask_0/o_pointer_reg[0]  ( .D(n5880), .CP(clk), .Q(
        \update_mask_0/N28 ) );
  dff_sg \update_mask_0/m_pointer_reg[1]  ( .D(n5883), .CP(clk), .Q(
        \update_mask_0/N24 ) );
  dff_sg \update_mask_0/m_pointer_reg[2]  ( .D(n5882), .CP(clk), .Q(
        \update_mask_0/N25 ) );
  dff_sg \update_mask_0/m_pointer_reg[3]  ( .D(n5884), .CP(clk), .Q(
        \update_mask_0/N26 ) );
  dff_sg \update_mask_0/reg_i_mask_reg[0]  ( .D(\update_mask_0/n1480 ), .CP(
        clk), .Q(\update_mask_0/reg_i_mask [0]) );
  dff_sg \update_mask_0/reg_i_mask_reg[1]  ( .D(\update_mask_0/n1479 ), .CP(
        clk), .Q(\update_mask_0/reg_i_mask [1]) );
  dff_sg \update_mask_0/reg_i_mask_reg[2]  ( .D(\update_mask_0/n1478 ), .CP(
        clk), .Q(\update_mask_0/reg_i_mask [2]) );
  dff_sg \update_mask_0/reg_i_mask_reg[3]  ( .D(\update_mask_0/n1477 ), .CP(
        clk), .Q(\update_mask_0/reg_i_mask [3]) );
  dff_sg \update_mask_0/reg_i_mask_reg[4]  ( .D(\update_mask_0/n1476 ), .CP(
        clk), .Q(\update_mask_0/reg_i_mask [4]) );
  dff_sg \update_mask_0/reg_i_mask_reg[5]  ( .D(\update_mask_0/n1475 ), .CP(
        clk), .Q(\update_mask_0/reg_i_mask [5]) );
  dff_sg \update_mask_0/reg_i_mask_reg[6]  ( .D(\update_mask_0/n1474 ), .CP(
        clk), .Q(\update_mask_0/reg_i_mask [6]) );
  dff_sg \update_mask_0/reg_i_mask_reg[7]  ( .D(\update_mask_0/n1473 ), .CP(
        clk), .Q(\update_mask_0/reg_i_mask [7]) );
  dff_sg \update_mask_0/reg_i_mask_reg[8]  ( .D(\update_mask_0/n1472 ), .CP(
        clk), .Q(\update_mask_0/reg_i_mask [8]) );
  dff_sg \update_mask_0/reg_i_mask_reg[9]  ( .D(\update_mask_0/n1471 ), .CP(
        clk), .Q(\update_mask_0/reg_i_mask [9]) );
  dff_sg \update_mask_0/reg_i_mask_reg[10]  ( .D(\update_mask_0/n1470 ), .CP(
        clk), .Q(\update_mask_0/reg_i_mask [10]) );
  dff_sg \update_mask_0/reg_i_mask_reg[11]  ( .D(\update_mask_0/n1469 ), .CP(
        clk), .Q(\update_mask_0/reg_i_mask [11]) );
  dff_sg \update_mask_0/reg_i_mask_reg[12]  ( .D(\update_mask_0/n1468 ), .CP(
        clk), .Q(\update_mask_0/reg_i_mask [12]) );
  dff_sg \update_mask_0/reg_i_mask_reg[13]  ( .D(\update_mask_0/n1467 ), .CP(
        clk), .Q(\update_mask_0/reg_i_mask [13]) );
  dff_sg \update_mask_0/reg_i_mask_reg[14]  ( .D(\update_mask_0/n1466 ), .CP(
        clk), .Q(\update_mask_0/reg_i_mask [14]) );
  dff_sg \update_mask_0/reg_i_mask_reg[15]  ( .D(\update_mask_0/n1465 ), .CP(
        clk), .Q(\update_mask_0/reg_i_mask [15]) );
  dff_sg \update_mask_0/reg_i_mask_reg[16]  ( .D(\update_mask_0/n1464 ), .CP(
        clk), .Q(\update_mask_0/reg_i_mask [16]) );
  dff_sg \update_mask_0/reg_i_mask_reg[17]  ( .D(\update_mask_0/n1463 ), .CP(
        clk), .Q(\update_mask_0/reg_i_mask [17]) );
  dff_sg \update_mask_0/reg_i_mask_reg[18]  ( .D(\update_mask_0/n1462 ), .CP(
        clk), .Q(\update_mask_0/reg_i_mask [18]) );
  dff_sg \update_mask_0/reg_i_mask_reg[19]  ( .D(\update_mask_0/n1461 ), .CP(
        clk), .Q(\update_mask_0/reg_i_mask [19]) );
  dff_sg \update_mask_0/reg_i_mask_reg[20]  ( .D(\update_mask_0/n1460 ), .CP(
        clk), .Q(\update_mask_0/reg_i_mask [20]) );
  dff_sg \update_mask_0/reg_i_mask_reg[21]  ( .D(\update_mask_0/n1459 ), .CP(
        clk), .Q(\update_mask_0/reg_i_mask [21]) );
  dff_sg \update_mask_0/reg_i_mask_reg[22]  ( .D(\update_mask_0/n1458 ), .CP(
        clk), .Q(\update_mask_0/reg_i_mask [22]) );
  dff_sg \update_mask_0/reg_i_mask_reg[23]  ( .D(\update_mask_0/n1457 ), .CP(
        clk), .Q(\update_mask_0/reg_i_mask [23]) );
  dff_sg \update_mask_0/reg_i_mask_reg[24]  ( .D(\update_mask_0/n1456 ), .CP(
        clk), .Q(\update_mask_0/reg_i_mask [24]) );
  dff_sg \update_mask_0/reg_i_mask_reg[25]  ( .D(\update_mask_0/n1455 ), .CP(
        clk), .Q(\update_mask_0/reg_i_mask [25]) );
  dff_sg \update_mask_0/reg_i_mask_reg[26]  ( .D(\update_mask_0/n1454 ), .CP(
        clk), .Q(\update_mask_0/reg_i_mask [26]) );
  dff_sg \update_mask_0/reg_i_mask_reg[27]  ( .D(\update_mask_0/n1453 ), .CP(
        clk), .Q(\update_mask_0/reg_i_mask [27]) );
  dff_sg \update_mask_0/reg_i_mask_reg[28]  ( .D(\update_mask_0/n1452 ), .CP(
        clk), .Q(\update_mask_0/reg_i_mask [28]) );
  dff_sg \update_mask_0/reg_i_mask_reg[29]  ( .D(\update_mask_0/n1451 ), .CP(
        clk), .Q(\update_mask_0/reg_i_mask [29]) );
  dff_sg \update_mask_0/reg_i_mask_reg[30]  ( .D(\update_mask_0/n1450 ), .CP(
        clk), .Q(\update_mask_0/reg_i_mask [30]) );
  dff_sg \update_mask_0/reg_i_mask_reg[31]  ( .D(\update_mask_0/n1449 ), .CP(
        clk), .Q(\update_mask_0/reg_i_mask [31]) );
  dff_sg \update_mask_0/reg_out_reg[0][0]  ( .D(\update_mask_0/n1448 ), .CP(
        clk), .Q(\update_mask_0/reg_out[0][0] ) );
  dff_sg \update_mask_0/reg_out_reg[0][1]  ( .D(\update_mask_0/n1447 ), .CP(
        clk), .Q(\update_mask_0/reg_out[0][1] ) );
  dff_sg \update_mask_0/reg_out_reg[0][2]  ( .D(\update_mask_0/n1446 ), .CP(
        clk), .Q(\update_mask_0/reg_out[0][2] ) );
  dff_sg \update_mask_0/reg_out_reg[0][3]  ( .D(\update_mask_0/n1445 ), .CP(
        clk), .Q(\update_mask_0/reg_out[0][3] ) );
  dff_sg \update_mask_0/reg_out_reg[0][4]  ( .D(\update_mask_0/n1444 ), .CP(
        clk), .Q(\update_mask_0/reg_out[0][4] ) );
  dff_sg \update_mask_0/reg_out_reg[0][5]  ( .D(\update_mask_0/n1443 ), .CP(
        clk), .Q(\update_mask_0/reg_out[0][5] ) );
  dff_sg \update_mask_0/reg_out_reg[0][6]  ( .D(\update_mask_0/n1442 ), .CP(
        clk), .Q(\update_mask_0/reg_out[0][6] ) );
  dff_sg \update_mask_0/reg_out_reg[0][7]  ( .D(\update_mask_0/n1441 ), .CP(
        clk), .Q(\update_mask_0/reg_out[0][7] ) );
  dff_sg \update_mask_0/reg_out_reg[0][8]  ( .D(\update_mask_0/n1440 ), .CP(
        clk), .Q(\update_mask_0/reg_out[0][8] ) );
  dff_sg \update_mask_0/reg_out_reg[0][9]  ( .D(\update_mask_0/n1439 ), .CP(
        clk), .Q(\update_mask_0/reg_out[0][9] ) );
  dff_sg \update_mask_0/reg_out_reg[0][10]  ( .D(\update_mask_0/n1438 ), .CP(
        clk), .Q(\update_mask_0/reg_out[0][10] ) );
  dff_sg \update_mask_0/reg_out_reg[0][11]  ( .D(\update_mask_0/n1437 ), .CP(
        clk), .Q(\update_mask_0/reg_out[0][11] ) );
  dff_sg \update_mask_0/reg_out_reg[0][12]  ( .D(\update_mask_0/n1436 ), .CP(
        clk), .Q(\update_mask_0/reg_out[0][12] ) );
  dff_sg \update_mask_0/reg_out_reg[0][13]  ( .D(\update_mask_0/n1435 ), .CP(
        clk), .Q(\update_mask_0/reg_out[0][13] ) );
  dff_sg \update_mask_0/reg_out_reg[0][14]  ( .D(\update_mask_0/n1434 ), .CP(
        clk), .Q(\update_mask_0/reg_out[0][14] ) );
  dff_sg \update_mask_0/reg_out_reg[0][15]  ( .D(\update_mask_0/n1433 ), .CP(
        clk), .Q(\update_mask_0/reg_out[0][15] ) );
  dff_sg \update_mask_0/reg_out_reg[0][16]  ( .D(\update_mask_0/n1432 ), .CP(
        clk), .Q(\update_mask_0/reg_out[0][16] ) );
  dff_sg \update_mask_0/reg_out_reg[0][17]  ( .D(\update_mask_0/n1431 ), .CP(
        clk), .Q(\update_mask_0/reg_out[0][17] ) );
  dff_sg \update_mask_0/reg_out_reg[0][18]  ( .D(\update_mask_0/n1430 ), .CP(
        clk), .Q(\update_mask_0/reg_out[0][18] ) );
  dff_sg \update_mask_0/reg_out_reg[0][19]  ( .D(\update_mask_0/n1429 ), .CP(
        clk), .Q(\update_mask_0/reg_out[0][19] ) );
  dff_sg \update_mask_0/reg_out_reg[1][0]  ( .D(\update_mask_0/n1428 ), .CP(
        clk), .Q(\update_mask_0/reg_out[1][0] ) );
  dff_sg \update_mask_0/reg_out_reg[1][1]  ( .D(\update_mask_0/n1427 ), .CP(
        clk), .Q(\update_mask_0/reg_out[1][1] ) );
  dff_sg \update_mask_0/reg_out_reg[1][2]  ( .D(\update_mask_0/n1426 ), .CP(
        clk), .Q(\update_mask_0/reg_out[1][2] ) );
  dff_sg \update_mask_0/reg_out_reg[1][3]  ( .D(\update_mask_0/n1425 ), .CP(
        clk), .Q(\update_mask_0/reg_out[1][3] ) );
  dff_sg \update_mask_0/reg_out_reg[1][4]  ( .D(\update_mask_0/n1424 ), .CP(
        clk), .Q(\update_mask_0/reg_out[1][4] ) );
  dff_sg \update_mask_0/reg_out_reg[1][5]  ( .D(\update_mask_0/n1423 ), .CP(
        clk), .Q(\update_mask_0/reg_out[1][5] ) );
  dff_sg \update_mask_0/reg_out_reg[1][6]  ( .D(\update_mask_0/n1422 ), .CP(
        clk), .Q(\update_mask_0/reg_out[1][6] ) );
  dff_sg \update_mask_0/reg_out_reg[1][7]  ( .D(\update_mask_0/n1421 ), .CP(
        clk), .Q(\update_mask_0/reg_out[1][7] ) );
  dff_sg \update_mask_0/reg_out_reg[1][8]  ( .D(\update_mask_0/n1420 ), .CP(
        clk), .Q(\update_mask_0/reg_out[1][8] ) );
  dff_sg \update_mask_0/reg_out_reg[1][9]  ( .D(\update_mask_0/n1419 ), .CP(
        clk), .Q(\update_mask_0/reg_out[1][9] ) );
  dff_sg \update_mask_0/reg_out_reg[1][10]  ( .D(\update_mask_0/n1418 ), .CP(
        clk), .Q(\update_mask_0/reg_out[1][10] ) );
  dff_sg \update_mask_0/reg_out_reg[1][11]  ( .D(\update_mask_0/n1417 ), .CP(
        clk), .Q(\update_mask_0/reg_out[1][11] ) );
  dff_sg \update_mask_0/reg_out_reg[1][12]  ( .D(\update_mask_0/n1416 ), .CP(
        clk), .Q(\update_mask_0/reg_out[1][12] ) );
  dff_sg \update_mask_0/reg_out_reg[1][13]  ( .D(\update_mask_0/n1415 ), .CP(
        clk), .Q(\update_mask_0/reg_out[1][13] ) );
  dff_sg \update_mask_0/reg_out_reg[1][14]  ( .D(\update_mask_0/n1414 ), .CP(
        clk), .Q(\update_mask_0/reg_out[1][14] ) );
  dff_sg \update_mask_0/reg_out_reg[1][15]  ( .D(\update_mask_0/n1413 ), .CP(
        clk), .Q(\update_mask_0/reg_out[1][15] ) );
  dff_sg \update_mask_0/reg_out_reg[1][16]  ( .D(\update_mask_0/n1412 ), .CP(
        clk), .Q(\update_mask_0/reg_out[1][16] ) );
  dff_sg \update_mask_0/reg_out_reg[1][17]  ( .D(\update_mask_0/n1411 ), .CP(
        clk), .Q(\update_mask_0/reg_out[1][17] ) );
  dff_sg \update_mask_0/reg_out_reg[1][18]  ( .D(\update_mask_0/n1410 ), .CP(
        clk), .Q(\update_mask_0/reg_out[1][18] ) );
  dff_sg \update_mask_0/reg_out_reg[1][19]  ( .D(\update_mask_0/n1409 ), .CP(
        clk), .Q(\update_mask_0/reg_out[1][19] ) );
  dff_sg \update_mask_0/reg_out_reg[2][0]  ( .D(\update_mask_0/n1408 ), .CP(
        clk), .Q(\update_mask_0/reg_out[2][0] ) );
  dff_sg \update_mask_0/reg_out_reg[2][1]  ( .D(\update_mask_0/n1407 ), .CP(
        clk), .Q(\update_mask_0/reg_out[2][1] ) );
  dff_sg \update_mask_0/reg_out_reg[2][2]  ( .D(\update_mask_0/n1406 ), .CP(
        clk), .Q(\update_mask_0/reg_out[2][2] ) );
  dff_sg \update_mask_0/reg_out_reg[2][3]  ( .D(\update_mask_0/n1405 ), .CP(
        clk), .Q(\update_mask_0/reg_out[2][3] ) );
  dff_sg \update_mask_0/reg_out_reg[2][4]  ( .D(\update_mask_0/n1404 ), .CP(
        clk), .Q(\update_mask_0/reg_out[2][4] ) );
  dff_sg \update_mask_0/reg_out_reg[2][5]  ( .D(\update_mask_0/n1403 ), .CP(
        clk), .Q(\update_mask_0/reg_out[2][5] ) );
  dff_sg \update_mask_0/reg_out_reg[2][6]  ( .D(\update_mask_0/n1402 ), .CP(
        clk), .Q(\update_mask_0/reg_out[2][6] ) );
  dff_sg \update_mask_0/reg_out_reg[2][7]  ( .D(\update_mask_0/n1401 ), .CP(
        clk), .Q(\update_mask_0/reg_out[2][7] ) );
  dff_sg \update_mask_0/reg_out_reg[2][8]  ( .D(\update_mask_0/n1400 ), .CP(
        clk), .Q(\update_mask_0/reg_out[2][8] ) );
  dff_sg \update_mask_0/reg_out_reg[2][9]  ( .D(\update_mask_0/n1399 ), .CP(
        clk), .Q(\update_mask_0/reg_out[2][9] ) );
  dff_sg \update_mask_0/reg_out_reg[2][10]  ( .D(\update_mask_0/n1398 ), .CP(
        clk), .Q(\update_mask_0/reg_out[2][10] ) );
  dff_sg \update_mask_0/reg_out_reg[2][11]  ( .D(\update_mask_0/n1397 ), .CP(
        clk), .Q(\update_mask_0/reg_out[2][11] ) );
  dff_sg \update_mask_0/reg_out_reg[2][12]  ( .D(\update_mask_0/n1396 ), .CP(
        clk), .Q(\update_mask_0/reg_out[2][12] ) );
  dff_sg \update_mask_0/reg_out_reg[2][13]  ( .D(\update_mask_0/n1395 ), .CP(
        clk), .Q(\update_mask_0/reg_out[2][13] ) );
  dff_sg \update_mask_0/reg_out_reg[2][14]  ( .D(\update_mask_0/n1394 ), .CP(
        clk), .Q(\update_mask_0/reg_out[2][14] ) );
  dff_sg \update_mask_0/reg_out_reg[2][15]  ( .D(\update_mask_0/n1393 ), .CP(
        clk), .Q(\update_mask_0/reg_out[2][15] ) );
  dff_sg \update_mask_0/reg_out_reg[2][16]  ( .D(\update_mask_0/n1392 ), .CP(
        clk), .Q(\update_mask_0/reg_out[2][16] ) );
  dff_sg \update_mask_0/reg_out_reg[2][17]  ( .D(\update_mask_0/n1391 ), .CP(
        clk), .Q(\update_mask_0/reg_out[2][17] ) );
  dff_sg \update_mask_0/reg_out_reg[2][18]  ( .D(\update_mask_0/n1390 ), .CP(
        clk), .Q(\update_mask_0/reg_out[2][18] ) );
  dff_sg \update_mask_0/reg_out_reg[2][19]  ( .D(\update_mask_0/n1389 ), .CP(
        clk), .Q(\update_mask_0/reg_out[2][19] ) );
  dff_sg \update_mask_0/reg_out_reg[3][0]  ( .D(\update_mask_0/n1388 ), .CP(
        clk), .Q(\update_mask_0/reg_out[3][0] ) );
  dff_sg \update_mask_0/reg_out_reg[3][1]  ( .D(\update_mask_0/n1387 ), .CP(
        clk), .Q(\update_mask_0/reg_out[3][1] ) );
  dff_sg \update_mask_0/reg_out_reg[3][2]  ( .D(\update_mask_0/n1386 ), .CP(
        clk), .Q(\update_mask_0/reg_out[3][2] ) );
  dff_sg \update_mask_0/reg_out_reg[3][3]  ( .D(\update_mask_0/n1385 ), .CP(
        clk), .Q(\update_mask_0/reg_out[3][3] ) );
  dff_sg \update_mask_0/reg_out_reg[3][4]  ( .D(\update_mask_0/n1384 ), .CP(
        clk), .Q(\update_mask_0/reg_out[3][4] ) );
  dff_sg \update_mask_0/reg_out_reg[3][5]  ( .D(\update_mask_0/n1383 ), .CP(
        clk), .Q(\update_mask_0/reg_out[3][5] ) );
  dff_sg \update_mask_0/reg_out_reg[3][6]  ( .D(\update_mask_0/n1382 ), .CP(
        clk), .Q(\update_mask_0/reg_out[3][6] ) );
  dff_sg \update_mask_0/reg_out_reg[3][7]  ( .D(\update_mask_0/n1381 ), .CP(
        clk), .Q(\update_mask_0/reg_out[3][7] ) );
  dff_sg \update_mask_0/reg_out_reg[3][8]  ( .D(\update_mask_0/n1380 ), .CP(
        clk), .Q(\update_mask_0/reg_out[3][8] ) );
  dff_sg \update_mask_0/reg_out_reg[3][9]  ( .D(\update_mask_0/n1379 ), .CP(
        clk), .Q(\update_mask_0/reg_out[3][9] ) );
  dff_sg \update_mask_0/reg_out_reg[3][10]  ( .D(\update_mask_0/n1378 ), .CP(
        clk), .Q(\update_mask_0/reg_out[3][10] ) );
  dff_sg \update_mask_0/reg_out_reg[3][11]  ( .D(\update_mask_0/n1377 ), .CP(
        clk), .Q(\update_mask_0/reg_out[3][11] ) );
  dff_sg \update_mask_0/reg_out_reg[3][12]  ( .D(\update_mask_0/n1376 ), .CP(
        clk), .Q(\update_mask_0/reg_out[3][12] ) );
  dff_sg \update_mask_0/reg_out_reg[3][13]  ( .D(\update_mask_0/n1375 ), .CP(
        clk), .Q(\update_mask_0/reg_out[3][13] ) );
  dff_sg \update_mask_0/reg_out_reg[3][14]  ( .D(\update_mask_0/n1374 ), .CP(
        clk), .Q(\update_mask_0/reg_out[3][14] ) );
  dff_sg \update_mask_0/reg_out_reg[3][15]  ( .D(\update_mask_0/n1373 ), .CP(
        clk), .Q(\update_mask_0/reg_out[3][15] ) );
  dff_sg \update_mask_0/reg_out_reg[3][16]  ( .D(\update_mask_0/n1372 ), .CP(
        clk), .Q(\update_mask_0/reg_out[3][16] ) );
  dff_sg \update_mask_0/reg_out_reg[3][17]  ( .D(\update_mask_0/n1371 ), .CP(
        clk), .Q(\update_mask_0/reg_out[3][17] ) );
  dff_sg \update_mask_0/reg_out_reg[3][18]  ( .D(\update_mask_0/n1370 ), .CP(
        clk), .Q(\update_mask_0/reg_out[3][18] ) );
  dff_sg \update_mask_0/reg_out_reg[3][19]  ( .D(\update_mask_0/n1369 ), .CP(
        clk), .Q(\update_mask_0/reg_out[3][19] ) );
  dff_sg \update_mask_0/reg_out_reg[4][0]  ( .D(\update_mask_0/n1368 ), .CP(
        clk), .Q(\update_mask_0/reg_out[4][0] ) );
  dff_sg \update_mask_0/reg_out_reg[4][1]  ( .D(\update_mask_0/n1367 ), .CP(
        clk), .Q(\update_mask_0/reg_out[4][1] ) );
  dff_sg \update_mask_0/reg_out_reg[4][2]  ( .D(\update_mask_0/n1366 ), .CP(
        clk), .Q(\update_mask_0/reg_out[4][2] ) );
  dff_sg \update_mask_0/reg_out_reg[4][3]  ( .D(\update_mask_0/n1365 ), .CP(
        clk), .Q(\update_mask_0/reg_out[4][3] ) );
  dff_sg \update_mask_0/reg_out_reg[4][4]  ( .D(\update_mask_0/n1364 ), .CP(
        clk), .Q(\update_mask_0/reg_out[4][4] ) );
  dff_sg \update_mask_0/reg_out_reg[4][5]  ( .D(\update_mask_0/n1363 ), .CP(
        clk), .Q(\update_mask_0/reg_out[4][5] ) );
  dff_sg \update_mask_0/reg_out_reg[4][6]  ( .D(\update_mask_0/n1362 ), .CP(
        clk), .Q(\update_mask_0/reg_out[4][6] ) );
  dff_sg \update_mask_0/reg_out_reg[4][7]  ( .D(\update_mask_0/n1361 ), .CP(
        clk), .Q(\update_mask_0/reg_out[4][7] ) );
  dff_sg \update_mask_0/reg_out_reg[4][8]  ( .D(\update_mask_0/n1360 ), .CP(
        clk), .Q(\update_mask_0/reg_out[4][8] ) );
  dff_sg \update_mask_0/reg_out_reg[4][9]  ( .D(\update_mask_0/n1359 ), .CP(
        clk), .Q(\update_mask_0/reg_out[4][9] ) );
  dff_sg \update_mask_0/reg_out_reg[4][10]  ( .D(\update_mask_0/n1358 ), .CP(
        clk), .Q(\update_mask_0/reg_out[4][10] ) );
  dff_sg \update_mask_0/reg_out_reg[4][11]  ( .D(\update_mask_0/n1357 ), .CP(
        clk), .Q(\update_mask_0/reg_out[4][11] ) );
  dff_sg \update_mask_0/reg_out_reg[4][12]  ( .D(\update_mask_0/n1356 ), .CP(
        clk), .Q(\update_mask_0/reg_out[4][12] ) );
  dff_sg \update_mask_0/reg_out_reg[4][13]  ( .D(\update_mask_0/n1355 ), .CP(
        clk), .Q(\update_mask_0/reg_out[4][13] ) );
  dff_sg \update_mask_0/reg_out_reg[4][14]  ( .D(\update_mask_0/n1354 ), .CP(
        clk), .Q(\update_mask_0/reg_out[4][14] ) );
  dff_sg \update_mask_0/reg_out_reg[4][15]  ( .D(\update_mask_0/n1353 ), .CP(
        clk), .Q(\update_mask_0/reg_out[4][15] ) );
  dff_sg \update_mask_0/reg_out_reg[4][16]  ( .D(\update_mask_0/n1352 ), .CP(
        clk), .Q(\update_mask_0/reg_out[4][16] ) );
  dff_sg \update_mask_0/reg_out_reg[4][17]  ( .D(\update_mask_0/n1351 ), .CP(
        clk), .Q(\update_mask_0/reg_out[4][17] ) );
  dff_sg \update_mask_0/reg_out_reg[4][18]  ( .D(\update_mask_0/n1350 ), .CP(
        clk), .Q(\update_mask_0/reg_out[4][18] ) );
  dff_sg \update_mask_0/reg_out_reg[4][19]  ( .D(\update_mask_0/n1349 ), .CP(
        clk), .Q(\update_mask_0/reg_out[4][19] ) );
  dff_sg \update_mask_0/reg_out_reg[5][0]  ( .D(\update_mask_0/n1348 ), .CP(
        clk), .Q(\update_mask_0/reg_out[5][0] ) );
  dff_sg \update_mask_0/reg_out_reg[5][1]  ( .D(\update_mask_0/n1347 ), .CP(
        clk), .Q(\update_mask_0/reg_out[5][1] ) );
  dff_sg \update_mask_0/reg_out_reg[5][2]  ( .D(\update_mask_0/n1346 ), .CP(
        clk), .Q(\update_mask_0/reg_out[5][2] ) );
  dff_sg \update_mask_0/reg_out_reg[5][3]  ( .D(\update_mask_0/n1345 ), .CP(
        clk), .Q(\update_mask_0/reg_out[5][3] ) );
  dff_sg \update_mask_0/reg_out_reg[5][4]  ( .D(\update_mask_0/n1344 ), .CP(
        clk), .Q(\update_mask_0/reg_out[5][4] ) );
  dff_sg \update_mask_0/reg_out_reg[5][5]  ( .D(\update_mask_0/n1343 ), .CP(
        clk), .Q(\update_mask_0/reg_out[5][5] ) );
  dff_sg \update_mask_0/reg_out_reg[5][6]  ( .D(\update_mask_0/n1342 ), .CP(
        clk), .Q(\update_mask_0/reg_out[5][6] ) );
  dff_sg \update_mask_0/reg_out_reg[5][7]  ( .D(\update_mask_0/n1341 ), .CP(
        clk), .Q(\update_mask_0/reg_out[5][7] ) );
  dff_sg \update_mask_0/reg_out_reg[5][8]  ( .D(\update_mask_0/n1340 ), .CP(
        clk), .Q(\update_mask_0/reg_out[5][8] ) );
  dff_sg \update_mask_0/reg_out_reg[5][9]  ( .D(\update_mask_0/n1339 ), .CP(
        clk), .Q(\update_mask_0/reg_out[5][9] ) );
  dff_sg \update_mask_0/reg_out_reg[5][10]  ( .D(\update_mask_0/n1338 ), .CP(
        clk), .Q(\update_mask_0/reg_out[5][10] ) );
  dff_sg \update_mask_0/reg_out_reg[5][11]  ( .D(\update_mask_0/n1337 ), .CP(
        clk), .Q(\update_mask_0/reg_out[5][11] ) );
  dff_sg \update_mask_0/reg_out_reg[5][12]  ( .D(\update_mask_0/n1336 ), .CP(
        clk), .Q(\update_mask_0/reg_out[5][12] ) );
  dff_sg \update_mask_0/reg_out_reg[5][13]  ( .D(\update_mask_0/n1335 ), .CP(
        clk), .Q(\update_mask_0/reg_out[5][13] ) );
  dff_sg \update_mask_0/reg_out_reg[5][14]  ( .D(\update_mask_0/n1334 ), .CP(
        clk), .Q(\update_mask_0/reg_out[5][14] ) );
  dff_sg \update_mask_0/reg_out_reg[5][15]  ( .D(\update_mask_0/n1333 ), .CP(
        clk), .Q(\update_mask_0/reg_out[5][15] ) );
  dff_sg \update_mask_0/reg_out_reg[5][16]  ( .D(\update_mask_0/n1332 ), .CP(
        clk), .Q(\update_mask_0/reg_out[5][16] ) );
  dff_sg \update_mask_0/reg_out_reg[5][17]  ( .D(\update_mask_0/n1331 ), .CP(
        clk), .Q(\update_mask_0/reg_out[5][17] ) );
  dff_sg \update_mask_0/reg_out_reg[5][18]  ( .D(\update_mask_0/n1330 ), .CP(
        clk), .Q(\update_mask_0/reg_out[5][18] ) );
  dff_sg \update_mask_0/reg_out_reg[5][19]  ( .D(\update_mask_0/n1329 ), .CP(
        clk), .Q(\update_mask_0/reg_out[5][19] ) );
  dff_sg \update_mask_0/reg_out_reg[6][0]  ( .D(\update_mask_0/n1328 ), .CP(
        clk), .Q(\update_mask_0/reg_out[6][0] ) );
  dff_sg \update_mask_0/reg_out_reg[6][1]  ( .D(\update_mask_0/n1327 ), .CP(
        clk), .Q(\update_mask_0/reg_out[6][1] ) );
  dff_sg \update_mask_0/reg_out_reg[6][2]  ( .D(\update_mask_0/n1326 ), .CP(
        clk), .Q(\update_mask_0/reg_out[6][2] ) );
  dff_sg \update_mask_0/reg_out_reg[6][3]  ( .D(\update_mask_0/n1325 ), .CP(
        clk), .Q(\update_mask_0/reg_out[6][3] ) );
  dff_sg \update_mask_0/reg_out_reg[6][4]  ( .D(\update_mask_0/n1324 ), .CP(
        clk), .Q(\update_mask_0/reg_out[6][4] ) );
  dff_sg \update_mask_0/reg_out_reg[6][5]  ( .D(\update_mask_0/n1323 ), .CP(
        clk), .Q(\update_mask_0/reg_out[6][5] ) );
  dff_sg \update_mask_0/reg_out_reg[6][6]  ( .D(\update_mask_0/n1322 ), .CP(
        clk), .Q(\update_mask_0/reg_out[6][6] ) );
  dff_sg \update_mask_0/reg_out_reg[6][7]  ( .D(\update_mask_0/n1321 ), .CP(
        clk), .Q(\update_mask_0/reg_out[6][7] ) );
  dff_sg \update_mask_0/reg_out_reg[6][8]  ( .D(\update_mask_0/n1320 ), .CP(
        clk), .Q(\update_mask_0/reg_out[6][8] ) );
  dff_sg \update_mask_0/reg_out_reg[6][9]  ( .D(\update_mask_0/n1319 ), .CP(
        clk), .Q(\update_mask_0/reg_out[6][9] ) );
  dff_sg \update_mask_0/reg_out_reg[6][10]  ( .D(\update_mask_0/n1318 ), .CP(
        clk), .Q(\update_mask_0/reg_out[6][10] ) );
  dff_sg \update_mask_0/reg_out_reg[6][11]  ( .D(\update_mask_0/n1317 ), .CP(
        clk), .Q(\update_mask_0/reg_out[6][11] ) );
  dff_sg \update_mask_0/reg_out_reg[6][12]  ( .D(\update_mask_0/n1316 ), .CP(
        clk), .Q(\update_mask_0/reg_out[6][12] ) );
  dff_sg \update_mask_0/reg_out_reg[6][13]  ( .D(\update_mask_0/n1315 ), .CP(
        clk), .Q(\update_mask_0/reg_out[6][13] ) );
  dff_sg \update_mask_0/reg_out_reg[6][14]  ( .D(\update_mask_0/n1314 ), .CP(
        clk), .Q(\update_mask_0/reg_out[6][14] ) );
  dff_sg \update_mask_0/reg_out_reg[6][15]  ( .D(\update_mask_0/n1313 ), .CP(
        clk), .Q(\update_mask_0/reg_out[6][15] ) );
  dff_sg \update_mask_0/reg_out_reg[6][16]  ( .D(\update_mask_0/n1312 ), .CP(
        clk), .Q(\update_mask_0/reg_out[6][16] ) );
  dff_sg \update_mask_0/reg_out_reg[6][17]  ( .D(\update_mask_0/n1311 ), .CP(
        clk), .Q(\update_mask_0/reg_out[6][17] ) );
  dff_sg \update_mask_0/reg_out_reg[6][18]  ( .D(\update_mask_0/n1310 ), .CP(
        clk), .Q(\update_mask_0/reg_out[6][18] ) );
  dff_sg \update_mask_0/reg_out_reg[6][19]  ( .D(\update_mask_0/n1309 ), .CP(
        clk), .Q(\update_mask_0/reg_out[6][19] ) );
  dff_sg \update_mask_0/reg_out_reg[7][0]  ( .D(\update_mask_0/n1308 ), .CP(
        clk), .Q(\update_mask_0/reg_out[7][0] ) );
  dff_sg \update_mask_0/reg_out_reg[7][1]  ( .D(\update_mask_0/n1307 ), .CP(
        clk), .Q(\update_mask_0/reg_out[7][1] ) );
  dff_sg \update_mask_0/reg_out_reg[7][2]  ( .D(\update_mask_0/n1306 ), .CP(
        clk), .Q(\update_mask_0/reg_out[7][2] ) );
  dff_sg \update_mask_0/reg_out_reg[7][3]  ( .D(\update_mask_0/n1305 ), .CP(
        clk), .Q(\update_mask_0/reg_out[7][3] ) );
  dff_sg \update_mask_0/reg_out_reg[7][4]  ( .D(\update_mask_0/n1304 ), .CP(
        clk), .Q(\update_mask_0/reg_out[7][4] ) );
  dff_sg \update_mask_0/reg_out_reg[7][5]  ( .D(\update_mask_0/n1303 ), .CP(
        clk), .Q(\update_mask_0/reg_out[7][5] ) );
  dff_sg \update_mask_0/reg_out_reg[7][6]  ( .D(\update_mask_0/n1302 ), .CP(
        clk), .Q(\update_mask_0/reg_out[7][6] ) );
  dff_sg \update_mask_0/reg_out_reg[7][7]  ( .D(\update_mask_0/n1301 ), .CP(
        clk), .Q(\update_mask_0/reg_out[7][7] ) );
  dff_sg \update_mask_0/reg_out_reg[7][8]  ( .D(\update_mask_0/n1300 ), .CP(
        clk), .Q(\update_mask_0/reg_out[7][8] ) );
  dff_sg \update_mask_0/reg_out_reg[7][9]  ( .D(\update_mask_0/n1299 ), .CP(
        clk), .Q(\update_mask_0/reg_out[7][9] ) );
  dff_sg \update_mask_0/reg_out_reg[7][10]  ( .D(\update_mask_0/n1298 ), .CP(
        clk), .Q(\update_mask_0/reg_out[7][10] ) );
  dff_sg \update_mask_0/reg_out_reg[7][11]  ( .D(\update_mask_0/n1297 ), .CP(
        clk), .Q(\update_mask_0/reg_out[7][11] ) );
  dff_sg \update_mask_0/reg_out_reg[7][12]  ( .D(\update_mask_0/n1296 ), .CP(
        clk), .Q(\update_mask_0/reg_out[7][12] ) );
  dff_sg \update_mask_0/reg_out_reg[7][13]  ( .D(\update_mask_0/n1295 ), .CP(
        clk), .Q(\update_mask_0/reg_out[7][13] ) );
  dff_sg \update_mask_0/reg_out_reg[7][14]  ( .D(\update_mask_0/n1294 ), .CP(
        clk), .Q(\update_mask_0/reg_out[7][14] ) );
  dff_sg \update_mask_0/reg_out_reg[7][15]  ( .D(\update_mask_0/n1293 ), .CP(
        clk), .Q(\update_mask_0/reg_out[7][15] ) );
  dff_sg \update_mask_0/reg_out_reg[7][16]  ( .D(\update_mask_0/n1292 ), .CP(
        clk), .Q(\update_mask_0/reg_out[7][16] ) );
  dff_sg \update_mask_0/reg_out_reg[7][17]  ( .D(\update_mask_0/n1291 ), .CP(
        clk), .Q(\update_mask_0/reg_out[7][17] ) );
  dff_sg \update_mask_0/reg_out_reg[7][18]  ( .D(\update_mask_0/n1290 ), .CP(
        clk), .Q(\update_mask_0/reg_out[7][18] ) );
  dff_sg \update_mask_0/reg_out_reg[7][19]  ( .D(\update_mask_0/n1289 ), .CP(
        clk), .Q(\update_mask_0/reg_out[7][19] ) );
  dff_sg \update_mask_0/reg_out_reg[8][0]  ( .D(\update_mask_0/n1288 ), .CP(
        clk), .Q(\update_mask_0/reg_out[8][0] ) );
  dff_sg \update_mask_0/reg_out_reg[8][1]  ( .D(\update_mask_0/n1287 ), .CP(
        clk), .Q(\update_mask_0/reg_out[8][1] ) );
  dff_sg \update_mask_0/reg_out_reg[8][2]  ( .D(\update_mask_0/n1286 ), .CP(
        clk), .Q(\update_mask_0/reg_out[8][2] ) );
  dff_sg \update_mask_0/reg_out_reg[8][3]  ( .D(\update_mask_0/n1285 ), .CP(
        clk), .Q(\update_mask_0/reg_out[8][3] ) );
  dff_sg \update_mask_0/reg_out_reg[8][4]  ( .D(\update_mask_0/n1284 ), .CP(
        clk), .Q(\update_mask_0/reg_out[8][4] ) );
  dff_sg \update_mask_0/reg_out_reg[8][5]  ( .D(\update_mask_0/n1283 ), .CP(
        clk), .Q(\update_mask_0/reg_out[8][5] ) );
  dff_sg \update_mask_0/reg_out_reg[8][6]  ( .D(\update_mask_0/n1282 ), .CP(
        clk), .Q(\update_mask_0/reg_out[8][6] ) );
  dff_sg \update_mask_0/reg_out_reg[8][7]  ( .D(\update_mask_0/n1281 ), .CP(
        clk), .Q(\update_mask_0/reg_out[8][7] ) );
  dff_sg \update_mask_0/reg_out_reg[8][8]  ( .D(\update_mask_0/n1280 ), .CP(
        clk), .Q(\update_mask_0/reg_out[8][8] ) );
  dff_sg \update_mask_0/reg_out_reg[8][9]  ( .D(\update_mask_0/n1279 ), .CP(
        clk), .Q(\update_mask_0/reg_out[8][9] ) );
  dff_sg \update_mask_0/reg_out_reg[8][10]  ( .D(\update_mask_0/n1278 ), .CP(
        clk), .Q(\update_mask_0/reg_out[8][10] ) );
  dff_sg \update_mask_0/reg_out_reg[8][11]  ( .D(\update_mask_0/n1277 ), .CP(
        clk), .Q(\update_mask_0/reg_out[8][11] ) );
  dff_sg \update_mask_0/reg_out_reg[8][12]  ( .D(\update_mask_0/n1276 ), .CP(
        clk), .Q(\update_mask_0/reg_out[8][12] ) );
  dff_sg \update_mask_0/reg_out_reg[8][13]  ( .D(\update_mask_0/n1275 ), .CP(
        clk), .Q(\update_mask_0/reg_out[8][13] ) );
  dff_sg \update_mask_0/reg_out_reg[8][14]  ( .D(\update_mask_0/n1274 ), .CP(
        clk), .Q(\update_mask_0/reg_out[8][14] ) );
  dff_sg \update_mask_0/reg_out_reg[8][15]  ( .D(\update_mask_0/n1273 ), .CP(
        clk), .Q(\update_mask_0/reg_out[8][15] ) );
  dff_sg \update_mask_0/reg_out_reg[8][16]  ( .D(\update_mask_0/n1272 ), .CP(
        clk), .Q(\update_mask_0/reg_out[8][16] ) );
  dff_sg \update_mask_0/reg_out_reg[8][17]  ( .D(\update_mask_0/n1271 ), .CP(
        clk), .Q(\update_mask_0/reg_out[8][17] ) );
  dff_sg \update_mask_0/reg_out_reg[8][18]  ( .D(\update_mask_0/n1270 ), .CP(
        clk), .Q(\update_mask_0/reg_out[8][18] ) );
  dff_sg \update_mask_0/reg_out_reg[8][19]  ( .D(\update_mask_0/n1269 ), .CP(
        clk), .Q(\update_mask_0/reg_out[8][19] ) );
  dff_sg \update_mask_0/reg_out_reg[9][0]  ( .D(\update_mask_0/n1268 ), .CP(
        clk), .Q(\update_mask_0/reg_out[9][0] ) );
  dff_sg \update_mask_0/reg_out_reg[9][1]  ( .D(\update_mask_0/n1267 ), .CP(
        clk), .Q(\update_mask_0/reg_out[9][1] ) );
  dff_sg \update_mask_0/reg_out_reg[9][2]  ( .D(\update_mask_0/n1266 ), .CP(
        clk), .Q(\update_mask_0/reg_out[9][2] ) );
  dff_sg \update_mask_0/reg_out_reg[9][3]  ( .D(\update_mask_0/n1265 ), .CP(
        clk), .Q(\update_mask_0/reg_out[9][3] ) );
  dff_sg \update_mask_0/reg_out_reg[9][4]  ( .D(\update_mask_0/n1264 ), .CP(
        clk), .Q(\update_mask_0/reg_out[9][4] ) );
  dff_sg \update_mask_0/reg_out_reg[9][5]  ( .D(\update_mask_0/n1263 ), .CP(
        clk), .Q(\update_mask_0/reg_out[9][5] ) );
  dff_sg \update_mask_0/reg_out_reg[9][6]  ( .D(\update_mask_0/n1262 ), .CP(
        clk), .Q(\update_mask_0/reg_out[9][6] ) );
  dff_sg \update_mask_0/reg_out_reg[9][7]  ( .D(\update_mask_0/n1261 ), .CP(
        clk), .Q(\update_mask_0/reg_out[9][7] ) );
  dff_sg \update_mask_0/reg_out_reg[9][8]  ( .D(\update_mask_0/n1260 ), .CP(
        clk), .Q(\update_mask_0/reg_out[9][8] ) );
  dff_sg \update_mask_0/reg_out_reg[9][9]  ( .D(\update_mask_0/n1259 ), .CP(
        clk), .Q(\update_mask_0/reg_out[9][9] ) );
  dff_sg \update_mask_0/reg_out_reg[9][10]  ( .D(\update_mask_0/n1258 ), .CP(
        clk), .Q(\update_mask_0/reg_out[9][10] ) );
  dff_sg \update_mask_0/reg_out_reg[9][11]  ( .D(\update_mask_0/n1257 ), .CP(
        clk), .Q(\update_mask_0/reg_out[9][11] ) );
  dff_sg \update_mask_0/reg_out_reg[9][12]  ( .D(\update_mask_0/n1256 ), .CP(
        clk), .Q(\update_mask_0/reg_out[9][12] ) );
  dff_sg \update_mask_0/reg_out_reg[9][13]  ( .D(\update_mask_0/n1255 ), .CP(
        clk), .Q(\update_mask_0/reg_out[9][13] ) );
  dff_sg \update_mask_0/reg_out_reg[9][14]  ( .D(\update_mask_0/n1254 ), .CP(
        clk), .Q(\update_mask_0/reg_out[9][14] ) );
  dff_sg \update_mask_0/reg_out_reg[9][15]  ( .D(\update_mask_0/n1253 ), .CP(
        clk), .Q(\update_mask_0/reg_out[9][15] ) );
  dff_sg \update_mask_0/reg_out_reg[9][16]  ( .D(\update_mask_0/n1252 ), .CP(
        clk), .Q(\update_mask_0/reg_out[9][16] ) );
  dff_sg \update_mask_0/reg_out_reg[9][17]  ( .D(\update_mask_0/n1251 ), .CP(
        clk), .Q(\update_mask_0/reg_out[9][17] ) );
  dff_sg \update_mask_0/reg_out_reg[9][18]  ( .D(\update_mask_0/n1250 ), .CP(
        clk), .Q(\update_mask_0/reg_out[9][18] ) );
  dff_sg \update_mask_0/reg_out_reg[9][19]  ( .D(\update_mask_0/n1249 ), .CP(
        clk), .Q(\update_mask_0/reg_out[9][19] ) );
  dff_sg \update_mask_0/reg_out_reg[10][0]  ( .D(\update_mask_0/n1248 ), .CP(
        clk), .Q(\update_mask_0/reg_out[10][0] ) );
  dff_sg \update_mask_0/reg_out_reg[10][1]  ( .D(\update_mask_0/n1247 ), .CP(
        clk), .Q(\update_mask_0/reg_out[10][1] ) );
  dff_sg \update_mask_0/reg_out_reg[10][2]  ( .D(\update_mask_0/n1246 ), .CP(
        clk), .Q(\update_mask_0/reg_out[10][2] ) );
  dff_sg \update_mask_0/reg_out_reg[10][3]  ( .D(\update_mask_0/n1245 ), .CP(
        clk), .Q(\update_mask_0/reg_out[10][3] ) );
  dff_sg \update_mask_0/reg_out_reg[10][4]  ( .D(\update_mask_0/n1244 ), .CP(
        clk), .Q(\update_mask_0/reg_out[10][4] ) );
  dff_sg \update_mask_0/reg_out_reg[10][5]  ( .D(\update_mask_0/n1243 ), .CP(
        clk), .Q(\update_mask_0/reg_out[10][5] ) );
  dff_sg \update_mask_0/reg_out_reg[10][6]  ( .D(\update_mask_0/n1242 ), .CP(
        clk), .Q(\update_mask_0/reg_out[10][6] ) );
  dff_sg \update_mask_0/reg_out_reg[10][7]  ( .D(\update_mask_0/n1241 ), .CP(
        clk), .Q(\update_mask_0/reg_out[10][7] ) );
  dff_sg \update_mask_0/reg_out_reg[10][8]  ( .D(\update_mask_0/n1240 ), .CP(
        clk), .Q(\update_mask_0/reg_out[10][8] ) );
  dff_sg \update_mask_0/reg_out_reg[10][9]  ( .D(\update_mask_0/n1239 ), .CP(
        clk), .Q(\update_mask_0/reg_out[10][9] ) );
  dff_sg \update_mask_0/reg_out_reg[10][10]  ( .D(\update_mask_0/n1238 ), .CP(
        clk), .Q(\update_mask_0/reg_out[10][10] ) );
  dff_sg \update_mask_0/reg_out_reg[10][11]  ( .D(\update_mask_0/n1237 ), .CP(
        clk), .Q(\update_mask_0/reg_out[10][11] ) );
  dff_sg \update_mask_0/reg_out_reg[10][12]  ( .D(\update_mask_0/n1236 ), .CP(
        clk), .Q(\update_mask_0/reg_out[10][12] ) );
  dff_sg \update_mask_0/reg_out_reg[10][13]  ( .D(\update_mask_0/n1235 ), .CP(
        clk), .Q(\update_mask_0/reg_out[10][13] ) );
  dff_sg \update_mask_0/reg_out_reg[10][14]  ( .D(\update_mask_0/n1234 ), .CP(
        clk), .Q(\update_mask_0/reg_out[10][14] ) );
  dff_sg \update_mask_0/reg_out_reg[10][15]  ( .D(\update_mask_0/n1233 ), .CP(
        clk), .Q(\update_mask_0/reg_out[10][15] ) );
  dff_sg \update_mask_0/reg_out_reg[10][16]  ( .D(\update_mask_0/n1232 ), .CP(
        clk), .Q(\update_mask_0/reg_out[10][16] ) );
  dff_sg \update_mask_0/reg_out_reg[10][17]  ( .D(\update_mask_0/n1231 ), .CP(
        clk), .Q(\update_mask_0/reg_out[10][17] ) );
  dff_sg \update_mask_0/reg_out_reg[10][18]  ( .D(\update_mask_0/n1230 ), .CP(
        clk), .Q(\update_mask_0/reg_out[10][18] ) );
  dff_sg \update_mask_0/reg_out_reg[10][19]  ( .D(\update_mask_0/n1229 ), .CP(
        clk), .Q(\update_mask_0/reg_out[10][19] ) );
  dff_sg \update_mask_0/reg_out_reg[11][0]  ( .D(\update_mask_0/n1228 ), .CP(
        clk), .Q(\update_mask_0/reg_out[11][0] ) );
  dff_sg \update_mask_0/reg_out_reg[11][1]  ( .D(\update_mask_0/n1227 ), .CP(
        clk), .Q(\update_mask_0/reg_out[11][1] ) );
  dff_sg \update_mask_0/reg_out_reg[11][2]  ( .D(\update_mask_0/n1226 ), .CP(
        clk), .Q(\update_mask_0/reg_out[11][2] ) );
  dff_sg \update_mask_0/reg_out_reg[11][3]  ( .D(\update_mask_0/n1225 ), .CP(
        clk), .Q(\update_mask_0/reg_out[11][3] ) );
  dff_sg \update_mask_0/reg_out_reg[11][4]  ( .D(\update_mask_0/n1224 ), .CP(
        clk), .Q(\update_mask_0/reg_out[11][4] ) );
  dff_sg \update_mask_0/reg_out_reg[11][5]  ( .D(\update_mask_0/n1223 ), .CP(
        clk), .Q(\update_mask_0/reg_out[11][5] ) );
  dff_sg \update_mask_0/reg_out_reg[11][6]  ( .D(\update_mask_0/n1222 ), .CP(
        clk), .Q(\update_mask_0/reg_out[11][6] ) );
  dff_sg \update_mask_0/reg_out_reg[11][7]  ( .D(\update_mask_0/n1221 ), .CP(
        clk), .Q(\update_mask_0/reg_out[11][7] ) );
  dff_sg \update_mask_0/reg_out_reg[11][8]  ( .D(\update_mask_0/n1220 ), .CP(
        clk), .Q(\update_mask_0/reg_out[11][8] ) );
  dff_sg \update_mask_0/reg_out_reg[11][9]  ( .D(\update_mask_0/n1219 ), .CP(
        clk), .Q(\update_mask_0/reg_out[11][9] ) );
  dff_sg \update_mask_0/reg_out_reg[11][10]  ( .D(\update_mask_0/n1218 ), .CP(
        clk), .Q(\update_mask_0/reg_out[11][10] ) );
  dff_sg \update_mask_0/reg_out_reg[11][11]  ( .D(\update_mask_0/n1217 ), .CP(
        clk), .Q(\update_mask_0/reg_out[11][11] ) );
  dff_sg \update_mask_0/reg_out_reg[11][12]  ( .D(\update_mask_0/n1216 ), .CP(
        clk), .Q(\update_mask_0/reg_out[11][12] ) );
  dff_sg \update_mask_0/reg_out_reg[11][13]  ( .D(\update_mask_0/n1215 ), .CP(
        clk), .Q(\update_mask_0/reg_out[11][13] ) );
  dff_sg \update_mask_0/reg_out_reg[11][14]  ( .D(\update_mask_0/n1214 ), .CP(
        clk), .Q(\update_mask_0/reg_out[11][14] ) );
  dff_sg \update_mask_0/reg_out_reg[11][15]  ( .D(\update_mask_0/n1213 ), .CP(
        clk), .Q(\update_mask_0/reg_out[11][15] ) );
  dff_sg \update_mask_0/reg_out_reg[11][16]  ( .D(\update_mask_0/n1212 ), .CP(
        clk), .Q(\update_mask_0/reg_out[11][16] ) );
  dff_sg \update_mask_0/reg_out_reg[11][17]  ( .D(\update_mask_0/n1211 ), .CP(
        clk), .Q(\update_mask_0/reg_out[11][17] ) );
  dff_sg \update_mask_0/reg_out_reg[11][18]  ( .D(\update_mask_0/n1210 ), .CP(
        clk), .Q(\update_mask_0/reg_out[11][18] ) );
  dff_sg \update_mask_0/reg_out_reg[11][19]  ( .D(\update_mask_0/n1209 ), .CP(
        clk), .Q(\update_mask_0/reg_out[11][19] ) );
  dff_sg \update_mask_0/reg_out_reg[12][0]  ( .D(\update_mask_0/n1208 ), .CP(
        clk), .Q(\update_mask_0/reg_out[12][0] ) );
  dff_sg \update_mask_0/reg_out_reg[12][1]  ( .D(\update_mask_0/n1207 ), .CP(
        clk), .Q(\update_mask_0/reg_out[12][1] ) );
  dff_sg \update_mask_0/reg_out_reg[12][2]  ( .D(\update_mask_0/n1206 ), .CP(
        clk), .Q(\update_mask_0/reg_out[12][2] ) );
  dff_sg \update_mask_0/reg_out_reg[12][3]  ( .D(\update_mask_0/n1205 ), .CP(
        clk), .Q(\update_mask_0/reg_out[12][3] ) );
  dff_sg \update_mask_0/reg_out_reg[12][4]  ( .D(\update_mask_0/n1204 ), .CP(
        clk), .Q(\update_mask_0/reg_out[12][4] ) );
  dff_sg \update_mask_0/reg_out_reg[12][5]  ( .D(\update_mask_0/n1203 ), .CP(
        clk), .Q(\update_mask_0/reg_out[12][5] ) );
  dff_sg \update_mask_0/reg_out_reg[12][6]  ( .D(\update_mask_0/n1202 ), .CP(
        clk), .Q(\update_mask_0/reg_out[12][6] ) );
  dff_sg \update_mask_0/reg_out_reg[12][7]  ( .D(\update_mask_0/n1201 ), .CP(
        clk), .Q(\update_mask_0/reg_out[12][7] ) );
  dff_sg \update_mask_0/reg_out_reg[12][8]  ( .D(\update_mask_0/n1200 ), .CP(
        clk), .Q(\update_mask_0/reg_out[12][8] ) );
  dff_sg \update_mask_0/reg_out_reg[12][9]  ( .D(\update_mask_0/n1199 ), .CP(
        clk), .Q(\update_mask_0/reg_out[12][9] ) );
  dff_sg \update_mask_0/reg_out_reg[12][10]  ( .D(\update_mask_0/n1198 ), .CP(
        clk), .Q(\update_mask_0/reg_out[12][10] ) );
  dff_sg \update_mask_0/reg_out_reg[12][11]  ( .D(\update_mask_0/n1197 ), .CP(
        clk), .Q(\update_mask_0/reg_out[12][11] ) );
  dff_sg \update_mask_0/reg_out_reg[12][12]  ( .D(\update_mask_0/n1196 ), .CP(
        clk), .Q(\update_mask_0/reg_out[12][12] ) );
  dff_sg \update_mask_0/reg_out_reg[12][13]  ( .D(\update_mask_0/n1195 ), .CP(
        clk), .Q(\update_mask_0/reg_out[12][13] ) );
  dff_sg \update_mask_0/reg_out_reg[12][14]  ( .D(\update_mask_0/n1194 ), .CP(
        clk), .Q(\update_mask_0/reg_out[12][14] ) );
  dff_sg \update_mask_0/reg_out_reg[12][15]  ( .D(\update_mask_0/n1193 ), .CP(
        clk), .Q(\update_mask_0/reg_out[12][15] ) );
  dff_sg \update_mask_0/reg_out_reg[12][16]  ( .D(\update_mask_0/n1192 ), .CP(
        clk), .Q(\update_mask_0/reg_out[12][16] ) );
  dff_sg \update_mask_0/reg_out_reg[12][17]  ( .D(\update_mask_0/n1191 ), .CP(
        clk), .Q(\update_mask_0/reg_out[12][17] ) );
  dff_sg \update_mask_0/reg_out_reg[12][18]  ( .D(\update_mask_0/n1190 ), .CP(
        clk), .Q(\update_mask_0/reg_out[12][18] ) );
  dff_sg \update_mask_0/reg_out_reg[12][19]  ( .D(\update_mask_0/n1189 ), .CP(
        clk), .Q(\update_mask_0/reg_out[12][19] ) );
  dff_sg \update_mask_0/reg_out_reg[13][0]  ( .D(\update_mask_0/n1188 ), .CP(
        clk), .Q(\update_mask_0/reg_out[13][0] ) );
  dff_sg \update_mask_0/reg_out_reg[13][1]  ( .D(\update_mask_0/n1187 ), .CP(
        clk), .Q(\update_mask_0/reg_out[13][1] ) );
  dff_sg \update_mask_0/reg_out_reg[13][2]  ( .D(\update_mask_0/n1186 ), .CP(
        clk), .Q(\update_mask_0/reg_out[13][2] ) );
  dff_sg \update_mask_0/reg_out_reg[13][3]  ( .D(\update_mask_0/n1185 ), .CP(
        clk), .Q(\update_mask_0/reg_out[13][3] ) );
  dff_sg \update_mask_0/reg_out_reg[13][4]  ( .D(\update_mask_0/n1184 ), .CP(
        clk), .Q(\update_mask_0/reg_out[13][4] ) );
  dff_sg \update_mask_0/reg_out_reg[13][5]  ( .D(\update_mask_0/n1183 ), .CP(
        clk), .Q(\update_mask_0/reg_out[13][5] ) );
  dff_sg \update_mask_0/reg_out_reg[13][6]  ( .D(\update_mask_0/n1182 ), .CP(
        clk), .Q(\update_mask_0/reg_out[13][6] ) );
  dff_sg \update_mask_0/reg_out_reg[13][7]  ( .D(\update_mask_0/n1181 ), .CP(
        clk), .Q(\update_mask_0/reg_out[13][7] ) );
  dff_sg \update_mask_0/reg_out_reg[13][8]  ( .D(\update_mask_0/n1180 ), .CP(
        clk), .Q(\update_mask_0/reg_out[13][8] ) );
  dff_sg \update_mask_0/reg_out_reg[13][9]  ( .D(\update_mask_0/n1179 ), .CP(
        clk), .Q(\update_mask_0/reg_out[13][9] ) );
  dff_sg \update_mask_0/reg_out_reg[13][10]  ( .D(\update_mask_0/n1178 ), .CP(
        clk), .Q(\update_mask_0/reg_out[13][10] ) );
  dff_sg \update_mask_0/reg_out_reg[13][11]  ( .D(\update_mask_0/n1177 ), .CP(
        clk), .Q(\update_mask_0/reg_out[13][11] ) );
  dff_sg \update_mask_0/reg_out_reg[13][12]  ( .D(\update_mask_0/n1176 ), .CP(
        clk), .Q(\update_mask_0/reg_out[13][12] ) );
  dff_sg \update_mask_0/reg_out_reg[13][13]  ( .D(\update_mask_0/n1175 ), .CP(
        clk), .Q(\update_mask_0/reg_out[13][13] ) );
  dff_sg \update_mask_0/reg_out_reg[13][14]  ( .D(\update_mask_0/n1174 ), .CP(
        clk), .Q(\update_mask_0/reg_out[13][14] ) );
  dff_sg \update_mask_0/reg_out_reg[13][15]  ( .D(\update_mask_0/n1173 ), .CP(
        clk), .Q(\update_mask_0/reg_out[13][15] ) );
  dff_sg \update_mask_0/reg_out_reg[13][16]  ( .D(\update_mask_0/n1172 ), .CP(
        clk), .Q(\update_mask_0/reg_out[13][16] ) );
  dff_sg \update_mask_0/reg_out_reg[13][17]  ( .D(\update_mask_0/n1171 ), .CP(
        clk), .Q(\update_mask_0/reg_out[13][17] ) );
  dff_sg \update_mask_0/reg_out_reg[13][18]  ( .D(\update_mask_0/n1170 ), .CP(
        clk), .Q(\update_mask_0/reg_out[13][18] ) );
  dff_sg \update_mask_0/reg_out_reg[13][19]  ( .D(\update_mask_0/n1169 ), .CP(
        clk), .Q(\update_mask_0/reg_out[13][19] ) );
  dff_sg \update_mask_0/reg_out_reg[14][0]  ( .D(\update_mask_0/n1168 ), .CP(
        clk), .Q(\update_mask_0/reg_out[14][0] ) );
  dff_sg \update_mask_0/reg_out_reg[14][1]  ( .D(\update_mask_0/n1167 ), .CP(
        clk), .Q(\update_mask_0/reg_out[14][1] ) );
  dff_sg \update_mask_0/reg_out_reg[14][2]  ( .D(\update_mask_0/n1166 ), .CP(
        clk), .Q(\update_mask_0/reg_out[14][2] ) );
  dff_sg \update_mask_0/reg_out_reg[14][3]  ( .D(\update_mask_0/n1165 ), .CP(
        clk), .Q(\update_mask_0/reg_out[14][3] ) );
  dff_sg \update_mask_0/reg_out_reg[14][4]  ( .D(\update_mask_0/n1164 ), .CP(
        clk), .Q(\update_mask_0/reg_out[14][4] ) );
  dff_sg \update_mask_0/reg_out_reg[14][5]  ( .D(\update_mask_0/n1163 ), .CP(
        clk), .Q(\update_mask_0/reg_out[14][5] ) );
  dff_sg \update_mask_0/reg_out_reg[14][6]  ( .D(\update_mask_0/n1162 ), .CP(
        clk), .Q(\update_mask_0/reg_out[14][6] ) );
  dff_sg \update_mask_0/reg_out_reg[14][7]  ( .D(\update_mask_0/n1161 ), .CP(
        clk), .Q(\update_mask_0/reg_out[14][7] ) );
  dff_sg \update_mask_0/reg_out_reg[14][8]  ( .D(\update_mask_0/n1160 ), .CP(
        clk), .Q(\update_mask_0/reg_out[14][8] ) );
  dff_sg \update_mask_0/reg_out_reg[14][9]  ( .D(\update_mask_0/n1159 ), .CP(
        clk), .Q(\update_mask_0/reg_out[14][9] ) );
  dff_sg \update_mask_0/reg_out_reg[14][10]  ( .D(\update_mask_0/n1158 ), .CP(
        clk), .Q(\update_mask_0/reg_out[14][10] ) );
  dff_sg \update_mask_0/reg_out_reg[14][11]  ( .D(\update_mask_0/n1157 ), .CP(
        clk), .Q(\update_mask_0/reg_out[14][11] ) );
  dff_sg \update_mask_0/reg_out_reg[14][12]  ( .D(\update_mask_0/n1156 ), .CP(
        clk), .Q(\update_mask_0/reg_out[14][12] ) );
  dff_sg \update_mask_0/reg_out_reg[14][13]  ( .D(\update_mask_0/n1155 ), .CP(
        clk), .Q(\update_mask_0/reg_out[14][13] ) );
  dff_sg \update_mask_0/reg_out_reg[14][14]  ( .D(\update_mask_0/n1154 ), .CP(
        clk), .Q(\update_mask_0/reg_out[14][14] ) );
  dff_sg \update_mask_0/reg_out_reg[14][15]  ( .D(\update_mask_0/n1153 ), .CP(
        clk), .Q(\update_mask_0/reg_out[14][15] ) );
  dff_sg \update_mask_0/reg_out_reg[14][16]  ( .D(\update_mask_0/n1152 ), .CP(
        clk), .Q(\update_mask_0/reg_out[14][16] ) );
  dff_sg \update_mask_0/reg_out_reg[14][17]  ( .D(\update_mask_0/n1151 ), .CP(
        clk), .Q(\update_mask_0/reg_out[14][17] ) );
  dff_sg \update_mask_0/reg_out_reg[14][18]  ( .D(\update_mask_0/n1150 ), .CP(
        clk), .Q(\update_mask_0/reg_out[14][18] ) );
  dff_sg \update_mask_0/reg_out_reg[14][19]  ( .D(\update_mask_0/n1149 ), .CP(
        clk), .Q(\update_mask_0/reg_out[14][19] ) );
  dff_sg \update_mask_0/reg_out_reg[15][0]  ( .D(\update_mask_0/n1148 ), .CP(
        clk), .Q(\update_mask_0/reg_out[15][0] ) );
  dff_sg \update_mask_0/reg_out_reg[15][1]  ( .D(\update_mask_0/n1147 ), .CP(
        clk), .Q(\update_mask_0/reg_out[15][1] ) );
  dff_sg \update_mask_0/reg_out_reg[15][2]  ( .D(\update_mask_0/n1146 ), .CP(
        clk), .Q(\update_mask_0/reg_out[15][2] ) );
  dff_sg \update_mask_0/reg_out_reg[15][3]  ( .D(\update_mask_0/n1145 ), .CP(
        clk), .Q(\update_mask_0/reg_out[15][3] ) );
  dff_sg \update_mask_0/reg_out_reg[15][4]  ( .D(\update_mask_0/n1144 ), .CP(
        clk), .Q(\update_mask_0/reg_out[15][4] ) );
  dff_sg \update_mask_0/reg_out_reg[15][5]  ( .D(\update_mask_0/n1143 ), .CP(
        clk), .Q(\update_mask_0/reg_out[15][5] ) );
  dff_sg \update_mask_0/reg_out_reg[15][6]  ( .D(\update_mask_0/n1142 ), .CP(
        clk), .Q(\update_mask_0/reg_out[15][6] ) );
  dff_sg \update_mask_0/reg_out_reg[15][7]  ( .D(\update_mask_0/n1141 ), .CP(
        clk), .Q(\update_mask_0/reg_out[15][7] ) );
  dff_sg \update_mask_0/reg_out_reg[15][8]  ( .D(\update_mask_0/n1140 ), .CP(
        clk), .Q(\update_mask_0/reg_out[15][8] ) );
  dff_sg \update_mask_0/reg_out_reg[15][9]  ( .D(\update_mask_0/n1139 ), .CP(
        clk), .Q(\update_mask_0/reg_out[15][9] ) );
  dff_sg \update_mask_0/reg_out_reg[15][10]  ( .D(\update_mask_0/n1138 ), .CP(
        clk), .Q(\update_mask_0/reg_out[15][10] ) );
  dff_sg \update_mask_0/reg_out_reg[15][11]  ( .D(\update_mask_0/n1137 ), .CP(
        clk), .Q(\update_mask_0/reg_out[15][11] ) );
  dff_sg \update_mask_0/reg_out_reg[15][12]  ( .D(\update_mask_0/n1136 ), .CP(
        clk), .Q(\update_mask_0/reg_out[15][12] ) );
  dff_sg \update_mask_0/reg_out_reg[15][13]  ( .D(\update_mask_0/n1135 ), .CP(
        clk), .Q(\update_mask_0/reg_out[15][13] ) );
  dff_sg \update_mask_0/reg_out_reg[15][14]  ( .D(\update_mask_0/n1134 ), .CP(
        clk), .Q(\update_mask_0/reg_out[15][14] ) );
  dff_sg \update_mask_0/reg_out_reg[15][15]  ( .D(\update_mask_0/n1133 ), .CP(
        clk), .Q(\update_mask_0/reg_out[15][15] ) );
  dff_sg \update_mask_0/reg_out_reg[15][16]  ( .D(\update_mask_0/n1132 ), .CP(
        clk), .Q(\update_mask_0/reg_out[15][16] ) );
  dff_sg \update_mask_0/reg_out_reg[15][17]  ( .D(\update_mask_0/n1131 ), .CP(
        clk), .Q(\update_mask_0/reg_out[15][17] ) );
  dff_sg \update_mask_0/reg_out_reg[15][18]  ( .D(\update_mask_0/n1130 ), .CP(
        clk), .Q(\update_mask_0/reg_out[15][18] ) );
  dff_sg \update_mask_0/reg_out_reg[15][19]  ( .D(\update_mask_0/n1129 ), .CP(
        clk), .Q(\update_mask_0/reg_out[15][19] ) );
  dff_sg \update_mask_0/state_reg[0]  ( .D(\update_mask_0/n1127 ), .CP(clk), 
        .Q(\update_mask_0/n4206 ) );
  dff_sg \update_mask_0/state_reg[1]  ( .D(n5885), .CP(clk), .Q(
        \update_mask_0/n4205 ) );
  dff_sg \update_mask_0/m_pointer_reg[4]  ( .D(n5877), .CP(clk), .Q(
        \update_mask_0/N27 ) );
  dff_sg \update_mask_0/m_pointer_reg[0]  ( .D(n5881), .CP(clk), .Q(
        \update_mask_0/N23 ) );
  dff_sg \update_output_0/o_im_reg[13][19]  ( .D(n5852), .CP(clk), .Q(n9288)
         );
  dff_sg \update_output_0/o_im_reg[13][18]  ( .D(n5833), .CP(clk), .Q(n9289)
         );
  dff_sg \update_output_0/o_im_reg[13][17]  ( .D(n5829), .CP(clk), .Q(n9290)
         );
  dff_sg \update_output_0/o_im_reg[13][16]  ( .D(n5840), .CP(clk), .Q(n9291)
         );
  dff_sg \update_output_0/o_im_reg[13][15]  ( .D(n5837), .CP(clk), .Q(n9292)
         );
  dff_sg \update_output_0/o_im_reg[13][14]  ( .D(n5870), .CP(clk), .Q(n9293)
         );
  dff_sg \update_output_0/o_im_reg[13][13]  ( .D(n5872), .CP(clk), .Q(n9294)
         );
  dff_sg \update_output_0/o_im_reg[13][12]  ( .D(n5875), .CP(clk), .Q(n9295)
         );
  dff_sg \update_output_0/o_im_reg[13][11]  ( .D(n5873), .CP(clk), .Q(n9296)
         );
  dff_sg \update_output_0/o_im_reg[13][10]  ( .D(n5848), .CP(clk), .Q(n9297)
         );
  dff_sg \update_output_0/o_im_reg[13][9]  ( .D(n5845), .CP(clk), .Q(n9298) );
  dff_sg \update_output_0/o_im_reg[13][8]  ( .D(n5812), .CP(clk), .Q(n9299) );
  dff_sg \update_output_0/o_im_reg[13][7]  ( .D(n5815), .CP(clk), .Q(n9300) );
  dff_sg \update_output_0/o_im_reg[13][6]  ( .D(n5825), .CP(clk), .Q(n9301) );
  dff_sg \update_output_0/o_im_reg[13][5]  ( .D(n5819), .CP(clk), .Q(n9302) );
  dff_sg \update_output_0/o_im_reg[13][4]  ( .D(n5799), .CP(clk), .Q(n9303) );
  dff_sg \update_output_0/o_im_reg[13][3]  ( .D(n5797), .CP(clk), .Q(n9304) );
  dff_sg \update_output_0/o_im_reg[13][2]  ( .D(n5803), .CP(clk), .Q(n9305) );
  dff_sg \update_output_0/o_im_reg[13][1]  ( .D(n5807), .CP(clk), .Q(n9306) );
  dff_sg \update_output_0/o_im_reg[13][0]  ( .D(n5876), .CP(clk), .Q(n9307) );
  dff_sg \update_output_0/o_im_reg[5][19]  ( .D(n5643), .CP(clk), .Q(n9448) );
  dff_sg \update_output_0/o_im_reg[5][18]  ( .D(n5634), .CP(clk), .Q(n9449) );
  dff_sg \update_output_0/o_im_reg[5][17]  ( .D(n5642), .CP(clk), .Q(n9450) );
  dff_sg \update_output_0/o_im_reg[5][16]  ( .D(n5633), .CP(clk), .Q(n9451) );
  dff_sg \update_output_0/o_im_reg[5][15]  ( .D(n5645), .CP(clk), .Q(n9452) );
  dff_sg \update_output_0/o_im_reg[5][14]  ( .D(n5635), .CP(clk), .Q(n9453) );
  dff_sg \update_output_0/o_im_reg[5][13]  ( .D(n5632), .CP(clk), .Q(n9454) );
  dff_sg \update_output_0/o_im_reg[5][12]  ( .D(n5874), .CP(clk), .Q(n9455) );
  dff_sg \update_output_0/o_im_reg[5][11]  ( .D(n5641), .CP(clk), .Q(n9456) );
  dff_sg \update_output_0/o_im_reg[5][10]  ( .D(n5631), .CP(clk), .Q(n9457) );
  dff_sg \update_output_0/o_im_reg[5][9]  ( .D(n5637), .CP(clk), .Q(n9458) );
  dff_sg \update_output_0/o_im_reg[5][8]  ( .D(n5640), .CP(clk), .Q(n9459) );
  dff_sg \update_output_0/o_im_reg[5][7]  ( .D(n5630), .CP(clk), .Q(n9460) );
  dff_sg \update_output_0/o_im_reg[5][6]  ( .D(n5644), .CP(clk), .Q(n9461) );
  dff_sg \update_output_0/o_im_reg[5][5]  ( .D(n5639), .CP(clk), .Q(n9462) );
  dff_sg \update_output_0/o_im_reg[5][4]  ( .D(n5629), .CP(clk), .Q(n9463) );
  dff_sg \update_output_0/o_im_reg[5][3]  ( .D(n5636), .CP(clk), .Q(n9464) );
  dff_sg \update_output_0/o_im_reg[5][2]  ( .D(n5638), .CP(clk), .Q(n9465) );
  dff_sg \update_output_0/o_im_reg[5][1]  ( .D(n5628), .CP(clk), .Q(n9466) );
  dff_sg \update_output_0/o_im_reg[5][0]  ( .D(n5646), .CP(clk), .Q(n9467) );
  dff_sg \update_output_0/o_im_reg[14][19]  ( .D(n5585), .CP(clk), .Q(n9268)
         );
  dff_sg \update_output_0/o_im_reg[14][18]  ( .D(n5568), .CP(clk), .Q(n9269)
         );
  dff_sg \update_output_0/o_im_reg[14][17]  ( .D(n5576), .CP(clk), .Q(n9270)
         );
  dff_sg \update_output_0/o_im_reg[14][16]  ( .D(n5580), .CP(clk), .Q(n9271)
         );
  dff_sg \update_output_0/o_im_reg[14][15]  ( .D(n5573), .CP(clk), .Q(n9272)
         );
  dff_sg \update_output_0/o_im_reg[14][14]  ( .D(n5575), .CP(clk), .Q(n9273)
         );
  dff_sg \update_output_0/o_im_reg[14][13]  ( .D(n5574), .CP(clk), .Q(n9274)
         );
  dff_sg \update_output_0/o_im_reg[14][12]  ( .D(n5577), .CP(clk), .Q(n9275)
         );
  dff_sg \update_output_0/o_im_reg[14][11]  ( .D(n5582), .CP(clk), .Q(n9276)
         );
  dff_sg \update_output_0/o_im_reg[14][10]  ( .D(n5570), .CP(clk), .Q(n9277)
         );
  dff_sg \update_output_0/o_im_reg[14][9]  ( .D(n5584), .CP(clk), .Q(n9278) );
  dff_sg \update_output_0/o_im_reg[14][8]  ( .D(n5571), .CP(clk), .Q(n9279) );
  dff_sg \update_output_0/o_im_reg[14][7]  ( .D(n5578), .CP(clk), .Q(n9280) );
  dff_sg \update_output_0/o_im_reg[14][6]  ( .D(n5581), .CP(clk), .Q(n9281) );
  dff_sg \update_output_0/o_im_reg[14][5]  ( .D(n5572), .CP(clk), .Q(n9282) );
  dff_sg \update_output_0/o_im_reg[14][4]  ( .D(n5586), .CP(clk), .Q(n9283) );
  dff_sg \update_output_0/o_im_reg[14][3]  ( .D(n5569), .CP(clk), .Q(n9284) );
  dff_sg \update_output_0/o_im_reg[14][2]  ( .D(n5583), .CP(clk), .Q(n9285) );
  dff_sg \update_output_0/o_im_reg[14][1]  ( .D(n5579), .CP(clk), .Q(n9286) );
  dff_sg \update_output_0/o_im_reg[14][0]  ( .D(n5587), .CP(clk), .Q(n9287) );
  dff_sg \update_output_0/o_im_reg[6][19]  ( .D(n5565), .CP(clk), .Q(n9428) );
  dff_sg \update_output_0/o_im_reg[6][18]  ( .D(n5548), .CP(clk), .Q(n9429) );
  dff_sg \update_output_0/o_im_reg[6][17]  ( .D(n5561), .CP(clk), .Q(n9430) );
  dff_sg \update_output_0/o_im_reg[6][16]  ( .D(n5552), .CP(clk), .Q(n9431) );
  dff_sg \update_output_0/o_im_reg[6][15]  ( .D(n5557), .CP(clk), .Q(n9432) );
  dff_sg \update_output_0/o_im_reg[6][14]  ( .D(n5554), .CP(clk), .Q(n9433) );
  dff_sg \update_output_0/o_im_reg[6][13]  ( .D(n5558), .CP(clk), .Q(n9434) );
  dff_sg \update_output_0/o_im_reg[6][12]  ( .D(n5562), .CP(clk), .Q(n9435) );
  dff_sg \update_output_0/o_im_reg[6][11]  ( .D(n5555), .CP(clk), .Q(n9436) );
  dff_sg \update_output_0/o_im_reg[6][10]  ( .D(n5550), .CP(clk), .Q(n9437) );
  dff_sg \update_output_0/o_im_reg[6][9]  ( .D(n5564), .CP(clk), .Q(n9438) );
  dff_sg \update_output_0/o_im_reg[6][8]  ( .D(n5559), .CP(clk), .Q(n9439) );
  dff_sg \update_output_0/o_im_reg[6][7]  ( .D(n5563), .CP(clk), .Q(n9440) );
  dff_sg \update_output_0/o_im_reg[6][6]  ( .D(n5553), .CP(clk), .Q(n9441) );
  dff_sg \update_output_0/o_im_reg[6][5]  ( .D(n5556), .CP(clk), .Q(n9442) );
  dff_sg \update_output_0/o_im_reg[6][4]  ( .D(n5566), .CP(clk), .Q(n9443) );
  dff_sg \update_output_0/o_im_reg[6][3]  ( .D(n5549), .CP(clk), .Q(n9444) );
  dff_sg \update_output_0/o_im_reg[6][2]  ( .D(n5567), .CP(clk), .Q(n9445) );
  dff_sg \update_output_0/o_im_reg[6][1]  ( .D(n5551), .CP(clk), .Q(n9446) );
  dff_sg \update_output_0/o_im_reg[6][0]  ( .D(n5560), .CP(clk), .Q(n9447) );
  dff_sg \update_output_0/o_im_reg[4][19]  ( .D(n5698), .CP(clk), .Q(n9468) );
  dff_sg \update_output_0/o_im_reg[4][18]  ( .D(n5703), .CP(clk), .Q(n9469) );
  dff_sg \update_output_0/o_im_reg[4][17]  ( .D(n5693), .CP(clk), .Q(n9470) );
  dff_sg \update_output_0/o_im_reg[4][16]  ( .D(n5686), .CP(clk), .Q(n9471) );
  dff_sg \update_output_0/o_im_reg[4][15]  ( .D(n5697), .CP(clk), .Q(n9472) );
  dff_sg \update_output_0/o_im_reg[4][14]  ( .D(n5704), .CP(clk), .Q(n9473) );
  dff_sg \update_output_0/o_im_reg[4][13]  ( .D(n5696), .CP(clk), .Q(n9474) );
  dff_sg \update_output_0/o_im_reg[4][12]  ( .D(n5691), .CP(clk), .Q(n9475) );
  dff_sg \update_output_0/o_im_reg[4][11]  ( .D(n5702), .CP(clk), .Q(n9476) );
  dff_sg \update_output_0/o_im_reg[4][10]  ( .D(n5690), .CP(clk), .Q(n9477) );
  dff_sg \update_output_0/o_im_reg[4][9]  ( .D(n5699), .CP(clk), .Q(n9478) );
  dff_sg \update_output_0/o_im_reg[4][8]  ( .D(n5701), .CP(clk), .Q(n9479) );
  dff_sg \update_output_0/o_im_reg[4][7]  ( .D(n5700), .CP(clk), .Q(n9480) );
  dff_sg \update_output_0/o_im_reg[4][6]  ( .D(n5695), .CP(clk), .Q(n9481) );
  dff_sg \update_output_0/o_im_reg[4][5]  ( .D(n5685), .CP(clk), .Q(n9482) );
  dff_sg \update_output_0/o_im_reg[4][4]  ( .D(n5687), .CP(clk), .Q(n9483) );
  dff_sg \update_output_0/o_im_reg[4][3]  ( .D(n5694), .CP(clk), .Q(n9484) );
  dff_sg \update_output_0/o_im_reg[4][2]  ( .D(n5689), .CP(clk), .Q(n9485) );
  dff_sg \update_output_0/o_im_reg[4][1]  ( .D(n5692), .CP(clk), .Q(n9486) );
  dff_sg \update_output_0/o_im_reg[4][0]  ( .D(n5688), .CP(clk), .Q(n9487) );
  dff_sg \update_output_0/o_im_reg[12][19]  ( .D(n5766), .CP(clk), .Q(n9308)
         );
  dff_sg \update_output_0/o_im_reg[12][18]  ( .D(n5771), .CP(clk), .Q(n9309)
         );
  dff_sg \update_output_0/o_im_reg[12][17]  ( .D(n5761), .CP(clk), .Q(n9310)
         );
  dff_sg \update_output_0/o_im_reg[12][16]  ( .D(n5754), .CP(clk), .Q(n9311)
         );
  dff_sg \update_output_0/o_im_reg[12][15]  ( .D(n5765), .CP(clk), .Q(n9312)
         );
  dff_sg \update_output_0/o_im_reg[12][14]  ( .D(n5772), .CP(clk), .Q(n9313)
         );
  dff_sg \update_output_0/o_im_reg[12][13]  ( .D(n5764), .CP(clk), .Q(n9314)
         );
  dff_sg \update_output_0/o_im_reg[12][12]  ( .D(n5759), .CP(clk), .Q(n9315)
         );
  dff_sg \update_output_0/o_im_reg[12][11]  ( .D(n5770), .CP(clk), .Q(n9316)
         );
  dff_sg \update_output_0/o_im_reg[12][10]  ( .D(n5758), .CP(clk), .Q(n9317)
         );
  dff_sg \update_output_0/o_im_reg[12][9]  ( .D(n5767), .CP(clk), .Q(n9318) );
  dff_sg \update_output_0/o_im_reg[12][8]  ( .D(n5769), .CP(clk), .Q(n9319) );
  dff_sg \update_output_0/o_im_reg[12][7]  ( .D(n5768), .CP(clk), .Q(n9320) );
  dff_sg \update_output_0/o_im_reg[12][6]  ( .D(n5763), .CP(clk), .Q(n9321) );
  dff_sg \update_output_0/o_im_reg[12][5]  ( .D(n5753), .CP(clk), .Q(n9322) );
  dff_sg \update_output_0/o_im_reg[12][4]  ( .D(n5755), .CP(clk), .Q(n9323) );
  dff_sg \update_output_0/o_im_reg[12][3]  ( .D(n5762), .CP(clk), .Q(n9324) );
  dff_sg \update_output_0/o_im_reg[12][2]  ( .D(n5757), .CP(clk), .Q(n9325) );
  dff_sg \update_output_0/o_im_reg[12][1]  ( .D(n5760), .CP(clk), .Q(n9326) );
  dff_sg \update_output_0/o_im_reg[12][0]  ( .D(n5756), .CP(clk), .Q(n9327) );
  dff_sg \update_output_0/o_im_reg[3][19]  ( .D(n5625), .CP(clk), .Q(n9488) );
  dff_sg \update_output_0/o_im_reg[3][18]  ( .D(n5620), .CP(clk), .Q(n9489) );
  dff_sg \update_output_0/o_im_reg[3][17]  ( .D(n5623), .CP(clk), .Q(n9490) );
  dff_sg \update_output_0/o_im_reg[3][16]  ( .D(n5619), .CP(clk), .Q(n9491) );
  dff_sg \update_output_0/o_im_reg[3][15]  ( .D(n5610), .CP(clk), .Q(n9492) );
  dff_sg \update_output_0/o_im_reg[3][14]  ( .D(n5612), .CP(clk), .Q(n9493) );
  dff_sg \update_output_0/o_im_reg[3][13]  ( .D(n5617), .CP(clk), .Q(n9494) );
  dff_sg \update_output_0/o_im_reg[3][12]  ( .D(n5609), .CP(clk), .Q(n9495) );
  dff_sg \update_output_0/o_im_reg[3][11]  ( .D(n5613), .CP(clk), .Q(n9496) );
  dff_sg \update_output_0/o_im_reg[3][10]  ( .D(n5616), .CP(clk), .Q(n9497) );
  dff_sg \update_output_0/o_im_reg[3][9]  ( .D(n5626), .CP(clk), .Q(n9498) );
  dff_sg \update_output_0/o_im_reg[3][8]  ( .D(n5621), .CP(clk), .Q(n9499) );
  dff_sg \update_output_0/o_im_reg[3][7]  ( .D(n5624), .CP(clk), .Q(n9500) );
  dff_sg \update_output_0/o_im_reg[3][6]  ( .D(n5611), .CP(clk), .Q(n9501) );
  dff_sg \update_output_0/o_im_reg[3][5]  ( .D(n5615), .CP(clk), .Q(n9502) );
  dff_sg \update_output_0/o_im_reg[3][4]  ( .D(n5608), .CP(clk), .Q(n9503) );
  dff_sg \update_output_0/o_im_reg[3][3]  ( .D(n5614), .CP(clk), .Q(n9504) );
  dff_sg \update_output_0/o_im_reg[3][2]  ( .D(n5627), .CP(clk), .Q(n9505) );
  dff_sg \update_output_0/o_im_reg[3][1]  ( .D(n5618), .CP(clk), .Q(n9506) );
  dff_sg \update_output_0/o_im_reg[3][0]  ( .D(n5622), .CP(clk), .Q(n9507) );
  dff_sg \update_output_0/o_im_reg[11][19]  ( .D(n5605), .CP(clk), .Q(n9328)
         );
  dff_sg \update_output_0/o_im_reg[11][18]  ( .D(n5594), .CP(clk), .Q(n9329)
         );
  dff_sg \update_output_0/o_im_reg[11][17]  ( .D(n5599), .CP(clk), .Q(n9330)
         );
  dff_sg \update_output_0/o_im_reg[11][16]  ( .D(n5593), .CP(clk), .Q(n9331)
         );
  dff_sg \update_output_0/o_im_reg[11][15]  ( .D(n5590), .CP(clk), .Q(n9332)
         );
  dff_sg \update_output_0/o_im_reg[11][14]  ( .D(n5607), .CP(clk), .Q(n9333)
         );
  dff_sg \update_output_0/o_im_reg[11][13]  ( .D(n5595), .CP(clk), .Q(n9334)
         );
  dff_sg \update_output_0/o_im_reg[11][12]  ( .D(n5600), .CP(clk), .Q(n9335)
         );
  dff_sg \update_output_0/o_im_reg[11][11]  ( .D(n5596), .CP(clk), .Q(n9336)
         );
  dff_sg \update_output_0/o_im_reg[11][10]  ( .D(n5597), .CP(clk), .Q(n9337)
         );
  dff_sg \update_output_0/o_im_reg[11][9]  ( .D(n5604), .CP(clk), .Q(n9338) );
  dff_sg \update_output_0/o_im_reg[11][8]  ( .D(n5603), .CP(clk), .Q(n9339) );
  dff_sg \update_output_0/o_im_reg[11][7]  ( .D(n5601), .CP(clk), .Q(n9340) );
  dff_sg \update_output_0/o_im_reg[11][6]  ( .D(n5588), .CP(clk), .Q(n9341) );
  dff_sg \update_output_0/o_im_reg[11][5]  ( .D(n5598), .CP(clk), .Q(n9342) );
  dff_sg \update_output_0/o_im_reg[11][4]  ( .D(n5606), .CP(clk), .Q(n9343) );
  dff_sg \update_output_0/o_im_reg[11][3]  ( .D(n5602), .CP(clk), .Q(n9344) );
  dff_sg \update_output_0/o_im_reg[11][2]  ( .D(n5589), .CP(clk), .Q(n9345) );
  dff_sg \update_output_0/o_im_reg[11][1]  ( .D(n5592), .CP(clk), .Q(n9346) );
  dff_sg \update_output_0/o_im_reg[11][0]  ( .D(n5591), .CP(clk), .Q(n9347) );
  dff_sg \update_output_0/o_im_reg[9][19]  ( .D(n5666), .CP(clk), .Q(n9368) );
  dff_sg \update_output_0/o_im_reg[9][18]  ( .D(n5665), .CP(clk), .Q(n9369) );
  dff_sg \update_output_0/o_im_reg[9][17]  ( .D(n5651), .CP(clk), .Q(n9370) );
  dff_sg \update_output_0/o_im_reg[9][16]  ( .D(n5649), .CP(clk), .Q(n9371) );
  dff_sg \update_output_0/o_im_reg[9][15]  ( .D(n5664), .CP(clk), .Q(n9372) );
  dff_sg \update_output_0/o_im_reg[9][14]  ( .D(n5658), .CP(clk), .Q(n9373) );
  dff_sg \update_output_0/o_im_reg[9][13]  ( .D(n5663), .CP(clk), .Q(n9374) );
  dff_sg \update_output_0/o_im_reg[9][12]  ( .D(n5662), .CP(clk), .Q(n9375) );
  dff_sg \update_output_0/o_im_reg[9][11]  ( .D(n5661), .CP(clk), .Q(n9376) );
  dff_sg \update_output_0/o_im_reg[9][10]  ( .D(n5657), .CP(clk), .Q(n9377) );
  dff_sg \update_output_0/o_im_reg[9][9]  ( .D(n5652), .CP(clk), .Q(n9378) );
  dff_sg \update_output_0/o_im_reg[9][8]  ( .D(n5654), .CP(clk), .Q(n9379) );
  dff_sg \update_output_0/o_im_reg[9][7]  ( .D(n5660), .CP(clk), .Q(n9380) );
  dff_sg \update_output_0/o_im_reg[9][6]  ( .D(n5659), .CP(clk), .Q(n9381) );
  dff_sg \update_output_0/o_im_reg[9][5]  ( .D(n5647), .CP(clk), .Q(n9382) );
  dff_sg \update_output_0/o_im_reg[9][4]  ( .D(n5656), .CP(clk), .Q(n9383) );
  dff_sg \update_output_0/o_im_reg[9][3]  ( .D(n5655), .CP(clk), .Q(n9384) );
  dff_sg \update_output_0/o_im_reg[9][2]  ( .D(n5650), .CP(clk), .Q(n9385) );
  dff_sg \update_output_0/o_im_reg[9][1]  ( .D(n5648), .CP(clk), .Q(n9386) );
  dff_sg \update_output_0/o_im_reg[9][0]  ( .D(n5653), .CP(clk), .Q(n9387) );
  dff_sg \update_output_0/o_im_reg[1][19]  ( .D(n5683), .CP(clk), .Q(n9528) );
  dff_sg \update_output_0/o_im_reg[1][18]  ( .D(n5673), .CP(clk), .Q(n9529) );
  dff_sg \update_output_0/o_im_reg[1][17]  ( .D(n5678), .CP(clk), .Q(n9530) );
  dff_sg \update_output_0/o_im_reg[1][16]  ( .D(n5671), .CP(clk), .Q(n9531) );
  dff_sg \update_output_0/o_im_reg[1][15]  ( .D(n5675), .CP(clk), .Q(n9532) );
  dff_sg \update_output_0/o_im_reg[1][14]  ( .D(n5871), .CP(clk), .Q(n9533) );
  dff_sg \update_output_0/o_im_reg[1][13]  ( .D(n5672), .CP(clk), .Q(n9534) );
  dff_sg \update_output_0/o_im_reg[1][12]  ( .D(n5682), .CP(clk), .Q(n9535) );
  dff_sg \update_output_0/o_im_reg[1][11]  ( .D(n5676), .CP(clk), .Q(n9536) );
  dff_sg \update_output_0/o_im_reg[1][10]  ( .D(n5670), .CP(clk), .Q(n9537) );
  dff_sg \update_output_0/o_im_reg[1][9]  ( .D(n5681), .CP(clk), .Q(n9538) );
  dff_sg \update_output_0/o_im_reg[1][8]  ( .D(n5684), .CP(clk), .Q(n9539) );
  dff_sg \update_output_0/o_im_reg[1][7]  ( .D(n5668), .CP(clk), .Q(n9540) );
  dff_sg \update_output_0/o_im_reg[1][6]  ( .D(n5674), .CP(clk), .Q(n9541) );
  dff_sg \update_output_0/o_im_reg[1][5]  ( .D(n5821), .CP(clk), .Q(n9542) );
  dff_sg \update_output_0/o_im_reg[1][4]  ( .D(n5669), .CP(clk), .Q(n9543) );
  dff_sg \update_output_0/o_im_reg[1][3]  ( .D(n5680), .CP(clk), .Q(n9544) );
  dff_sg \update_output_0/o_im_reg[1][2]  ( .D(n5677), .CP(clk), .Q(n9545) );
  dff_sg \update_output_0/o_im_reg[1][1]  ( .D(n5667), .CP(clk), .Q(n9546) );
  dff_sg \update_output_0/o_im_reg[1][0]  ( .D(n5679), .CP(clk), .Q(n9547) );
  dff_sg \update_output_0/o_im_reg[10][19]  ( .D(n5851), .CP(clk), .Q(n9348)
         );
  dff_sg \update_output_0/o_im_reg[10][18]  ( .D(n5834), .CP(clk), .Q(n9349)
         );
  dff_sg \update_output_0/o_im_reg[10][17]  ( .D(n5830), .CP(clk), .Q(n9350)
         );
  dff_sg \update_output_0/o_im_reg[10][16]  ( .D(n5839), .CP(clk), .Q(n9351)
         );
  dff_sg \update_output_0/o_im_reg[10][15]  ( .D(n5838), .CP(clk), .Q(n9352)
         );
  dff_sg \update_output_0/o_im_reg[10][14]  ( .D(n5868), .CP(clk), .Q(n9353)
         );
  dff_sg \update_output_0/o_im_reg[10][13]  ( .D(n5867), .CP(clk), .Q(n9354)
         );
  dff_sg \update_output_0/o_im_reg[10][12]  ( .D(n5865), .CP(clk), .Q(n9355)
         );
  dff_sg \update_output_0/o_im_reg[10][11]  ( .D(n5869), .CP(clk), .Q(n9356)
         );
  dff_sg \update_output_0/o_im_reg[10][10]  ( .D(n5847), .CP(clk), .Q(n9357)
         );
  dff_sg \update_output_0/o_im_reg[10][9]  ( .D(n5846), .CP(clk), .Q(n9358) );
  dff_sg \update_output_0/o_im_reg[10][8]  ( .D(n5813), .CP(clk), .Q(n9359) );
  dff_sg \update_output_0/o_im_reg[10][7]  ( .D(n5814), .CP(clk), .Q(n9360) );
  dff_sg \update_output_0/o_im_reg[10][6]  ( .D(n5826), .CP(clk), .Q(n9361) );
  dff_sg \update_output_0/o_im_reg[10][5]  ( .D(n5822), .CP(clk), .Q(n9362) );
  dff_sg \update_output_0/o_im_reg[10][4]  ( .D(n5798), .CP(clk), .Q(n9363) );
  dff_sg \update_output_0/o_im_reg[10][3]  ( .D(n5794), .CP(clk), .Q(n9364) );
  dff_sg \update_output_0/o_im_reg[10][2]  ( .D(n5805), .CP(clk), .Q(n9365) );
  dff_sg \update_output_0/o_im_reg[10][1]  ( .D(n5806), .CP(clk), .Q(n9366) );
  dff_sg \update_output_0/o_im_reg[10][0]  ( .D(n5866), .CP(clk), .Q(n9367) );
  dff_sg \update_output_0/o_im_reg[2][19]  ( .D(n5854), .CP(clk), .Q(n9508) );
  dff_sg \update_output_0/o_im_reg[2][18]  ( .D(n5832), .CP(clk), .Q(n9509) );
  dff_sg \update_output_0/o_im_reg[2][17]  ( .D(n5828), .CP(clk), .Q(n9510) );
  dff_sg \update_output_0/o_im_reg[2][16]  ( .D(n5842), .CP(clk), .Q(n9511) );
  dff_sg \update_output_0/o_im_reg[2][15]  ( .D(n5836), .CP(clk), .Q(n9512) );
  dff_sg \update_output_0/o_im_reg[2][14]  ( .D(n5864), .CP(clk), .Q(n9513) );
  dff_sg \update_output_0/o_im_reg[2][13]  ( .D(n5862), .CP(clk), .Q(n9514) );
  dff_sg \update_output_0/o_im_reg[2][12]  ( .D(n5863), .CP(clk), .Q(n9515) );
  dff_sg \update_output_0/o_im_reg[2][11]  ( .D(n5860), .CP(clk), .Q(n9516) );
  dff_sg \update_output_0/o_im_reg[2][10]  ( .D(n5850), .CP(clk), .Q(n9517) );
  dff_sg \update_output_0/o_im_reg[2][9]  ( .D(n5844), .CP(clk), .Q(n9518) );
  dff_sg \update_output_0/o_im_reg[2][8]  ( .D(n5811), .CP(clk), .Q(n9519) );
  dff_sg \update_output_0/o_im_reg[2][7]  ( .D(n5817), .CP(clk), .Q(n9520) );
  dff_sg \update_output_0/o_im_reg[2][6]  ( .D(n5824), .CP(clk), .Q(n9521) );
  dff_sg \update_output_0/o_im_reg[2][5]  ( .D(n5820), .CP(clk), .Q(n9522) );
  dff_sg \update_output_0/o_im_reg[2][4]  ( .D(n5801), .CP(clk), .Q(n9523) );
  dff_sg \update_output_0/o_im_reg[2][3]  ( .D(n5796), .CP(clk), .Q(n9524) );
  dff_sg \update_output_0/o_im_reg[2][2]  ( .D(n5804), .CP(clk), .Q(n9525) );
  dff_sg \update_output_0/o_im_reg[2][1]  ( .D(n5809), .CP(clk), .Q(n9526) );
  dff_sg \update_output_0/o_im_reg[2][0]  ( .D(n5861), .CP(clk), .Q(n9527) );
  dff_sg \update_output_0/o_im_reg[0][19]  ( .D(n5853), .CP(clk), .Q(n9548) );
  dff_sg \update_output_0/o_im_reg[0][18]  ( .D(n5831), .CP(clk), .Q(n9549) );
  dff_sg \update_output_0/o_im_reg[0][17]  ( .D(n5827), .CP(clk), .Q(n9550) );
  dff_sg \update_output_0/o_im_reg[0][16]  ( .D(n5841), .CP(clk), .Q(n9551) );
  dff_sg \update_output_0/o_im_reg[0][15]  ( .D(n5835), .CP(clk), .Q(n9552) );
  dff_sg \update_output_0/o_im_reg[0][14]  ( .D(n5855), .CP(clk), .Q(n9553) );
  dff_sg \update_output_0/o_im_reg[0][13]  ( .D(n5858), .CP(clk), .Q(n9554) );
  dff_sg \update_output_0/o_im_reg[0][12]  ( .D(n5856), .CP(clk), .Q(n9555) );
  dff_sg \update_output_0/o_im_reg[0][11]  ( .D(n5859), .CP(clk), .Q(n9556) );
  dff_sg \update_output_0/o_im_reg[0][10]  ( .D(n5849), .CP(clk), .Q(n9557) );
  dff_sg \update_output_0/o_im_reg[0][9]  ( .D(n5843), .CP(clk), .Q(n9558) );
  dff_sg \update_output_0/o_im_reg[0][8]  ( .D(n5810), .CP(clk), .Q(n9559) );
  dff_sg \update_output_0/o_im_reg[0][7]  ( .D(n5816), .CP(clk), .Q(n9560) );
  dff_sg \update_output_0/o_im_reg[0][6]  ( .D(n5823), .CP(clk), .Q(n9561) );
  dff_sg \update_output_0/o_im_reg[0][5]  ( .D(n5818), .CP(clk), .Q(n9562) );
  dff_sg \update_output_0/o_im_reg[0][4]  ( .D(n5800), .CP(clk), .Q(n9563) );
  dff_sg \update_output_0/o_im_reg[0][3]  ( .D(n5795), .CP(clk), .Q(n9564) );
  dff_sg \update_output_0/o_im_reg[0][2]  ( .D(n5802), .CP(clk), .Q(n9565) );
  dff_sg \update_output_0/o_im_reg[0][1]  ( .D(n5808), .CP(clk), .Q(n9566) );
  dff_sg \update_output_0/o_im_reg[0][0]  ( .D(n5857), .CP(clk), .Q(n9567) );
  dff_sg \update_output_0/o_im_reg[8][19]  ( .D(n5787), .CP(clk), .Q(n9388) );
  dff_sg \update_output_0/o_im_reg[8][18]  ( .D(n5792), .CP(clk), .Q(n9389) );
  dff_sg \update_output_0/o_im_reg[8][17]  ( .D(n5782), .CP(clk), .Q(n9390) );
  dff_sg \update_output_0/o_im_reg[8][16]  ( .D(n5773), .CP(clk), .Q(n9391) );
  dff_sg \update_output_0/o_im_reg[8][15]  ( .D(n5786), .CP(clk), .Q(n9392) );
  dff_sg \update_output_0/o_im_reg[8][14]  ( .D(n5781), .CP(clk), .Q(n9393) );
  dff_sg \update_output_0/o_im_reg[8][13]  ( .D(n5785), .CP(clk), .Q(n9394) );
  dff_sg \update_output_0/o_im_reg[8][12]  ( .D(n5780), .CP(clk), .Q(n9395) );
  dff_sg \update_output_0/o_im_reg[8][11]  ( .D(n5775), .CP(clk), .Q(n9396) );
  dff_sg \update_output_0/o_im_reg[8][10]  ( .D(n5778), .CP(clk), .Q(n9397) );
  dff_sg \update_output_0/o_im_reg[8][9]  ( .D(n5788), .CP(clk), .Q(n9398) );
  dff_sg \update_output_0/o_im_reg[8][8]  ( .D(n5774), .CP(clk), .Q(n9399) );
  dff_sg \update_output_0/o_im_reg[8][7]  ( .D(n5789), .CP(clk), .Q(n9400) );
  dff_sg \update_output_0/o_im_reg[8][6]  ( .D(n5776), .CP(clk), .Q(n9401) );
  dff_sg \update_output_0/o_im_reg[8][5]  ( .D(n5784), .CP(clk), .Q(n9402) );
  dff_sg \update_output_0/o_im_reg[8][4]  ( .D(n5783), .CP(clk), .Q(n9403) );
  dff_sg \update_output_0/o_im_reg[8][3]  ( .D(n5777), .CP(clk), .Q(n9404) );
  dff_sg \update_output_0/o_im_reg[8][2]  ( .D(n5779), .CP(clk), .Q(n9405) );
  dff_sg \update_output_0/o_im_reg[8][1]  ( .D(n5790), .CP(clk), .Q(n9406) );
  dff_sg \update_output_0/o_im_reg[8][0]  ( .D(n5791), .CP(clk), .Q(n9407) );
  dff_sg \update_output_0/o_im_reg[7][19]  ( .D(n5727), .CP(clk), .Q(n9408) );
  dff_sg \update_output_0/o_im_reg[7][18]  ( .D(n5724), .CP(clk), .Q(n9409) );
  dff_sg \update_output_0/o_im_reg[7][17]  ( .D(n5717), .CP(clk), .Q(n9410) );
  dff_sg \update_output_0/o_im_reg[7][16]  ( .D(n5721), .CP(clk), .Q(n9411) );
  dff_sg \update_output_0/o_im_reg[7][15]  ( .D(n5716), .CP(clk), .Q(n9412) );
  dff_sg \update_output_0/o_im_reg[7][14]  ( .D(n5725), .CP(clk), .Q(n9413) );
  dff_sg \update_output_0/o_im_reg[7][13]  ( .D(n5711), .CP(clk), .Q(n9414) );
  dff_sg \update_output_0/o_im_reg[7][12]  ( .D(n5723), .CP(clk), .Q(n9415) );
  dff_sg \update_output_0/o_im_reg[7][11]  ( .D(n5713), .CP(clk), .Q(n9416) );
  dff_sg \update_output_0/o_im_reg[7][10]  ( .D(n5714), .CP(clk), .Q(n9417) );
  dff_sg \update_output_0/o_im_reg[7][9]  ( .D(n5729), .CP(clk), .Q(n9418) );
  dff_sg \update_output_0/o_im_reg[7][8]  ( .D(n5710), .CP(clk), .Q(n9419) );
  dff_sg \update_output_0/o_im_reg[7][7]  ( .D(n5715), .CP(clk), .Q(n9420) );
  dff_sg \update_output_0/o_im_reg[7][6]  ( .D(n5719), .CP(clk), .Q(n9421) );
  dff_sg \update_output_0/o_im_reg[7][5]  ( .D(n5726), .CP(clk), .Q(n9422) );
  dff_sg \update_output_0/o_im_reg[7][4]  ( .D(n5728), .CP(clk), .Q(n9423) );
  dff_sg \update_output_0/o_im_reg[7][3]  ( .D(n5722), .CP(clk), .Q(n9424) );
  dff_sg \update_output_0/o_im_reg[7][2]  ( .D(n5718), .CP(clk), .Q(n9425) );
  dff_sg \update_output_0/o_im_reg[7][1]  ( .D(n5720), .CP(clk), .Q(n9426) );
  dff_sg \update_output_0/o_im_reg[7][0]  ( .D(n5712), .CP(clk), .Q(n9427) );
  dff_sg \update_output_0/o_im_reg[15][19]  ( .D(n5747), .CP(clk), .Q(n9248)
         );
  dff_sg \update_output_0/o_im_reg[15][18]  ( .D(n5739), .CP(clk), .Q(n9249)
         );
  dff_sg \update_output_0/o_im_reg[15][17]  ( .D(n5745), .CP(clk), .Q(n9250)
         );
  dff_sg \update_output_0/o_im_reg[15][16]  ( .D(n5742), .CP(clk), .Q(n9251)
         );
  dff_sg \update_output_0/o_im_reg[15][15]  ( .D(n5732), .CP(clk), .Q(n9252)
         );
  dff_sg \update_output_0/o_im_reg[15][14]  ( .D(n5734), .CP(clk), .Q(n9253)
         );
  dff_sg \update_output_0/o_im_reg[15][13]  ( .D(n5740), .CP(clk), .Q(n9254)
         );
  dff_sg \update_output_0/o_im_reg[15][12]  ( .D(n5731), .CP(clk), .Q(n9255)
         );
  dff_sg \update_output_0/o_im_reg[15][11]  ( .D(n5735), .CP(clk), .Q(n9256)
         );
  dff_sg \update_output_0/o_im_reg[15][10]  ( .D(n5736), .CP(clk), .Q(n9257)
         );
  dff_sg \update_output_0/o_im_reg[15][9]  ( .D(n5748), .CP(clk), .Q(n9258) );
  dff_sg \update_output_0/o_im_reg[15][8]  ( .D(n5744), .CP(clk), .Q(n9259) );
  dff_sg \update_output_0/o_im_reg[15][7]  ( .D(n5746), .CP(clk), .Q(n9260) );
  dff_sg \update_output_0/o_im_reg[15][6]  ( .D(n5733), .CP(clk), .Q(n9261) );
  dff_sg \update_output_0/o_im_reg[15][5]  ( .D(n5738), .CP(clk), .Q(n9262) );
  dff_sg \update_output_0/o_im_reg[15][4]  ( .D(n5730), .CP(clk), .Q(n9263) );
  dff_sg \update_output_0/o_im_reg[15][3]  ( .D(n5743), .CP(clk), .Q(n9264) );
  dff_sg \update_output_0/o_im_reg[15][2]  ( .D(n5749), .CP(clk), .Q(n9265) );
  dff_sg \update_output_0/o_im_reg[15][1]  ( .D(n5741), .CP(clk), .Q(n9266) );
  dff_sg \update_output_0/o_im_reg[15][0]  ( .D(n5737), .CP(clk), .Q(n9267) );
  dff_sg \update_output_0/o_pointer_reg[3]  ( .D(n5751), .CP(clk), .Q(
        \update_output_0/N34 ) );
  dff_sg \update_output_0/o_pointer_reg[2]  ( .D(n5750), .CP(clk), .Q(
        \update_output_0/N33 ) );
  dff_sg \update_output_0/o_pointer_reg[1]  ( .D(\update_output_0/n3549 ), 
        .CP(clk), .Q(\update_output_0/N32 ) );
  dff_sg \update_output_0/o_pointer_reg[0]  ( .D(n5752), .CP(clk), .Q(
        \update_output_0/N31 ) );
  dff_sg \update_output_0/i_pointer_reg[3]  ( .D(n5705), .CP(clk), .Q(
        \update_output_0/N30 ) );
  dff_sg \update_output_0/state_reg[1]  ( .D(n5708), .CP(clk), .Q(
        \update_output_0/n9019 ) );
  dff_sg \update_output_0/state_reg[0]  ( .D(n5709), .CP(clk), .Q(
        \update_output_0/n9020 ) );
  dff_sg \update_output_0/i_pointer_reg[2]  ( .D(n5706), .CP(clk), .Q(
        \update_output_0/N29 ) );
  dff_sg \update_output_0/i_pointer_reg[1]  ( .D(n5707), .CP(clk), .Q(
        \update_output_0/N28 ) );
  dff_sg \update_output_0/i_pointer_reg[0]  ( .D(n5793), .CP(clk), .Q(
        \update_output_0/N27 ) );
  nor_x2_sg U3714 ( .A(n3092), .B(n3095), .X(n3094) );
  nand_x8_sg U4846 ( .A(n9195), .B(n3886), .X(n3828) );
  nand_x8_sg U4907 ( .A(n9195), .B(n3928), .X(n3889) );
  nand_x8_sg U4970 ( .A(n3974), .B(n3928), .X(n3935) );
  nand_x8_sg U5031 ( .A(n3974), .B(n3886), .X(n3977) );
  nand_x8_sg U5032 ( .A(n7419), .B(n4016), .X(n3974) );
  nor_x2_sg U5292 ( .A(reset), .B(n4202), .X(n4203) );
  nand_x8_sg U5355 ( .A(n3886), .B(n4249), .X(n4210) );
  nand_x8_sg U5416 ( .A(n3928), .B(n4249), .X(n4252) );
  nand_x8_sg U5417 ( .A(n7419), .B(n9193), .X(n4249) );
  nand_x8_sg U5434 ( .A(n9192), .B(n4307), .X(n3092) );
  nor_x2_sg U5498 ( .A(n4306), .B(n7571), .X(n4179) );
  nor_x2_sg U5585 ( .A(\update_output_0/n6687 ), .B(n7435), .X(n4421) );
  nor_x2_sg U5586 ( .A(\update_output_0/n6667 ), .B(n7433), .X(n4420) );
  nor_x2_sg U5596 ( .A(\update_output_0/n6547 ), .B(n7429), .X(n4432) );
  nor_x2_sg U5598 ( .A(n4440), .B(n7570), .X(n4439) );
  nor_x2_sg U5599 ( .A(n4441), .B(n4442), .X(n4440) );
  nor_x2_sg U5603 ( .A(n4446), .B(n4447), .X(n4441) );
  nor_x2_sg U5606 ( .A(n7541), .B(n5514), .X(n4446) );
  nor_x2_sg U5607 ( .A(\update_output_0/n6567 ), .B(n7428), .X(n4438) );
  nor_x2_sg U5632 ( .A(\update_output_0/n6688 ), .B(n7434), .X(n4471) );
  nor_x2_sg U5633 ( .A(\update_output_0/n6668 ), .B(n7432), .X(n4470) );
  nor_x2_sg U5643 ( .A(\update_output_0/n6548 ), .B(n7429), .X(n4479) );
  nor_x2_sg U5645 ( .A(n4485), .B(n7570), .X(n4484) );
  nor_x2_sg U5646 ( .A(n4486), .B(n4487), .X(n4485) );
  nor_x2_sg U5650 ( .A(n4490), .B(n4491), .X(n4486) );
  nor_x2_sg U5653 ( .A(n7541), .B(n5503), .X(n4490) );
  nor_x2_sg U5654 ( .A(\update_output_0/n6568 ), .B(n7427), .X(n4483) );
  nor_x2_sg U5679 ( .A(\update_output_0/n6686 ), .B(n4422), .X(n4513) );
  nor_x2_sg U5680 ( .A(\update_output_0/n6666 ), .B(n4423), .X(n4512) );
  nor_x2_sg U5690 ( .A(\update_output_0/n6546 ), .B(n7429), .X(n4521) );
  nor_x2_sg U5692 ( .A(n4527), .B(n7570), .X(n4526) );
  nor_x2_sg U5693 ( .A(n4528), .B(n4529), .X(n4527) );
  nor_x2_sg U5697 ( .A(n4532), .B(n4533), .X(n4528) );
  nor_x2_sg U5700 ( .A(n7540), .B(n5525), .X(n4532) );
  nor_x2_sg U5701 ( .A(\update_output_0/n6566 ), .B(n4303), .X(n4525) );
  nor_x2_sg U5726 ( .A(\update_output_0/n6685 ), .B(n7435), .X(n4555) );
  nor_x2_sg U5727 ( .A(\update_output_0/n6665 ), .B(n7433), .X(n4554) );
  nor_x2_sg U5737 ( .A(\update_output_0/n6545 ), .B(n7429), .X(n4563) );
  nor_x2_sg U5739 ( .A(n4569), .B(n7570), .X(n4568) );
  nor_x2_sg U5740 ( .A(n4570), .B(n4571), .X(n4569) );
  nor_x2_sg U5744 ( .A(n4574), .B(n4575), .X(n4570) );
  nor_x2_sg U5747 ( .A(n7540), .B(n5536), .X(n4574) );
  nor_x2_sg U5748 ( .A(\update_output_0/n6565 ), .B(n7428), .X(n4567) );
  nor_x2_sg U5773 ( .A(\update_output_0/n6692 ), .B(n7434), .X(n4597) );
  nor_x2_sg U5774 ( .A(\update_output_0/n6672 ), .B(n7432), .X(n4596) );
  nor_x2_sg U5784 ( .A(\update_output_0/n6552 ), .B(n7429), .X(n4605) );
  nor_x2_sg U5786 ( .A(n4611), .B(n7570), .X(n4610) );
  nor_x2_sg U5787 ( .A(n4612), .B(n4613), .X(n4611) );
  nor_x2_sg U5791 ( .A(n4616), .B(n4617), .X(n4612) );
  nor_x2_sg U5794 ( .A(n7540), .B(n5459), .X(n4616) );
  nor_x2_sg U5795 ( .A(\update_output_0/n6572 ), .B(n7427), .X(n4609) );
  nor_x2_sg U5820 ( .A(\update_output_0/n6691 ), .B(n4422), .X(n4639) );
  nor_x2_sg U5821 ( .A(\update_output_0/n6671 ), .B(n4423), .X(n4638) );
  nor_x2_sg U5831 ( .A(\update_output_0/n6551 ), .B(n7429), .X(n4647) );
  nor_x2_sg U5833 ( .A(n4653), .B(n7570), .X(n4652) );
  nor_x2_sg U5834 ( .A(n4654), .B(n4655), .X(n4653) );
  nor_x2_sg U5838 ( .A(n4658), .B(n4659), .X(n4654) );
  nor_x2_sg U5841 ( .A(n7541), .B(n5470), .X(n4658) );
  nor_x2_sg U5842 ( .A(\update_output_0/n6571 ), .B(n4303), .X(n4651) );
  nor_x2_sg U5870 ( .A(\update_output_0/n6689 ), .B(n7435), .X(n4683) );
  nor_x2_sg U5871 ( .A(\update_output_0/n6669 ), .B(n7433), .X(n4682) );
  nor_x2_sg U5881 ( .A(\update_output_0/n6549 ), .B(n7429), .X(n4691) );
  nor_x2_sg U5883 ( .A(n4697), .B(n7570), .X(n4696) );
  nor_x2_sg U5884 ( .A(n4698), .B(n4699), .X(n4697) );
  nor_x2_sg U5888 ( .A(n4702), .B(n4703), .X(n4698) );
  nor_x2_sg U5891 ( .A(n7540), .B(n5492), .X(n4702) );
  nor_x2_sg U5892 ( .A(\update_output_0/n6569 ), .B(n7428), .X(n4695) );
  nor_x2_sg U5917 ( .A(\update_output_0/n6690 ), .B(n7434), .X(n4725) );
  nor_x2_sg U5918 ( .A(\update_output_0/n6670 ), .B(n7432), .X(n4724) );
  nor_x2_sg U5928 ( .A(\update_output_0/n6550 ), .B(n7429), .X(n4733) );
  nor_x2_sg U5930 ( .A(n4739), .B(n7570), .X(n4738) );
  nor_x2_sg U5931 ( .A(n4740), .B(n4741), .X(n4739) );
  nor_x2_sg U5935 ( .A(n4744), .B(n4745), .X(n4740) );
  nor_x2_sg U5938 ( .A(n7541), .B(n5481), .X(n4744) );
  nor_x2_sg U5939 ( .A(\update_output_0/n6570 ), .B(n7427), .X(n4737) );
  nor_x2_sg U5964 ( .A(\update_output_0/n6701 ), .B(n4422), .X(n4767) );
  nor_x2_sg U5965 ( .A(\update_output_0/n6681 ), .B(n4423), .X(n4766) );
  nor_x2_sg U5975 ( .A(\update_output_0/n6561 ), .B(n7429), .X(n4775) );
  nor_x2_sg U5977 ( .A(n4781), .B(n7570), .X(n4780) );
  nor_x2_sg U5978 ( .A(n4782), .B(n4783), .X(n4781) );
  nor_x2_sg U5982 ( .A(n4786), .B(n4787), .X(n4782) );
  nor_x2_sg U5985 ( .A(n7541), .B(n5360), .X(n4786) );
  nor_x2_sg U5986 ( .A(\update_output_0/n6581 ), .B(n4303), .X(n4779) );
  nor_x2_sg U6011 ( .A(\update_output_0/n6702 ), .B(n7435), .X(n4809) );
  nor_x2_sg U6012 ( .A(\update_output_0/n6682 ), .B(n7433), .X(n4808) );
  nor_x2_sg U6022 ( .A(\update_output_0/n6562 ), .B(n7429), .X(n4817) );
  nor_x2_sg U6024 ( .A(n4823), .B(n7570), .X(n4822) );
  nor_x2_sg U6025 ( .A(n4824), .B(n4825), .X(n4823) );
  nor_x2_sg U6029 ( .A(n4828), .B(n4829), .X(n4824) );
  nor_x2_sg U6032 ( .A(n7541), .B(n5349), .X(n4828) );
  nor_x2_sg U6033 ( .A(\update_output_0/n6582 ), .B(n7428), .X(n4821) );
  nor_x2_sg U6058 ( .A(\update_output_0/n6699 ), .B(n7434), .X(n4851) );
  nor_x2_sg U6059 ( .A(\update_output_0/n6679 ), .B(n7432), .X(n4850) );
  nor_x2_sg U6069 ( .A(\update_output_0/n6559 ), .B(n7429), .X(n4859) );
  nor_x2_sg U6071 ( .A(n4865), .B(n7570), .X(n4864) );
  nor_x2_sg U6072 ( .A(n4866), .B(n4867), .X(n4865) );
  nor_x2_sg U6076 ( .A(n4870), .B(n4871), .X(n4866) );
  nor_x2_sg U6079 ( .A(n7541), .B(n5382), .X(n4870) );
  nor_x2_sg U6080 ( .A(\update_output_0/n6579 ), .B(n7427), .X(n4863) );
  nor_x2_sg U6105 ( .A(\update_output_0/n6700 ), .B(n4422), .X(n4893) );
  nor_x2_sg U6106 ( .A(\update_output_0/n6680 ), .B(n4423), .X(n4892) );
  nor_x2_sg U6116 ( .A(\update_output_0/n6560 ), .B(n7429), .X(n4901) );
  nor_x2_sg U6118 ( .A(n4907), .B(n7570), .X(n4906) );
  nor_x2_sg U6119 ( .A(n4908), .B(n4909), .X(n4907) );
  nor_x2_sg U6123 ( .A(n4912), .B(n4913), .X(n4908) );
  nor_x2_sg U6126 ( .A(n7540), .B(n5371), .X(n4912) );
  nor_x2_sg U6127 ( .A(\update_output_0/n6580 ), .B(n4303), .X(n4905) );
  nor_x2_sg U6152 ( .A(\update_output_0/n6693 ), .B(n7435), .X(n4935) );
  nor_x2_sg U6153 ( .A(\update_output_0/n6673 ), .B(n7433), .X(n4934) );
  nor_x2_sg U6163 ( .A(\update_output_0/n6553 ), .B(n3932), .X(n4943) );
  nor_x2_sg U6165 ( .A(n4949), .B(n7570), .X(n4948) );
  nor_x2_sg U6166 ( .A(n4950), .B(n4951), .X(n4949) );
  nor_x2_sg U6170 ( .A(n4954), .B(n4955), .X(n4950) );
  nor_x2_sg U6173 ( .A(n7540), .B(n5448), .X(n4954) );
  nor_x2_sg U6174 ( .A(\update_output_0/n6573 ), .B(n7428), .X(n4947) );
  nor_x2_sg U6199 ( .A(\update_output_0/n6694 ), .B(n7434), .X(n4977) );
  nor_x2_sg U6200 ( .A(\update_output_0/n6674 ), .B(n7432), .X(n4976) );
  nor_x2_sg U6210 ( .A(\update_output_0/n6554 ), .B(n7429), .X(n4985) );
  nor_x2_sg U6212 ( .A(n4991), .B(n7570), .X(n4990) );
  nor_x2_sg U6213 ( .A(n4992), .B(n4993), .X(n4991) );
  nor_x2_sg U6217 ( .A(n4996), .B(n4997), .X(n4992) );
  nor_x2_sg U6220 ( .A(n7540), .B(n5437), .X(n4996) );
  nor_x2_sg U6221 ( .A(\update_output_0/n6574 ), .B(n7427), .X(n4989) );
  nor_x2_sg U6246 ( .A(\update_output_0/n6703 ), .B(n4422), .X(n5019) );
  nor_x2_sg U6247 ( .A(\update_output_0/n6683 ), .B(n4423), .X(n5018) );
  nor_x2_sg U6257 ( .A(\update_output_0/n6563 ), .B(n3932), .X(n5027) );
  nor_x2_sg U6259 ( .A(n5033), .B(n7570), .X(n5032) );
  nor_x2_sg U6260 ( .A(n5034), .B(n5035), .X(n5033) );
  nor_x2_sg U6264 ( .A(n5038), .B(n5039), .X(n5034) );
  nor_x2_sg U6267 ( .A(n7541), .B(n5338), .X(n5038) );
  nor_x2_sg U6268 ( .A(\update_output_0/n6583 ), .B(n4303), .X(n5031) );
  nor_x2_sg U6290 ( .A(n4306), .B(n7570), .X(n4392) );
  nand_x8_sg U6291 ( .A(n4182), .B(n7540), .X(n4306) );
  nand_x8_sg U6307 ( .A(n5064), .B(n3886), .X(n4404) );
  nand_x8_sg U6308 ( .A(n7419), .B(n3098), .X(n3886) );
  nand_x8_sg U6324 ( .A(n5064), .B(n3928), .X(n4398) );
  nand_x8_sg U6325 ( .A(n7419), .B(n4393), .X(n3928) );
  nand_x8_sg U6326 ( .A(n7419), .B(n5075), .X(n5064) );
  nor_x2_sg U6337 ( .A(n7570), .B(n3095), .X(n4099) );
  nor_x2_sg U6347 ( .A(\update_output_0/n6698 ), .B(n7435), .X(n5091) );
  nor_x2_sg U6348 ( .A(\update_output_0/n6678 ), .B(n7433), .X(n5090) );
  nor_x2_sg U6358 ( .A(\update_output_0/n6558 ), .B(n7429), .X(n5099) );
  nor_x2_sg U6360 ( .A(n5105), .B(n7570), .X(n5104) );
  nor_x2_sg U6361 ( .A(n5106), .B(n5107), .X(n5105) );
  nor_x2_sg U6365 ( .A(n5110), .B(n5111), .X(n5106) );
  nor_x2_sg U6368 ( .A(n7541), .B(n5393), .X(n5110) );
  nor_x2_sg U6369 ( .A(\update_output_0/n6578 ), .B(n7428), .X(n5103) );
  nor_x2_sg U6384 ( .A(\update_output_0/n6697 ), .B(n7434), .X(n5127) );
  nor_x2_sg U6385 ( .A(\update_output_0/n6677 ), .B(n7432), .X(n5126) );
  nor_x2_sg U6395 ( .A(\update_output_0/n6557 ), .B(n3932), .X(n5135) );
  nor_x2_sg U6397 ( .A(n5141), .B(n7570), .X(n5140) );
  nor_x2_sg U6398 ( .A(n5142), .B(n5143), .X(n5141) );
  nor_x2_sg U6402 ( .A(n5146), .B(n5147), .X(n5142) );
  nor_x2_sg U6405 ( .A(n7541), .B(n5404), .X(n5146) );
  nor_x2_sg U6406 ( .A(\update_output_0/n6577 ), .B(n7427), .X(n5139) );
  nor_x2_sg U6422 ( .A(\update_output_0/n6695 ), .B(n4422), .X(n5163) );
  nor_x2_sg U6423 ( .A(\update_output_0/n6675 ), .B(n4423), .X(n5162) );
  nor_x2_sg U6433 ( .A(\update_output_0/n6555 ), .B(n7429), .X(n5171) );
  nor_x2_sg U6435 ( .A(n5177), .B(n7570), .X(n5176) );
  nor_x2_sg U6436 ( .A(n5178), .B(n5179), .X(n5177) );
  nor_x2_sg U6440 ( .A(n5182), .B(n5183), .X(n5178) );
  nor_x2_sg U6443 ( .A(n7541), .B(n5426), .X(n5182) );
  nor_x2_sg U6444 ( .A(\update_output_0/n6575 ), .B(n4303), .X(n5175) );
  nor_x2_sg U6466 ( .A(\update_output_0/n6696 ), .B(n7435), .X(n5203) );
  nor_x2_sg U6467 ( .A(\update_output_0/n6676 ), .B(n7433), .X(n5202) );
  nor_x2_sg U6477 ( .A(\update_output_0/n6556 ), .B(n3932), .X(n5211) );
  nor_x2_sg U6479 ( .A(n5217), .B(n7570), .X(n5216) );
  nor_x2_sg U6480 ( .A(n5218), .B(n5219), .X(n5217) );
  nor_x2_sg U6484 ( .A(n5222), .B(n5223), .X(n5218) );
  nor_x2_sg U6487 ( .A(n7540), .B(n5415), .X(n5222) );
  nor_x2_sg U6488 ( .A(\update_output_0/n6576 ), .B(n7428), .X(n5215) );
  nor_x2_sg U6507 ( .A(\update_output_0/n6684 ), .B(n7434), .X(n5240) );
  nand_x8_sg U6508 ( .A(n9240), .B(n5241), .X(n4422) );
  nor_x2_sg U6509 ( .A(\update_output_0/n6664 ), .B(n7432), .X(n5239) );
  nand_x8_sg U6510 ( .A(n9240), .B(n5242), .X(n4423) );
  nor_x2_sg U6524 ( .A(\update_output_0/n6544 ), .B(n7429), .X(n5250) );
  nand_x8_sg U6525 ( .A(n7570), .B(n7323), .X(n3932) );
  nor_x2_sg U6527 ( .A(n5256), .B(n7570), .X(n5255) );
  nor_x2_sg U6528 ( .A(n5257), .B(n5258), .X(n5256) );
  nor_x2_sg U6532 ( .A(n5261), .B(n5262), .X(n5257) );
  nor_x2_sg U6535 ( .A(n7541), .B(n5547), .X(n5261) );
  nor_x2_sg U6536 ( .A(\update_output_0/n6564 ), .B(n7427), .X(n5254) );
  nand_x8_sg U6537 ( .A(n7570), .B(n7558), .X(n4303) );
  nand_x8_sg U6541 ( .A(n6381), .B(n7571), .X(n4297) );
  nand_x8_sg U6544 ( .A(n6381), .B(n7570), .X(n5236) );
  nand_x8_sg U6549 ( .A(n5241), .B(n4182), .X(n3095) );
  nand_x8_sg U6552 ( .A(n9197), .B(n5268), .X(n3930) );
  nor_x2_sg U6568 ( .A(n5283), .B(n5284), .X(n3816) );
  nor_x2_sg U6571 ( .A(n5286), .B(n5274), .X(n5285) );
  nand_x8_sg U6577 ( .A(n5290), .B(n5291), .X(n5283) );
  nand_x8_sg U6597 ( .A(n5292), .B(n5274), .X(n5290) );
  nand_x8_sg U6598 ( .A(n5292), .B(n5307), .X(n5274) );
  nor_x2_sg U6618 ( .A(n5323), .B(n5324), .X(n5322) );
  \**FFGEN**  \update_mask_0/increment_reg  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(\update_mask_0/n991 ), .force_10(
        n5928), .force_11(1'b0), .QN(\update_mask_0/n919 ) );
  \**FFGEN**  \update_mask_0/o_mask_reg[31]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(n756), .force_10(
        \update_mask_0/n996 ), .force_11(1'b0), .Q(o_mask[31]) );
  \**FFGEN**  \update_mask_0/o_mask_reg[30]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(n759), .force_10(
        \update_mask_0/n1000 ), .force_11(1'b0), .Q(o_mask[30]) );
  \**FFGEN**  \update_mask_0/o_mask_reg[29]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(n762), .force_10(
        \update_mask_0/n1004 ), .force_11(1'b0), .Q(o_mask[29]) );
  \**FFGEN**  \update_mask_0/o_mask_reg[28]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(n765), .force_10(
        \update_mask_0/n1008 ), .force_11(1'b0), .Q(o_mask[28]) );
  \**FFGEN**  \update_mask_0/o_mask_reg[27]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(n768), .force_10(
        \update_mask_0/n1012 ), .force_11(1'b0), .Q(o_mask[27]) );
  \**FFGEN**  \update_mask_0/o_mask_reg[26]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(n771), .force_10(
        \update_mask_0/n1016 ), .force_11(1'b0), .Q(o_mask[26]) );
  \**FFGEN**  \update_mask_0/o_mask_reg[25]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(n769), .force_10(
        \update_mask_0/n1020 ), .force_11(1'b0), .Q(o_mask[25]) );
  \**FFGEN**  \update_mask_0/o_mask_reg[24]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(n770), .force_10(
        \update_mask_0/n1024 ), .force_11(1'b0), .Q(o_mask[24]) );
  \**FFGEN**  \update_mask_0/o_mask_reg[23]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(n766), .force_10(
        \update_mask_0/n1028 ), .force_11(1'b0), .Q(o_mask[23]) );
  \**FFGEN**  \update_mask_0/o_mask_reg[22]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(n767), .force_10(
        \update_mask_0/n1032 ), .force_11(1'b0), .Q(o_mask[22]) );
  \**FFGEN**  \update_mask_0/o_mask_reg[21]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(n763), .force_10(
        \update_mask_0/n1036 ), .force_11(1'b0), .Q(o_mask[21]) );
  \**FFGEN**  \update_mask_0/o_mask_reg[20]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(n764), .force_10(
        \update_mask_0/n1040 ), .force_11(1'b0), .Q(o_mask[20]) );
  \**FFGEN**  \update_mask_0/o_mask_reg[19]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(n760), .force_10(
        \update_mask_0/n1044 ), .force_11(1'b0), .Q(o_mask[19]) );
  \**FFGEN**  \update_mask_0/o_mask_reg[18]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(n761), .force_10(
        \update_mask_0/n1048 ), .force_11(1'b0), .Q(o_mask[18]) );
  \**FFGEN**  \update_mask_0/o_mask_reg[17]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(n746), .force_10(
        \update_mask_0/n1052 ), .force_11(1'b0), .Q(o_mask[17]) );
  \**FFGEN**  \update_mask_0/o_mask_reg[16]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(n753), .force_10(
        \update_mask_0/n1056 ), .force_11(1'b0), .Q(o_mask[16]) );
  \**FFGEN**  \update_mask_0/o_mask_reg[15]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(n751), .force_10(
        \update_mask_0/n1060 ), .force_11(1'b0), .Q(o_mask[15]) );
  \**FFGEN**  \update_mask_0/o_mask_reg[14]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(n752), .force_10(
        \update_mask_0/n1064 ), .force_11(1'b0), .Q(o_mask[14]) );
  \**FFGEN**  \update_mask_0/o_mask_reg[13]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(n741), .force_10(
        \update_mask_0/n1068 ), .force_11(1'b0), .Q(o_mask[13]) );
  \**FFGEN**  \update_mask_0/o_mask_reg[12]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(n742), .force_10(
        \update_mask_0/n1072 ), .force_11(1'b0), .Q(o_mask[12]) );
  \**FFGEN**  \update_mask_0/o_mask_reg[11]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(n740), .force_10(
        \update_mask_0/n1076 ), .force_11(1'b0), .Q(o_mask[11]) );
  \**FFGEN**  \update_mask_0/o_mask_reg[10]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(n744), .force_10(
        \update_mask_0/n1080 ), .force_11(1'b0), .Q(o_mask[10]) );
  \**FFGEN**  \update_mask_0/o_mask_reg[9]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(n743), .force_10(
        \update_mask_0/n1084 ), .force_11(1'b0), .Q(o_mask[9]) );
  \**FFGEN**  \update_mask_0/o_mask_reg[8]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(n745), .force_10(
        \update_mask_0/n1088 ), .force_11(1'b0), .Q(o_mask[8]) );
  \**FFGEN**  \update_mask_0/o_mask_reg[7]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(n750), .force_10(
        \update_mask_0/n1092 ), .force_11(1'b0), .Q(o_mask[7]) );
  \**FFGEN**  \update_mask_0/o_mask_reg[6]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(n748), .force_10(
        \update_mask_0/n1096 ), .force_11(1'b0), .Q(o_mask[6]) );
  \**FFGEN**  \update_mask_0/o_mask_reg[5]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(n757), .force_10(
        \update_mask_0/n1100 ), .force_11(1'b0), .Q(o_mask[5]) );
  \**FFGEN**  \update_mask_0/o_mask_reg[4]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(n758), .force_10(
        \update_mask_0/n1104 ), .force_11(1'b0), .Q(o_mask[4]) );
  \**FFGEN**  \update_mask_0/o_mask_reg[3]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(n754), .force_10(
        \update_mask_0/n1108 ), .force_11(1'b0), .Q(o_mask[3]) );
  \**FFGEN**  \update_mask_0/o_mask_reg[2]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(n755), .force_10(
        \update_mask_0/n1112 ), .force_11(1'b0), .Q(o_mask[2]) );
  \**FFGEN**  \update_mask_0/o_mask_reg[1]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(n747), .force_10(
        \update_mask_0/n1116 ), .force_11(1'b0), .Q(o_mask[1]) );
  \**FFGEN**  \update_mask_0/o_mask_reg[0]  ( .next_state(1'b0), .clocked_on(
        1'b0), .force_00(1'b0), .force_01(n749), .force_10(
        \update_mask_0/n988 ), .force_11(1'b0), .Q(o_mask[0]) );
  \**FFGEN**  \update_output_0/increment_reg  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2183 ), 
        .force_10(n9182), .force_11(1'b0), .QN(\update_output_0/n1535 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[15][19]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2187 ), 
        .force_10(\update_output_0/n2188 ), .force_11(1'b0), .Q(n5328) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[15][18]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2191 ), 
        .force_10(\update_output_0/n2192 ), .force_11(1'b0), .Q(n5339) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[15][17]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2195 ), 
        .force_10(\update_output_0/n2196 ), .force_11(1'b0), .Q(n5350) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[15][16]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2199 ), 
        .force_10(\update_output_0/n2200 ), .force_11(1'b0), .Q(n5361) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[15][15]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2203 ), 
        .force_10(\update_output_0/n2204 ), .force_11(1'b0), .Q(n5372) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[15][14]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2207 ), 
        .force_10(\update_output_0/n2208 ), .force_11(1'b0), .Q(n5383) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[15][13]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2211 ), 
        .force_10(\update_output_0/n2212 ), .force_11(1'b0), .Q(n5394) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[15][12]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2215 ), 
        .force_10(\update_output_0/n2216 ), .force_11(1'b0), .Q(n5405) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[15][11]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2219 ), 
        .force_10(\update_output_0/n2220 ), .force_11(1'b0), .Q(n5416) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[15][10]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2223 ), 
        .force_10(\update_output_0/n2224 ), .force_11(1'b0), .Q(n5427) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[15][9]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2227 ), 
        .force_10(\update_output_0/n2228 ), .force_11(1'b0), .Q(n5438) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[15][8]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2231 ), 
        .force_10(\update_output_0/n2232 ), .force_11(1'b0), .Q(n5449) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[15][7]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2235 ), 
        .force_10(\update_output_0/n2236 ), .force_11(1'b0), .Q(n5460) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[15][6]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2239 ), 
        .force_10(\update_output_0/n2240 ), .force_11(1'b0), .Q(n5471) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[15][5]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2243 ), 
        .force_10(\update_output_0/n2244 ), .force_11(1'b0), .Q(n5482) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[15][4]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2247 ), 
        .force_10(\update_output_0/n2248 ), .force_11(1'b0), .Q(n5493) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[15][3]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2251 ), 
        .force_10(\update_output_0/n2252 ), .force_11(1'b0), .Q(n5504) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[15][2]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2255 ), 
        .force_10(\update_output_0/n2256 ), .force_11(1'b0), .Q(n5515) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[15][1]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2259 ), 
        .force_10(\update_output_0/n2260 ), .force_11(1'b0), .Q(n5526) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[15][0]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2263 ), 
        .force_10(\update_output_0/n2264 ), .force_11(1'b0), .Q(n5537) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[14][19]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2267 ), 
        .force_10(\update_output_0/n2268 ), .force_11(1'b0), .Q(n5329) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[14][18]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2271 ), 
        .force_10(\update_output_0/n2272 ), .force_11(1'b0), .Q(n5340) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[14][17]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2275 ), 
        .force_10(\update_output_0/n2276 ), .force_11(1'b0), .Q(n5351) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[14][16]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2279 ), 
        .force_10(\update_output_0/n2280 ), .force_11(1'b0), .Q(n5362) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[14][15]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2283 ), 
        .force_10(\update_output_0/n2284 ), .force_11(1'b0), .Q(n5373) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[14][14]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2287 ), 
        .force_10(\update_output_0/n2288 ), .force_11(1'b0), .Q(n5384) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[14][13]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2291 ), 
        .force_10(\update_output_0/n2292 ), .force_11(1'b0), .Q(n5395) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[14][12]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2295 ), 
        .force_10(\update_output_0/n2296 ), .force_11(1'b0), .Q(n5406) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[14][11]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2299 ), 
        .force_10(\update_output_0/n2300 ), .force_11(1'b0), .Q(n5417) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[14][10]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2303 ), 
        .force_10(\update_output_0/n2304 ), .force_11(1'b0), .Q(n5428) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[14][9]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2307 ), 
        .force_10(\update_output_0/n2308 ), .force_11(1'b0), .Q(n5439) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[14][8]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2311 ), 
        .force_10(\update_output_0/n2312 ), .force_11(1'b0), .Q(n5450) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[14][7]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2315 ), 
        .force_10(\update_output_0/n2316 ), .force_11(1'b0), .Q(n5461) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[14][6]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2319 ), 
        .force_10(\update_output_0/n2320 ), .force_11(1'b0), .Q(n5472) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[14][5]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2323 ), 
        .force_10(\update_output_0/n2324 ), .force_11(1'b0), .Q(n5483) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[14][4]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2327 ), 
        .force_10(\update_output_0/n2328 ), .force_11(1'b0), .Q(n5494) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[14][3]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2331 ), 
        .force_10(\update_output_0/n2332 ), .force_11(1'b0), .Q(n5505) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[14][2]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2335 ), 
        .force_10(\update_output_0/n2336 ), .force_11(1'b0), .Q(n5516) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[14][1]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2339 ), 
        .force_10(\update_output_0/n2340 ), .force_11(1'b0), .Q(n5527) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[14][0]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2343 ), 
        .force_10(\update_output_0/n2344 ), .force_11(1'b0), .Q(n5538) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[13][19]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2347 ), 
        .force_10(\update_output_0/n2348 ), .force_11(1'b0), .QN(
        \update_output_0/n6703 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[13][18]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2351 ), 
        .force_10(\update_output_0/n2352 ), .force_11(1'b0), .QN(
        \update_output_0/n6702 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[13][17]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2355 ), 
        .force_10(\update_output_0/n2356 ), .force_11(1'b0), .QN(
        \update_output_0/n6701 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[13][16]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2359 ), 
        .force_10(\update_output_0/n2360 ), .force_11(1'b0), .QN(
        \update_output_0/n6700 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[13][15]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2363 ), 
        .force_10(\update_output_0/n2364 ), .force_11(1'b0), .QN(
        \update_output_0/n6699 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[13][14]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2367 ), 
        .force_10(\update_output_0/n2368 ), .force_11(1'b0), .QN(
        \update_output_0/n6698 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[13][13]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2371 ), 
        .force_10(\update_output_0/n2372 ), .force_11(1'b0), .QN(
        \update_output_0/n6697 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[13][12]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2375 ), 
        .force_10(\update_output_0/n2376 ), .force_11(1'b0), .QN(
        \update_output_0/n6696 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[13][11]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2379 ), 
        .force_10(\update_output_0/n2380 ), .force_11(1'b0), .QN(
        \update_output_0/n6695 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[13][10]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2383 ), 
        .force_10(\update_output_0/n2384 ), .force_11(1'b0), .QN(
        \update_output_0/n6694 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[13][9]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2387 ), 
        .force_10(\update_output_0/n2388 ), .force_11(1'b0), .QN(
        \update_output_0/n6693 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[13][8]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2391 ), 
        .force_10(\update_output_0/n2392 ), .force_11(1'b0), .QN(
        \update_output_0/n6692 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[13][7]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2395 ), 
        .force_10(\update_output_0/n2396 ), .force_11(1'b0), .QN(
        \update_output_0/n6691 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[13][6]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2399 ), 
        .force_10(\update_output_0/n2400 ), .force_11(1'b0), .QN(
        \update_output_0/n6690 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[13][5]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2403 ), 
        .force_10(\update_output_0/n2404 ), .force_11(1'b0), .QN(
        \update_output_0/n6689 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[13][4]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2407 ), 
        .force_10(\update_output_0/n2408 ), .force_11(1'b0), .QN(
        \update_output_0/n6688 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[13][3]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2411 ), 
        .force_10(\update_output_0/n2412 ), .force_11(1'b0), .QN(
        \update_output_0/n6687 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[13][2]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2415 ), 
        .force_10(\update_output_0/n2416 ), .force_11(1'b0), .QN(
        \update_output_0/n6686 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[13][1]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2419 ), 
        .force_10(\update_output_0/n2420 ), .force_11(1'b0), .QN(
        \update_output_0/n6685 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[13][0]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2423 ), 
        .force_10(\update_output_0/n2424 ), .force_11(1'b0), .QN(
        \update_output_0/n6684 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[12][19]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2427 ), 
        .force_10(\update_output_0/n2428 ), .force_11(1'b0), .QN(
        \update_output_0/n6683 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[12][18]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2431 ), 
        .force_10(\update_output_0/n2432 ), .force_11(1'b0), .QN(
        \update_output_0/n6682 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[12][17]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2435 ), 
        .force_10(\update_output_0/n2436 ), .force_11(1'b0), .QN(
        \update_output_0/n6681 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[12][16]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2439 ), 
        .force_10(\update_output_0/n2440 ), .force_11(1'b0), .QN(
        \update_output_0/n6680 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[12][15]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2443 ), 
        .force_10(\update_output_0/n2444 ), .force_11(1'b0), .QN(
        \update_output_0/n6679 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[12][14]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2447 ), 
        .force_10(\update_output_0/n2448 ), .force_11(1'b0), .QN(
        \update_output_0/n6678 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[12][13]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2451 ), 
        .force_10(\update_output_0/n2452 ), .force_11(1'b0), .QN(
        \update_output_0/n6677 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[12][12]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2455 ), 
        .force_10(\update_output_0/n2456 ), .force_11(1'b0), .QN(
        \update_output_0/n6676 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[12][11]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2459 ), 
        .force_10(\update_output_0/n2460 ), .force_11(1'b0), .QN(
        \update_output_0/n6675 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[12][10]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2463 ), 
        .force_10(\update_output_0/n2464 ), .force_11(1'b0), .QN(
        \update_output_0/n6674 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[12][9]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2467 ), 
        .force_10(\update_output_0/n2468 ), .force_11(1'b0), .QN(
        \update_output_0/n6673 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[12][8]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2471 ), 
        .force_10(\update_output_0/n2472 ), .force_11(1'b0), .QN(
        \update_output_0/n6672 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[12][7]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2475 ), 
        .force_10(\update_output_0/n2476 ), .force_11(1'b0), .QN(
        \update_output_0/n6671 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[12][6]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2479 ), 
        .force_10(\update_output_0/n2480 ), .force_11(1'b0), .QN(
        \update_output_0/n6670 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[12][5]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2483 ), 
        .force_10(\update_output_0/n2484 ), .force_11(1'b0), .QN(
        \update_output_0/n6669 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[12][4]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2487 ), 
        .force_10(\update_output_0/n2488 ), .force_11(1'b0), .QN(
        \update_output_0/n6668 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[12][3]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2491 ), 
        .force_10(\update_output_0/n2492 ), .force_11(1'b0), .QN(
        \update_output_0/n6667 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[12][2]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2495 ), 
        .force_10(\update_output_0/n2496 ), .force_11(1'b0), .QN(
        \update_output_0/n6666 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[12][1]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2499 ), 
        .force_10(\update_output_0/n2500 ), .force_11(1'b0), .QN(
        \update_output_0/n6665 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[12][0]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2503 ), 
        .force_10(\update_output_0/n2504 ), .force_11(1'b0), .QN(
        \update_output_0/n6664 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[11][19]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2507 ), 
        .force_10(\update_output_0/n2508 ), .force_11(1'b0), .Q(n5330) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[11][18]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2511 ), 
        .force_10(\update_output_0/n2512 ), .force_11(1'b0), .Q(n5341) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[11][17]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2515 ), 
        .force_10(\update_output_0/n2516 ), .force_11(1'b0), .Q(n5352) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[11][16]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2519 ), 
        .force_10(\update_output_0/n2520 ), .force_11(1'b0), .Q(n5363) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[11][15]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2523 ), 
        .force_10(\update_output_0/n2524 ), .force_11(1'b0), .Q(n5374) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[11][14]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2527 ), 
        .force_10(\update_output_0/n2528 ), .force_11(1'b0), .Q(n5385) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[11][13]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2531 ), 
        .force_10(\update_output_0/n2532 ), .force_11(1'b0), .Q(n5396) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[11][12]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2535 ), 
        .force_10(\update_output_0/n2536 ), .force_11(1'b0), .Q(n5407) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[11][11]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2539 ), 
        .force_10(\update_output_0/n2540 ), .force_11(1'b0), .Q(n5418) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[11][10]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2543 ), 
        .force_10(\update_output_0/n2544 ), .force_11(1'b0), .Q(n5429) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[11][9]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2547 ), 
        .force_10(\update_output_0/n2548 ), .force_11(1'b0), .Q(n5440) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[11][8]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2551 ), 
        .force_10(\update_output_0/n2552 ), .force_11(1'b0), .Q(n5451) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[11][7]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2555 ), 
        .force_10(\update_output_0/n2556 ), .force_11(1'b0), .Q(n5462) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[11][6]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2559 ), 
        .force_10(\update_output_0/n2560 ), .force_11(1'b0), .Q(n5473) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[11][5]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2563 ), 
        .force_10(\update_output_0/n2564 ), .force_11(1'b0), .Q(n5484) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[11][4]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2567 ), 
        .force_10(\update_output_0/n2568 ), .force_11(1'b0), .Q(n5495) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[11][3]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2571 ), 
        .force_10(\update_output_0/n2572 ), .force_11(1'b0), .Q(n5506) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[11][2]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2575 ), 
        .force_10(\update_output_0/n2576 ), .force_11(1'b0), .Q(n5517) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[11][1]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2579 ), 
        .force_10(\update_output_0/n2580 ), .force_11(1'b0), .Q(n5528) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[11][0]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2583 ), 
        .force_10(\update_output_0/n2584 ), .force_11(1'b0), .Q(n5539) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[10][19]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2587 ), 
        .force_10(\update_output_0/n2588 ), .force_11(1'b0), .Q(n5331) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[10][18]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2591 ), 
        .force_10(\update_output_0/n2592 ), .force_11(1'b0), .Q(n5342) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[10][17]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2595 ), 
        .force_10(\update_output_0/n2596 ), .force_11(1'b0), .Q(n5353) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[10][16]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2599 ), 
        .force_10(\update_output_0/n2600 ), .force_11(1'b0), .Q(n5364) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[10][15]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2603 ), 
        .force_10(\update_output_0/n2604 ), .force_11(1'b0), .Q(n5375) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[10][14]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2607 ), 
        .force_10(\update_output_0/n2608 ), .force_11(1'b0), .Q(n5386) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[10][13]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2611 ), 
        .force_10(\update_output_0/n2612 ), .force_11(1'b0), .Q(n5397) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[10][12]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2615 ), 
        .force_10(\update_output_0/n2616 ), .force_11(1'b0), .Q(n5408) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[10][11]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2619 ), 
        .force_10(\update_output_0/n2620 ), .force_11(1'b0), .Q(n5419) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[10][10]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2623 ), 
        .force_10(\update_output_0/n2624 ), .force_11(1'b0), .Q(n5430) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[10][9]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2627 ), 
        .force_10(\update_output_0/n2628 ), .force_11(1'b0), .Q(n5441) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[10][8]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2631 ), 
        .force_10(\update_output_0/n2632 ), .force_11(1'b0), .Q(n5452) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[10][7]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2635 ), 
        .force_10(\update_output_0/n2636 ), .force_11(1'b0), .Q(n5463) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[10][6]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2639 ), 
        .force_10(\update_output_0/n2640 ), .force_11(1'b0), .Q(n5474) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[10][5]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2643 ), 
        .force_10(\update_output_0/n2644 ), .force_11(1'b0), .Q(n5485) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[10][4]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2647 ), 
        .force_10(\update_output_0/n2648 ), .force_11(1'b0), .Q(n5496) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[10][3]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2651 ), 
        .force_10(\update_output_0/n2652 ), .force_11(1'b0), .Q(n5507) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[10][2]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2655 ), 
        .force_10(\update_output_0/n2656 ), .force_11(1'b0), .Q(n5518) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[10][1]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2659 ), 
        .force_10(\update_output_0/n2660 ), .force_11(1'b0), .Q(n5529) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[10][0]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2663 ), 
        .force_10(\update_output_0/n2664 ), .force_11(1'b0), .Q(n5540) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[9][19]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2667 ), 
        .force_10(\update_output_0/n2668 ), .force_11(1'b0), .Q(n5332) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[9][18]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2671 ), 
        .force_10(\update_output_0/n2672 ), .force_11(1'b0), .Q(n5343) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[9][17]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2675 ), 
        .force_10(\update_output_0/n2676 ), .force_11(1'b0), .Q(n5354) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[9][16]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2679 ), 
        .force_10(\update_output_0/n2680 ), .force_11(1'b0), .Q(n5365) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[9][15]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2683 ), 
        .force_10(\update_output_0/n2684 ), .force_11(1'b0), .Q(n5376) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[9][14]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2687 ), 
        .force_10(\update_output_0/n2688 ), .force_11(1'b0), .Q(n5387) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[9][13]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2691 ), 
        .force_10(\update_output_0/n2692 ), .force_11(1'b0), .Q(n5398) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[9][12]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2695 ), 
        .force_10(\update_output_0/n2696 ), .force_11(1'b0), .Q(n5409) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[9][11]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2699 ), 
        .force_10(\update_output_0/n2700 ), .force_11(1'b0), .Q(n5420) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[9][10]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2703 ), 
        .force_10(\update_output_0/n2704 ), .force_11(1'b0), .Q(n5431) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[9][9]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2707 ), 
        .force_10(\update_output_0/n2708 ), .force_11(1'b0), .Q(n5442) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[9][8]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2711 ), 
        .force_10(\update_output_0/n2712 ), .force_11(1'b0), .Q(n5453) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[9][7]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2715 ), 
        .force_10(\update_output_0/n2716 ), .force_11(1'b0), .Q(n5464) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[9][6]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2719 ), 
        .force_10(\update_output_0/n2720 ), .force_11(1'b0), .Q(n5475) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[9][5]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2723 ), 
        .force_10(\update_output_0/n2724 ), .force_11(1'b0), .Q(n5486) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[9][4]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2727 ), 
        .force_10(\update_output_0/n2728 ), .force_11(1'b0), .Q(n5497) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[9][3]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2731 ), 
        .force_10(\update_output_0/n2732 ), .force_11(1'b0), .Q(n5508) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[9][2]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2735 ), 
        .force_10(\update_output_0/n2736 ), .force_11(1'b0), .Q(n5519) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[9][1]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2739 ), 
        .force_10(\update_output_0/n2740 ), .force_11(1'b0), .Q(n5530) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[9][0]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2743 ), 
        .force_10(\update_output_0/n2744 ), .force_11(1'b0), .Q(n5541) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[8][19]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2747 ), 
        .force_10(\update_output_0/n2748 ), .force_11(1'b0), .Q(n5333) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[8][18]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2751 ), 
        .force_10(\update_output_0/n2752 ), .force_11(1'b0), .Q(n5344) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[8][17]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2755 ), 
        .force_10(\update_output_0/n2756 ), .force_11(1'b0), .Q(n5355) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[8][16]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2759 ), 
        .force_10(\update_output_0/n2760 ), .force_11(1'b0), .Q(n5366) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[8][15]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2763 ), 
        .force_10(\update_output_0/n2764 ), .force_11(1'b0), .Q(n5377) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[8][14]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2767 ), 
        .force_10(\update_output_0/n2768 ), .force_11(1'b0), .Q(n5388) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[8][13]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2771 ), 
        .force_10(\update_output_0/n2772 ), .force_11(1'b0), .Q(n5399) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[8][12]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2775 ), 
        .force_10(\update_output_0/n2776 ), .force_11(1'b0), .Q(n5410) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[8][11]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2779 ), 
        .force_10(\update_output_0/n2780 ), .force_11(1'b0), .Q(n5421) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[8][10]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2783 ), 
        .force_10(\update_output_0/n2784 ), .force_11(1'b0), .Q(n5432) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[8][9]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2787 ), 
        .force_10(\update_output_0/n2788 ), .force_11(1'b0), .Q(n5443) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[8][8]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2791 ), 
        .force_10(\update_output_0/n2792 ), .force_11(1'b0), .Q(n5454) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[8][7]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2795 ), 
        .force_10(\update_output_0/n2796 ), .force_11(1'b0), .Q(n5465) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[8][6]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2799 ), 
        .force_10(\update_output_0/n2800 ), .force_11(1'b0), .Q(n5476) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[8][5]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2803 ), 
        .force_10(\update_output_0/n2804 ), .force_11(1'b0), .Q(n5487) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[8][4]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2807 ), 
        .force_10(\update_output_0/n2808 ), .force_11(1'b0), .Q(n5498) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[8][3]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2811 ), 
        .force_10(\update_output_0/n2812 ), .force_11(1'b0), .Q(n5509) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[8][2]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2815 ), 
        .force_10(\update_output_0/n2816 ), .force_11(1'b0), .Q(n5520) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[8][1]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2819 ), 
        .force_10(\update_output_0/n2820 ), .force_11(1'b0), .Q(n5531) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[8][0]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2823 ), 
        .force_10(\update_output_0/n2824 ), .force_11(1'b0), .Q(n5542) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[7][19]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2827 ), 
        .force_10(\update_output_0/n2828 ), .force_11(1'b0), .QN(
        \update_output_0/n6583 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[7][18]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2831 ), 
        .force_10(\update_output_0/n2832 ), .force_11(1'b0), .QN(
        \update_output_0/n6582 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[7][17]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2835 ), 
        .force_10(\update_output_0/n2836 ), .force_11(1'b0), .QN(
        \update_output_0/n6581 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[7][16]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2839 ), 
        .force_10(\update_output_0/n2840 ), .force_11(1'b0), .QN(
        \update_output_0/n6580 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[7][15]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2843 ), 
        .force_10(\update_output_0/n2844 ), .force_11(1'b0), .QN(
        \update_output_0/n6579 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[7][14]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2847 ), 
        .force_10(\update_output_0/n2848 ), .force_11(1'b0), .QN(
        \update_output_0/n6578 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[7][13]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2851 ), 
        .force_10(\update_output_0/n2852 ), .force_11(1'b0), .QN(
        \update_output_0/n6577 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[7][12]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2855 ), 
        .force_10(\update_output_0/n2856 ), .force_11(1'b0), .QN(
        \update_output_0/n6576 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[7][11]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2859 ), 
        .force_10(\update_output_0/n2860 ), .force_11(1'b0), .QN(
        \update_output_0/n6575 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[7][10]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2863 ), 
        .force_10(\update_output_0/n2864 ), .force_11(1'b0), .QN(
        \update_output_0/n6574 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[7][9]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2867 ), 
        .force_10(\update_output_0/n2868 ), .force_11(1'b0), .QN(
        \update_output_0/n6573 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[7][8]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2871 ), 
        .force_10(\update_output_0/n2872 ), .force_11(1'b0), .QN(
        \update_output_0/n6572 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[7][7]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2875 ), 
        .force_10(\update_output_0/n2876 ), .force_11(1'b0), .QN(
        \update_output_0/n6571 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[7][6]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2879 ), 
        .force_10(\update_output_0/n2880 ), .force_11(1'b0), .QN(
        \update_output_0/n6570 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[7][5]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2883 ), 
        .force_10(\update_output_0/n2884 ), .force_11(1'b0), .QN(
        \update_output_0/n6569 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[7][4]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2887 ), 
        .force_10(\update_output_0/n2888 ), .force_11(1'b0), .QN(
        \update_output_0/n6568 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[7][3]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2891 ), 
        .force_10(\update_output_0/n2892 ), .force_11(1'b0), .QN(
        \update_output_0/n6567 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[7][2]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2895 ), 
        .force_10(\update_output_0/n2896 ), .force_11(1'b0), .QN(
        \update_output_0/n6566 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[7][1]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2899 ), 
        .force_10(\update_output_0/n2900 ), .force_11(1'b0), .QN(
        \update_output_0/n6565 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[7][0]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2903 ), 
        .force_10(\update_output_0/n2904 ), .force_11(1'b0), .QN(
        \update_output_0/n6564 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[6][19]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2907 ), 
        .force_10(\update_output_0/n2908 ), .force_11(1'b0), .QN(
        \update_output_0/n6563 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[6][18]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2911 ), 
        .force_10(\update_output_0/n2912 ), .force_11(1'b0), .QN(
        \update_output_0/n6562 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[6][17]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2915 ), 
        .force_10(\update_output_0/n2916 ), .force_11(1'b0), .QN(
        \update_output_0/n6561 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[6][16]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2919 ), 
        .force_10(\update_output_0/n2920 ), .force_11(1'b0), .QN(
        \update_output_0/n6560 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[6][15]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2923 ), 
        .force_10(\update_output_0/n2924 ), .force_11(1'b0), .QN(
        \update_output_0/n6559 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[6][14]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2927 ), 
        .force_10(\update_output_0/n2928 ), .force_11(1'b0), .QN(
        \update_output_0/n6558 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[6][13]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2931 ), 
        .force_10(\update_output_0/n2932 ), .force_11(1'b0), .QN(
        \update_output_0/n6557 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[6][12]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2935 ), 
        .force_10(\update_output_0/n2936 ), .force_11(1'b0), .QN(
        \update_output_0/n6556 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[6][11]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2939 ), 
        .force_10(\update_output_0/n2940 ), .force_11(1'b0), .QN(
        \update_output_0/n6555 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[6][10]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2943 ), 
        .force_10(\update_output_0/n2944 ), .force_11(1'b0), .QN(
        \update_output_0/n6554 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[6][9]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2947 ), 
        .force_10(\update_output_0/n2948 ), .force_11(1'b0), .QN(
        \update_output_0/n6553 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[6][8]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2951 ), 
        .force_10(\update_output_0/n2952 ), .force_11(1'b0), .QN(
        \update_output_0/n6552 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[6][7]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2955 ), 
        .force_10(\update_output_0/n2956 ), .force_11(1'b0), .QN(
        \update_output_0/n6551 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[6][6]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2959 ), 
        .force_10(\update_output_0/n2960 ), .force_11(1'b0), .QN(
        \update_output_0/n6550 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[6][5]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2963 ), 
        .force_10(\update_output_0/n2964 ), .force_11(1'b0), .QN(
        \update_output_0/n6549 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[6][4]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2967 ), 
        .force_10(\update_output_0/n2968 ), .force_11(1'b0), .QN(
        \update_output_0/n6548 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[6][3]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2971 ), 
        .force_10(\update_output_0/n2972 ), .force_11(1'b0), .QN(
        \update_output_0/n6547 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[6][2]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2975 ), 
        .force_10(\update_output_0/n2976 ), .force_11(1'b0), .QN(
        \update_output_0/n6546 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[6][1]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2979 ), 
        .force_10(\update_output_0/n2980 ), .force_11(1'b0), .QN(
        \update_output_0/n6545 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[6][0]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2983 ), 
        .force_10(\update_output_0/n2984 ), .force_11(1'b0), .QN(
        \update_output_0/n6544 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[5][19]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2987 ), 
        .force_10(\update_output_0/n2988 ), .force_11(1'b0), .Q(n5334) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[5][18]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2991 ), 
        .force_10(\update_output_0/n2992 ), .force_11(1'b0), .Q(n5345) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[5][17]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2995 ), 
        .force_10(\update_output_0/n2996 ), .force_11(1'b0), .Q(n5356) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[5][16]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2999 ), 
        .force_10(\update_output_0/n3000 ), .force_11(1'b0), .Q(n5367) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[5][15]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3003 ), 
        .force_10(\update_output_0/n3004 ), .force_11(1'b0), .Q(n5378) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[5][14]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3007 ), 
        .force_10(\update_output_0/n3008 ), .force_11(1'b0), .Q(n5389) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[5][13]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3011 ), 
        .force_10(\update_output_0/n3012 ), .force_11(1'b0), .Q(n5400) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[5][12]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3015 ), 
        .force_10(\update_output_0/n3016 ), .force_11(1'b0), .Q(n5411) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[5][11]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3019 ), 
        .force_10(\update_output_0/n3020 ), .force_11(1'b0), .Q(n5422) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[5][10]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3023 ), 
        .force_10(\update_output_0/n3024 ), .force_11(1'b0), .Q(n5433) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[5][9]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3027 ), 
        .force_10(\update_output_0/n3028 ), .force_11(1'b0), .Q(n5444) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[5][8]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3031 ), 
        .force_10(\update_output_0/n3032 ), .force_11(1'b0), .Q(n5455) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[5][7]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3035 ), 
        .force_10(\update_output_0/n3036 ), .force_11(1'b0), .Q(n5466) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[5][6]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3039 ), 
        .force_10(\update_output_0/n3040 ), .force_11(1'b0), .Q(n5477) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[5][5]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3043 ), 
        .force_10(\update_output_0/n3044 ), .force_11(1'b0), .Q(n5488) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[5][4]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3047 ), 
        .force_10(\update_output_0/n3048 ), .force_11(1'b0), .Q(n5499) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[5][3]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3051 ), 
        .force_10(\update_output_0/n3052 ), .force_11(1'b0), .Q(n5510) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[5][2]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3055 ), 
        .force_10(\update_output_0/n3056 ), .force_11(1'b0), .Q(n5521) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[5][1]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3059 ), 
        .force_10(\update_output_0/n3060 ), .force_11(1'b0), .Q(n5532) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[5][0]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3063 ), 
        .force_10(\update_output_0/n3064 ), .force_11(1'b0), .Q(n5543) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[4][19]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3067 ), 
        .force_10(\update_output_0/n3068 ), .force_11(1'b0), .Q(n5335) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[4][18]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3071 ), 
        .force_10(\update_output_0/n3072 ), .force_11(1'b0), .Q(n5346) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[4][17]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3075 ), 
        .force_10(\update_output_0/n3076 ), .force_11(1'b0), .Q(n5357) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[4][16]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3079 ), 
        .force_10(\update_output_0/n3080 ), .force_11(1'b0), .Q(n5368) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[4][15]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3083 ), 
        .force_10(\update_output_0/n3084 ), .force_11(1'b0), .Q(n5379) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[4][14]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3087 ), 
        .force_10(\update_output_0/n3088 ), .force_11(1'b0), .Q(n5390) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[4][13]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3091 ), 
        .force_10(\update_output_0/n3092 ), .force_11(1'b0), .Q(n5401) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[4][12]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3095 ), 
        .force_10(\update_output_0/n3096 ), .force_11(1'b0), .Q(n5412) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[4][11]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3099 ), 
        .force_10(\update_output_0/n3100 ), .force_11(1'b0), .Q(n5423) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[4][10]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3103 ), 
        .force_10(\update_output_0/n3104 ), .force_11(1'b0), .Q(n5434) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[4][9]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3107 ), 
        .force_10(\update_output_0/n3108 ), .force_11(1'b0), .Q(n5445) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[4][8]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3111 ), 
        .force_10(\update_output_0/n3112 ), .force_11(1'b0), .Q(n5456) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[4][7]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3115 ), 
        .force_10(\update_output_0/n3116 ), .force_11(1'b0), .Q(n5467) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[4][6]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3119 ), 
        .force_10(\update_output_0/n3120 ), .force_11(1'b0), .Q(n5478) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[4][5]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3123 ), 
        .force_10(\update_output_0/n3124 ), .force_11(1'b0), .Q(n5489) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[4][4]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3127 ), 
        .force_10(\update_output_0/n3128 ), .force_11(1'b0), .Q(n5500) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[4][3]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3131 ), 
        .force_10(\update_output_0/n3132 ), .force_11(1'b0), .Q(n5511) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[4][2]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3135 ), 
        .force_10(\update_output_0/n3136 ), .force_11(1'b0), .Q(n5522) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[4][1]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3139 ), 
        .force_10(\update_output_0/n3140 ), .force_11(1'b0), .Q(n5533) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[4][0]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3143 ), 
        .force_10(\update_output_0/n3144 ), .force_11(1'b0), .Q(n5544) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[3][19]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3147 ), 
        .force_10(\update_output_0/n3148 ), .force_11(1'b0), .Q(n5336) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[3][18]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3151 ), 
        .force_10(\update_output_0/n3152 ), .force_11(1'b0), .Q(n5347) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[3][17]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3155 ), 
        .force_10(\update_output_0/n3156 ), .force_11(1'b0), .Q(n5358) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[3][16]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3159 ), 
        .force_10(\update_output_0/n3160 ), .force_11(1'b0), .Q(n5369) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[3][15]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3163 ), 
        .force_10(\update_output_0/n3164 ), .force_11(1'b0), .Q(n5380) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[3][14]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3167 ), 
        .force_10(\update_output_0/n3168 ), .force_11(1'b0), .Q(n5391) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[3][13]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3171 ), 
        .force_10(\update_output_0/n3172 ), .force_11(1'b0), .Q(n5402) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[3][12]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3175 ), 
        .force_10(\update_output_0/n3176 ), .force_11(1'b0), .Q(n5413) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[3][11]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3179 ), 
        .force_10(\update_output_0/n3180 ), .force_11(1'b0), .Q(n5424) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[3][10]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3183 ), 
        .force_10(\update_output_0/n3184 ), .force_11(1'b0), .Q(n5435) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[3][9]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3187 ), 
        .force_10(\update_output_0/n3188 ), .force_11(1'b0), .Q(n5446) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[3][8]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3191 ), 
        .force_10(\update_output_0/n3192 ), .force_11(1'b0), .Q(n5457) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[3][7]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3195 ), 
        .force_10(\update_output_0/n3196 ), .force_11(1'b0), .Q(n5468) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[3][6]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3199 ), 
        .force_10(\update_output_0/n3200 ), .force_11(1'b0), .Q(n5479) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[3][5]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3203 ), 
        .force_10(\update_output_0/n3204 ), .force_11(1'b0), .Q(n5490) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[3][4]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3207 ), 
        .force_10(\update_output_0/n3208 ), .force_11(1'b0), .Q(n5501) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[3][3]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3211 ), 
        .force_10(\update_output_0/n3212 ), .force_11(1'b0), .Q(n5512) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[3][2]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3215 ), 
        .force_10(\update_output_0/n3216 ), .force_11(1'b0), .Q(n5523) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[3][1]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3219 ), 
        .force_10(\update_output_0/n3220 ), .force_11(1'b0), .Q(n5534) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[3][0]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3223 ), 
        .force_10(\update_output_0/n3224 ), .force_11(1'b0), .Q(n5545) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[2][19]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3227 ), 
        .force_10(\update_output_0/n3228 ), .force_11(1'b0), .Q(n5337) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[2][18]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3231 ), 
        .force_10(\update_output_0/n3232 ), .force_11(1'b0), .Q(n5348) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[2][17]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3235 ), 
        .force_10(\update_output_0/n3236 ), .force_11(1'b0), .Q(n5359) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[2][16]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3239 ), 
        .force_10(\update_output_0/n3240 ), .force_11(1'b0), .Q(n5370) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[2][15]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3243 ), 
        .force_10(\update_output_0/n3244 ), .force_11(1'b0), .Q(n5381) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[2][14]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3247 ), 
        .force_10(\update_output_0/n3248 ), .force_11(1'b0), .Q(n5392) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[2][13]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3251 ), 
        .force_10(\update_output_0/n3252 ), .force_11(1'b0), .Q(n5403) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[2][12]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3255 ), 
        .force_10(\update_output_0/n3256 ), .force_11(1'b0), .Q(n5414) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[2][11]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3259 ), 
        .force_10(\update_output_0/n3260 ), .force_11(1'b0), .Q(n5425) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[2][10]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3263 ), 
        .force_10(\update_output_0/n3264 ), .force_11(1'b0), .Q(n5436) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[2][9]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3267 ), 
        .force_10(\update_output_0/n3268 ), .force_11(1'b0), .Q(n5447) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[2][8]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3271 ), 
        .force_10(\update_output_0/n3272 ), .force_11(1'b0), .Q(n5458) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[2][7]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3275 ), 
        .force_10(\update_output_0/n3276 ), .force_11(1'b0), .Q(n5469) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[2][6]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3279 ), 
        .force_10(\update_output_0/n3280 ), .force_11(1'b0), .Q(n5480) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[2][5]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3283 ), 
        .force_10(\update_output_0/n3284 ), .force_11(1'b0), .Q(n5491) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[2][4]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3287 ), 
        .force_10(\update_output_0/n3288 ), .force_11(1'b0), .Q(n5502) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[2][3]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3291 ), 
        .force_10(\update_output_0/n3292 ), .force_11(1'b0), .Q(n5513) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[2][2]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3295 ), 
        .force_10(\update_output_0/n3296 ), .force_11(1'b0), .Q(n5524) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[2][1]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3299 ), 
        .force_10(\update_output_0/n3300 ), .force_11(1'b0), .Q(n5535) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[2][0]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3303 ), 
        .force_10(\update_output_0/n3304 ), .force_11(1'b0), .Q(n5546) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[1][19]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3307 ), 
        .force_10(\update_output_0/n3308 ), .force_11(1'b0), .Q(n5338) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[1][18]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3311 ), 
        .force_10(\update_output_0/n3312 ), .force_11(1'b0), .Q(n5349) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[1][17]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3315 ), 
        .force_10(\update_output_0/n3316 ), .force_11(1'b0), .Q(n5360) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[1][16]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3319 ), 
        .force_10(\update_output_0/n3320 ), .force_11(1'b0), .Q(n5371) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[1][15]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3323 ), 
        .force_10(\update_output_0/n3324 ), .force_11(1'b0), .Q(n5382) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[1][14]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3327 ), 
        .force_10(\update_output_0/n3328 ), .force_11(1'b0), .Q(n5393) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[1][13]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3331 ), 
        .force_10(\update_output_0/n3332 ), .force_11(1'b0), .Q(n5404) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[1][12]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3335 ), 
        .force_10(\update_output_0/n3336 ), .force_11(1'b0), .Q(n5415) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[1][11]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3339 ), 
        .force_10(\update_output_0/n3340 ), .force_11(1'b0), .Q(n5426) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[1][10]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3343 ), 
        .force_10(\update_output_0/n3344 ), .force_11(1'b0), .Q(n5437) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[1][9]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3347 ), 
        .force_10(\update_output_0/n3348 ), .force_11(1'b0), .Q(n5448) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[1][8]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3351 ), 
        .force_10(\update_output_0/n3352 ), .force_11(1'b0), .Q(n5459) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[1][7]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3355 ), 
        .force_10(\update_output_0/n3356 ), .force_11(1'b0), .Q(n5470) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[1][6]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3359 ), 
        .force_10(\update_output_0/n3360 ), .force_11(1'b0), .Q(n5481) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[1][5]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3363 ), 
        .force_10(\update_output_0/n3364 ), .force_11(1'b0), .Q(n5492) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[1][4]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3367 ), 
        .force_10(\update_output_0/n3368 ), .force_11(1'b0), .Q(n5503) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[1][3]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3371 ), 
        .force_10(\update_output_0/n3372 ), .force_11(1'b0), .Q(n5514) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[1][2]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3375 ), 
        .force_10(\update_output_0/n3376 ), .force_11(1'b0), .Q(n5525) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[1][1]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3379 ), 
        .force_10(\update_output_0/n3380 ), .force_11(1'b0), .Q(n5536) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[1][0]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3383 ), 
        .force_10(\update_output_0/n3384 ), .force_11(1'b0), .Q(n5547) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[0][19]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3387 ), 
        .force_10(\update_output_0/n3388 ), .force_11(1'b0), .QN(
        \update_output_0/n6443 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[0][18]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3391 ), 
        .force_10(\update_output_0/n3392 ), .force_11(1'b0), .QN(
        \update_output_0/n6442 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[0][17]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3395 ), 
        .force_10(\update_output_0/n3396 ), .force_11(1'b0), .QN(
        \update_output_0/n6441 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[0][16]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3399 ), 
        .force_10(\update_output_0/n3400 ), .force_11(1'b0), .QN(
        \update_output_0/n6440 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[0][15]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3403 ), 
        .force_10(\update_output_0/n3404 ), .force_11(1'b0), .QN(
        \update_output_0/n6439 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[0][14]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3407 ), 
        .force_10(\update_output_0/n3408 ), .force_11(1'b0), .QN(
        \update_output_0/n6438 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[0][13]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3411 ), 
        .force_10(\update_output_0/n3412 ), .force_11(1'b0), .QN(
        \update_output_0/n6437 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[0][12]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3415 ), 
        .force_10(\update_output_0/n3416 ), .force_11(1'b0), .QN(
        \update_output_0/n6436 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[0][11]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3419 ), 
        .force_10(\update_output_0/n3420 ), .force_11(1'b0), .QN(
        \update_output_0/n6435 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[0][10]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3423 ), 
        .force_10(\update_output_0/n3424 ), .force_11(1'b0), .QN(
        \update_output_0/n6434 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[0][9]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3427 ), 
        .force_10(\update_output_0/n3428 ), .force_11(1'b0), .QN(
        \update_output_0/n6433 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[0][8]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3431 ), 
        .force_10(\update_output_0/n3432 ), .force_11(1'b0), .QN(
        \update_output_0/n6432 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[0][7]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3435 ), 
        .force_10(\update_output_0/n3436 ), .force_11(1'b0), .QN(
        \update_output_0/n6431 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[0][6]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3439 ), 
        .force_10(\update_output_0/n3440 ), .force_11(1'b0), .QN(
        \update_output_0/n6430 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[0][5]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3443 ), 
        .force_10(\update_output_0/n3444 ), .force_11(1'b0), .QN(
        \update_output_0/n6429 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[0][4]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3447 ), 
        .force_10(\update_output_0/n3448 ), .force_11(1'b0), .QN(
        \update_output_0/n6428 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[0][3]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3451 ), 
        .force_10(\update_output_0/n3452 ), .force_11(1'b0), .QN(
        \update_output_0/n6427 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[0][2]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3455 ), 
        .force_10(\update_output_0/n3456 ), .force_11(1'b0), .QN(
        \update_output_0/n6426 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[0][1]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n3459 ), 
        .force_10(\update_output_0/n3460 ), .force_11(1'b0), .QN(
        \update_output_0/n6425 ) );
  \**FFGEN**  \update_output_0/pre_o_im_reg[0][0]  ( .next_state(1'b0), 
        .clocked_on(1'b0), .force_00(1'b0), .force_01(\update_output_0/n2179 ), 
        .force_10(\update_output_0/n2180 ), .force_11(1'b0), .QN(
        \update_output_0/n6424 ) );
  nand_x8_sg U2963 ( .A(n7564), .B(n7561), .X(n4192) );
  nand_x8_sg U2956 ( .A(n6152), .B(n7569), .X(n4184) );
  nand_x8_sg U2955 ( .A(n7564), .B(n7563), .X(n4196) );
  nor_x2_sg U2167 ( .A(n883), .B(n7568), .X(n882) );
  nor_x2_sg U2166 ( .A(n884), .B(n885), .X(n883) );
  nor_x2_sg U2165 ( .A(n888), .B(n9082), .X(n884) );
  nor_x2_sg U2164 ( .A(\i_im[1][0] ), .B(n7560), .X(n888) );
  nor_x2_sg U2161 ( .A(\i_im[0][0] ), .B(n7561), .X(n890) );
  nor_x2_sg U2156 ( .A(n7391), .B(n9102), .X(n875) );
  nand_x8_sg U2932 ( .A(n7392), .B(n7568), .X(n881) );
  nor_x2_sg U2147 ( .A(n7383), .B(n9142), .X(n863) );
  nand_x8_sg U2915 ( .A(n1511), .B(n1512), .X(n866) );
  nor_x2_sg U2145 ( .A(n7381), .B(n9162), .X(n864) );
  nand_x8_sg U2912 ( .A(n1510), .B(n1511), .X(n865) );
  nand_x8_sg U1478 ( .A(n809), .B(n3096), .X(n772) );
  nand_x8_sg U1772 ( .A(n7375), .B(n824), .X(n3098) );
  nand_x8_sg U2972 ( .A(n845), .B(n846), .X(n824) );
  nor_x2_sg U2971 ( .A(n1195), .B(n1196), .X(n845) );
  nor_x2_sg U2946 ( .A(n1525), .B(n7568), .X(n1524) );
  nor_x2_sg U2945 ( .A(n1526), .B(n1527), .X(n1525) );
  nor_x2_sg U2944 ( .A(n1530), .B(n9101), .X(n1526) );
  nor_x2_sg U2943 ( .A(\i_im[1][19] ), .B(n7560), .X(n1530) );
  nor_x2_sg U2940 ( .A(\i_im[0][19] ), .B(n7562), .X(n1532) );
  nor_x2_sg U2933 ( .A(n7390), .B(n9121), .X(n1520) );
  nor_x2_sg U2916 ( .A(n7382), .B(n9161), .X(n1508) );
  nor_x2_sg U2913 ( .A(n7380), .B(n9181), .X(n1509) );
  nor_x2_sg U2892 ( .A(n1489), .B(n7568), .X(n1488) );
  nor_x2_sg U2891 ( .A(n1490), .B(n1491), .X(n1489) );
  nor_x2_sg U2890 ( .A(n1494), .B(n9100), .X(n1490) );
  nor_x2_sg U2889 ( .A(\i_im[1][18] ), .B(n7560), .X(n1494) );
  nor_x2_sg U2886 ( .A(\i_im[0][18] ), .B(n7562), .X(n1496) );
  nor_x2_sg U2881 ( .A(n7391), .B(n9120), .X(n1484) );
  nor_x2_sg U2872 ( .A(n7383), .B(n9160), .X(n1475) );
  nor_x2_sg U2870 ( .A(n7381), .B(n9180), .X(n1476) );
  nor_x2_sg U2852 ( .A(n1456), .B(n7568), .X(n1455) );
  nor_x2_sg U2851 ( .A(n1457), .B(n1458), .X(n1456) );
  nor_x2_sg U2850 ( .A(n1461), .B(n9099), .X(n1457) );
  nor_x2_sg U2849 ( .A(\i_im[1][17] ), .B(n7563), .X(n1461) );
  nor_x2_sg U2846 ( .A(\i_im[0][17] ), .B(n7562), .X(n1463) );
  nor_x2_sg U2841 ( .A(n881), .B(n9119), .X(n1451) );
  nor_x2_sg U2832 ( .A(n866), .B(n9159), .X(n1442) );
  nor_x2_sg U2830 ( .A(n865), .B(n9179), .X(n1443) );
  nor_x2_sg U2811 ( .A(n1423), .B(n7568), .X(n1422) );
  nor_x2_sg U2810 ( .A(n1424), .B(n1425), .X(n1423) );
  nor_x2_sg U2809 ( .A(n1428), .B(n9098), .X(n1424) );
  nor_x2_sg U2808 ( .A(\i_im[1][16] ), .B(n7563), .X(n1428) );
  nor_x2_sg U2805 ( .A(\i_im[0][16] ), .B(n7562), .X(n1430) );
  nor_x2_sg U2800 ( .A(n7390), .B(n9118), .X(n1418) );
  nor_x2_sg U2791 ( .A(n7382), .B(n9158), .X(n1409) );
  nor_x2_sg U2789 ( .A(n7380), .B(n9178), .X(n1410) );
  nor_x2_sg U2771 ( .A(n1390), .B(n7568), .X(n1389) );
  nor_x2_sg U2770 ( .A(n1391), .B(n1392), .X(n1390) );
  nor_x2_sg U2769 ( .A(n1395), .B(n9097), .X(n1391) );
  nor_x2_sg U2768 ( .A(\i_im[1][15] ), .B(n7563), .X(n1395) );
  nor_x2_sg U2765 ( .A(\i_im[0][15] ), .B(n7562), .X(n1397) );
  nor_x2_sg U2760 ( .A(n7391), .B(n9117), .X(n1385) );
  nor_x2_sg U2751 ( .A(n7383), .B(n9157), .X(n1376) );
  nor_x2_sg U2749 ( .A(n7381), .B(n9177), .X(n1377) );
  nor_x2_sg U2730 ( .A(n1354), .B(n7568), .X(n1353) );
  nor_x2_sg U2729 ( .A(n1355), .B(n1356), .X(n1354) );
  nor_x2_sg U2728 ( .A(n1359), .B(n9096), .X(n1355) );
  nor_x2_sg U2727 ( .A(\i_im[1][14] ), .B(n7563), .X(n1359) );
  nor_x2_sg U2724 ( .A(\i_im[0][14] ), .B(n7562), .X(n1361) );
  nor_x2_sg U2719 ( .A(n881), .B(n9116), .X(n1349) );
  nor_x2_sg U2710 ( .A(n866), .B(n9156), .X(n1340) );
  nor_x2_sg U2708 ( .A(n865), .B(n9176), .X(n1341) );
  nor_x2_sg U2691 ( .A(n1321), .B(n7568), .X(n1320) );
  nor_x2_sg U2690 ( .A(n1322), .B(n1323), .X(n1321) );
  nor_x2_sg U2689 ( .A(n1326), .B(n9095), .X(n1322) );
  nor_x2_sg U2688 ( .A(\i_im[1][13] ), .B(n7560), .X(n1326) );
  nor_x2_sg U2685 ( .A(\i_im[0][13] ), .B(n7562), .X(n1328) );
  nor_x2_sg U2680 ( .A(n7390), .B(n9115), .X(n1316) );
  nor_x2_sg U2671 ( .A(n7382), .B(n9155), .X(n1307) );
  nor_x2_sg U2669 ( .A(n7380), .B(n9175), .X(n1308) );
  nor_x2_sg U2651 ( .A(n1288), .B(n7568), .X(n1287) );
  nor_x2_sg U2650 ( .A(n1289), .B(n1290), .X(n1288) );
  nor_x2_sg U2649 ( .A(n1293), .B(n9094), .X(n1289) );
  nor_x2_sg U2648 ( .A(\i_im[1][12] ), .B(n7563), .X(n1293) );
  nor_x2_sg U2645 ( .A(\i_im[0][12] ), .B(n7562), .X(n1295) );
  nor_x2_sg U2640 ( .A(n7391), .B(n9114), .X(n1283) );
  nor_x2_sg U2631 ( .A(n7383), .B(n9154), .X(n1274) );
  nor_x2_sg U2629 ( .A(n7381), .B(n9174), .X(n1275) );
  nor_x2_sg U2610 ( .A(n1255), .B(n7568), .X(n1254) );
  nor_x2_sg U2609 ( .A(n1256), .B(n1257), .X(n1255) );
  nor_x2_sg U2608 ( .A(n1260), .B(n9093), .X(n1256) );
  nor_x2_sg U2607 ( .A(\i_im[1][11] ), .B(n7563), .X(n1260) );
  nor_x2_sg U2604 ( .A(\i_im[0][11] ), .B(n7561), .X(n1262) );
  nor_x2_sg U2599 ( .A(n881), .B(n9113), .X(n1250) );
  nor_x2_sg U2590 ( .A(n866), .B(n9153), .X(n1241) );
  nor_x2_sg U2588 ( .A(n865), .B(n9173), .X(n1242) );
  nor_x2_sg U2570 ( .A(n1222), .B(n7568), .X(n1221) );
  nor_x2_sg U2569 ( .A(n1223), .B(n1224), .X(n1222) );
  nor_x2_sg U2568 ( .A(n1227), .B(n9092), .X(n1223) );
  nor_x2_sg U2567 ( .A(\i_im[1][10] ), .B(n7563), .X(n1227) );
  nor_x2_sg U2564 ( .A(\i_im[0][10] ), .B(n7561), .X(n1229) );
  nor_x2_sg U2559 ( .A(n7390), .B(n9112), .X(n1217) );
  nor_x2_sg U2550 ( .A(n7382), .B(n9152), .X(n1208) );
  nor_x2_sg U2548 ( .A(n7380), .B(n9172), .X(n1209) );
  nor_x2_sg U2542 ( .A(n847), .B(n848), .X(n846) );
  nor_x2_sg U2528 ( .A(n1184), .B(n7568), .X(n1183) );
  nor_x2_sg U2527 ( .A(n1185), .B(n1186), .X(n1184) );
  nor_x2_sg U2526 ( .A(n1189), .B(n9091), .X(n1185) );
  nor_x2_sg U2525 ( .A(\i_im[1][9] ), .B(n7563), .X(n1189) );
  nor_x2_sg U2522 ( .A(\i_im[0][9] ), .B(n7561), .X(n1191) );
  nor_x2_sg U2517 ( .A(n7391), .B(n9111), .X(n1179) );
  nor_x2_sg U2508 ( .A(n7383), .B(n9151), .X(n1170) );
  nor_x2_sg U2506 ( .A(n7381), .B(n9171), .X(n1171) );
  nor_x2_sg U2489 ( .A(n1151), .B(n7568), .X(n1150) );
  nor_x2_sg U2488 ( .A(n1152), .B(n1153), .X(n1151) );
  nor_x2_sg U2487 ( .A(n1156), .B(n9090), .X(n1152) );
  nor_x2_sg U2486 ( .A(\i_im[1][8] ), .B(n7560), .X(n1156) );
  nor_x2_sg U2483 ( .A(\i_im[0][8] ), .B(n7562), .X(n1158) );
  nor_x2_sg U2478 ( .A(n881), .B(n9110), .X(n1146) );
  nor_x2_sg U2469 ( .A(n866), .B(n9150), .X(n1137) );
  nor_x2_sg U2467 ( .A(n865), .B(n9170), .X(n1138) );
  nor_x2_sg U2449 ( .A(n1118), .B(n7568), .X(n1117) );
  nor_x2_sg U2448 ( .A(n1119), .B(n1120), .X(n1118) );
  nor_x2_sg U2447 ( .A(n1123), .B(n9089), .X(n1119) );
  nor_x2_sg U2446 ( .A(\i_im[1][7] ), .B(n7560), .X(n1123) );
  nor_x2_sg U2443 ( .A(\i_im[0][7] ), .B(n7562), .X(n1125) );
  nor_x2_sg U2438 ( .A(n7390), .B(n9109), .X(n1113) );
  nor_x2_sg U2429 ( .A(n7382), .B(n9149), .X(n1104) );
  nor_x2_sg U2427 ( .A(n7380), .B(n9169), .X(n1105) );
  nor_x2_sg U2408 ( .A(n1085), .B(n7568), .X(n1084) );
  nor_x2_sg U2407 ( .A(n1086), .B(n1087), .X(n1085) );
  nor_x2_sg U2406 ( .A(n1090), .B(n9088), .X(n1086) );
  nor_x2_sg U2405 ( .A(\i_im[1][6] ), .B(n7560), .X(n1090) );
  nor_x2_sg U2402 ( .A(\i_im[0][6] ), .B(n7562), .X(n1092) );
  nor_x2_sg U2397 ( .A(n7391), .B(n9108), .X(n1080) );
  nor_x2_sg U2388 ( .A(n7383), .B(n9148), .X(n1071) );
  nor_x2_sg U2386 ( .A(n7381), .B(n9168), .X(n1072) );
  nor_x2_sg U2368 ( .A(n1052), .B(n7568), .X(n1051) );
  nor_x2_sg U2367 ( .A(n1053), .B(n1054), .X(n1052) );
  nor_x2_sg U2366 ( .A(n1057), .B(n9087), .X(n1053) );
  nor_x2_sg U2365 ( .A(\i_im[1][5] ), .B(n7560), .X(n1057) );
  nor_x2_sg U2362 ( .A(\i_im[0][5] ), .B(n7561), .X(n1059) );
  nor_x2_sg U2357 ( .A(n881), .B(n9107), .X(n1047) );
  nor_x2_sg U2348 ( .A(n866), .B(n9147), .X(n1038) );
  nor_x2_sg U2346 ( .A(n865), .B(n9167), .X(n1039) );
  nor_x2_sg U2327 ( .A(n1016), .B(n7568), .X(n1015) );
  nor_x2_sg U2326 ( .A(n1017), .B(n1018), .X(n1016) );
  nor_x2_sg U2325 ( .A(n1021), .B(n9086), .X(n1017) );
  nor_x2_sg U2324 ( .A(\i_im[1][4] ), .B(n7560), .X(n1021) );
  nor_x2_sg U2321 ( .A(\i_im[0][4] ), .B(n7562), .X(n1023) );
  nor_x2_sg U2316 ( .A(n7390), .B(n9106), .X(n1011) );
  nor_x2_sg U2307 ( .A(n7382), .B(n9146), .X(n1002) );
  nor_x2_sg U2305 ( .A(n7380), .B(n9166), .X(n1003) );
  nor_x2_sg U2288 ( .A(n983), .B(n7568), .X(n982) );
  nor_x2_sg U2287 ( .A(n984), .B(n985), .X(n983) );
  nor_x2_sg U2286 ( .A(n988), .B(n9085), .X(n984) );
  nor_x2_sg U2285 ( .A(\i_im[1][3] ), .B(n7560), .X(n988) );
  nor_x2_sg U2282 ( .A(\i_im[0][3] ), .B(n7561), .X(n990) );
  nor_x2_sg U2277 ( .A(n7391), .B(n9105), .X(n978) );
  nor_x2_sg U2268 ( .A(n7383), .B(n9145), .X(n969) );
  nor_x2_sg U2266 ( .A(n7381), .B(n9165), .X(n970) );
  nor_x2_sg U2248 ( .A(n950), .B(n7568), .X(n949) );
  nor_x2_sg U2247 ( .A(n951), .B(n952), .X(n950) );
  nor_x2_sg U2246 ( .A(n955), .B(n9084), .X(n951) );
  nor_x2_sg U2245 ( .A(\i_im[1][2] ), .B(n7560), .X(n955) );
  nor_x2_sg U2242 ( .A(\i_im[0][2] ), .B(n7562), .X(n957) );
  nor_x2_sg U2237 ( .A(n881), .B(n9104), .X(n945) );
  nor_x2_sg U2228 ( .A(n866), .B(n9144), .X(n936) );
  nor_x2_sg U2226 ( .A(n865), .B(n9164), .X(n937) );
  nor_x2_sg U2207 ( .A(n917), .B(n7568), .X(n916) );
  nor_x2_sg U2206 ( .A(n918), .B(n919), .X(n917) );
  nor_x2_sg U2205 ( .A(n922), .B(n9083), .X(n918) );
  nor_x2_sg U2204 ( .A(\i_im[1][1] ), .B(n7560), .X(n922) );
  nor_x2_sg U2201 ( .A(\i_im[0][1] ), .B(n7562), .X(n924) );
  nor_x2_sg U2196 ( .A(n7390), .B(n9103), .X(n912) );
  nor_x2_sg U2187 ( .A(n7382), .B(n9143), .X(n903) );
  nor_x2_sg U2185 ( .A(n7380), .B(n9163), .X(n904) );
  nand_x8_sg U1519 ( .A(n794), .B(n3096), .X(n792) );
  nand_x8_sg U1560 ( .A(n796), .B(n797), .X(n795) );
  nand_x8_sg U1602 ( .A(n799), .B(n7558), .X(n798) );
  nand_x8_sg U1644 ( .A(n801), .B(n802), .X(n800) );
  nand_x8_sg U1688 ( .A(n804), .B(n802), .X(n803) );
  nand_x8_sg U1730 ( .A(n796), .B(n802), .X(n805) );
  nand_x8_sg U1774 ( .A(n807), .B(n802), .X(n806) );
  nor_x2_sg U1773 ( .A(n3098), .B(n7559), .X(n807) );
  nand_x8_sg U1816 ( .A(n809), .B(n3099), .X(n808) );
  nand_x8_sg U1858 ( .A(n794), .B(n3099), .X(n810) );
  nand_x8_sg U1900 ( .A(n812), .B(n9205), .X(n811) );
  nand_x8_sg U1944 ( .A(n814), .B(n9205), .X(n813) );
  nand_x8_sg U1986 ( .A(n816), .B(n3099), .X(n815) );
  nand_x8_sg U2029 ( .A(n818), .B(n3099), .X(n817) );
  nand_x8_sg U2073 ( .A(n820), .B(n9205), .X(n819) );
  nand_x8_sg U2136 ( .A(n5893), .B(n9205), .X(n821) );
  nand_x8_sg U3590 ( .A(n9185), .B(n1576), .X(n838) );
  nand_x8_sg U3709 ( .A(n7523), .B(n5307), .X(n826) );
  nand_x8_sg U3689 ( .A(n5302), .B(n7522), .X(n834) );
  nor_x2_sg U3686 ( .A(n2060), .B(n7522), .X(n2059) );
  nor_x2_sg U3685 ( .A(n2061), .B(n9059), .X(n2060) );
  nor_x2_sg U3684 ( .A(n2066), .B(n2067), .X(n2061) );
  nand_x8_sg U3669 ( .A(n2058), .B(n7522), .X(n833) );
  nand_x8_sg U3664 ( .A(n2056), .B(n7522), .X(n835) );
  nand_x8_sg U3660 ( .A(n2055), .B(n7522), .X(n3101) );
  nand_x8_sg U3651 ( .A(n2038), .B(n7316), .X(n830) );
  nand_x8_sg U3646 ( .A(n2046), .B(n6383), .X(n832) );
  nand_x8_sg U3636 ( .A(n2039), .B(n6383), .X(n831) );
  nand_x8_sg U3632 ( .A(n2038), .B(n9219), .X(n828) );
  nand_x8_sg U3568 ( .A(n7310), .B(n9066), .X(n5286) );
  nand_x8_sg U3559 ( .A(n1838), .B(n7310), .X(n3814) );
  nor_x2_sg U3398 ( .A(n1805), .B(n1806), .X(n1801) );
  nor_x2_sg U3395 ( .A(n1851), .B(n9072), .X(n1846) );
  nor_x2_sg U3389 ( .A(n1848), .B(n9069), .X(n1847) );
  nor_x2_sg U3370 ( .A(n1831), .B(n9079), .X(n1825) );
  nor_x2_sg U3364 ( .A(n1827), .B(n9080), .X(n1826) );
  nor_x2_sg U3357 ( .A(n1821), .B(n1822), .X(n1815) );
  nor_x2_sg U3351 ( .A(n1817), .B(n1818), .X(n1816) );
  nand_x8_sg U2999 ( .A(n836), .B(n837), .X(n829) );
  nor_x2_sg U2998 ( .A(n7520), .B(n838), .X(n836) );
  nand_x8_sg U3089 ( .A(n9184), .B(n7318), .X(n841) );
  nand_x8_sg U3028 ( .A(n840), .B(n9186), .X(n839) );
  nor_x2_sg U3027 ( .A(n7520), .B(n841), .X(n840) );
  nand_x8_sg U3056 ( .A(n843), .B(n837), .X(n842) );
  nand_x8_sg U3087 ( .A(n844), .B(n9186), .X(n825) );
  inv_x4_sg U6688 ( .A(n7556), .X(n7555) );
  inv_x2_sg U6689 ( .A(n3104), .X(n7557) );
  nor_x1_sg U6690 ( .A(n7538), .B(reset), .X(n3104) );
  inv_x4_sg U6691 ( .A(n7539), .X(n7538) );
  inv_x2_sg U6692 ( .A(n9204), .X(n7539) );
  inv_x1_sg U6693 ( .A(n3807), .X(n9204) );
  nand_x2_sg U6694 ( .A(n928), .B(n929), .X(n774) );
  nand_x2_sg U6695 ( .A(n961), .B(n962), .X(n775) );
  nand_x2_sg U6696 ( .A(n994), .B(n995), .X(n776) );
  nand_x2_sg U6697 ( .A(n1096), .B(n1097), .X(n779) );
  nand_x2_sg U6698 ( .A(n1129), .B(n1130), .X(n780) );
  nand_x2_sg U6699 ( .A(n1162), .B(n1163), .X(n781) );
  nand_x2_sg U6700 ( .A(n1266), .B(n1267), .X(n784) );
  nand_x2_sg U6701 ( .A(n1299), .B(n1300), .X(n785) );
  nand_x2_sg U6702 ( .A(n1332), .B(n1333), .X(n786) );
  nand_x2_sg U6703 ( .A(n1434), .B(n1435), .X(n789) );
  nand_x2_sg U6704 ( .A(n1467), .B(n1468), .X(n790) );
  nand_x2_sg U6705 ( .A(n1500), .B(n1501), .X(n791) );
  inv_x2_sg U6706 ( .A(n3819), .X(n5924) );
  nor_x1_sg U6707 ( .A(n5310), .B(n5311), .X(n3819) );
  nand_x2_sg U6708 ( .A(n5290), .B(n5306), .X(n5277) );
  inv_x2_sg U6709 ( .A(n7036), .X(n7037) );
  inv_x1_sg U6710 ( .A(\update_mask_0/N25 ), .X(n7036) );
  inv_x4_sg U6711 ( .A(n7525), .X(n7524) );
  inv_x4_sg U6712 ( .A(n781), .X(n7353) );
  inv_x4_sg U6713 ( .A(n784), .X(n7359) );
  inv_x4_sg U6714 ( .A(n774), .X(n7338) );
  inv_x4_sg U6715 ( .A(n785), .X(n7361) );
  inv_x4_sg U6716 ( .A(n775), .X(n7340) );
  inv_x4_sg U6717 ( .A(n779), .X(n7349) );
  inv_x4_sg U6718 ( .A(n780), .X(n7351) );
  inv_x4_sg U6719 ( .A(n786), .X(n7363) );
  inv_x4_sg U6720 ( .A(n789), .X(n7369) );
  inv_x4_sg U6721 ( .A(n790), .X(n7371) );
  inv_x4_sg U6722 ( .A(n791), .X(n7373) );
  inv_x4_sg U6723 ( .A(n776), .X(n7342) );
  inv_x4_sg U6724 ( .A(n7557), .X(n7556) );
  inv_x4_sg U6725 ( .A(n777), .X(n7344) );
  inv_x4_sg U6726 ( .A(n7566), .X(n7565) );
  inv_x4_sg U6727 ( .A(n6048), .X(n7388) );
  inv_x4_sg U6728 ( .A(n879), .X(n7386) );
  inv_x4_sg U6729 ( .A(n4207), .X(n7399) );
  inv_x4_sg U6730 ( .A(n862), .X(n7378) );
  inv_x4_sg U6731 ( .A(n858), .X(n7376) );
  inv_x4_sg U6732 ( .A(n3827), .X(n7475) );
  inv_x4_sg U6733 ( .A(n3852), .X(n7481) );
  inv_x4_sg U6734 ( .A(n3876), .X(n7469) );
  inv_x4_sg U6735 ( .A(n3867), .X(n7477) );
  inv_x4_sg U6736 ( .A(n3873), .X(n7483) );
  inv_x4_sg U6737 ( .A(n3840), .X(n7471) );
  inv_x4_sg U6738 ( .A(n3843), .X(n7479) );
  inv_x4_sg U6739 ( .A(n3861), .X(n7485) );
  inv_x4_sg U6740 ( .A(n3855), .X(n7473) );
  inv_x4_sg U6741 ( .A(n4416), .X(n7438) );
  inv_x4_sg U6742 ( .A(n4451), .X(n7425) );
  inv_x4_sg U6743 ( .A(n4445), .X(n7322) );
  inv_x4_sg U6744 ( .A(n4415), .X(n7440) );
  inv_x4_sg U6745 ( .A(n4419), .X(n7436) );
  inv_x4_sg U6746 ( .A(n3864), .X(n7442) );
  inv_x4_sg U6747 ( .A(n3834), .X(n7467) );
  inv_x4_sg U6748 ( .A(n3849), .X(n7449) );
  inv_x4_sg U6749 ( .A(n3870), .X(n7444) );
  inv_x4_sg U6750 ( .A(n3858), .X(n7451) );
  inv_x4_sg U6751 ( .A(n3846), .X(n7453) );
  inv_x4_sg U6752 ( .A(n3879), .X(n7465) );
  inv_x4_sg U6753 ( .A(n3837), .X(n7487) );
  inv_x4_sg U6754 ( .A(n3885), .X(n7489) );
  inv_x4_sg U6755 ( .A(n3831), .X(n7493) );
  inv_x4_sg U6756 ( .A(n3882), .X(n7491) );
  inv_x1_sg U6757 ( .A(n5926), .X(n5927) );
  inv_x4_sg U6758 ( .A(n7037), .X(n7521) );
  nor_x2_sg U6759 ( .A(n5889), .B(n5891), .X(n5314) );
  inv_x1_sg U6760 ( .A(n5321), .X(n5886) );
  inv_x2_sg U6761 ( .A(n5886), .X(n5887) );
  inv_x1_sg U6762 ( .A(n5315), .X(n5888) );
  inv_x2_sg U6763 ( .A(n5888), .X(n5889) );
  inv_x1_sg U6764 ( .A(n5316), .X(n5890) );
  inv_x2_sg U6765 ( .A(n5890), .X(n5891) );
  inv_x1_sg U6766 ( .A(n822), .X(n5892) );
  inv_x2_sg U6767 ( .A(n5892), .X(n5893) );
  inv_x1_sg U6768 ( .A(\update_output_0/N28 ), .X(n5894) );
  inv_x2_sg U6769 ( .A(n5894), .X(n5895) );
  inv_x1_sg U6770 ( .A(\update_output_0/n9020 ), .X(n5896) );
  inv_x2_sg U6771 ( .A(n5896), .X(n5897) );
  inv_x1_sg U6772 ( .A(\update_output_0/n9019 ), .X(n5898) );
  inv_x2_sg U6773 ( .A(n5898), .X(n5899) );
  inv_x1_sg U6774 ( .A(\update_output_0/N30 ), .X(n5900) );
  inv_x2_sg U6775 ( .A(n5900), .X(n5901) );
  inv_x1_sg U6776 ( .A(\update_output_0/N31 ), .X(n5902) );
  inv_x2_sg U6777 ( .A(n5902), .X(n5903) );
  inv_x1_sg U6778 ( .A(\update_output_0/N32 ), .X(n5904) );
  inv_x2_sg U6779 ( .A(n5904), .X(n5905) );
  inv_x1_sg U6780 ( .A(\update_output_0/N34 ), .X(n5906) );
  inv_x2_sg U6781 ( .A(n5906), .X(n5907) );
  inv_x1_sg U6782 ( .A(\update_mask_0/N23 ), .X(n5908) );
  inv_x2_sg U6783 ( .A(n5908), .X(n5909) );
  inv_x1_sg U6784 ( .A(\update_mask_0/n4205 ), .X(n5910) );
  inv_x2_sg U6785 ( .A(n5910), .X(n5911) );
  inv_x1_sg U6786 ( .A(\update_mask_0/n4206 ), .X(n5912) );
  inv_x2_sg U6787 ( .A(n5912), .X(n5913) );
  inv_x1_sg U6788 ( .A(\update_mask_0/N26 ), .X(n5914) );
  inv_x2_sg U6789 ( .A(n5914), .X(n5915) );
  inv_x1_sg U6790 ( .A(\update_mask_0/N24 ), .X(n5916) );
  inv_x2_sg U6791 ( .A(n5916), .X(n5917) );
  inv_x1_sg U6792 ( .A(\update_mask_0/N28 ), .X(n5918) );
  inv_x2_sg U6793 ( .A(n5918), .X(n5919) );
  inv_x1_sg U6794 ( .A(\update_mask_0/N30 ), .X(n5920) );
  inv_x2_sg U6795 ( .A(n5920), .X(n5921) );
  inv_x1_sg U6796 ( .A(\update_mask_0/N31 ), .X(n5922) );
  inv_x2_sg U6797 ( .A(n5922), .X(n5923) );
  nor_x2_sg U6798 ( .A(n9218), .B(n3824), .X(n3821) );
  nor_x2_sg U6799 ( .A(n3821), .B(n3822), .X(n3820) );
  nor_x2_sg U6800 ( .A(n9198), .B(n3823), .X(n3822) );
  inv_x1_sg U6801 ( .A(\update_mask_0/reg_i_mask [9]), .X(n5931) );
  inv_x1_sg U6802 ( .A(\update_mask_0/reg_i_mask [11]), .X(n5933) );
  inv_x1_sg U6803 ( .A(\update_mask_0/reg_i_mask [16]), .X(n5935) );
  inv_x1_sg U6804 ( .A(\update_mask_0/reg_i_mask [17]), .X(n5937) );
  inv_x1_sg U6805 ( .A(\update_mask_0/reg_i_mask [19]), .X(n5939) );
  inv_x1_sg U6806 ( .A(\update_mask_0/reg_i_mask [24]), .X(n5941) );
  inv_x1_sg U6807 ( .A(\update_mask_0/reg_i_mask [25]), .X(n5943) );
  inv_x1_sg U6808 ( .A(\update_mask_0/reg_i_mask [27]), .X(n5945) );
  inv_x4_sg U6809 ( .A(n5924), .X(n5925) );
  inv_x1_sg U6810 ( .A(\update_mask_0/reg_i_mask [12]), .X(n5963) );
  inv_x1_sg U6811 ( .A(\update_mask_0/reg_i_mask [13]), .X(n5965) );
  inv_x1_sg U6812 ( .A(\update_mask_0/reg_i_mask [18]), .X(n5969) );
  inv_x1_sg U6813 ( .A(\update_mask_0/reg_i_mask [20]), .X(n5971) );
  inv_x1_sg U6814 ( .A(\update_mask_0/reg_i_mask [21]), .X(n5973) );
  inv_x1_sg U6815 ( .A(\update_mask_0/reg_i_mask [26]), .X(n5977) );
  inv_x1_sg U6816 ( .A(\update_mask_0/reg_i_mask [28]), .X(n5979) );
  inv_x1_sg U6817 ( .A(\update_mask_0/reg_i_mask [29]), .X(n5981) );
  nand_x4_sg U6818 ( .A(n2070), .B(n5988), .X(n5312) );
  nor_x2_sg U6819 ( .A(n7316), .B(n9215), .X(n2056) );
  nor_x2_sg U6820 ( .A(n9241), .B(n8990), .X(n812) );
  inv_x4_sg U6821 ( .A(n3824), .X(n9198) );
  nand_x4_sg U6822 ( .A(n5292), .B(n5312), .X(n3824) );
  inv_x1_sg U6823 ( .A(n5325), .X(n5929) );
  inv_x4_sg U6824 ( .A(n3816), .X(n5926) );
  nor_x2_sg U6825 ( .A(n5274), .B(n7308), .X(n5284) );
  inv_x1_sg U6826 ( .A(n1992), .X(n5928) );
  nand_x4_sg U6827 ( .A(n9184), .B(n827), .X(n1992) );
  inv_x8_sg U6828 ( .A(n7312), .X(n7541) );
  nand_x4_sg U6829 ( .A(n7400), .B(n3100), .X(n4206) );
  nor_x2_sg U6830 ( .A(n5952), .B(n5988), .X(n3809) );
  inv_x8_sg U6831 ( .A(n831), .X(n9064) );
  inv_x8_sg U6832 ( .A(n830), .X(n9063) );
  inv_x8_sg U6833 ( .A(n832), .X(n9216) );
  nor_x2_sg U6834 ( .A(n5318), .B(n5319), .X(n5317) );
  inv_x2_sg U6835 ( .A(n4202), .X(n9196) );
  inv_x1_sg U6836 ( .A(\update_mask_0/reg_out[10][19] ), .X(n5947) );
  inv_x2_sg U6837 ( .A(n5929), .X(n5930) );
  nor_x2_sg U6838 ( .A(n5327), .B(n5319), .X(n5326) );
  nor_x4_sg U6839 ( .A(n4297), .B(n9243), .X(n4419) );
  inv_x4_sg U6840 ( .A(n826), .X(n9184) );
  nor_x2_sg U6841 ( .A(n5990), .B(n9209), .X(n4201) );
  inv_x4_sg U6842 ( .A(output_taken), .X(n9209) );
  nor_x4_sg U6843 ( .A(n7541), .B(n8990), .X(n794) );
  inv_x8_sg U6844 ( .A(n5313), .X(n9207) );
  nand_x4_sg U6845 ( .A(n3809), .B(input_ready), .X(n5313) );
  nand_x2_sg U6846 ( .A(n9218), .B(n9246), .X(n5327) );
  inv_x8_sg U6847 ( .A(n5952), .X(n9218) );
  nor_x8_sg U6848 ( .A(n9246), .B(n5950), .X(n3100) );
  inv_x8_sg U6849 ( .A(n5990), .X(n9246) );
  inv_x8_sg U6850 ( .A(n828), .X(n9062) );
  inv_x8_sg U6851 ( .A(n835), .X(n9065) );
  inv_x8_sg U6852 ( .A(n834), .X(n9057) );
  inv_x8_sg U6853 ( .A(n833), .X(n9060) );
  nor_x2_sg U6854 ( .A(n6383), .B(n7316), .X(n2058) );
  nor_x2_sg U6855 ( .A(n7522), .B(n9219), .X(n2046) );
  nand_x2_sg U6856 ( .A(\update_mask_0/n919 ), .B(n5292), .X(n5291) );
  nor_x8_sg U6857 ( .A(reset), .B(n9207), .X(n5292) );
  nor_x2_sg U6858 ( .A(n3098), .B(n8990), .X(n799) );
  inv_x1_sg U6859 ( .A(\update_mask_0/reg_i_mask [4]), .X(n5953) );
  inv_x1_sg U6860 ( .A(\update_mask_0/reg_i_mask [5]), .X(n5955) );
  inv_x1_sg U6861 ( .A(\update_mask_0/reg_i_mask [6]), .X(n5957) );
  inv_x1_sg U6862 ( .A(\update_mask_0/reg_i_mask [8]), .X(n5959) );
  inv_x1_sg U6863 ( .A(\update_mask_0/reg_i_mask [10]), .X(n5961) );
  inv_x1_sg U6864 ( .A(\update_mask_0/reg_i_mask [14]), .X(n5967) );
  inv_x1_sg U6865 ( .A(\update_mask_0/reg_i_mask [22]), .X(n5975) );
  inv_x1_sg U6866 ( .A(\update_mask_0/reg_i_mask [30]), .X(n5983) );
  inv_x1_sg U6867 ( .A(\update_mask_0/reg_out[6][19] ), .X(n5985) );
  nor_x4_sg U6868 ( .A(n4297), .B(n9242), .X(n4415) );
  nor_x8_sg U6869 ( .A(n7571), .B(n9242), .X(n4437) );
  inv_x8_sg U6870 ( .A(n5241), .X(n9242) );
  nor_x8_sg U6871 ( .A(n9243), .B(n7571), .X(n4436) );
  inv_x8_sg U6872 ( .A(n5242), .X(n9243) );
  inv_x2_sg U6873 ( .A(n5931), .X(n5932) );
  inv_x2_sg U6874 ( .A(n5933), .X(n5934) );
  inv_x2_sg U6875 ( .A(n5935), .X(n5936) );
  inv_x2_sg U6876 ( .A(n5937), .X(n5938) );
  inv_x2_sg U6877 ( .A(n5939), .X(n5940) );
  inv_x2_sg U6878 ( .A(n5941), .X(n5942) );
  inv_x2_sg U6879 ( .A(n5943), .X(n5944) );
  inv_x2_sg U6880 ( .A(n5945), .X(n5946) );
  inv_x2_sg U6881 ( .A(n5947), .X(n5948) );
  inv_x8_sg U6882 ( .A(n7312), .X(n7540) );
  nor_x8_sg U6883 ( .A(n9218), .B(n5988), .X(n5307) );
  inv_x4_sg U6884 ( .A(n5899), .X(n5949) );
  inv_x8_sg U6885 ( .A(n5949), .X(n5950) );
  nand_x4_sg U6886 ( .A(n5950), .B(n5988), .X(n5319) );
  inv_x4_sg U6887 ( .A(n5913), .X(n5951) );
  inv_x8_sg U6888 ( .A(n5951), .X(n5952) );
  nor_x8_sg U6889 ( .A(n1553), .B(n841), .X(n1537) );
  nand_x8_sg U6890 ( .A(n838), .B(n7520), .X(n1553) );
  inv_x8_sg U6891 ( .A(n1567), .X(n9188) );
  nand_x4_sg U6892 ( .A(n1568), .B(n837), .X(n1567) );
  nor_x2_sg U6893 ( .A(n7522), .B(n7316), .X(n2039) );
  inv_x2_sg U6894 ( .A(n880), .X(n6047) );
  inv_x4_sg U6895 ( .A(input_ready), .X(n9208) );
  nor_x2_sg U6896 ( .A(n7312), .B(n9183), .X(n801) );
  nor_x2_sg U6897 ( .A(n7541), .B(n9183), .X(n804) );
  inv_x4_sg U6898 ( .A(n3096), .X(n9183) );
  nor_x4_sg U6899 ( .A(n3930), .B(n9244), .X(n4202) );
  inv_x4_sg U6900 ( .A(n4206), .X(n9244) );
  inv_x2_sg U6901 ( .A(n5953), .X(n5954) );
  inv_x2_sg U6902 ( .A(n5955), .X(n5956) );
  inv_x2_sg U6903 ( .A(n5957), .X(n5958) );
  inv_x2_sg U6904 ( .A(n5959), .X(n5960) );
  inv_x2_sg U6905 ( .A(n5961), .X(n5962) );
  inv_x2_sg U6906 ( .A(n5963), .X(n5964) );
  inv_x2_sg U6907 ( .A(n5965), .X(n5966) );
  inv_x2_sg U6908 ( .A(n5967), .X(n5968) );
  inv_x2_sg U6909 ( .A(n5969), .X(n5970) );
  inv_x2_sg U6910 ( .A(n5971), .X(n5972) );
  inv_x2_sg U6911 ( .A(n5973), .X(n5974) );
  inv_x2_sg U6912 ( .A(n5975), .X(n5976) );
  inv_x2_sg U6913 ( .A(n5977), .X(n5978) );
  inv_x2_sg U6914 ( .A(n5979), .X(n5980) );
  inv_x2_sg U6915 ( .A(n5981), .X(n5982) );
  inv_x2_sg U6916 ( .A(n5983), .X(n5984) );
  inv_x2_sg U6917 ( .A(n5985), .X(n5986) );
  nor_x4_sg U6918 ( .A(n7312), .B(n8990), .X(n809) );
  nor_x4_sg U6919 ( .A(n9241), .B(n3098), .X(n796) );
  nor_x4_sg U6920 ( .A(n5274), .B(n5283), .X(n3813) );
  nor_x2_sg U6921 ( .A(n7312), .B(n8991), .X(n816) );
  nor_x2_sg U6922 ( .A(n7540), .B(n8991), .X(n818) );
  nor_x2_sg U6923 ( .A(n9241), .B(n8991), .X(n820) );
  inv_x8_sg U6924 ( .A(n802), .X(n8991) );
  inv_x4_sg U6925 ( .A(n5911), .X(n5987) );
  inv_x8_sg U6926 ( .A(n5987), .X(n5988) );
  inv_x4_sg U6927 ( .A(n5897), .X(n5989) );
  inv_x8_sg U6928 ( .A(n5989), .X(n5990) );
  inv_x8_sg U6929 ( .A(n1833), .X(n9078) );
  nand_x8_sg U6930 ( .A(n1839), .B(n9077), .X(n1833) );
  nor_x8_sg U6931 ( .A(n9245), .B(n7570), .X(n797) );
  nor_x8_sg U6932 ( .A(n7571), .B(n9245), .X(n802) );
  inv_x8_sg U6933 ( .A(n3100), .X(n9245) );
  nor_x8_sg U6934 ( .A(n1575), .B(n841), .X(n1558) );
  nand_x8_sg U6935 ( .A(n7519), .B(n838), .X(n1575) );
  inv_x8_sg U6936 ( .A(n1564), .X(n9187) );
  nand_x4_sg U6937 ( .A(n1565), .B(n837), .X(n1564) );
  inv_x4_sg U6938 ( .A(n5905), .X(n5991) );
  inv_x8_sg U6939 ( .A(n5991), .X(n5992) );
  nor_x8_sg U6940 ( .A(n7312), .B(n5992), .X(n5242) );
  nor_x8_sg U6941 ( .A(n3098), .B(n5992), .X(n3096) );
  nor_x8_sg U6942 ( .A(n4393), .B(n5992), .X(n3099) );
  nor_x8_sg U6943 ( .A(n7540), .B(n5992), .X(n5241) );
  nand_x1_sg U6944 ( .A(\i_im[3][0] ), .B(n7393), .X(n886) );
  nand_x1_sg U6945 ( .A(\i_im[2][0] ), .B(n7392), .X(n887) );
  nand_x1_sg U6946 ( .A(\i_im[3][1] ), .B(n7393), .X(n920) );
  nand_x1_sg U6947 ( .A(\i_im[2][1] ), .B(n7392), .X(n921) );
  nand_x1_sg U6948 ( .A(\i_im[3][2] ), .B(n7393), .X(n953) );
  nand_x1_sg U6949 ( .A(\i_im[2][2] ), .B(n7392), .X(n954) );
  nand_x1_sg U6950 ( .A(\i_im[3][3] ), .B(n7393), .X(n986) );
  nand_x1_sg U6951 ( .A(\i_im[2][3] ), .B(n7392), .X(n987) );
  nand_x1_sg U6952 ( .A(\i_im[3][4] ), .B(n7393), .X(n1019) );
  nand_x1_sg U6953 ( .A(\i_im[2][4] ), .B(n7392), .X(n1020) );
  nand_x1_sg U6954 ( .A(\i_im[3][5] ), .B(n7393), .X(n1055) );
  nand_x1_sg U6955 ( .A(\i_im[2][5] ), .B(n7392), .X(n1056) );
  nand_x1_sg U6956 ( .A(\i_im[3][6] ), .B(n7393), .X(n1088) );
  nand_x1_sg U6957 ( .A(\i_im[2][6] ), .B(n7392), .X(n1089) );
  nand_x1_sg U6958 ( .A(\i_im[3][7] ), .B(n7393), .X(n1121) );
  nand_x1_sg U6959 ( .A(\i_im[2][7] ), .B(n7392), .X(n1122) );
  nand_x1_sg U6960 ( .A(\i_im[3][8] ), .B(n7393), .X(n1154) );
  nand_x1_sg U6961 ( .A(\i_im[2][8] ), .B(n7392), .X(n1155) );
  nand_x1_sg U6962 ( .A(\i_im[3][9] ), .B(n7393), .X(n1187) );
  nand_x1_sg U6963 ( .A(\i_im[2][9] ), .B(n7392), .X(n1188) );
  nand_x1_sg U6964 ( .A(\i_im[3][10] ), .B(n7393), .X(n1225) );
  nand_x1_sg U6965 ( .A(\i_im[2][10] ), .B(n7392), .X(n1226) );
  nand_x1_sg U6966 ( .A(\i_im[3][11] ), .B(n7393), .X(n1258) );
  nand_x1_sg U6967 ( .A(\i_im[2][11] ), .B(n7392), .X(n1259) );
  nand_x1_sg U6968 ( .A(\i_im[3][12] ), .B(n7393), .X(n1291) );
  nand_x1_sg U6969 ( .A(\i_im[2][12] ), .B(n7392), .X(n1292) );
  nand_x1_sg U6970 ( .A(\i_im[3][13] ), .B(n7393), .X(n1324) );
  nand_x1_sg U6971 ( .A(\i_im[2][13] ), .B(n7392), .X(n1325) );
  nand_x1_sg U6972 ( .A(\i_im[3][14] ), .B(n7393), .X(n1357) );
  nand_x1_sg U6973 ( .A(\i_im[2][14] ), .B(n7392), .X(n1358) );
  nand_x1_sg U6974 ( .A(\i_im[3][15] ), .B(n7393), .X(n1393) );
  nand_x1_sg U6975 ( .A(\i_im[2][15] ), .B(n7392), .X(n1394) );
  nand_x1_sg U6976 ( .A(\i_im[3][16] ), .B(n7393), .X(n1426) );
  nand_x1_sg U6977 ( .A(\i_im[2][16] ), .B(n7392), .X(n1427) );
  nand_x1_sg U6978 ( .A(\i_im[3][17] ), .B(n7393), .X(n1459) );
  nand_x1_sg U6979 ( .A(\i_im[2][17] ), .B(n7392), .X(n1460) );
  nand_x1_sg U6980 ( .A(\i_im[3][18] ), .B(n7393), .X(n1492) );
  nand_x1_sg U6981 ( .A(\i_im[2][18] ), .B(n7392), .X(n1493) );
  nand_x1_sg U6982 ( .A(\i_im[3][19] ), .B(n7393), .X(n1528) );
  nand_x1_sg U6983 ( .A(\i_im[2][19] ), .B(n7392), .X(n1529) );
  nand_x1_sg U6984 ( .A(n1591), .B(n1592), .X(n1590) );
  nand_x1_sg U6985 ( .A(n1602), .B(n1603), .X(n1601) );
  nand_x1_sg U6986 ( .A(n1625), .B(n1626), .X(n1624) );
  nand_x1_sg U6987 ( .A(n1836), .B(n1837), .X(n1835) );
  nand_x1_sg U6988 ( .A(n1813), .B(n1814), .X(n1812) );
  nand_x1_sg U6989 ( .A(n1755), .B(n1756), .X(n1754) );
  nand_x1_sg U6990 ( .A(n1765), .B(n1766), .X(n1764) );
  nand_x1_sg U6991 ( .A(n1787), .B(n1788), .X(n1786) );
  nand_x1_sg U6992 ( .A(n1905), .B(n1906), .X(n1904) );
  nand_x1_sg U6993 ( .A(n1915), .B(n1916), .X(n1914) );
  nand_x1_sg U6994 ( .A(n1937), .B(n1938), .X(n1936) );
  nand_x1_sg U6995 ( .A(n7558), .B(n5545), .X(n5259) );
  nand_x1_sg U6996 ( .A(n7323), .B(n5546), .X(n5260) );
  nand_x1_sg U6997 ( .A(\update_output_0/n6424 ), .B(n7540), .X(n5263) );
  nand_x1_sg U6998 ( .A(n7558), .B(n5534), .X(n4572) );
  nand_x1_sg U6999 ( .A(n7323), .B(n5535), .X(n4573) );
  nand_x1_sg U7000 ( .A(\update_output_0/n6425 ), .B(n7540), .X(n4576) );
  nand_x1_sg U7001 ( .A(n7558), .B(n5523), .X(n4530) );
  nand_x1_sg U7002 ( .A(n7323), .B(n5524), .X(n4531) );
  nand_x1_sg U7003 ( .A(\update_output_0/n6426 ), .B(n7541), .X(n4534) );
  nand_x1_sg U7004 ( .A(n7558), .B(n5512), .X(n4443) );
  nand_x1_sg U7005 ( .A(n7323), .B(n5513), .X(n4444) );
  nand_x1_sg U7006 ( .A(\update_output_0/n6427 ), .B(n7541), .X(n4448) );
  nand_x1_sg U7007 ( .A(n7558), .B(n5501), .X(n4488) );
  nand_x1_sg U7008 ( .A(n7323), .B(n5502), .X(n4489) );
  nand_x1_sg U7009 ( .A(\update_output_0/n6428 ), .B(n7541), .X(n4492) );
  nand_x1_sg U7010 ( .A(n7558), .B(n5490), .X(n4700) );
  nand_x1_sg U7011 ( .A(n7323), .B(n5491), .X(n4701) );
  nand_x1_sg U7012 ( .A(\update_output_0/n6429 ), .B(n7540), .X(n4704) );
  nand_x1_sg U7013 ( .A(n7558), .B(n5479), .X(n4742) );
  nand_x1_sg U7014 ( .A(n7323), .B(n5480), .X(n4743) );
  nand_x1_sg U7015 ( .A(\update_output_0/n6430 ), .B(n7540), .X(n4746) );
  nand_x1_sg U7016 ( .A(n7558), .B(n5468), .X(n4656) );
  nand_x1_sg U7017 ( .A(n7323), .B(n5469), .X(n4657) );
  nand_x1_sg U7018 ( .A(\update_output_0/n6431 ), .B(n7540), .X(n4660) );
  nand_x1_sg U7019 ( .A(n7558), .B(n5457), .X(n4614) );
  nand_x1_sg U7020 ( .A(n7323), .B(n5458), .X(n4615) );
  nand_x1_sg U7021 ( .A(\update_output_0/n6432 ), .B(n7541), .X(n4618) );
  nand_x1_sg U7022 ( .A(n7558), .B(n5446), .X(n4952) );
  nand_x1_sg U7023 ( .A(n7323), .B(n5447), .X(n4953) );
  nand_x1_sg U7024 ( .A(\update_output_0/n6433 ), .B(n7540), .X(n4956) );
  nand_x1_sg U7025 ( .A(n7558), .B(n5435), .X(n4994) );
  nand_x1_sg U7026 ( .A(n7323), .B(n5436), .X(n4995) );
  nand_x1_sg U7027 ( .A(\update_output_0/n6434 ), .B(n7541), .X(n4998) );
  nand_x1_sg U7028 ( .A(n7558), .B(n5424), .X(n5180) );
  nand_x1_sg U7029 ( .A(n7323), .B(n5425), .X(n5181) );
  nand_x1_sg U7030 ( .A(\update_output_0/n6435 ), .B(n7541), .X(n5184) );
  nand_x1_sg U7031 ( .A(n7558), .B(n5413), .X(n5220) );
  nand_x1_sg U7032 ( .A(n7323), .B(n5414), .X(n5221) );
  nand_x1_sg U7033 ( .A(\update_output_0/n6436 ), .B(n7541), .X(n5224) );
  nand_x1_sg U7034 ( .A(n7558), .B(n5402), .X(n5144) );
  nand_x1_sg U7035 ( .A(n7323), .B(n5403), .X(n5145) );
  nand_x1_sg U7036 ( .A(\update_output_0/n6437 ), .B(n7541), .X(n5148) );
  nand_x1_sg U7037 ( .A(n7558), .B(n5391), .X(n5108) );
  nand_x1_sg U7038 ( .A(n4445), .B(n5392), .X(n5109) );
  nand_x1_sg U7039 ( .A(\update_output_0/n6438 ), .B(n7541), .X(n5112) );
  nand_x1_sg U7040 ( .A(n7558), .B(n5380), .X(n4868) );
  nand_x1_sg U7041 ( .A(n7323), .B(n5381), .X(n4869) );
  nand_x1_sg U7042 ( .A(\update_output_0/n6439 ), .B(n7541), .X(n4872) );
  nand_x1_sg U7043 ( .A(n5994), .B(n5369), .X(n4910) );
  nand_x1_sg U7044 ( .A(n7323), .B(n5370), .X(n4911) );
  nand_x1_sg U7045 ( .A(\update_output_0/n6440 ), .B(n7541), .X(n4914) );
  nand_x1_sg U7046 ( .A(n7558), .B(n5358), .X(n4784) );
  nand_x1_sg U7047 ( .A(n7323), .B(n5359), .X(n4785) );
  nand_x1_sg U7048 ( .A(\update_output_0/n6441 ), .B(n7541), .X(n4788) );
  nand_x1_sg U7049 ( .A(n7558), .B(n5347), .X(n4826) );
  nand_x1_sg U7050 ( .A(n7323), .B(n5348), .X(n4827) );
  nand_x1_sg U7051 ( .A(\update_output_0/n6442 ), .B(n7540), .X(n4830) );
  nand_x1_sg U7052 ( .A(n7558), .B(n5336), .X(n5036) );
  nand_x1_sg U7053 ( .A(n7323), .B(n5337), .X(n5037) );
  nand_x1_sg U7054 ( .A(\update_output_0/n6443 ), .B(n7540), .X(n5040) );
  nand_x1_sg U7055 ( .A(\i_im[5][0] ), .B(n7389), .X(n877) );
  nand_x1_sg U7056 ( .A(\i_im[4][0] ), .B(n7387), .X(n878) );
  nand_x1_sg U7057 ( .A(\i_im[5][1] ), .B(n7389), .X(n914) );
  nand_x1_sg U7058 ( .A(\i_im[4][1] ), .B(n7387), .X(n915) );
  nand_x1_sg U7059 ( .A(\i_im[5][2] ), .B(n7389), .X(n947) );
  nand_x1_sg U7060 ( .A(\i_im[4][2] ), .B(n7387), .X(n948) );
  nand_x1_sg U7061 ( .A(\i_im[5][3] ), .B(n7389), .X(n980) );
  nand_x1_sg U7062 ( .A(\i_im[4][3] ), .B(n7387), .X(n981) );
  nand_x1_sg U7063 ( .A(\i_im[5][4] ), .B(n7389), .X(n1013) );
  nand_x1_sg U7064 ( .A(\i_im[4][4] ), .B(n7387), .X(n1014) );
  nand_x1_sg U7065 ( .A(\i_im[5][5] ), .B(n7389), .X(n1049) );
  nand_x1_sg U7066 ( .A(\i_im[4][5] ), .B(n7387), .X(n1050) );
  nand_x1_sg U7067 ( .A(\i_im[5][6] ), .B(n7389), .X(n1082) );
  nand_x1_sg U7068 ( .A(\i_im[4][6] ), .B(n7387), .X(n1083) );
  nand_x1_sg U7069 ( .A(\i_im[5][7] ), .B(n7389), .X(n1115) );
  nand_x1_sg U7070 ( .A(\i_im[4][7] ), .B(n7387), .X(n1116) );
  nand_x1_sg U7071 ( .A(\i_im[5][8] ), .B(n6048), .X(n1148) );
  nand_x1_sg U7072 ( .A(\i_im[4][8] ), .B(n879), .X(n1149) );
  nand_x1_sg U7073 ( .A(\i_im[5][9] ), .B(n7389), .X(n1181) );
  nand_x1_sg U7074 ( .A(\i_im[4][9] ), .B(n7387), .X(n1182) );
  nand_x1_sg U7075 ( .A(\i_im[5][10] ), .B(n7389), .X(n1219) );
  nand_x1_sg U7076 ( .A(\i_im[4][10] ), .B(n7387), .X(n1220) );
  nand_x1_sg U7077 ( .A(\i_im[5][11] ), .B(n7389), .X(n1252) );
  nand_x1_sg U7078 ( .A(\i_im[4][11] ), .B(n7387), .X(n1253) );
  nand_x1_sg U7079 ( .A(\i_im[5][12] ), .B(n7389), .X(n1285) );
  nand_x1_sg U7080 ( .A(\i_im[4][12] ), .B(n7387), .X(n1286) );
  nand_x1_sg U7081 ( .A(\i_im[5][13] ), .B(n7389), .X(n1318) );
  nand_x1_sg U7082 ( .A(\i_im[4][13] ), .B(n7387), .X(n1319) );
  nand_x1_sg U7083 ( .A(\i_im[5][14] ), .B(n7389), .X(n1351) );
  nand_x1_sg U7084 ( .A(\i_im[4][14] ), .B(n7387), .X(n1352) );
  nand_x1_sg U7085 ( .A(\i_im[5][15] ), .B(n7389), .X(n1387) );
  nand_x1_sg U7086 ( .A(\i_im[4][15] ), .B(n7387), .X(n1388) );
  nand_x1_sg U7087 ( .A(\i_im[5][16] ), .B(n7389), .X(n1420) );
  nand_x1_sg U7088 ( .A(\i_im[4][16] ), .B(n7387), .X(n1421) );
  nand_x1_sg U7089 ( .A(\i_im[5][17] ), .B(n7389), .X(n1453) );
  nand_x1_sg U7090 ( .A(\i_im[4][17] ), .B(n7387), .X(n1454) );
  nand_x1_sg U7091 ( .A(\i_im[5][18] ), .B(n7389), .X(n1486) );
  nand_x1_sg U7092 ( .A(\i_im[4][18] ), .B(n7387), .X(n1487) );
  nand_x1_sg U7093 ( .A(\i_im[5][19] ), .B(n7389), .X(n1522) );
  nand_x1_sg U7094 ( .A(\i_im[4][19] ), .B(n7387), .X(n1523) );
  nand_x1_sg U7095 ( .A(n1654), .B(n1655), .X(n1653) );
  nand_x1_sg U7096 ( .A(n1640), .B(n1641), .X(n1639) );
  nand_x1_sg U7097 ( .A(n7320), .B(n1643), .X(n1637) );
  nand_x1_sg U7098 ( .A(n1644), .B(n1645), .X(n1643) );
  nand_x1_sg U7099 ( .A(n1650), .B(n1651), .X(n1649) );
  nand_x1_sg U7100 ( .A(n1662), .B(n1663), .X(n1661) );
  nand_x1_sg U7101 ( .A(n1672), .B(n1673), .X(n1671) );
  nand_x1_sg U7102 ( .A(n1676), .B(n1677), .X(n1675) );
  nand_x1_sg U7103 ( .A(n1666), .B(n1667), .X(n1665) );
  nand_x1_sg U7104 ( .A(n1618), .B(n1619), .X(n1617) );
  nand_x1_sg U7105 ( .A(n1614), .B(n1615), .X(n1613) );
  nand_x1_sg U7106 ( .A(n7320), .B(n1595), .X(n1588) );
  nand_x1_sg U7107 ( .A(n1596), .B(n1597), .X(n1595) );
  nand_x1_sg U7108 ( .A(n1606), .B(n1607), .X(n1605) );
  nand_x1_sg U7109 ( .A(n1629), .B(n1630), .X(n1628) );
  nand_x1_sg U7110 ( .A(n1718), .B(n1719), .X(n1717) );
  nand_x1_sg U7111 ( .A(n1704), .B(n1705), .X(n1703) );
  nand_x1_sg U7112 ( .A(n7320), .B(n1707), .X(n1701) );
  nand_x1_sg U7113 ( .A(n1708), .B(n1709), .X(n1707) );
  nand_x1_sg U7114 ( .A(n1714), .B(n1715), .X(n1713) );
  nand_x1_sg U7115 ( .A(n1726), .B(n1727), .X(n1725) );
  nand_x1_sg U7116 ( .A(n1736), .B(n1737), .X(n1735) );
  nand_x1_sg U7117 ( .A(n1740), .B(n1741), .X(n1739) );
  nand_x1_sg U7118 ( .A(n1730), .B(n1731), .X(n1729) );
  nand_x1_sg U7119 ( .A(n1842), .B(n1843), .X(n1841) );
  nand_x1_sg U7120 ( .A(n9067), .B(n1812), .X(n1807) );
  nand_x1_sg U7121 ( .A(n1809), .B(n1810), .X(n1808) );
  inv_x1_sg U7122 ( .A(n1835), .X(n9067) );
  nand_x1_sg U7123 ( .A(n1781), .B(n1782), .X(n1780) );
  nand_x1_sg U7124 ( .A(n1777), .B(n1778), .X(n1776) );
  nand_x1_sg U7125 ( .A(n7320), .B(n1758), .X(n1752) );
  nand_x1_sg U7126 ( .A(n1759), .B(n1760), .X(n1758) );
  nand_x1_sg U7127 ( .A(n1769), .B(n1770), .X(n1768) );
  nand_x1_sg U7128 ( .A(n1791), .B(n1792), .X(n1790) );
  nand_x1_sg U7129 ( .A(n1864), .B(n1865), .X(n1859) );
  nand_x1_sg U7130 ( .A(n1861), .B(n1862), .X(n1860) );
  nand_x1_sg U7131 ( .A(n1873), .B(n1874), .X(n1867) );
  nand_x1_sg U7132 ( .A(n1869), .B(n1870), .X(n1868) );
  nand_x1_sg U7133 ( .A(n1881), .B(n1882), .X(n1880) );
  nand_x1_sg U7134 ( .A(n1884), .B(n1885), .X(n1879) );
  nand_x1_sg U7135 ( .A(n1889), .B(n1890), .X(n1888) );
  nand_x1_sg U7136 ( .A(n1892), .B(n1893), .X(n1887) );
  nand_x1_sg U7137 ( .A(n1967), .B(n1968), .X(n1966) );
  nand_x1_sg U7138 ( .A(n1952), .B(n1953), .X(n1951) );
  nand_x1_sg U7139 ( .A(n7320), .B(n1955), .X(n1949) );
  nand_x1_sg U7140 ( .A(n1956), .B(n1957), .X(n1955) );
  nand_x1_sg U7141 ( .A(n1962), .B(n1963), .X(n1961) );
  nand_x1_sg U7142 ( .A(n1975), .B(n1976), .X(n1974) );
  nand_x1_sg U7143 ( .A(n1985), .B(n1986), .X(n1984) );
  nand_x1_sg U7144 ( .A(n1989), .B(n1990), .X(n1988) );
  nand_x1_sg U7145 ( .A(n1979), .B(n1980), .X(n1978) );
  nand_x1_sg U7146 ( .A(n1931), .B(n1932), .X(n1930) );
  nand_x1_sg U7147 ( .A(n1927), .B(n1928), .X(n1926) );
  nand_x1_sg U7148 ( .A(n7320), .B(n1908), .X(n1902) );
  nand_x1_sg U7149 ( .A(n1909), .B(n1910), .X(n1908) );
  nand_x1_sg U7150 ( .A(n1919), .B(n1920), .X(n1918) );
  nand_x1_sg U7151 ( .A(n1941), .B(n1942), .X(n1940) );
  nand_x1_sg U7152 ( .A(n4436), .B(n5544), .X(n5253) );
  nand_x1_sg U7153 ( .A(n4437), .B(n5543), .X(n5252) );
  nand_x1_sg U7154 ( .A(n4436), .B(n5533), .X(n4566) );
  nand_x1_sg U7155 ( .A(n4437), .B(n5532), .X(n4565) );
  nand_x1_sg U7156 ( .A(n4436), .B(n5522), .X(n4524) );
  nand_x1_sg U7157 ( .A(n4437), .B(n5521), .X(n4523) );
  nand_x1_sg U7158 ( .A(n4436), .B(n5511), .X(n4435) );
  nand_x1_sg U7159 ( .A(n4437), .B(n5510), .X(n4434) );
  nand_x1_sg U7160 ( .A(n4436), .B(n5500), .X(n4482) );
  nand_x1_sg U7161 ( .A(n4437), .B(n5499), .X(n4481) );
  nand_x1_sg U7162 ( .A(n4436), .B(n5489), .X(n4694) );
  nand_x1_sg U7163 ( .A(n4437), .B(n5488), .X(n4693) );
  nand_x1_sg U7164 ( .A(n4436), .B(n5478), .X(n4736) );
  nand_x1_sg U7165 ( .A(n4437), .B(n5477), .X(n4735) );
  nand_x1_sg U7166 ( .A(n4436), .B(n5467), .X(n4650) );
  nand_x1_sg U7167 ( .A(n4437), .B(n5466), .X(n4649) );
  nand_x1_sg U7168 ( .A(n4436), .B(n5456), .X(n4608) );
  nand_x1_sg U7169 ( .A(n4437), .B(n5455), .X(n4607) );
  nand_x1_sg U7170 ( .A(n4436), .B(n5445), .X(n4946) );
  nand_x1_sg U7171 ( .A(n4437), .B(n5444), .X(n4945) );
  nand_x1_sg U7172 ( .A(n4436), .B(n5434), .X(n4988) );
  nand_x1_sg U7173 ( .A(n4437), .B(n5433), .X(n4987) );
  nand_x1_sg U7174 ( .A(n4436), .B(n5423), .X(n5174) );
  nand_x1_sg U7175 ( .A(n4437), .B(n5422), .X(n5173) );
  nand_x1_sg U7176 ( .A(n4436), .B(n5412), .X(n5214) );
  nand_x1_sg U7177 ( .A(n4437), .B(n5411), .X(n5213) );
  nand_x1_sg U7178 ( .A(n4436), .B(n5401), .X(n5138) );
  nand_x1_sg U7179 ( .A(n4437), .B(n5400), .X(n5137) );
  nand_x1_sg U7180 ( .A(n4436), .B(n5390), .X(n5102) );
  nand_x1_sg U7181 ( .A(n4437), .B(n5389), .X(n5101) );
  nand_x1_sg U7182 ( .A(n4436), .B(n5379), .X(n4862) );
  nand_x1_sg U7183 ( .A(n4437), .B(n5378), .X(n4861) );
  nand_x1_sg U7184 ( .A(n4436), .B(n5368), .X(n4904) );
  nand_x1_sg U7185 ( .A(n4437), .B(n5367), .X(n4903) );
  nand_x1_sg U7186 ( .A(n4436), .B(n5357), .X(n4778) );
  nand_x1_sg U7187 ( .A(n4437), .B(n5356), .X(n4777) );
  nand_x1_sg U7188 ( .A(n4436), .B(n5346), .X(n4820) );
  nand_x1_sg U7189 ( .A(n4437), .B(n5345), .X(n4819) );
  nand_x1_sg U7190 ( .A(n4437), .B(n5334), .X(n5029) );
  nand_x1_sg U7191 ( .A(n4436), .B(n5335), .X(n5030) );
  nor_x1_sg U7192 ( .A(n9122), .B(n882), .X(n873) );
  nand_x1_sg U7193 ( .A(n7395), .B(\i_im[7][0] ), .X(n891) );
  nor_x1_sg U7194 ( .A(n875), .B(n876), .X(n874) );
  nor_x1_sg U7195 ( .A(n9123), .B(n916), .X(n910) );
  nand_x1_sg U7196 ( .A(n7394), .B(\i_im[7][1] ), .X(n925) );
  nor_x1_sg U7197 ( .A(n912), .B(n913), .X(n911) );
  nor_x1_sg U7198 ( .A(n9124), .B(n949), .X(n943) );
  nand_x1_sg U7199 ( .A(n4186), .B(\i_im[7][2] ), .X(n958) );
  nor_x1_sg U7200 ( .A(n945), .B(n946), .X(n944) );
  nor_x1_sg U7201 ( .A(n9125), .B(n982), .X(n976) );
  nand_x1_sg U7202 ( .A(n7395), .B(\i_im[7][3] ), .X(n991) );
  nor_x1_sg U7203 ( .A(n9126), .B(n1015), .X(n1009) );
  nand_x1_sg U7204 ( .A(n7394), .B(\i_im[7][4] ), .X(n1024) );
  nor_x1_sg U7205 ( .A(n9127), .B(n1051), .X(n1045) );
  nand_x1_sg U7206 ( .A(n4186), .B(\i_im[7][5] ), .X(n1060) );
  nor_x1_sg U7207 ( .A(n1047), .B(n1048), .X(n1046) );
  nor_x1_sg U7208 ( .A(n9128), .B(n1084), .X(n1078) );
  nand_x1_sg U7209 ( .A(n7395), .B(\i_im[7][6] ), .X(n1093) );
  nor_x1_sg U7210 ( .A(n1080), .B(n1081), .X(n1079) );
  nor_x1_sg U7211 ( .A(n9129), .B(n1117), .X(n1111) );
  nand_x1_sg U7212 ( .A(n7394), .B(\i_im[7][7] ), .X(n1126) );
  nor_x1_sg U7213 ( .A(n9130), .B(n1150), .X(n1144) );
  nand_x1_sg U7214 ( .A(n4186), .B(\i_im[7][8] ), .X(n1159) );
  nor_x1_sg U7215 ( .A(n9131), .B(n1183), .X(n1177) );
  nand_x1_sg U7216 ( .A(n7395), .B(\i_im[7][9] ), .X(n1192) );
  nor_x1_sg U7217 ( .A(n1179), .B(n1180), .X(n1178) );
  nor_x1_sg U7218 ( .A(n9132), .B(n1221), .X(n1215) );
  nand_x1_sg U7219 ( .A(n7394), .B(\i_im[7][10] ), .X(n1230) );
  nor_x1_sg U7220 ( .A(n9133), .B(n1254), .X(n1248) );
  nand_x1_sg U7221 ( .A(n4186), .B(\i_im[7][11] ), .X(n1263) );
  nor_x1_sg U7222 ( .A(n9134), .B(n1287), .X(n1281) );
  nand_x1_sg U7223 ( .A(n7395), .B(\i_im[7][12] ), .X(n1296) );
  nor_x1_sg U7224 ( .A(n1283), .B(n1284), .X(n1282) );
  nor_x1_sg U7225 ( .A(n9135), .B(n1320), .X(n1314) );
  nand_x1_sg U7226 ( .A(n7394), .B(\i_im[7][13] ), .X(n1329) );
  nor_x1_sg U7227 ( .A(n1316), .B(n1317), .X(n1315) );
  nor_x1_sg U7228 ( .A(n9136), .B(n1353), .X(n1347) );
  nand_x1_sg U7229 ( .A(n4186), .B(\i_im[7][14] ), .X(n1362) );
  nor_x1_sg U7230 ( .A(n9137), .B(n1389), .X(n1383) );
  nand_x1_sg U7231 ( .A(n7395), .B(\i_im[7][15] ), .X(n1398) );
  nor_x1_sg U7232 ( .A(n9138), .B(n1422), .X(n1416) );
  nand_x1_sg U7233 ( .A(n7394), .B(\i_im[7][16] ), .X(n1431) );
  nor_x1_sg U7234 ( .A(n9139), .B(n1455), .X(n1449) );
  nand_x1_sg U7235 ( .A(n4186), .B(\i_im[7][17] ), .X(n1464) );
  nor_x1_sg U7236 ( .A(n9140), .B(n1488), .X(n1482) );
  nand_x1_sg U7237 ( .A(n7395), .B(\i_im[7][18] ), .X(n1497) );
  nor_x1_sg U7238 ( .A(n1484), .B(n1485), .X(n1483) );
  nor_x1_sg U7239 ( .A(n9141), .B(n1524), .X(n1518) );
  nand_x1_sg U7240 ( .A(n7394), .B(\i_im[7][19] ), .X(n1533) );
  nand_x1_sg U7241 ( .A(n1584), .B(n1585), .X(n1583) );
  nand_x1_sg U7242 ( .A(n1682), .B(n1683), .X(n1681) );
  nor_x1_sg U7243 ( .A(n9070), .B(n1798), .X(n1797) );
  nand_x1_sg U7244 ( .A(n1748), .B(n1749), .X(n1747) );
  nand_x1_sg U7245 ( .A(n1855), .B(n1856), .X(n1854) );
  nand_x1_sg U7246 ( .A(n1898), .B(n1899), .X(n1897) );
  inv_x1_sg U7247 ( .A(n2068), .X(n9056) );
  nand_x1_sg U7248 ( .A(n7375), .B(n5247), .X(n5245) );
  nand_x1_sg U7249 ( .A(n5248), .B(n5249), .X(n5247) );
  nand_x1_sg U7250 ( .A(n7430), .B(n5539), .X(n5246) );
  nand_x1_sg U7251 ( .A(n7439), .B(n5538), .X(n5234) );
  nand_x1_sg U7252 ( .A(n7441), .B(n5541), .X(n5235) );
  nand_x1_sg U7253 ( .A(n7437), .B(n5542), .X(n5238) );
  nand_x1_sg U7254 ( .A(n7375), .B(n4560), .X(n4558) );
  nand_x1_sg U7255 ( .A(n4561), .B(n4562), .X(n4560) );
  nand_x1_sg U7256 ( .A(n7431), .B(n5528), .X(n4559) );
  nand_x1_sg U7257 ( .A(n7439), .B(n5527), .X(n4550) );
  nand_x1_sg U7258 ( .A(n7441), .B(n5530), .X(n4551) );
  nand_x1_sg U7259 ( .A(n7437), .B(n5531), .X(n4553) );
  nand_x1_sg U7260 ( .A(n7375), .B(n4518), .X(n4516) );
  nand_x1_sg U7261 ( .A(n4519), .B(n4520), .X(n4518) );
  nand_x1_sg U7262 ( .A(n4428), .B(n5517), .X(n4517) );
  nand_x1_sg U7263 ( .A(n7439), .B(n5516), .X(n4508) );
  nand_x1_sg U7264 ( .A(n7441), .B(n5519), .X(n4509) );
  nand_x1_sg U7265 ( .A(n7437), .B(n5520), .X(n4511) );
  nand_x1_sg U7266 ( .A(n7375), .B(n4429), .X(n4426) );
  nand_x1_sg U7267 ( .A(n4430), .B(n4431), .X(n4429) );
  nand_x1_sg U7268 ( .A(n7431), .B(n5506), .X(n4427) );
  nand_x1_sg U7269 ( .A(n7439), .B(n5505), .X(n4413) );
  nand_x1_sg U7270 ( .A(n7441), .B(n5508), .X(n4414) );
  nand_x1_sg U7271 ( .A(n7437), .B(n5509), .X(n4418) );
  nand_x1_sg U7272 ( .A(n7375), .B(n4476), .X(n4474) );
  nand_x1_sg U7273 ( .A(n4477), .B(n4478), .X(n4476) );
  nand_x1_sg U7274 ( .A(n7430), .B(n5495), .X(n4475) );
  nand_x1_sg U7275 ( .A(n7439), .B(n5494), .X(n4466) );
  nand_x1_sg U7276 ( .A(n7441), .B(n5497), .X(n4467) );
  nand_x1_sg U7277 ( .A(n7437), .B(n5498), .X(n4469) );
  nand_x1_sg U7278 ( .A(n7375), .B(n4688), .X(n4686) );
  nand_x1_sg U7279 ( .A(n4689), .B(n4690), .X(n4688) );
  nand_x1_sg U7280 ( .A(n7431), .B(n5484), .X(n4687) );
  nand_x1_sg U7281 ( .A(n7439), .B(n5483), .X(n4678) );
  nand_x1_sg U7282 ( .A(n7441), .B(n5486), .X(n4679) );
  nand_x1_sg U7283 ( .A(n7437), .B(n5487), .X(n4681) );
  nand_x1_sg U7284 ( .A(n7375), .B(n4730), .X(n4728) );
  nand_x1_sg U7285 ( .A(n4731), .B(n4732), .X(n4730) );
  nand_x1_sg U7286 ( .A(n7430), .B(n5473), .X(n4729) );
  nand_x1_sg U7287 ( .A(n7439), .B(n5472), .X(n4720) );
  nand_x1_sg U7288 ( .A(n7441), .B(n5475), .X(n4721) );
  nand_x1_sg U7289 ( .A(n7437), .B(n5476), .X(n4723) );
  nand_x1_sg U7290 ( .A(n7375), .B(n4644), .X(n4642) );
  nand_x1_sg U7291 ( .A(n4645), .B(n4646), .X(n4644) );
  nand_x1_sg U7292 ( .A(n4428), .B(n5462), .X(n4643) );
  nand_x1_sg U7293 ( .A(n7439), .B(n5461), .X(n4634) );
  nand_x1_sg U7294 ( .A(n7441), .B(n5464), .X(n4635) );
  nand_x1_sg U7295 ( .A(n7437), .B(n5465), .X(n4637) );
  nand_x1_sg U7296 ( .A(n7375), .B(n4602), .X(n4600) );
  nand_x1_sg U7297 ( .A(n4603), .B(n4604), .X(n4602) );
  nand_x1_sg U7298 ( .A(n7430), .B(n5451), .X(n4601) );
  nand_x1_sg U7299 ( .A(n7439), .B(n5450), .X(n4592) );
  nand_x1_sg U7300 ( .A(n7441), .B(n5453), .X(n4593) );
  nand_x1_sg U7301 ( .A(n7437), .B(n5454), .X(n4595) );
  nand_x1_sg U7302 ( .A(n7375), .B(n4940), .X(n4938) );
  nand_x1_sg U7303 ( .A(n4941), .B(n4942), .X(n4940) );
  nand_x1_sg U7304 ( .A(n7431), .B(n5440), .X(n4939) );
  nand_x1_sg U7305 ( .A(n7439), .B(n5439), .X(n4930) );
  nand_x1_sg U7306 ( .A(n7441), .B(n5442), .X(n4931) );
  nand_x1_sg U7307 ( .A(n7437), .B(n5443), .X(n4933) );
  nand_x1_sg U7308 ( .A(n7375), .B(n4982), .X(n4980) );
  nand_x1_sg U7309 ( .A(n4983), .B(n4984), .X(n4982) );
  nand_x1_sg U7310 ( .A(n7430), .B(n5429), .X(n4981) );
  nand_x1_sg U7311 ( .A(n7439), .B(n5428), .X(n4972) );
  nand_x1_sg U7312 ( .A(n7441), .B(n5431), .X(n4973) );
  nand_x1_sg U7313 ( .A(n7437), .B(n5432), .X(n4975) );
  nand_x1_sg U7314 ( .A(n7375), .B(n5168), .X(n5166) );
  nand_x1_sg U7315 ( .A(n5169), .B(n5170), .X(n5168) );
  nand_x1_sg U7316 ( .A(n4428), .B(n5418), .X(n5167) );
  nand_x1_sg U7317 ( .A(n4416), .B(n5417), .X(n5158) );
  nand_x1_sg U7318 ( .A(n4415), .B(n5420), .X(n5159) );
  nand_x1_sg U7319 ( .A(n4419), .B(n5421), .X(n5161) );
  nand_x1_sg U7320 ( .A(n7375), .B(n5208), .X(n5206) );
  nand_x1_sg U7321 ( .A(n5209), .B(n5210), .X(n5208) );
  nand_x1_sg U7322 ( .A(n7431), .B(n5407), .X(n5207) );
  nand_x1_sg U7323 ( .A(n7439), .B(n5406), .X(n5198) );
  nand_x1_sg U7324 ( .A(n7441), .B(n5409), .X(n5199) );
  nand_x1_sg U7325 ( .A(n7437), .B(n5410), .X(n5201) );
  nand_x1_sg U7326 ( .A(n6380), .B(n5132), .X(n5130) );
  nand_x1_sg U7327 ( .A(n5133), .B(n5134), .X(n5132) );
  nand_x1_sg U7328 ( .A(n7430), .B(n5396), .X(n5131) );
  nand_x1_sg U7329 ( .A(n7439), .B(n5395), .X(n5122) );
  nand_x1_sg U7330 ( .A(n7441), .B(n5398), .X(n5123) );
  nand_x1_sg U7331 ( .A(n7437), .B(n5399), .X(n5125) );
  nand_x1_sg U7332 ( .A(n7375), .B(n5096), .X(n5094) );
  nand_x1_sg U7333 ( .A(n5097), .B(n5098), .X(n5096) );
  nand_x1_sg U7334 ( .A(n7431), .B(n5385), .X(n5095) );
  nand_x1_sg U7335 ( .A(n7439), .B(n5384), .X(n5086) );
  nand_x1_sg U7336 ( .A(n7441), .B(n5387), .X(n5087) );
  nand_x1_sg U7337 ( .A(n7437), .B(n5388), .X(n5089) );
  nand_x1_sg U7338 ( .A(n7375), .B(n4856), .X(n4854) );
  nand_x1_sg U7339 ( .A(n4857), .B(n4858), .X(n4856) );
  nand_x1_sg U7340 ( .A(n7430), .B(n5374), .X(n4855) );
  nand_x1_sg U7341 ( .A(n7439), .B(n5373), .X(n4846) );
  nand_x1_sg U7342 ( .A(n7441), .B(n5376), .X(n4847) );
  nand_x1_sg U7343 ( .A(n7437), .B(n5377), .X(n4849) );
  nand_x1_sg U7344 ( .A(n7375), .B(n4898), .X(n4896) );
  nand_x1_sg U7345 ( .A(n4899), .B(n4900), .X(n4898) );
  nand_x1_sg U7346 ( .A(n4428), .B(n5363), .X(n4897) );
  nand_x1_sg U7347 ( .A(n7439), .B(n5362), .X(n4888) );
  nand_x1_sg U7348 ( .A(n7441), .B(n5365), .X(n4889) );
  nand_x1_sg U7349 ( .A(n7437), .B(n5366), .X(n4891) );
  nand_x1_sg U7350 ( .A(n7375), .B(n4772), .X(n4770) );
  nand_x1_sg U7351 ( .A(n4773), .B(n4774), .X(n4772) );
  nand_x1_sg U7352 ( .A(n4428), .B(n5352), .X(n4771) );
  nand_x1_sg U7353 ( .A(n7439), .B(n5351), .X(n4762) );
  nand_x1_sg U7354 ( .A(n7441), .B(n5354), .X(n4763) );
  nand_x1_sg U7355 ( .A(n7437), .B(n5355), .X(n4765) );
  nand_x1_sg U7356 ( .A(n7375), .B(n4814), .X(n4812) );
  nand_x1_sg U7357 ( .A(n4815), .B(n4816), .X(n4814) );
  nand_x1_sg U7358 ( .A(n7431), .B(n5341), .X(n4813) );
  nand_x1_sg U7359 ( .A(n7439), .B(n5340), .X(n4804) );
  nand_x1_sg U7360 ( .A(n7441), .B(n5343), .X(n4805) );
  nand_x1_sg U7361 ( .A(n7437), .B(n5344), .X(n4807) );
  nand_x1_sg U7362 ( .A(n7375), .B(n5024), .X(n5022) );
  nand_x1_sg U7363 ( .A(n5025), .B(n5026), .X(n5024) );
  nand_x1_sg U7364 ( .A(n4428), .B(n5330), .X(n5023) );
  nand_x1_sg U7365 ( .A(n7439), .B(n5329), .X(n5014) );
  nand_x1_sg U7366 ( .A(n7441), .B(n5332), .X(n5015) );
  nand_x1_sg U7367 ( .A(n7437), .B(n5333), .X(n5017) );
  nand_x1_sg U7368 ( .A(\i_im[8][0] ), .B(n7377), .X(n857) );
  nand_x1_sg U7369 ( .A(\i_im[9][0] ), .B(n859), .X(n856) );
  nand_x1_sg U7370 ( .A(\i_im[14][0] ), .B(n7379), .X(n861) );
  nand_x1_sg U7371 ( .A(n7398), .B(n872), .X(n869) );
  nand_x1_sg U7372 ( .A(n873), .B(n874), .X(n872) );
  nand_x1_sg U7373 ( .A(\i_im[10][0] ), .B(n7397), .X(n893) );
  nand_x1_sg U7374 ( .A(\i_im[15][0] ), .B(n7400), .X(n892) );
  nand_x1_sg U7375 ( .A(\i_im[8][1] ), .B(n7377), .X(n900) );
  nand_x1_sg U7376 ( .A(\i_im[9][1] ), .B(n859), .X(n899) );
  nand_x1_sg U7377 ( .A(\i_im[14][1] ), .B(n7379), .X(n902) );
  nand_x1_sg U7378 ( .A(n7398), .B(n909), .X(n907) );
  nand_x1_sg U7379 ( .A(n910), .B(n911), .X(n909) );
  nand_x1_sg U7380 ( .A(\i_im[10][1] ), .B(n7396), .X(n927) );
  nand_x1_sg U7381 ( .A(\i_im[15][1] ), .B(n7400), .X(n926) );
  nand_x1_sg U7382 ( .A(\i_im[8][2] ), .B(n7377), .X(n933) );
  nand_x1_sg U7383 ( .A(\i_im[9][2] ), .B(n859), .X(n932) );
  nand_x1_sg U7384 ( .A(\i_im[14][2] ), .B(n7379), .X(n935) );
  nand_x1_sg U7385 ( .A(n7398), .B(n942), .X(n940) );
  nand_x1_sg U7386 ( .A(n943), .B(n944), .X(n942) );
  nand_x1_sg U7387 ( .A(\i_im[10][2] ), .B(n894), .X(n960) );
  nand_x1_sg U7388 ( .A(\i_im[15][2] ), .B(n7400), .X(n959) );
  nand_x1_sg U7389 ( .A(\i_im[8][3] ), .B(n7377), .X(n966) );
  nand_x1_sg U7390 ( .A(\i_im[9][3] ), .B(n859), .X(n965) );
  nand_x1_sg U7391 ( .A(\i_im[14][3] ), .B(n7379), .X(n968) );
  nand_x1_sg U7392 ( .A(n7398), .B(n975), .X(n973) );
  nand_x1_sg U7393 ( .A(n976), .B(n977), .X(n975) );
  nand_x1_sg U7394 ( .A(\i_im[10][3] ), .B(n7397), .X(n993) );
  nand_x1_sg U7395 ( .A(\i_im[15][3] ), .B(n7400), .X(n992) );
  nand_x1_sg U7396 ( .A(\i_im[8][4] ), .B(n7377), .X(n999) );
  nand_x1_sg U7397 ( .A(\i_im[9][4] ), .B(n859), .X(n998) );
  nand_x1_sg U7398 ( .A(\i_im[14][4] ), .B(n7379), .X(n1001) );
  nand_x1_sg U7399 ( .A(n7398), .B(n1008), .X(n1006) );
  nand_x1_sg U7400 ( .A(n1009), .B(n1010), .X(n1008) );
  nand_x1_sg U7401 ( .A(\i_im[10][4] ), .B(n7396), .X(n1026) );
  nand_x1_sg U7402 ( .A(\i_im[15][4] ), .B(n7400), .X(n1025) );
  nand_x1_sg U7403 ( .A(\i_im[8][5] ), .B(n7377), .X(n1035) );
  nand_x1_sg U7404 ( .A(\i_im[9][5] ), .B(n859), .X(n1034) );
  nand_x1_sg U7405 ( .A(\i_im[14][5] ), .B(n7379), .X(n1037) );
  nand_x1_sg U7406 ( .A(n7398), .B(n1044), .X(n1042) );
  nand_x1_sg U7407 ( .A(n1045), .B(n1046), .X(n1044) );
  nand_x1_sg U7408 ( .A(\i_im[10][5] ), .B(n894), .X(n1062) );
  nand_x1_sg U7409 ( .A(\i_im[15][5] ), .B(n7400), .X(n1061) );
  nand_x1_sg U7410 ( .A(\i_im[8][6] ), .B(n7377), .X(n1068) );
  nand_x1_sg U7411 ( .A(\i_im[9][6] ), .B(n859), .X(n1067) );
  nand_x1_sg U7412 ( .A(\i_im[14][6] ), .B(n7379), .X(n1070) );
  nand_x1_sg U7413 ( .A(n7398), .B(n1077), .X(n1075) );
  nand_x1_sg U7414 ( .A(n1078), .B(n1079), .X(n1077) );
  nand_x1_sg U7415 ( .A(\i_im[10][6] ), .B(n7397), .X(n1095) );
  nand_x1_sg U7416 ( .A(\i_im[15][6] ), .B(n7400), .X(n1094) );
  nand_x1_sg U7417 ( .A(\i_im[8][7] ), .B(n7377), .X(n1101) );
  nand_x1_sg U7418 ( .A(\i_im[9][7] ), .B(n859), .X(n1100) );
  nand_x1_sg U7419 ( .A(\i_im[14][7] ), .B(n7379), .X(n1103) );
  nand_x1_sg U7420 ( .A(n7398), .B(n1110), .X(n1108) );
  nand_x1_sg U7421 ( .A(n1111), .B(n1112), .X(n1110) );
  nand_x1_sg U7422 ( .A(\i_im[10][7] ), .B(n7396), .X(n1128) );
  nand_x1_sg U7423 ( .A(\i_im[15][7] ), .B(n4207), .X(n1127) );
  nand_x1_sg U7424 ( .A(\i_im[8][8] ), .B(n7377), .X(n1134) );
  nand_x1_sg U7425 ( .A(\i_im[9][8] ), .B(n859), .X(n1133) );
  nand_x1_sg U7426 ( .A(\i_im[14][8] ), .B(n7379), .X(n1136) );
  nand_x1_sg U7427 ( .A(n6151), .B(n1143), .X(n1141) );
  nand_x1_sg U7428 ( .A(n1144), .B(n1145), .X(n1143) );
  nand_x1_sg U7429 ( .A(\i_im[10][8] ), .B(n894), .X(n1161) );
  nand_x1_sg U7430 ( .A(\i_im[15][8] ), .B(n7400), .X(n1160) );
  nand_x1_sg U7431 ( .A(\i_im[8][9] ), .B(n7377), .X(n1167) );
  nand_x1_sg U7432 ( .A(\i_im[9][9] ), .B(n859), .X(n1166) );
  nand_x1_sg U7433 ( .A(\i_im[14][9] ), .B(n7379), .X(n1169) );
  nand_x1_sg U7434 ( .A(n7398), .B(n1176), .X(n1174) );
  nand_x1_sg U7435 ( .A(n1177), .B(n1178), .X(n1176) );
  nand_x1_sg U7436 ( .A(\i_im[10][9] ), .B(n7397), .X(n1194) );
  nand_x1_sg U7437 ( .A(\i_im[15][9] ), .B(n7400), .X(n1193) );
  nand_x1_sg U7438 ( .A(\i_im[8][10] ), .B(n7377), .X(n1205) );
  nand_x1_sg U7439 ( .A(\i_im[9][10] ), .B(n859), .X(n1204) );
  nand_x1_sg U7440 ( .A(\i_im[14][10] ), .B(n7379), .X(n1207) );
  nand_x1_sg U7441 ( .A(n7398), .B(n1214), .X(n1212) );
  nand_x1_sg U7442 ( .A(n1215), .B(n1216), .X(n1214) );
  nand_x1_sg U7443 ( .A(\i_im[10][10] ), .B(n7396), .X(n1232) );
  nand_x1_sg U7444 ( .A(\i_im[15][10] ), .B(n7400), .X(n1231) );
  nand_x1_sg U7445 ( .A(\i_im[8][11] ), .B(n7377), .X(n1238) );
  nand_x1_sg U7446 ( .A(\i_im[9][11] ), .B(n859), .X(n1237) );
  nand_x1_sg U7447 ( .A(\i_im[14][11] ), .B(n7379), .X(n1240) );
  nand_x1_sg U7448 ( .A(n7398), .B(n1247), .X(n1245) );
  nand_x1_sg U7449 ( .A(n1248), .B(n1249), .X(n1247) );
  nand_x1_sg U7450 ( .A(\i_im[10][11] ), .B(n894), .X(n1265) );
  nand_x1_sg U7451 ( .A(\i_im[15][11] ), .B(n7400), .X(n1264) );
  nand_x1_sg U7452 ( .A(\i_im[8][12] ), .B(n858), .X(n1271) );
  nand_x1_sg U7453 ( .A(\i_im[9][12] ), .B(n859), .X(n1270) );
  nand_x1_sg U7454 ( .A(\i_im[14][12] ), .B(n862), .X(n1273) );
  nand_x1_sg U7455 ( .A(n7398), .B(n1280), .X(n1278) );
  nand_x1_sg U7456 ( .A(n1281), .B(n1282), .X(n1280) );
  nand_x1_sg U7457 ( .A(\i_im[10][12] ), .B(n7397), .X(n1298) );
  nand_x1_sg U7458 ( .A(\i_im[15][12] ), .B(n7400), .X(n1297) );
  nand_x1_sg U7459 ( .A(\i_im[8][13] ), .B(n7377), .X(n1304) );
  nand_x1_sg U7460 ( .A(\i_im[9][13] ), .B(n859), .X(n1303) );
  nand_x1_sg U7461 ( .A(\i_im[14][13] ), .B(n7379), .X(n1306) );
  nand_x1_sg U7462 ( .A(n7398), .B(n1313), .X(n1311) );
  nand_x1_sg U7463 ( .A(n1314), .B(n1315), .X(n1313) );
  nand_x1_sg U7464 ( .A(\i_im[10][13] ), .B(n7396), .X(n1331) );
  nand_x1_sg U7465 ( .A(\i_im[15][13] ), .B(n7400), .X(n1330) );
  nand_x1_sg U7466 ( .A(\i_im[8][14] ), .B(n7377), .X(n1337) );
  nand_x1_sg U7467 ( .A(\i_im[9][14] ), .B(n859), .X(n1336) );
  nand_x1_sg U7468 ( .A(\i_im[14][14] ), .B(n7379), .X(n1339) );
  nand_x1_sg U7469 ( .A(n7398), .B(n1346), .X(n1344) );
  nand_x1_sg U7470 ( .A(n1347), .B(n1348), .X(n1346) );
  nand_x1_sg U7471 ( .A(\i_im[10][14] ), .B(n894), .X(n1364) );
  nand_x1_sg U7472 ( .A(\i_im[15][14] ), .B(n7400), .X(n1363) );
  nand_x1_sg U7473 ( .A(\i_im[8][15] ), .B(n7377), .X(n1373) );
  nand_x1_sg U7474 ( .A(\i_im[9][15] ), .B(n859), .X(n1372) );
  nand_x1_sg U7475 ( .A(\i_im[14][15] ), .B(n7379), .X(n1375) );
  nand_x1_sg U7476 ( .A(n7398), .B(n1382), .X(n1380) );
  nand_x1_sg U7477 ( .A(n1383), .B(n1384), .X(n1382) );
  nand_x1_sg U7478 ( .A(\i_im[10][15] ), .B(n7397), .X(n1400) );
  nand_x1_sg U7479 ( .A(\i_im[15][15] ), .B(n7400), .X(n1399) );
  nand_x1_sg U7480 ( .A(\i_im[8][16] ), .B(n7377), .X(n1406) );
  nand_x1_sg U7481 ( .A(\i_im[9][16] ), .B(n859), .X(n1405) );
  nand_x1_sg U7482 ( .A(\i_im[14][16] ), .B(n7379), .X(n1408) );
  nand_x1_sg U7483 ( .A(n7398), .B(n1415), .X(n1413) );
  nand_x1_sg U7484 ( .A(n1416), .B(n1417), .X(n1415) );
  nand_x1_sg U7485 ( .A(\i_im[10][16] ), .B(n7396), .X(n1433) );
  nand_x1_sg U7486 ( .A(\i_im[15][16] ), .B(n7400), .X(n1432) );
  nand_x1_sg U7487 ( .A(\i_im[8][17] ), .B(n7377), .X(n1439) );
  nand_x1_sg U7488 ( .A(\i_im[9][17] ), .B(n859), .X(n1438) );
  nand_x1_sg U7489 ( .A(\i_im[14][17] ), .B(n7379), .X(n1441) );
  nand_x1_sg U7490 ( .A(n7398), .B(n1448), .X(n1446) );
  nand_x1_sg U7491 ( .A(n1449), .B(n1450), .X(n1448) );
  nand_x1_sg U7492 ( .A(\i_im[10][17] ), .B(n894), .X(n1466) );
  nand_x1_sg U7493 ( .A(\i_im[15][17] ), .B(n7400), .X(n1465) );
  nand_x1_sg U7494 ( .A(\i_im[8][18] ), .B(n7377), .X(n1472) );
  nand_x1_sg U7495 ( .A(\i_im[9][18] ), .B(n859), .X(n1471) );
  nand_x1_sg U7496 ( .A(\i_im[14][18] ), .B(n7379), .X(n1474) );
  nand_x1_sg U7497 ( .A(n7398), .B(n1481), .X(n1479) );
  nand_x1_sg U7498 ( .A(n1482), .B(n1483), .X(n1481) );
  nand_x1_sg U7499 ( .A(\i_im[10][18] ), .B(n7397), .X(n1499) );
  nand_x1_sg U7500 ( .A(\i_im[15][18] ), .B(n7400), .X(n1498) );
  nand_x1_sg U7501 ( .A(\i_im[8][19] ), .B(n7377), .X(n1505) );
  nand_x1_sg U7502 ( .A(\i_im[9][19] ), .B(n859), .X(n1504) );
  nand_x1_sg U7503 ( .A(\i_im[14][19] ), .B(n7379), .X(n1507) );
  nand_x1_sg U7504 ( .A(n7398), .B(n1517), .X(n1515) );
  nand_x1_sg U7505 ( .A(n1518), .B(n1519), .X(n1517) );
  nand_x1_sg U7506 ( .A(\i_im[10][19] ), .B(n7396), .X(n1535) );
  nand_x1_sg U7507 ( .A(\i_im[15][19] ), .B(n7400), .X(n1534) );
  nand_x1_sg U7508 ( .A(n1633), .B(n1634), .X(n1632) );
  nand_x1_sg U7509 ( .A(n1697), .B(n1698), .X(n1696) );
  nand_x1_sg U7510 ( .A(n1794), .B(n1795), .X(n1745) );
  nand_x1_sg U7511 ( .A(n1796), .B(n1797), .X(n1795) );
  nand_x1_sg U7512 ( .A(n1945), .B(n1946), .X(n1944) );
  nor_x1_sg U7513 ( .A(n9061), .B(n2052), .X(n2051) );
  nand_x1_sg U7514 ( .A(n2032), .B(n2033), .X(n2031) );
  inv_x2_sg U7515 ( .A(n3097), .X(n5993) );
  nor_x1_sg U7516 ( .A(n7540), .B(n7321), .X(n3097) );
  nor_x1_sg U7517 ( .A(n5243), .B(n5244), .X(n5230) );
  nand_x1_sg U7518 ( .A(n7426), .B(n5540), .X(n5265) );
  nor_x1_sg U7519 ( .A(n5232), .B(n5233), .X(n5231) );
  nor_x1_sg U7520 ( .A(n5239), .B(n5240), .X(n5237) );
  nor_x1_sg U7521 ( .A(n4556), .B(n4557), .X(n4546) );
  nand_x1_sg U7522 ( .A(n7426), .B(n5529), .X(n4578) );
  nor_x1_sg U7523 ( .A(n4548), .B(n4549), .X(n4547) );
  nor_x1_sg U7524 ( .A(n4554), .B(n4555), .X(n4552) );
  nor_x1_sg U7525 ( .A(n4514), .B(n4515), .X(n4504) );
  nand_x1_sg U7526 ( .A(n7426), .B(n5518), .X(n4536) );
  nor_x1_sg U7527 ( .A(n4506), .B(n4507), .X(n4505) );
  nor_x1_sg U7528 ( .A(n4512), .B(n4513), .X(n4510) );
  nor_x1_sg U7529 ( .A(n4424), .B(n4425), .X(n4409) );
  nand_x1_sg U7530 ( .A(n7426), .B(n5507), .X(n4450) );
  nor_x1_sg U7531 ( .A(n4411), .B(n4412), .X(n4410) );
  nor_x1_sg U7532 ( .A(n4420), .B(n4421), .X(n4417) );
  nor_x1_sg U7533 ( .A(n4472), .B(n4473), .X(n4462) );
  nand_x1_sg U7534 ( .A(n7426), .B(n5496), .X(n4494) );
  nor_x1_sg U7535 ( .A(n4464), .B(n4465), .X(n4463) );
  nor_x1_sg U7536 ( .A(n4470), .B(n4471), .X(n4468) );
  nor_x1_sg U7537 ( .A(n4684), .B(n4685), .X(n4674) );
  nand_x1_sg U7538 ( .A(n7426), .B(n5485), .X(n4706) );
  nor_x1_sg U7539 ( .A(n4676), .B(n4677), .X(n4675) );
  nor_x1_sg U7540 ( .A(n4682), .B(n4683), .X(n4680) );
  nor_x1_sg U7541 ( .A(n4726), .B(n4727), .X(n4716) );
  nand_x1_sg U7542 ( .A(n7426), .B(n5474), .X(n4748) );
  nor_x1_sg U7543 ( .A(n4718), .B(n4719), .X(n4717) );
  nor_x1_sg U7544 ( .A(n4724), .B(n4725), .X(n4722) );
  nor_x1_sg U7545 ( .A(n4640), .B(n4641), .X(n4630) );
  nand_x1_sg U7546 ( .A(n7426), .B(n5463), .X(n4662) );
  nor_x1_sg U7547 ( .A(n4632), .B(n4633), .X(n4631) );
  nor_x1_sg U7548 ( .A(n4638), .B(n4639), .X(n4636) );
  nor_x1_sg U7549 ( .A(n4598), .B(n4599), .X(n4588) );
  nand_x1_sg U7550 ( .A(n7426), .B(n5452), .X(n4620) );
  nor_x1_sg U7551 ( .A(n4590), .B(n4591), .X(n4589) );
  nor_x1_sg U7552 ( .A(n4596), .B(n4597), .X(n4594) );
  nor_x1_sg U7553 ( .A(n4936), .B(n4937), .X(n4926) );
  nand_x1_sg U7554 ( .A(n7426), .B(n5441), .X(n4958) );
  nor_x1_sg U7555 ( .A(n4928), .B(n4929), .X(n4927) );
  nor_x1_sg U7556 ( .A(n4934), .B(n4935), .X(n4932) );
  nor_x1_sg U7557 ( .A(n4978), .B(n4979), .X(n4968) );
  nand_x1_sg U7558 ( .A(n7426), .B(n5430), .X(n5000) );
  nor_x1_sg U7559 ( .A(n4970), .B(n4971), .X(n4969) );
  nor_x1_sg U7560 ( .A(n4976), .B(n4977), .X(n4974) );
  nor_x1_sg U7561 ( .A(n5164), .B(n5165), .X(n5154) );
  nand_x1_sg U7562 ( .A(n4451), .B(n5419), .X(n5186) );
  nor_x1_sg U7563 ( .A(n5156), .B(n5157), .X(n5155) );
  nor_x1_sg U7564 ( .A(n5162), .B(n5163), .X(n5160) );
  nor_x1_sg U7565 ( .A(n5204), .B(n5205), .X(n5194) );
  nand_x1_sg U7566 ( .A(n7426), .B(n5408), .X(n5226) );
  nor_x1_sg U7567 ( .A(n5196), .B(n5197), .X(n5195) );
  nor_x1_sg U7568 ( .A(n5202), .B(n5203), .X(n5200) );
  nor_x1_sg U7569 ( .A(n5128), .B(n5129), .X(n5118) );
  nand_x1_sg U7570 ( .A(n7426), .B(n5397), .X(n5150) );
  nor_x1_sg U7571 ( .A(n5120), .B(n5121), .X(n5119) );
  nor_x1_sg U7572 ( .A(n5126), .B(n5127), .X(n5124) );
  nor_x1_sg U7573 ( .A(n5092), .B(n5093), .X(n5082) );
  nand_x1_sg U7574 ( .A(n7426), .B(n5386), .X(n5114) );
  nor_x1_sg U7575 ( .A(n5084), .B(n5085), .X(n5083) );
  nor_x1_sg U7576 ( .A(n5090), .B(n5091), .X(n5088) );
  nor_x1_sg U7577 ( .A(n4852), .B(n4853), .X(n4842) );
  nand_x1_sg U7578 ( .A(n7426), .B(n5375), .X(n4874) );
  nor_x1_sg U7579 ( .A(n4844), .B(n4845), .X(n4843) );
  nor_x1_sg U7580 ( .A(n4850), .B(n4851), .X(n4848) );
  nor_x1_sg U7581 ( .A(n4894), .B(n4895), .X(n4884) );
  nand_x1_sg U7582 ( .A(n7426), .B(n5364), .X(n4916) );
  nor_x1_sg U7583 ( .A(n4886), .B(n4887), .X(n4885) );
  nor_x1_sg U7584 ( .A(n4892), .B(n4893), .X(n4890) );
  nor_x1_sg U7585 ( .A(n4768), .B(n4769), .X(n4758) );
  nand_x1_sg U7586 ( .A(n7426), .B(n5353), .X(n4790) );
  nor_x1_sg U7587 ( .A(n4760), .B(n4761), .X(n4759) );
  nor_x1_sg U7588 ( .A(n4766), .B(n4767), .X(n4764) );
  nor_x1_sg U7589 ( .A(n4810), .B(n4811), .X(n4800) );
  nand_x1_sg U7590 ( .A(n7426), .B(n5342), .X(n4832) );
  nor_x1_sg U7591 ( .A(n4802), .B(n4803), .X(n4801) );
  nor_x1_sg U7592 ( .A(n4808), .B(n4809), .X(n4806) );
  nor_x1_sg U7593 ( .A(n5020), .B(n5021), .X(n5010) );
  nand_x1_sg U7594 ( .A(n7426), .B(n5331), .X(n5042) );
  nor_x1_sg U7595 ( .A(n5012), .B(n5013), .X(n5011) );
  nor_x1_sg U7596 ( .A(n5018), .B(n5019), .X(n5016) );
  nor_x1_sg U7597 ( .A(n7374), .B(n7372), .X(n1365) );
  nor_x1_sg U7598 ( .A(n7370), .B(n1367), .X(n1366) );
  nand_x1_sg U7599 ( .A(n1999), .B(n2000), .X(n1998) );
  nand_x1_sg U7600 ( .A(n2014), .B(n2015), .X(n2013) );
  nand_x1_sg U7601 ( .A(n2029), .B(n2030), .X(n2028) );
  nand_x1_sg U7602 ( .A(n2050), .B(n2051), .X(n2049) );
  nand_x1_sg U7603 ( .A(n4099), .B(n9206), .X(n5080) );
  inv_x1_sg U7604 ( .A(n3098), .X(n9206) );
  nand_x1_sg U7605 ( .A(n5190), .B(n6156), .X(n5189) );
  nand_x1_sg U7606 ( .A(n7520), .B(n1995), .X(n1994) );
  nand_x1_sg U7607 ( .A(n1996), .B(n1997), .X(n1995) );
  nand_x1_sg U7608 ( .A(n4186), .B(n7398), .X(n4185) );
  nand_x1_sg U7609 ( .A(n4182), .B(n4192), .X(n4191) );
  nand_x1_sg U7610 ( .A(n9199), .B(n5276), .X(n5275) );
  inv_x1_sg U7611 ( .A(n5277), .X(n9199) );
  inv_x1_sg U7612 ( .A(\update_mask_0/reg_out[15][19] ), .X(n6009) );
  inv_x1_sg U7613 ( .A(\update_mask_0/reg_out[14][19] ), .X(n5999) );
  inv_x1_sg U7614 ( .A(\update_mask_0/reg_out[13][19] ), .X(n6045) );
  inv_x1_sg U7615 ( .A(\update_mask_0/reg_out[12][19] ), .X(n7034) );
  inv_x1_sg U7616 ( .A(\update_mask_0/reg_out[11][19] ), .X(n6007) );
  inv_x1_sg U7617 ( .A(\update_mask_0/reg_out[9][19] ), .X(n6005) );
  inv_x1_sg U7618 ( .A(\update_mask_0/reg_out[8][19] ), .X(n5997) );
  inv_x1_sg U7619 ( .A(\update_mask_0/reg_out[7][19] ), .X(n6043) );
  inv_x1_sg U7620 ( .A(\update_mask_0/reg_out[5][19] ), .X(n6041) );
  inv_x2_sg U7621 ( .A(\update_mask_0/reg_out[5][16] ), .X(n9032) );
  inv_x1_sg U7622 ( .A(\update_mask_0/reg_out[4][19] ), .X(n7032) );
  inv_x2_sg U7623 ( .A(\update_mask_0/reg_out[4][16] ), .X(n9036) );
  inv_x1_sg U7624 ( .A(\update_mask_0/reg_out[3][19] ), .X(n6003) );
  inv_x2_sg U7625 ( .A(\update_mask_0/reg_out[3][16] ), .X(n9040) );
  inv_x1_sg U7626 ( .A(\update_mask_0/reg_out[2][19] ), .X(n5995) );
  inv_x2_sg U7627 ( .A(\update_mask_0/reg_out[2][16] ), .X(n9044) );
  inv_x2_sg U7628 ( .A(\update_mask_0/reg_out[1][17] ), .X(n9048) );
  inv_x2_sg U7629 ( .A(\update_mask_0/reg_out[0][17] ), .X(n9052) );
  inv_x1_sg U7630 ( .A(\update_mask_0/reg_i_mask [31]), .X(n7030) );
  inv_x1_sg U7631 ( .A(\update_mask_0/reg_i_mask [23]), .X(n7028) );
  inv_x1_sg U7632 ( .A(\update_mask_0/reg_i_mask [15]), .X(n7026) );
  inv_x1_sg U7633 ( .A(\update_mask_0/reg_i_mask [7]), .X(n7024) );
  inv_x1_sg U7634 ( .A(n9567), .X(n6902) );
  inv_x1_sg U7635 ( .A(n9566), .X(n6900) );
  inv_x1_sg U7636 ( .A(n9565), .X(n6898) );
  inv_x1_sg U7637 ( .A(n9564), .X(n6896) );
  inv_x1_sg U7638 ( .A(n9563), .X(n6894) );
  inv_x1_sg U7639 ( .A(n9562), .X(n6892) );
  inv_x1_sg U7640 ( .A(n9561), .X(n6890) );
  inv_x1_sg U7641 ( .A(n9560), .X(n6888) );
  inv_x1_sg U7642 ( .A(n9559), .X(n6886) );
  inv_x1_sg U7643 ( .A(n9558), .X(n6884) );
  inv_x1_sg U7644 ( .A(n9557), .X(n6882) );
  inv_x1_sg U7645 ( .A(n9556), .X(n6880) );
  inv_x1_sg U7646 ( .A(n9555), .X(n6878) );
  inv_x1_sg U7647 ( .A(n9554), .X(n6876) );
  inv_x1_sg U7648 ( .A(n9553), .X(n6874) );
  inv_x1_sg U7649 ( .A(n9552), .X(n6872) );
  inv_x1_sg U7650 ( .A(n9551), .X(n6870) );
  inv_x1_sg U7651 ( .A(n9550), .X(n6868) );
  inv_x1_sg U7652 ( .A(n9549), .X(n6866) );
  inv_x1_sg U7653 ( .A(n9548), .X(n6864) );
  inv_x1_sg U7654 ( .A(n9547), .X(n6782) );
  inv_x1_sg U7655 ( .A(n9546), .X(n6780) );
  inv_x1_sg U7656 ( .A(n9545), .X(n6778) );
  inv_x1_sg U7657 ( .A(n9544), .X(n6776) );
  inv_x1_sg U7658 ( .A(n9543), .X(n6774) );
  inv_x1_sg U7659 ( .A(n9542), .X(n6772) );
  inv_x1_sg U7660 ( .A(n9541), .X(n6770) );
  inv_x1_sg U7661 ( .A(n9540), .X(n6768) );
  inv_x1_sg U7662 ( .A(n9539), .X(n6766) );
  inv_x1_sg U7663 ( .A(n9538), .X(n6764) );
  inv_x1_sg U7664 ( .A(n9537), .X(n6762) );
  inv_x1_sg U7665 ( .A(n9536), .X(n6760) );
  inv_x1_sg U7666 ( .A(n9535), .X(n6758) );
  inv_x1_sg U7667 ( .A(n9534), .X(n6756) );
  inv_x1_sg U7668 ( .A(n9533), .X(n6754) );
  inv_x1_sg U7669 ( .A(n9532), .X(n6752) );
  inv_x1_sg U7670 ( .A(n9531), .X(n6750) );
  inv_x1_sg U7671 ( .A(n9530), .X(n6748) );
  inv_x1_sg U7672 ( .A(n9529), .X(n6746) );
  inv_x1_sg U7673 ( .A(n9528), .X(n6744) );
  inv_x1_sg U7674 ( .A(n9527), .X(n6862) );
  inv_x1_sg U7675 ( .A(n9526), .X(n6860) );
  inv_x1_sg U7676 ( .A(n9525), .X(n6858) );
  inv_x1_sg U7677 ( .A(n9524), .X(n6856) );
  inv_x1_sg U7678 ( .A(n9523), .X(n6854) );
  inv_x1_sg U7679 ( .A(n9522), .X(n6852) );
  inv_x1_sg U7680 ( .A(n9521), .X(n6850) );
  inv_x1_sg U7681 ( .A(n9520), .X(n6848) );
  inv_x1_sg U7682 ( .A(n9519), .X(n6846) );
  inv_x1_sg U7683 ( .A(n9518), .X(n6844) );
  inv_x1_sg U7684 ( .A(n9517), .X(n6842) );
  inv_x1_sg U7685 ( .A(n9516), .X(n6840) );
  inv_x1_sg U7686 ( .A(n9515), .X(n6838) );
  inv_x1_sg U7687 ( .A(n9514), .X(n6836) );
  inv_x1_sg U7688 ( .A(n9513), .X(n6834) );
  inv_x1_sg U7689 ( .A(n9512), .X(n6832) );
  inv_x1_sg U7690 ( .A(n9511), .X(n6830) );
  inv_x1_sg U7691 ( .A(n9510), .X(n6828) );
  inv_x1_sg U7692 ( .A(n9509), .X(n6826) );
  inv_x1_sg U7693 ( .A(n9508), .X(n6824) );
  inv_x1_sg U7694 ( .A(n9507), .X(n6662) );
  inv_x1_sg U7695 ( .A(n9506), .X(n6660) );
  inv_x1_sg U7696 ( .A(n9505), .X(n6658) );
  inv_x1_sg U7697 ( .A(n9504), .X(n6656) );
  inv_x1_sg U7698 ( .A(n9503), .X(n6654) );
  inv_x1_sg U7699 ( .A(n9502), .X(n6652) );
  inv_x1_sg U7700 ( .A(n9501), .X(n6650) );
  inv_x1_sg U7701 ( .A(n9500), .X(n6648) );
  inv_x1_sg U7702 ( .A(n9499), .X(n6646) );
  inv_x1_sg U7703 ( .A(n9498), .X(n6644) );
  inv_x1_sg U7704 ( .A(n9497), .X(n6642) );
  inv_x1_sg U7705 ( .A(n9496), .X(n6640) );
  inv_x1_sg U7706 ( .A(n9495), .X(n6638) );
  inv_x1_sg U7707 ( .A(n9494), .X(n6636) );
  inv_x1_sg U7708 ( .A(n9493), .X(n6634) );
  inv_x1_sg U7709 ( .A(n9492), .X(n6632) );
  inv_x1_sg U7710 ( .A(n9491), .X(n6630) );
  inv_x1_sg U7711 ( .A(n9490), .X(n6628) );
  inv_x1_sg U7712 ( .A(n9489), .X(n6626) );
  inv_x1_sg U7713 ( .A(n9488), .X(n6624) );
  inv_x1_sg U7714 ( .A(n9487), .X(n6582) );
  inv_x1_sg U7715 ( .A(n9486), .X(n6580) );
  inv_x1_sg U7716 ( .A(n9485), .X(n6578) );
  inv_x1_sg U7717 ( .A(n9484), .X(n6576) );
  inv_x1_sg U7718 ( .A(n9483), .X(n6574) );
  inv_x1_sg U7719 ( .A(n9482), .X(n6572) );
  inv_x1_sg U7720 ( .A(n9481), .X(n6570) );
  inv_x1_sg U7721 ( .A(n9480), .X(n6568) );
  inv_x1_sg U7722 ( .A(n9479), .X(n6566) );
  inv_x1_sg U7723 ( .A(n9478), .X(n6564) );
  inv_x1_sg U7724 ( .A(n9477), .X(n6562) );
  inv_x1_sg U7725 ( .A(n9476), .X(n6560) );
  inv_x1_sg U7726 ( .A(n9475), .X(n6558) );
  inv_x1_sg U7727 ( .A(n9474), .X(n6556) );
  inv_x1_sg U7728 ( .A(n9473), .X(n6554) );
  inv_x1_sg U7729 ( .A(n9472), .X(n6552) );
  inv_x1_sg U7730 ( .A(n9471), .X(n6550) );
  inv_x1_sg U7731 ( .A(n9470), .X(n6548) );
  inv_x1_sg U7732 ( .A(n9469), .X(n6546) );
  inv_x1_sg U7733 ( .A(n9468), .X(n6544) );
  inv_x1_sg U7734 ( .A(n9467), .X(n6462) );
  inv_x1_sg U7735 ( .A(n9466), .X(n6460) );
  inv_x1_sg U7736 ( .A(n9465), .X(n6458) );
  inv_x1_sg U7737 ( .A(n9464), .X(n6456) );
  inv_x1_sg U7738 ( .A(n9463), .X(n6454) );
  inv_x1_sg U7739 ( .A(n9462), .X(n6452) );
  inv_x1_sg U7740 ( .A(n9461), .X(n6450) );
  inv_x1_sg U7741 ( .A(n9460), .X(n6448) );
  inv_x1_sg U7742 ( .A(n9459), .X(n6446) );
  inv_x1_sg U7743 ( .A(n9458), .X(n6444) );
  inv_x1_sg U7744 ( .A(n9457), .X(n6442) );
  inv_x1_sg U7745 ( .A(n9456), .X(n6440) );
  inv_x1_sg U7746 ( .A(n9455), .X(n6438) );
  inv_x1_sg U7747 ( .A(n9454), .X(n6436) );
  inv_x1_sg U7748 ( .A(n9453), .X(n6434) );
  inv_x1_sg U7749 ( .A(n9452), .X(n6432) );
  inv_x1_sg U7750 ( .A(n9451), .X(n6430) );
  inv_x1_sg U7751 ( .A(n9450), .X(n6428) );
  inv_x1_sg U7752 ( .A(n9449), .X(n6426) );
  inv_x1_sg U7753 ( .A(n9448), .X(n6424) );
  inv_x1_sg U7754 ( .A(n9447), .X(n6542) );
  inv_x1_sg U7755 ( .A(n9446), .X(n6540) );
  inv_x1_sg U7756 ( .A(n9445), .X(n6538) );
  inv_x1_sg U7757 ( .A(n9444), .X(n6536) );
  inv_x1_sg U7758 ( .A(n9443), .X(n6534) );
  inv_x1_sg U7759 ( .A(n9442), .X(n6532) );
  inv_x1_sg U7760 ( .A(n9441), .X(n6530) );
  inv_x1_sg U7761 ( .A(n9440), .X(n6528) );
  inv_x1_sg U7762 ( .A(n9439), .X(n6526) );
  inv_x1_sg U7763 ( .A(n9438), .X(n6524) );
  inv_x1_sg U7764 ( .A(n9437), .X(n6522) );
  inv_x1_sg U7765 ( .A(n9436), .X(n6520) );
  inv_x1_sg U7766 ( .A(n9435), .X(n6518) );
  inv_x1_sg U7767 ( .A(n9434), .X(n6516) );
  inv_x1_sg U7768 ( .A(n9433), .X(n6514) );
  inv_x1_sg U7769 ( .A(n9432), .X(n6512) );
  inv_x1_sg U7770 ( .A(n9431), .X(n6510) );
  inv_x1_sg U7771 ( .A(n9430), .X(n6508) );
  inv_x1_sg U7772 ( .A(n9429), .X(n6506) );
  inv_x1_sg U7773 ( .A(n9428), .X(n6504) );
  inv_x1_sg U7774 ( .A(n9427), .X(n6982) );
  inv_x1_sg U7775 ( .A(n9426), .X(n6980) );
  inv_x1_sg U7776 ( .A(n9425), .X(n6978) );
  inv_x1_sg U7777 ( .A(n9424), .X(n6976) );
  inv_x1_sg U7778 ( .A(n9423), .X(n6974) );
  inv_x1_sg U7779 ( .A(n9422), .X(n6972) );
  inv_x1_sg U7780 ( .A(n9421), .X(n6970) );
  inv_x1_sg U7781 ( .A(n9420), .X(n6968) );
  inv_x1_sg U7782 ( .A(n9419), .X(n6966) );
  inv_x1_sg U7783 ( .A(n9418), .X(n6964) );
  inv_x1_sg U7784 ( .A(n9417), .X(n6962) );
  inv_x1_sg U7785 ( .A(n9416), .X(n6960) );
  inv_x1_sg U7786 ( .A(n9415), .X(n6958) );
  inv_x1_sg U7787 ( .A(n9414), .X(n6956) );
  inv_x1_sg U7788 ( .A(n9413), .X(n6954) );
  inv_x1_sg U7789 ( .A(n9412), .X(n6952) );
  inv_x1_sg U7790 ( .A(n9411), .X(n6950) );
  inv_x1_sg U7791 ( .A(n9410), .X(n6948) );
  inv_x1_sg U7792 ( .A(n9409), .X(n6946) );
  inv_x1_sg U7793 ( .A(n9408), .X(n6944) );
  inv_x1_sg U7794 ( .A(n9407), .X(n6942) );
  inv_x1_sg U7795 ( .A(n9406), .X(n6940) );
  inv_x1_sg U7796 ( .A(n9405), .X(n6938) );
  inv_x1_sg U7797 ( .A(n9404), .X(n6936) );
  inv_x1_sg U7798 ( .A(n9403), .X(n6934) );
  inv_x1_sg U7799 ( .A(n9402), .X(n6932) );
  inv_x1_sg U7800 ( .A(n9401), .X(n6930) );
  inv_x1_sg U7801 ( .A(n9400), .X(n6928) );
  inv_x1_sg U7802 ( .A(n9399), .X(n6926) );
  inv_x1_sg U7803 ( .A(n9398), .X(n6924) );
  inv_x1_sg U7804 ( .A(n9397), .X(n6922) );
  inv_x1_sg U7805 ( .A(n9396), .X(n6920) );
  inv_x1_sg U7806 ( .A(n9395), .X(n6918) );
  inv_x1_sg U7807 ( .A(n9394), .X(n6916) );
  inv_x1_sg U7808 ( .A(n9393), .X(n6914) );
  inv_x1_sg U7809 ( .A(n9392), .X(n6912) );
  inv_x1_sg U7810 ( .A(n9391), .X(n6910) );
  inv_x1_sg U7811 ( .A(n9390), .X(n6908) );
  inv_x1_sg U7812 ( .A(n9389), .X(n6906) );
  inv_x1_sg U7813 ( .A(n9388), .X(n6904) );
  inv_x1_sg U7814 ( .A(n9387), .X(n6742) );
  inv_x1_sg U7815 ( .A(n9386), .X(n6740) );
  inv_x1_sg U7816 ( .A(n9385), .X(n6738) );
  inv_x1_sg U7817 ( .A(n9384), .X(n6736) );
  inv_x1_sg U7818 ( .A(n9383), .X(n6734) );
  inv_x1_sg U7819 ( .A(n9382), .X(n6732) );
  inv_x1_sg U7820 ( .A(n9381), .X(n6730) );
  inv_x1_sg U7821 ( .A(n9380), .X(n6728) );
  inv_x1_sg U7822 ( .A(n9379), .X(n6726) );
  inv_x1_sg U7823 ( .A(n9378), .X(n6724) );
  inv_x1_sg U7824 ( .A(n9377), .X(n6722) );
  inv_x1_sg U7825 ( .A(n9376), .X(n6720) );
  inv_x1_sg U7826 ( .A(n9375), .X(n6718) );
  inv_x1_sg U7827 ( .A(n9374), .X(n6716) );
  inv_x1_sg U7828 ( .A(n9373), .X(n6714) );
  inv_x1_sg U7829 ( .A(n9372), .X(n6712) );
  inv_x1_sg U7830 ( .A(n9371), .X(n6710) );
  inv_x1_sg U7831 ( .A(n9370), .X(n6708) );
  inv_x1_sg U7832 ( .A(n9369), .X(n6706) );
  inv_x1_sg U7833 ( .A(n9368), .X(n6704) );
  inv_x1_sg U7834 ( .A(n9367), .X(n6822) );
  inv_x1_sg U7835 ( .A(n9366), .X(n6820) );
  inv_x1_sg U7836 ( .A(n9365), .X(n6818) );
  inv_x1_sg U7837 ( .A(n9364), .X(n6816) );
  inv_x1_sg U7838 ( .A(n9363), .X(n6814) );
  inv_x1_sg U7839 ( .A(n9362), .X(n6812) );
  inv_x1_sg U7840 ( .A(n9361), .X(n6810) );
  inv_x1_sg U7841 ( .A(n9360), .X(n6808) );
  inv_x1_sg U7842 ( .A(n9359), .X(n6806) );
  inv_x1_sg U7843 ( .A(n9358), .X(n6804) );
  inv_x1_sg U7844 ( .A(n9357), .X(n6802) );
  inv_x1_sg U7845 ( .A(n9356), .X(n6800) );
  inv_x1_sg U7846 ( .A(n9355), .X(n6798) );
  inv_x1_sg U7847 ( .A(n9354), .X(n6796) );
  inv_x1_sg U7848 ( .A(n9353), .X(n6794) );
  inv_x1_sg U7849 ( .A(n9352), .X(n6792) );
  inv_x1_sg U7850 ( .A(n9351), .X(n6790) );
  inv_x1_sg U7851 ( .A(n9350), .X(n6788) );
  inv_x1_sg U7852 ( .A(n9349), .X(n6786) );
  inv_x1_sg U7853 ( .A(n9348), .X(n6784) );
  inv_x1_sg U7854 ( .A(n9347), .X(n6702) );
  inv_x1_sg U7855 ( .A(n9346), .X(n6700) );
  inv_x1_sg U7856 ( .A(n9345), .X(n6698) );
  inv_x1_sg U7857 ( .A(n9344), .X(n6696) );
  inv_x1_sg U7858 ( .A(n9343), .X(n6694) );
  inv_x1_sg U7859 ( .A(n9342), .X(n6692) );
  inv_x1_sg U7860 ( .A(n9341), .X(n6690) );
  inv_x1_sg U7861 ( .A(n9340), .X(n6688) );
  inv_x1_sg U7862 ( .A(n9339), .X(n6686) );
  inv_x1_sg U7863 ( .A(n9338), .X(n6684) );
  inv_x1_sg U7864 ( .A(n9337), .X(n6682) );
  inv_x1_sg U7865 ( .A(n9336), .X(n6680) );
  inv_x1_sg U7866 ( .A(n9335), .X(n6678) );
  inv_x1_sg U7867 ( .A(n9334), .X(n6676) );
  inv_x1_sg U7868 ( .A(n9333), .X(n6674) );
  inv_x1_sg U7869 ( .A(n9332), .X(n6672) );
  inv_x1_sg U7870 ( .A(n9331), .X(n6670) );
  inv_x1_sg U7871 ( .A(n9330), .X(n6668) );
  inv_x1_sg U7872 ( .A(n9329), .X(n6666) );
  inv_x1_sg U7873 ( .A(n9328), .X(n6664) );
  inv_x1_sg U7874 ( .A(n9327), .X(n6622) );
  inv_x1_sg U7875 ( .A(n9326), .X(n6620) );
  inv_x1_sg U7876 ( .A(n9325), .X(n6618) );
  inv_x1_sg U7877 ( .A(n9324), .X(n6616) );
  inv_x1_sg U7878 ( .A(n9323), .X(n6614) );
  inv_x1_sg U7879 ( .A(n9322), .X(n6612) );
  inv_x1_sg U7880 ( .A(n9321), .X(n6610) );
  inv_x1_sg U7881 ( .A(n9320), .X(n6608) );
  inv_x1_sg U7882 ( .A(n9319), .X(n6606) );
  inv_x1_sg U7883 ( .A(n9318), .X(n6604) );
  inv_x1_sg U7884 ( .A(n9317), .X(n6602) );
  inv_x1_sg U7885 ( .A(n9316), .X(n6600) );
  inv_x1_sg U7886 ( .A(n9315), .X(n6598) );
  inv_x1_sg U7887 ( .A(n9314), .X(n6596) );
  inv_x1_sg U7888 ( .A(n9313), .X(n6594) );
  inv_x1_sg U7889 ( .A(n9312), .X(n6592) );
  inv_x1_sg U7890 ( .A(n9311), .X(n6590) );
  inv_x1_sg U7891 ( .A(n9310), .X(n6588) );
  inv_x1_sg U7892 ( .A(n9309), .X(n6586) );
  inv_x1_sg U7893 ( .A(n9308), .X(n6584) );
  inv_x1_sg U7894 ( .A(n9307), .X(n6422) );
  inv_x1_sg U7895 ( .A(n9306), .X(n6420) );
  inv_x1_sg U7896 ( .A(n9305), .X(n6418) );
  inv_x1_sg U7897 ( .A(n9304), .X(n6416) );
  inv_x1_sg U7898 ( .A(n9303), .X(n6414) );
  inv_x1_sg U7899 ( .A(n9302), .X(n6412) );
  inv_x1_sg U7900 ( .A(n9301), .X(n6410) );
  inv_x1_sg U7901 ( .A(n9300), .X(n6408) );
  inv_x1_sg U7902 ( .A(n9299), .X(n6406) );
  inv_x1_sg U7903 ( .A(n9298), .X(n6404) );
  inv_x1_sg U7904 ( .A(n9297), .X(n6402) );
  inv_x1_sg U7905 ( .A(n9296), .X(n6400) );
  inv_x1_sg U7906 ( .A(n9295), .X(n6398) );
  inv_x1_sg U7907 ( .A(n9294), .X(n6396) );
  inv_x1_sg U7908 ( .A(n9293), .X(n6394) );
  inv_x1_sg U7909 ( .A(n9292), .X(n6392) );
  inv_x1_sg U7910 ( .A(n9291), .X(n6390) );
  inv_x1_sg U7911 ( .A(n9290), .X(n6388) );
  inv_x1_sg U7912 ( .A(n9289), .X(n6386) );
  inv_x1_sg U7913 ( .A(n9288), .X(n6384) );
  inv_x1_sg U7914 ( .A(n9287), .X(n6502) );
  inv_x1_sg U7915 ( .A(n9286), .X(n6500) );
  inv_x1_sg U7916 ( .A(n9285), .X(n6498) );
  inv_x1_sg U7917 ( .A(n9284), .X(n6496) );
  inv_x1_sg U7918 ( .A(n9283), .X(n6494) );
  inv_x1_sg U7919 ( .A(n9282), .X(n6492) );
  inv_x1_sg U7920 ( .A(n9281), .X(n6490) );
  inv_x1_sg U7921 ( .A(n9280), .X(n6488) );
  inv_x1_sg U7922 ( .A(n9279), .X(n6486) );
  inv_x1_sg U7923 ( .A(n9278), .X(n6484) );
  inv_x1_sg U7924 ( .A(n9277), .X(n6482) );
  inv_x1_sg U7925 ( .A(n9276), .X(n6480) );
  inv_x1_sg U7926 ( .A(n9275), .X(n6478) );
  inv_x1_sg U7927 ( .A(n9274), .X(n6476) );
  inv_x1_sg U7928 ( .A(n9273), .X(n6474) );
  inv_x1_sg U7929 ( .A(n9272), .X(n6472) );
  inv_x1_sg U7930 ( .A(n9271), .X(n6470) );
  inv_x1_sg U7931 ( .A(n9270), .X(n6468) );
  inv_x1_sg U7932 ( .A(n9269), .X(n6466) );
  inv_x1_sg U7933 ( .A(n9268), .X(n6464) );
  inv_x1_sg U7934 ( .A(n9267), .X(n7022) );
  inv_x1_sg U7935 ( .A(n9266), .X(n7020) );
  inv_x1_sg U7936 ( .A(n9265), .X(n7018) );
  inv_x1_sg U7937 ( .A(n9264), .X(n7016) );
  inv_x1_sg U7938 ( .A(n9263), .X(n7014) );
  inv_x1_sg U7939 ( .A(n9262), .X(n7012) );
  inv_x1_sg U7940 ( .A(n9261), .X(n7010) );
  inv_x1_sg U7941 ( .A(n9260), .X(n7008) );
  inv_x1_sg U7942 ( .A(n9259), .X(n7006) );
  inv_x1_sg U7943 ( .A(n9258), .X(n7004) );
  inv_x1_sg U7944 ( .A(n9257), .X(n7002) );
  inv_x1_sg U7945 ( .A(n9256), .X(n7000) );
  inv_x1_sg U7946 ( .A(n9255), .X(n6998) );
  inv_x1_sg U7947 ( .A(n9254), .X(n6996) );
  inv_x1_sg U7948 ( .A(n9253), .X(n6994) );
  inv_x1_sg U7949 ( .A(n9252), .X(n6992) );
  inv_x1_sg U7950 ( .A(n9251), .X(n6990) );
  inv_x1_sg U7951 ( .A(n9250), .X(n6988) );
  inv_x1_sg U7952 ( .A(n9249), .X(n6986) );
  inv_x1_sg U7953 ( .A(n9248), .X(n6984) );
  inv_x1_sg U7954 ( .A(n823), .X(n9182) );
  nand_x1_sg U7955 ( .A(n7523), .B(n1561), .X(n749) );
  nand_x1_sg U7956 ( .A(n7523), .B(n1563), .X(n747) );
  nand_x1_sg U7957 ( .A(n7523), .B(n1554), .X(n755) );
  nand_x1_sg U7958 ( .A(n7523), .B(n1555), .X(n754) );
  nand_x1_sg U7959 ( .A(n7523), .B(n1550), .X(n758) );
  nand_x1_sg U7960 ( .A(n7523), .B(n1551), .X(n757) );
  nand_x1_sg U7961 ( .A(n7523), .B(n1562), .X(n748) );
  nand_x1_sg U7962 ( .A(n7523), .B(n1560), .X(n750) );
  nand_x1_sg U7963 ( .A(n7523), .B(n1569), .X(n745) );
  nand_x1_sg U7964 ( .A(n7523), .B(n1571), .X(n743) );
  nand_x1_sg U7965 ( .A(n7523), .B(n1570), .X(n744) );
  nand_x1_sg U7966 ( .A(n7523), .B(n1574), .X(n740) );
  nand_x1_sg U7967 ( .A(n7523), .B(n1572), .X(n742) );
  nand_x1_sg U7968 ( .A(n7523), .B(n1573), .X(n741) );
  nand_x1_sg U7969 ( .A(n7523), .B(n1557), .X(n752) );
  nand_x1_sg U7970 ( .A(n7523), .B(n1559), .X(n751) );
  nand_x1_sg U7971 ( .A(n7523), .B(n1556), .X(n753) );
  nand_x1_sg U7972 ( .A(n7523), .B(n1566), .X(n746) );
  nand_x1_sg U7973 ( .A(n7523), .B(n1547), .X(n761) );
  nand_x1_sg U7974 ( .A(n7523), .B(n1548), .X(n760) );
  nand_x1_sg U7975 ( .A(n7523), .B(n1544), .X(n764) );
  nand_x1_sg U7976 ( .A(n7523), .B(n1545), .X(n763) );
  nand_x1_sg U7977 ( .A(n7523), .B(n1541), .X(n767) );
  nand_x1_sg U7978 ( .A(n7523), .B(n1542), .X(n766) );
  nand_x1_sg U7979 ( .A(n7523), .B(n1538), .X(n770) );
  nand_x1_sg U7980 ( .A(n7523), .B(n1539), .X(n769) );
  nand_x1_sg U7981 ( .A(n7523), .B(n1536), .X(n771) );
  nand_x1_sg U7982 ( .A(n7523), .B(n1540), .X(n768) );
  nand_x1_sg U7983 ( .A(n7523), .B(n1543), .X(n765) );
  nand_x1_sg U7984 ( .A(n7523), .B(n1546), .X(n762) );
  nand_x1_sg U7985 ( .A(n7523), .B(n1549), .X(n759) );
  nand_x1_sg U7986 ( .A(n7523), .B(n1552), .X(n756) );
  nand_x1_sg U7987 ( .A(n4394), .B(n4395), .X(n5793) );
  nand_x1_sg U7988 ( .A(n4182), .B(n7560), .X(n4394) );
  nand_x1_sg U7989 ( .A(n4193), .B(n4194), .X(n5707) );
  nand_x1_sg U7990 ( .A(n4182), .B(n4195), .X(n4194) );
  nand_x1_sg U7991 ( .A(n4188), .B(n4189), .X(n5706) );
  nand_x1_sg U7992 ( .A(n7568), .B(n4187), .X(n4188) );
  nand_x1_sg U7993 ( .A(n4190), .B(n7393), .X(n4189) );
  nand_x1_sg U7994 ( .A(n4204), .B(n4205), .X(n5709) );
  nand_x1_sg U7995 ( .A(n4198), .B(n4199), .X(n5708) );
  nand_x1_sg U7996 ( .A(n4180), .B(n4181), .X(n5705) );
  nand_x1_sg U7997 ( .A(n4182), .B(n4183), .X(n4181) );
  nand_x1_sg U7998 ( .A(n4184), .B(n4185), .X(n4183) );
  nand_x1_sg U7999 ( .A(n4304), .B(n9189), .X(n5752) );
  inv_x1_sg U8000 ( .A(n4305), .X(n9189) );
  nand_x1_sg U8001 ( .A(n3090), .B(n3091), .X(\update_output_0/n3549 ) );
  nand_x1_sg U8002 ( .A(n4291), .B(n4292), .X(n5750) );
  nand_x1_sg U8003 ( .A(n7570), .B(n4294), .X(n4291) );
  nand_x1_sg U8004 ( .A(n4295), .B(n9194), .X(n5751) );
  inv_x1_sg U8005 ( .A(n4296), .X(n9194) );
  nand_x1_sg U8006 ( .A(n4265), .B(n4266), .X(n5737) );
  nand_x1_sg U8007 ( .A(n7415), .B(n7443), .X(n4266) );
  nand_x1_sg U8008 ( .A(n4273), .B(n4274), .X(n5741) );
  nand_x1_sg U8009 ( .A(n7415), .B(n7488), .X(n4274) );
  nand_x1_sg U8010 ( .A(n4289), .B(n4290), .X(n5749) );
  nand_x1_sg U8011 ( .A(n7415), .B(n7490), .X(n4290) );
  nand_x1_sg U8012 ( .A(n4277), .B(n4278), .X(n5743) );
  nand_x1_sg U8013 ( .A(n7415), .B(n7494), .X(n4278) );
  nand_x1_sg U8014 ( .A(n4250), .B(n4251), .X(n5730) );
  nand_x1_sg U8015 ( .A(n7415), .B(n7492), .X(n4251) );
  nand_x1_sg U8016 ( .A(n4267), .B(n4268), .X(n5738) );
  nand_x1_sg U8017 ( .A(n7415), .B(n7482), .X(n4268) );
  nand_x1_sg U8018 ( .A(n4257), .B(n4258), .X(n5733) );
  nand_x1_sg U8019 ( .A(n7415), .B(n7480), .X(n4258) );
  nand_x1_sg U8020 ( .A(n4283), .B(n4284), .X(n5746) );
  nand_x1_sg U8021 ( .A(n7415), .B(n7484), .X(n4284) );
  nand_x1_sg U8022 ( .A(n4279), .B(n4280), .X(n5744) );
  nand_x1_sg U8023 ( .A(n7415), .B(n7486), .X(n4280) );
  nand_x1_sg U8024 ( .A(n4287), .B(n4288), .X(n5748) );
  nand_x1_sg U8025 ( .A(n7415), .B(n7470), .X(n4288) );
  nand_x1_sg U8026 ( .A(n4263), .B(n4264), .X(n5736) );
  nand_x1_sg U8027 ( .A(n7415), .B(n7468), .X(n4264) );
  nand_x1_sg U8028 ( .A(n4261), .B(n4262), .X(n5735) );
  nand_x1_sg U8029 ( .A(n7415), .B(n7450), .X(n4262) );
  nand_x1_sg U8030 ( .A(n4253), .B(n4254), .X(n5731) );
  nand_x1_sg U8031 ( .A(n7415), .B(n7445), .X(n4254) );
  nand_x1_sg U8032 ( .A(n4271), .B(n4272), .X(n5740) );
  nand_x1_sg U8033 ( .A(n7415), .B(n7452), .X(n4272) );
  nand_x1_sg U8034 ( .A(n4259), .B(n4260), .X(n5734) );
  nand_x1_sg U8035 ( .A(n7415), .B(n7454), .X(n4260) );
  nand_x1_sg U8036 ( .A(n4255), .B(n4256), .X(n5732) );
  nand_x1_sg U8037 ( .A(n7415), .B(n7474), .X(n4256) );
  nand_x1_sg U8038 ( .A(n4275), .B(n4276), .X(n5742) );
  nand_x1_sg U8039 ( .A(n7415), .B(n7472), .X(n4276) );
  nand_x1_sg U8040 ( .A(n4281), .B(n4282), .X(n5745) );
  nand_x1_sg U8041 ( .A(n7415), .B(n7478), .X(n4282) );
  nand_x1_sg U8042 ( .A(n4269), .B(n4270), .X(n5739) );
  nand_x1_sg U8043 ( .A(n7415), .B(n7476), .X(n4270) );
  nand_x1_sg U8044 ( .A(n4285), .B(n4286), .X(n5747) );
  nand_x1_sg U8045 ( .A(n7415), .B(n7466), .X(n4286) );
  nand_x1_sg U8046 ( .A(n4213), .B(n4214), .X(n5712) );
  nand_x1_sg U8047 ( .A(n7416), .B(n7443), .X(n4214) );
  nand_x1_sg U8048 ( .A(n4229), .B(n4230), .X(n5720) );
  nand_x1_sg U8049 ( .A(n7416), .B(n7488), .X(n4230) );
  nand_x1_sg U8050 ( .A(n4225), .B(n4226), .X(n5718) );
  nand_x1_sg U8051 ( .A(n7416), .B(n7490), .X(n4226) );
  nand_x1_sg U8052 ( .A(n4233), .B(n4234), .X(n5722) );
  nand_x1_sg U8053 ( .A(n7416), .B(n7494), .X(n4234) );
  nand_x1_sg U8054 ( .A(n4245), .B(n4246), .X(n5728) );
  nand_x1_sg U8055 ( .A(n7416), .B(n7492), .X(n4246) );
  nand_x1_sg U8056 ( .A(n4241), .B(n4242), .X(n5726) );
  nand_x1_sg U8057 ( .A(n7416), .B(n7482), .X(n4242) );
  nand_x1_sg U8058 ( .A(n4227), .B(n4228), .X(n5719) );
  nand_x1_sg U8059 ( .A(n7416), .B(n7480), .X(n4228) );
  nand_x1_sg U8060 ( .A(n4219), .B(n4220), .X(n5715) );
  nand_x1_sg U8061 ( .A(n7416), .B(n7484), .X(n4220) );
  nand_x1_sg U8062 ( .A(n4208), .B(n4209), .X(n5710) );
  nand_x1_sg U8063 ( .A(n7416), .B(n7486), .X(n4209) );
  nand_x1_sg U8064 ( .A(n4247), .B(n4248), .X(n5729) );
  nand_x1_sg U8065 ( .A(n7416), .B(n7470), .X(n4248) );
  nand_x1_sg U8066 ( .A(n4217), .B(n4218), .X(n5714) );
  nand_x1_sg U8067 ( .A(n7416), .B(n7468), .X(n4218) );
  nand_x1_sg U8068 ( .A(n4215), .B(n4216), .X(n5713) );
  nand_x1_sg U8069 ( .A(n7416), .B(n7450), .X(n4216) );
  nand_x1_sg U8070 ( .A(n4235), .B(n4236), .X(n5723) );
  nand_x1_sg U8071 ( .A(n7416), .B(n7445), .X(n4236) );
  nand_x1_sg U8072 ( .A(n4211), .B(n4212), .X(n5711) );
  nand_x1_sg U8073 ( .A(n7416), .B(n7452), .X(n4212) );
  nand_x1_sg U8074 ( .A(n4239), .B(n4240), .X(n5725) );
  nand_x1_sg U8075 ( .A(n7416), .B(n7454), .X(n4240) );
  nand_x1_sg U8076 ( .A(n4221), .B(n4222), .X(n5716) );
  nand_x1_sg U8077 ( .A(n7416), .B(n7474), .X(n4222) );
  nand_x1_sg U8078 ( .A(n4231), .B(n4232), .X(n5721) );
  nand_x1_sg U8079 ( .A(n7416), .B(n7472), .X(n4232) );
  nand_x1_sg U8080 ( .A(n4223), .B(n4224), .X(n5717) );
  nand_x1_sg U8081 ( .A(n7416), .B(n7478), .X(n4224) );
  nand_x1_sg U8082 ( .A(n4237), .B(n4238), .X(n5724) );
  nand_x1_sg U8083 ( .A(n7416), .B(n7476), .X(n4238) );
  nand_x1_sg U8084 ( .A(n4243), .B(n4244), .X(n5727) );
  nand_x1_sg U8085 ( .A(n7416), .B(n7466), .X(n4244) );
  nand_x1_sg U8086 ( .A(n4387), .B(n4388), .X(n5791) );
  nand_x1_sg U8087 ( .A(n7443), .B(n7497), .X(n4388) );
  nand_x1_sg U8088 ( .A(n4385), .B(n4386), .X(n5790) );
  nand_x1_sg U8089 ( .A(n7488), .B(n7496), .X(n4386) );
  nand_x1_sg U8090 ( .A(n4363), .B(n4364), .X(n5779) );
  nand_x1_sg U8091 ( .A(n7490), .B(n7497), .X(n4364) );
  nand_x1_sg U8092 ( .A(n4359), .B(n4360), .X(n5777) );
  nand_x1_sg U8093 ( .A(n7494), .B(n7496), .X(n4360) );
  nand_x1_sg U8094 ( .A(n4371), .B(n4372), .X(n5783) );
  nand_x1_sg U8095 ( .A(n7492), .B(n7496), .X(n4372) );
  nand_x1_sg U8096 ( .A(n4373), .B(n4374), .X(n5784) );
  nand_x1_sg U8097 ( .A(n7482), .B(n7497), .X(n4374) );
  nand_x1_sg U8098 ( .A(n4357), .B(n4358), .X(n5776) );
  nand_x1_sg U8099 ( .A(n7480), .B(n7497), .X(n4358) );
  nand_x1_sg U8100 ( .A(n4383), .B(n4384), .X(n5789) );
  nand_x1_sg U8101 ( .A(n3873), .B(n7496), .X(n4384) );
  nand_x1_sg U8102 ( .A(n4353), .B(n4354), .X(n5774) );
  nand_x1_sg U8103 ( .A(n3861), .B(n7496), .X(n4354) );
  nand_x1_sg U8104 ( .A(n4381), .B(n4382), .X(n5788) );
  nand_x1_sg U8105 ( .A(n7470), .B(n7497), .X(n4382) );
  nand_x1_sg U8106 ( .A(n4361), .B(n4362), .X(n5778) );
  nand_x1_sg U8107 ( .A(n3834), .B(n7497), .X(n4362) );
  nand_x1_sg U8108 ( .A(n4355), .B(n4356), .X(n5775) );
  nand_x1_sg U8109 ( .A(n7450), .B(n4352), .X(n4356) );
  nand_x1_sg U8110 ( .A(n4365), .B(n4366), .X(n5780) );
  nand_x1_sg U8111 ( .A(n7445), .B(n7496), .X(n4366) );
  nand_x1_sg U8112 ( .A(n4375), .B(n4376), .X(n5785) );
  nand_x1_sg U8113 ( .A(n7452), .B(n7497), .X(n4376) );
  nand_x1_sg U8114 ( .A(n4367), .B(n4368), .X(n5781) );
  nand_x1_sg U8115 ( .A(n7454), .B(n7496), .X(n4368) );
  nand_x1_sg U8116 ( .A(n4377), .B(n4378), .X(n5786) );
  nand_x1_sg U8117 ( .A(n7474), .B(n7496), .X(n4378) );
  nand_x1_sg U8118 ( .A(n4350), .B(n4351), .X(n5773) );
  nand_x1_sg U8119 ( .A(n7472), .B(n7497), .X(n4351) );
  nand_x1_sg U8120 ( .A(n4369), .B(n4370), .X(n5782) );
  nand_x1_sg U8121 ( .A(n7478), .B(n7497), .X(n4370) );
  nand_x1_sg U8122 ( .A(n4389), .B(n4390), .X(n5792) );
  nand_x1_sg U8123 ( .A(n3827), .B(n7496), .X(n4390) );
  nand_x1_sg U8124 ( .A(n4379), .B(n4380), .X(n5787) );
  nand_x1_sg U8125 ( .A(n3879), .B(n7496), .X(n4380) );
  nand_x1_sg U8126 ( .A(n5047), .B(n5048), .X(n5857) );
  nand_x1_sg U8127 ( .A(n7443), .B(n7464), .X(n5048) );
  nand_x1_sg U8128 ( .A(n4541), .B(n4542), .X(n5808) );
  nand_x1_sg U8129 ( .A(n7488), .B(n7463), .X(n4542) );
  nand_x1_sg U8130 ( .A(n4495), .B(n4496), .X(n5802) );
  nand_x1_sg U8131 ( .A(n7490), .B(n7464), .X(n4496) );
  nand_x1_sg U8132 ( .A(n4399), .B(n4400), .X(n5795) );
  nand_x1_sg U8133 ( .A(n7494), .B(n7463), .X(n4400) );
  nand_x1_sg U8134 ( .A(n4457), .B(n4458), .X(n5800) );
  nand_x1_sg U8135 ( .A(n7492), .B(n7463), .X(n4458) );
  nand_x1_sg U8136 ( .A(n4663), .B(n4664), .X(n5818) );
  nand_x1_sg U8137 ( .A(n7482), .B(n7463), .X(n4664) );
  nand_x1_sg U8138 ( .A(n4707), .B(n4708), .X(n5823) );
  nand_x1_sg U8139 ( .A(n7480), .B(n7463), .X(n4708) );
  nand_x1_sg U8140 ( .A(n4625), .B(n4626), .X(n5816) );
  nand_x1_sg U8141 ( .A(n7484), .B(n7464), .X(n4626) );
  nand_x1_sg U8142 ( .A(n4579), .B(n4580), .X(n5810) );
  nand_x1_sg U8143 ( .A(n7486), .B(n7463), .X(n4580) );
  nand_x1_sg U8144 ( .A(n4917), .B(n4918), .X(n5843) );
  nand_x1_sg U8145 ( .A(n7470), .B(n7463), .X(n4918) );
  nand_x1_sg U8146 ( .A(n4963), .B(n4964), .X(n5849) );
  nand_x1_sg U8147 ( .A(n7468), .B(n7463), .X(n4964) );
  nand_x1_sg U8148 ( .A(n5051), .B(n5052), .X(n5859) );
  nand_x1_sg U8149 ( .A(n7450), .B(n7463), .X(n5052) );
  nand_x1_sg U8150 ( .A(n5045), .B(n5046), .X(n5856) );
  nand_x1_sg U8151 ( .A(n7445), .B(n7463), .X(n5046) );
  nand_x1_sg U8152 ( .A(n5049), .B(n5050), .X(n5858) );
  nand_x1_sg U8153 ( .A(n7452), .B(n7463), .X(n5050) );
  nand_x1_sg U8154 ( .A(n5043), .B(n5044), .X(n5855) );
  nand_x1_sg U8155 ( .A(n7454), .B(n7463), .X(n5044) );
  nand_x1_sg U8156 ( .A(n4833), .B(n4834), .X(n5835) );
  nand_x1_sg U8157 ( .A(n7474), .B(n7463), .X(n4834) );
  nand_x1_sg U8158 ( .A(n4879), .B(n4880), .X(n5841) );
  nand_x1_sg U8159 ( .A(n7472), .B(n7464), .X(n4880) );
  nand_x1_sg U8160 ( .A(n4749), .B(n4750), .X(n5827) );
  nand_x1_sg U8161 ( .A(n7478), .B(n7464), .X(n4750) );
  nand_x1_sg U8162 ( .A(n4791), .B(n4792), .X(n5831) );
  nand_x1_sg U8163 ( .A(n7476), .B(n7463), .X(n4792) );
  nand_x1_sg U8164 ( .A(n5005), .B(n5006), .X(n5853) );
  nand_x1_sg U8165 ( .A(n7466), .B(n7464), .X(n5006) );
  nand_x1_sg U8166 ( .A(n5056), .B(n5057), .X(n5861) );
  nand_x1_sg U8167 ( .A(n7412), .B(n7443), .X(n5057) );
  nand_x1_sg U8168 ( .A(n4543), .B(n4544), .X(n5809) );
  nand_x1_sg U8169 ( .A(n7412), .B(n7488), .X(n4544) );
  nand_x1_sg U8170 ( .A(n4499), .B(n4500), .X(n5804) );
  nand_x1_sg U8171 ( .A(n7412), .B(n7490), .X(n4500) );
  nand_x1_sg U8172 ( .A(n4402), .B(n4403), .X(n5796) );
  nand_x1_sg U8173 ( .A(n7412), .B(n7494), .X(n4403) );
  nand_x1_sg U8174 ( .A(n4459), .B(n4460), .X(n5801) );
  nand_x1_sg U8175 ( .A(n7412), .B(n7492), .X(n4460) );
  nand_x1_sg U8176 ( .A(n4667), .B(n4668), .X(n5820) );
  nand_x1_sg U8177 ( .A(n7412), .B(n7482), .X(n4668) );
  nand_x1_sg U8178 ( .A(n4709), .B(n4710), .X(n5824) );
  nand_x1_sg U8179 ( .A(n7412), .B(n7480), .X(n4710) );
  nand_x1_sg U8180 ( .A(n4627), .B(n4628), .X(n5817) );
  nand_x1_sg U8181 ( .A(n7412), .B(n7484), .X(n4628) );
  nand_x1_sg U8182 ( .A(n4581), .B(n4582), .X(n5811) );
  nand_x1_sg U8183 ( .A(n7412), .B(n7486), .X(n4582) );
  nand_x1_sg U8184 ( .A(n4919), .B(n4920), .X(n5844) );
  nand_x1_sg U8185 ( .A(n7412), .B(n7470), .X(n4920) );
  nand_x1_sg U8186 ( .A(n4965), .B(n4966), .X(n5850) );
  nand_x1_sg U8187 ( .A(n7412), .B(n7468), .X(n4966) );
  nand_x1_sg U8188 ( .A(n5054), .B(n5055), .X(n5860) );
  nand_x1_sg U8189 ( .A(n7412), .B(n7450), .X(n5055) );
  nand_x1_sg U8190 ( .A(n5060), .B(n5061), .X(n5863) );
  nand_x1_sg U8191 ( .A(n7412), .B(n7445), .X(n5061) );
  nand_x1_sg U8192 ( .A(n5058), .B(n5059), .X(n5862) );
  nand_x1_sg U8193 ( .A(n7412), .B(n7452), .X(n5059) );
  nand_x1_sg U8194 ( .A(n5062), .B(n5063), .X(n5864) );
  nand_x1_sg U8195 ( .A(n7412), .B(n7454), .X(n5063) );
  nand_x1_sg U8196 ( .A(n4835), .B(n4836), .X(n5836) );
  nand_x1_sg U8197 ( .A(n7412), .B(n7474), .X(n4836) );
  nand_x1_sg U8198 ( .A(n4881), .B(n4882), .X(n5842) );
  nand_x1_sg U8199 ( .A(n7412), .B(n7472), .X(n4882) );
  nand_x1_sg U8200 ( .A(n4751), .B(n4752), .X(n5828) );
  nand_x1_sg U8201 ( .A(n7412), .B(n7478), .X(n4752) );
  nand_x1_sg U8202 ( .A(n4793), .B(n4794), .X(n5832) );
  nand_x1_sg U8203 ( .A(n7412), .B(n7476), .X(n4794) );
  nand_x1_sg U8204 ( .A(n5007), .B(n5008), .X(n5854) );
  nand_x1_sg U8205 ( .A(n7412), .B(n7466), .X(n5008) );
  nand_x1_sg U8206 ( .A(n5067), .B(n5068), .X(n5866) );
  nand_x1_sg U8207 ( .A(n7411), .B(n7443), .X(n5068) );
  nand_x1_sg U8208 ( .A(n4537), .B(n4538), .X(n5806) );
  nand_x1_sg U8209 ( .A(n7411), .B(n7488), .X(n4538) );
  nand_x1_sg U8210 ( .A(n4501), .B(n4502), .X(n5805) );
  nand_x1_sg U8211 ( .A(n7411), .B(n7490), .X(n4502) );
  nand_x1_sg U8212 ( .A(n4396), .B(n4397), .X(n5794) );
  nand_x1_sg U8213 ( .A(n7411), .B(n7494), .X(n4397) );
  nand_x1_sg U8214 ( .A(n4453), .B(n4454), .X(n5798) );
  nand_x1_sg U8215 ( .A(n7411), .B(n7492), .X(n4454) );
  nand_x1_sg U8216 ( .A(n4671), .B(n4672), .X(n5822) );
  nand_x1_sg U8217 ( .A(n7411), .B(n7482), .X(n4672) );
  nand_x1_sg U8218 ( .A(n4713), .B(n4714), .X(n5826) );
  nand_x1_sg U8219 ( .A(n7411), .B(n7480), .X(n4714) );
  nand_x1_sg U8220 ( .A(n4621), .B(n4622), .X(n5814) );
  nand_x1_sg U8221 ( .A(n7411), .B(n7484), .X(n4622) );
  nand_x1_sg U8222 ( .A(n4585), .B(n4586), .X(n5813) );
  nand_x1_sg U8223 ( .A(n7411), .B(n7486), .X(n4586) );
  nand_x1_sg U8224 ( .A(n4923), .B(n4924), .X(n5846) );
  nand_x1_sg U8225 ( .A(n7411), .B(n7470), .X(n4924) );
  nand_x1_sg U8226 ( .A(n4959), .B(n4960), .X(n5847) );
  nand_x1_sg U8227 ( .A(n7411), .B(n7468), .X(n4960) );
  nand_x1_sg U8228 ( .A(n5073), .B(n5074), .X(n5869) );
  nand_x1_sg U8229 ( .A(n7411), .B(n7450), .X(n5074) );
  nand_x1_sg U8230 ( .A(n5065), .B(n5066), .X(n5865) );
  nand_x1_sg U8231 ( .A(n7411), .B(n7445), .X(n5066) );
  nand_x1_sg U8232 ( .A(n5069), .B(n5070), .X(n5867) );
  nand_x1_sg U8233 ( .A(n7411), .B(n7452), .X(n5070) );
  nand_x1_sg U8234 ( .A(n5071), .B(n5072), .X(n5868) );
  nand_x1_sg U8235 ( .A(n7411), .B(n7454), .X(n5072) );
  nand_x1_sg U8236 ( .A(n4839), .B(n4840), .X(n5838) );
  nand_x1_sg U8237 ( .A(n7411), .B(n7474), .X(n4840) );
  nand_x1_sg U8238 ( .A(n4875), .B(n4876), .X(n5839) );
  nand_x1_sg U8239 ( .A(n7411), .B(n7472), .X(n4876) );
  nand_x1_sg U8240 ( .A(n4755), .B(n4756), .X(n5830) );
  nand_x1_sg U8241 ( .A(n7411), .B(n7478), .X(n4756) );
  nand_x1_sg U8242 ( .A(n4797), .B(n4798), .X(n5834) );
  nand_x1_sg U8243 ( .A(n7411), .B(n7476), .X(n4798) );
  nand_x1_sg U8244 ( .A(n5001), .B(n5002), .X(n5851) );
  nand_x1_sg U8245 ( .A(n7411), .B(n7466), .X(n5002) );
  nand_x1_sg U8246 ( .A(n4125), .B(n4126), .X(n5679) );
  nand_x1_sg U8247 ( .A(n7443), .B(n7456), .X(n4125) );
  nand_x1_sg U8248 ( .A(n4100), .B(n4101), .X(n5667) );
  nand_x1_sg U8249 ( .A(n7488), .B(n7456), .X(n4100) );
  nand_x1_sg U8250 ( .A(n4121), .B(n4122), .X(n5677) );
  nand_x1_sg U8251 ( .A(n7490), .B(n7456), .X(n4121) );
  nand_x1_sg U8252 ( .A(n4127), .B(n4128), .X(n5680) );
  nand_x1_sg U8253 ( .A(n7494), .B(n7456), .X(n4127) );
  nand_x1_sg U8254 ( .A(n4105), .B(n4106), .X(n5669) );
  nand_x1_sg U8255 ( .A(n7492), .B(n7457), .X(n4105) );
  nand_x1_sg U8256 ( .A(n4669), .B(n4670), .X(n5821) );
  nand_x1_sg U8257 ( .A(n7482), .B(n7456), .X(n4669) );
  nand_x1_sg U8258 ( .A(n4115), .B(n4116), .X(n5674) );
  nand_x1_sg U8259 ( .A(n7480), .B(n7456), .X(n4115) );
  nand_x1_sg U8260 ( .A(n4103), .B(n4104), .X(n5668) );
  nand_x1_sg U8261 ( .A(n7484), .B(n7456), .X(n4103) );
  nand_x1_sg U8262 ( .A(n4135), .B(n4136), .X(n5684) );
  nand_x1_sg U8263 ( .A(n7486), .B(n7457), .X(n4135) );
  nand_x1_sg U8264 ( .A(n4129), .B(n4130), .X(n5681) );
  nand_x1_sg U8265 ( .A(n7470), .B(n7457), .X(n4129) );
  nand_x1_sg U8266 ( .A(n4107), .B(n4108), .X(n5670) );
  nand_x1_sg U8267 ( .A(n7468), .B(n7456), .X(n4107) );
  nand_x1_sg U8268 ( .A(n4119), .B(n4120), .X(n5676) );
  nand_x1_sg U8269 ( .A(n7450), .B(n7456), .X(n4119) );
  nand_x1_sg U8270 ( .A(n4131), .B(n4132), .X(n5682) );
  nand_x1_sg U8271 ( .A(n7445), .B(n7456), .X(n4131) );
  nand_x1_sg U8272 ( .A(n4111), .B(n4112), .X(n5672) );
  nand_x1_sg U8273 ( .A(n7452), .B(n7457), .X(n4111) );
  nand_x1_sg U8274 ( .A(n5078), .B(n5079), .X(n5871) );
  nand_x1_sg U8275 ( .A(n7454), .B(n7456), .X(n5078) );
  nand_x1_sg U8276 ( .A(n4117), .B(n4118), .X(n5675) );
  nand_x1_sg U8277 ( .A(n3855), .B(n7457), .X(n4117) );
  nand_x1_sg U8278 ( .A(n4109), .B(n4110), .X(n5671) );
  nand_x1_sg U8279 ( .A(n7472), .B(n7456), .X(n4109) );
  nand_x1_sg U8280 ( .A(n4123), .B(n4124), .X(n5678) );
  nand_x1_sg U8281 ( .A(n7478), .B(n7457), .X(n4123) );
  nand_x1_sg U8282 ( .A(n4113), .B(n4114), .X(n5673) );
  nand_x1_sg U8283 ( .A(n7476), .B(n7456), .X(n4113) );
  nand_x1_sg U8284 ( .A(n4133), .B(n4134), .X(n5683) );
  nand_x1_sg U8285 ( .A(n7466), .B(n7456), .X(n4133) );
  nand_x1_sg U8286 ( .A(n4070), .B(n4071), .X(n5653) );
  nand_x1_sg U8287 ( .A(n7443), .B(n7509), .X(n4070) );
  nand_x1_sg U8288 ( .A(n4060), .B(n4061), .X(n5648) );
  nand_x1_sg U8289 ( .A(n3837), .B(n7509), .X(n4060) );
  nand_x1_sg U8290 ( .A(n4064), .B(n4065), .X(n5650) );
  nand_x1_sg U8291 ( .A(n3885), .B(n7509), .X(n4064) );
  nand_x1_sg U8292 ( .A(n4074), .B(n4075), .X(n5655) );
  nand_x1_sg U8293 ( .A(n7494), .B(n7510), .X(n4074) );
  nand_x1_sg U8294 ( .A(n4076), .B(n4077), .X(n5656) );
  nand_x1_sg U8295 ( .A(n3882), .B(n7509), .X(n4076) );
  nand_x1_sg U8296 ( .A(n4057), .B(n4058), .X(n5647) );
  nand_x1_sg U8297 ( .A(n7482), .B(n7509), .X(n4057) );
  nand_x1_sg U8298 ( .A(n4082), .B(n4083), .X(n5659) );
  nand_x1_sg U8299 ( .A(n7480), .B(n7509), .X(n4082) );
  nand_x1_sg U8300 ( .A(n4084), .B(n4085), .X(n5660) );
  nand_x1_sg U8301 ( .A(n7484), .B(n7509), .X(n4084) );
  nand_x1_sg U8302 ( .A(n4072), .B(n4073), .X(n5654) );
  nand_x1_sg U8303 ( .A(n7486), .B(n7509), .X(n4072) );
  nand_x1_sg U8304 ( .A(n4068), .B(n4069), .X(n5652) );
  nand_x1_sg U8305 ( .A(n7470), .B(n7510), .X(n4068) );
  nand_x1_sg U8306 ( .A(n4078), .B(n4079), .X(n5657) );
  nand_x1_sg U8307 ( .A(n7468), .B(n7509), .X(n4078) );
  nand_x1_sg U8308 ( .A(n4086), .B(n4087), .X(n5661) );
  nand_x1_sg U8309 ( .A(n7450), .B(n7510), .X(n4086) );
  nand_x1_sg U8310 ( .A(n4088), .B(n4089), .X(n5662) );
  nand_x1_sg U8311 ( .A(n7445), .B(n7509), .X(n4088) );
  nand_x1_sg U8312 ( .A(n4090), .B(n4091), .X(n5663) );
  nand_x1_sg U8313 ( .A(n3858), .B(n7509), .X(n4090) );
  nand_x1_sg U8314 ( .A(n4080), .B(n4081), .X(n5658) );
  nand_x1_sg U8315 ( .A(n7454), .B(n7510), .X(n4080) );
  nand_x1_sg U8316 ( .A(n4092), .B(n4093), .X(n5664) );
  nand_x1_sg U8317 ( .A(n7474), .B(n7510), .X(n4092) );
  nand_x1_sg U8318 ( .A(n4062), .B(n4063), .X(n5649) );
  nand_x1_sg U8319 ( .A(n7472), .B(n7510), .X(n4062) );
  nand_x1_sg U8320 ( .A(n4066), .B(n4067), .X(n5651) );
  nand_x1_sg U8321 ( .A(n7478), .B(n7509), .X(n4066) );
  nand_x1_sg U8322 ( .A(n4094), .B(n4095), .X(n5665) );
  nand_x1_sg U8323 ( .A(n7476), .B(n7509), .X(n4094) );
  nand_x1_sg U8324 ( .A(n4096), .B(n4097), .X(n5666) );
  nand_x1_sg U8325 ( .A(n7466), .B(n7509), .X(n4096) );
  nand_x1_sg U8326 ( .A(n3940), .B(n3941), .X(n5591) );
  nand_x1_sg U8327 ( .A(n7414), .B(n7443), .X(n3941) );
  nand_x1_sg U8328 ( .A(n3942), .B(n3943), .X(n5592) );
  nand_x1_sg U8329 ( .A(n7414), .B(n7488), .X(n3943) );
  nand_x1_sg U8330 ( .A(n3936), .B(n3937), .X(n5589) );
  nand_x1_sg U8331 ( .A(n7414), .B(n7490), .X(n3937) );
  nand_x1_sg U8332 ( .A(n3962), .B(n3963), .X(n5602) );
  nand_x1_sg U8333 ( .A(n7414), .B(n7494), .X(n3963) );
  nand_x1_sg U8334 ( .A(n3970), .B(n3971), .X(n5606) );
  nand_x1_sg U8335 ( .A(n7414), .B(n7492), .X(n3971) );
  nand_x1_sg U8336 ( .A(n3954), .B(n3955), .X(n5598) );
  nand_x1_sg U8337 ( .A(n7414), .B(n7482), .X(n3955) );
  nand_x1_sg U8338 ( .A(n3933), .B(n3934), .X(n5588) );
  nand_x1_sg U8339 ( .A(n7414), .B(n7480), .X(n3934) );
  nand_x1_sg U8340 ( .A(n3960), .B(n3961), .X(n5601) );
  nand_x1_sg U8341 ( .A(n7414), .B(n7484), .X(n3961) );
  nand_x1_sg U8342 ( .A(n3964), .B(n3965), .X(n5603) );
  nand_x1_sg U8343 ( .A(n7414), .B(n7486), .X(n3965) );
  nand_x1_sg U8344 ( .A(n3966), .B(n3967), .X(n5604) );
  nand_x1_sg U8345 ( .A(n7414), .B(n7470), .X(n3967) );
  nand_x1_sg U8346 ( .A(n3952), .B(n3953), .X(n5597) );
  nand_x1_sg U8347 ( .A(n7414), .B(n7468), .X(n3953) );
  nand_x1_sg U8348 ( .A(n3950), .B(n3951), .X(n5596) );
  nand_x1_sg U8349 ( .A(n7414), .B(n7450), .X(n3951) );
  nand_x1_sg U8350 ( .A(n3958), .B(n3959), .X(n5600) );
  nand_x1_sg U8351 ( .A(n7414), .B(n7445), .X(n3959) );
  nand_x1_sg U8352 ( .A(n3948), .B(n3949), .X(n5595) );
  nand_x1_sg U8353 ( .A(n7414), .B(n7452), .X(n3949) );
  nand_x1_sg U8354 ( .A(n3972), .B(n3973), .X(n5607) );
  nand_x1_sg U8355 ( .A(n7414), .B(n7454), .X(n3973) );
  nand_x1_sg U8356 ( .A(n3938), .B(n3939), .X(n5590) );
  nand_x1_sg U8357 ( .A(n7414), .B(n7474), .X(n3939) );
  nand_x1_sg U8358 ( .A(n3944), .B(n3945), .X(n5593) );
  nand_x1_sg U8359 ( .A(n7414), .B(n7472), .X(n3945) );
  nand_x1_sg U8360 ( .A(n3956), .B(n3957), .X(n5599) );
  nand_x1_sg U8361 ( .A(n7414), .B(n7478), .X(n3957) );
  nand_x1_sg U8362 ( .A(n3946), .B(n3947), .X(n5594) );
  nand_x1_sg U8363 ( .A(n7414), .B(n7476), .X(n3947) );
  nand_x1_sg U8364 ( .A(n3968), .B(n3969), .X(n5605) );
  nand_x1_sg U8365 ( .A(n7414), .B(n7466), .X(n3969) );
  nand_x1_sg U8366 ( .A(n4004), .B(n4005), .X(n5622) );
  nand_x1_sg U8367 ( .A(n7413), .B(n7443), .X(n4005) );
  nand_x1_sg U8368 ( .A(n3996), .B(n3997), .X(n5618) );
  nand_x1_sg U8369 ( .A(n7413), .B(n7488), .X(n3997) );
  nand_x1_sg U8370 ( .A(n4014), .B(n4015), .X(n5627) );
  nand_x1_sg U8371 ( .A(n7413), .B(n7490), .X(n4015) );
  nand_x1_sg U8372 ( .A(n3988), .B(n3989), .X(n5614) );
  nand_x1_sg U8373 ( .A(n7413), .B(n7494), .X(n3989) );
  nand_x1_sg U8374 ( .A(n3975), .B(n3976), .X(n5608) );
  nand_x1_sg U8375 ( .A(n7413), .B(n7492), .X(n3976) );
  nand_x1_sg U8376 ( .A(n3990), .B(n3991), .X(n5615) );
  nand_x1_sg U8377 ( .A(n7413), .B(n7482), .X(n3991) );
  nand_x1_sg U8378 ( .A(n3982), .B(n3983), .X(n5611) );
  nand_x1_sg U8379 ( .A(n7413), .B(n7480), .X(n3983) );
  nand_x1_sg U8380 ( .A(n4008), .B(n4009), .X(n5624) );
  nand_x1_sg U8381 ( .A(n7413), .B(n7484), .X(n4009) );
  nand_x1_sg U8382 ( .A(n4002), .B(n4003), .X(n5621) );
  nand_x1_sg U8383 ( .A(n7413), .B(n7486), .X(n4003) );
  nand_x1_sg U8384 ( .A(n4012), .B(n4013), .X(n5626) );
  nand_x1_sg U8385 ( .A(n7413), .B(n7470), .X(n4013) );
  nand_x1_sg U8386 ( .A(n3992), .B(n3993), .X(n5616) );
  nand_x1_sg U8387 ( .A(n7413), .B(n7468), .X(n3993) );
  nand_x1_sg U8388 ( .A(n3986), .B(n3987), .X(n5613) );
  nand_x1_sg U8389 ( .A(n7413), .B(n7450), .X(n3987) );
  nand_x1_sg U8390 ( .A(n3978), .B(n3979), .X(n5609) );
  nand_x1_sg U8391 ( .A(n7413), .B(n7445), .X(n3979) );
  nand_x1_sg U8392 ( .A(n3994), .B(n3995), .X(n5617) );
  nand_x1_sg U8393 ( .A(n7413), .B(n7452), .X(n3995) );
  nand_x1_sg U8394 ( .A(n3984), .B(n3985), .X(n5612) );
  nand_x1_sg U8395 ( .A(n7413), .B(n7454), .X(n3985) );
  nand_x1_sg U8396 ( .A(n3980), .B(n3981), .X(n5610) );
  nand_x1_sg U8397 ( .A(n7413), .B(n7474), .X(n3981) );
  nand_x1_sg U8398 ( .A(n3998), .B(n3999), .X(n5619) );
  nand_x1_sg U8399 ( .A(n7413), .B(n7472), .X(n3999) );
  nand_x1_sg U8400 ( .A(n4006), .B(n4007), .X(n5623) );
  nand_x1_sg U8401 ( .A(n7413), .B(n7478), .X(n4007) );
  nand_x1_sg U8402 ( .A(n4000), .B(n4001), .X(n5620) );
  nand_x1_sg U8403 ( .A(n7413), .B(n7476), .X(n4001) );
  nand_x1_sg U8404 ( .A(n4010), .B(n4011), .X(n5625) );
  nand_x1_sg U8405 ( .A(n7413), .B(n7466), .X(n4011) );
  nand_x1_sg U8406 ( .A(n4315), .B(n4316), .X(n5756) );
  nand_x1_sg U8407 ( .A(n7443), .B(n7499), .X(n4316) );
  nand_x1_sg U8408 ( .A(n4323), .B(n4324), .X(n5760) );
  nand_x1_sg U8409 ( .A(n7488), .B(n7499), .X(n4324) );
  nand_x1_sg U8410 ( .A(n4317), .B(n4318), .X(n5757) );
  nand_x1_sg U8411 ( .A(n7490), .B(n7499), .X(n4318) );
  nand_x1_sg U8412 ( .A(n4327), .B(n4328), .X(n5762) );
  nand_x1_sg U8413 ( .A(n7494), .B(n7499), .X(n4328) );
  nand_x1_sg U8414 ( .A(n4313), .B(n4314), .X(n5755) );
  nand_x1_sg U8415 ( .A(n7492), .B(n7500), .X(n4314) );
  nand_x1_sg U8416 ( .A(n4308), .B(n4309), .X(n5753) );
  nand_x1_sg U8417 ( .A(n7482), .B(n7499), .X(n4309) );
  nand_x1_sg U8418 ( .A(n4329), .B(n4330), .X(n5763) );
  nand_x1_sg U8419 ( .A(n7480), .B(n7499), .X(n4330) );
  nand_x1_sg U8420 ( .A(n4339), .B(n4340), .X(n5768) );
  nand_x1_sg U8421 ( .A(n7484), .B(n7499), .X(n4340) );
  nand_x1_sg U8422 ( .A(n4341), .B(n4342), .X(n5769) );
  nand_x1_sg U8423 ( .A(n7486), .B(n7499), .X(n4342) );
  nand_x1_sg U8424 ( .A(n4337), .B(n4338), .X(n5767) );
  nand_x1_sg U8425 ( .A(n7470), .B(n7500), .X(n4338) );
  nand_x1_sg U8426 ( .A(n4319), .B(n4320), .X(n5758) );
  nand_x1_sg U8427 ( .A(n7468), .B(n7500), .X(n4320) );
  nand_x1_sg U8428 ( .A(n4343), .B(n4344), .X(n5770) );
  nand_x1_sg U8429 ( .A(n7450), .B(n7500), .X(n4344) );
  nand_x1_sg U8430 ( .A(n4321), .B(n4322), .X(n5759) );
  nand_x1_sg U8431 ( .A(n7445), .B(n7499), .X(n4322) );
  nand_x1_sg U8432 ( .A(n4331), .B(n4332), .X(n5764) );
  nand_x1_sg U8433 ( .A(n7452), .B(n7500), .X(n4332) );
  nand_x1_sg U8434 ( .A(n4347), .B(n4348), .X(n5772) );
  nand_x1_sg U8435 ( .A(n7454), .B(n7499), .X(n4348) );
  nand_x1_sg U8436 ( .A(n4333), .B(n4334), .X(n5765) );
  nand_x1_sg U8437 ( .A(n7474), .B(n7499), .X(n4334) );
  nand_x1_sg U8438 ( .A(n4311), .B(n4312), .X(n5754) );
  nand_x1_sg U8439 ( .A(n7472), .B(n7499), .X(n4312) );
  nand_x1_sg U8440 ( .A(n4325), .B(n4326), .X(n5761) );
  nand_x1_sg U8441 ( .A(n7478), .B(n7500), .X(n4326) );
  nand_x1_sg U8442 ( .A(n4345), .B(n4346), .X(n5771) );
  nand_x1_sg U8443 ( .A(n7476), .B(n7499), .X(n4346) );
  nand_x1_sg U8444 ( .A(n4335), .B(n4336), .X(n5766) );
  nand_x1_sg U8445 ( .A(n7466), .B(n7499), .X(n4336) );
  nand_x1_sg U8446 ( .A(n4144), .B(n4145), .X(n5688) );
  nand_x1_sg U8447 ( .A(n7443), .B(n7507), .X(n4145) );
  nand_x1_sg U8448 ( .A(n4152), .B(n4153), .X(n5692) );
  nand_x1_sg U8449 ( .A(n7488), .B(n7506), .X(n4153) );
  nand_x1_sg U8450 ( .A(n4146), .B(n4147), .X(n5689) );
  nand_x1_sg U8451 ( .A(n7490), .B(n7506), .X(n4147) );
  nand_x1_sg U8452 ( .A(n4156), .B(n4157), .X(n5694) );
  nand_x1_sg U8453 ( .A(n7494), .B(n7507), .X(n4157) );
  nand_x1_sg U8454 ( .A(n4142), .B(n4143), .X(n5687) );
  nand_x1_sg U8455 ( .A(n7492), .B(n7507), .X(n4143) );
  nand_x1_sg U8456 ( .A(n4137), .B(n4138), .X(n5685) );
  nand_x1_sg U8457 ( .A(n7482), .B(n7507), .X(n4138) );
  nand_x1_sg U8458 ( .A(n4158), .B(n4159), .X(n5695) );
  nand_x1_sg U8459 ( .A(n3843), .B(n7506), .X(n4159) );
  nand_x1_sg U8460 ( .A(n4168), .B(n4169), .X(n5700) );
  nand_x1_sg U8461 ( .A(n7484), .B(n7507), .X(n4169) );
  nand_x1_sg U8462 ( .A(n4170), .B(n4171), .X(n5701) );
  nand_x1_sg U8463 ( .A(n7486), .B(n7506), .X(n4171) );
  nand_x1_sg U8464 ( .A(n4166), .B(n4167), .X(n5699) );
  nand_x1_sg U8465 ( .A(n3876), .B(n7506), .X(n4167) );
  nand_x1_sg U8466 ( .A(n4148), .B(n4149), .X(n5690) );
  nand_x1_sg U8467 ( .A(n7468), .B(n7506), .X(n4149) );
  nand_x1_sg U8468 ( .A(n4172), .B(n4173), .X(n5702) );
  nand_x1_sg U8469 ( .A(n7450), .B(n4139), .X(n4173) );
  nand_x1_sg U8470 ( .A(n4150), .B(n4151), .X(n5691) );
  nand_x1_sg U8471 ( .A(n7445), .B(n7507), .X(n4151) );
  nand_x1_sg U8472 ( .A(n4160), .B(n4161), .X(n5696) );
  nand_x1_sg U8473 ( .A(n7452), .B(n7507), .X(n4161) );
  nand_x1_sg U8474 ( .A(n4176), .B(n4177), .X(n5704) );
  nand_x1_sg U8475 ( .A(n7454), .B(n7506), .X(n4177) );
  nand_x1_sg U8476 ( .A(n4162), .B(n4163), .X(n5697) );
  nand_x1_sg U8477 ( .A(n7474), .B(n7507), .X(n4163) );
  nand_x1_sg U8478 ( .A(n4140), .B(n4141), .X(n5686) );
  nand_x1_sg U8479 ( .A(n7472), .B(n7506), .X(n4141) );
  nand_x1_sg U8480 ( .A(n4154), .B(n4155), .X(n5693) );
  nand_x1_sg U8481 ( .A(n3867), .B(n7507), .X(n4155) );
  nand_x1_sg U8482 ( .A(n4174), .B(n4175), .X(n5703) );
  nand_x1_sg U8483 ( .A(n7476), .B(n7507), .X(n4175) );
  nand_x1_sg U8484 ( .A(n4164), .B(n4165), .X(n5698) );
  nand_x1_sg U8485 ( .A(n7466), .B(n7506), .X(n4165) );
  nand_x1_sg U8486 ( .A(n3862), .B(n3863), .X(n5560) );
  nand_x1_sg U8487 ( .A(n7443), .B(n7418), .X(n3863) );
  nand_x1_sg U8488 ( .A(n3835), .B(n3836), .X(n5551) );
  nand_x1_sg U8489 ( .A(n7488), .B(n7418), .X(n3836) );
  nand_x1_sg U8490 ( .A(n3883), .B(n3884), .X(n5567) );
  nand_x1_sg U8491 ( .A(n7490), .B(n7418), .X(n3884) );
  nand_x1_sg U8492 ( .A(n3829), .B(n3830), .X(n5549) );
  nand_x1_sg U8493 ( .A(n7494), .B(n7418), .X(n3830) );
  nand_x1_sg U8494 ( .A(n3880), .B(n3881), .X(n5566) );
  nand_x1_sg U8495 ( .A(n7492), .B(n7418), .X(n3881) );
  nand_x1_sg U8496 ( .A(n3850), .B(n3851), .X(n5556) );
  nand_x1_sg U8497 ( .A(n3852), .B(n7418), .X(n3851) );
  nand_x1_sg U8498 ( .A(n3841), .B(n3842), .X(n5553) );
  nand_x1_sg U8499 ( .A(n7480), .B(n7418), .X(n3842) );
  nand_x1_sg U8500 ( .A(n3871), .B(n3872), .X(n5563) );
  nand_x1_sg U8501 ( .A(n7484), .B(n7418), .X(n3872) );
  nand_x1_sg U8502 ( .A(n3859), .B(n3860), .X(n5559) );
  nand_x1_sg U8503 ( .A(n7486), .B(n7418), .X(n3860) );
  nand_x1_sg U8504 ( .A(n3874), .B(n3875), .X(n5564) );
  nand_x1_sg U8505 ( .A(n7470), .B(n7418), .X(n3875) );
  nand_x1_sg U8506 ( .A(n3832), .B(n3833), .X(n5550) );
  nand_x1_sg U8507 ( .A(n7468), .B(n7418), .X(n3833) );
  nand_x1_sg U8508 ( .A(n3847), .B(n3848), .X(n5555) );
  nand_x1_sg U8509 ( .A(n7450), .B(n7418), .X(n3848) );
  nand_x1_sg U8510 ( .A(n3868), .B(n3869), .X(n5562) );
  nand_x1_sg U8511 ( .A(n7445), .B(n7418), .X(n3869) );
  nand_x1_sg U8512 ( .A(n3856), .B(n3857), .X(n5558) );
  nand_x1_sg U8513 ( .A(n7452), .B(n7418), .X(n3857) );
  nand_x1_sg U8514 ( .A(n3844), .B(n3845), .X(n5554) );
  nand_x1_sg U8515 ( .A(n7454), .B(n7418), .X(n3845) );
  nand_x1_sg U8516 ( .A(n3853), .B(n3854), .X(n5557) );
  nand_x1_sg U8517 ( .A(n7474), .B(n7418), .X(n3854) );
  nand_x1_sg U8518 ( .A(n3838), .B(n3839), .X(n5552) );
  nand_x1_sg U8519 ( .A(n7472), .B(n7418), .X(n3839) );
  nand_x1_sg U8520 ( .A(n3865), .B(n3866), .X(n5561) );
  nand_x1_sg U8521 ( .A(n7478), .B(n7418), .X(n3866) );
  nand_x1_sg U8522 ( .A(n3825), .B(n3826), .X(n5548) );
  nand_x1_sg U8523 ( .A(n7476), .B(n7418), .X(n3826) );
  nand_x1_sg U8524 ( .A(n3877), .B(n3878), .X(n5565) );
  nand_x1_sg U8525 ( .A(n7466), .B(n7418), .X(n3878) );
  nand_x1_sg U8526 ( .A(n3926), .B(n3927), .X(n5587) );
  nand_x1_sg U8527 ( .A(n7417), .B(n7443), .X(n3927) );
  nand_x1_sg U8528 ( .A(n3910), .B(n3911), .X(n5579) );
  nand_x1_sg U8529 ( .A(n7417), .B(n7488), .X(n3911) );
  nand_x1_sg U8530 ( .A(n3918), .B(n3919), .X(n5583) );
  nand_x1_sg U8531 ( .A(n7417), .B(n7490), .X(n3919) );
  nand_x1_sg U8532 ( .A(n3890), .B(n3891), .X(n5569) );
  nand_x1_sg U8533 ( .A(n7417), .B(n7494), .X(n3891) );
  nand_x1_sg U8534 ( .A(n3924), .B(n3925), .X(n5586) );
  nand_x1_sg U8535 ( .A(n7417), .B(n7492), .X(n3925) );
  nand_x1_sg U8536 ( .A(n3896), .B(n3897), .X(n5572) );
  nand_x1_sg U8537 ( .A(n7417), .B(n7482), .X(n3897) );
  nand_x1_sg U8538 ( .A(n3914), .B(n3915), .X(n5581) );
  nand_x1_sg U8539 ( .A(n7417), .B(n7480), .X(n3915) );
  nand_x1_sg U8540 ( .A(n3908), .B(n3909), .X(n5578) );
  nand_x1_sg U8541 ( .A(n7417), .B(n7484), .X(n3909) );
  nand_x1_sg U8542 ( .A(n3894), .B(n3895), .X(n5571) );
  nand_x1_sg U8543 ( .A(n7417), .B(n7486), .X(n3895) );
  nand_x1_sg U8544 ( .A(n3920), .B(n3921), .X(n5584) );
  nand_x1_sg U8545 ( .A(n7417), .B(n7470), .X(n3921) );
  nand_x1_sg U8546 ( .A(n3892), .B(n3893), .X(n5570) );
  nand_x1_sg U8547 ( .A(n7417), .B(n7468), .X(n3893) );
  nand_x1_sg U8548 ( .A(n3916), .B(n3917), .X(n5582) );
  nand_x1_sg U8549 ( .A(n7417), .B(n7450), .X(n3917) );
  nand_x1_sg U8550 ( .A(n3906), .B(n3907), .X(n5577) );
  nand_x1_sg U8551 ( .A(n7417), .B(n7445), .X(n3907) );
  nand_x1_sg U8552 ( .A(n3900), .B(n3901), .X(n5574) );
  nand_x1_sg U8553 ( .A(n7417), .B(n7452), .X(n3901) );
  nand_x1_sg U8554 ( .A(n3902), .B(n3903), .X(n5575) );
  nand_x1_sg U8555 ( .A(n7417), .B(n7454), .X(n3903) );
  nand_x1_sg U8556 ( .A(n3898), .B(n3899), .X(n5573) );
  nand_x1_sg U8557 ( .A(n7417), .B(n7474), .X(n3899) );
  nand_x1_sg U8558 ( .A(n3912), .B(n3913), .X(n5580) );
  nand_x1_sg U8559 ( .A(n7417), .B(n7472), .X(n3913) );
  nand_x1_sg U8560 ( .A(n3904), .B(n3905), .X(n5576) );
  nand_x1_sg U8561 ( .A(n7417), .B(n7478), .X(n3905) );
  nand_x1_sg U8562 ( .A(n3887), .B(n3888), .X(n5568) );
  nand_x1_sg U8563 ( .A(n7417), .B(n7476), .X(n3888) );
  nand_x1_sg U8564 ( .A(n3922), .B(n3923), .X(n5585) );
  nand_x1_sg U8565 ( .A(n7417), .B(n7466), .X(n3923) );
  nand_x1_sg U8566 ( .A(n4055), .B(n4056), .X(n5646) );
  nand_x1_sg U8567 ( .A(n7443), .B(n7447), .X(n4055) );
  nand_x1_sg U8568 ( .A(n4018), .B(n4019), .X(n5628) );
  nand_x1_sg U8569 ( .A(n7488), .B(n7447), .X(n4018) );
  nand_x1_sg U8570 ( .A(n4039), .B(n4040), .X(n5638) );
  nand_x1_sg U8571 ( .A(n7490), .B(n7447), .X(n4039) );
  nand_x1_sg U8572 ( .A(n4035), .B(n4036), .X(n5636) );
  nand_x1_sg U8573 ( .A(n7494), .B(n7448), .X(n4035) );
  nand_x1_sg U8574 ( .A(n4021), .B(n4022), .X(n5629) );
  nand_x1_sg U8575 ( .A(n7492), .B(n7447), .X(n4021) );
  nand_x1_sg U8576 ( .A(n4041), .B(n4042), .X(n5639) );
  nand_x1_sg U8577 ( .A(n7482), .B(n7448), .X(n4041) );
  nand_x1_sg U8578 ( .A(n4051), .B(n4052), .X(n5644) );
  nand_x1_sg U8579 ( .A(n7480), .B(n7447), .X(n4051) );
  nand_x1_sg U8580 ( .A(n4023), .B(n4024), .X(n5630) );
  nand_x1_sg U8581 ( .A(n7484), .B(n7448), .X(n4023) );
  nand_x1_sg U8582 ( .A(n4043), .B(n4044), .X(n5640) );
  nand_x1_sg U8583 ( .A(n7486), .B(n7447), .X(n4043) );
  nand_x1_sg U8584 ( .A(n4037), .B(n4038), .X(n5637) );
  nand_x1_sg U8585 ( .A(n7470), .B(n7447), .X(n4037) );
  nand_x1_sg U8586 ( .A(n4025), .B(n4026), .X(n5631) );
  nand_x1_sg U8587 ( .A(n7468), .B(n7447), .X(n4025) );
  nand_x1_sg U8588 ( .A(n4045), .B(n4046), .X(n5641) );
  nand_x1_sg U8589 ( .A(n7450), .B(n7447), .X(n4045) );
  nand_x1_sg U8590 ( .A(n5187), .B(n5188), .X(n5874) );
  nand_x1_sg U8591 ( .A(n7445), .B(n7447), .X(n5187) );
  nand_x1_sg U8592 ( .A(n4027), .B(n4028), .X(n5632) );
  nand_x1_sg U8593 ( .A(n7452), .B(n7447), .X(n4027) );
  nand_x1_sg U8594 ( .A(n4033), .B(n4034), .X(n5635) );
  nand_x1_sg U8595 ( .A(n3846), .B(n7447), .X(n4033) );
  nand_x1_sg U8596 ( .A(n4053), .B(n4054), .X(n5645) );
  nand_x1_sg U8597 ( .A(n7474), .B(n7448), .X(n4053) );
  nand_x1_sg U8598 ( .A(n4029), .B(n4030), .X(n5633) );
  nand_x1_sg U8599 ( .A(n7472), .B(n7448), .X(n4029) );
  nand_x1_sg U8600 ( .A(n4047), .B(n4048), .X(n5642) );
  nand_x1_sg U8601 ( .A(n7478), .B(n7448), .X(n4047) );
  nand_x1_sg U8602 ( .A(n4031), .B(n4032), .X(n5634) );
  nand_x1_sg U8603 ( .A(n7476), .B(n7447), .X(n4031) );
  nand_x1_sg U8604 ( .A(n4049), .B(n4050), .X(n5643) );
  nand_x1_sg U8605 ( .A(n7466), .B(n7447), .X(n4049) );
  nand_x1_sg U8606 ( .A(n5227), .B(n5228), .X(n5876) );
  nand_x1_sg U8607 ( .A(n3864), .B(n7421), .X(n5228) );
  nand_x1_sg U8608 ( .A(n4539), .B(n4540), .X(n5807) );
  nand_x1_sg U8609 ( .A(n7488), .B(n7421), .X(n4540) );
  nand_x1_sg U8610 ( .A(n4497), .B(n4498), .X(n5803) );
  nand_x1_sg U8611 ( .A(n7490), .B(n7422), .X(n4498) );
  nand_x1_sg U8612 ( .A(n4405), .B(n4406), .X(n5797) );
  nand_x1_sg U8613 ( .A(n3831), .B(n7421), .X(n4406) );
  nand_x1_sg U8614 ( .A(n4455), .B(n4456), .X(n5799) );
  nand_x1_sg U8615 ( .A(n7492), .B(n7421), .X(n4456) );
  nand_x1_sg U8616 ( .A(n4665), .B(n4666), .X(n5819) );
  nand_x1_sg U8617 ( .A(n7482), .B(n7421), .X(n4666) );
  nand_x1_sg U8618 ( .A(n4711), .B(n4712), .X(n5825) );
  nand_x1_sg U8619 ( .A(n7480), .B(n7421), .X(n4712) );
  nand_x1_sg U8620 ( .A(n4623), .B(n4624), .X(n5815) );
  nand_x1_sg U8621 ( .A(n7484), .B(n7422), .X(n4624) );
  nand_x1_sg U8622 ( .A(n4583), .B(n4584), .X(n5812) );
  nand_x1_sg U8623 ( .A(n7486), .B(n7421), .X(n4584) );
  nand_x1_sg U8624 ( .A(n4921), .B(n4922), .X(n5845) );
  nand_x1_sg U8625 ( .A(n7470), .B(n7421), .X(n4922) );
  nand_x1_sg U8626 ( .A(n4961), .B(n4962), .X(n5848) );
  nand_x1_sg U8627 ( .A(n7468), .B(n7421), .X(n4962) );
  nand_x1_sg U8628 ( .A(n5151), .B(n5152), .X(n5873) );
  nand_x1_sg U8629 ( .A(n3849), .B(n7422), .X(n5152) );
  nand_x1_sg U8630 ( .A(n5191), .B(n5192), .X(n5875) );
  nand_x1_sg U8631 ( .A(n3870), .B(n7421), .X(n5192) );
  nand_x1_sg U8632 ( .A(n5115), .B(n5116), .X(n5872) );
  nand_x1_sg U8633 ( .A(n7452), .B(n7421), .X(n5116) );
  nand_x1_sg U8634 ( .A(n5076), .B(n5077), .X(n5870) );
  nand_x1_sg U8635 ( .A(n7454), .B(n7421), .X(n5077) );
  nand_x1_sg U8636 ( .A(n4837), .B(n4838), .X(n5837) );
  nand_x1_sg U8637 ( .A(n7474), .B(n7421), .X(n4838) );
  nand_x1_sg U8638 ( .A(n4877), .B(n4878), .X(n5840) );
  nand_x1_sg U8639 ( .A(n3840), .B(n7422), .X(n4878) );
  nand_x1_sg U8640 ( .A(n4753), .B(n4754), .X(n5829) );
  nand_x1_sg U8641 ( .A(n7478), .B(n7422), .X(n4754) );
  nand_x1_sg U8642 ( .A(n4795), .B(n4796), .X(n5833) );
  nand_x1_sg U8643 ( .A(n7476), .B(n7421), .X(n4796) );
  nand_x1_sg U8644 ( .A(n5003), .B(n5004), .X(n5852) );
  nand_x1_sg U8645 ( .A(n7466), .B(n7422), .X(n5004) );
  nand_x1_sg U8646 ( .A(n5293), .B(n9201), .X(n5881) );
  inv_x1_sg U8647 ( .A(n5294), .X(n9201) );
  nand_x1_sg U8648 ( .A(n5270), .B(n5271), .X(n5877) );
  nand_x1_sg U8649 ( .A(n5272), .B(n5273), .X(n5271) );
  nand_x1_sg U8650 ( .A(n7520), .B(n5275), .X(n5270) );
  nand_x1_sg U8651 ( .A(n5308), .B(n5309), .X(n5885) );
  nand_x1_sg U8652 ( .A(n3805), .B(n3806), .X(\update_mask_0/n1129 ) );
  nand_x1_sg U8653 ( .A(n7530), .B(\i_im[15][19] ), .X(n3805) );
  nand_x1_sg U8654 ( .A(n3803), .B(n3804), .X(\update_mask_0/n1130 ) );
  nand_x1_sg U8655 ( .A(n7531), .B(\i_im[15][18] ), .X(n3803) );
  nand_x1_sg U8656 ( .A(n3801), .B(n3802), .X(\update_mask_0/n1131 ) );
  nand_x1_sg U8657 ( .A(n7529), .B(\i_im[15][17] ), .X(n3801) );
  nand_x1_sg U8658 ( .A(n3799), .B(n3800), .X(\update_mask_0/n1132 ) );
  nand_x1_sg U8659 ( .A(n7531), .B(\i_im[15][16] ), .X(n3799) );
  nand_x1_sg U8660 ( .A(n3797), .B(n3798), .X(\update_mask_0/n1133 ) );
  nand_x1_sg U8661 ( .A(n7530), .B(\i_im[15][15] ), .X(n3797) );
  nand_x1_sg U8662 ( .A(n3795), .B(n3796), .X(\update_mask_0/n1134 ) );
  nand_x1_sg U8663 ( .A(n7528), .B(\i_im[15][14] ), .X(n3795) );
  nand_x1_sg U8664 ( .A(n3793), .B(n3794), .X(\update_mask_0/n1135 ) );
  nand_x1_sg U8665 ( .A(n7534), .B(\i_im[15][13] ), .X(n3793) );
  nand_x1_sg U8666 ( .A(n3791), .B(n3792), .X(\update_mask_0/n1136 ) );
  nand_x1_sg U8667 ( .A(n7534), .B(\i_im[15][12] ), .X(n3791) );
  nand_x1_sg U8668 ( .A(n3789), .B(n3790), .X(\update_mask_0/n1137 ) );
  nand_x1_sg U8669 ( .A(n7534), .B(\i_im[15][11] ), .X(n3789) );
  nand_x1_sg U8670 ( .A(n3787), .B(n3788), .X(\update_mask_0/n1138 ) );
  nand_x1_sg U8671 ( .A(n7534), .B(\i_im[15][10] ), .X(n3787) );
  nand_x1_sg U8672 ( .A(n3785), .B(n3786), .X(\update_mask_0/n1139 ) );
  nand_x1_sg U8673 ( .A(n7534), .B(\i_im[15][9] ), .X(n3785) );
  nand_x1_sg U8674 ( .A(n3783), .B(n3784), .X(\update_mask_0/n1140 ) );
  nand_x1_sg U8675 ( .A(n7533), .B(\i_im[15][8] ), .X(n3783) );
  nand_x1_sg U8676 ( .A(n3781), .B(n3782), .X(\update_mask_0/n1141 ) );
  nand_x1_sg U8677 ( .A(n7530), .B(\i_im[15][7] ), .X(n3781) );
  nand_x1_sg U8678 ( .A(n3779), .B(n3780), .X(\update_mask_0/n1142 ) );
  nand_x1_sg U8679 ( .A(n7527), .B(\i_im[15][6] ), .X(n3779) );
  nand_x1_sg U8680 ( .A(n3777), .B(n3778), .X(\update_mask_0/n1143 ) );
  nand_x1_sg U8681 ( .A(n7528), .B(\i_im[15][5] ), .X(n3777) );
  nand_x1_sg U8682 ( .A(n3775), .B(n3776), .X(\update_mask_0/n1144 ) );
  nand_x1_sg U8683 ( .A(n7531), .B(\i_im[15][4] ), .X(n3775) );
  nand_x1_sg U8684 ( .A(n3773), .B(n3774), .X(\update_mask_0/n1145 ) );
  nand_x1_sg U8685 ( .A(n7533), .B(\i_im[15][3] ), .X(n3773) );
  nand_x1_sg U8686 ( .A(n3771), .B(n3772), .X(\update_mask_0/n1146 ) );
  nand_x1_sg U8687 ( .A(n7529), .B(\i_im[15][2] ), .X(n3771) );
  nand_x1_sg U8688 ( .A(n3769), .B(n3770), .X(\update_mask_0/n1147 ) );
  nand_x1_sg U8689 ( .A(n7529), .B(\i_im[15][1] ), .X(n3769) );
  nand_x1_sg U8690 ( .A(n3767), .B(n3768), .X(\update_mask_0/n1148 ) );
  nand_x1_sg U8691 ( .A(n7530), .B(\i_im[15][0] ), .X(n3767) );
  nand_x1_sg U8692 ( .A(n3765), .B(n3766), .X(\update_mask_0/n1149 ) );
  nand_x1_sg U8693 ( .A(n7531), .B(\i_im[14][19] ), .X(n3765) );
  nand_x1_sg U8694 ( .A(n3763), .B(n3764), .X(\update_mask_0/n1150 ) );
  nand_x1_sg U8695 ( .A(n7535), .B(\i_im[14][18] ), .X(n3763) );
  nand_x1_sg U8696 ( .A(n3761), .B(n3762), .X(\update_mask_0/n1151 ) );
  nand_x1_sg U8697 ( .A(n7530), .B(\i_im[14][17] ), .X(n3761) );
  nand_x1_sg U8698 ( .A(n3759), .B(n3760), .X(\update_mask_0/n1152 ) );
  nand_x1_sg U8699 ( .A(n7535), .B(\i_im[14][16] ), .X(n3759) );
  nand_x1_sg U8700 ( .A(n3757), .B(n3758), .X(\update_mask_0/n1153 ) );
  nand_x1_sg U8701 ( .A(n7534), .B(\i_im[14][15] ), .X(n3757) );
  nand_x1_sg U8702 ( .A(n3755), .B(n3756), .X(\update_mask_0/n1154 ) );
  nand_x1_sg U8703 ( .A(n7529), .B(\i_im[14][14] ), .X(n3755) );
  nand_x1_sg U8704 ( .A(n3753), .B(n3754), .X(\update_mask_0/n1155 ) );
  nand_x1_sg U8705 ( .A(n7534), .B(\i_im[14][13] ), .X(n3753) );
  nand_x1_sg U8706 ( .A(n3751), .B(n3752), .X(\update_mask_0/n1156 ) );
  nand_x1_sg U8707 ( .A(n7534), .B(\i_im[14][12] ), .X(n3751) );
  nand_x1_sg U8708 ( .A(n3749), .B(n3750), .X(\update_mask_0/n1157 ) );
  nand_x1_sg U8709 ( .A(n7527), .B(\i_im[14][11] ), .X(n3749) );
  nand_x1_sg U8710 ( .A(n3747), .B(n3748), .X(\update_mask_0/n1158 ) );
  nand_x1_sg U8711 ( .A(n7528), .B(\i_im[14][10] ), .X(n3747) );
  nand_x1_sg U8712 ( .A(n3745), .B(n3746), .X(\update_mask_0/n1159 ) );
  nand_x1_sg U8713 ( .A(n7531), .B(\i_im[14][9] ), .X(n3745) );
  nand_x1_sg U8714 ( .A(n3743), .B(n3744), .X(\update_mask_0/n1160 ) );
  nand_x1_sg U8715 ( .A(n7538), .B(\i_im[14][8] ), .X(n3743) );
  nand_x1_sg U8716 ( .A(n3741), .B(n3742), .X(\update_mask_0/n1161 ) );
  nand_x1_sg U8717 ( .A(n7533), .B(\i_im[14][7] ), .X(n3741) );
  nand_x1_sg U8718 ( .A(n3739), .B(n3740), .X(\update_mask_0/n1162 ) );
  nand_x1_sg U8719 ( .A(n7528), .B(\i_im[14][6] ), .X(n3739) );
  nand_x1_sg U8720 ( .A(n3737), .B(n3738), .X(\update_mask_0/n1163 ) );
  nand_x1_sg U8721 ( .A(n7528), .B(\i_im[14][5] ), .X(n3737) );
  nand_x1_sg U8722 ( .A(n3735), .B(n3736), .X(\update_mask_0/n1164 ) );
  nand_x1_sg U8723 ( .A(n7528), .B(\i_im[14][4] ), .X(n3735) );
  nand_x1_sg U8724 ( .A(n3733), .B(n3734), .X(\update_mask_0/n1165 ) );
  nand_x1_sg U8725 ( .A(n7528), .B(\i_im[14][3] ), .X(n3733) );
  nand_x1_sg U8726 ( .A(n3731), .B(n3732), .X(\update_mask_0/n1166 ) );
  nand_x1_sg U8727 ( .A(n7528), .B(\i_im[14][2] ), .X(n3731) );
  nand_x1_sg U8728 ( .A(n3729), .B(n3730), .X(\update_mask_0/n1167 ) );
  nand_x1_sg U8729 ( .A(n7528), .B(\i_im[14][1] ), .X(n3729) );
  nand_x1_sg U8730 ( .A(n3727), .B(n3728), .X(\update_mask_0/n1168 ) );
  nand_x1_sg U8731 ( .A(n7528), .B(\i_im[14][0] ), .X(n3727) );
  nand_x1_sg U8732 ( .A(n3725), .B(n3726), .X(\update_mask_0/n1169 ) );
  nand_x1_sg U8733 ( .A(n7528), .B(\i_im[13][19] ), .X(n3725) );
  nand_x1_sg U8734 ( .A(n3723), .B(n3724), .X(\update_mask_0/n1170 ) );
  nand_x1_sg U8735 ( .A(n7528), .B(\i_im[13][18] ), .X(n3723) );
  nand_x1_sg U8736 ( .A(n3721), .B(n3722), .X(\update_mask_0/n1171 ) );
  nand_x1_sg U8737 ( .A(n7534), .B(\i_im[13][17] ), .X(n3721) );
  nand_x1_sg U8738 ( .A(n3719), .B(n3720), .X(\update_mask_0/n1172 ) );
  nand_x1_sg U8739 ( .A(n7535), .B(\i_im[13][16] ), .X(n3719) );
  nand_x1_sg U8740 ( .A(n3717), .B(n3718), .X(\update_mask_0/n1173 ) );
  nand_x1_sg U8741 ( .A(n7534), .B(\i_im[13][15] ), .X(n3717) );
  nand_x1_sg U8742 ( .A(n3715), .B(n3716), .X(\update_mask_0/n1174 ) );
  nand_x1_sg U8743 ( .A(n7535), .B(\i_im[13][14] ), .X(n3715) );
  nand_x1_sg U8744 ( .A(n3713), .B(n3714), .X(\update_mask_0/n1175 ) );
  nand_x1_sg U8745 ( .A(n7536), .B(\i_im[13][13] ), .X(n3713) );
  nand_x1_sg U8746 ( .A(n3711), .B(n3712), .X(\update_mask_0/n1176 ) );
  nand_x1_sg U8747 ( .A(n7528), .B(\i_im[13][12] ), .X(n3711) );
  nand_x1_sg U8748 ( .A(n3709), .B(n3710), .X(\update_mask_0/n1177 ) );
  nand_x1_sg U8749 ( .A(n7534), .B(\i_im[13][11] ), .X(n3709) );
  nand_x1_sg U8750 ( .A(n3707), .B(n3708), .X(\update_mask_0/n1178 ) );
  nand_x1_sg U8751 ( .A(n7535), .B(\i_im[13][10] ), .X(n3707) );
  nand_x1_sg U8752 ( .A(n3705), .B(n3706), .X(\update_mask_0/n1179 ) );
  nand_x1_sg U8753 ( .A(n7536), .B(\i_im[13][9] ), .X(n3705) );
  nand_x1_sg U8754 ( .A(n3703), .B(n3704), .X(\update_mask_0/n1180 ) );
  nand_x1_sg U8755 ( .A(n7527), .B(\i_im[13][8] ), .X(n3703) );
  nand_x1_sg U8756 ( .A(n3701), .B(n3702), .X(\update_mask_0/n1181 ) );
  nand_x1_sg U8757 ( .A(n7529), .B(\i_im[13][7] ), .X(n3701) );
  nand_x1_sg U8758 ( .A(n3699), .B(n3700), .X(\update_mask_0/n1182 ) );
  nand_x1_sg U8759 ( .A(n7533), .B(\i_im[13][6] ), .X(n3699) );
  nand_x1_sg U8760 ( .A(n3697), .B(n3698), .X(\update_mask_0/n1183 ) );
  nand_x1_sg U8761 ( .A(n7535), .B(\i_im[13][5] ), .X(n3697) );
  nand_x1_sg U8762 ( .A(n3695), .B(n3696), .X(\update_mask_0/n1184 ) );
  nand_x1_sg U8763 ( .A(n7531), .B(\i_im[13][4] ), .X(n3695) );
  nand_x1_sg U8764 ( .A(n3693), .B(n3694), .X(\update_mask_0/n1185 ) );
  nand_x1_sg U8765 ( .A(n7534), .B(\i_im[13][3] ), .X(n3693) );
  nand_x1_sg U8766 ( .A(n3691), .B(n3692), .X(\update_mask_0/n1186 ) );
  nand_x1_sg U8767 ( .A(n7535), .B(\i_im[13][2] ), .X(n3691) );
  nand_x1_sg U8768 ( .A(n3689), .B(n3690), .X(\update_mask_0/n1187 ) );
  nand_x1_sg U8769 ( .A(n7533), .B(\i_im[13][1] ), .X(n3689) );
  nand_x1_sg U8770 ( .A(n3687), .B(n3688), .X(\update_mask_0/n1188 ) );
  nand_x1_sg U8771 ( .A(n7535), .B(\i_im[13][0] ), .X(n3687) );
  nand_x1_sg U8772 ( .A(n3685), .B(n3686), .X(\update_mask_0/n1189 ) );
  nand_x1_sg U8773 ( .A(n7533), .B(\i_im[12][19] ), .X(n3685) );
  nand_x1_sg U8774 ( .A(n3683), .B(n3684), .X(\update_mask_0/n1190 ) );
  nand_x1_sg U8775 ( .A(n7533), .B(\i_im[12][18] ), .X(n3683) );
  nand_x1_sg U8776 ( .A(n3681), .B(n3682), .X(\update_mask_0/n1191 ) );
  nand_x1_sg U8777 ( .A(n7533), .B(\i_im[12][17] ), .X(n3681) );
  nand_x1_sg U8778 ( .A(n3679), .B(n3680), .X(\update_mask_0/n1192 ) );
  nand_x1_sg U8779 ( .A(n7528), .B(\i_im[12][16] ), .X(n3679) );
  nand_x1_sg U8780 ( .A(n3677), .B(n3678), .X(\update_mask_0/n1193 ) );
  nand_x1_sg U8781 ( .A(n7533), .B(\i_im[12][15] ), .X(n3677) );
  nand_x1_sg U8782 ( .A(n3675), .B(n3676), .X(\update_mask_0/n1194 ) );
  nand_x1_sg U8783 ( .A(n7535), .B(\i_im[12][14] ), .X(n3675) );
  nand_x1_sg U8784 ( .A(n3673), .B(n3674), .X(\update_mask_0/n1195 ) );
  nand_x1_sg U8785 ( .A(n7534), .B(\i_im[12][13] ), .X(n3673) );
  nand_x1_sg U8786 ( .A(n3671), .B(n3672), .X(\update_mask_0/n1196 ) );
  nand_x1_sg U8787 ( .A(n7527), .B(\i_im[12][12] ), .X(n3671) );
  nand_x1_sg U8788 ( .A(n3669), .B(n3670), .X(\update_mask_0/n1197 ) );
  nand_x1_sg U8789 ( .A(n7536), .B(\i_im[12][11] ), .X(n3669) );
  nand_x1_sg U8790 ( .A(n3667), .B(n3668), .X(\update_mask_0/n1198 ) );
  nand_x1_sg U8791 ( .A(n7528), .B(\i_im[12][10] ), .X(n3667) );
  nand_x1_sg U8792 ( .A(n3665), .B(n3666), .X(\update_mask_0/n1199 ) );
  nand_x1_sg U8793 ( .A(n7535), .B(\i_im[12][9] ), .X(n3665) );
  nand_x1_sg U8794 ( .A(n3663), .B(n3664), .X(\update_mask_0/n1200 ) );
  nand_x1_sg U8795 ( .A(n7534), .B(\i_im[12][8] ), .X(n3663) );
  nand_x1_sg U8796 ( .A(n3661), .B(n3662), .X(\update_mask_0/n1201 ) );
  nand_x1_sg U8797 ( .A(n7533), .B(\i_im[12][7] ), .X(n3661) );
  nand_x1_sg U8798 ( .A(n3659), .B(n3660), .X(\update_mask_0/n1202 ) );
  nand_x1_sg U8799 ( .A(n7528), .B(\i_im[12][6] ), .X(n3659) );
  nand_x1_sg U8800 ( .A(n3657), .B(n3658), .X(\update_mask_0/n1203 ) );
  nand_x1_sg U8801 ( .A(n7535), .B(\i_im[12][5] ), .X(n3657) );
  nand_x1_sg U8802 ( .A(n3655), .B(n3656), .X(\update_mask_0/n1204 ) );
  nand_x1_sg U8803 ( .A(n7534), .B(\i_im[12][4] ), .X(n3655) );
  nand_x1_sg U8804 ( .A(n3653), .B(n3654), .X(\update_mask_0/n1205 ) );
  nand_x1_sg U8805 ( .A(n7533), .B(\i_im[12][3] ), .X(n3653) );
  nand_x1_sg U8806 ( .A(n3651), .B(n3652), .X(\update_mask_0/n1206 ) );
  nand_x1_sg U8807 ( .A(n7528), .B(\i_im[12][2] ), .X(n3651) );
  nand_x1_sg U8808 ( .A(n3649), .B(n3650), .X(\update_mask_0/n1207 ) );
  nand_x1_sg U8809 ( .A(n7528), .B(\i_im[12][1] ), .X(n3649) );
  nand_x1_sg U8810 ( .A(n3647), .B(n3648), .X(\update_mask_0/n1208 ) );
  nand_x1_sg U8811 ( .A(n7534), .B(\i_im[12][0] ), .X(n3647) );
  nand_x1_sg U8812 ( .A(n3645), .B(n3646), .X(\update_mask_0/n1209 ) );
  nand_x1_sg U8813 ( .A(n7535), .B(\i_im[11][19] ), .X(n3645) );
  nand_x1_sg U8814 ( .A(n3643), .B(n3644), .X(\update_mask_0/n1210 ) );
  nand_x1_sg U8815 ( .A(n7533), .B(\i_im[11][18] ), .X(n3643) );
  nand_x1_sg U8816 ( .A(n3641), .B(n3642), .X(\update_mask_0/n1211 ) );
  nand_x1_sg U8817 ( .A(n7528), .B(\i_im[11][17] ), .X(n3641) );
  nand_x1_sg U8818 ( .A(n3639), .B(n3640), .X(\update_mask_0/n1212 ) );
  nand_x1_sg U8819 ( .A(n7534), .B(\i_im[11][16] ), .X(n3639) );
  nand_x1_sg U8820 ( .A(n3637), .B(n3638), .X(\update_mask_0/n1213 ) );
  nand_x1_sg U8821 ( .A(n7535), .B(\i_im[11][15] ), .X(n3637) );
  nand_x1_sg U8822 ( .A(n3635), .B(n3636), .X(\update_mask_0/n1214 ) );
  nand_x1_sg U8823 ( .A(n7536), .B(\i_im[11][14] ), .X(n3635) );
  nand_x1_sg U8824 ( .A(n3633), .B(n3634), .X(\update_mask_0/n1215 ) );
  nand_x1_sg U8825 ( .A(n7536), .B(\i_im[11][13] ), .X(n3633) );
  nand_x1_sg U8826 ( .A(n3631), .B(n3632), .X(\update_mask_0/n1216 ) );
  nand_x1_sg U8827 ( .A(n7536), .B(\i_im[11][12] ), .X(n3631) );
  nand_x1_sg U8828 ( .A(n3629), .B(n3630), .X(\update_mask_0/n1217 ) );
  nand_x1_sg U8829 ( .A(n7530), .B(\i_im[11][11] ), .X(n3629) );
  nand_x1_sg U8830 ( .A(n3627), .B(n3628), .X(\update_mask_0/n1218 ) );
  nand_x1_sg U8831 ( .A(n7536), .B(\i_im[11][10] ), .X(n3627) );
  nand_x1_sg U8832 ( .A(n3625), .B(n3626), .X(\update_mask_0/n1219 ) );
  nand_x1_sg U8833 ( .A(n7527), .B(\i_im[11][9] ), .X(n3625) );
  nand_x1_sg U8834 ( .A(n3623), .B(n3624), .X(\update_mask_0/n1220 ) );
  nand_x1_sg U8835 ( .A(n7536), .B(\i_im[11][8] ), .X(n3623) );
  nand_x1_sg U8836 ( .A(n3621), .B(n3622), .X(\update_mask_0/n1221 ) );
  nand_x1_sg U8837 ( .A(n7535), .B(\i_im[11][7] ), .X(n3621) );
  nand_x1_sg U8838 ( .A(n3619), .B(n3620), .X(\update_mask_0/n1222 ) );
  nand_x1_sg U8839 ( .A(n7536), .B(\i_im[11][6] ), .X(n3619) );
  nand_x1_sg U8840 ( .A(n3617), .B(n3618), .X(\update_mask_0/n1223 ) );
  nand_x1_sg U8841 ( .A(n7528), .B(\i_im[11][5] ), .X(n3617) );
  nand_x1_sg U8842 ( .A(n3615), .B(n3616), .X(\update_mask_0/n1224 ) );
  nand_x1_sg U8843 ( .A(n7527), .B(\i_im[11][4] ), .X(n3615) );
  nand_x1_sg U8844 ( .A(n3613), .B(n3614), .X(\update_mask_0/n1225 ) );
  nand_x1_sg U8845 ( .A(n7527), .B(\i_im[11][3] ), .X(n3613) );
  nand_x1_sg U8846 ( .A(n3611), .B(n3612), .X(\update_mask_0/n1226 ) );
  nand_x1_sg U8847 ( .A(n7527), .B(\i_im[11][2] ), .X(n3611) );
  nand_x1_sg U8848 ( .A(n3609), .B(n3610), .X(\update_mask_0/n1227 ) );
  nand_x1_sg U8849 ( .A(n7527), .B(\i_im[11][1] ), .X(n3609) );
  nand_x1_sg U8850 ( .A(n3607), .B(n3608), .X(\update_mask_0/n1228 ) );
  nand_x1_sg U8851 ( .A(n7527), .B(\i_im[11][0] ), .X(n3607) );
  nand_x1_sg U8852 ( .A(n3605), .B(n3606), .X(\update_mask_0/n1229 ) );
  nand_x1_sg U8853 ( .A(n7527), .B(\i_im[10][19] ), .X(n3605) );
  nand_x1_sg U8854 ( .A(n3603), .B(n3604), .X(\update_mask_0/n1230 ) );
  nand_x1_sg U8855 ( .A(n7527), .B(\i_im[10][18] ), .X(n3603) );
  nand_x1_sg U8856 ( .A(n3601), .B(n3602), .X(\update_mask_0/n1231 ) );
  nand_x1_sg U8857 ( .A(n7527), .B(\i_im[10][17] ), .X(n3601) );
  nand_x1_sg U8858 ( .A(n3599), .B(n3600), .X(\update_mask_0/n1232 ) );
  nand_x1_sg U8859 ( .A(n7527), .B(\i_im[10][16] ), .X(n3599) );
  nand_x1_sg U8860 ( .A(n3597), .B(n3598), .X(\update_mask_0/n1233 ) );
  nand_x1_sg U8861 ( .A(n7533), .B(\i_im[10][15] ), .X(n3597) );
  nand_x1_sg U8862 ( .A(n3595), .B(n3596), .X(\update_mask_0/n1234 ) );
  nand_x1_sg U8863 ( .A(n7536), .B(\i_im[10][14] ), .X(n3595) );
  nand_x1_sg U8864 ( .A(n3593), .B(n3594), .X(\update_mask_0/n1235 ) );
  nand_x1_sg U8865 ( .A(n7530), .B(\i_im[10][13] ), .X(n3593) );
  nand_x1_sg U8866 ( .A(n3591), .B(n3592), .X(\update_mask_0/n1236 ) );
  nand_x1_sg U8867 ( .A(n7533), .B(\i_im[10][12] ), .X(n3591) );
  nand_x1_sg U8868 ( .A(n3589), .B(n3590), .X(\update_mask_0/n1237 ) );
  nand_x1_sg U8869 ( .A(n7536), .B(\i_im[10][11] ), .X(n3589) );
  nand_x1_sg U8870 ( .A(n3587), .B(n3588), .X(\update_mask_0/n1238 ) );
  nand_x1_sg U8871 ( .A(n7531), .B(\i_im[10][10] ), .X(n3587) );
  nand_x1_sg U8872 ( .A(n3585), .B(n3586), .X(\update_mask_0/n1239 ) );
  nand_x1_sg U8873 ( .A(n7534), .B(\i_im[10][9] ), .X(n3585) );
  nand_x1_sg U8874 ( .A(n3583), .B(n3584), .X(\update_mask_0/n1240 ) );
  nand_x1_sg U8875 ( .A(n7533), .B(\i_im[10][8] ), .X(n3583) );
  nand_x1_sg U8876 ( .A(n3581), .B(n3582), .X(\update_mask_0/n1241 ) );
  nand_x1_sg U8877 ( .A(n7527), .B(\i_im[10][7] ), .X(n3581) );
  nand_x1_sg U8878 ( .A(n3579), .B(n3580), .X(\update_mask_0/n1242 ) );
  nand_x1_sg U8879 ( .A(n7531), .B(\i_im[10][6] ), .X(n3579) );
  nand_x1_sg U8880 ( .A(n3577), .B(n3578), .X(\update_mask_0/n1243 ) );
  nand_x1_sg U8881 ( .A(n7527), .B(\i_im[10][5] ), .X(n3577) );
  nand_x1_sg U8882 ( .A(n3575), .B(n3576), .X(\update_mask_0/n1244 ) );
  nand_x1_sg U8883 ( .A(n7530), .B(\i_im[10][4] ), .X(n3575) );
  nand_x1_sg U8884 ( .A(n3573), .B(n3574), .X(\update_mask_0/n1245 ) );
  nand_x1_sg U8885 ( .A(n7534), .B(\i_im[10][3] ), .X(n3573) );
  nand_x1_sg U8886 ( .A(n3571), .B(n3572), .X(\update_mask_0/n1246 ) );
  nand_x1_sg U8887 ( .A(n7527), .B(\i_im[10][2] ), .X(n3571) );
  nand_x1_sg U8888 ( .A(n3569), .B(n3570), .X(\update_mask_0/n1247 ) );
  nand_x1_sg U8889 ( .A(n7533), .B(\i_im[10][1] ), .X(n3569) );
  nand_x1_sg U8890 ( .A(n3567), .B(n3568), .X(\update_mask_0/n1248 ) );
  nand_x1_sg U8891 ( .A(n7528), .B(\i_im[10][0] ), .X(n3567) );
  nand_x1_sg U8892 ( .A(n3565), .B(n3566), .X(\update_mask_0/n1249 ) );
  nand_x1_sg U8893 ( .A(n7530), .B(\i_im[9][19] ), .X(n3565) );
  nand_x1_sg U8894 ( .A(n3563), .B(n3564), .X(\update_mask_0/n1250 ) );
  nand_x1_sg U8895 ( .A(n7527), .B(\i_im[9][18] ), .X(n3563) );
  nand_x1_sg U8896 ( .A(n3561), .B(n3562), .X(\update_mask_0/n1251 ) );
  nand_x1_sg U8897 ( .A(n7530), .B(\i_im[9][17] ), .X(n3561) );
  nand_x1_sg U8898 ( .A(n3559), .B(n3560), .X(\update_mask_0/n1252 ) );
  nand_x1_sg U8899 ( .A(n7531), .B(\i_im[9][16] ), .X(n3559) );
  nand_x1_sg U8900 ( .A(n3557), .B(n3558), .X(\update_mask_0/n1253 ) );
  nand_x1_sg U8901 ( .A(n7530), .B(\i_im[9][15] ), .X(n3557) );
  nand_x1_sg U8902 ( .A(n3555), .B(n3556), .X(\update_mask_0/n1254 ) );
  nand_x1_sg U8903 ( .A(n7527), .B(\i_im[9][14] ), .X(n3555) );
  nand_x1_sg U8904 ( .A(n3553), .B(n3554), .X(\update_mask_0/n1255 ) );
  nand_x1_sg U8905 ( .A(n7535), .B(\i_im[9][13] ), .X(n3553) );
  nand_x1_sg U8906 ( .A(n3551), .B(n3552), .X(\update_mask_0/n1256 ) );
  nand_x1_sg U8907 ( .A(n7527), .B(\i_im[9][12] ), .X(n3551) );
  nand_x1_sg U8908 ( .A(n3549), .B(n3550), .X(\update_mask_0/n1257 ) );
  nand_x1_sg U8909 ( .A(n7528), .B(\i_im[9][11] ), .X(n3549) );
  nand_x1_sg U8910 ( .A(n3547), .B(n3548), .X(\update_mask_0/n1258 ) );
  nand_x1_sg U8911 ( .A(n7535), .B(\i_im[9][10] ), .X(n3547) );
  nand_x1_sg U8912 ( .A(n3545), .B(n3546), .X(\update_mask_0/n1259 ) );
  nand_x1_sg U8913 ( .A(n7528), .B(\i_im[9][9] ), .X(n3545) );
  nand_x1_sg U8914 ( .A(n3543), .B(n3544), .X(\update_mask_0/n1260 ) );
  nand_x1_sg U8915 ( .A(n7535), .B(\i_im[9][8] ), .X(n3543) );
  nand_x1_sg U8916 ( .A(n3541), .B(n3542), .X(\update_mask_0/n1261 ) );
  nand_x1_sg U8917 ( .A(n7527), .B(\i_im[9][7] ), .X(n3541) );
  nand_x1_sg U8918 ( .A(n3539), .B(n3540), .X(\update_mask_0/n1262 ) );
  nand_x1_sg U8919 ( .A(n7528), .B(\i_im[9][6] ), .X(n3539) );
  nand_x1_sg U8920 ( .A(n3537), .B(n3538), .X(\update_mask_0/n1263 ) );
  nand_x1_sg U8921 ( .A(n7531), .B(\i_im[9][5] ), .X(n3537) );
  nand_x1_sg U8922 ( .A(n3535), .B(n3536), .X(\update_mask_0/n1264 ) );
  nand_x1_sg U8923 ( .A(n7531), .B(\i_im[9][4] ), .X(n3535) );
  nand_x1_sg U8924 ( .A(n3533), .B(n3534), .X(\update_mask_0/n1265 ) );
  nand_x1_sg U8925 ( .A(n7527), .B(\i_im[9][3] ), .X(n3533) );
  nand_x1_sg U8926 ( .A(n3531), .B(n3532), .X(\update_mask_0/n1266 ) );
  nand_x1_sg U8927 ( .A(n7534), .B(\i_im[9][2] ), .X(n3531) );
  nand_x1_sg U8928 ( .A(n3529), .B(n3530), .X(\update_mask_0/n1267 ) );
  nand_x1_sg U8929 ( .A(n7534), .B(\i_im[9][1] ), .X(n3529) );
  nand_x1_sg U8930 ( .A(n3527), .B(n3528), .X(\update_mask_0/n1268 ) );
  nand_x1_sg U8931 ( .A(n7535), .B(\i_im[9][0] ), .X(n3527) );
  nand_x1_sg U8932 ( .A(n3525), .B(n3526), .X(\update_mask_0/n1269 ) );
  nand_x1_sg U8933 ( .A(n7529), .B(\i_im[8][19] ), .X(n3525) );
  nand_x1_sg U8934 ( .A(n3523), .B(n3524), .X(\update_mask_0/n1270 ) );
  nand_x1_sg U8935 ( .A(n7529), .B(\i_im[8][18] ), .X(n3523) );
  nand_x1_sg U8936 ( .A(n3521), .B(n3522), .X(\update_mask_0/n1271 ) );
  nand_x1_sg U8937 ( .A(n7530), .B(\i_im[8][17] ), .X(n3521) );
  nand_x1_sg U8938 ( .A(n3519), .B(n3520), .X(\update_mask_0/n1272 ) );
  nand_x1_sg U8939 ( .A(n7527), .B(\i_im[8][16] ), .X(n3519) );
  nand_x1_sg U8940 ( .A(n3517), .B(n3518), .X(\update_mask_0/n1273 ) );
  nand_x1_sg U8941 ( .A(n7534), .B(\i_im[8][15] ), .X(n3517) );
  nand_x1_sg U8942 ( .A(n3515), .B(n3516), .X(\update_mask_0/n1274 ) );
  nand_x1_sg U8943 ( .A(n7531), .B(\i_im[8][14] ), .X(n3515) );
  nand_x1_sg U8944 ( .A(n3513), .B(n3514), .X(\update_mask_0/n1275 ) );
  nand_x1_sg U8945 ( .A(n7536), .B(\i_im[8][13] ), .X(n3513) );
  nand_x1_sg U8946 ( .A(n3511), .B(n3512), .X(\update_mask_0/n1276 ) );
  nand_x1_sg U8947 ( .A(n7528), .B(\i_im[8][12] ), .X(n3511) );
  nand_x1_sg U8948 ( .A(n3509), .B(n3510), .X(\update_mask_0/n1277 ) );
  nand_x1_sg U8949 ( .A(n7536), .B(\i_im[8][11] ), .X(n3509) );
  nand_x1_sg U8950 ( .A(n3507), .B(n3508), .X(\update_mask_0/n1278 ) );
  nand_x1_sg U8951 ( .A(n7535), .B(\i_im[8][10] ), .X(n3507) );
  nand_x1_sg U8952 ( .A(n3505), .B(n3506), .X(\update_mask_0/n1279 ) );
  nand_x1_sg U8953 ( .A(n7536), .B(\i_im[8][9] ), .X(n3505) );
  nand_x1_sg U8954 ( .A(n3503), .B(n3504), .X(\update_mask_0/n1280 ) );
  nand_x1_sg U8955 ( .A(n7534), .B(\i_im[8][8] ), .X(n3503) );
  nand_x1_sg U8956 ( .A(n3501), .B(n3502), .X(\update_mask_0/n1281 ) );
  nand_x1_sg U8957 ( .A(n7535), .B(\i_im[8][7] ), .X(n3501) );
  nand_x1_sg U8958 ( .A(n3499), .B(n3500), .X(\update_mask_0/n1282 ) );
  nand_x1_sg U8959 ( .A(n7527), .B(\i_im[8][6] ), .X(n3499) );
  nand_x1_sg U8960 ( .A(n3497), .B(n3498), .X(\update_mask_0/n1283 ) );
  nand_x1_sg U8961 ( .A(n7533), .B(\i_im[8][5] ), .X(n3497) );
  nand_x1_sg U8962 ( .A(n3495), .B(n3496), .X(\update_mask_0/n1284 ) );
  nand_x1_sg U8963 ( .A(n7534), .B(\i_im[8][4] ), .X(n3495) );
  nand_x1_sg U8964 ( .A(n3493), .B(n3494), .X(\update_mask_0/n1285 ) );
  nand_x1_sg U8965 ( .A(n7531), .B(\i_im[8][3] ), .X(n3493) );
  nand_x1_sg U8966 ( .A(n3491), .B(n3492), .X(\update_mask_0/n1286 ) );
  nand_x1_sg U8967 ( .A(n7536), .B(\i_im[8][2] ), .X(n3491) );
  nand_x1_sg U8968 ( .A(n3489), .B(n3490), .X(\update_mask_0/n1287 ) );
  nand_x1_sg U8969 ( .A(n7533), .B(\i_im[8][1] ), .X(n3489) );
  nand_x1_sg U8970 ( .A(n3487), .B(n3488), .X(\update_mask_0/n1288 ) );
  nand_x1_sg U8971 ( .A(n7536), .B(\i_im[8][0] ), .X(n3487) );
  nand_x1_sg U8972 ( .A(n3485), .B(n3486), .X(\update_mask_0/n1289 ) );
  nand_x1_sg U8973 ( .A(n7530), .B(\i_im[7][19] ), .X(n3485) );
  nand_x1_sg U8974 ( .A(n3483), .B(n3484), .X(\update_mask_0/n1290 ) );
  nand_x1_sg U8975 ( .A(n7533), .B(\i_im[7][18] ), .X(n3483) );
  nand_x1_sg U8976 ( .A(n3481), .B(n3482), .X(\update_mask_0/n1291 ) );
  nand_x1_sg U8977 ( .A(n7533), .B(\i_im[7][17] ), .X(n3481) );
  nand_x1_sg U8978 ( .A(n3479), .B(n3480), .X(\update_mask_0/n1292 ) );
  nand_x1_sg U8979 ( .A(n7527), .B(\i_im[7][16] ), .X(n3479) );
  nand_x1_sg U8980 ( .A(n3477), .B(n3478), .X(\update_mask_0/n1293 ) );
  nand_x1_sg U8981 ( .A(n7533), .B(\i_im[7][15] ), .X(n3477) );
  nand_x1_sg U8982 ( .A(n3475), .B(n3476), .X(\update_mask_0/n1294 ) );
  nand_x1_sg U8983 ( .A(n7533), .B(\i_im[7][14] ), .X(n3475) );
  nand_x1_sg U8984 ( .A(n3473), .B(n3474), .X(\update_mask_0/n1295 ) );
  nand_x1_sg U8985 ( .A(n7528), .B(\i_im[7][13] ), .X(n3473) );
  nand_x1_sg U8986 ( .A(n3471), .B(n3472), .X(\update_mask_0/n1296 ) );
  nand_x1_sg U8987 ( .A(n7533), .B(\i_im[7][12] ), .X(n3471) );
  nand_x1_sg U8988 ( .A(n3469), .B(n3470), .X(\update_mask_0/n1297 ) );
  nand_x1_sg U8989 ( .A(n7528), .B(\i_im[7][11] ), .X(n3469) );
  nand_x1_sg U8990 ( .A(n3467), .B(n3468), .X(\update_mask_0/n1298 ) );
  nand_x1_sg U8991 ( .A(n7535), .B(\i_im[7][10] ), .X(n3467) );
  nand_x1_sg U8992 ( .A(n3465), .B(n3466), .X(\update_mask_0/n1299 ) );
  nand_x1_sg U8993 ( .A(n7528), .B(\i_im[7][9] ), .X(n3465) );
  nand_x1_sg U8994 ( .A(n3463), .B(n3464), .X(\update_mask_0/n1300 ) );
  nand_x1_sg U8995 ( .A(n7535), .B(\i_im[7][8] ), .X(n3463) );
  nand_x1_sg U8996 ( .A(n3461), .B(n3462), .X(\update_mask_0/n1301 ) );
  nand_x1_sg U8997 ( .A(n7533), .B(\i_im[7][7] ), .X(n3461) );
  nand_x1_sg U8998 ( .A(n3459), .B(n3460), .X(\update_mask_0/n1302 ) );
  nand_x1_sg U8999 ( .A(n7529), .B(\i_im[7][6] ), .X(n3459) );
  nand_x1_sg U9000 ( .A(n3457), .B(n3458), .X(\update_mask_0/n1303 ) );
  nand_x1_sg U9001 ( .A(n7528), .B(\i_im[7][5] ), .X(n3457) );
  nand_x1_sg U9002 ( .A(n3455), .B(n3456), .X(\update_mask_0/n1304 ) );
  nand_x1_sg U9003 ( .A(n7529), .B(\i_im[7][4] ), .X(n3455) );
  nand_x1_sg U9004 ( .A(n3453), .B(n3454), .X(\update_mask_0/n1305 ) );
  nand_x1_sg U9005 ( .A(n7531), .B(\i_im[7][3] ), .X(n3453) );
  nand_x1_sg U9006 ( .A(n3451), .B(n3452), .X(\update_mask_0/n1306 ) );
  nand_x1_sg U9007 ( .A(n7536), .B(\i_im[7][2] ), .X(n3451) );
  nand_x1_sg U9008 ( .A(n3449), .B(n3450), .X(\update_mask_0/n1307 ) );
  nand_x1_sg U9009 ( .A(n7531), .B(\i_im[7][1] ), .X(n3449) );
  nand_x1_sg U9010 ( .A(n3447), .B(n3448), .X(\update_mask_0/n1308 ) );
  nand_x1_sg U9011 ( .A(n7533), .B(\i_im[7][0] ), .X(n3447) );
  nand_x1_sg U9012 ( .A(n3445), .B(n3446), .X(\update_mask_0/n1309 ) );
  nand_x1_sg U9013 ( .A(n7533), .B(\i_im[6][19] ), .X(n3445) );
  nand_x1_sg U9014 ( .A(n3443), .B(n3444), .X(\update_mask_0/n1310 ) );
  nand_x1_sg U9015 ( .A(n7533), .B(\i_im[6][18] ), .X(n3443) );
  nand_x1_sg U9016 ( .A(n3441), .B(n3442), .X(\update_mask_0/n1311 ) );
  nand_x1_sg U9017 ( .A(n7536), .B(\i_im[6][17] ), .X(n3441) );
  nand_x1_sg U9018 ( .A(n3439), .B(n3440), .X(\update_mask_0/n1312 ) );
  nand_x1_sg U9019 ( .A(n7533), .B(\i_im[6][16] ), .X(n3439) );
  nand_x1_sg U9020 ( .A(n3437), .B(n3438), .X(\update_mask_0/n1313 ) );
  nand_x1_sg U9021 ( .A(n7536), .B(\i_im[6][15] ), .X(n3437) );
  nand_x1_sg U9022 ( .A(n3435), .B(n3436), .X(\update_mask_0/n1314 ) );
  nand_x1_sg U9023 ( .A(n7534), .B(\i_im[6][14] ), .X(n3435) );
  nand_x1_sg U9024 ( .A(n3433), .B(n3434), .X(\update_mask_0/n1315 ) );
  nand_x1_sg U9025 ( .A(n7529), .B(\i_im[6][13] ), .X(n3433) );
  nand_x1_sg U9026 ( .A(n3431), .B(n3432), .X(\update_mask_0/n1316 ) );
  nand_x1_sg U9027 ( .A(n7531), .B(\i_im[6][12] ), .X(n3431) );
  nand_x1_sg U9028 ( .A(n3429), .B(n3430), .X(\update_mask_0/n1317 ) );
  nand_x1_sg U9029 ( .A(n7530), .B(\i_im[6][11] ), .X(n3429) );
  nand_x1_sg U9030 ( .A(n3427), .B(n3428), .X(\update_mask_0/n1318 ) );
  nand_x1_sg U9031 ( .A(n7529), .B(\i_im[6][10] ), .X(n3427) );
  nand_x1_sg U9032 ( .A(n3425), .B(n3426), .X(\update_mask_0/n1319 ) );
  nand_x1_sg U9033 ( .A(n7531), .B(\i_im[6][9] ), .X(n3425) );
  nand_x1_sg U9034 ( .A(n3423), .B(n3424), .X(\update_mask_0/n1320 ) );
  nand_x1_sg U9035 ( .A(n7530), .B(\i_im[6][8] ), .X(n3423) );
  nand_x1_sg U9036 ( .A(n3421), .B(n3422), .X(\update_mask_0/n1321 ) );
  nand_x1_sg U9037 ( .A(n7529), .B(\i_im[6][7] ), .X(n3421) );
  nand_x1_sg U9038 ( .A(n3419), .B(n3420), .X(\update_mask_0/n1322 ) );
  nand_x1_sg U9039 ( .A(n7529), .B(\i_im[6][6] ), .X(n3419) );
  nand_x1_sg U9040 ( .A(n3417), .B(n3418), .X(\update_mask_0/n1323 ) );
  nand_x1_sg U9041 ( .A(n7531), .B(\i_im[6][5] ), .X(n3417) );
  nand_x1_sg U9042 ( .A(n3415), .B(n3416), .X(\update_mask_0/n1324 ) );
  nand_x1_sg U9043 ( .A(n7536), .B(\i_im[6][4] ), .X(n3415) );
  nand_x1_sg U9044 ( .A(n3413), .B(n3414), .X(\update_mask_0/n1325 ) );
  nand_x1_sg U9045 ( .A(n7536), .B(\i_im[6][3] ), .X(n3413) );
  nand_x1_sg U9046 ( .A(n3411), .B(n3412), .X(\update_mask_0/n1326 ) );
  nand_x1_sg U9047 ( .A(n7536), .B(\i_im[6][2] ), .X(n3411) );
  nand_x1_sg U9048 ( .A(n3409), .B(n3410), .X(\update_mask_0/n1327 ) );
  nand_x1_sg U9049 ( .A(n7536), .B(\i_im[6][1] ), .X(n3409) );
  nand_x1_sg U9050 ( .A(n3407), .B(n3408), .X(\update_mask_0/n1328 ) );
  nand_x1_sg U9051 ( .A(n7536), .B(\i_im[6][0] ), .X(n3407) );
  nand_x1_sg U9052 ( .A(n3405), .B(n3406), .X(\update_mask_0/n1329 ) );
  nand_x1_sg U9053 ( .A(n7536), .B(\i_im[5][19] ), .X(n3405) );
  nand_x1_sg U9054 ( .A(n3403), .B(n3404), .X(\update_mask_0/n1330 ) );
  nand_x1_sg U9055 ( .A(n7536), .B(\i_im[5][18] ), .X(n3403) );
  nand_x1_sg U9056 ( .A(n3401), .B(n3402), .X(\update_mask_0/n1331 ) );
  nand_x1_sg U9057 ( .A(n7536), .B(\i_im[5][17] ), .X(n3401) );
  nand_x1_sg U9058 ( .A(n3399), .B(n3400), .X(\update_mask_0/n1332 ) );
  nand_x1_sg U9059 ( .A(n7536), .B(\i_im[5][16] ), .X(n3399) );
  inv_x1_sg U9060 ( .A(n9032), .X(n7046) );
  nand_x1_sg U9061 ( .A(n3397), .B(n3398), .X(\update_mask_0/n1333 ) );
  nand_x1_sg U9062 ( .A(n7536), .B(\i_im[5][15] ), .X(n3397) );
  nand_x1_sg U9063 ( .A(n3395), .B(n3396), .X(\update_mask_0/n1334 ) );
  nand_x1_sg U9064 ( .A(n7536), .B(\i_im[5][14] ), .X(n3395) );
  nand_x1_sg U9065 ( .A(n3393), .B(n3394), .X(\update_mask_0/n1335 ) );
  nand_x1_sg U9066 ( .A(n7534), .B(\i_im[5][13] ), .X(n3393) );
  nand_x1_sg U9067 ( .A(n3391), .B(n3392), .X(\update_mask_0/n1336 ) );
  nand_x1_sg U9068 ( .A(n7535), .B(\i_im[5][12] ), .X(n3391) );
  nand_x1_sg U9069 ( .A(n3389), .B(n3390), .X(\update_mask_0/n1337 ) );
  nand_x1_sg U9070 ( .A(n7536), .B(\i_im[5][11] ), .X(n3389) );
  nand_x1_sg U9071 ( .A(n3387), .B(n3388), .X(\update_mask_0/n1338 ) );
  nand_x1_sg U9072 ( .A(n7534), .B(\i_im[5][10] ), .X(n3387) );
  nand_x1_sg U9073 ( .A(n3385), .B(n3386), .X(\update_mask_0/n1339 ) );
  nand_x1_sg U9074 ( .A(n7535), .B(\i_im[5][9] ), .X(n3385) );
  nand_x1_sg U9075 ( .A(n3383), .B(n3384), .X(\update_mask_0/n1340 ) );
  nand_x1_sg U9076 ( .A(n7536), .B(\i_im[5][8] ), .X(n3383) );
  nand_x1_sg U9077 ( .A(n3381), .B(n3382), .X(\update_mask_0/n1341 ) );
  nand_x1_sg U9078 ( .A(n7534), .B(\i_im[5][7] ), .X(n3381) );
  nand_x1_sg U9079 ( .A(n3379), .B(n3380), .X(\update_mask_0/n1342 ) );
  nand_x1_sg U9080 ( .A(n7535), .B(\i_im[5][6] ), .X(n3379) );
  nand_x1_sg U9081 ( .A(n3377), .B(n3378), .X(\update_mask_0/n1343 ) );
  nand_x1_sg U9082 ( .A(n7533), .B(\i_im[5][5] ), .X(n3377) );
  nand_x1_sg U9083 ( .A(n3375), .B(n3376), .X(\update_mask_0/n1344 ) );
  nand_x1_sg U9084 ( .A(n7528), .B(\i_im[5][4] ), .X(n3375) );
  nand_x1_sg U9085 ( .A(n3373), .B(n3374), .X(\update_mask_0/n1345 ) );
  nand_x1_sg U9086 ( .A(n7536), .B(\i_im[5][3] ), .X(n3373) );
  nand_x1_sg U9087 ( .A(n3371), .B(n3372), .X(\update_mask_0/n1346 ) );
  nand_x1_sg U9088 ( .A(n7535), .B(\i_im[5][2] ), .X(n3371) );
  nand_x1_sg U9089 ( .A(n3369), .B(n3370), .X(\update_mask_0/n1347 ) );
  nand_x1_sg U9090 ( .A(n7534), .B(\i_im[5][1] ), .X(n3369) );
  nand_x1_sg U9091 ( .A(n3367), .B(n3368), .X(\update_mask_0/n1348 ) );
  nand_x1_sg U9092 ( .A(n7528), .B(\i_im[5][0] ), .X(n3367) );
  nand_x1_sg U9093 ( .A(n3365), .B(n3366), .X(\update_mask_0/n1349 ) );
  nand_x1_sg U9094 ( .A(n7536), .B(\i_im[4][19] ), .X(n3365) );
  nand_x1_sg U9095 ( .A(n3363), .B(n3364), .X(\update_mask_0/n1350 ) );
  nand_x1_sg U9096 ( .A(n7529), .B(\i_im[4][18] ), .X(n3363) );
  nand_x1_sg U9097 ( .A(n3361), .B(n3362), .X(\update_mask_0/n1351 ) );
  nand_x1_sg U9098 ( .A(n7536), .B(\i_im[4][17] ), .X(n3361) );
  nand_x1_sg U9099 ( .A(n3359), .B(n3360), .X(\update_mask_0/n1352 ) );
  nand_x1_sg U9100 ( .A(n7534), .B(\i_im[4][16] ), .X(n3359) );
  inv_x1_sg U9101 ( .A(n9036), .X(n7045) );
  nand_x1_sg U9102 ( .A(n3357), .B(n3358), .X(\update_mask_0/n1353 ) );
  nand_x1_sg U9103 ( .A(n7535), .B(\i_im[4][15] ), .X(n3357) );
  nand_x1_sg U9104 ( .A(n3355), .B(n3356), .X(\update_mask_0/n1354 ) );
  nand_x1_sg U9105 ( .A(n7527), .B(\i_im[4][14] ), .X(n3355) );
  nand_x1_sg U9106 ( .A(n3353), .B(n3354), .X(\update_mask_0/n1355 ) );
  nand_x1_sg U9107 ( .A(n7533), .B(\i_im[4][13] ), .X(n3353) );
  nand_x1_sg U9108 ( .A(n3351), .B(n3352), .X(\update_mask_0/n1356 ) );
  nand_x1_sg U9109 ( .A(n7529), .B(\i_im[4][12] ), .X(n3351) );
  nand_x1_sg U9110 ( .A(n3349), .B(n3350), .X(\update_mask_0/n1357 ) );
  nand_x1_sg U9111 ( .A(n7536), .B(\i_im[4][11] ), .X(n3349) );
  nand_x1_sg U9112 ( .A(n3347), .B(n3348), .X(\update_mask_0/n1358 ) );
  nand_x1_sg U9113 ( .A(n7536), .B(\i_im[4][10] ), .X(n3347) );
  nand_x1_sg U9114 ( .A(n3345), .B(n3346), .X(\update_mask_0/n1359 ) );
  nand_x1_sg U9115 ( .A(n7536), .B(\i_im[4][9] ), .X(n3345) );
  nand_x1_sg U9116 ( .A(n3343), .B(n3344), .X(\update_mask_0/n1360 ) );
  nand_x1_sg U9117 ( .A(n7536), .B(\i_im[4][8] ), .X(n3343) );
  nand_x1_sg U9118 ( .A(n3341), .B(n3342), .X(\update_mask_0/n1361 ) );
  nand_x1_sg U9119 ( .A(n7533), .B(\i_im[4][7] ), .X(n3341) );
  nand_x1_sg U9120 ( .A(n3339), .B(n3340), .X(\update_mask_0/n1362 ) );
  nand_x1_sg U9121 ( .A(n7536), .B(\i_im[4][6] ), .X(n3339) );
  nand_x1_sg U9122 ( .A(n3337), .B(n3338), .X(\update_mask_0/n1363 ) );
  nand_x1_sg U9123 ( .A(n7536), .B(\i_im[4][5] ), .X(n3337) );
  nand_x1_sg U9124 ( .A(n3335), .B(n3336), .X(\update_mask_0/n1364 ) );
  nand_x1_sg U9125 ( .A(n7533), .B(\i_im[4][4] ), .X(n3335) );
  nand_x1_sg U9126 ( .A(n3333), .B(n3334), .X(\update_mask_0/n1365 ) );
  nand_x1_sg U9127 ( .A(n7536), .B(\i_im[4][3] ), .X(n3333) );
  nand_x1_sg U9128 ( .A(n3331), .B(n3332), .X(\update_mask_0/n1366 ) );
  nand_x1_sg U9129 ( .A(n7534), .B(\i_im[4][2] ), .X(n3331) );
  nand_x1_sg U9130 ( .A(n3329), .B(n3330), .X(\update_mask_0/n1367 ) );
  nand_x1_sg U9131 ( .A(n7536), .B(\i_im[4][1] ), .X(n3329) );
  nand_x1_sg U9132 ( .A(n3327), .B(n3328), .X(\update_mask_0/n1368 ) );
  nand_x1_sg U9133 ( .A(n7531), .B(\i_im[4][0] ), .X(n3327) );
  nand_x1_sg U9134 ( .A(n3325), .B(n3326), .X(\update_mask_0/n1369 ) );
  nand_x1_sg U9135 ( .A(n7530), .B(\i_im[3][19] ), .X(n3325) );
  nand_x1_sg U9136 ( .A(n3323), .B(n3324), .X(\update_mask_0/n1370 ) );
  nand_x1_sg U9137 ( .A(n7527), .B(\i_im[3][18] ), .X(n3323) );
  nand_x1_sg U9138 ( .A(n3321), .B(n3322), .X(\update_mask_0/n1371 ) );
  nand_x1_sg U9139 ( .A(n7534), .B(\i_im[3][17] ), .X(n3321) );
  nand_x1_sg U9140 ( .A(n3319), .B(n3320), .X(\update_mask_0/n1372 ) );
  nand_x1_sg U9141 ( .A(n7534), .B(\i_im[3][16] ), .X(n3319) );
  inv_x1_sg U9142 ( .A(n9040), .X(n7044) );
  nand_x1_sg U9143 ( .A(n3317), .B(n3318), .X(\update_mask_0/n1373 ) );
  nand_x1_sg U9144 ( .A(n7528), .B(\i_im[3][15] ), .X(n3317) );
  nand_x1_sg U9145 ( .A(n3315), .B(n3316), .X(\update_mask_0/n1374 ) );
  nand_x1_sg U9146 ( .A(n7531), .B(\i_im[3][14] ), .X(n3315) );
  nand_x1_sg U9147 ( .A(n3313), .B(n3314), .X(\update_mask_0/n1375 ) );
  nand_x1_sg U9148 ( .A(n7527), .B(\i_im[3][13] ), .X(n3313) );
  nand_x1_sg U9149 ( .A(n3311), .B(n3312), .X(\update_mask_0/n1376 ) );
  nand_x1_sg U9150 ( .A(n7533), .B(\i_im[3][12] ), .X(n3311) );
  nand_x1_sg U9151 ( .A(n3309), .B(n3310), .X(\update_mask_0/n1377 ) );
  nand_x1_sg U9152 ( .A(n7527), .B(\i_im[3][11] ), .X(n3309) );
  nand_x1_sg U9153 ( .A(n3307), .B(n3308), .X(\update_mask_0/n1378 ) );
  nand_x1_sg U9154 ( .A(n7530), .B(\i_im[3][10] ), .X(n3307) );
  nand_x1_sg U9155 ( .A(n3305), .B(n3306), .X(\update_mask_0/n1379 ) );
  nand_x1_sg U9156 ( .A(n7527), .B(\i_im[3][9] ), .X(n3305) );
  nand_x1_sg U9157 ( .A(n3303), .B(n3304), .X(\update_mask_0/n1380 ) );
  nand_x1_sg U9158 ( .A(n7528), .B(\i_im[3][8] ), .X(n3303) );
  nand_x1_sg U9159 ( .A(n3301), .B(n3302), .X(\update_mask_0/n1381 ) );
  nand_x1_sg U9160 ( .A(n7535), .B(\i_im[3][7] ), .X(n3301) );
  nand_x1_sg U9161 ( .A(n3299), .B(n3300), .X(\update_mask_0/n1382 ) );
  nand_x1_sg U9162 ( .A(n7527), .B(\i_im[3][6] ), .X(n3299) );
  nand_x1_sg U9163 ( .A(n3297), .B(n3298), .X(\update_mask_0/n1383 ) );
  nand_x1_sg U9164 ( .A(n7529), .B(\i_im[3][5] ), .X(n3297) );
  nand_x1_sg U9165 ( .A(n3295), .B(n3296), .X(\update_mask_0/n1384 ) );
  nand_x1_sg U9166 ( .A(n7528), .B(\i_im[3][4] ), .X(n3295) );
  nand_x1_sg U9167 ( .A(n3293), .B(n3294), .X(\update_mask_0/n1385 ) );
  nand_x1_sg U9168 ( .A(n7530), .B(\i_im[3][3] ), .X(n3293) );
  nand_x1_sg U9169 ( .A(n3291), .B(n3292), .X(\update_mask_0/n1386 ) );
  nand_x1_sg U9170 ( .A(n7529), .B(\i_im[3][2] ), .X(n3291) );
  nand_x1_sg U9171 ( .A(n3289), .B(n3290), .X(\update_mask_0/n1387 ) );
  nand_x1_sg U9172 ( .A(n7529), .B(\i_im[3][1] ), .X(n3289) );
  nand_x1_sg U9173 ( .A(n3287), .B(n3288), .X(\update_mask_0/n1388 ) );
  nand_x1_sg U9174 ( .A(n7530), .B(\i_im[3][0] ), .X(n3287) );
  nand_x1_sg U9175 ( .A(n3285), .B(n3286), .X(\update_mask_0/n1389 ) );
  nand_x1_sg U9176 ( .A(n7531), .B(\i_im[2][19] ), .X(n3285) );
  nand_x1_sg U9177 ( .A(n3283), .B(n3284), .X(\update_mask_0/n1390 ) );
  nand_x1_sg U9178 ( .A(n7535), .B(\i_im[2][18] ), .X(n3283) );
  nand_x1_sg U9179 ( .A(n3281), .B(n3282), .X(\update_mask_0/n1391 ) );
  nand_x1_sg U9180 ( .A(n7529), .B(\i_im[2][17] ), .X(n3281) );
  nand_x1_sg U9181 ( .A(n3279), .B(n3280), .X(\update_mask_0/n1392 ) );
  nand_x1_sg U9182 ( .A(n7530), .B(\i_im[2][16] ), .X(n3279) );
  inv_x1_sg U9183 ( .A(n9044), .X(n7043) );
  nand_x1_sg U9184 ( .A(n3277), .B(n3278), .X(\update_mask_0/n1393 ) );
  nand_x1_sg U9185 ( .A(n7531), .B(\i_im[2][15] ), .X(n3277) );
  nand_x1_sg U9186 ( .A(n3275), .B(n3276), .X(\update_mask_0/n1394 ) );
  nand_x1_sg U9187 ( .A(n7535), .B(\i_im[2][14] ), .X(n3275) );
  nand_x1_sg U9188 ( .A(n3273), .B(n3274), .X(\update_mask_0/n1395 ) );
  nand_x1_sg U9189 ( .A(n7533), .B(\i_im[2][13] ), .X(n3273) );
  nand_x1_sg U9190 ( .A(n3271), .B(n3272), .X(\update_mask_0/n1396 ) );
  nand_x1_sg U9191 ( .A(n7535), .B(\i_im[2][12] ), .X(n3271) );
  nand_x1_sg U9192 ( .A(n3269), .B(n3270), .X(\update_mask_0/n1397 ) );
  nand_x1_sg U9193 ( .A(n7534), .B(\i_im[2][11] ), .X(n3269) );
  nand_x1_sg U9194 ( .A(n3267), .B(n3268), .X(\update_mask_0/n1398 ) );
  nand_x1_sg U9195 ( .A(n7531), .B(\i_im[2][10] ), .X(n3267) );
  nand_x1_sg U9196 ( .A(n3265), .B(n3266), .X(\update_mask_0/n1399 ) );
  nand_x1_sg U9197 ( .A(n7530), .B(\i_im[2][9] ), .X(n3265) );
  nand_x1_sg U9198 ( .A(n3263), .B(n3264), .X(\update_mask_0/n1400 ) );
  nand_x1_sg U9199 ( .A(n7527), .B(\i_im[2][8] ), .X(n3263) );
  nand_x1_sg U9200 ( .A(n3261), .B(n3262), .X(\update_mask_0/n1401 ) );
  nand_x1_sg U9201 ( .A(n7535), .B(\i_im[2][7] ), .X(n3261) );
  nand_x1_sg U9202 ( .A(n3259), .B(n3260), .X(\update_mask_0/n1402 ) );
  nand_x1_sg U9203 ( .A(n7535), .B(\i_im[2][6] ), .X(n3259) );
  nand_x1_sg U9204 ( .A(n3257), .B(n3258), .X(\update_mask_0/n1403 ) );
  nand_x1_sg U9205 ( .A(n7533), .B(\i_im[2][5] ), .X(n3257) );
  nand_x1_sg U9206 ( .A(n3255), .B(n3256), .X(\update_mask_0/n1404 ) );
  nand_x1_sg U9207 ( .A(n7530), .B(\i_im[2][4] ), .X(n3255) );
  nand_x1_sg U9208 ( .A(n3253), .B(n3254), .X(\update_mask_0/n1405 ) );
  nand_x1_sg U9209 ( .A(n7529), .B(\i_im[2][3] ), .X(n3253) );
  nand_x1_sg U9210 ( .A(n3251), .B(n3252), .X(\update_mask_0/n1406 ) );
  nand_x1_sg U9211 ( .A(n7527), .B(\i_im[2][2] ), .X(n3251) );
  nand_x1_sg U9212 ( .A(n3249), .B(n3250), .X(\update_mask_0/n1407 ) );
  nand_x1_sg U9213 ( .A(n7533), .B(\i_im[2][1] ), .X(n3249) );
  nand_x1_sg U9214 ( .A(n3247), .B(n3248), .X(\update_mask_0/n1408 ) );
  nand_x1_sg U9215 ( .A(n7533), .B(\i_im[2][0] ), .X(n3247) );
  nand_x1_sg U9216 ( .A(n3245), .B(n3246), .X(\update_mask_0/n1409 ) );
  nand_x1_sg U9217 ( .A(\i_im[1][19] ), .B(n7535), .X(n3245) );
  nand_x1_sg U9218 ( .A(n3243), .B(n3244), .X(\update_mask_0/n1410 ) );
  nand_x1_sg U9219 ( .A(\i_im[1][18] ), .B(n7529), .X(n3243) );
  nand_x1_sg U9220 ( .A(n3241), .B(n3242), .X(\update_mask_0/n1411 ) );
  nand_x1_sg U9221 ( .A(\i_im[1][17] ), .B(n7530), .X(n3241) );
  inv_x1_sg U9222 ( .A(n9048), .X(n7042) );
  nand_x1_sg U9223 ( .A(n3239), .B(n3240), .X(\update_mask_0/n1412 ) );
  nand_x1_sg U9224 ( .A(\i_im[1][16] ), .B(n7527), .X(n3239) );
  nand_x1_sg U9225 ( .A(n3237), .B(n3238), .X(\update_mask_0/n1413 ) );
  nand_x1_sg U9226 ( .A(\i_im[1][15] ), .B(n7536), .X(n3237) );
  nand_x1_sg U9227 ( .A(n3235), .B(n3236), .X(\update_mask_0/n1414 ) );
  nand_x1_sg U9228 ( .A(\i_im[1][14] ), .B(n7529), .X(n3235) );
  nand_x1_sg U9229 ( .A(n3233), .B(n3234), .X(\update_mask_0/n1415 ) );
  nand_x1_sg U9230 ( .A(\i_im[1][13] ), .B(n7533), .X(n3233) );
  nand_x1_sg U9231 ( .A(n3231), .B(n3232), .X(\update_mask_0/n1416 ) );
  nand_x1_sg U9232 ( .A(\i_im[1][12] ), .B(n7528), .X(n3231) );
  nand_x1_sg U9233 ( .A(n3229), .B(n3230), .X(\update_mask_0/n1417 ) );
  nand_x1_sg U9234 ( .A(\i_im[1][11] ), .B(n7536), .X(n3229) );
  nand_x1_sg U9235 ( .A(n3227), .B(n3228), .X(\update_mask_0/n1418 ) );
  nand_x1_sg U9236 ( .A(\i_im[1][10] ), .B(n7536), .X(n3227) );
  nand_x1_sg U9237 ( .A(n3225), .B(n3226), .X(\update_mask_0/n1419 ) );
  nand_x1_sg U9238 ( .A(\i_im[1][9] ), .B(n7536), .X(n3225) );
  nand_x1_sg U9239 ( .A(n3223), .B(n3224), .X(\update_mask_0/n1420 ) );
  nand_x1_sg U9240 ( .A(\i_im[1][8] ), .B(n7536), .X(n3223) );
  nand_x1_sg U9241 ( .A(n3221), .B(n3222), .X(\update_mask_0/n1421 ) );
  nand_x1_sg U9242 ( .A(\i_im[1][7] ), .B(n7536), .X(n3221) );
  nand_x1_sg U9243 ( .A(n3219), .B(n3220), .X(\update_mask_0/n1422 ) );
  nand_x1_sg U9244 ( .A(\i_im[1][6] ), .B(n7529), .X(n3219) );
  nand_x1_sg U9245 ( .A(n3217), .B(n3218), .X(\update_mask_0/n1423 ) );
  nand_x1_sg U9246 ( .A(\i_im[1][5] ), .B(n7535), .X(n3217) );
  nand_x1_sg U9247 ( .A(n3215), .B(n3216), .X(\update_mask_0/n1424 ) );
  nand_x1_sg U9248 ( .A(\i_im[1][4] ), .B(n7534), .X(n3215) );
  nand_x1_sg U9249 ( .A(n3213), .B(n3214), .X(\update_mask_0/n1425 ) );
  nand_x1_sg U9250 ( .A(\i_im[1][3] ), .B(n7531), .X(n3213) );
  nand_x1_sg U9251 ( .A(n3211), .B(n3212), .X(\update_mask_0/n1426 ) );
  nand_x1_sg U9252 ( .A(\i_im[1][2] ), .B(n7527), .X(n3211) );
  nand_x1_sg U9253 ( .A(n3209), .B(n3210), .X(\update_mask_0/n1427 ) );
  nand_x1_sg U9254 ( .A(\i_im[1][1] ), .B(n7535), .X(n3209) );
  nand_x1_sg U9255 ( .A(n3207), .B(n3208), .X(\update_mask_0/n1428 ) );
  nand_x1_sg U9256 ( .A(\i_im[1][0] ), .B(n7529), .X(n3207) );
  nand_x1_sg U9257 ( .A(n3205), .B(n3206), .X(\update_mask_0/n1429 ) );
  nand_x1_sg U9258 ( .A(\i_im[0][19] ), .B(n7530), .X(n3205) );
  nand_x1_sg U9259 ( .A(n3203), .B(n3204), .X(\update_mask_0/n1430 ) );
  nand_x1_sg U9260 ( .A(\i_im[0][18] ), .B(n7534), .X(n3203) );
  nand_x1_sg U9261 ( .A(n3201), .B(n3202), .X(\update_mask_0/n1431 ) );
  nand_x1_sg U9262 ( .A(\i_im[0][17] ), .B(n7528), .X(n3201) );
  inv_x1_sg U9263 ( .A(n9052), .X(n6049) );
  nand_x1_sg U9264 ( .A(n3199), .B(n3200), .X(\update_mask_0/n1432 ) );
  nand_x1_sg U9265 ( .A(\i_im[0][16] ), .B(n7530), .X(n3199) );
  nand_x1_sg U9266 ( .A(n3197), .B(n3198), .X(\update_mask_0/n1433 ) );
  nand_x1_sg U9267 ( .A(\i_im[0][15] ), .B(n7530), .X(n3197) );
  nand_x1_sg U9268 ( .A(n3195), .B(n3196), .X(\update_mask_0/n1434 ) );
  nand_x1_sg U9269 ( .A(\i_im[0][14] ), .B(n7528), .X(n3195) );
  nand_x1_sg U9270 ( .A(n3193), .B(n3194), .X(\update_mask_0/n1435 ) );
  nand_x1_sg U9271 ( .A(\i_im[0][13] ), .B(n7529), .X(n3193) );
  nand_x1_sg U9272 ( .A(n3191), .B(n3192), .X(\update_mask_0/n1436 ) );
  nand_x1_sg U9273 ( .A(\i_im[0][12] ), .B(n7528), .X(n3191) );
  nand_x1_sg U9274 ( .A(n3189), .B(n3190), .X(\update_mask_0/n1437 ) );
  nand_x1_sg U9275 ( .A(\i_im[0][11] ), .B(n7527), .X(n3189) );
  nand_x1_sg U9276 ( .A(n3187), .B(n3188), .X(\update_mask_0/n1438 ) );
  nand_x1_sg U9277 ( .A(\i_im[0][10] ), .B(n7531), .X(n3187) );
  nand_x1_sg U9278 ( .A(n3185), .B(n3186), .X(\update_mask_0/n1439 ) );
  nand_x1_sg U9279 ( .A(\i_im[0][9] ), .B(n7535), .X(n3185) );
  nand_x1_sg U9280 ( .A(n3183), .B(n3184), .X(\update_mask_0/n1440 ) );
  nand_x1_sg U9281 ( .A(\i_im[0][8] ), .B(n7531), .X(n3183) );
  nand_x1_sg U9282 ( .A(n3181), .B(n3182), .X(\update_mask_0/n1441 ) );
  nand_x1_sg U9283 ( .A(\i_im[0][7] ), .B(n7529), .X(n3181) );
  nand_x1_sg U9284 ( .A(n3179), .B(n3180), .X(\update_mask_0/n1442 ) );
  nand_x1_sg U9285 ( .A(\i_im[0][6] ), .B(n7530), .X(n3179) );
  nand_x1_sg U9286 ( .A(n3177), .B(n3178), .X(\update_mask_0/n1443 ) );
  nand_x1_sg U9287 ( .A(\i_im[0][5] ), .B(n7531), .X(n3177) );
  nand_x1_sg U9288 ( .A(n3175), .B(n3176), .X(\update_mask_0/n1444 ) );
  nand_x1_sg U9289 ( .A(\i_im[0][4] ), .B(n7529), .X(n3175) );
  nand_x1_sg U9290 ( .A(n3173), .B(n3174), .X(\update_mask_0/n1445 ) );
  nand_x1_sg U9291 ( .A(\i_im[0][3] ), .B(n7530), .X(n3173) );
  nand_x1_sg U9292 ( .A(n3171), .B(n3172), .X(\update_mask_0/n1446 ) );
  nand_x1_sg U9293 ( .A(\i_im[0][2] ), .B(n7531), .X(n3171) );
  nand_x1_sg U9294 ( .A(n3169), .B(n3170), .X(\update_mask_0/n1447 ) );
  nand_x1_sg U9295 ( .A(\i_im[0][1] ), .B(n7529), .X(n3169) );
  nand_x1_sg U9296 ( .A(n3167), .B(n3168), .X(\update_mask_0/n1448 ) );
  nand_x1_sg U9297 ( .A(\i_im[0][0] ), .B(n7530), .X(n3167) );
  nand_x1_sg U9298 ( .A(n3165), .B(n3166), .X(\update_mask_0/n1449 ) );
  nand_x1_sg U9299 ( .A(i_mask[31]), .B(n7531), .X(n3165) );
  nand_x1_sg U9300 ( .A(n3163), .B(n3164), .X(\update_mask_0/n1450 ) );
  nand_x1_sg U9301 ( .A(i_mask[30]), .B(n7531), .X(n3163) );
  nand_x1_sg U9302 ( .A(n3161), .B(n3162), .X(\update_mask_0/n1451 ) );
  nand_x1_sg U9303 ( .A(i_mask[29]), .B(n7531), .X(n3161) );
  nand_x1_sg U9304 ( .A(n3159), .B(n3160), .X(\update_mask_0/n1452 ) );
  nand_x1_sg U9305 ( .A(i_mask[28]), .B(n7531), .X(n3159) );
  nand_x1_sg U9306 ( .A(n3157), .B(n3158), .X(\update_mask_0/n1453 ) );
  nand_x1_sg U9307 ( .A(i_mask[27]), .B(n7531), .X(n3157) );
  nand_x1_sg U9308 ( .A(n3155), .B(n3156), .X(\update_mask_0/n1454 ) );
  nand_x1_sg U9309 ( .A(i_mask[26]), .B(n7531), .X(n3155) );
  nand_x1_sg U9310 ( .A(n3153), .B(n3154), .X(\update_mask_0/n1455 ) );
  nand_x1_sg U9311 ( .A(i_mask[25]), .B(n7531), .X(n3153) );
  nand_x1_sg U9312 ( .A(n3151), .B(n3152), .X(\update_mask_0/n1456 ) );
  nand_x1_sg U9313 ( .A(i_mask[24]), .B(n7531), .X(n3151) );
  nand_x1_sg U9314 ( .A(n3149), .B(n3150), .X(\update_mask_0/n1457 ) );
  nand_x1_sg U9315 ( .A(i_mask[23]), .B(n7531), .X(n3149) );
  nand_x1_sg U9316 ( .A(n3147), .B(n3148), .X(\update_mask_0/n1458 ) );
  nand_x1_sg U9317 ( .A(i_mask[22]), .B(n7530), .X(n3147) );
  nand_x1_sg U9318 ( .A(n3145), .B(n3146), .X(\update_mask_0/n1459 ) );
  nand_x1_sg U9319 ( .A(i_mask[21]), .B(n7530), .X(n3145) );
  nand_x1_sg U9320 ( .A(n3143), .B(n3144), .X(\update_mask_0/n1460 ) );
  nand_x1_sg U9321 ( .A(i_mask[20]), .B(n7530), .X(n3143) );
  nand_x1_sg U9322 ( .A(n3141), .B(n3142), .X(\update_mask_0/n1461 ) );
  nand_x1_sg U9323 ( .A(i_mask[19]), .B(n7530), .X(n3141) );
  nand_x1_sg U9324 ( .A(n3139), .B(n3140), .X(\update_mask_0/n1462 ) );
  nand_x1_sg U9325 ( .A(i_mask[18]), .B(n7530), .X(n3139) );
  nand_x1_sg U9326 ( .A(n3137), .B(n3138), .X(\update_mask_0/n1463 ) );
  nand_x1_sg U9327 ( .A(i_mask[17]), .B(n7530), .X(n3137) );
  nand_x1_sg U9328 ( .A(n3135), .B(n3136), .X(\update_mask_0/n1464 ) );
  nand_x1_sg U9329 ( .A(i_mask[16]), .B(n7530), .X(n3135) );
  nand_x1_sg U9330 ( .A(n3133), .B(n3134), .X(\update_mask_0/n1465 ) );
  nand_x1_sg U9331 ( .A(i_mask[15]), .B(n7530), .X(n3133) );
  nand_x1_sg U9332 ( .A(n3131), .B(n3132), .X(\update_mask_0/n1466 ) );
  nand_x1_sg U9333 ( .A(i_mask[14]), .B(n7530), .X(n3131) );
  nand_x1_sg U9334 ( .A(n3129), .B(n3130), .X(\update_mask_0/n1467 ) );
  nand_x1_sg U9335 ( .A(i_mask[13]), .B(n7529), .X(n3129) );
  nand_x1_sg U9336 ( .A(n3127), .B(n3128), .X(\update_mask_0/n1468 ) );
  nand_x1_sg U9337 ( .A(i_mask[12]), .B(n7529), .X(n3127) );
  nand_x1_sg U9338 ( .A(n3125), .B(n3126), .X(\update_mask_0/n1469 ) );
  nand_x1_sg U9339 ( .A(i_mask[11]), .B(n7529), .X(n3125) );
  nand_x1_sg U9340 ( .A(n3123), .B(n3124), .X(\update_mask_0/n1470 ) );
  nand_x1_sg U9341 ( .A(i_mask[10]), .B(n7529), .X(n3123) );
  nand_x1_sg U9342 ( .A(n3121), .B(n3122), .X(\update_mask_0/n1471 ) );
  nand_x1_sg U9343 ( .A(i_mask[9]), .B(n7529), .X(n3121) );
  nand_x1_sg U9344 ( .A(n3119), .B(n3120), .X(\update_mask_0/n1472 ) );
  nand_x1_sg U9345 ( .A(i_mask[8]), .B(n7529), .X(n3119) );
  nand_x1_sg U9346 ( .A(n3117), .B(n3118), .X(\update_mask_0/n1473 ) );
  nand_x1_sg U9347 ( .A(i_mask[7]), .B(n7529), .X(n3117) );
  nand_x1_sg U9348 ( .A(n3115), .B(n3116), .X(\update_mask_0/n1474 ) );
  nand_x1_sg U9349 ( .A(i_mask[6]), .B(n7529), .X(n3115) );
  nand_x1_sg U9350 ( .A(n3113), .B(n3114), .X(\update_mask_0/n1475 ) );
  nand_x1_sg U9351 ( .A(i_mask[5]), .B(n7529), .X(n3113) );
  nand_x1_sg U9352 ( .A(n3111), .B(n3112), .X(\update_mask_0/n1476 ) );
  nand_x1_sg U9353 ( .A(i_mask[4]), .B(n7534), .X(n3111) );
  nand_x1_sg U9354 ( .A(n3109), .B(n3110), .X(\update_mask_0/n1477 ) );
  nand_x1_sg U9355 ( .A(i_mask[3]), .B(n7534), .X(n3109) );
  nand_x1_sg U9356 ( .A(n3107), .B(n3108), .X(\update_mask_0/n1478 ) );
  nand_x1_sg U9357 ( .A(i_mask[2]), .B(n7527), .X(n3107) );
  nand_x1_sg U9358 ( .A(n3105), .B(n3106), .X(\update_mask_0/n1479 ) );
  nand_x1_sg U9359 ( .A(i_mask[1]), .B(n7529), .X(n3105) );
  nand_x1_sg U9360 ( .A(n3102), .B(n3103), .X(\update_mask_0/n1480 ) );
  nand_x1_sg U9361 ( .A(i_mask[0]), .B(n7527), .X(n3102) );
  nand_x1_sg U9362 ( .A(n5303), .B(n5304), .X(n5884) );
  nand_x1_sg U9363 ( .A(n5295), .B(n5296), .X(n5882) );
  nand_x1_sg U9364 ( .A(n7522), .B(n5297), .X(n5296) );
  nand_x1_sg U9365 ( .A(n9200), .B(n5298), .X(n5297) );
  nand_x1_sg U9366 ( .A(n5300), .B(n5301), .X(n5883) );
  nand_x1_sg U9367 ( .A(n5288), .B(n5289), .X(n5880) );
  nand_x1_sg U9368 ( .A(n5278), .B(n5279), .X(n5878) );
  nand_x1_sg U9369 ( .A(n5281), .B(n5282), .X(n5879) );
  nand_x1_sg U9370 ( .A(n3810), .B(n3811), .X(\update_mask_0/n1128 ) );
  nor_x4_sg U9371 ( .A(n7526), .B(n9230), .X(n3827) );
  inv_x4_sg U9372 ( .A(n4799), .X(n9230) );
  inv_x2_sg U9373 ( .A(\update_output_0/N29 ), .X(n6001) );
  nor_x4_sg U9374 ( .A(n7526), .B(n9225), .X(n3879) );
  inv_x4_sg U9375 ( .A(n5009), .X(n9225) );
  nor_x4_sg U9376 ( .A(n7526), .B(n9231), .X(n3867) );
  inv_x4_sg U9377 ( .A(n4757), .X(n9231) );
  nor_x2_sg U9378 ( .A(n9241), .B(n7526), .X(n3093) );
  nand_x1_sg U9379 ( .A(n4182), .B(n7559), .X(n4300) );
  inv_x2_sg U9380 ( .A(\update_mask_0/reg_out[0][0] ), .X(n6011) );
  inv_x2_sg U9381 ( .A(\update_mask_0/reg_out[0][5] ), .X(n6013) );
  inv_x2_sg U9382 ( .A(\update_mask_0/reg_out[0][10] ), .X(n6015) );
  inv_x2_sg U9383 ( .A(\update_mask_0/reg_out[1][0] ), .X(n6017) );
  inv_x2_sg U9384 ( .A(\update_mask_0/reg_out[1][5] ), .X(n6019) );
  inv_x2_sg U9385 ( .A(\update_mask_0/reg_out[1][10] ), .X(n6021) );
  inv_x2_sg U9386 ( .A(\update_mask_0/reg_out[3][0] ), .X(n6023) );
  inv_x2_sg U9387 ( .A(\update_mask_0/reg_out[3][5] ), .X(n6025) );
  inv_x2_sg U9388 ( .A(\update_mask_0/reg_out[3][10] ), .X(n6027) );
  inv_x2_sg U9389 ( .A(\update_mask_0/reg_out[6][0] ), .X(n6029) );
  inv_x2_sg U9390 ( .A(\update_mask_0/reg_out[6][5] ), .X(n6031) );
  inv_x2_sg U9391 ( .A(\update_mask_0/reg_out[6][10] ), .X(n6033) );
  inv_x2_sg U9392 ( .A(\update_mask_0/reg_out[7][0] ), .X(n6035) );
  inv_x2_sg U9393 ( .A(\update_mask_0/reg_out[7][5] ), .X(n6037) );
  inv_x2_sg U9394 ( .A(\update_mask_0/reg_out[7][10] ), .X(n6039) );
  inv_x2_sg U9395 ( .A(\update_mask_0/reg_out[12][0] ), .X(n6105) );
  inv_x2_sg U9396 ( .A(\update_mask_0/reg_out[12][5] ), .X(n6107) );
  inv_x2_sg U9397 ( .A(\update_mask_0/reg_out[12][10] ), .X(n6109) );
  nor_x4_sg U9398 ( .A(n7526), .B(n9228), .X(n3840) );
  inv_x4_sg U9399 ( .A(n4883), .X(n9228) );
  nor_x4_sg U9400 ( .A(n7526), .B(n9224), .X(n3846) );
  inv_x4_sg U9401 ( .A(n5081), .X(n9224) );
  nor_x4_sg U9402 ( .A(n4184), .B(n8988), .X(n858) );
  inv_x8_sg U9403 ( .A(n1512), .X(n8988) );
  nor_x2_sg U9404 ( .A(n9219), .B(n7048), .X(n2064) );
  inv_x2_sg U9405 ( .A(\update_mask_0/reg_out[0][1] ), .X(n6157) );
  inv_x2_sg U9406 ( .A(\update_mask_0/reg_out[0][6] ), .X(n6159) );
  inv_x2_sg U9407 ( .A(\update_mask_0/reg_out[0][11] ), .X(n6161) );
  inv_x2_sg U9408 ( .A(\update_mask_0/reg_out[1][1] ), .X(n6051) );
  inv_x2_sg U9409 ( .A(\update_mask_0/reg_out[1][6] ), .X(n6053) );
  inv_x2_sg U9410 ( .A(\update_mask_0/reg_out[1][11] ), .X(n6055) );
  inv_x2_sg U9411 ( .A(\update_mask_0/reg_out[2][0] ), .X(n6057) );
  inv_x2_sg U9412 ( .A(\update_mask_0/reg_out[2][5] ), .X(n6059) );
  inv_x2_sg U9413 ( .A(\update_mask_0/reg_out[2][10] ), .X(n6061) );
  inv_x2_sg U9414 ( .A(\update_mask_0/reg_out[3][1] ), .X(n6063) );
  inv_x2_sg U9415 ( .A(\update_mask_0/reg_out[3][6] ), .X(n6065) );
  inv_x2_sg U9416 ( .A(\update_mask_0/reg_out[3][11] ), .X(n6067) );
  inv_x2_sg U9417 ( .A(\update_mask_0/reg_out[4][0] ), .X(n6069) );
  inv_x2_sg U9418 ( .A(\update_mask_0/reg_out[4][5] ), .X(n6071) );
  inv_x2_sg U9419 ( .A(\update_mask_0/reg_out[4][10] ), .X(n6073) );
  inv_x2_sg U9420 ( .A(\update_mask_0/reg_out[5][0] ), .X(n6075) );
  inv_x2_sg U9421 ( .A(\update_mask_0/reg_out[5][5] ), .X(n6077) );
  inv_x2_sg U9422 ( .A(\update_mask_0/reg_out[5][10] ), .X(n6079) );
  inv_x2_sg U9423 ( .A(\update_mask_0/reg_out[6][1] ), .X(n6195) );
  inv_x2_sg U9424 ( .A(\update_mask_0/reg_out[6][6] ), .X(n6197) );
  inv_x2_sg U9425 ( .A(\update_mask_0/reg_out[6][11] ), .X(n6199) );
  inv_x2_sg U9426 ( .A(\update_mask_0/reg_out[7][1] ), .X(n6081) );
  inv_x2_sg U9427 ( .A(\update_mask_0/reg_out[7][6] ), .X(n6083) );
  inv_x2_sg U9428 ( .A(\update_mask_0/reg_out[7][11] ), .X(n6085) );
  inv_x2_sg U9429 ( .A(\update_mask_0/reg_out[9][0] ), .X(n6087) );
  inv_x2_sg U9430 ( .A(\update_mask_0/reg_out[9][5] ), .X(n6089) );
  inv_x2_sg U9431 ( .A(\update_mask_0/reg_out[9][10] ), .X(n6091) );
  inv_x2_sg U9432 ( .A(\update_mask_0/reg_out[10][0] ), .X(n6093) );
  inv_x2_sg U9433 ( .A(\update_mask_0/reg_out[10][5] ), .X(n6095) );
  inv_x2_sg U9434 ( .A(\update_mask_0/reg_out[10][10] ), .X(n6097) );
  inv_x2_sg U9435 ( .A(\update_mask_0/reg_out[11][0] ), .X(n6099) );
  inv_x2_sg U9436 ( .A(\update_mask_0/reg_out[11][5] ), .X(n6101) );
  inv_x2_sg U9437 ( .A(\update_mask_0/reg_out[11][10] ), .X(n6103) );
  inv_x2_sg U9438 ( .A(\update_mask_0/reg_out[12][1] ), .X(n6221) );
  inv_x2_sg U9439 ( .A(\update_mask_0/reg_out[12][6] ), .X(n6223) );
  inv_x2_sg U9440 ( .A(\update_mask_0/reg_out[12][11] ), .X(n6225) );
  inv_x2_sg U9441 ( .A(\update_mask_0/reg_out[15][0] ), .X(n6111) );
  inv_x2_sg U9442 ( .A(\update_mask_0/reg_out[15][5] ), .X(n6113) );
  inv_x2_sg U9443 ( .A(\update_mask_0/reg_out[15][10] ), .X(n6115) );
  nor_x2_sg U9444 ( .A(n4303), .B(n7526), .X(n4302) );
  inv_x2_sg U9445 ( .A(\update_mask_0/reg_out[8][2] ), .X(n6119) );
  inv_x2_sg U9446 ( .A(\update_mask_0/reg_out[8][7] ), .X(n6121) );
  inv_x2_sg U9447 ( .A(\update_mask_0/reg_out[8][12] ), .X(n6123) );
  inv_x2_sg U9448 ( .A(\update_mask_0/reg_out[8][16] ), .X(n6125) );
  inv_x2_sg U9449 ( .A(\update_mask_0/reg_out[9][16] ), .X(n6127) );
  inv_x2_sg U9450 ( .A(\update_mask_0/reg_out[10][16] ), .X(n6129) );
  inv_x2_sg U9451 ( .A(\update_mask_0/reg_out[11][16] ), .X(n6131) );
  inv_x2_sg U9452 ( .A(\update_mask_0/reg_out[12][16] ), .X(n6133) );
  inv_x2_sg U9453 ( .A(\update_mask_0/reg_out[13][2] ), .X(n6135) );
  inv_x2_sg U9454 ( .A(\update_mask_0/reg_out[13][7] ), .X(n6137) );
  inv_x2_sg U9455 ( .A(\update_mask_0/reg_out[13][12] ), .X(n6139) );
  inv_x2_sg U9456 ( .A(\update_mask_0/reg_out[13][16] ), .X(n6141) );
  inv_x2_sg U9457 ( .A(\update_mask_0/reg_out[14][2] ), .X(n6143) );
  inv_x2_sg U9458 ( .A(\update_mask_0/reg_out[14][7] ), .X(n6145) );
  inv_x2_sg U9459 ( .A(\update_mask_0/reg_out[14][12] ), .X(n6147) );
  inv_x2_sg U9460 ( .A(\update_mask_0/reg_out[15][16] ), .X(n6149) );
  nor_x4_sg U9461 ( .A(n7526), .B(n9229), .X(n3855) );
  inv_x4_sg U9462 ( .A(n4841), .X(n9229) );
  nor_x4_sg U9463 ( .A(n7526), .B(n9223), .X(n3858) );
  inv_x4_sg U9464 ( .A(n5117), .X(n9223) );
  inv_x4_sg U9465 ( .A(n5993), .X(n5994) );
  nor_x8_sg U9466 ( .A(n4184), .B(n9247), .X(n859) );
  inv_x8_sg U9467 ( .A(n1510), .X(n9247) );
  nor_x4_sg U9468 ( .A(n5236), .B(n9241), .X(n4416) );
  nor_x2_sg U9469 ( .A(n9219), .B(n9215), .X(n2055) );
  nand_x8_sg U9470 ( .A(n6050), .B(n9213), .X(n1872) );
  nor_x2_sg U9471 ( .A(n6377), .B(n7310), .X(n6050) );
  nand_x8_sg U9472 ( .A(n7308), .B(n1965), .X(n1876) );
  nor_x2_sg U9473 ( .A(n6377), .B(n7310), .X(n1965) );
  inv_x2_sg U9474 ( .A(\update_mask_0/reg_out[0][2] ), .X(n7049) );
  inv_x2_sg U9475 ( .A(\update_mask_0/reg_out[0][7] ), .X(n7051) );
  inv_x2_sg U9476 ( .A(\update_mask_0/reg_out[0][12] ), .X(n7053) );
  inv_x2_sg U9477 ( .A(\update_mask_0/reg_out[1][2] ), .X(n7055) );
  inv_x2_sg U9478 ( .A(\update_mask_0/reg_out[1][7] ), .X(n7057) );
  inv_x2_sg U9479 ( .A(\update_mask_0/reg_out[1][12] ), .X(n7059) );
  inv_x2_sg U9480 ( .A(\update_mask_0/reg_out[2][1] ), .X(n6163) );
  inv_x2_sg U9481 ( .A(\update_mask_0/reg_out[2][6] ), .X(n6165) );
  inv_x2_sg U9482 ( .A(\update_mask_0/reg_out[2][11] ), .X(n6167) );
  inv_x2_sg U9483 ( .A(\update_mask_0/reg_out[3][2] ), .X(n6171) );
  inv_x2_sg U9484 ( .A(\update_mask_0/reg_out[3][7] ), .X(n6173) );
  inv_x2_sg U9485 ( .A(\update_mask_0/reg_out[3][12] ), .X(n6175) );
  inv_x2_sg U9486 ( .A(\update_mask_0/reg_out[4][1] ), .X(n6179) );
  inv_x2_sg U9487 ( .A(\update_mask_0/reg_out[4][6] ), .X(n6181) );
  inv_x2_sg U9488 ( .A(\update_mask_0/reg_out[4][11] ), .X(n6183) );
  inv_x2_sg U9489 ( .A(\update_mask_0/reg_out[5][1] ), .X(n6187) );
  inv_x2_sg U9490 ( .A(\update_mask_0/reg_out[5][6] ), .X(n6189) );
  inv_x2_sg U9491 ( .A(\update_mask_0/reg_out[5][11] ), .X(n6191) );
  inv_x2_sg U9492 ( .A(\update_mask_0/reg_out[6][2] ), .X(n7095) );
  inv_x2_sg U9493 ( .A(\update_mask_0/reg_out[6][7] ), .X(n7097) );
  inv_x2_sg U9494 ( .A(\update_mask_0/reg_out[6][12] ), .X(n7099) );
  inv_x2_sg U9495 ( .A(\update_mask_0/reg_out[7][2] ), .X(n7105) );
  inv_x2_sg U9496 ( .A(\update_mask_0/reg_out[7][7] ), .X(n7107) );
  inv_x2_sg U9497 ( .A(\update_mask_0/reg_out[7][12] ), .X(n7109) );
  inv_x2_sg U9498 ( .A(\update_mask_0/reg_out[9][1] ), .X(n6203) );
  inv_x2_sg U9499 ( .A(\update_mask_0/reg_out[9][6] ), .X(n6205) );
  inv_x2_sg U9500 ( .A(\update_mask_0/reg_out[9][11] ), .X(n6207) );
  inv_x2_sg U9501 ( .A(\update_mask_0/reg_out[10][1] ), .X(n6209) );
  inv_x2_sg U9502 ( .A(\update_mask_0/reg_out[10][6] ), .X(n6211) );
  inv_x2_sg U9503 ( .A(\update_mask_0/reg_out[10][11] ), .X(n6213) );
  inv_x2_sg U9504 ( .A(\update_mask_0/reg_out[11][1] ), .X(n6215) );
  inv_x2_sg U9505 ( .A(\update_mask_0/reg_out[11][6] ), .X(n6217) );
  inv_x2_sg U9506 ( .A(\update_mask_0/reg_out[11][11] ), .X(n6219) );
  inv_x2_sg U9507 ( .A(\update_mask_0/reg_out[12][2] ), .X(n7139) );
  inv_x2_sg U9508 ( .A(\update_mask_0/reg_out[12][7] ), .X(n7141) );
  inv_x2_sg U9509 ( .A(\update_mask_0/reg_out[12][12] ), .X(n7143) );
  inv_x2_sg U9510 ( .A(\update_mask_0/reg_out[15][1] ), .X(n6227) );
  inv_x2_sg U9511 ( .A(\update_mask_0/reg_out[15][6] ), .X(n6229) );
  inv_x2_sg U9512 ( .A(\update_mask_0/reg_out[15][11] ), .X(n6231) );
  inv_x2_sg U9513 ( .A(\update_mask_0/reg_out[0][15] ), .X(n6341) );
  inv_x2_sg U9514 ( .A(\update_mask_0/reg_out[1][15] ), .X(n6117) );
  inv_x2_sg U9515 ( .A(\update_mask_0/reg_out[8][3] ), .X(n6345) );
  inv_x2_sg U9516 ( .A(\update_mask_0/reg_out[8][8] ), .X(n6347) );
  inv_x2_sg U9517 ( .A(\update_mask_0/reg_out[8][13] ), .X(n6349) );
  inv_x2_sg U9518 ( .A(\update_mask_0/reg_out[8][17] ), .X(n6351) );
  inv_x2_sg U9519 ( .A(\update_mask_0/reg_out[9][17] ), .X(n6353) );
  inv_x2_sg U9520 ( .A(\update_mask_0/reg_out[10][17] ), .X(n6355) );
  inv_x2_sg U9521 ( .A(\update_mask_0/reg_out[11][17] ), .X(n6357) );
  inv_x2_sg U9522 ( .A(\update_mask_0/reg_out[12][17] ), .X(n6359) );
  inv_x2_sg U9523 ( .A(\update_mask_0/reg_out[13][3] ), .X(n6361) );
  inv_x2_sg U9524 ( .A(\update_mask_0/reg_out[13][8] ), .X(n6363) );
  inv_x2_sg U9525 ( .A(\update_mask_0/reg_out[13][13] ), .X(n6365) );
  inv_x2_sg U9526 ( .A(\update_mask_0/reg_out[13][17] ), .X(n6367) );
  inv_x2_sg U9527 ( .A(\update_mask_0/reg_out[14][3] ), .X(n6369) );
  inv_x2_sg U9528 ( .A(\update_mask_0/reg_out[14][8] ), .X(n6371) );
  inv_x2_sg U9529 ( .A(\update_mask_0/reg_out[14][13] ), .X(n6373) );
  inv_x2_sg U9530 ( .A(\update_mask_0/reg_out[15][17] ), .X(n6375) );
  nor_x4_sg U9531 ( .A(n7526), .B(n9221), .X(n3870) );
  inv_x4_sg U9532 ( .A(n5193), .X(n9221) );
  nor_x4_sg U9533 ( .A(n7526), .B(n9227), .X(n3876) );
  inv_x4_sg U9534 ( .A(n4925), .X(n9227) );
  nor_x4_sg U9535 ( .A(n7526), .B(n9239), .X(n3831) );
  inv_x4_sg U9536 ( .A(n4408), .X(n9239) );
  inv_x2_sg U9537 ( .A(n5995), .X(n5996) );
  inv_x2_sg U9538 ( .A(n5997), .X(n5998) );
  inv_x2_sg U9539 ( .A(n5999), .X(n6000) );
  inv_x4_sg U9540 ( .A(n6001), .X(n6002) );
  nor_x8_sg U9541 ( .A(n5236), .B(n7559), .X(n4452) );
  nor_x2_sg U9542 ( .A(n7316), .B(n6340), .X(n2065) );
  inv_x2_sg U9543 ( .A(\update_mask_0/reg_out[2][2] ), .X(n7061) );
  inv_x2_sg U9544 ( .A(\update_mask_0/reg_out[2][7] ), .X(n7063) );
  inv_x2_sg U9545 ( .A(\update_mask_0/reg_out[2][12] ), .X(n7065) );
  inv_x2_sg U9546 ( .A(\update_mask_0/reg_out[2][17] ), .X(n6169) );
  inv_x2_sg U9547 ( .A(\update_mask_0/reg_out[3][17] ), .X(n6177) );
  inv_x2_sg U9548 ( .A(\update_mask_0/reg_out[4][2] ), .X(n7075) );
  inv_x2_sg U9549 ( .A(\update_mask_0/reg_out[4][7] ), .X(n7077) );
  inv_x2_sg U9550 ( .A(\update_mask_0/reg_out[4][12] ), .X(n7079) );
  inv_x2_sg U9551 ( .A(\update_mask_0/reg_out[4][17] ), .X(n6185) );
  inv_x2_sg U9552 ( .A(\update_mask_0/reg_out[5][2] ), .X(n7085) );
  inv_x2_sg U9553 ( .A(\update_mask_0/reg_out[5][7] ), .X(n7087) );
  inv_x2_sg U9554 ( .A(\update_mask_0/reg_out[5][12] ), .X(n7089) );
  inv_x2_sg U9555 ( .A(\update_mask_0/reg_out[5][17] ), .X(n6193) );
  inv_x2_sg U9556 ( .A(\update_mask_0/reg_out[7][15] ), .X(n6201) );
  inv_x2_sg U9557 ( .A(\update_mask_0/reg_out[9][2] ), .X(n7115) );
  inv_x2_sg U9558 ( .A(\update_mask_0/reg_out[9][7] ), .X(n7117) );
  inv_x2_sg U9559 ( .A(\update_mask_0/reg_out[9][12] ), .X(n7119) );
  inv_x2_sg U9560 ( .A(\update_mask_0/reg_out[10][2] ), .X(n7123) );
  inv_x2_sg U9561 ( .A(\update_mask_0/reg_out[10][7] ), .X(n7125) );
  inv_x2_sg U9562 ( .A(\update_mask_0/reg_out[10][12] ), .X(n7127) );
  inv_x2_sg U9563 ( .A(\update_mask_0/reg_out[11][2] ), .X(n7131) );
  inv_x2_sg U9564 ( .A(\update_mask_0/reg_out[11][7] ), .X(n7133) );
  inv_x2_sg U9565 ( .A(\update_mask_0/reg_out[11][12] ), .X(n7135) );
  inv_x2_sg U9566 ( .A(\update_mask_0/reg_out[15][2] ), .X(n7151) );
  inv_x2_sg U9567 ( .A(\update_mask_0/reg_out[15][7] ), .X(n7153) );
  inv_x2_sg U9568 ( .A(\update_mask_0/reg_out[15][12] ), .X(n7155) );
  inv_x2_sg U9569 ( .A(\update_mask_0/reg_i_mask [0]), .X(n6233) );
  inv_x2_sg U9570 ( .A(\update_mask_0/reg_out[4][3] ), .X(n6235) );
  inv_x2_sg U9571 ( .A(\update_mask_0/reg_out[4][8] ), .X(n6237) );
  inv_x2_sg U9572 ( .A(\update_mask_0/reg_out[4][13] ), .X(n6239) );
  inv_x2_sg U9573 ( .A(\update_mask_0/reg_out[5][3] ), .X(n6241) );
  inv_x2_sg U9574 ( .A(\update_mask_0/reg_out[5][8] ), .X(n6243) );
  inv_x2_sg U9575 ( .A(\update_mask_0/reg_out[5][13] ), .X(n6245) );
  inv_x2_sg U9576 ( .A(\update_mask_0/reg_out[9][3] ), .X(n6247) );
  inv_x2_sg U9577 ( .A(\update_mask_0/reg_out[9][8] ), .X(n6249) );
  inv_x2_sg U9578 ( .A(\update_mask_0/reg_out[9][13] ), .X(n6251) );
  inv_x2_sg U9579 ( .A(\update_mask_0/reg_out[11][3] ), .X(n6253) );
  inv_x2_sg U9580 ( .A(\update_mask_0/reg_out[11][8] ), .X(n6255) );
  inv_x2_sg U9581 ( .A(\update_mask_0/reg_out[11][13] ), .X(n6257) );
  inv_x2_sg U9582 ( .A(\update_mask_0/reg_out[15][3] ), .X(n6259) );
  inv_x2_sg U9583 ( .A(\update_mask_0/reg_out[15][8] ), .X(n6261) );
  inv_x2_sg U9584 ( .A(\update_mask_0/reg_out[15][13] ), .X(n6263) );
  inv_x2_sg U9585 ( .A(\update_mask_0/reg_out[1][18] ), .X(n6265) );
  inv_x2_sg U9586 ( .A(\update_mask_0/reg_out[8][0] ), .X(n6267) );
  inv_x2_sg U9587 ( .A(\update_mask_0/reg_out[8][5] ), .X(n6269) );
  inv_x2_sg U9588 ( .A(\update_mask_0/reg_out[8][10] ), .X(n6271) );
  inv_x2_sg U9589 ( .A(\update_mask_0/reg_out[13][0] ), .X(n6273) );
  inv_x2_sg U9590 ( .A(\update_mask_0/reg_out[13][5] ), .X(n6275) );
  inv_x2_sg U9591 ( .A(\update_mask_0/reg_out[13][10] ), .X(n6277) );
  inv_x2_sg U9592 ( .A(\update_mask_0/reg_out[14][0] ), .X(n6279) );
  inv_x2_sg U9593 ( .A(\update_mask_0/reg_out[14][5] ), .X(n6281) );
  inv_x2_sg U9594 ( .A(\update_mask_0/reg_out[14][10] ), .X(n6283) );
  inv_x2_sg U9595 ( .A(\update_mask_0/reg_out[0][3] ), .X(n6285) );
  inv_x2_sg U9596 ( .A(\update_mask_0/reg_out[0][8] ), .X(n6287) );
  inv_x2_sg U9597 ( .A(\update_mask_0/reg_out[0][13] ), .X(n6289) );
  inv_x2_sg U9598 ( .A(\update_mask_0/reg_out[1][3] ), .X(n6291) );
  inv_x2_sg U9599 ( .A(\update_mask_0/reg_out[1][8] ), .X(n6293) );
  inv_x2_sg U9600 ( .A(\update_mask_0/reg_out[1][13] ), .X(n6295) );
  inv_x2_sg U9601 ( .A(\update_mask_0/reg_out[2][3] ), .X(n6297) );
  inv_x2_sg U9602 ( .A(\update_mask_0/reg_out[2][8] ), .X(n6299) );
  inv_x2_sg U9603 ( .A(\update_mask_0/reg_out[2][13] ), .X(n6301) );
  inv_x2_sg U9604 ( .A(\update_mask_0/reg_out[3][3] ), .X(n6303) );
  inv_x2_sg U9605 ( .A(\update_mask_0/reg_out[3][8] ), .X(n6305) );
  inv_x2_sg U9606 ( .A(\update_mask_0/reg_out[3][13] ), .X(n6307) );
  inv_x2_sg U9607 ( .A(\update_mask_0/reg_out[6][3] ), .X(n6309) );
  inv_x2_sg U9608 ( .A(\update_mask_0/reg_out[6][8] ), .X(n6311) );
  inv_x2_sg U9609 ( .A(\update_mask_0/reg_out[6][13] ), .X(n6313) );
  inv_x2_sg U9610 ( .A(\update_mask_0/reg_out[6][17] ), .X(n6315) );
  inv_x2_sg U9611 ( .A(\update_mask_0/reg_out[7][3] ), .X(n6317) );
  inv_x2_sg U9612 ( .A(\update_mask_0/reg_out[7][8] ), .X(n6319) );
  inv_x2_sg U9613 ( .A(\update_mask_0/reg_out[7][13] ), .X(n6321) );
  inv_x2_sg U9614 ( .A(\update_mask_0/reg_out[7][17] ), .X(n6323) );
  inv_x2_sg U9615 ( .A(\update_mask_0/reg_out[10][3] ), .X(n6325) );
  inv_x2_sg U9616 ( .A(\update_mask_0/reg_out[10][8] ), .X(n6327) );
  inv_x2_sg U9617 ( .A(\update_mask_0/reg_out[10][13] ), .X(n6329) );
  inv_x2_sg U9618 ( .A(\update_mask_0/reg_out[12][3] ), .X(n6331) );
  inv_x2_sg U9619 ( .A(\update_mask_0/reg_out[12][8] ), .X(n6333) );
  inv_x2_sg U9620 ( .A(\update_mask_0/reg_out[12][13] ), .X(n6335) );
  inv_x2_sg U9621 ( .A(\update_mask_0/reg_out[14][17] ), .X(n6337) );
  inv_x2_sg U9622 ( .A(\update_mask_0/reg_out[0][16] ), .X(n7267) );
  inv_x2_sg U9623 ( .A(\update_mask_0/reg_out[1][16] ), .X(n7269) );
  inv_x2_sg U9624 ( .A(\update_mask_0/reg_out[0][18] ), .X(n6343) );
  inv_x2_sg U9625 ( .A(\update_mask_0/reg_out[8][4] ), .X(n7273) );
  inv_x2_sg U9626 ( .A(\update_mask_0/reg_out[8][9] ), .X(n7275) );
  inv_x2_sg U9627 ( .A(\update_mask_0/reg_out[8][14] ), .X(n7277) );
  inv_x2_sg U9628 ( .A(\update_mask_0/reg_out[8][18] ), .X(n7279) );
  inv_x2_sg U9629 ( .A(\update_mask_0/reg_out[9][18] ), .X(n7281) );
  inv_x2_sg U9630 ( .A(\update_mask_0/reg_out[10][18] ), .X(n7283) );
  inv_x2_sg U9631 ( .A(\update_mask_0/reg_out[11][18] ), .X(n7285) );
  inv_x2_sg U9632 ( .A(\update_mask_0/reg_out[12][18] ), .X(n7287) );
  inv_x2_sg U9633 ( .A(\update_mask_0/reg_out[13][4] ), .X(n7289) );
  inv_x2_sg U9634 ( .A(\update_mask_0/reg_out[13][9] ), .X(n7291) );
  inv_x2_sg U9635 ( .A(\update_mask_0/reg_out[13][14] ), .X(n7293) );
  inv_x2_sg U9636 ( .A(\update_mask_0/reg_out[13][18] ), .X(n7295) );
  inv_x2_sg U9637 ( .A(\update_mask_0/reg_out[14][4] ), .X(n7297) );
  inv_x2_sg U9638 ( .A(\update_mask_0/reg_out[14][9] ), .X(n7299) );
  inv_x2_sg U9639 ( .A(\update_mask_0/reg_out[14][14] ), .X(n7301) );
  inv_x2_sg U9640 ( .A(\update_mask_0/reg_out[15][18] ), .X(n7303) );
  nor_x2_sg U9641 ( .A(n5286), .B(n7308), .X(n1594) );
  inv_x2_sg U9642 ( .A(\update_mask_0/N29 ), .X(n6378) );
  inv_x2_sg U9643 ( .A(\update_output_0/N27 ), .X(n7038) );
  nor_x4_sg U9644 ( .A(n7526), .B(n9226), .X(n3834) );
  inv_x4_sg U9645 ( .A(n4967), .X(n9226) );
  nor_x4_sg U9646 ( .A(n7526), .B(n9235), .X(n3861) );
  inv_x4_sg U9647 ( .A(n4587), .X(n9235) );
  nor_x4_sg U9648 ( .A(n7526), .B(n9238), .X(n3882) );
  inv_x4_sg U9649 ( .A(n4461), .X(n9238) );
  inv_x8_sg U9650 ( .A(n6151), .X(n6152) );
  inv_x4_sg U9651 ( .A(n7310), .X(n9077) );
  inv_x2_sg U9652 ( .A(n6003), .X(n6004) );
  inv_x2_sg U9653 ( .A(n6005), .X(n6006) );
  inv_x2_sg U9654 ( .A(n6007), .X(n6008) );
  inv_x2_sg U9655 ( .A(n6009), .X(n6010) );
  inv_x4_sg U9656 ( .A(n6011), .X(n6012) );
  inv_x4_sg U9657 ( .A(n6013), .X(n6014) );
  inv_x4_sg U9658 ( .A(n6015), .X(n6016) );
  inv_x4_sg U9659 ( .A(n6017), .X(n6018) );
  inv_x4_sg U9660 ( .A(n6019), .X(n6020) );
  inv_x4_sg U9661 ( .A(n6021), .X(n6022) );
  inv_x4_sg U9662 ( .A(n6023), .X(n6024) );
  inv_x4_sg U9663 ( .A(n6025), .X(n6026) );
  inv_x4_sg U9664 ( .A(n6027), .X(n6028) );
  inv_x4_sg U9665 ( .A(n6029), .X(n6030) );
  inv_x4_sg U9666 ( .A(n6031), .X(n6032) );
  inv_x4_sg U9667 ( .A(n6033), .X(n6034) );
  inv_x4_sg U9668 ( .A(n6035), .X(n6036) );
  inv_x4_sg U9669 ( .A(n6037), .X(n6038) );
  inv_x4_sg U9670 ( .A(n6039), .X(n6040) );
  nor_x4_sg U9671 ( .A(n6383), .B(n9219), .X(n5302) );
  nor_x8_sg U9672 ( .A(n4192), .B(n4184), .X(n871) );
  nor_x8_sg U9673 ( .A(n5236), .B(n7559), .X(n7424) );
  inv_x2_sg U9674 ( .A(\update_mask_0/reg_i_mask [3]), .X(n7047) );
  inv_x2_sg U9675 ( .A(\update_mask_0/reg_out[2][18] ), .X(n7069) );
  inv_x2_sg U9676 ( .A(\update_mask_0/reg_out[3][18] ), .X(n7073) );
  inv_x2_sg U9677 ( .A(\update_mask_0/reg_out[4][15] ), .X(n7081) );
  inv_x2_sg U9678 ( .A(\update_mask_0/reg_out[4][18] ), .X(n7083) );
  inv_x2_sg U9679 ( .A(\update_mask_0/reg_out[5][18] ), .X(n7093) );
  inv_x2_sg U9680 ( .A(\update_mask_0/reg_out[7][16] ), .X(n7111) );
  inv_x2_sg U9681 ( .A(\update_mask_0/reg_out[12][15] ), .X(n7145) );
  inv_x2_sg U9682 ( .A(\update_mask_0/reg_out[4][4] ), .X(n7161) );
  inv_x2_sg U9683 ( .A(\update_mask_0/reg_out[4][9] ), .X(n7163) );
  inv_x2_sg U9684 ( .A(\update_mask_0/reg_out[4][14] ), .X(n7165) );
  inv_x2_sg U9685 ( .A(\update_mask_0/reg_out[5][4] ), .X(n7167) );
  inv_x2_sg U9686 ( .A(\update_mask_0/reg_out[5][9] ), .X(n7169) );
  inv_x2_sg U9687 ( .A(\update_mask_0/reg_out[5][14] ), .X(n7171) );
  inv_x2_sg U9688 ( .A(\update_mask_0/reg_out[9][4] ), .X(n7173) );
  inv_x2_sg U9689 ( .A(\update_mask_0/reg_out[9][9] ), .X(n7175) );
  inv_x2_sg U9690 ( .A(\update_mask_0/reg_out[9][14] ), .X(n7177) );
  inv_x2_sg U9691 ( .A(\update_mask_0/reg_out[11][4] ), .X(n7179) );
  inv_x2_sg U9692 ( .A(\update_mask_0/reg_out[11][9] ), .X(n7181) );
  inv_x2_sg U9693 ( .A(\update_mask_0/reg_out[11][14] ), .X(n7183) );
  inv_x2_sg U9694 ( .A(\update_mask_0/reg_out[15][4] ), .X(n7185) );
  inv_x2_sg U9695 ( .A(\update_mask_0/reg_out[15][9] ), .X(n7187) );
  inv_x2_sg U9696 ( .A(\update_mask_0/reg_out[15][14] ), .X(n7189) );
  inv_x2_sg U9697 ( .A(n9569), .X(n7040) );
  inv_x2_sg U9698 ( .A(\update_mask_0/reg_out[1][19] ), .X(n7191) );
  inv_x2_sg U9699 ( .A(\update_mask_0/reg_out[8][1] ), .X(n7193) );
  inv_x2_sg U9700 ( .A(\update_mask_0/reg_out[8][6] ), .X(n7195) );
  inv_x2_sg U9701 ( .A(\update_mask_0/reg_out[8][11] ), .X(n7197) );
  inv_x2_sg U9702 ( .A(\update_mask_0/reg_out[13][1] ), .X(n7199) );
  inv_x2_sg U9703 ( .A(\update_mask_0/reg_out[13][6] ), .X(n7201) );
  inv_x2_sg U9704 ( .A(\update_mask_0/reg_out[13][11] ), .X(n7203) );
  inv_x2_sg U9705 ( .A(\update_mask_0/reg_out[14][1] ), .X(n7207) );
  inv_x2_sg U9706 ( .A(\update_mask_0/reg_out[14][6] ), .X(n7209) );
  inv_x2_sg U9707 ( .A(\update_mask_0/reg_out[14][11] ), .X(n7211) );
  inv_x2_sg U9708 ( .A(\update_mask_0/reg_out[0][4] ), .X(n7213) );
  inv_x2_sg U9709 ( .A(\update_mask_0/reg_out[0][9] ), .X(n7215) );
  inv_x2_sg U9710 ( .A(\update_mask_0/reg_out[0][14] ), .X(n7217) );
  inv_x2_sg U9711 ( .A(\update_mask_0/reg_out[1][4] ), .X(n7219) );
  inv_x2_sg U9712 ( .A(\update_mask_0/reg_out[1][9] ), .X(n7221) );
  inv_x2_sg U9713 ( .A(\update_mask_0/reg_out[1][14] ), .X(n7223) );
  inv_x2_sg U9714 ( .A(\update_mask_0/reg_out[2][4] ), .X(n7225) );
  inv_x2_sg U9715 ( .A(\update_mask_0/reg_out[2][9] ), .X(n7227) );
  inv_x2_sg U9716 ( .A(\update_mask_0/reg_out[2][14] ), .X(n7229) );
  inv_x2_sg U9717 ( .A(\update_mask_0/reg_out[3][4] ), .X(n7231) );
  inv_x2_sg U9718 ( .A(\update_mask_0/reg_out[3][9] ), .X(n7233) );
  inv_x2_sg U9719 ( .A(\update_mask_0/reg_out[3][14] ), .X(n7235) );
  inv_x2_sg U9720 ( .A(\update_mask_0/reg_out[6][4] ), .X(n7237) );
  inv_x2_sg U9721 ( .A(\update_mask_0/reg_out[6][9] ), .X(n7239) );
  inv_x2_sg U9722 ( .A(\update_mask_0/reg_out[6][14] ), .X(n7241) );
  inv_x2_sg U9723 ( .A(\update_mask_0/reg_out[6][18] ), .X(n7243) );
  inv_x2_sg U9724 ( .A(\update_mask_0/reg_out[7][4] ), .X(n7245) );
  inv_x2_sg U9725 ( .A(\update_mask_0/reg_out[7][9] ), .X(n7247) );
  inv_x2_sg U9726 ( .A(\update_mask_0/reg_out[7][14] ), .X(n7249) );
  inv_x2_sg U9727 ( .A(\update_mask_0/reg_out[7][18] ), .X(n7251) );
  inv_x2_sg U9728 ( .A(\update_mask_0/reg_out[10][4] ), .X(n7253) );
  inv_x2_sg U9729 ( .A(\update_mask_0/reg_out[10][9] ), .X(n7255) );
  inv_x2_sg U9730 ( .A(\update_mask_0/reg_out[10][14] ), .X(n7257) );
  inv_x2_sg U9731 ( .A(\update_mask_0/reg_out[12][4] ), .X(n7259) );
  inv_x2_sg U9732 ( .A(\update_mask_0/reg_out[12][9] ), .X(n7261) );
  inv_x2_sg U9733 ( .A(\update_mask_0/reg_out[12][14] ), .X(n7263) );
  inv_x2_sg U9734 ( .A(\update_mask_0/reg_out[14][18] ), .X(n7265) );
  inv_x2_sg U9735 ( .A(n9568), .X(n7305) );
  inv_x2_sg U9736 ( .A(\update_mask_0/reg_i_mask [2]), .X(n6339) );
  inv_x2_sg U9737 ( .A(\update_mask_0/reg_out[0][19] ), .X(n7271) );
  inv_x2_sg U9738 ( .A(\update_mask_0/N27 ), .X(n6153) );
  inv_x2_sg U9739 ( .A(\update_output_0/N33 ), .X(n6155) );
  nor_x2_sg U9740 ( .A(n7160), .B(n9219), .X(n2066) );
  nor_x4_sg U9741 ( .A(n7526), .B(n9222), .X(n3849) );
  inv_x4_sg U9742 ( .A(n5153), .X(n9222) );
  nor_x4_sg U9743 ( .A(n7526), .B(n9234), .X(n3873) );
  inv_x4_sg U9744 ( .A(n4629), .X(n9234) );
  nor_x4_sg U9745 ( .A(n7526), .B(n9237), .X(n3885) );
  inv_x4_sg U9746 ( .A(n4503), .X(n9237) );
  inv_x2_sg U9747 ( .A(n6041), .X(n6042) );
  inv_x2_sg U9748 ( .A(n6043), .X(n6044) );
  inv_x2_sg U9749 ( .A(n6045), .X(n6046) );
  inv_x4_sg U9750 ( .A(n6047), .X(n6048) );
  inv_x8_sg U9751 ( .A(n9066), .X(n6377) );
  inv_x4_sg U9752 ( .A(n6051), .X(n6052) );
  inv_x4_sg U9753 ( .A(n6053), .X(n6054) );
  inv_x4_sg U9754 ( .A(n6055), .X(n6056) );
  inv_x4_sg U9755 ( .A(n6057), .X(n6058) );
  inv_x4_sg U9756 ( .A(n6059), .X(n6060) );
  inv_x4_sg U9757 ( .A(n6061), .X(n6062) );
  inv_x4_sg U9758 ( .A(n6063), .X(n6064) );
  inv_x4_sg U9759 ( .A(n6065), .X(n6066) );
  inv_x4_sg U9760 ( .A(n6067), .X(n6068) );
  inv_x4_sg U9761 ( .A(n6069), .X(n6070) );
  inv_x4_sg U9762 ( .A(n6071), .X(n6072) );
  inv_x4_sg U9763 ( .A(n6073), .X(n6074) );
  inv_x4_sg U9764 ( .A(n6075), .X(n6076) );
  inv_x4_sg U9765 ( .A(n6077), .X(n6078) );
  inv_x4_sg U9766 ( .A(n6079), .X(n6080) );
  inv_x4_sg U9767 ( .A(n6081), .X(n6082) );
  inv_x4_sg U9768 ( .A(n6083), .X(n6084) );
  inv_x4_sg U9769 ( .A(n6085), .X(n6086) );
  inv_x4_sg U9770 ( .A(n6087), .X(n6088) );
  inv_x4_sg U9771 ( .A(n6089), .X(n6090) );
  inv_x4_sg U9772 ( .A(n6091), .X(n6092) );
  inv_x4_sg U9773 ( .A(n6093), .X(n6094) );
  inv_x4_sg U9774 ( .A(n6095), .X(n6096) );
  inv_x4_sg U9775 ( .A(n6097), .X(n6098) );
  inv_x4_sg U9776 ( .A(n6099), .X(n6100) );
  inv_x4_sg U9777 ( .A(n6101), .X(n6102) );
  inv_x4_sg U9778 ( .A(n6103), .X(n6104) );
  inv_x4_sg U9779 ( .A(n6105), .X(n6106) );
  inv_x4_sg U9780 ( .A(n6107), .X(n6108) );
  inv_x4_sg U9781 ( .A(n6109), .X(n6110) );
  inv_x4_sg U9782 ( .A(n6111), .X(n6112) );
  inv_x4_sg U9783 ( .A(n6113), .X(n6114) );
  inv_x4_sg U9784 ( .A(n6115), .X(n6116) );
  inv_x4_sg U9785 ( .A(n6117), .X(n6118) );
  inv_x4_sg U9786 ( .A(n6119), .X(n6120) );
  inv_x4_sg U9787 ( .A(n6121), .X(n6122) );
  inv_x4_sg U9788 ( .A(n6123), .X(n6124) );
  inv_x4_sg U9789 ( .A(n6125), .X(n6126) );
  inv_x4_sg U9790 ( .A(n6127), .X(n6128) );
  inv_x4_sg U9791 ( .A(n6129), .X(n6130) );
  inv_x4_sg U9792 ( .A(n6131), .X(n6132) );
  inv_x4_sg U9793 ( .A(n6133), .X(n6134) );
  inv_x4_sg U9794 ( .A(n6135), .X(n6136) );
  inv_x4_sg U9795 ( .A(n6137), .X(n6138) );
  inv_x4_sg U9796 ( .A(n6139), .X(n6140) );
  inv_x4_sg U9797 ( .A(n6141), .X(n6142) );
  inv_x4_sg U9798 ( .A(n6143), .X(n6144) );
  inv_x4_sg U9799 ( .A(n6145), .X(n6146) );
  inv_x4_sg U9800 ( .A(n6147), .X(n6148) );
  inv_x4_sg U9801 ( .A(n6149), .X(n6150) );
  nor_x4_sg U9802 ( .A(n7522), .B(n6383), .X(n2038) );
  inv_x4_sg U9803 ( .A(n5901), .X(n6151) );
  nor_x4_sg U9804 ( .A(n9066), .B(n9213), .X(n1838) );
  nor_x8_sg U9805 ( .A(n826), .B(n7318), .X(n837) );
  nor_x8_sg U9806 ( .A(n5236), .B(n7559), .X(n7423) );
  nor_x8_sg U9807 ( .A(n7563), .B(n7564), .X(n1510) );
  inv_x8_sg U9808 ( .A(n1845), .X(n9074) );
  nand_x8_sg U9809 ( .A(n7310), .B(n1839), .X(n1845) );
  inv_x8_sg U9810 ( .A(n5274), .X(n9203) );
  inv_x8_sg U9811 ( .A(n1872), .X(n9075) );
  nor_x2_sg U9812 ( .A(n8990), .B(n7559), .X(n814) );
  inv_x8_sg U9813 ( .A(n797), .X(n8990) );
  inv_x2_sg U9814 ( .A(\update_mask_0/reg_out[2][15] ), .X(n7067) );
  inv_x2_sg U9815 ( .A(\update_mask_0/reg_out[3][15] ), .X(n7071) );
  inv_x2_sg U9816 ( .A(\update_mask_0/reg_out[5][15] ), .X(n7091) );
  inv_x2_sg U9817 ( .A(\update_mask_0/reg_out[6][15] ), .X(n7101) );
  inv_x2_sg U9818 ( .A(\update_mask_0/reg_out[6][16] ), .X(n7103) );
  inv_x2_sg U9819 ( .A(\update_mask_0/reg_out[8][15] ), .X(n7113) );
  inv_x2_sg U9820 ( .A(\update_mask_0/reg_out[9][15] ), .X(n7121) );
  inv_x2_sg U9821 ( .A(\update_mask_0/reg_out[10][15] ), .X(n7129) );
  inv_x2_sg U9822 ( .A(\update_mask_0/reg_out[11][15] ), .X(n7137) );
  inv_x2_sg U9823 ( .A(\update_mask_0/reg_out[14][15] ), .X(n7147) );
  inv_x2_sg U9824 ( .A(\update_mask_0/reg_out[14][16] ), .X(n7149) );
  inv_x2_sg U9825 ( .A(\update_mask_0/reg_out[15][15] ), .X(n7157) );
  inv_x2_sg U9826 ( .A(\update_mask_0/reg_i_mask [1]), .X(n7159) );
  inv_x2_sg U9827 ( .A(\update_mask_0/reg_out[13][15] ), .X(n7205) );
  nor_x2_sg U9828 ( .A(output_taken), .B(n9211), .X(n5324) );
  nor_x2_sg U9829 ( .A(n5930), .B(n9210), .X(n5323) );
  nor_x4_sg U9830 ( .A(n7526), .B(n9232), .X(n3843) );
  inv_x4_sg U9831 ( .A(n4715), .X(n9232) );
  nor_x4_sg U9832 ( .A(n7526), .B(n9236), .X(n3837) );
  inv_x4_sg U9833 ( .A(n4545), .X(n9236) );
  nor_x4_sg U9834 ( .A(n7526), .B(n9220), .X(n3864) );
  inv_x4_sg U9835 ( .A(n5229), .X(n9220) );
  nor_x4_sg U9836 ( .A(n8988), .B(n7569), .X(n879) );
  nor_x4_sg U9837 ( .A(n4192), .B(n8989), .X(n4207) );
  inv_x8_sg U9838 ( .A(n1511), .X(n8989) );
  inv_x4_sg U9839 ( .A(n7320), .X(n9071) );
  inv_x4_sg U9840 ( .A(reset), .X(n9197) );
  inv_x4_sg U9841 ( .A(n6153), .X(n6154) );
  nor_x4_sg U9842 ( .A(n7321), .B(n7312), .X(n4445) );
  inv_x4_sg U9843 ( .A(n6155), .X(n6156) );
  inv_x4_sg U9844 ( .A(n6157), .X(n6158) );
  inv_x4_sg U9845 ( .A(n6159), .X(n6160) );
  inv_x4_sg U9846 ( .A(n6161), .X(n6162) );
  inv_x4_sg U9847 ( .A(n6163), .X(n6164) );
  inv_x4_sg U9848 ( .A(n6165), .X(n6166) );
  inv_x4_sg U9849 ( .A(n6167), .X(n6168) );
  inv_x4_sg U9850 ( .A(n6169), .X(n6170) );
  inv_x4_sg U9851 ( .A(n6171), .X(n6172) );
  inv_x4_sg U9852 ( .A(n6173), .X(n6174) );
  inv_x4_sg U9853 ( .A(n6175), .X(n6176) );
  inv_x4_sg U9854 ( .A(n6177), .X(n6178) );
  inv_x4_sg U9855 ( .A(n6179), .X(n6180) );
  inv_x4_sg U9856 ( .A(n6181), .X(n6182) );
  inv_x4_sg U9857 ( .A(n6183), .X(n6184) );
  inv_x4_sg U9858 ( .A(n6185), .X(n6186) );
  inv_x4_sg U9859 ( .A(n6187), .X(n6188) );
  inv_x4_sg U9860 ( .A(n6189), .X(n6190) );
  inv_x4_sg U9861 ( .A(n6191), .X(n6192) );
  inv_x4_sg U9862 ( .A(n6193), .X(n6194) );
  inv_x4_sg U9863 ( .A(n6195), .X(n6196) );
  inv_x4_sg U9864 ( .A(n6197), .X(n6198) );
  inv_x4_sg U9865 ( .A(n6199), .X(n6200) );
  inv_x4_sg U9866 ( .A(n6201), .X(n6202) );
  inv_x4_sg U9867 ( .A(n6203), .X(n6204) );
  inv_x4_sg U9868 ( .A(n6205), .X(n6206) );
  inv_x4_sg U9869 ( .A(n6207), .X(n6208) );
  inv_x4_sg U9870 ( .A(n6209), .X(n6210) );
  inv_x4_sg U9871 ( .A(n6211), .X(n6212) );
  inv_x4_sg U9872 ( .A(n6213), .X(n6214) );
  inv_x4_sg U9873 ( .A(n6215), .X(n6216) );
  inv_x4_sg U9874 ( .A(n6217), .X(n6218) );
  inv_x4_sg U9875 ( .A(n6219), .X(n6220) );
  inv_x4_sg U9876 ( .A(n6221), .X(n6222) );
  inv_x4_sg U9877 ( .A(n6223), .X(n6224) );
  inv_x4_sg U9878 ( .A(n6225), .X(n6226) );
  inv_x4_sg U9879 ( .A(n6227), .X(n6228) );
  inv_x4_sg U9880 ( .A(n6229), .X(n6230) );
  inv_x4_sg U9881 ( .A(n6231), .X(n6232) );
  inv_x4_sg U9882 ( .A(n6233), .X(n6234) );
  inv_x4_sg U9883 ( .A(n6235), .X(n6236) );
  inv_x4_sg U9884 ( .A(n6237), .X(n6238) );
  inv_x4_sg U9885 ( .A(n6239), .X(n6240) );
  inv_x4_sg U9886 ( .A(n6241), .X(n6242) );
  inv_x4_sg U9887 ( .A(n6243), .X(n6244) );
  inv_x4_sg U9888 ( .A(n6245), .X(n6246) );
  inv_x4_sg U9889 ( .A(n6247), .X(n6248) );
  inv_x4_sg U9890 ( .A(n6249), .X(n6250) );
  inv_x4_sg U9891 ( .A(n6251), .X(n6252) );
  inv_x4_sg U9892 ( .A(n6253), .X(n6254) );
  inv_x4_sg U9893 ( .A(n6255), .X(n6256) );
  inv_x4_sg U9894 ( .A(n6257), .X(n6258) );
  inv_x4_sg U9895 ( .A(n6259), .X(n6260) );
  inv_x4_sg U9896 ( .A(n6261), .X(n6262) );
  inv_x4_sg U9897 ( .A(n6263), .X(n6264) );
  inv_x4_sg U9898 ( .A(n6265), .X(n6266) );
  inv_x4_sg U9899 ( .A(n6267), .X(n6268) );
  inv_x4_sg U9900 ( .A(n6269), .X(n6270) );
  inv_x4_sg U9901 ( .A(n6271), .X(n6272) );
  inv_x4_sg U9902 ( .A(n6273), .X(n6274) );
  inv_x4_sg U9903 ( .A(n6275), .X(n6276) );
  inv_x4_sg U9904 ( .A(n6277), .X(n6278) );
  inv_x4_sg U9905 ( .A(n6279), .X(n6280) );
  inv_x4_sg U9906 ( .A(n6281), .X(n6282) );
  inv_x4_sg U9907 ( .A(n6283), .X(n6284) );
  inv_x4_sg U9908 ( .A(n6285), .X(n6286) );
  inv_x4_sg U9909 ( .A(n6287), .X(n6288) );
  inv_x4_sg U9910 ( .A(n6289), .X(n6290) );
  inv_x4_sg U9911 ( .A(n6291), .X(n6292) );
  inv_x4_sg U9912 ( .A(n6293), .X(n6294) );
  inv_x4_sg U9913 ( .A(n6295), .X(n6296) );
  inv_x4_sg U9914 ( .A(n6297), .X(n6298) );
  inv_x4_sg U9915 ( .A(n6299), .X(n6300) );
  inv_x4_sg U9916 ( .A(n6301), .X(n6302) );
  inv_x4_sg U9917 ( .A(n6303), .X(n6304) );
  inv_x4_sg U9918 ( .A(n6305), .X(n6306) );
  inv_x4_sg U9919 ( .A(n6307), .X(n6308) );
  inv_x4_sg U9920 ( .A(n6309), .X(n6310) );
  inv_x4_sg U9921 ( .A(n6311), .X(n6312) );
  inv_x4_sg U9922 ( .A(n6313), .X(n6314) );
  inv_x4_sg U9923 ( .A(n6315), .X(n6316) );
  inv_x4_sg U9924 ( .A(n6317), .X(n6318) );
  inv_x4_sg U9925 ( .A(n6319), .X(n6320) );
  inv_x4_sg U9926 ( .A(n6321), .X(n6322) );
  inv_x4_sg U9927 ( .A(n6323), .X(n6324) );
  inv_x4_sg U9928 ( .A(n6325), .X(n6326) );
  inv_x4_sg U9929 ( .A(n6327), .X(n6328) );
  inv_x4_sg U9930 ( .A(n6329), .X(n6330) );
  inv_x4_sg U9931 ( .A(n6331), .X(n6332) );
  inv_x4_sg U9932 ( .A(n6333), .X(n6334) );
  inv_x4_sg U9933 ( .A(n6335), .X(n6336) );
  inv_x4_sg U9934 ( .A(n6337), .X(n6338) );
  inv_x4_sg U9935 ( .A(n6339), .X(n6340) );
  inv_x4_sg U9936 ( .A(n6341), .X(n6342) );
  inv_x4_sg U9937 ( .A(n6343), .X(n6344) );
  inv_x4_sg U9938 ( .A(n6345), .X(n6346) );
  inv_x4_sg U9939 ( .A(n6347), .X(n6348) );
  inv_x4_sg U9940 ( .A(n6349), .X(n6350) );
  inv_x4_sg U9941 ( .A(n6351), .X(n6352) );
  inv_x4_sg U9942 ( .A(n6353), .X(n6354) );
  inv_x4_sg U9943 ( .A(n6355), .X(n6356) );
  inv_x4_sg U9944 ( .A(n6357), .X(n6358) );
  inv_x4_sg U9945 ( .A(n6359), .X(n6360) );
  inv_x4_sg U9946 ( .A(n6361), .X(n6362) );
  inv_x4_sg U9947 ( .A(n6363), .X(n6364) );
  inv_x4_sg U9948 ( .A(n6365), .X(n6366) );
  inv_x4_sg U9949 ( .A(n6367), .X(n6368) );
  inv_x4_sg U9950 ( .A(n6369), .X(n6370) );
  inv_x4_sg U9951 ( .A(n6371), .X(n6372) );
  inv_x4_sg U9952 ( .A(n6373), .X(n6374) );
  inv_x4_sg U9953 ( .A(n6375), .X(n6376) );
  nor_x4_sg U9954 ( .A(n9066), .B(n7308), .X(n1839) );
  nor_x8_sg U9955 ( .A(n4192), .B(n4184), .X(n7384) );
  inv_x8_sg U9956 ( .A(n838), .X(n9186) );
  nor_x8_sg U9957 ( .A(n7562), .B(n7564), .X(n1512) );
  inv_x4_sg U9958 ( .A(n6378), .X(n6379) );
  inv_x8_sg U9959 ( .A(n6379), .X(n9066) );
  inv_x4_sg U9960 ( .A(n5907), .X(n6380) );
  inv_x8_sg U9961 ( .A(n6380), .X(n6381) );
  inv_x4_sg U9962 ( .A(n1623), .X(n9068) );
  nor_x8_sg U9963 ( .A(n5286), .B(n9213), .X(n1623) );
  inv_x8_sg U9964 ( .A(n3814), .X(n9073) );
  inv_x8_sg U9965 ( .A(n1876), .X(n9076) );
  inv_x4_sg U9966 ( .A(n5917), .X(n6382) );
  inv_x8_sg U9967 ( .A(n6382), .X(n6383) );
  inv_x8_sg U9968 ( .A(n6383), .X(n9215) );
  nor_x2_sg U9969 ( .A(n9193), .B(n4301), .X(n4298) );
  inv_x4_sg U9970 ( .A(n4302), .X(n9193) );
  inv_x1_sg U9971 ( .A(n5299), .X(n9200) );
  nor_x4_sg U9972 ( .A(n7526), .B(n9233), .X(n3852) );
  inv_x4_sg U9973 ( .A(n4673), .X(n9233) );
  nand_x4_sg U9974 ( .A(n9197), .B(n5312), .X(n3823) );
  inv_x4_sg U9975 ( .A(n4197), .X(n9192) );
  nor_x4_sg U9976 ( .A(n3930), .B(n4182), .X(n4197) );
  inv_x2_sg U9977 ( .A(n6384), .X(\o_im[13][19] ) );
  inv_x2_sg U9978 ( .A(n6386), .X(\o_im[13][18] ) );
  inv_x2_sg U9979 ( .A(n6388), .X(\o_im[13][17] ) );
  inv_x2_sg U9980 ( .A(n6390), .X(\o_im[13][16] ) );
  inv_x2_sg U9981 ( .A(n6392), .X(\o_im[13][15] ) );
  inv_x2_sg U9982 ( .A(n6394), .X(\o_im[13][14] ) );
  inv_x2_sg U9983 ( .A(n6396), .X(\o_im[13][13] ) );
  inv_x2_sg U9984 ( .A(n6398), .X(\o_im[13][12] ) );
  inv_x2_sg U9985 ( .A(n6400), .X(\o_im[13][11] ) );
  inv_x2_sg U9986 ( .A(n6402), .X(\o_im[13][10] ) );
  inv_x2_sg U9987 ( .A(n6404), .X(\o_im[13][9] ) );
  inv_x2_sg U9988 ( .A(n6406), .X(\o_im[13][8] ) );
  inv_x2_sg U9989 ( .A(n6408), .X(\o_im[13][7] ) );
  inv_x2_sg U9990 ( .A(n6410), .X(\o_im[13][6] ) );
  inv_x2_sg U9991 ( .A(n6412), .X(\o_im[13][5] ) );
  inv_x2_sg U9992 ( .A(n6414), .X(\o_im[13][4] ) );
  inv_x2_sg U9993 ( .A(n6416), .X(\o_im[13][3] ) );
  inv_x2_sg U9994 ( .A(n6418), .X(\o_im[13][2] ) );
  inv_x2_sg U9995 ( .A(n6420), .X(\o_im[13][1] ) );
  inv_x2_sg U9996 ( .A(n6422), .X(\o_im[13][0] ) );
  inv_x2_sg U9997 ( .A(n6424), .X(\o_im[5][19] ) );
  inv_x2_sg U9998 ( .A(n6426), .X(\o_im[5][18] ) );
  inv_x2_sg U9999 ( .A(n6428), .X(\o_im[5][17] ) );
  inv_x2_sg U10000 ( .A(n6430), .X(\o_im[5][16] ) );
  inv_x2_sg U10001 ( .A(n6432), .X(\o_im[5][15] ) );
  inv_x2_sg U10002 ( .A(n6434), .X(\o_im[5][14] ) );
  inv_x2_sg U10003 ( .A(n6436), .X(\o_im[5][13] ) );
  inv_x2_sg U10004 ( .A(n6438), .X(\o_im[5][12] ) );
  inv_x2_sg U10005 ( .A(n6440), .X(\o_im[5][11] ) );
  inv_x2_sg U10006 ( .A(n6442), .X(\o_im[5][10] ) );
  inv_x2_sg U10007 ( .A(n6444), .X(\o_im[5][9] ) );
  inv_x2_sg U10008 ( .A(n6446), .X(\o_im[5][8] ) );
  inv_x2_sg U10009 ( .A(n6448), .X(\o_im[5][7] ) );
  inv_x2_sg U10010 ( .A(n6450), .X(\o_im[5][6] ) );
  inv_x2_sg U10011 ( .A(n6452), .X(\o_im[5][5] ) );
  inv_x2_sg U10012 ( .A(n6454), .X(\o_im[5][4] ) );
  inv_x2_sg U10013 ( .A(n6456), .X(\o_im[5][3] ) );
  inv_x2_sg U10014 ( .A(n6458), .X(\o_im[5][2] ) );
  inv_x2_sg U10015 ( .A(n6460), .X(\o_im[5][1] ) );
  inv_x2_sg U10016 ( .A(n6462), .X(\o_im[5][0] ) );
  inv_x2_sg U10017 ( .A(n6464), .X(\o_im[14][19] ) );
  inv_x2_sg U10018 ( .A(n6466), .X(\o_im[14][18] ) );
  inv_x2_sg U10019 ( .A(n6468), .X(\o_im[14][17] ) );
  inv_x2_sg U10020 ( .A(n6470), .X(\o_im[14][16] ) );
  inv_x2_sg U10021 ( .A(n6472), .X(\o_im[14][15] ) );
  inv_x2_sg U10022 ( .A(n6474), .X(\o_im[14][14] ) );
  inv_x2_sg U10023 ( .A(n6476), .X(\o_im[14][13] ) );
  inv_x2_sg U10024 ( .A(n6478), .X(\o_im[14][12] ) );
  inv_x2_sg U10025 ( .A(n6480), .X(\o_im[14][11] ) );
  inv_x2_sg U10026 ( .A(n6482), .X(\o_im[14][10] ) );
  inv_x2_sg U10027 ( .A(n6484), .X(\o_im[14][9] ) );
  inv_x2_sg U10028 ( .A(n6486), .X(\o_im[14][8] ) );
  inv_x2_sg U10029 ( .A(n6488), .X(\o_im[14][7] ) );
  inv_x2_sg U10030 ( .A(n6490), .X(\o_im[14][6] ) );
  inv_x2_sg U10031 ( .A(n6492), .X(\o_im[14][5] ) );
  inv_x2_sg U10032 ( .A(n6494), .X(\o_im[14][4] ) );
  inv_x2_sg U10033 ( .A(n6496), .X(\o_im[14][3] ) );
  inv_x2_sg U10034 ( .A(n6498), .X(\o_im[14][2] ) );
  inv_x2_sg U10035 ( .A(n6500), .X(\o_im[14][1] ) );
  inv_x2_sg U10036 ( .A(n6502), .X(\o_im[14][0] ) );
  inv_x2_sg U10037 ( .A(n6504), .X(\o_im[6][19] ) );
  inv_x2_sg U10038 ( .A(n6506), .X(\o_im[6][18] ) );
  inv_x2_sg U10039 ( .A(n6508), .X(\o_im[6][17] ) );
  inv_x2_sg U10040 ( .A(n6510), .X(\o_im[6][16] ) );
  inv_x2_sg U10041 ( .A(n6512), .X(\o_im[6][15] ) );
  inv_x2_sg U10042 ( .A(n6514), .X(\o_im[6][14] ) );
  inv_x2_sg U10043 ( .A(n6516), .X(\o_im[6][13] ) );
  inv_x2_sg U10044 ( .A(n6518), .X(\o_im[6][12] ) );
  inv_x2_sg U10045 ( .A(n6520), .X(\o_im[6][11] ) );
  inv_x2_sg U10046 ( .A(n6522), .X(\o_im[6][10] ) );
  inv_x2_sg U10047 ( .A(n6524), .X(\o_im[6][9] ) );
  inv_x2_sg U10048 ( .A(n6526), .X(\o_im[6][8] ) );
  inv_x2_sg U10049 ( .A(n6528), .X(\o_im[6][7] ) );
  inv_x2_sg U10050 ( .A(n6530), .X(\o_im[6][6] ) );
  inv_x2_sg U10051 ( .A(n6532), .X(\o_im[6][5] ) );
  inv_x2_sg U10052 ( .A(n6534), .X(\o_im[6][4] ) );
  inv_x2_sg U10053 ( .A(n6536), .X(\o_im[6][3] ) );
  inv_x2_sg U10054 ( .A(n6538), .X(\o_im[6][2] ) );
  inv_x2_sg U10055 ( .A(n6540), .X(\o_im[6][1] ) );
  inv_x2_sg U10056 ( .A(n6542), .X(\o_im[6][0] ) );
  inv_x2_sg U10057 ( .A(n6544), .X(\o_im[4][19] ) );
  inv_x2_sg U10058 ( .A(n6546), .X(\o_im[4][18] ) );
  inv_x2_sg U10059 ( .A(n6548), .X(\o_im[4][17] ) );
  inv_x2_sg U10060 ( .A(n6550), .X(\o_im[4][16] ) );
  inv_x2_sg U10061 ( .A(n6552), .X(\o_im[4][15] ) );
  inv_x2_sg U10062 ( .A(n6554), .X(\o_im[4][14] ) );
  inv_x2_sg U10063 ( .A(n6556), .X(\o_im[4][13] ) );
  inv_x2_sg U10064 ( .A(n6558), .X(\o_im[4][12] ) );
  inv_x2_sg U10065 ( .A(n6560), .X(\o_im[4][11] ) );
  inv_x2_sg U10066 ( .A(n6562), .X(\o_im[4][10] ) );
  inv_x2_sg U10067 ( .A(n6564), .X(\o_im[4][9] ) );
  inv_x2_sg U10068 ( .A(n6566), .X(\o_im[4][8] ) );
  inv_x2_sg U10069 ( .A(n6568), .X(\o_im[4][7] ) );
  inv_x2_sg U10070 ( .A(n6570), .X(\o_im[4][6] ) );
  inv_x2_sg U10071 ( .A(n6572), .X(\o_im[4][5] ) );
  inv_x2_sg U10072 ( .A(n6574), .X(\o_im[4][4] ) );
  inv_x2_sg U10073 ( .A(n6576), .X(\o_im[4][3] ) );
  inv_x2_sg U10074 ( .A(n6578), .X(\o_im[4][2] ) );
  inv_x2_sg U10075 ( .A(n6580), .X(\o_im[4][1] ) );
  inv_x2_sg U10076 ( .A(n6582), .X(\o_im[4][0] ) );
  inv_x2_sg U10077 ( .A(n6584), .X(\o_im[12][19] ) );
  inv_x2_sg U10078 ( .A(n6586), .X(\o_im[12][18] ) );
  inv_x2_sg U10079 ( .A(n6588), .X(\o_im[12][17] ) );
  inv_x2_sg U10080 ( .A(n6590), .X(\o_im[12][16] ) );
  inv_x2_sg U10081 ( .A(n6592), .X(\o_im[12][15] ) );
  inv_x2_sg U10082 ( .A(n6594), .X(\o_im[12][14] ) );
  inv_x2_sg U10083 ( .A(n6596), .X(\o_im[12][13] ) );
  inv_x2_sg U10084 ( .A(n6598), .X(\o_im[12][12] ) );
  inv_x2_sg U10085 ( .A(n6600), .X(\o_im[12][11] ) );
  inv_x2_sg U10086 ( .A(n6602), .X(\o_im[12][10] ) );
  inv_x2_sg U10087 ( .A(n6604), .X(\o_im[12][9] ) );
  inv_x2_sg U10088 ( .A(n6606), .X(\o_im[12][8] ) );
  inv_x2_sg U10089 ( .A(n6608), .X(\o_im[12][7] ) );
  inv_x2_sg U10090 ( .A(n6610), .X(\o_im[12][6] ) );
  inv_x2_sg U10091 ( .A(n6612), .X(\o_im[12][5] ) );
  inv_x2_sg U10092 ( .A(n6614), .X(\o_im[12][4] ) );
  inv_x2_sg U10093 ( .A(n6616), .X(\o_im[12][3] ) );
  inv_x2_sg U10094 ( .A(n6618), .X(\o_im[12][2] ) );
  inv_x2_sg U10095 ( .A(n6620), .X(\o_im[12][1] ) );
  inv_x2_sg U10096 ( .A(n6622), .X(\o_im[12][0] ) );
  inv_x2_sg U10097 ( .A(n6624), .X(\o_im[3][19] ) );
  inv_x2_sg U10098 ( .A(n6626), .X(\o_im[3][18] ) );
  inv_x2_sg U10099 ( .A(n6628), .X(\o_im[3][17] ) );
  inv_x2_sg U10100 ( .A(n6630), .X(\o_im[3][16] ) );
  inv_x2_sg U10101 ( .A(n6632), .X(\o_im[3][15] ) );
  inv_x2_sg U10102 ( .A(n6634), .X(\o_im[3][14] ) );
  inv_x2_sg U10103 ( .A(n6636), .X(\o_im[3][13] ) );
  inv_x2_sg U10104 ( .A(n6638), .X(\o_im[3][12] ) );
  inv_x2_sg U10105 ( .A(n6640), .X(\o_im[3][11] ) );
  inv_x2_sg U10106 ( .A(n6642), .X(\o_im[3][10] ) );
  inv_x2_sg U10107 ( .A(n6644), .X(\o_im[3][9] ) );
  inv_x2_sg U10108 ( .A(n6646), .X(\o_im[3][8] ) );
  inv_x2_sg U10109 ( .A(n6648), .X(\o_im[3][7] ) );
  inv_x2_sg U10110 ( .A(n6650), .X(\o_im[3][6] ) );
  inv_x2_sg U10111 ( .A(n6652), .X(\o_im[3][5] ) );
  inv_x2_sg U10112 ( .A(n6654), .X(\o_im[3][4] ) );
  inv_x2_sg U10113 ( .A(n6656), .X(\o_im[3][3] ) );
  inv_x2_sg U10114 ( .A(n6658), .X(\o_im[3][2] ) );
  inv_x2_sg U10115 ( .A(n6660), .X(\o_im[3][1] ) );
  inv_x2_sg U10116 ( .A(n6662), .X(\o_im[3][0] ) );
  inv_x2_sg U10117 ( .A(n6664), .X(\o_im[11][19] ) );
  inv_x2_sg U10118 ( .A(n6666), .X(\o_im[11][18] ) );
  inv_x2_sg U10119 ( .A(n6668), .X(\o_im[11][17] ) );
  inv_x2_sg U10120 ( .A(n6670), .X(\o_im[11][16] ) );
  inv_x2_sg U10121 ( .A(n6672), .X(\o_im[11][15] ) );
  inv_x2_sg U10122 ( .A(n6674), .X(\o_im[11][14] ) );
  inv_x2_sg U10123 ( .A(n6676), .X(\o_im[11][13] ) );
  inv_x2_sg U10124 ( .A(n6678), .X(\o_im[11][12] ) );
  inv_x2_sg U10125 ( .A(n6680), .X(\o_im[11][11] ) );
  inv_x2_sg U10126 ( .A(n6682), .X(\o_im[11][10] ) );
  inv_x2_sg U10127 ( .A(n6684), .X(\o_im[11][9] ) );
  inv_x2_sg U10128 ( .A(n6686), .X(\o_im[11][8] ) );
  inv_x2_sg U10129 ( .A(n6688), .X(\o_im[11][7] ) );
  inv_x2_sg U10130 ( .A(n6690), .X(\o_im[11][6] ) );
  inv_x2_sg U10131 ( .A(n6692), .X(\o_im[11][5] ) );
  inv_x2_sg U10132 ( .A(n6694), .X(\o_im[11][4] ) );
  inv_x2_sg U10133 ( .A(n6696), .X(\o_im[11][3] ) );
  inv_x2_sg U10134 ( .A(n6698), .X(\o_im[11][2] ) );
  inv_x2_sg U10135 ( .A(n6700), .X(\o_im[11][1] ) );
  inv_x2_sg U10136 ( .A(n6702), .X(\o_im[11][0] ) );
  inv_x2_sg U10137 ( .A(n6704), .X(\o_im[9][19] ) );
  inv_x2_sg U10138 ( .A(n6706), .X(\o_im[9][18] ) );
  inv_x2_sg U10139 ( .A(n6708), .X(\o_im[9][17] ) );
  inv_x2_sg U10140 ( .A(n6710), .X(\o_im[9][16] ) );
  inv_x2_sg U10141 ( .A(n6712), .X(\o_im[9][15] ) );
  inv_x2_sg U10142 ( .A(n6714), .X(\o_im[9][14] ) );
  inv_x2_sg U10143 ( .A(n6716), .X(\o_im[9][13] ) );
  inv_x2_sg U10144 ( .A(n6718), .X(\o_im[9][12] ) );
  inv_x2_sg U10145 ( .A(n6720), .X(\o_im[9][11] ) );
  inv_x2_sg U10146 ( .A(n6722), .X(\o_im[9][10] ) );
  inv_x2_sg U10147 ( .A(n6724), .X(\o_im[9][9] ) );
  inv_x2_sg U10148 ( .A(n6726), .X(\o_im[9][8] ) );
  inv_x2_sg U10149 ( .A(n6728), .X(\o_im[9][7] ) );
  inv_x2_sg U10150 ( .A(n6730), .X(\o_im[9][6] ) );
  inv_x2_sg U10151 ( .A(n6732), .X(\o_im[9][5] ) );
  inv_x2_sg U10152 ( .A(n6734), .X(\o_im[9][4] ) );
  inv_x2_sg U10153 ( .A(n6736), .X(\o_im[9][3] ) );
  inv_x2_sg U10154 ( .A(n6738), .X(\o_im[9][2] ) );
  inv_x2_sg U10155 ( .A(n6740), .X(\o_im[9][1] ) );
  inv_x2_sg U10156 ( .A(n6742), .X(\o_im[9][0] ) );
  inv_x2_sg U10157 ( .A(n6744), .X(\o_im[1][19] ) );
  inv_x2_sg U10158 ( .A(n6746), .X(\o_im[1][18] ) );
  inv_x2_sg U10159 ( .A(n6748), .X(\o_im[1][17] ) );
  inv_x2_sg U10160 ( .A(n6750), .X(\o_im[1][16] ) );
  inv_x2_sg U10161 ( .A(n6752), .X(\o_im[1][15] ) );
  inv_x2_sg U10162 ( .A(n6754), .X(\o_im[1][14] ) );
  inv_x2_sg U10163 ( .A(n6756), .X(\o_im[1][13] ) );
  inv_x2_sg U10164 ( .A(n6758), .X(\o_im[1][12] ) );
  inv_x2_sg U10165 ( .A(n6760), .X(\o_im[1][11] ) );
  inv_x2_sg U10166 ( .A(n6762), .X(\o_im[1][10] ) );
  inv_x2_sg U10167 ( .A(n6764), .X(\o_im[1][9] ) );
  inv_x2_sg U10168 ( .A(n6766), .X(\o_im[1][8] ) );
  inv_x2_sg U10169 ( .A(n6768), .X(\o_im[1][7] ) );
  inv_x2_sg U10170 ( .A(n6770), .X(\o_im[1][6] ) );
  inv_x2_sg U10171 ( .A(n6772), .X(\o_im[1][5] ) );
  inv_x2_sg U10172 ( .A(n6774), .X(\o_im[1][4] ) );
  inv_x2_sg U10173 ( .A(n6776), .X(\o_im[1][3] ) );
  inv_x2_sg U10174 ( .A(n6778), .X(\o_im[1][2] ) );
  inv_x2_sg U10175 ( .A(n6780), .X(\o_im[1][1] ) );
  inv_x2_sg U10176 ( .A(n6782), .X(\o_im[1][0] ) );
  inv_x2_sg U10177 ( .A(n6784), .X(\o_im[10][19] ) );
  inv_x2_sg U10178 ( .A(n6786), .X(\o_im[10][18] ) );
  inv_x2_sg U10179 ( .A(n6788), .X(\o_im[10][17] ) );
  inv_x2_sg U10180 ( .A(n6790), .X(\o_im[10][16] ) );
  inv_x2_sg U10181 ( .A(n6792), .X(\o_im[10][15] ) );
  inv_x2_sg U10182 ( .A(n6794), .X(\o_im[10][14] ) );
  inv_x2_sg U10183 ( .A(n6796), .X(\o_im[10][13] ) );
  inv_x2_sg U10184 ( .A(n6798), .X(\o_im[10][12] ) );
  inv_x2_sg U10185 ( .A(n6800), .X(\o_im[10][11] ) );
  inv_x2_sg U10186 ( .A(n6802), .X(\o_im[10][10] ) );
  inv_x2_sg U10187 ( .A(n6804), .X(\o_im[10][9] ) );
  inv_x2_sg U10188 ( .A(n6806), .X(\o_im[10][8] ) );
  inv_x2_sg U10189 ( .A(n6808), .X(\o_im[10][7] ) );
  inv_x2_sg U10190 ( .A(n6810), .X(\o_im[10][6] ) );
  inv_x2_sg U10191 ( .A(n6812), .X(\o_im[10][5] ) );
  inv_x2_sg U10192 ( .A(n6814), .X(\o_im[10][4] ) );
  inv_x2_sg U10193 ( .A(n6816), .X(\o_im[10][3] ) );
  inv_x2_sg U10194 ( .A(n6818), .X(\o_im[10][2] ) );
  inv_x2_sg U10195 ( .A(n6820), .X(\o_im[10][1] ) );
  inv_x2_sg U10196 ( .A(n6822), .X(\o_im[10][0] ) );
  inv_x2_sg U10197 ( .A(n6824), .X(\o_im[2][19] ) );
  inv_x2_sg U10198 ( .A(n6826), .X(\o_im[2][18] ) );
  inv_x2_sg U10199 ( .A(n6828), .X(\o_im[2][17] ) );
  inv_x2_sg U10200 ( .A(n6830), .X(\o_im[2][16] ) );
  inv_x2_sg U10201 ( .A(n6832), .X(\o_im[2][15] ) );
  inv_x2_sg U10202 ( .A(n6834), .X(\o_im[2][14] ) );
  inv_x2_sg U10203 ( .A(n6836), .X(\o_im[2][13] ) );
  inv_x2_sg U10204 ( .A(n6838), .X(\o_im[2][12] ) );
  inv_x2_sg U10205 ( .A(n6840), .X(\o_im[2][11] ) );
  inv_x2_sg U10206 ( .A(n6842), .X(\o_im[2][10] ) );
  inv_x2_sg U10207 ( .A(n6844), .X(\o_im[2][9] ) );
  inv_x2_sg U10208 ( .A(n6846), .X(\o_im[2][8] ) );
  inv_x2_sg U10209 ( .A(n6848), .X(\o_im[2][7] ) );
  inv_x2_sg U10210 ( .A(n6850), .X(\o_im[2][6] ) );
  inv_x2_sg U10211 ( .A(n6852), .X(\o_im[2][5] ) );
  inv_x2_sg U10212 ( .A(n6854), .X(\o_im[2][4] ) );
  inv_x2_sg U10213 ( .A(n6856), .X(\o_im[2][3] ) );
  inv_x2_sg U10214 ( .A(n6858), .X(\o_im[2][2] ) );
  inv_x2_sg U10215 ( .A(n6860), .X(\o_im[2][1] ) );
  inv_x2_sg U10216 ( .A(n6862), .X(\o_im[2][0] ) );
  inv_x2_sg U10217 ( .A(n6864), .X(\o_im[0][19] ) );
  inv_x2_sg U10218 ( .A(n6866), .X(\o_im[0][18] ) );
  inv_x2_sg U10219 ( .A(n6868), .X(\o_im[0][17] ) );
  inv_x2_sg U10220 ( .A(n6870), .X(\o_im[0][16] ) );
  inv_x2_sg U10221 ( .A(n6872), .X(\o_im[0][15] ) );
  inv_x2_sg U10222 ( .A(n6874), .X(\o_im[0][14] ) );
  inv_x2_sg U10223 ( .A(n6876), .X(\o_im[0][13] ) );
  inv_x2_sg U10224 ( .A(n6878), .X(\o_im[0][12] ) );
  inv_x2_sg U10225 ( .A(n6880), .X(\o_im[0][11] ) );
  inv_x2_sg U10226 ( .A(n6882), .X(\o_im[0][10] ) );
  inv_x2_sg U10227 ( .A(n6884), .X(\o_im[0][9] ) );
  inv_x2_sg U10228 ( .A(n6886), .X(\o_im[0][8] ) );
  inv_x2_sg U10229 ( .A(n6888), .X(\o_im[0][7] ) );
  inv_x2_sg U10230 ( .A(n6890), .X(\o_im[0][6] ) );
  inv_x2_sg U10231 ( .A(n6892), .X(\o_im[0][5] ) );
  inv_x2_sg U10232 ( .A(n6894), .X(\o_im[0][4] ) );
  inv_x2_sg U10233 ( .A(n6896), .X(\o_im[0][3] ) );
  inv_x2_sg U10234 ( .A(n6898), .X(\o_im[0][2] ) );
  inv_x2_sg U10235 ( .A(n6900), .X(\o_im[0][1] ) );
  inv_x2_sg U10236 ( .A(n6902), .X(\o_im[0][0] ) );
  inv_x2_sg U10237 ( .A(n6904), .X(\o_im[8][19] ) );
  inv_x2_sg U10238 ( .A(n6906), .X(\o_im[8][18] ) );
  inv_x2_sg U10239 ( .A(n6908), .X(\o_im[8][17] ) );
  inv_x2_sg U10240 ( .A(n6910), .X(\o_im[8][16] ) );
  inv_x2_sg U10241 ( .A(n6912), .X(\o_im[8][15] ) );
  inv_x2_sg U10242 ( .A(n6914), .X(\o_im[8][14] ) );
  inv_x2_sg U10243 ( .A(n6916), .X(\o_im[8][13] ) );
  inv_x2_sg U10244 ( .A(n6918), .X(\o_im[8][12] ) );
  inv_x2_sg U10245 ( .A(n6920), .X(\o_im[8][11] ) );
  inv_x2_sg U10246 ( .A(n6922), .X(\o_im[8][10] ) );
  inv_x2_sg U10247 ( .A(n6924), .X(\o_im[8][9] ) );
  inv_x2_sg U10248 ( .A(n6926), .X(\o_im[8][8] ) );
  inv_x2_sg U10249 ( .A(n6928), .X(\o_im[8][7] ) );
  inv_x2_sg U10250 ( .A(n6930), .X(\o_im[8][6] ) );
  inv_x2_sg U10251 ( .A(n6932), .X(\o_im[8][5] ) );
  inv_x2_sg U10252 ( .A(n6934), .X(\o_im[8][4] ) );
  inv_x2_sg U10253 ( .A(n6936), .X(\o_im[8][3] ) );
  inv_x2_sg U10254 ( .A(n6938), .X(\o_im[8][2] ) );
  inv_x2_sg U10255 ( .A(n6940), .X(\o_im[8][1] ) );
  inv_x2_sg U10256 ( .A(n6942), .X(\o_im[8][0] ) );
  inv_x2_sg U10257 ( .A(n6944), .X(\o_im[7][19] ) );
  inv_x2_sg U10258 ( .A(n6946), .X(\o_im[7][18] ) );
  inv_x2_sg U10259 ( .A(n6948), .X(\o_im[7][17] ) );
  inv_x2_sg U10260 ( .A(n6950), .X(\o_im[7][16] ) );
  inv_x2_sg U10261 ( .A(n6952), .X(\o_im[7][15] ) );
  inv_x2_sg U10262 ( .A(n6954), .X(\o_im[7][14] ) );
  inv_x2_sg U10263 ( .A(n6956), .X(\o_im[7][13] ) );
  inv_x2_sg U10264 ( .A(n6958), .X(\o_im[7][12] ) );
  inv_x2_sg U10265 ( .A(n6960), .X(\o_im[7][11] ) );
  inv_x2_sg U10266 ( .A(n6962), .X(\o_im[7][10] ) );
  inv_x2_sg U10267 ( .A(n6964), .X(\o_im[7][9] ) );
  inv_x2_sg U10268 ( .A(n6966), .X(\o_im[7][8] ) );
  inv_x2_sg U10269 ( .A(n6968), .X(\o_im[7][7] ) );
  inv_x2_sg U10270 ( .A(n6970), .X(\o_im[7][6] ) );
  inv_x2_sg U10271 ( .A(n6972), .X(\o_im[7][5] ) );
  inv_x2_sg U10272 ( .A(n6974), .X(\o_im[7][4] ) );
  inv_x2_sg U10273 ( .A(n6976), .X(\o_im[7][3] ) );
  inv_x2_sg U10274 ( .A(n6978), .X(\o_im[7][2] ) );
  inv_x2_sg U10275 ( .A(n6980), .X(\o_im[7][1] ) );
  inv_x2_sg U10276 ( .A(n6982), .X(\o_im[7][0] ) );
  inv_x2_sg U10277 ( .A(n6984), .X(\o_im[15][19] ) );
  inv_x2_sg U10278 ( .A(n6986), .X(\o_im[15][18] ) );
  inv_x2_sg U10279 ( .A(n6988), .X(\o_im[15][17] ) );
  inv_x2_sg U10280 ( .A(n6990), .X(\o_im[15][16] ) );
  inv_x2_sg U10281 ( .A(n6992), .X(\o_im[15][15] ) );
  inv_x2_sg U10282 ( .A(n6994), .X(\o_im[15][14] ) );
  inv_x2_sg U10283 ( .A(n6996), .X(\o_im[15][13] ) );
  inv_x2_sg U10284 ( .A(n6998), .X(\o_im[15][12] ) );
  inv_x2_sg U10285 ( .A(n7000), .X(\o_im[15][11] ) );
  inv_x2_sg U10286 ( .A(n7002), .X(\o_im[15][10] ) );
  inv_x2_sg U10287 ( .A(n7004), .X(\o_im[15][9] ) );
  inv_x2_sg U10288 ( .A(n7006), .X(\o_im[15][8] ) );
  inv_x2_sg U10289 ( .A(n7008), .X(\o_im[15][7] ) );
  inv_x2_sg U10290 ( .A(n7010), .X(\o_im[15][6] ) );
  inv_x2_sg U10291 ( .A(n7012), .X(\o_im[15][5] ) );
  inv_x2_sg U10292 ( .A(n7014), .X(\o_im[15][4] ) );
  inv_x2_sg U10293 ( .A(n7016), .X(\o_im[15][3] ) );
  inv_x2_sg U10294 ( .A(n7018), .X(\o_im[15][2] ) );
  inv_x2_sg U10295 ( .A(n7020), .X(\o_im[15][1] ) );
  inv_x2_sg U10296 ( .A(n7022), .X(\o_im[15][0] ) );
  inv_x2_sg U10297 ( .A(n7024), .X(n7025) );
  inv_x2_sg U10298 ( .A(n7026), .X(n7027) );
  inv_x2_sg U10299 ( .A(n7028), .X(n7029) );
  inv_x2_sg U10300 ( .A(n7030), .X(n7031) );
  inv_x2_sg U10301 ( .A(n7032), .X(n7033) );
  inv_x2_sg U10302 ( .A(n7034), .X(n7035) );
  nand_x1_sg U10303 ( .A(n7035), .B(n7320), .X(n1686) );
  nor_x4_sg U10304 ( .A(n4297), .B(n9241), .X(n4451) );
  inv_x8_sg U10305 ( .A(n7323), .X(n9241) );
  nor_x4_sg U10306 ( .A(n4196), .B(n8989), .X(n862) );
  inv_x4_sg U10307 ( .A(n7038), .X(n7039) );
  inv_x4_sg U10308 ( .A(n7040), .X(state[0]) );
  inv_x4_sg U10309 ( .A(state[0]), .X(n9210) );
  inv_x4_sg U10310 ( .A(n7047), .X(n7048) );
  inv_x4_sg U10311 ( .A(n7049), .X(n7050) );
  inv_x4_sg U10312 ( .A(n7051), .X(n7052) );
  inv_x4_sg U10313 ( .A(n7053), .X(n7054) );
  inv_x4_sg U10314 ( .A(n7055), .X(n7056) );
  inv_x4_sg U10315 ( .A(n7057), .X(n7058) );
  inv_x4_sg U10316 ( .A(n7059), .X(n7060) );
  inv_x4_sg U10317 ( .A(n7061), .X(n7062) );
  inv_x4_sg U10318 ( .A(n7063), .X(n7064) );
  inv_x4_sg U10319 ( .A(n7065), .X(n7066) );
  inv_x4_sg U10320 ( .A(n7067), .X(n7068) );
  inv_x4_sg U10321 ( .A(n7069), .X(n7070) );
  inv_x4_sg U10322 ( .A(n7071), .X(n7072) );
  inv_x4_sg U10323 ( .A(n7073), .X(n7074) );
  inv_x4_sg U10324 ( .A(n7075), .X(n7076) );
  inv_x4_sg U10325 ( .A(n7077), .X(n7078) );
  inv_x4_sg U10326 ( .A(n7079), .X(n7080) );
  inv_x4_sg U10327 ( .A(n7081), .X(n7082) );
  inv_x4_sg U10328 ( .A(n7083), .X(n7084) );
  inv_x4_sg U10329 ( .A(n7085), .X(n7086) );
  inv_x4_sg U10330 ( .A(n7087), .X(n7088) );
  inv_x4_sg U10331 ( .A(n7089), .X(n7090) );
  inv_x4_sg U10332 ( .A(n7091), .X(n7092) );
  inv_x4_sg U10333 ( .A(n7093), .X(n7094) );
  inv_x4_sg U10334 ( .A(n7095), .X(n7096) );
  inv_x4_sg U10335 ( .A(n7097), .X(n7098) );
  inv_x4_sg U10336 ( .A(n7099), .X(n7100) );
  inv_x4_sg U10337 ( .A(n7101), .X(n7102) );
  inv_x4_sg U10338 ( .A(n7103), .X(n7104) );
  inv_x4_sg U10339 ( .A(n7105), .X(n7106) );
  inv_x4_sg U10340 ( .A(n7107), .X(n7108) );
  inv_x4_sg U10341 ( .A(n7109), .X(n7110) );
  inv_x4_sg U10342 ( .A(n7111), .X(n7112) );
  inv_x4_sg U10343 ( .A(n7113), .X(n7114) );
  inv_x4_sg U10344 ( .A(n7115), .X(n7116) );
  inv_x4_sg U10345 ( .A(n7117), .X(n7118) );
  inv_x4_sg U10346 ( .A(n7119), .X(n7120) );
  inv_x4_sg U10347 ( .A(n7121), .X(n7122) );
  inv_x4_sg U10348 ( .A(n7123), .X(n7124) );
  inv_x4_sg U10349 ( .A(n7125), .X(n7126) );
  inv_x4_sg U10350 ( .A(n7127), .X(n7128) );
  inv_x4_sg U10351 ( .A(n7129), .X(n7130) );
  inv_x4_sg U10352 ( .A(n7131), .X(n7132) );
  inv_x4_sg U10353 ( .A(n7133), .X(n7134) );
  inv_x4_sg U10354 ( .A(n7135), .X(n7136) );
  inv_x4_sg U10355 ( .A(n7137), .X(n7138) );
  inv_x4_sg U10356 ( .A(n7139), .X(n7140) );
  inv_x4_sg U10357 ( .A(n7141), .X(n7142) );
  inv_x4_sg U10358 ( .A(n7143), .X(n7144) );
  inv_x4_sg U10359 ( .A(n7145), .X(n7146) );
  inv_x4_sg U10360 ( .A(n7147), .X(n7148) );
  inv_x4_sg U10361 ( .A(n7149), .X(n7150) );
  inv_x4_sg U10362 ( .A(n7151), .X(n7152) );
  inv_x4_sg U10363 ( .A(n7153), .X(n7154) );
  inv_x4_sg U10364 ( .A(n7155), .X(n7156) );
  inv_x4_sg U10365 ( .A(n7157), .X(n7158) );
  inv_x4_sg U10366 ( .A(n7159), .X(n7160) );
  inv_x4_sg U10367 ( .A(n7161), .X(n7162) );
  inv_x4_sg U10368 ( .A(n7163), .X(n7164) );
  inv_x4_sg U10369 ( .A(n7165), .X(n7166) );
  inv_x4_sg U10370 ( .A(n7167), .X(n7168) );
  inv_x4_sg U10371 ( .A(n7169), .X(n7170) );
  inv_x4_sg U10372 ( .A(n7171), .X(n7172) );
  inv_x4_sg U10373 ( .A(n7173), .X(n7174) );
  inv_x4_sg U10374 ( .A(n7175), .X(n7176) );
  inv_x4_sg U10375 ( .A(n7177), .X(n7178) );
  inv_x4_sg U10376 ( .A(n7179), .X(n7180) );
  inv_x4_sg U10377 ( .A(n7181), .X(n7182) );
  inv_x4_sg U10378 ( .A(n7183), .X(n7184) );
  inv_x4_sg U10379 ( .A(n7185), .X(n7186) );
  inv_x4_sg U10380 ( .A(n7187), .X(n7188) );
  inv_x4_sg U10381 ( .A(n7189), .X(n7190) );
  inv_x4_sg U10382 ( .A(n7191), .X(n7192) );
  inv_x4_sg U10383 ( .A(n7193), .X(n7194) );
  inv_x4_sg U10384 ( .A(n7195), .X(n7196) );
  inv_x4_sg U10385 ( .A(n7197), .X(n7198) );
  inv_x4_sg U10386 ( .A(n7199), .X(n7200) );
  inv_x4_sg U10387 ( .A(n7201), .X(n7202) );
  inv_x4_sg U10388 ( .A(n7203), .X(n7204) );
  inv_x4_sg U10389 ( .A(n7205), .X(n7206) );
  inv_x4_sg U10390 ( .A(n7207), .X(n7208) );
  inv_x4_sg U10391 ( .A(n7209), .X(n7210) );
  inv_x4_sg U10392 ( .A(n7211), .X(n7212) );
  inv_x4_sg U10393 ( .A(n7213), .X(n7214) );
  inv_x4_sg U10394 ( .A(n7215), .X(n7216) );
  inv_x4_sg U10395 ( .A(n7217), .X(n7218) );
  inv_x4_sg U10396 ( .A(n7219), .X(n7220) );
  inv_x4_sg U10397 ( .A(n7221), .X(n7222) );
  inv_x4_sg U10398 ( .A(n7223), .X(n7224) );
  inv_x4_sg U10399 ( .A(n7225), .X(n7226) );
  inv_x4_sg U10400 ( .A(n7227), .X(n7228) );
  inv_x4_sg U10401 ( .A(n7229), .X(n7230) );
  inv_x4_sg U10402 ( .A(n7231), .X(n7232) );
  inv_x4_sg U10403 ( .A(n7233), .X(n7234) );
  inv_x4_sg U10404 ( .A(n7235), .X(n7236) );
  inv_x4_sg U10405 ( .A(n7237), .X(n7238) );
  inv_x4_sg U10406 ( .A(n7239), .X(n7240) );
  inv_x4_sg U10407 ( .A(n7241), .X(n7242) );
  inv_x4_sg U10408 ( .A(n7243), .X(n7244) );
  inv_x4_sg U10409 ( .A(n7245), .X(n7246) );
  inv_x4_sg U10410 ( .A(n7247), .X(n7248) );
  inv_x4_sg U10411 ( .A(n7249), .X(n7250) );
  inv_x4_sg U10412 ( .A(n7251), .X(n7252) );
  inv_x4_sg U10413 ( .A(n7253), .X(n7254) );
  inv_x4_sg U10414 ( .A(n7255), .X(n7256) );
  inv_x4_sg U10415 ( .A(n7257), .X(n7258) );
  inv_x4_sg U10416 ( .A(n7259), .X(n7260) );
  inv_x4_sg U10417 ( .A(n7261), .X(n7262) );
  inv_x4_sg U10418 ( .A(n7263), .X(n7264) );
  inv_x4_sg U10419 ( .A(n7265), .X(n7266) );
  inv_x4_sg U10420 ( .A(n7267), .X(n7268) );
  inv_x4_sg U10421 ( .A(n7269), .X(n7270) );
  inv_x4_sg U10422 ( .A(n7271), .X(n7272) );
  inv_x4_sg U10423 ( .A(n7273), .X(n7274) );
  inv_x4_sg U10424 ( .A(n7275), .X(n7276) );
  inv_x4_sg U10425 ( .A(n7277), .X(n7278) );
  inv_x4_sg U10426 ( .A(n7279), .X(n7280) );
  inv_x4_sg U10427 ( .A(n7281), .X(n7282) );
  inv_x4_sg U10428 ( .A(n7283), .X(n7284) );
  inv_x4_sg U10429 ( .A(n7285), .X(n7286) );
  inv_x4_sg U10430 ( .A(n7287), .X(n7288) );
  inv_x4_sg U10431 ( .A(n7289), .X(n7290) );
  inv_x4_sg U10432 ( .A(n7291), .X(n7292) );
  inv_x4_sg U10433 ( .A(n7293), .X(n7294) );
  inv_x4_sg U10434 ( .A(n7295), .X(n7296) );
  inv_x4_sg U10435 ( .A(n7297), .X(n7298) );
  inv_x4_sg U10436 ( .A(n7299), .X(n7300) );
  inv_x4_sg U10437 ( .A(n7301), .X(n7302) );
  inv_x4_sg U10438 ( .A(n7303), .X(n7304) );
  nor_x4_sg U10439 ( .A(n7526), .B(n7570), .X(n4017) );
  inv_x4_sg U10440 ( .A(n7305), .X(state[1]) );
  inv_x4_sg U10441 ( .A(state[1]), .X(n9211) );
  nor_x8_sg U10442 ( .A(n4192), .B(n4184), .X(n7385) );
  nor_x2_sg U10443 ( .A(n7519), .B(n841), .X(n844) );
  nor_x2_sg U10444 ( .A(n7519), .B(n838), .X(n843) );
  inv_x8_sg U10445 ( .A(n4393), .X(n9205) );
  nand_x8_sg U10446 ( .A(n6381), .B(n824), .X(n4393) );
  inv_x4_sg U10447 ( .A(n5919), .X(n7307) );
  inv_x8_sg U10448 ( .A(n7307), .X(n7308) );
  inv_x8_sg U10449 ( .A(n7308), .X(n9213) );
  inv_x8_sg U10450 ( .A(n1829), .X(n9212) );
  nand_x8_sg U10451 ( .A(n1838), .B(n9077), .X(n1829) );
  inv_x8_sg U10452 ( .A(n3929), .X(n9195) );
  nor_x4_sg U10453 ( .A(n3930), .B(n3931), .X(n3929) );
  nor_x4_sg U10454 ( .A(n3932), .B(n7526), .X(n3931) );
  inv_x8_sg U10455 ( .A(n5236), .X(n9240) );
  inv_x4_sg U10456 ( .A(n5921), .X(n7309) );
  inv_x8_sg U10457 ( .A(n7309), .X(n7310) );
  inv_x4_sg U10458 ( .A(n5903), .X(n7311) );
  inv_x8_sg U10459 ( .A(n7311), .X(n7312) );
  inv_x4_sg U10460 ( .A(n5923), .X(n7313) );
  inv_x8_sg U10461 ( .A(n7313), .X(n7314) );
  inv_x4_sg U10462 ( .A(n7314), .X(n9081) );
  inv_x4_sg U10463 ( .A(n5909), .X(n7315) );
  inv_x8_sg U10464 ( .A(n7315), .X(n7316) );
  inv_x8_sg U10465 ( .A(n7316), .X(n9219) );
  nor_x8_sg U10466 ( .A(n7398), .B(n7569), .X(n1511) );
  inv_x4_sg U10467 ( .A(n5915), .X(n7317) );
  inv_x8_sg U10468 ( .A(n7317), .X(n7318) );
  inv_x4_sg U10469 ( .A(n7318), .X(n9217) );
  nor_x1_sg U10470 ( .A(n7346), .B(n811), .X(\update_output_0/n2644 ) );
  nor_x1_sg U10471 ( .A(n7347), .B(n811), .X(\update_output_0/n2640 ) );
  nor_x1_sg U10472 ( .A(n7332), .B(n811), .X(\update_output_0/n2636 ) );
  nor_x1_sg U10473 ( .A(n7331), .B(n811), .X(\update_output_0/n2632 ) );
  nor_x1_sg U10474 ( .A(n7330), .B(n811), .X(\update_output_0/n2628 ) );
  nor_x1_sg U10475 ( .A(n7355), .B(n811), .X(\update_output_0/n2624 ) );
  nor_x1_sg U10476 ( .A(n7357), .B(n811), .X(\update_output_0/n2620 ) );
  nor_x1_sg U10477 ( .A(n7329), .B(n811), .X(\update_output_0/n2616 ) );
  nor_x1_sg U10478 ( .A(n7328), .B(n811), .X(\update_output_0/n2612 ) );
  nor_x1_sg U10479 ( .A(n7327), .B(n811), .X(\update_output_0/n2608 ) );
  nor_x1_sg U10480 ( .A(n7365), .B(n811), .X(\update_output_0/n2604 ) );
  nor_x1_sg U10481 ( .A(n7367), .B(n811), .X(\update_output_0/n2600 ) );
  nor_x1_sg U10482 ( .A(n7326), .B(n811), .X(\update_output_0/n2596 ) );
  nor_x1_sg U10483 ( .A(n7346), .B(n813), .X(\update_output_0/n2564 ) );
  nor_x1_sg U10484 ( .A(n7347), .B(n813), .X(\update_output_0/n2560 ) );
  nor_x1_sg U10485 ( .A(n7332), .B(n813), .X(\update_output_0/n2556 ) );
  nor_x1_sg U10486 ( .A(n7331), .B(n813), .X(\update_output_0/n2552 ) );
  nor_x1_sg U10487 ( .A(n7330), .B(n813), .X(\update_output_0/n2548 ) );
  nor_x1_sg U10488 ( .A(n7355), .B(n813), .X(\update_output_0/n2544 ) );
  nor_x1_sg U10489 ( .A(n7357), .B(n813), .X(\update_output_0/n2540 ) );
  nor_x1_sg U10490 ( .A(n7329), .B(n813), .X(\update_output_0/n2536 ) );
  nor_x1_sg U10491 ( .A(n7328), .B(n813), .X(\update_output_0/n2532 ) );
  nor_x1_sg U10492 ( .A(n7327), .B(n813), .X(\update_output_0/n2528 ) );
  nor_x1_sg U10493 ( .A(n7365), .B(n813), .X(\update_output_0/n2524 ) );
  nor_x1_sg U10494 ( .A(n7367), .B(n813), .X(\update_output_0/n2520 ) );
  nor_x1_sg U10495 ( .A(n7326), .B(n813), .X(\update_output_0/n2516 ) );
  nor_x1_sg U10496 ( .A(n7346), .B(n819), .X(\update_output_0/n2324 ) );
  nor_x1_sg U10497 ( .A(n7347), .B(n819), .X(\update_output_0/n2320 ) );
  nor_x1_sg U10498 ( .A(n7332), .B(n819), .X(\update_output_0/n2316 ) );
  nor_x1_sg U10499 ( .A(n7331), .B(n819), .X(\update_output_0/n2312 ) );
  nor_x1_sg U10500 ( .A(n7330), .B(n819), .X(\update_output_0/n2308 ) );
  nor_x1_sg U10501 ( .A(n7355), .B(n819), .X(\update_output_0/n2304 ) );
  nor_x1_sg U10502 ( .A(n7357), .B(n819), .X(\update_output_0/n2300 ) );
  nor_x1_sg U10503 ( .A(n7329), .B(n819), .X(\update_output_0/n2296 ) );
  nor_x1_sg U10504 ( .A(n7328), .B(n819), .X(\update_output_0/n2292 ) );
  nor_x1_sg U10505 ( .A(n7327), .B(n819), .X(\update_output_0/n2288 ) );
  nor_x1_sg U10506 ( .A(n7365), .B(n819), .X(\update_output_0/n2284 ) );
  nor_x1_sg U10507 ( .A(n7367), .B(n819), .X(\update_output_0/n2280 ) );
  nor_x1_sg U10508 ( .A(n7326), .B(n819), .X(\update_output_0/n2276 ) );
  nor_x1_sg U10509 ( .A(n7346), .B(n821), .X(\update_output_0/n2244 ) );
  nor_x1_sg U10510 ( .A(n7347), .B(n821), .X(\update_output_0/n2240 ) );
  nor_x1_sg U10511 ( .A(n7332), .B(n821), .X(\update_output_0/n2236 ) );
  nor_x1_sg U10512 ( .A(n7331), .B(n821), .X(\update_output_0/n2232 ) );
  nor_x1_sg U10513 ( .A(n7330), .B(n821), .X(\update_output_0/n2228 ) );
  nor_x1_sg U10514 ( .A(n7355), .B(n821), .X(\update_output_0/n2224 ) );
  nor_x1_sg U10515 ( .A(n7357), .B(n821), .X(\update_output_0/n2220 ) );
  nor_x1_sg U10516 ( .A(n7329), .B(n821), .X(\update_output_0/n2216 ) );
  nor_x1_sg U10517 ( .A(n7328), .B(n821), .X(\update_output_0/n2212 ) );
  nor_x1_sg U10518 ( .A(n7327), .B(n821), .X(\update_output_0/n2208 ) );
  nor_x1_sg U10519 ( .A(n7365), .B(n821), .X(\update_output_0/n2204 ) );
  nor_x1_sg U10520 ( .A(n7367), .B(n821), .X(\update_output_0/n2200 ) );
  nor_x1_sg U10521 ( .A(n7326), .B(n821), .X(\update_output_0/n2196 ) );
  nor_x1_sg U10522 ( .A(n7346), .B(n803), .X(\update_output_0/n3044 ) );
  nor_x1_sg U10523 ( .A(n7347), .B(n803), .X(\update_output_0/n3040 ) );
  nor_x1_sg U10524 ( .A(n7332), .B(n803), .X(\update_output_0/n3036 ) );
  nor_x1_sg U10525 ( .A(n7331), .B(n803), .X(\update_output_0/n3032 ) );
  nor_x1_sg U10526 ( .A(n7330), .B(n803), .X(\update_output_0/n3028 ) );
  nor_x1_sg U10527 ( .A(n7355), .B(n803), .X(\update_output_0/n3024 ) );
  nor_x1_sg U10528 ( .A(n7357), .B(n803), .X(\update_output_0/n3020 ) );
  nor_x1_sg U10529 ( .A(n7329), .B(n803), .X(\update_output_0/n3016 ) );
  nor_x1_sg U10530 ( .A(n7328), .B(n803), .X(\update_output_0/n3012 ) );
  nor_x1_sg U10531 ( .A(n7327), .B(n803), .X(\update_output_0/n3008 ) );
  nor_x1_sg U10532 ( .A(n7365), .B(n803), .X(\update_output_0/n3004 ) );
  nor_x1_sg U10533 ( .A(n7367), .B(n803), .X(\update_output_0/n3000 ) );
  nor_x1_sg U10534 ( .A(n7326), .B(n803), .X(\update_output_0/n2996 ) );
  nor_x1_sg U10535 ( .A(n7346), .B(n805), .X(\update_output_0/n2964 ) );
  nor_x1_sg U10536 ( .A(n7347), .B(n805), .X(\update_output_0/n2960 ) );
  nor_x1_sg U10537 ( .A(n7332), .B(n805), .X(\update_output_0/n2956 ) );
  nor_x1_sg U10538 ( .A(n7331), .B(n805), .X(\update_output_0/n2952 ) );
  nor_x1_sg U10539 ( .A(n7330), .B(n805), .X(\update_output_0/n2948 ) );
  nor_x1_sg U10540 ( .A(n7355), .B(n805), .X(\update_output_0/n2944 ) );
  nor_x1_sg U10541 ( .A(n7357), .B(n805), .X(\update_output_0/n2940 ) );
  nor_x1_sg U10542 ( .A(n7329), .B(n805), .X(\update_output_0/n2936 ) );
  nor_x1_sg U10543 ( .A(n7328), .B(n805), .X(\update_output_0/n2932 ) );
  nor_x1_sg U10544 ( .A(n7327), .B(n805), .X(\update_output_0/n2928 ) );
  nor_x1_sg U10545 ( .A(n7365), .B(n805), .X(\update_output_0/n2924 ) );
  nor_x1_sg U10546 ( .A(n7367), .B(n805), .X(\update_output_0/n2920 ) );
  nor_x1_sg U10547 ( .A(n7326), .B(n805), .X(\update_output_0/n2916 ) );
  nor_x1_sg U10548 ( .A(n7346), .B(n806), .X(\update_output_0/n2884 ) );
  nor_x1_sg U10549 ( .A(n7347), .B(n806), .X(\update_output_0/n2880 ) );
  nor_x1_sg U10550 ( .A(n7332), .B(n806), .X(\update_output_0/n2876 ) );
  nor_x1_sg U10551 ( .A(n7331), .B(n806), .X(\update_output_0/n2872 ) );
  nor_x1_sg U10552 ( .A(n7330), .B(n806), .X(\update_output_0/n2868 ) );
  nor_x1_sg U10553 ( .A(n7355), .B(n806), .X(\update_output_0/n2864 ) );
  nor_x1_sg U10554 ( .A(n7357), .B(n806), .X(\update_output_0/n2860 ) );
  nor_x1_sg U10555 ( .A(n7329), .B(n806), .X(\update_output_0/n2856 ) );
  nor_x1_sg U10556 ( .A(n7328), .B(n806), .X(\update_output_0/n2852 ) );
  nor_x1_sg U10557 ( .A(n7327), .B(n806), .X(\update_output_0/n2848 ) );
  nor_x1_sg U10558 ( .A(n7365), .B(n806), .X(\update_output_0/n2844 ) );
  nor_x1_sg U10559 ( .A(n7367), .B(n806), .X(\update_output_0/n2840 ) );
  nor_x1_sg U10560 ( .A(n7326), .B(n806), .X(\update_output_0/n2836 ) );
  nor_x1_sg U10561 ( .A(n7346), .B(n798), .X(\update_output_0/n3204 ) );
  nor_x1_sg U10562 ( .A(n7347), .B(n798), .X(\update_output_0/n3200 ) );
  nor_x1_sg U10563 ( .A(n7332), .B(n798), .X(\update_output_0/n3196 ) );
  nor_x1_sg U10564 ( .A(n7331), .B(n798), .X(\update_output_0/n3192 ) );
  nor_x1_sg U10565 ( .A(n7330), .B(n798), .X(\update_output_0/n3188 ) );
  nor_x1_sg U10566 ( .A(n7355), .B(n798), .X(\update_output_0/n3184 ) );
  nor_x1_sg U10567 ( .A(n7357), .B(n798), .X(\update_output_0/n3180 ) );
  nor_x1_sg U10568 ( .A(n7329), .B(n798), .X(\update_output_0/n3176 ) );
  nor_x1_sg U10569 ( .A(n7328), .B(n798), .X(\update_output_0/n3172 ) );
  nor_x1_sg U10570 ( .A(n7327), .B(n798), .X(\update_output_0/n3168 ) );
  nor_x1_sg U10571 ( .A(n7365), .B(n798), .X(\update_output_0/n3164 ) );
  nor_x1_sg U10572 ( .A(n7367), .B(n798), .X(\update_output_0/n3160 ) );
  nor_x1_sg U10573 ( .A(n7326), .B(n798), .X(\update_output_0/n3156 ) );
  nor_x1_sg U10574 ( .A(n7346), .B(n795), .X(\update_output_0/n3284 ) );
  nor_x1_sg U10575 ( .A(n7347), .B(n795), .X(\update_output_0/n3280 ) );
  nor_x1_sg U10576 ( .A(n7332), .B(n795), .X(\update_output_0/n3276 ) );
  nor_x1_sg U10577 ( .A(n7331), .B(n795), .X(\update_output_0/n3272 ) );
  nor_x1_sg U10578 ( .A(n7330), .B(n795), .X(\update_output_0/n3268 ) );
  nor_x1_sg U10579 ( .A(n7355), .B(n795), .X(\update_output_0/n3264 ) );
  nor_x1_sg U10580 ( .A(n7357), .B(n795), .X(\update_output_0/n3260 ) );
  nor_x1_sg U10581 ( .A(n7329), .B(n795), .X(\update_output_0/n3256 ) );
  nor_x1_sg U10582 ( .A(n7328), .B(n795), .X(\update_output_0/n3252 ) );
  nor_x1_sg U10583 ( .A(n7327), .B(n795), .X(\update_output_0/n3248 ) );
  nor_x1_sg U10584 ( .A(n7365), .B(n795), .X(\update_output_0/n3244 ) );
  nor_x1_sg U10585 ( .A(n7367), .B(n795), .X(\update_output_0/n3240 ) );
  nor_x1_sg U10586 ( .A(n7326), .B(n795), .X(\update_output_0/n3236 ) );
  nor_x1_sg U10587 ( .A(n7401), .B(n805), .X(\update_output_0/n2984 ) );
  nor_x1_sg U10588 ( .A(n7336), .B(n805), .X(\update_output_0/n2980 ) );
  nor_x1_sg U10589 ( .A(n7335), .B(n805), .X(\update_output_0/n2976 ) );
  nor_x1_sg U10590 ( .A(n7334), .B(n805), .X(\update_output_0/n2972 ) );
  nor_x1_sg U10591 ( .A(n7333), .B(n805), .X(\update_output_0/n2968 ) );
  nor_x1_sg U10592 ( .A(n7401), .B(n806), .X(\update_output_0/n2904 ) );
  nor_x1_sg U10593 ( .A(n7336), .B(n806), .X(\update_output_0/n2900 ) );
  nor_x1_sg U10594 ( .A(n7335), .B(n806), .X(\update_output_0/n2896 ) );
  nor_x1_sg U10595 ( .A(n7334), .B(n806), .X(\update_output_0/n2892 ) );
  nor_x1_sg U10596 ( .A(n7333), .B(n806), .X(\update_output_0/n2888 ) );
  nor_x1_sg U10597 ( .A(n7401), .B(n798), .X(\update_output_0/n3224 ) );
  nor_x1_sg U10598 ( .A(n7336), .B(n798), .X(\update_output_0/n3220 ) );
  nor_x1_sg U10599 ( .A(n7335), .B(n798), .X(\update_output_0/n3216 ) );
  nor_x1_sg U10600 ( .A(n7334), .B(n798), .X(\update_output_0/n3212 ) );
  nor_x1_sg U10601 ( .A(n7333), .B(n798), .X(\update_output_0/n3208 ) );
  nor_x1_sg U10602 ( .A(n7401), .B(n795), .X(\update_output_0/n3304 ) );
  nor_x1_sg U10603 ( .A(n7336), .B(n795), .X(\update_output_0/n3300 ) );
  nor_x1_sg U10604 ( .A(n7335), .B(n795), .X(\update_output_0/n3296 ) );
  nor_x1_sg U10605 ( .A(n7334), .B(n795), .X(\update_output_0/n3292 ) );
  nor_x1_sg U10606 ( .A(n7333), .B(n795), .X(\update_output_0/n3288 ) );
  nor_x1_sg U10607 ( .A(n7325), .B(n795), .X(\update_output_0/n3232 ) );
  nor_x1_sg U10608 ( .A(n7324), .B(n795), .X(\update_output_0/n3228 ) );
  nor_x1_sg U10609 ( .A(n7325), .B(n798), .X(\update_output_0/n3152 ) );
  nor_x1_sg U10610 ( .A(n7324), .B(n798), .X(\update_output_0/n3148 ) );
  nor_x1_sg U10611 ( .A(n7325), .B(n803), .X(\update_output_0/n2992 ) );
  nor_x1_sg U10612 ( .A(n7324), .B(n803), .X(\update_output_0/n2988 ) );
  nor_x1_sg U10613 ( .A(n7325), .B(n805), .X(\update_output_0/n2912 ) );
  nor_x1_sg U10614 ( .A(n7324), .B(n805), .X(\update_output_0/n2908 ) );
  nor_x1_sg U10615 ( .A(n7325), .B(n806), .X(\update_output_0/n2832 ) );
  nor_x1_sg U10616 ( .A(n7324), .B(n806), .X(\update_output_0/n2828 ) );
  nor_x1_sg U10617 ( .A(n7325), .B(n811), .X(\update_output_0/n2592 ) );
  nor_x1_sg U10618 ( .A(n7324), .B(n811), .X(\update_output_0/n2588 ) );
  nor_x1_sg U10619 ( .A(n7325), .B(n813), .X(\update_output_0/n2512 ) );
  nor_x1_sg U10620 ( .A(n7324), .B(n813), .X(\update_output_0/n2508 ) );
  nor_x1_sg U10621 ( .A(n7325), .B(n819), .X(\update_output_0/n2272 ) );
  nor_x1_sg U10622 ( .A(n7324), .B(n819), .X(\update_output_0/n2268 ) );
  nor_x1_sg U10623 ( .A(n7325), .B(n821), .X(\update_output_0/n2192 ) );
  nor_x1_sg U10624 ( .A(n7324), .B(n821), .X(\update_output_0/n2188 ) );
  nand_x2_sg U10625 ( .A(n1365), .B(n1366), .X(n1195) );
  nor_x1_sg U10626 ( .A(n7346), .B(n808), .X(\update_output_0/n2804 ) );
  nor_x1_sg U10627 ( .A(n7347), .B(n808), .X(\update_output_0/n2800 ) );
  nor_x1_sg U10628 ( .A(n7332), .B(n808), .X(\update_output_0/n2796 ) );
  nor_x1_sg U10629 ( .A(n7331), .B(n808), .X(\update_output_0/n2792 ) );
  nor_x1_sg U10630 ( .A(n7330), .B(n808), .X(\update_output_0/n2788 ) );
  nor_x1_sg U10631 ( .A(n7355), .B(n808), .X(\update_output_0/n2784 ) );
  nor_x1_sg U10632 ( .A(n7357), .B(n808), .X(\update_output_0/n2780 ) );
  nor_x1_sg U10633 ( .A(n7329), .B(n808), .X(\update_output_0/n2776 ) );
  nor_x1_sg U10634 ( .A(n7328), .B(n808), .X(\update_output_0/n2772 ) );
  nor_x1_sg U10635 ( .A(n7327), .B(n808), .X(\update_output_0/n2768 ) );
  nor_x1_sg U10636 ( .A(n7365), .B(n808), .X(\update_output_0/n2764 ) );
  nor_x1_sg U10637 ( .A(n7367), .B(n808), .X(\update_output_0/n2760 ) );
  nor_x1_sg U10638 ( .A(n7326), .B(n808), .X(\update_output_0/n2756 ) );
  nor_x1_sg U10639 ( .A(n7346), .B(n810), .X(\update_output_0/n2724 ) );
  nor_x1_sg U10640 ( .A(n7347), .B(n810), .X(\update_output_0/n2720 ) );
  nor_x1_sg U10641 ( .A(n7332), .B(n810), .X(\update_output_0/n2716 ) );
  nor_x1_sg U10642 ( .A(n7331), .B(n810), .X(\update_output_0/n2712 ) );
  nor_x1_sg U10643 ( .A(n7330), .B(n810), .X(\update_output_0/n2708 ) );
  nor_x1_sg U10644 ( .A(n7355), .B(n810), .X(\update_output_0/n2704 ) );
  nor_x1_sg U10645 ( .A(n7357), .B(n810), .X(\update_output_0/n2700 ) );
  nor_x1_sg U10646 ( .A(n7329), .B(n810), .X(\update_output_0/n2696 ) );
  nor_x1_sg U10647 ( .A(n7328), .B(n810), .X(\update_output_0/n2692 ) );
  nor_x1_sg U10648 ( .A(n7327), .B(n810), .X(\update_output_0/n2688 ) );
  nor_x1_sg U10649 ( .A(n7365), .B(n810), .X(\update_output_0/n2684 ) );
  nor_x1_sg U10650 ( .A(n7367), .B(n810), .X(\update_output_0/n2680 ) );
  nor_x1_sg U10651 ( .A(n7326), .B(n810), .X(\update_output_0/n2676 ) );
  nor_x1_sg U10652 ( .A(n7346), .B(n817), .X(\update_output_0/n2404 ) );
  nor_x1_sg U10653 ( .A(n7347), .B(n817), .X(\update_output_0/n2400 ) );
  nor_x1_sg U10654 ( .A(n7332), .B(n817), .X(\update_output_0/n2396 ) );
  nor_x1_sg U10655 ( .A(n7331), .B(n817), .X(\update_output_0/n2392 ) );
  nor_x1_sg U10656 ( .A(n7330), .B(n817), .X(\update_output_0/n2388 ) );
  nor_x1_sg U10657 ( .A(n7355), .B(n817), .X(\update_output_0/n2384 ) );
  nor_x1_sg U10658 ( .A(n7357), .B(n817), .X(\update_output_0/n2380 ) );
  nor_x1_sg U10659 ( .A(n7329), .B(n817), .X(\update_output_0/n2376 ) );
  nor_x1_sg U10660 ( .A(n7328), .B(n817), .X(\update_output_0/n2372 ) );
  nor_x1_sg U10661 ( .A(n7327), .B(n817), .X(\update_output_0/n2368 ) );
  nor_x1_sg U10662 ( .A(n7365), .B(n817), .X(\update_output_0/n2364 ) );
  nor_x1_sg U10663 ( .A(n7367), .B(n817), .X(\update_output_0/n2360 ) );
  nor_x1_sg U10664 ( .A(n7326), .B(n817), .X(\update_output_0/n2356 ) );
  nor_x1_sg U10665 ( .A(n7347), .B(n772), .X(\update_output_0/n3440 ) );
  nor_x1_sg U10666 ( .A(n7332), .B(n772), .X(\update_output_0/n3436 ) );
  nor_x1_sg U10667 ( .A(n7331), .B(n772), .X(\update_output_0/n3432 ) );
  nor_x1_sg U10668 ( .A(n7330), .B(n772), .X(\update_output_0/n3428 ) );
  nor_x1_sg U10669 ( .A(n7355), .B(n772), .X(\update_output_0/n3424 ) );
  nor_x1_sg U10670 ( .A(n7357), .B(n772), .X(\update_output_0/n3420 ) );
  nor_x1_sg U10671 ( .A(n7329), .B(n772), .X(\update_output_0/n3416 ) );
  nor_x1_sg U10672 ( .A(n7328), .B(n772), .X(\update_output_0/n3412 ) );
  nor_x1_sg U10673 ( .A(n7327), .B(n772), .X(\update_output_0/n3408 ) );
  nor_x1_sg U10674 ( .A(n7365), .B(n772), .X(\update_output_0/n3404 ) );
  nor_x1_sg U10675 ( .A(n7367), .B(n772), .X(\update_output_0/n3400 ) );
  nor_x1_sg U10676 ( .A(n7326), .B(n772), .X(\update_output_0/n3396 ) );
  nor_x1_sg U10677 ( .A(n7325), .B(n772), .X(\update_output_0/n3392 ) );
  nor_x1_sg U10678 ( .A(n7346), .B(n792), .X(\update_output_0/n3364 ) );
  nor_x1_sg U10679 ( .A(n7347), .B(n792), .X(\update_output_0/n3360 ) );
  nor_x1_sg U10680 ( .A(n7332), .B(n792), .X(\update_output_0/n3356 ) );
  nor_x1_sg U10681 ( .A(n7331), .B(n792), .X(\update_output_0/n3352 ) );
  nor_x1_sg U10682 ( .A(n7330), .B(n792), .X(\update_output_0/n3348 ) );
  nor_x1_sg U10683 ( .A(n7355), .B(n792), .X(\update_output_0/n3344 ) );
  nor_x1_sg U10684 ( .A(n7357), .B(n792), .X(\update_output_0/n3340 ) );
  nor_x1_sg U10685 ( .A(n7329), .B(n792), .X(\update_output_0/n3336 ) );
  nor_x1_sg U10686 ( .A(n7328), .B(n792), .X(\update_output_0/n3332 ) );
  nor_x1_sg U10687 ( .A(n7327), .B(n792), .X(\update_output_0/n3328 ) );
  nor_x1_sg U10688 ( .A(n7365), .B(n792), .X(\update_output_0/n3324 ) );
  nor_x1_sg U10689 ( .A(n7367), .B(n792), .X(\update_output_0/n3320 ) );
  nor_x1_sg U10690 ( .A(n7326), .B(n792), .X(\update_output_0/n3316 ) );
  nor_x1_sg U10691 ( .A(n7401), .B(n811), .X(\update_output_0/n2664 ) );
  nor_x1_sg U10692 ( .A(n7336), .B(n811), .X(\update_output_0/n2660 ) );
  nor_x1_sg U10693 ( .A(n7335), .B(n811), .X(\update_output_0/n2656 ) );
  nor_x1_sg U10694 ( .A(n7334), .B(n811), .X(\update_output_0/n2652 ) );
  nor_x1_sg U10695 ( .A(n7333), .B(n811), .X(\update_output_0/n2648 ) );
  nor_x1_sg U10696 ( .A(n7401), .B(n813), .X(\update_output_0/n2584 ) );
  nor_x1_sg U10697 ( .A(n7336), .B(n813), .X(\update_output_0/n2580 ) );
  nor_x1_sg U10698 ( .A(n7335), .B(n813), .X(\update_output_0/n2576 ) );
  nor_x1_sg U10699 ( .A(n7334), .B(n813), .X(\update_output_0/n2572 ) );
  nor_x1_sg U10700 ( .A(n7333), .B(n813), .X(\update_output_0/n2568 ) );
  nor_x1_sg U10701 ( .A(n7401), .B(n819), .X(\update_output_0/n2344 ) );
  nor_x1_sg U10702 ( .A(n7336), .B(n819), .X(\update_output_0/n2340 ) );
  nor_x1_sg U10703 ( .A(n7335), .B(n819), .X(\update_output_0/n2336 ) );
  nor_x1_sg U10704 ( .A(n7334), .B(n819), .X(\update_output_0/n2332 ) );
  nor_x1_sg U10705 ( .A(n7333), .B(n819), .X(\update_output_0/n2328 ) );
  nor_x1_sg U10706 ( .A(n7401), .B(n821), .X(\update_output_0/n2264 ) );
  nor_x1_sg U10707 ( .A(n7336), .B(n821), .X(\update_output_0/n2260 ) );
  nor_x1_sg U10708 ( .A(n7335), .B(n821), .X(\update_output_0/n2256 ) );
  nor_x1_sg U10709 ( .A(n7334), .B(n821), .X(\update_output_0/n2252 ) );
  nor_x1_sg U10710 ( .A(n7333), .B(n821), .X(\update_output_0/n2248 ) );
  nor_x1_sg U10711 ( .A(n7401), .B(n803), .X(\update_output_0/n3064 ) );
  nor_x1_sg U10712 ( .A(n7336), .B(n803), .X(\update_output_0/n3060 ) );
  nor_x1_sg U10713 ( .A(n7335), .B(n803), .X(\update_output_0/n3056 ) );
  nor_x1_sg U10714 ( .A(n7334), .B(n803), .X(\update_output_0/n3052 ) );
  nor_x1_sg U10715 ( .A(n7333), .B(n803), .X(\update_output_0/n3048 ) );
  nor_x1_sg U10716 ( .A(n7324), .B(n772), .X(\update_output_0/n3388 ) );
  nor_x1_sg U10717 ( .A(n7325), .B(n792), .X(\update_output_0/n3312 ) );
  nor_x1_sg U10718 ( .A(n7324), .B(n792), .X(\update_output_0/n3308 ) );
  nor_x1_sg U10719 ( .A(n7325), .B(n808), .X(\update_output_0/n2752 ) );
  nor_x1_sg U10720 ( .A(n7324), .B(n808), .X(\update_output_0/n2748 ) );
  nor_x1_sg U10721 ( .A(n7325), .B(n810), .X(\update_output_0/n2672 ) );
  nor_x1_sg U10722 ( .A(n7324), .B(n810), .X(\update_output_0/n2668 ) );
  nor_x1_sg U10723 ( .A(n7325), .B(n817), .X(\update_output_0/n2352 ) );
  nor_x1_sg U10724 ( .A(n7324), .B(n817), .X(\update_output_0/n2348 ) );
  nor_x1_sg U10725 ( .A(n7401), .B(n772), .X(\update_output_0/n2180 ) );
  nand_x2_sg U10726 ( .A(n7367), .B(n7365), .X(n1367) );
  nand_x2_sg U10727 ( .A(n849), .B(n850), .X(n848) );
  nor_x1_sg U10728 ( .A(n7343), .B(n7341), .X(n849) );
  nor_x1_sg U10729 ( .A(n7339), .B(n851), .X(n850) );
  nand_x2_sg U10730 ( .A(n7336), .B(n7401), .X(n851) );
  nand_x2_sg U10731 ( .A(n1027), .B(n1028), .X(n847) );
  nor_x1_sg U10732 ( .A(n7354), .B(n7352), .X(n1027) );
  nor_x1_sg U10733 ( .A(n7350), .B(n1029), .X(n1028) );
  nand_x2_sg U10734 ( .A(n7347), .B(n7344), .X(n1029) );
  nand_x2_sg U10735 ( .A(n1197), .B(n1198), .X(n1196) );
  nor_x1_sg U10736 ( .A(n7364), .B(n7362), .X(n1197) );
  nor_x1_sg U10737 ( .A(n7360), .B(n1199), .X(n1198) );
  nand_x2_sg U10738 ( .A(n7357), .B(n7355), .X(n1199) );
  nor_x1_sg U10739 ( .A(n9247), .B(n7569), .X(n880) );
  nand_x4_sg U10740 ( .A(n7419), .B(n5080), .X(n4102) );
  nand_x2_sg U10741 ( .A(n4017), .B(n7558), .X(n4016) );
  nor_x1_sg U10742 ( .A(n7568), .B(n7526), .X(n4190) );
  inv_x4_sg U10743 ( .A(n3823), .X(n7525) );
  nor_x1_sg U10744 ( .A(n7343), .B(n808), .X(\update_output_0/n2807 ) );
  nor_x1_sg U10745 ( .A(n7345), .B(n808), .X(\update_output_0/n2803 ) );
  nor_x1_sg U10746 ( .A(n7348), .B(n808), .X(\update_output_0/n2799 ) );
  nor_x1_sg U10747 ( .A(n7350), .B(n808), .X(\update_output_0/n2795 ) );
  nor_x1_sg U10748 ( .A(n7352), .B(n808), .X(\update_output_0/n2791 ) );
  nor_x1_sg U10749 ( .A(n7354), .B(n808), .X(\update_output_0/n2787 ) );
  nor_x1_sg U10750 ( .A(n7356), .B(n808), .X(\update_output_0/n2783 ) );
  nor_x1_sg U10751 ( .A(n7358), .B(n808), .X(\update_output_0/n2779 ) );
  nor_x1_sg U10752 ( .A(n7360), .B(n808), .X(\update_output_0/n2775 ) );
  nor_x1_sg U10753 ( .A(n7362), .B(n808), .X(\update_output_0/n2771 ) );
  nor_x1_sg U10754 ( .A(n7364), .B(n808), .X(\update_output_0/n2767 ) );
  nor_x1_sg U10755 ( .A(n7366), .B(n808), .X(\update_output_0/n2763 ) );
  nor_x1_sg U10756 ( .A(n7368), .B(n808), .X(\update_output_0/n2759 ) );
  nor_x1_sg U10757 ( .A(n7370), .B(n808), .X(\update_output_0/n2755 ) );
  nor_x1_sg U10758 ( .A(n7343), .B(n810), .X(\update_output_0/n2727 ) );
  nor_x1_sg U10759 ( .A(n7345), .B(n810), .X(\update_output_0/n2723 ) );
  nor_x1_sg U10760 ( .A(n7348), .B(n810), .X(\update_output_0/n2719 ) );
  nor_x1_sg U10761 ( .A(n7350), .B(n810), .X(\update_output_0/n2715 ) );
  nor_x1_sg U10762 ( .A(n7352), .B(n810), .X(\update_output_0/n2711 ) );
  nor_x1_sg U10763 ( .A(n7354), .B(n810), .X(\update_output_0/n2707 ) );
  nor_x1_sg U10764 ( .A(n7356), .B(n810), .X(\update_output_0/n2703 ) );
  nor_x1_sg U10765 ( .A(n7358), .B(n810), .X(\update_output_0/n2699 ) );
  nor_x1_sg U10766 ( .A(n7360), .B(n810), .X(\update_output_0/n2695 ) );
  nor_x1_sg U10767 ( .A(n7362), .B(n810), .X(\update_output_0/n2691 ) );
  nor_x1_sg U10768 ( .A(n7364), .B(n810), .X(\update_output_0/n2687 ) );
  nor_x1_sg U10769 ( .A(n7366), .B(n810), .X(\update_output_0/n2683 ) );
  nor_x1_sg U10770 ( .A(n7368), .B(n810), .X(\update_output_0/n2679 ) );
  nor_x1_sg U10771 ( .A(n7370), .B(n810), .X(\update_output_0/n2675 ) );
  nor_x1_sg U10772 ( .A(n7343), .B(n815), .X(\update_output_0/n2487 ) );
  nor_x1_sg U10773 ( .A(n7346), .B(n815), .X(\update_output_0/n2484 ) );
  nor_x1_sg U10774 ( .A(n7345), .B(n815), .X(\update_output_0/n2483 ) );
  nor_x1_sg U10775 ( .A(n7347), .B(n815), .X(\update_output_0/n2480 ) );
  nor_x1_sg U10776 ( .A(n7348), .B(n815), .X(\update_output_0/n2479 ) );
  nor_x1_sg U10777 ( .A(n7332), .B(n815), .X(\update_output_0/n2476 ) );
  nor_x1_sg U10778 ( .A(n7350), .B(n815), .X(\update_output_0/n2475 ) );
  nor_x1_sg U10779 ( .A(n7331), .B(n815), .X(\update_output_0/n2472 ) );
  nor_x1_sg U10780 ( .A(n7352), .B(n815), .X(\update_output_0/n2471 ) );
  nor_x1_sg U10781 ( .A(n7330), .B(n815), .X(\update_output_0/n2468 ) );
  nor_x1_sg U10782 ( .A(n7354), .B(n815), .X(\update_output_0/n2467 ) );
  nor_x1_sg U10783 ( .A(n7355), .B(n815), .X(\update_output_0/n2464 ) );
  nor_x1_sg U10784 ( .A(n7356), .B(n815), .X(\update_output_0/n2463 ) );
  nor_x1_sg U10785 ( .A(n7357), .B(n815), .X(\update_output_0/n2460 ) );
  nor_x1_sg U10786 ( .A(n7358), .B(n815), .X(\update_output_0/n2459 ) );
  nor_x1_sg U10787 ( .A(n7329), .B(n815), .X(\update_output_0/n2456 ) );
  nor_x1_sg U10788 ( .A(n7360), .B(n815), .X(\update_output_0/n2455 ) );
  nor_x1_sg U10789 ( .A(n7328), .B(n815), .X(\update_output_0/n2452 ) );
  nor_x1_sg U10790 ( .A(n7362), .B(n815), .X(\update_output_0/n2451 ) );
  nor_x1_sg U10791 ( .A(n7327), .B(n815), .X(\update_output_0/n2448 ) );
  nor_x1_sg U10792 ( .A(n7364), .B(n815), .X(\update_output_0/n2447 ) );
  nor_x1_sg U10793 ( .A(n7365), .B(n815), .X(\update_output_0/n2444 ) );
  nor_x1_sg U10794 ( .A(n7366), .B(n815), .X(\update_output_0/n2443 ) );
  nor_x1_sg U10795 ( .A(n7367), .B(n815), .X(\update_output_0/n2440 ) );
  nor_x1_sg U10796 ( .A(n7368), .B(n815), .X(\update_output_0/n2439 ) );
  nor_x1_sg U10797 ( .A(n7326), .B(n815), .X(\update_output_0/n2436 ) );
  nor_x1_sg U10798 ( .A(n7370), .B(n815), .X(\update_output_0/n2435 ) );
  nor_x1_sg U10799 ( .A(n7343), .B(n817), .X(\update_output_0/n2407 ) );
  nor_x1_sg U10800 ( .A(n7345), .B(n817), .X(\update_output_0/n2403 ) );
  nor_x1_sg U10801 ( .A(n7348), .B(n817), .X(\update_output_0/n2399 ) );
  nor_x1_sg U10802 ( .A(n7350), .B(n817), .X(\update_output_0/n2395 ) );
  nor_x1_sg U10803 ( .A(n7352), .B(n817), .X(\update_output_0/n2391 ) );
  nor_x1_sg U10804 ( .A(n7354), .B(n817), .X(\update_output_0/n2387 ) );
  nor_x1_sg U10805 ( .A(n7356), .B(n817), .X(\update_output_0/n2383 ) );
  nor_x1_sg U10806 ( .A(n7358), .B(n817), .X(\update_output_0/n2379 ) );
  nor_x1_sg U10807 ( .A(n7360), .B(n817), .X(\update_output_0/n2375 ) );
  nor_x1_sg U10808 ( .A(n7362), .B(n817), .X(\update_output_0/n2371 ) );
  nor_x1_sg U10809 ( .A(n7364), .B(n817), .X(\update_output_0/n2367 ) );
  nor_x1_sg U10810 ( .A(n7366), .B(n817), .X(\update_output_0/n2363 ) );
  nor_x1_sg U10811 ( .A(n7368), .B(n817), .X(\update_output_0/n2359 ) );
  nor_x1_sg U10812 ( .A(n7370), .B(n817), .X(\update_output_0/n2355 ) );
  nor_x1_sg U10813 ( .A(n7345), .B(n772), .X(\update_output_0/n3443 ) );
  nor_x1_sg U10814 ( .A(n7348), .B(n772), .X(\update_output_0/n3439 ) );
  nor_x1_sg U10815 ( .A(n7350), .B(n772), .X(\update_output_0/n3435 ) );
  nor_x1_sg U10816 ( .A(n7352), .B(n772), .X(\update_output_0/n3431 ) );
  nor_x1_sg U10817 ( .A(n7354), .B(n772), .X(\update_output_0/n3427 ) );
  nor_x1_sg U10818 ( .A(n7356), .B(n772), .X(\update_output_0/n3423 ) );
  nor_x1_sg U10819 ( .A(n7358), .B(n772), .X(\update_output_0/n3419 ) );
  nor_x1_sg U10820 ( .A(n7360), .B(n772), .X(\update_output_0/n3415 ) );
  nor_x1_sg U10821 ( .A(n7362), .B(n772), .X(\update_output_0/n3411 ) );
  nor_x1_sg U10822 ( .A(n7364), .B(n772), .X(\update_output_0/n3407 ) );
  nor_x1_sg U10823 ( .A(n7366), .B(n772), .X(\update_output_0/n3403 ) );
  nor_x1_sg U10824 ( .A(n7368), .B(n772), .X(\update_output_0/n3399 ) );
  nor_x1_sg U10825 ( .A(n7370), .B(n772), .X(\update_output_0/n3395 ) );
  nor_x1_sg U10826 ( .A(n7372), .B(n772), .X(\update_output_0/n3391 ) );
  nor_x1_sg U10827 ( .A(n7343), .B(n792), .X(\update_output_0/n3367 ) );
  nor_x1_sg U10828 ( .A(n7345), .B(n792), .X(\update_output_0/n3363 ) );
  nor_x1_sg U10829 ( .A(n7348), .B(n792), .X(\update_output_0/n3359 ) );
  nor_x1_sg U10830 ( .A(n7350), .B(n792), .X(\update_output_0/n3355 ) );
  nor_x1_sg U10831 ( .A(n7352), .B(n792), .X(\update_output_0/n3351 ) );
  nor_x1_sg U10832 ( .A(n7354), .B(n792), .X(\update_output_0/n3347 ) );
  nor_x1_sg U10833 ( .A(n7356), .B(n792), .X(\update_output_0/n3343 ) );
  nor_x1_sg U10834 ( .A(n7358), .B(n792), .X(\update_output_0/n3339 ) );
  nor_x1_sg U10835 ( .A(n7360), .B(n792), .X(\update_output_0/n3335 ) );
  nor_x1_sg U10836 ( .A(n7362), .B(n792), .X(\update_output_0/n3331 ) );
  nor_x1_sg U10837 ( .A(n7364), .B(n792), .X(\update_output_0/n3327 ) );
  nor_x1_sg U10838 ( .A(n7366), .B(n792), .X(\update_output_0/n3323 ) );
  nor_x1_sg U10839 ( .A(n7368), .B(n792), .X(\update_output_0/n3319 ) );
  nor_x1_sg U10840 ( .A(n7370), .B(n792), .X(\update_output_0/n3315 ) );
  nor_x1_sg U10841 ( .A(n7343), .B(n811), .X(\update_output_0/n2647 ) );
  nor_x1_sg U10842 ( .A(n7345), .B(n811), .X(\update_output_0/n2643 ) );
  nor_x1_sg U10843 ( .A(n7348), .B(n811), .X(\update_output_0/n2639 ) );
  nor_x1_sg U10844 ( .A(n7350), .B(n811), .X(\update_output_0/n2635 ) );
  nor_x1_sg U10845 ( .A(n7352), .B(n811), .X(\update_output_0/n2631 ) );
  nor_x1_sg U10846 ( .A(n7354), .B(n811), .X(\update_output_0/n2627 ) );
  nor_x1_sg U10847 ( .A(n7356), .B(n811), .X(\update_output_0/n2623 ) );
  nor_x1_sg U10848 ( .A(n7358), .B(n811), .X(\update_output_0/n2619 ) );
  nor_x1_sg U10849 ( .A(n7360), .B(n811), .X(\update_output_0/n2615 ) );
  nor_x1_sg U10850 ( .A(n7362), .B(n811), .X(\update_output_0/n2611 ) );
  nor_x1_sg U10851 ( .A(n7364), .B(n811), .X(\update_output_0/n2607 ) );
  nor_x1_sg U10852 ( .A(n7366), .B(n811), .X(\update_output_0/n2603 ) );
  nor_x1_sg U10853 ( .A(n7368), .B(n811), .X(\update_output_0/n2599 ) );
  nor_x1_sg U10854 ( .A(n7370), .B(n811), .X(\update_output_0/n2595 ) );
  nor_x1_sg U10855 ( .A(n7343), .B(n813), .X(\update_output_0/n2567 ) );
  nor_x1_sg U10856 ( .A(n7345), .B(n813), .X(\update_output_0/n2563 ) );
  nor_x1_sg U10857 ( .A(n7348), .B(n813), .X(\update_output_0/n2559 ) );
  nor_x1_sg U10858 ( .A(n7350), .B(n813), .X(\update_output_0/n2555 ) );
  nor_x1_sg U10859 ( .A(n7352), .B(n813), .X(\update_output_0/n2551 ) );
  nor_x1_sg U10860 ( .A(n7354), .B(n813), .X(\update_output_0/n2547 ) );
  nor_x1_sg U10861 ( .A(n7356), .B(n813), .X(\update_output_0/n2543 ) );
  nor_x1_sg U10862 ( .A(n7358), .B(n813), .X(\update_output_0/n2539 ) );
  nor_x1_sg U10863 ( .A(n7360), .B(n813), .X(\update_output_0/n2535 ) );
  nor_x1_sg U10864 ( .A(n7362), .B(n813), .X(\update_output_0/n2531 ) );
  nor_x1_sg U10865 ( .A(n7364), .B(n813), .X(\update_output_0/n2527 ) );
  nor_x1_sg U10866 ( .A(n7366), .B(n813), .X(\update_output_0/n2523 ) );
  nor_x1_sg U10867 ( .A(n7368), .B(n813), .X(\update_output_0/n2519 ) );
  nor_x1_sg U10868 ( .A(n7370), .B(n813), .X(\update_output_0/n2515 ) );
  nor_x1_sg U10869 ( .A(n7343), .B(n819), .X(\update_output_0/n2327 ) );
  nor_x1_sg U10870 ( .A(n7345), .B(n819), .X(\update_output_0/n2323 ) );
  nor_x1_sg U10871 ( .A(n7348), .B(n819), .X(\update_output_0/n2319 ) );
  nor_x1_sg U10872 ( .A(n7350), .B(n819), .X(\update_output_0/n2315 ) );
  nor_x1_sg U10873 ( .A(n7352), .B(n819), .X(\update_output_0/n2311 ) );
  nor_x1_sg U10874 ( .A(n7354), .B(n819), .X(\update_output_0/n2307 ) );
  nor_x1_sg U10875 ( .A(n7356), .B(n819), .X(\update_output_0/n2303 ) );
  nor_x1_sg U10876 ( .A(n7358), .B(n819), .X(\update_output_0/n2299 ) );
  nor_x1_sg U10877 ( .A(n7360), .B(n819), .X(\update_output_0/n2295 ) );
  nor_x1_sg U10878 ( .A(n7362), .B(n819), .X(\update_output_0/n2291 ) );
  nor_x1_sg U10879 ( .A(n7364), .B(n819), .X(\update_output_0/n2287 ) );
  nor_x1_sg U10880 ( .A(n7366), .B(n819), .X(\update_output_0/n2283 ) );
  nor_x1_sg U10881 ( .A(n7368), .B(n819), .X(\update_output_0/n2279 ) );
  nor_x1_sg U10882 ( .A(n7370), .B(n819), .X(\update_output_0/n2275 ) );
  nor_x1_sg U10883 ( .A(n7343), .B(n821), .X(\update_output_0/n2247 ) );
  nor_x1_sg U10884 ( .A(n7345), .B(n821), .X(\update_output_0/n2243 ) );
  nor_x1_sg U10885 ( .A(n7348), .B(n821), .X(\update_output_0/n2239 ) );
  nor_x1_sg U10886 ( .A(n7350), .B(n821), .X(\update_output_0/n2235 ) );
  nor_x1_sg U10887 ( .A(n7352), .B(n821), .X(\update_output_0/n2231 ) );
  nor_x1_sg U10888 ( .A(n7354), .B(n821), .X(\update_output_0/n2227 ) );
  nor_x1_sg U10889 ( .A(n7356), .B(n821), .X(\update_output_0/n2223 ) );
  nor_x1_sg U10890 ( .A(n7358), .B(n821), .X(\update_output_0/n2219 ) );
  nor_x1_sg U10891 ( .A(n7360), .B(n821), .X(\update_output_0/n2215 ) );
  nor_x1_sg U10892 ( .A(n7362), .B(n821), .X(\update_output_0/n2211 ) );
  nor_x1_sg U10893 ( .A(n7364), .B(n821), .X(\update_output_0/n2207 ) );
  nor_x1_sg U10894 ( .A(n7366), .B(n821), .X(\update_output_0/n2203 ) );
  nor_x1_sg U10895 ( .A(n7368), .B(n821), .X(\update_output_0/n2199 ) );
  nor_x1_sg U10896 ( .A(n7370), .B(n821), .X(\update_output_0/n2195 ) );
  nor_x1_sg U10897 ( .A(n7343), .B(n800), .X(\update_output_0/n3127 ) );
  nor_x1_sg U10898 ( .A(n7346), .B(n800), .X(\update_output_0/n3124 ) );
  nor_x1_sg U10899 ( .A(n777), .B(n800), .X(\update_output_0/n3123 ) );
  nor_x1_sg U10900 ( .A(n7347), .B(n800), .X(\update_output_0/n3120 ) );
  nor_x1_sg U10901 ( .A(n7348), .B(n800), .X(\update_output_0/n3119 ) );
  nor_x1_sg U10902 ( .A(n7332), .B(n800), .X(\update_output_0/n3116 ) );
  nor_x1_sg U10903 ( .A(n7350), .B(n800), .X(\update_output_0/n3115 ) );
  nor_x1_sg U10904 ( .A(n7331), .B(n800), .X(\update_output_0/n3112 ) );
  nor_x1_sg U10905 ( .A(n7352), .B(n800), .X(\update_output_0/n3111 ) );
  nor_x1_sg U10906 ( .A(n7330), .B(n800), .X(\update_output_0/n3108 ) );
  nor_x1_sg U10907 ( .A(n7354), .B(n800), .X(\update_output_0/n3107 ) );
  nor_x1_sg U10908 ( .A(n7355), .B(n800), .X(\update_output_0/n3104 ) );
  nor_x1_sg U10909 ( .A(n7356), .B(n800), .X(\update_output_0/n3103 ) );
  nor_x1_sg U10910 ( .A(n7357), .B(n800), .X(\update_output_0/n3100 ) );
  nor_x1_sg U10911 ( .A(n7358), .B(n800), .X(\update_output_0/n3099 ) );
  nor_x1_sg U10912 ( .A(n7329), .B(n800), .X(\update_output_0/n3096 ) );
  nor_x1_sg U10913 ( .A(n7360), .B(n800), .X(\update_output_0/n3095 ) );
  nor_x1_sg U10914 ( .A(n7328), .B(n800), .X(\update_output_0/n3092 ) );
  nor_x1_sg U10915 ( .A(n7362), .B(n800), .X(\update_output_0/n3091 ) );
  nor_x1_sg U10916 ( .A(n7327), .B(n800), .X(\update_output_0/n3088 ) );
  nor_x1_sg U10917 ( .A(n7364), .B(n800), .X(\update_output_0/n3087 ) );
  nor_x1_sg U10918 ( .A(n7365), .B(n800), .X(\update_output_0/n3084 ) );
  nor_x1_sg U10919 ( .A(n7366), .B(n800), .X(\update_output_0/n3083 ) );
  nor_x1_sg U10920 ( .A(n7367), .B(n800), .X(\update_output_0/n3080 ) );
  nor_x1_sg U10921 ( .A(n7368), .B(n800), .X(\update_output_0/n3079 ) );
  nor_x1_sg U10922 ( .A(n7326), .B(n800), .X(\update_output_0/n3076 ) );
  nor_x1_sg U10923 ( .A(n7370), .B(n800), .X(\update_output_0/n3075 ) );
  nor_x1_sg U10924 ( .A(n7343), .B(n803), .X(\update_output_0/n3047 ) );
  nor_x1_sg U10925 ( .A(n7345), .B(n803), .X(\update_output_0/n3043 ) );
  nor_x1_sg U10926 ( .A(n7348), .B(n803), .X(\update_output_0/n3039 ) );
  nor_x1_sg U10927 ( .A(n7350), .B(n803), .X(\update_output_0/n3035 ) );
  nor_x1_sg U10928 ( .A(n7352), .B(n803), .X(\update_output_0/n3031 ) );
  nor_x1_sg U10929 ( .A(n7354), .B(n803), .X(\update_output_0/n3027 ) );
  nor_x1_sg U10930 ( .A(n7356), .B(n803), .X(\update_output_0/n3023 ) );
  nor_x1_sg U10931 ( .A(n7358), .B(n803), .X(\update_output_0/n3019 ) );
  nor_x1_sg U10932 ( .A(n7360), .B(n803), .X(\update_output_0/n3015 ) );
  nor_x1_sg U10933 ( .A(n7362), .B(n803), .X(\update_output_0/n3011 ) );
  nor_x1_sg U10934 ( .A(n7364), .B(n803), .X(\update_output_0/n3007 ) );
  nor_x1_sg U10935 ( .A(n7366), .B(n803), .X(\update_output_0/n3003 ) );
  nor_x1_sg U10936 ( .A(n7368), .B(n803), .X(\update_output_0/n2999 ) );
  nor_x1_sg U10937 ( .A(n7370), .B(n803), .X(\update_output_0/n2995 ) );
  nor_x1_sg U10938 ( .A(n7343), .B(n805), .X(\update_output_0/n2967 ) );
  nor_x1_sg U10939 ( .A(n7345), .B(n805), .X(\update_output_0/n2963 ) );
  nor_x1_sg U10940 ( .A(n7348), .B(n805), .X(\update_output_0/n2959 ) );
  nor_x1_sg U10941 ( .A(n7350), .B(n805), .X(\update_output_0/n2955 ) );
  nor_x1_sg U10942 ( .A(n7352), .B(n805), .X(\update_output_0/n2951 ) );
  nor_x1_sg U10943 ( .A(n7354), .B(n805), .X(\update_output_0/n2947 ) );
  nor_x1_sg U10944 ( .A(n7356), .B(n805), .X(\update_output_0/n2943 ) );
  nor_x1_sg U10945 ( .A(n7358), .B(n805), .X(\update_output_0/n2939 ) );
  nor_x1_sg U10946 ( .A(n7360), .B(n805), .X(\update_output_0/n2935 ) );
  nor_x1_sg U10947 ( .A(n7362), .B(n805), .X(\update_output_0/n2931 ) );
  nor_x1_sg U10948 ( .A(n7364), .B(n805), .X(\update_output_0/n2927 ) );
  nor_x1_sg U10949 ( .A(n7366), .B(n805), .X(\update_output_0/n2923 ) );
  nor_x1_sg U10950 ( .A(n7368), .B(n805), .X(\update_output_0/n2919 ) );
  nor_x1_sg U10951 ( .A(n7370), .B(n805), .X(\update_output_0/n2915 ) );
  nor_x1_sg U10952 ( .A(n7343), .B(n806), .X(\update_output_0/n2887 ) );
  nor_x1_sg U10953 ( .A(n7345), .B(n806), .X(\update_output_0/n2883 ) );
  nor_x1_sg U10954 ( .A(n7348), .B(n806), .X(\update_output_0/n2879 ) );
  nor_x1_sg U10955 ( .A(n7350), .B(n806), .X(\update_output_0/n2875 ) );
  nor_x1_sg U10956 ( .A(n7352), .B(n806), .X(\update_output_0/n2871 ) );
  nor_x1_sg U10957 ( .A(n7354), .B(n806), .X(\update_output_0/n2867 ) );
  nor_x1_sg U10958 ( .A(n7356), .B(n806), .X(\update_output_0/n2863 ) );
  nor_x1_sg U10959 ( .A(n7358), .B(n806), .X(\update_output_0/n2859 ) );
  nor_x1_sg U10960 ( .A(n7360), .B(n806), .X(\update_output_0/n2855 ) );
  nor_x1_sg U10961 ( .A(n7362), .B(n806), .X(\update_output_0/n2851 ) );
  nor_x1_sg U10962 ( .A(n7364), .B(n806), .X(\update_output_0/n2847 ) );
  nor_x1_sg U10963 ( .A(n7366), .B(n806), .X(\update_output_0/n2843 ) );
  nor_x1_sg U10964 ( .A(n7368), .B(n806), .X(\update_output_0/n2839 ) );
  nor_x1_sg U10965 ( .A(n7370), .B(n806), .X(\update_output_0/n2835 ) );
  nor_x1_sg U10966 ( .A(n7343), .B(n798), .X(\update_output_0/n3207 ) );
  nor_x1_sg U10967 ( .A(n7345), .B(n798), .X(\update_output_0/n3203 ) );
  nor_x1_sg U10968 ( .A(n7348), .B(n798), .X(\update_output_0/n3199 ) );
  nor_x1_sg U10969 ( .A(n7350), .B(n798), .X(\update_output_0/n3195 ) );
  nor_x1_sg U10970 ( .A(n7352), .B(n798), .X(\update_output_0/n3191 ) );
  nor_x1_sg U10971 ( .A(n7354), .B(n798), .X(\update_output_0/n3187 ) );
  nor_x1_sg U10972 ( .A(n7356), .B(n798), .X(\update_output_0/n3183 ) );
  nor_x1_sg U10973 ( .A(n7358), .B(n798), .X(\update_output_0/n3179 ) );
  nor_x1_sg U10974 ( .A(n7360), .B(n798), .X(\update_output_0/n3175 ) );
  nor_x1_sg U10975 ( .A(n7362), .B(n798), .X(\update_output_0/n3171 ) );
  nor_x1_sg U10976 ( .A(n7364), .B(n798), .X(\update_output_0/n3167 ) );
  nor_x1_sg U10977 ( .A(n7366), .B(n798), .X(\update_output_0/n3163 ) );
  nor_x1_sg U10978 ( .A(n7368), .B(n798), .X(\update_output_0/n3159 ) );
  nor_x1_sg U10979 ( .A(n7370), .B(n798), .X(\update_output_0/n3155 ) );
  nor_x1_sg U10980 ( .A(n7343), .B(n795), .X(\update_output_0/n3287 ) );
  nor_x1_sg U10981 ( .A(n7345), .B(n795), .X(\update_output_0/n3283 ) );
  nor_x1_sg U10982 ( .A(n7348), .B(n795), .X(\update_output_0/n3279 ) );
  nor_x1_sg U10983 ( .A(n7350), .B(n795), .X(\update_output_0/n3275 ) );
  nor_x1_sg U10984 ( .A(n7352), .B(n795), .X(\update_output_0/n3271 ) );
  nor_x1_sg U10985 ( .A(n7354), .B(n795), .X(\update_output_0/n3267 ) );
  nor_x1_sg U10986 ( .A(n7356), .B(n795), .X(\update_output_0/n3263 ) );
  nor_x1_sg U10987 ( .A(n7358), .B(n795), .X(\update_output_0/n3259 ) );
  nor_x1_sg U10988 ( .A(n7360), .B(n795), .X(\update_output_0/n3255 ) );
  nor_x1_sg U10989 ( .A(n7362), .B(n795), .X(\update_output_0/n3251 ) );
  nor_x1_sg U10990 ( .A(n7364), .B(n795), .X(\update_output_0/n3247 ) );
  nor_x1_sg U10991 ( .A(n7366), .B(n795), .X(\update_output_0/n3243 ) );
  nor_x1_sg U10992 ( .A(n7368), .B(n795), .X(\update_output_0/n3239 ) );
  nor_x1_sg U10993 ( .A(n7370), .B(n795), .X(\update_output_0/n3235 ) );
  nor_x1_sg U10994 ( .A(n7401), .B(n808), .X(\update_output_0/n2824 ) );
  nor_x1_sg U10995 ( .A(n7402), .B(n808), .X(\update_output_0/n2823 ) );
  nor_x1_sg U10996 ( .A(n7336), .B(n808), .X(\update_output_0/n2820 ) );
  nor_x1_sg U10997 ( .A(n7337), .B(n808), .X(\update_output_0/n2819 ) );
  nor_x1_sg U10998 ( .A(n7335), .B(n808), .X(\update_output_0/n2816 ) );
  nor_x1_sg U10999 ( .A(n7339), .B(n808), .X(\update_output_0/n2815 ) );
  nor_x1_sg U11000 ( .A(n7334), .B(n808), .X(\update_output_0/n2812 ) );
  nor_x1_sg U11001 ( .A(n7341), .B(n808), .X(\update_output_0/n2811 ) );
  nor_x1_sg U11002 ( .A(n7333), .B(n808), .X(\update_output_0/n2808 ) );
  nor_x1_sg U11003 ( .A(n7401), .B(n810), .X(\update_output_0/n2744 ) );
  nor_x1_sg U11004 ( .A(n7402), .B(n810), .X(\update_output_0/n2743 ) );
  nor_x1_sg U11005 ( .A(n7336), .B(n810), .X(\update_output_0/n2740 ) );
  nor_x1_sg U11006 ( .A(n7337), .B(n810), .X(\update_output_0/n2739 ) );
  nor_x1_sg U11007 ( .A(n7335), .B(n810), .X(\update_output_0/n2736 ) );
  nor_x1_sg U11008 ( .A(n7339), .B(n810), .X(\update_output_0/n2735 ) );
  nor_x1_sg U11009 ( .A(n7334), .B(n810), .X(\update_output_0/n2732 ) );
  nor_x1_sg U11010 ( .A(n7341), .B(n810), .X(\update_output_0/n2731 ) );
  nor_x1_sg U11011 ( .A(n7333), .B(n810), .X(\update_output_0/n2728 ) );
  nor_x1_sg U11012 ( .A(n7401), .B(n817), .X(\update_output_0/n2424 ) );
  nor_x1_sg U11013 ( .A(n7402), .B(n817), .X(\update_output_0/n2423 ) );
  nor_x1_sg U11014 ( .A(n7336), .B(n817), .X(\update_output_0/n2420 ) );
  nor_x1_sg U11015 ( .A(n7337), .B(n817), .X(\update_output_0/n2419 ) );
  nor_x1_sg U11016 ( .A(n7335), .B(n817), .X(\update_output_0/n2416 ) );
  nor_x1_sg U11017 ( .A(n7339), .B(n817), .X(\update_output_0/n2415 ) );
  nor_x1_sg U11018 ( .A(n7334), .B(n817), .X(\update_output_0/n2412 ) );
  nor_x1_sg U11019 ( .A(n7341), .B(n817), .X(\update_output_0/n2411 ) );
  nor_x1_sg U11020 ( .A(n7333), .B(n817), .X(\update_output_0/n2408 ) );
  nor_x1_sg U11021 ( .A(n7336), .B(n772), .X(\update_output_0/n3460 ) );
  nor_x1_sg U11022 ( .A(n7337), .B(n772), .X(\update_output_0/n3459 ) );
  nor_x1_sg U11023 ( .A(n7335), .B(n772), .X(\update_output_0/n3456 ) );
  nor_x1_sg U11024 ( .A(n7339), .B(n772), .X(\update_output_0/n3455 ) );
  nor_x1_sg U11025 ( .A(n7334), .B(n772), .X(\update_output_0/n3452 ) );
  nor_x1_sg U11026 ( .A(n7341), .B(n772), .X(\update_output_0/n3451 ) );
  nor_x1_sg U11027 ( .A(n7333), .B(n772), .X(\update_output_0/n3448 ) );
  nor_x1_sg U11028 ( .A(n7343), .B(n772), .X(\update_output_0/n3447 ) );
  nor_x1_sg U11029 ( .A(n7346), .B(n772), .X(\update_output_0/n3444 ) );
  nor_x1_sg U11030 ( .A(n7401), .B(n792), .X(\update_output_0/n3384 ) );
  nor_x1_sg U11031 ( .A(n7402), .B(n792), .X(\update_output_0/n3383 ) );
  nor_x1_sg U11032 ( .A(n7336), .B(n792), .X(\update_output_0/n3380 ) );
  nor_x1_sg U11033 ( .A(n7337), .B(n792), .X(\update_output_0/n3379 ) );
  nor_x1_sg U11034 ( .A(n7335), .B(n792), .X(\update_output_0/n3376 ) );
  nor_x1_sg U11035 ( .A(n7339), .B(n792), .X(\update_output_0/n3375 ) );
  nor_x1_sg U11036 ( .A(n7334), .B(n792), .X(\update_output_0/n3372 ) );
  nor_x1_sg U11037 ( .A(n7341), .B(n792), .X(\update_output_0/n3371 ) );
  nor_x1_sg U11038 ( .A(n7333), .B(n792), .X(\update_output_0/n3368 ) );
  nor_x1_sg U11039 ( .A(n7402), .B(n811), .X(\update_output_0/n2663 ) );
  nor_x1_sg U11040 ( .A(n7337), .B(n811), .X(\update_output_0/n2659 ) );
  nor_x1_sg U11041 ( .A(n7339), .B(n811), .X(\update_output_0/n2655 ) );
  nor_x1_sg U11042 ( .A(n7341), .B(n811), .X(\update_output_0/n2651 ) );
  nor_x1_sg U11043 ( .A(n7402), .B(n813), .X(\update_output_0/n2583 ) );
  nor_x1_sg U11044 ( .A(n7337), .B(n813), .X(\update_output_0/n2579 ) );
  nor_x1_sg U11045 ( .A(n7339), .B(n813), .X(\update_output_0/n2575 ) );
  nor_x1_sg U11046 ( .A(n7341), .B(n813), .X(\update_output_0/n2571 ) );
  nor_x1_sg U11047 ( .A(n7402), .B(n819), .X(\update_output_0/n2343 ) );
  nor_x1_sg U11048 ( .A(n7337), .B(n819), .X(\update_output_0/n2339 ) );
  nor_x1_sg U11049 ( .A(n7339), .B(n819), .X(\update_output_0/n2335 ) );
  nor_x1_sg U11050 ( .A(n7341), .B(n819), .X(\update_output_0/n2331 ) );
  nor_x1_sg U11051 ( .A(n7402), .B(n821), .X(\update_output_0/n2263 ) );
  nor_x1_sg U11052 ( .A(n7337), .B(n821), .X(\update_output_0/n2259 ) );
  nor_x1_sg U11053 ( .A(n7339), .B(n821), .X(\update_output_0/n2255 ) );
  nor_x1_sg U11054 ( .A(n7341), .B(n821), .X(\update_output_0/n2251 ) );
  nor_x1_sg U11055 ( .A(n7402), .B(n803), .X(\update_output_0/n3063 ) );
  nor_x1_sg U11056 ( .A(n7337), .B(n803), .X(\update_output_0/n3059 ) );
  nor_x1_sg U11057 ( .A(n7339), .B(n803), .X(\update_output_0/n3055 ) );
  nor_x1_sg U11058 ( .A(n7341), .B(n803), .X(\update_output_0/n3051 ) );
  nor_x1_sg U11059 ( .A(n7402), .B(n805), .X(\update_output_0/n2983 ) );
  nor_x1_sg U11060 ( .A(n7337), .B(n805), .X(\update_output_0/n2979 ) );
  nor_x1_sg U11061 ( .A(n7339), .B(n805), .X(\update_output_0/n2975 ) );
  nor_x1_sg U11062 ( .A(n7341), .B(n805), .X(\update_output_0/n2971 ) );
  nor_x1_sg U11063 ( .A(n7402), .B(n806), .X(\update_output_0/n2903 ) );
  nor_x1_sg U11064 ( .A(n7337), .B(n806), .X(\update_output_0/n2899 ) );
  nor_x1_sg U11065 ( .A(n7339), .B(n806), .X(\update_output_0/n2895 ) );
  nor_x1_sg U11066 ( .A(n7341), .B(n806), .X(\update_output_0/n2891 ) );
  nor_x1_sg U11067 ( .A(n7402), .B(n798), .X(\update_output_0/n3223 ) );
  nor_x1_sg U11068 ( .A(n7337), .B(n798), .X(\update_output_0/n3219 ) );
  nor_x1_sg U11069 ( .A(n7339), .B(n798), .X(\update_output_0/n3215 ) );
  nor_x1_sg U11070 ( .A(n7341), .B(n798), .X(\update_output_0/n3211 ) );
  nor_x1_sg U11071 ( .A(n7402), .B(n795), .X(\update_output_0/n3303 ) );
  nor_x1_sg U11072 ( .A(n7337), .B(n795), .X(\update_output_0/n3299 ) );
  nor_x1_sg U11073 ( .A(n7339), .B(n795), .X(\update_output_0/n3295 ) );
  nor_x1_sg U11074 ( .A(n7341), .B(n795), .X(\update_output_0/n3291 ) );
  nor_x1_sg U11075 ( .A(n7325), .B(n800), .X(\update_output_0/n3072 ) );
  nor_x1_sg U11076 ( .A(n7324), .B(n800), .X(\update_output_0/n3068 ) );
  nor_x1_sg U11077 ( .A(n7325), .B(n815), .X(\update_output_0/n2432 ) );
  nor_x1_sg U11078 ( .A(n7324), .B(n815), .X(\update_output_0/n2428 ) );
  nor_x1_sg U11079 ( .A(n7402), .B(n772), .X(\update_output_0/n2179 ) );
  nor_x1_sg U11080 ( .A(n7374), .B(n772), .X(\update_output_0/n3387 ) );
  nor_x1_sg U11081 ( .A(n7372), .B(n792), .X(\update_output_0/n3311 ) );
  nor_x1_sg U11082 ( .A(n7374), .B(n792), .X(\update_output_0/n3307 ) );
  nor_x1_sg U11083 ( .A(n7372), .B(n798), .X(\update_output_0/n3151 ) );
  nor_x1_sg U11084 ( .A(n7374), .B(n798), .X(\update_output_0/n3147 ) );
  nor_x1_sg U11085 ( .A(n7372), .B(n800), .X(\update_output_0/n3071 ) );
  nor_x1_sg U11086 ( .A(n7374), .B(n800), .X(\update_output_0/n3067 ) );
  nor_x1_sg U11087 ( .A(n7372), .B(n805), .X(\update_output_0/n2911 ) );
  nor_x1_sg U11088 ( .A(n7374), .B(n805), .X(\update_output_0/n2907 ) );
  nor_x1_sg U11089 ( .A(n7372), .B(n806), .X(\update_output_0/n2831 ) );
  nor_x1_sg U11090 ( .A(n7374), .B(n806), .X(\update_output_0/n2827 ) );
  nor_x1_sg U11091 ( .A(n7372), .B(n810), .X(\update_output_0/n2671 ) );
  nor_x1_sg U11092 ( .A(n7374), .B(n810), .X(\update_output_0/n2667 ) );
  nor_x1_sg U11093 ( .A(n7372), .B(n811), .X(\update_output_0/n2591 ) );
  nor_x1_sg U11094 ( .A(n7374), .B(n811), .X(\update_output_0/n2587 ) );
  nor_x1_sg U11095 ( .A(n7372), .B(n815), .X(\update_output_0/n2431 ) );
  nor_x1_sg U11096 ( .A(n7374), .B(n815), .X(\update_output_0/n2427 ) );
  nor_x1_sg U11097 ( .A(n7372), .B(n817), .X(\update_output_0/n2351 ) );
  nor_x1_sg U11098 ( .A(n7374), .B(n817), .X(\update_output_0/n2347 ) );
  nor_x1_sg U11099 ( .A(n7372), .B(n821), .X(\update_output_0/n2191 ) );
  nor_x1_sg U11100 ( .A(n7374), .B(n821), .X(\update_output_0/n2187 ) );
  nor_x1_sg U11101 ( .A(n7372), .B(n795), .X(\update_output_0/n3231 ) );
  nor_x1_sg U11102 ( .A(n7374), .B(n795), .X(\update_output_0/n3227 ) );
  nor_x1_sg U11103 ( .A(n7372), .B(n803), .X(\update_output_0/n2991 ) );
  nor_x1_sg U11104 ( .A(n7374), .B(n803), .X(\update_output_0/n2987 ) );
  nor_x1_sg U11105 ( .A(n7372), .B(n808), .X(\update_output_0/n2751 ) );
  nor_x1_sg U11106 ( .A(n7374), .B(n808), .X(\update_output_0/n2747 ) );
  nor_x1_sg U11107 ( .A(n7372), .B(n813), .X(\update_output_0/n2511 ) );
  nor_x1_sg U11108 ( .A(n7374), .B(n813), .X(\update_output_0/n2507 ) );
  nor_x1_sg U11109 ( .A(n7372), .B(n819), .X(\update_output_0/n2271 ) );
  nor_x1_sg U11110 ( .A(n7374), .B(n819), .X(\update_output_0/n2267 ) );
  nand_x4_sg U11111 ( .A(n7419), .B(n4098), .X(n4059) );
  nand_x1_sg U11112 ( .A(n4099), .B(n9205), .X(n4098) );
  nand_x4_sg U11113 ( .A(n7419), .B(n5266), .X(n4407) );
  nand_x1_sg U11114 ( .A(n5267), .B(n9205), .X(n5266) );
  nor_x1_sg U11115 ( .A(n3095), .B(n7571), .X(n5267) );
  nand_x4_sg U11116 ( .A(n7419), .B(n5189), .X(n4020) );
  nor_x1_sg U11117 ( .A(n3095), .B(n3098), .X(n5190) );
  nand_x2_sg U11118 ( .A(n4017), .B(n7323), .X(n5075) );
  nand_x2_sg U11119 ( .A(n9191), .B(n7375), .X(n4301) );
  nand_x2_sg U11120 ( .A(n9191), .B(n4300), .X(n4294) );
  nand_x1_sg U11121 ( .A(n9212), .B(n3813), .X(n5287) );
  inv_x4_sg U11122 ( .A(n7538), .X(n7537) );
  nand_x1_sg U11123 ( .A(n9203), .B(n9216), .X(n5295) );
  nand_x2_sg U11124 ( .A(n5290), .B(n5293), .X(n5299) );
  nand_x2_sg U11125 ( .A(n9192), .B(n4191), .X(n4187) );
  nand_x1_sg U11126 ( .A(n9203), .B(n3101), .X(n5306) );
  nand_x1_sg U11127 ( .A(n4197), .B(n7562), .X(n4395) );
  nand_x1_sg U11128 ( .A(n4197), .B(n7564), .X(n4193) );
  nand_x1_sg U11129 ( .A(n4196), .B(n9247), .X(n4195) );
  nor_x1_sg U11130 ( .A(n7520), .B(n3101), .X(n5273) );
  nor_x1_sg U11131 ( .A(n7559), .B(n8991), .X(n822) );
  nor_x1_sg U11132 ( .A(n9245), .B(n824), .X(\update_output_0/n2183 ) );
  nor_x1_sg U11133 ( .A(n828), .B(n829), .X(\update_mask_0/n988 ) );
  nor_x1_sg U11134 ( .A(n828), .B(n839), .X(\update_mask_0/n1088 ) );
  nor_x1_sg U11135 ( .A(n828), .B(n842), .X(\update_mask_0/n1056 ) );
  nor_x1_sg U11136 ( .A(n828), .B(n825), .X(\update_mask_0/n1024 ) );
  nor_x1_sg U11137 ( .A(n834), .B(n829), .X(\update_mask_0/n1100 ) );
  nor_x1_sg U11138 ( .A(n3101), .B(n829), .X(\update_mask_0/n1092 ) );
  nor_x1_sg U11139 ( .A(n834), .B(n842), .X(\update_mask_0/n1036 ) );
  nor_x1_sg U11140 ( .A(n3101), .B(n842), .X(\update_mask_0/n1028 ) );
  nor_x1_sg U11141 ( .A(n834), .B(n839), .X(\update_mask_0/n1068 ) );
  nor_x1_sg U11142 ( .A(n3101), .B(n839), .X(\update_mask_0/n1060 ) );
  nor_x1_sg U11143 ( .A(n834), .B(n825), .X(\update_mask_0/n1004 ) );
  nor_x1_sg U11144 ( .A(n3101), .B(n825), .X(\update_mask_0/n996 ) );
  nor_x1_sg U11145 ( .A(n7401), .B(n815), .X(\update_output_0/n2504 ) );
  nor_x1_sg U11146 ( .A(n7402), .B(n815), .X(\update_output_0/n2503 ) );
  nor_x1_sg U11147 ( .A(n7336), .B(n815), .X(\update_output_0/n2500 ) );
  nor_x1_sg U11148 ( .A(n7337), .B(n815), .X(\update_output_0/n2499 ) );
  nor_x1_sg U11149 ( .A(n7335), .B(n815), .X(\update_output_0/n2496 ) );
  nor_x1_sg U11150 ( .A(n7339), .B(n815), .X(\update_output_0/n2495 ) );
  nor_x1_sg U11151 ( .A(n7334), .B(n815), .X(\update_output_0/n2492 ) );
  nor_x1_sg U11152 ( .A(n7341), .B(n815), .X(\update_output_0/n2491 ) );
  nor_x1_sg U11153 ( .A(n7333), .B(n815), .X(\update_output_0/n2488 ) );
  nor_x1_sg U11154 ( .A(n7401), .B(n800), .X(\update_output_0/n3144 ) );
  nor_x1_sg U11155 ( .A(n7402), .B(n800), .X(\update_output_0/n3143 ) );
  nor_x1_sg U11156 ( .A(n7336), .B(n800), .X(\update_output_0/n3140 ) );
  nor_x1_sg U11157 ( .A(n7337), .B(n800), .X(\update_output_0/n3139 ) );
  nor_x1_sg U11158 ( .A(n7335), .B(n800), .X(\update_output_0/n3136 ) );
  nor_x1_sg U11159 ( .A(n7339), .B(n800), .X(\update_output_0/n3135 ) );
  nor_x1_sg U11160 ( .A(n7334), .B(n800), .X(\update_output_0/n3132 ) );
  nor_x1_sg U11161 ( .A(n7341), .B(n800), .X(\update_output_0/n3131 ) );
  nor_x1_sg U11162 ( .A(n7333), .B(n800), .X(\update_output_0/n3128 ) );
  nand_x1_sg U11163 ( .A(n9187), .B(n9216), .X(n1555) );
  nand_x1_sg U11164 ( .A(n1558), .B(n9216), .X(n1574) );
  nand_x1_sg U11165 ( .A(n9188), .B(n9216), .X(n1548) );
  nand_x1_sg U11166 ( .A(n1537), .B(n9216), .X(n1540) );
  nand_x1_sg U11167 ( .A(n9187), .B(n9057), .X(n1551) );
  nand_x1_sg U11168 ( .A(n1558), .B(n9057), .X(n1573) );
  nand_x1_sg U11169 ( .A(n9188), .B(n9057), .X(n1545) );
  nand_x1_sg U11170 ( .A(n1537), .B(n9057), .X(n1546) );
  nand_x1_sg U11171 ( .A(n9187), .B(n9062), .X(n1561) );
  nand_x1_sg U11172 ( .A(n9187), .B(n9063), .X(n1563) );
  nand_x1_sg U11173 ( .A(n9187), .B(n9064), .X(n1554) );
  nand_x1_sg U11174 ( .A(n9187), .B(n9060), .X(n1550) );
  nand_x1_sg U11175 ( .A(n9187), .B(n9065), .X(n1562) );
  nand_x1_sg U11176 ( .A(n9187), .B(n9214), .X(n1560) );
  nand_x1_sg U11177 ( .A(n9188), .B(n9062), .X(n1556) );
  nand_x1_sg U11178 ( .A(n9188), .B(n9063), .X(n1566) );
  nand_x1_sg U11179 ( .A(n9188), .B(n9064), .X(n1547) );
  nand_x1_sg U11180 ( .A(n9188), .B(n9060), .X(n1544) );
  nand_x1_sg U11181 ( .A(n9188), .B(n9065), .X(n1541) );
  nand_x1_sg U11182 ( .A(n9188), .B(n9214), .X(n1542) );
  nand_x1_sg U11183 ( .A(n1558), .B(n9060), .X(n1572) );
  nand_x1_sg U11184 ( .A(n1537), .B(n9060), .X(n1543) );
  nand_x1_sg U11185 ( .A(n1558), .B(n9065), .X(n1557) );
  nand_x1_sg U11186 ( .A(n1537), .B(n9065), .X(n1549) );
  nand_x1_sg U11187 ( .A(n1558), .B(n9062), .X(n1569) );
  nand_x1_sg U11188 ( .A(n1558), .B(n9063), .X(n1571) );
  nand_x1_sg U11189 ( .A(n1558), .B(n9064), .X(n1570) );
  nand_x1_sg U11190 ( .A(n1558), .B(n9214), .X(n1559) );
  nand_x1_sg U11191 ( .A(n1537), .B(n9062), .X(n1538) );
  nand_x1_sg U11192 ( .A(n1537), .B(n9063), .X(n1539) );
  nand_x1_sg U11193 ( .A(n1537), .B(n9064), .X(n1536) );
  nand_x1_sg U11194 ( .A(n1537), .B(n9214), .X(n1552) );
  nor_x1_sg U11195 ( .A(n826), .B(n827), .X(\update_mask_0/n991 ) );
  nand_x4_sg U11196 ( .A(n7419), .B(n4391), .X(n4352) );
  nand_x1_sg U11197 ( .A(n4392), .B(n3099), .X(n4391) );
  nand_x4_sg U11198 ( .A(n7419), .B(n4349), .X(n4310) );
  nand_x1_sg U11199 ( .A(n4179), .B(n3099), .X(n4349) );
  nand_x4_sg U11200 ( .A(n1030), .B(n1031), .X(n777) );
  nor_x1_sg U11201 ( .A(n1032), .B(n1033), .X(n1031) );
  nor_x1_sg U11202 ( .A(n1040), .B(n1041), .X(n1030) );
  nand_x4_sg U11203 ( .A(n1233), .B(n1234), .X(n783) );
  nor_x1_sg U11204 ( .A(n1235), .B(n1236), .X(n1234) );
  nor_x1_sg U11205 ( .A(n1243), .B(n1244), .X(n1233) );
  nand_x4_sg U11206 ( .A(n852), .B(n853), .X(n793) );
  nor_x1_sg U11207 ( .A(n854), .B(n855), .X(n853) );
  nor_x1_sg U11208 ( .A(n867), .B(n868), .X(n852) );
  nand_x4_sg U11209 ( .A(n895), .B(n896), .X(n773) );
  nor_x1_sg U11210 ( .A(n897), .B(n898), .X(n896) );
  nor_x1_sg U11211 ( .A(n905), .B(n906), .X(n895) );
  nand_x4_sg U11212 ( .A(n1063), .B(n1064), .X(n778) );
  nor_x1_sg U11213 ( .A(n1065), .B(n1066), .X(n1064) );
  nor_x1_sg U11214 ( .A(n1073), .B(n1074), .X(n1063) );
  nand_x4_sg U11215 ( .A(n1200), .B(n1201), .X(n782) );
  nor_x1_sg U11216 ( .A(n1202), .B(n1203), .X(n1201) );
  nor_x1_sg U11217 ( .A(n1210), .B(n1211), .X(n1200) );
  nand_x4_sg U11218 ( .A(n1368), .B(n1369), .X(n787) );
  nor_x1_sg U11219 ( .A(n1370), .B(n1371), .X(n1369) );
  nor_x1_sg U11220 ( .A(n1378), .B(n1379), .X(n1368) );
  nand_x4_sg U11221 ( .A(n1401), .B(n1402), .X(n788) );
  nor_x1_sg U11222 ( .A(n1403), .B(n1404), .X(n1402) );
  nor_x1_sg U11223 ( .A(n1411), .B(n1412), .X(n1401) );
  nand_x4_sg U11224 ( .A(n7419), .B(n5053), .X(n4401) );
  nand_x1_sg U11225 ( .A(n4392), .B(n3096), .X(n5053) );
  nand_x4_sg U11226 ( .A(n7419), .B(n4178), .X(n4139) );
  nand_x1_sg U11227 ( .A(n4179), .B(n3096), .X(n4178) );
  nand_x2_sg U11228 ( .A(n886), .B(n887), .X(n885) );
  nand_x2_sg U11229 ( .A(n1055), .B(n1056), .X(n1054) );
  nand_x2_sg U11230 ( .A(n1088), .B(n1089), .X(n1087) );
  nand_x2_sg U11231 ( .A(n920), .B(n921), .X(n919) );
  nand_x2_sg U11232 ( .A(n1225), .B(n1226), .X(n1224) );
  nand_x2_sg U11233 ( .A(n1258), .B(n1259), .X(n1257) );
  nand_x2_sg U11234 ( .A(n1393), .B(n1394), .X(n1392) );
  nand_x2_sg U11235 ( .A(n1426), .B(n1427), .X(n1425) );
  nor_x1_sg U11236 ( .A(n963), .B(n964), .X(n962) );
  nor_x1_sg U11237 ( .A(n971), .B(n972), .X(n961) );
  nor_x1_sg U11238 ( .A(n996), .B(n997), .X(n995) );
  nor_x1_sg U11239 ( .A(n1004), .B(n1005), .X(n994) );
  nor_x1_sg U11240 ( .A(n1098), .B(n1099), .X(n1097) );
  nor_x1_sg U11241 ( .A(n1106), .B(n1107), .X(n1096) );
  nor_x1_sg U11242 ( .A(n1164), .B(n1165), .X(n1163) );
  nor_x1_sg U11243 ( .A(n1172), .B(n1173), .X(n1162) );
  nor_x1_sg U11244 ( .A(n1268), .B(n1269), .X(n1267) );
  nor_x1_sg U11245 ( .A(n1276), .B(n1277), .X(n1266) );
  nor_x1_sg U11246 ( .A(n1301), .B(n1302), .X(n1300) );
  nor_x1_sg U11247 ( .A(n1309), .B(n1310), .X(n1299) );
  nor_x1_sg U11248 ( .A(n1469), .B(n1470), .X(n1468) );
  nor_x1_sg U11249 ( .A(n1477), .B(n1478), .X(n1467) );
  nor_x1_sg U11250 ( .A(n1502), .B(n1503), .X(n1501) );
  nor_x1_sg U11251 ( .A(n1513), .B(n1514), .X(n1500) );
  nor_x1_sg U11252 ( .A(n930), .B(n931), .X(n929) );
  nor_x1_sg U11253 ( .A(n938), .B(n939), .X(n928) );
  nor_x1_sg U11254 ( .A(n1131), .B(n1132), .X(n1130) );
  nor_x1_sg U11255 ( .A(n1139), .B(n1140), .X(n1129) );
  nor_x1_sg U11256 ( .A(n1334), .B(n1335), .X(n1333) );
  nor_x1_sg U11257 ( .A(n1342), .B(n1343), .X(n1332) );
  nor_x1_sg U11258 ( .A(n1436), .B(n1437), .X(n1435) );
  nor_x1_sg U11259 ( .A(n1444), .B(n1445), .X(n1434) );
  nand_x2_sg U11260 ( .A(n953), .B(n954), .X(n952) );
  nand_x2_sg U11261 ( .A(n986), .B(n987), .X(n985) );
  nand_x2_sg U11262 ( .A(n1019), .B(n1020), .X(n1018) );
  nand_x2_sg U11263 ( .A(n1121), .B(n1122), .X(n1120) );
  nand_x2_sg U11264 ( .A(n1324), .B(n1325), .X(n1323) );
  nand_x2_sg U11265 ( .A(n1291), .B(n1292), .X(n1290) );
  nand_x2_sg U11266 ( .A(n1528), .B(n1529), .X(n1527) );
  nand_x2_sg U11267 ( .A(n1357), .B(n1358), .X(n1356) );
  nand_x2_sg U11268 ( .A(n1459), .B(n1460), .X(n1458) );
  nand_x2_sg U11269 ( .A(n1154), .B(n1155), .X(n1153) );
  nand_x2_sg U11270 ( .A(n1187), .B(n1188), .X(n1186) );
  nand_x2_sg U11271 ( .A(n4674), .B(n4675), .X(n4673) );
  nand_x2_sg U11272 ( .A(n4716), .B(n4717), .X(n4715) );
  nand_x2_sg U11273 ( .A(n4630), .B(n4631), .X(n4629) );
  nand_x2_sg U11274 ( .A(n4588), .B(n4589), .X(n4587) );
  nand_x2_sg U11275 ( .A(n4926), .B(n4927), .X(n4925) );
  nand_x2_sg U11276 ( .A(n4842), .B(n4843), .X(n4841) );
  nand_x2_sg U11277 ( .A(n4884), .B(n4885), .X(n4883) );
  nand_x2_sg U11278 ( .A(n4758), .B(n4759), .X(n4757) );
  nand_x2_sg U11279 ( .A(n4800), .B(n4801), .X(n4799) );
  nand_x2_sg U11280 ( .A(n4546), .B(n4547), .X(n4545) );
  nand_x2_sg U11281 ( .A(n4504), .B(n4505), .X(n4503) );
  nand_x2_sg U11282 ( .A(n4409), .B(n4410), .X(n4408) );
  nand_x2_sg U11283 ( .A(n4462), .B(n4463), .X(n4461) );
  nand_x2_sg U11284 ( .A(n5230), .B(n5231), .X(n5229) );
  nand_x2_sg U11285 ( .A(n4968), .B(n4969), .X(n4967) );
  nand_x2_sg U11286 ( .A(n5154), .B(n5155), .X(n5153) );
  nand_x2_sg U11287 ( .A(n5194), .B(n5195), .X(n5193) );
  nand_x2_sg U11288 ( .A(n5118), .B(n5119), .X(n5117) );
  nand_x2_sg U11289 ( .A(n5082), .B(n5083), .X(n5081) );
  nor_x1_sg U11290 ( .A(n5250), .B(n5251), .X(n5249) );
  nor_x1_sg U11291 ( .A(n5254), .B(n5255), .X(n5248) );
  nor_x1_sg U11292 ( .A(n4479), .B(n4480), .X(n4478) );
  nor_x1_sg U11293 ( .A(n4483), .B(n4484), .X(n4477) );
  nor_x1_sg U11294 ( .A(n4733), .B(n4734), .X(n4732) );
  nor_x1_sg U11295 ( .A(n4737), .B(n4738), .X(n4731) );
  nor_x1_sg U11296 ( .A(n4605), .B(n4606), .X(n4604) );
  nor_x1_sg U11297 ( .A(n4609), .B(n4610), .X(n4603) );
  nor_x1_sg U11298 ( .A(n4985), .B(n4986), .X(n4984) );
  nor_x1_sg U11299 ( .A(n4989), .B(n4990), .X(n4983) );
  nor_x1_sg U11300 ( .A(n4859), .B(n4860), .X(n4858) );
  nor_x1_sg U11301 ( .A(n4863), .B(n4864), .X(n4857) );
  nor_x1_sg U11302 ( .A(n4563), .B(n4564), .X(n4562) );
  nor_x1_sg U11303 ( .A(n4567), .B(n4568), .X(n4561) );
  nor_x1_sg U11304 ( .A(n4521), .B(n4522), .X(n4520) );
  nor_x1_sg U11305 ( .A(n4525), .B(n4526), .X(n4519) );
  nor_x1_sg U11306 ( .A(n4432), .B(n4433), .X(n4431) );
  nor_x1_sg U11307 ( .A(n4438), .B(n4439), .X(n4430) );
  nor_x1_sg U11308 ( .A(n4691), .B(n4692), .X(n4690) );
  nor_x1_sg U11309 ( .A(n4695), .B(n4696), .X(n4689) );
  nor_x1_sg U11310 ( .A(n4647), .B(n4648), .X(n4646) );
  nor_x1_sg U11311 ( .A(n4651), .B(n4652), .X(n4645) );
  nor_x1_sg U11312 ( .A(n4943), .B(n4944), .X(n4942) );
  nor_x1_sg U11313 ( .A(n4947), .B(n4948), .X(n4941) );
  nor_x1_sg U11314 ( .A(n5171), .B(n5172), .X(n5170) );
  nor_x1_sg U11315 ( .A(n5175), .B(n5176), .X(n5169) );
  nor_x1_sg U11316 ( .A(n5099), .B(n5100), .X(n5098) );
  nor_x1_sg U11317 ( .A(n5103), .B(n5104), .X(n5097) );
  nor_x1_sg U11318 ( .A(n4901), .B(n4902), .X(n4900) );
  nor_x1_sg U11319 ( .A(n4905), .B(n4906), .X(n4899) );
  nor_x1_sg U11320 ( .A(n4775), .B(n4776), .X(n4774) );
  nor_x1_sg U11321 ( .A(n4779), .B(n4780), .X(n4773) );
  nor_x1_sg U11322 ( .A(n4817), .B(n4818), .X(n4816) );
  nor_x1_sg U11323 ( .A(n4821), .B(n4822), .X(n4815) );
  nor_x1_sg U11324 ( .A(n5211), .B(n5212), .X(n5210) );
  nor_x1_sg U11325 ( .A(n5215), .B(n5216), .X(n5209) );
  nor_x1_sg U11326 ( .A(n5135), .B(n5136), .X(n5134) );
  nor_x1_sg U11327 ( .A(n5139), .B(n5140), .X(n5133) );
  nand_x2_sg U11328 ( .A(n5259), .B(n5260), .X(n5258) );
  nand_x2_sg U11329 ( .A(n5144), .B(n5145), .X(n5143) );
  nand_x2_sg U11330 ( .A(n5108), .B(n5109), .X(n5107) );
  nand_x2_sg U11331 ( .A(n5010), .B(n5011), .X(n5009) );
  nand_x2_sg U11332 ( .A(n5180), .B(n5181), .X(n5179) );
  nor_x1_sg U11333 ( .A(n5027), .B(n5028), .X(n5026) );
  nor_x1_sg U11334 ( .A(n5031), .B(n5032), .X(n5025) );
  nand_x2_sg U11335 ( .A(n5220), .B(n5221), .X(n5219) );
  nand_x2_sg U11336 ( .A(n5036), .B(n5037), .X(n5035) );
  nand_x2_sg U11337 ( .A(n4742), .B(n4743), .X(n4741) );
  nand_x2_sg U11338 ( .A(n4952), .B(n4953), .X(n4951) );
  nand_x2_sg U11339 ( .A(n4994), .B(n4995), .X(n4993) );
  nand_x2_sg U11340 ( .A(n4868), .B(n4869), .X(n4867) );
  nand_x2_sg U11341 ( .A(n4910), .B(n4911), .X(n4909) );
  nand_x2_sg U11342 ( .A(n4784), .B(n4785), .X(n4783) );
  nand_x2_sg U11343 ( .A(n4826), .B(n4827), .X(n4825) );
  nand_x2_sg U11344 ( .A(n4700), .B(n4701), .X(n4699) );
  nand_x2_sg U11345 ( .A(n4572), .B(n4573), .X(n4571) );
  nand_x2_sg U11346 ( .A(n4443), .B(n4444), .X(n4442) );
  nand_x2_sg U11347 ( .A(n4488), .B(n4489), .X(n4487) );
  nand_x2_sg U11348 ( .A(n4614), .B(n4615), .X(n4613) );
  nand_x2_sg U11349 ( .A(n4656), .B(n4657), .X(n4655) );
  nand_x2_sg U11350 ( .A(n4530), .B(n4531), .X(n4529) );
  nor_x1_sg U11351 ( .A(n4298), .B(n9190), .X(n4295) );
  nor_x1_sg U11352 ( .A(n4297), .B(n7526), .X(n4296) );
  nand_x1_sg U11353 ( .A(n4293), .B(n4017), .X(n4292) );
  nor_x1_sg U11354 ( .A(n3092), .B(n7559), .X(n4293) );
  nand_x1_sg U11355 ( .A(n3808), .B(n3809), .X(n3807) );
  nor_x1_sg U11356 ( .A(n5925), .B(n3820), .X(\update_mask_0/n1127 ) );
  nand_x2_sg U11357 ( .A(n9203), .B(n9219), .X(n5293) );
  nand_x1_sg U11358 ( .A(n9203), .B(n9217), .X(n5276) );
  nor_x1_sg U11359 ( .A(n9217), .B(n5274), .X(n5272) );
  nand_x1_sg U11360 ( .A(n9203), .B(n9215), .X(n5298) );
  nor_x1_sg U11361 ( .A(n5290), .B(n9219), .X(n5294) );
  nand_x1_sg U11362 ( .A(n9211), .B(n9210), .X(n5321) );
  nor_x1_sg U11363 ( .A(n7520), .B(n9186), .X(n1565) );
  nor_x1_sg U11364 ( .A(n9186), .B(n7519), .X(n1568) );
  nand_x1_sg U11365 ( .A(n2013), .B(n9217), .X(n1996) );
  nor_x1_sg U11366 ( .A(n2016), .B(n2017), .X(n2015) );
  nor_x1_sg U11367 ( .A(n2022), .B(n2023), .X(n2014) );
  nand_x2_sg U11368 ( .A(n1577), .B(n1578), .X(n1576) );
  nor_x1_sg U11369 ( .A(n1743), .B(n1744), .X(n1577) );
  nor_x1_sg U11370 ( .A(n1579), .B(n1580), .X(n1578) );
  nor_x1_sg U11371 ( .A(n831), .B(n829), .X(\update_mask_0/n1112 ) );
  nor_x1_sg U11372 ( .A(n832), .B(n829), .X(\update_mask_0/n1108 ) );
  nor_x1_sg U11373 ( .A(n831), .B(n839), .X(\update_mask_0/n1080 ) );
  nor_x1_sg U11374 ( .A(n832), .B(n839), .X(\update_mask_0/n1076 ) );
  nor_x1_sg U11375 ( .A(n831), .B(n842), .X(\update_mask_0/n1048 ) );
  nor_x1_sg U11376 ( .A(n832), .B(n842), .X(\update_mask_0/n1044 ) );
  nor_x1_sg U11377 ( .A(n831), .B(n825), .X(\update_mask_0/n1016 ) );
  nor_x1_sg U11378 ( .A(n832), .B(n825), .X(\update_mask_0/n1012 ) );
  nor_x1_sg U11379 ( .A(n830), .B(n829), .X(\update_mask_0/n1116 ) );
  nor_x1_sg U11380 ( .A(n830), .B(n839), .X(\update_mask_0/n1084 ) );
  nor_x1_sg U11381 ( .A(n830), .B(n842), .X(\update_mask_0/n1052 ) );
  nor_x1_sg U11382 ( .A(n830), .B(n825), .X(\update_mask_0/n1020 ) );
  nor_x1_sg U11383 ( .A(n833), .B(n829), .X(\update_mask_0/n1104 ) );
  nor_x1_sg U11384 ( .A(n835), .B(n829), .X(\update_mask_0/n1096 ) );
  nor_x1_sg U11385 ( .A(n833), .B(n842), .X(\update_mask_0/n1040 ) );
  nor_x1_sg U11386 ( .A(n835), .B(n842), .X(\update_mask_0/n1032 ) );
  nand_x2_sg U11387 ( .A(n1611), .B(n1612), .X(n1610) );
  nand_x1_sg U11388 ( .A(n9074), .B(n1613), .X(n1612) );
  nand_x1_sg U11389 ( .A(n9073), .B(n1617), .X(n1611) );
  nand_x2_sg U11390 ( .A(n1774), .B(n1775), .X(n1773) );
  nand_x1_sg U11391 ( .A(n9074), .B(n1776), .X(n1775) );
  nand_x1_sg U11392 ( .A(n9073), .B(n1780), .X(n1774) );
  nand_x2_sg U11393 ( .A(n1924), .B(n1925), .X(n1923) );
  nand_x1_sg U11394 ( .A(n9074), .B(n1926), .X(n1925) );
  nand_x1_sg U11395 ( .A(n9073), .B(n1930), .X(n1924) );
  nor_x1_sg U11396 ( .A(n1815), .B(n1816), .X(n1814) );
  nand_x2_sg U11397 ( .A(n1820), .B(n9048), .X(n1817) );
  nand_x2_sg U11398 ( .A(n1599), .B(n1600), .X(n1586) );
  nand_x1_sg U11399 ( .A(n9075), .B(n1601), .X(n1600) );
  nand_x1_sg U11400 ( .A(n9076), .B(n1605), .X(n1599) );
  nand_x2_sg U11401 ( .A(n1762), .B(n1763), .X(n1750) );
  nand_x1_sg U11402 ( .A(n9075), .B(n1764), .X(n1763) );
  nand_x1_sg U11403 ( .A(n9076), .B(n1768), .X(n1762) );
  nand_x2_sg U11404 ( .A(n1912), .B(n1913), .X(n1900) );
  nand_x1_sg U11405 ( .A(n9075), .B(n1914), .X(n1913) );
  nand_x1_sg U11406 ( .A(n9076), .B(n1918), .X(n1912) );
  nor_x1_sg U11407 ( .A(n9058), .B(n2059), .X(n2050) );
  nand_x2_sg U11408 ( .A(n1621), .B(n1622), .X(n1609) );
  nand_x1_sg U11409 ( .A(n1623), .B(n1624), .X(n1622) );
  nand_x1_sg U11410 ( .A(n9212), .B(n1628), .X(n1621) );
  nand_x2_sg U11411 ( .A(n1784), .B(n1785), .X(n1772) );
  nand_x1_sg U11412 ( .A(n1623), .B(n1786), .X(n1785) );
  nand_x1_sg U11413 ( .A(n9212), .B(n1790), .X(n1784) );
  nand_x2_sg U11414 ( .A(n1934), .B(n1935), .X(n1922) );
  nand_x1_sg U11415 ( .A(n1623), .B(n1936), .X(n1935) );
  nand_x1_sg U11416 ( .A(n9212), .B(n1940), .X(n1934) );
  nor_x1_sg U11417 ( .A(n833), .B(n839), .X(\update_mask_0/n1072 ) );
  nor_x1_sg U11418 ( .A(n835), .B(n839), .X(\update_mask_0/n1064 ) );
  nor_x1_sg U11419 ( .A(n833), .B(n825), .X(\update_mask_0/n1008 ) );
  nor_x1_sg U11420 ( .A(n835), .B(n825), .X(\update_mask_0/n1000 ) );
  nand_x4_sg U11421 ( .A(n1993), .B(n1994), .X(n827) );
  nand_x1_sg U11422 ( .A(n7519), .B(n2028), .X(n1993) );
  nor_x1_sg U11423 ( .A(n1657), .B(n1658), .X(n1633) );
  nand_x2_sg U11424 ( .A(n1669), .B(n1670), .X(n1657) );
  nand_x2_sg U11425 ( .A(n1659), .B(n1660), .X(n1658) );
  nand_x1_sg U11426 ( .A(n1623), .B(n1671), .X(n1670) );
  nor_x1_sg U11427 ( .A(n1721), .B(n1722), .X(n1697) );
  nand_x2_sg U11428 ( .A(n1733), .B(n1734), .X(n1721) );
  nand_x2_sg U11429 ( .A(n1723), .B(n1724), .X(n1722) );
  nand_x1_sg U11430 ( .A(n1623), .B(n1735), .X(n1734) );
  nor_x1_sg U11431 ( .A(n1801), .B(n1802), .X(n1796) );
  nand_x2_sg U11432 ( .A(n1803), .B(n1804), .X(n1802) );
  nand_x2_sg U11433 ( .A(n1807), .B(n1808), .X(n1806) );
  nor_x1_sg U11434 ( .A(n1970), .B(n1971), .X(n1945) );
  nand_x2_sg U11435 ( .A(n1982), .B(n1983), .X(n1970) );
  nand_x2_sg U11436 ( .A(n1972), .B(n1973), .X(n1971) );
  nand_x1_sg U11437 ( .A(n1623), .B(n1984), .X(n1983) );
  nor_x1_sg U11438 ( .A(n1635), .B(n1636), .X(n1634) );
  nand_x2_sg U11439 ( .A(n1637), .B(n1638), .X(n1636) );
  nand_x2_sg U11440 ( .A(n1647), .B(n1648), .X(n1635) );
  nor_x1_sg U11441 ( .A(n1699), .B(n1700), .X(n1698) );
  nand_x2_sg U11442 ( .A(n1701), .B(n1702), .X(n1700) );
  nand_x2_sg U11443 ( .A(n1711), .B(n1712), .X(n1699) );
  nor_x1_sg U11444 ( .A(n1947), .B(n1948), .X(n1946) );
  nand_x2_sg U11445 ( .A(n1949), .B(n1950), .X(n1948) );
  nand_x2_sg U11446 ( .A(n1959), .B(n1960), .X(n1947) );
  nand_x1_sg U11447 ( .A(n824), .B(n3100), .X(n823) );
  nor_x1_sg U11448 ( .A(n2034), .B(n2035), .X(n2033) );
  nor_x1_sg U11449 ( .A(n2042), .B(n2043), .X(n2032) );
  nand_x2_sg U11450 ( .A(n2036), .B(n2037), .X(n2035) );
  nor_x1_sg U11451 ( .A(n1586), .B(n1587), .X(n1585) );
  nor_x1_sg U11452 ( .A(n1609), .B(n1610), .X(n1584) );
  nand_x2_sg U11453 ( .A(n1588), .B(n1589), .X(n1587) );
  nor_x1_sg U11454 ( .A(n1684), .B(n1685), .X(n1683) );
  nor_x1_sg U11455 ( .A(n1690), .B(n1691), .X(n1682) );
  nand_x2_sg U11456 ( .A(n1686), .B(n1687), .X(n1685) );
  nor_x1_sg U11457 ( .A(n1750), .B(n1751), .X(n1749) );
  nor_x1_sg U11458 ( .A(n1772), .B(n1773), .X(n1748) );
  nand_x2_sg U11459 ( .A(n1752), .B(n1753), .X(n1751) );
  nor_x1_sg U11460 ( .A(n1900), .B(n1901), .X(n1899) );
  nor_x1_sg U11461 ( .A(n1922), .B(n1923), .X(n1898) );
  nand_x2_sg U11462 ( .A(n1902), .B(n1903), .X(n1901) );
  nor_x1_sg U11463 ( .A(n1825), .B(n1826), .X(n1813) );
  nand_x1_sg U11464 ( .A(\o_im[8][0] ), .B(n7495), .X(n4387) );
  nand_x1_sg U11465 ( .A(\o_im[8][2] ), .B(n7495), .X(n4363) );
  nand_x1_sg U11466 ( .A(\o_im[8][3] ), .B(n7408), .X(n4359) );
  nand_x1_sg U11467 ( .A(\o_im[8][4] ), .B(n7408), .X(n4371) );
  nand_x1_sg U11468 ( .A(\o_im[8][6] ), .B(n7495), .X(n4357) );
  nand_x1_sg U11469 ( .A(\o_im[8][7] ), .B(n7408), .X(n4383) );
  nand_x1_sg U11470 ( .A(\o_im[8][8] ), .B(n7408), .X(n4353) );
  nand_x1_sg U11471 ( .A(\o_im[8][9] ), .B(n7495), .X(n4381) );
  nand_x1_sg U11472 ( .A(\o_im[8][12] ), .B(n7408), .X(n4365) );
  nand_x1_sg U11473 ( .A(\o_im[8][13] ), .B(n7495), .X(n4375) );
  nand_x1_sg U11474 ( .A(\o_im[8][15] ), .B(n7408), .X(n4377) );
  nand_x1_sg U11475 ( .A(\o_im[8][16] ), .B(n7495), .X(n4350) );
  nand_x1_sg U11476 ( .A(\o_im[8][17] ), .B(n7495), .X(n4369) );
  nand_x1_sg U11477 ( .A(\o_im[8][18] ), .B(n7408), .X(n4389) );
  nand_x1_sg U11478 ( .A(\o_im[12][0] ), .B(n7498), .X(n4315) );
  nand_x1_sg U11479 ( .A(\o_im[12][1] ), .B(n7409), .X(n4323) );
  nand_x1_sg U11480 ( .A(\o_im[12][2] ), .B(n7409), .X(n4317) );
  nand_x1_sg U11481 ( .A(\o_im[12][3] ), .B(n7498), .X(n4327) );
  nand_x1_sg U11482 ( .A(\o_im[12][5] ), .B(n7498), .X(n4308) );
  nand_x1_sg U11483 ( .A(\o_im[12][6] ), .B(n7409), .X(n4329) );
  nand_x1_sg U11484 ( .A(\o_im[12][7] ), .B(n7498), .X(n4339) );
  nand_x1_sg U11485 ( .A(\o_im[12][8] ), .B(n7409), .X(n4341) );
  nand_x1_sg U11486 ( .A(\o_im[12][12] ), .B(n7498), .X(n4321) );
  nand_x1_sg U11487 ( .A(\o_im[12][14] ), .B(n7409), .X(n4347) );
  nand_x1_sg U11488 ( .A(\o_im[12][15] ), .B(n7498), .X(n4333) );
  nand_x1_sg U11489 ( .A(\o_im[12][16] ), .B(n7409), .X(n4311) );
  nand_x1_sg U11490 ( .A(\o_im[12][18] ), .B(n7498), .X(n4345) );
  nand_x1_sg U11491 ( .A(\o_im[12][19] ), .B(n7409), .X(n4335) );
  nand_x2_sg U11492 ( .A(n892), .B(n893), .X(n867) );
  nand_x2_sg U11493 ( .A(n926), .B(n927), .X(n905) );
  nand_x2_sg U11494 ( .A(n1094), .B(n1095), .X(n1073) );
  nand_x2_sg U11495 ( .A(n1231), .B(n1232), .X(n1210) );
  nand_x2_sg U11496 ( .A(n1399), .B(n1400), .X(n1378) );
  nand_x2_sg U11497 ( .A(n1432), .B(n1433), .X(n1411) );
  nand_x2_sg U11498 ( .A(n1061), .B(n1062), .X(n1040) );
  nand_x2_sg U11499 ( .A(n1264), .B(n1265), .X(n1243) );
  nand_x1_sg U11500 ( .A(\o_im[8][1] ), .B(n7408), .X(n4385) );
  nand_x1_sg U11501 ( .A(\o_im[8][5] ), .B(n7495), .X(n4373) );
  nand_x1_sg U11502 ( .A(\o_im[8][10] ), .B(n7408), .X(n4361) );
  nand_x1_sg U11503 ( .A(\o_im[8][11] ), .B(n7495), .X(n4355) );
  nand_x1_sg U11504 ( .A(\o_im[8][14] ), .B(n7495), .X(n4367) );
  nand_x1_sg U11505 ( .A(\o_im[8][19] ), .B(n7495), .X(n4379) );
  nand_x1_sg U11506 ( .A(\o_im[12][4] ), .B(n7498), .X(n4313) );
  nand_x1_sg U11507 ( .A(\o_im[12][9] ), .B(n7409), .X(n4337) );
  nand_x1_sg U11508 ( .A(\o_im[12][10] ), .B(n7409), .X(n4319) );
  nand_x1_sg U11509 ( .A(\o_im[12][11] ), .B(n7409), .X(n4343) );
  nand_x1_sg U11510 ( .A(\o_im[12][13] ), .B(n7409), .X(n4331) );
  nand_x1_sg U11511 ( .A(\o_im[12][17] ), .B(n7409), .X(n4325) );
  nand_x1_sg U11512 ( .A(\o_im[9][5] ), .B(n7508), .X(n4058) );
  nand_x1_sg U11513 ( .A(\o_im[9][6] ), .B(n7508), .X(n4083) );
  nand_x1_sg U11514 ( .A(\o_im[9][7] ), .B(n7406), .X(n4085) );
  nand_x1_sg U11515 ( .A(\o_im[9][8] ), .B(n7406), .X(n4073) );
  nand_x1_sg U11516 ( .A(\o_im[9][17] ), .B(n7406), .X(n4067) );
  nand_x1_sg U11517 ( .A(\o_im[9][18] ), .B(n7508), .X(n4095) );
  nand_x1_sg U11518 ( .A(\o_im[13][5] ), .B(n7403), .X(n4665) );
  nand_x1_sg U11519 ( .A(\o_im[13][6] ), .B(n7420), .X(n4711) );
  nand_x1_sg U11520 ( .A(\o_im[13][8] ), .B(n7420), .X(n4583) );
  nand_x1_sg U11521 ( .A(\o_im[13][9] ), .B(n7403), .X(n4921) );
  nand_x1_sg U11522 ( .A(\o_im[13][15] ), .B(n7420), .X(n4837) );
  nand_x1_sg U11523 ( .A(\o_im[13][18] ), .B(n7403), .X(n4795) );
  nand_x1_sg U11524 ( .A(\o_im[9][1] ), .B(n7406), .X(n4061) );
  nand_x1_sg U11525 ( .A(\o_im[9][2] ), .B(n7406), .X(n4065) );
  nand_x1_sg U11526 ( .A(\o_im[9][4] ), .B(n7406), .X(n4077) );
  nand_x1_sg U11527 ( .A(\o_im[13][1] ), .B(n7403), .X(n4539) );
  nand_x1_sg U11528 ( .A(\o_im[13][3] ), .B(n7403), .X(n4405) );
  nand_x1_sg U11529 ( .A(\o_im[13][4] ), .B(n7420), .X(n4455) );
  nand_x1_sg U11530 ( .A(\o_im[9][0] ), .B(n7508), .X(n4071) );
  nand_x1_sg U11531 ( .A(\o_im[9][10] ), .B(n7406), .X(n4079) );
  nand_x1_sg U11532 ( .A(\o_im[9][12] ), .B(n7508), .X(n4089) );
  nand_x1_sg U11533 ( .A(\o_im[9][13] ), .B(n7406), .X(n4091) );
  nand_x1_sg U11534 ( .A(\o_im[9][19] ), .B(n7406), .X(n4097) );
  nand_x1_sg U11535 ( .A(\o_im[13][0] ), .B(n7403), .X(n5227) );
  nand_x1_sg U11536 ( .A(\o_im[13][10] ), .B(n7403), .X(n4961) );
  nand_x1_sg U11537 ( .A(\o_im[13][12] ), .B(n7403), .X(n5191) );
  nand_x1_sg U11538 ( .A(\o_im[13][13] ), .B(n7420), .X(n5115) );
  nand_x1_sg U11539 ( .A(\o_im[13][14] ), .B(n7403), .X(n5076) );
  nand_x1_sg U11540 ( .A(\o_im[0][5] ), .B(n7462), .X(n4663) );
  nand_x1_sg U11541 ( .A(\o_im[0][6] ), .B(n7407), .X(n4707) );
  nand_x1_sg U11542 ( .A(\o_im[0][8] ), .B(n7407), .X(n4579) );
  nand_x1_sg U11543 ( .A(\o_im[0][9] ), .B(n7462), .X(n4917) );
  nand_x1_sg U11544 ( .A(\o_im[0][15] ), .B(n7407), .X(n4833) );
  nand_x1_sg U11545 ( .A(\o_im[0][18] ), .B(n7462), .X(n4791) );
  nand_x1_sg U11546 ( .A(\o_im[4][5] ), .B(n7505), .X(n4137) );
  nand_x1_sg U11547 ( .A(\o_im[4][6] ), .B(n7410), .X(n4158) );
  nand_x1_sg U11548 ( .A(\o_im[4][7] ), .B(n7505), .X(n4168) );
  nand_x1_sg U11549 ( .A(\o_im[4][8] ), .B(n7410), .X(n4170) );
  nand_x1_sg U11550 ( .A(\o_im[4][15] ), .B(n7505), .X(n4162) );
  nand_x1_sg U11551 ( .A(\o_im[4][16] ), .B(n7410), .X(n4140) );
  nand_x1_sg U11552 ( .A(\o_im[4][18] ), .B(n7505), .X(n4174) );
  nand_x1_sg U11553 ( .A(\o_im[0][1] ), .B(n7462), .X(n4541) );
  nand_x1_sg U11554 ( .A(\o_im[0][3] ), .B(n7462), .X(n4399) );
  nand_x1_sg U11555 ( .A(\o_im[0][4] ), .B(n7407), .X(n4457) );
  nand_x1_sg U11556 ( .A(\o_im[4][1] ), .B(n7410), .X(n4152) );
  nand_x1_sg U11557 ( .A(\o_im[4][2] ), .B(n7410), .X(n4146) );
  nand_x1_sg U11558 ( .A(\o_im[4][3] ), .B(n7505), .X(n4156) );
  nand_x1_sg U11559 ( .A(\o_im[0][10] ), .B(n7407), .X(n4963) );
  nand_x1_sg U11560 ( .A(\o_im[0][11] ), .B(n7407), .X(n5051) );
  nand_x1_sg U11561 ( .A(\o_im[0][12] ), .B(n7407), .X(n5045) );
  nand_x1_sg U11562 ( .A(\o_im[0][13] ), .B(n7462), .X(n5049) );
  nand_x1_sg U11563 ( .A(\o_im[0][14] ), .B(n7462), .X(n5043) );
  nand_x1_sg U11564 ( .A(\o_im[4][0] ), .B(n7505), .X(n4144) );
  nand_x1_sg U11565 ( .A(\o_im[4][12] ), .B(n7505), .X(n4150) );
  nand_x1_sg U11566 ( .A(\o_im[4][14] ), .B(n7410), .X(n4176) );
  nand_x1_sg U11567 ( .A(\o_im[4][19] ), .B(n7410), .X(n4164) );
  nand_x1_sg U11568 ( .A(\o_im[9][3] ), .B(n7508), .X(n4075) );
  nand_x1_sg U11569 ( .A(\o_im[9][9] ), .B(n7406), .X(n4069) );
  nand_x1_sg U11570 ( .A(\o_im[9][11] ), .B(n7406), .X(n4087) );
  nand_x1_sg U11571 ( .A(\o_im[9][14] ), .B(n7406), .X(n4081) );
  nand_x1_sg U11572 ( .A(\o_im[9][15] ), .B(n7508), .X(n4093) );
  nand_x1_sg U11573 ( .A(\o_im[9][16] ), .B(n7406), .X(n4063) );
  nand_x1_sg U11574 ( .A(\o_im[13][2] ), .B(n7420), .X(n4497) );
  nand_x1_sg U11575 ( .A(\o_im[13][7] ), .B(n7420), .X(n4623) );
  nand_x1_sg U11576 ( .A(\o_im[13][11] ), .B(n7403), .X(n5151) );
  nand_x1_sg U11577 ( .A(\o_im[13][16] ), .B(n7403), .X(n4877) );
  nand_x1_sg U11578 ( .A(\o_im[13][17] ), .B(n7420), .X(n4753) );
  nand_x1_sg U11579 ( .A(\o_im[13][19] ), .B(n7403), .X(n5003) );
  nand_x1_sg U11580 ( .A(\o_im[0][0] ), .B(n7407), .X(n5047) );
  nand_x1_sg U11581 ( .A(\o_im[0][2] ), .B(n7407), .X(n4495) );
  nand_x1_sg U11582 ( .A(\o_im[0][7] ), .B(n7462), .X(n4625) );
  nand_x1_sg U11583 ( .A(\o_im[0][16] ), .B(n7407), .X(n4879) );
  nand_x1_sg U11584 ( .A(\o_im[0][17] ), .B(n7407), .X(n4749) );
  nand_x1_sg U11585 ( .A(\o_im[0][19] ), .B(n7407), .X(n5005) );
  nand_x1_sg U11586 ( .A(\o_im[4][4] ), .B(n7410), .X(n4142) );
  nand_x1_sg U11587 ( .A(\o_im[4][9] ), .B(n7505), .X(n4166) );
  nand_x1_sg U11588 ( .A(\o_im[4][10] ), .B(n7410), .X(n4148) );
  nand_x1_sg U11589 ( .A(\o_im[4][11] ), .B(n7505), .X(n4172) );
  nand_x1_sg U11590 ( .A(\o_im[4][13] ), .B(n7505), .X(n4160) );
  nand_x1_sg U11591 ( .A(\o_im[4][17] ), .B(n7505), .X(n4154) );
  nand_x2_sg U11592 ( .A(n1075), .B(n1076), .X(n1074) );
  nand_x1_sg U11593 ( .A(\i_im[11][6] ), .B(n7385), .X(n1076) );
  nand_x2_sg U11594 ( .A(n1082), .B(n1083), .X(n1081) );
  nor_x1_sg U11595 ( .A(n1217), .B(n1218), .X(n1216) );
  nand_x2_sg U11596 ( .A(n1219), .B(n1220), .X(n1218) );
  nor_x1_sg U11597 ( .A(n1385), .B(n1386), .X(n1384) );
  nand_x2_sg U11598 ( .A(n1387), .B(n1388), .X(n1386) );
  nor_x1_sg U11599 ( .A(n1250), .B(n1251), .X(n1249) );
  nand_x2_sg U11600 ( .A(n1252), .B(n1253), .X(n1251) );
  nand_x2_sg U11601 ( .A(n869), .B(n870), .X(n868) );
  nand_x1_sg U11602 ( .A(\i_im[11][0] ), .B(n7385), .X(n870) );
  nand_x2_sg U11603 ( .A(n907), .B(n908), .X(n906) );
  nand_x1_sg U11604 ( .A(\i_im[11][1] ), .B(n7384), .X(n908) );
  nand_x2_sg U11605 ( .A(n1212), .B(n1213), .X(n1211) );
  nand_x1_sg U11606 ( .A(\i_im[11][10] ), .B(n7384), .X(n1213) );
  nand_x2_sg U11607 ( .A(n1380), .B(n1381), .X(n1379) );
  nand_x1_sg U11608 ( .A(\i_im[11][15] ), .B(n7385), .X(n1381) );
  nand_x2_sg U11609 ( .A(n1042), .B(n1043), .X(n1041) );
  nand_x1_sg U11610 ( .A(\i_im[11][5] ), .B(n871), .X(n1043) );
  nand_x2_sg U11611 ( .A(n1245), .B(n1246), .X(n1244) );
  nand_x1_sg U11612 ( .A(\i_im[11][11] ), .B(n871), .X(n1246) );
  nand_x2_sg U11613 ( .A(n860), .B(n861), .X(n854) );
  nor_x1_sg U11614 ( .A(n863), .B(n864), .X(n860) );
  nand_x2_sg U11615 ( .A(n901), .B(n902), .X(n897) );
  nor_x1_sg U11616 ( .A(n903), .B(n904), .X(n901) );
  nand_x2_sg U11617 ( .A(n1069), .B(n1070), .X(n1065) );
  nor_x1_sg U11618 ( .A(n1071), .B(n1072), .X(n1069) );
  nand_x2_sg U11619 ( .A(n1206), .B(n1207), .X(n1202) );
  nor_x1_sg U11620 ( .A(n1208), .B(n1209), .X(n1206) );
  nand_x2_sg U11621 ( .A(n1374), .B(n1375), .X(n1370) );
  nor_x1_sg U11622 ( .A(n1376), .B(n1377), .X(n1374) );
  nand_x2_sg U11623 ( .A(n1036), .B(n1037), .X(n1032) );
  nor_x1_sg U11624 ( .A(n1038), .B(n1039), .X(n1036) );
  nand_x2_sg U11625 ( .A(n1239), .B(n1240), .X(n1235) );
  nor_x1_sg U11626 ( .A(n1241), .B(n1242), .X(n1239) );
  nand_x2_sg U11627 ( .A(n877), .B(n878), .X(n876) );
  nand_x2_sg U11628 ( .A(n914), .B(n915), .X(n913) );
  nand_x2_sg U11629 ( .A(n1049), .B(n1050), .X(n1048) );
  nor_x1_sg U11630 ( .A(n1418), .B(n1419), .X(n1417) );
  nand_x2_sg U11631 ( .A(n1420), .B(n1421), .X(n1419) );
  nand_x2_sg U11632 ( .A(n1413), .B(n1414), .X(n1412) );
  nand_x1_sg U11633 ( .A(\i_im[11][16] ), .B(n7384), .X(n1414) );
  nand_x2_sg U11634 ( .A(n1407), .B(n1408), .X(n1403) );
  nor_x1_sg U11635 ( .A(n1409), .B(n1410), .X(n1407) );
  nand_x1_sg U11636 ( .A(\o_im[6][0] ), .B(n7518), .X(n3862) );
  nand_x1_sg U11637 ( .A(\o_im[6][1] ), .B(n7518), .X(n3835) );
  nand_x1_sg U11638 ( .A(\o_im[6][2] ), .B(n7517), .X(n3883) );
  nand_x1_sg U11639 ( .A(\o_im[6][3] ), .B(n7517), .X(n3829) );
  nand_x1_sg U11640 ( .A(\o_im[6][4] ), .B(n7518), .X(n3880) );
  nand_x1_sg U11641 ( .A(\o_im[6][7] ), .B(n7518), .X(n3871) );
  nand_x1_sg U11642 ( .A(\o_im[6][9] ), .B(n7517), .X(n3874) );
  nand_x1_sg U11643 ( .A(\o_im[6][11] ), .B(n7517), .X(n3847) );
  nand_x1_sg U11644 ( .A(\o_im[6][13] ), .B(n7517), .X(n3856) );
  nand_x1_sg U11645 ( .A(\o_im[6][14] ), .B(n7518), .X(n3844) );
  nand_x1_sg U11646 ( .A(\o_im[6][15] ), .B(n7518), .X(n3853) );
  nand_x1_sg U11647 ( .A(\o_im[6][16] ), .B(n7517), .X(n3838) );
  nand_x1_sg U11648 ( .A(\o_im[6][17] ), .B(n7517), .X(n3865) );
  nand_x1_sg U11649 ( .A(\o_im[6][18] ), .B(n7518), .X(n3825) );
  nand_x1_sg U11650 ( .A(\o_im[7][1] ), .B(n7503), .X(n4229) );
  nand_x1_sg U11651 ( .A(\o_im[7][3] ), .B(n7504), .X(n4233) );
  nand_x1_sg U11652 ( .A(\o_im[7][4] ), .B(n7504), .X(n4245) );
  nand_x1_sg U11653 ( .A(\o_im[7][5] ), .B(n7503), .X(n4241) );
  nand_x1_sg U11654 ( .A(\o_im[7][6] ), .B(n7504), .X(n4227) );
  nand_x1_sg U11655 ( .A(\o_im[7][8] ), .B(n7504), .X(n4208) );
  nand_x1_sg U11656 ( .A(\o_im[7][9] ), .B(n7503), .X(n4247) );
  nand_x1_sg U11657 ( .A(\o_im[7][10] ), .B(n7503), .X(n4217) );
  nand_x1_sg U11658 ( .A(\o_im[7][11] ), .B(n7504), .X(n4215) );
  nand_x1_sg U11659 ( .A(\o_im[7][12] ), .B(n7503), .X(n4235) );
  nand_x1_sg U11660 ( .A(\o_im[7][13] ), .B(n7503), .X(n4211) );
  nand_x1_sg U11661 ( .A(\o_im[7][14] ), .B(n7504), .X(n4239) );
  nand_x1_sg U11662 ( .A(\o_im[7][15] ), .B(n7504), .X(n4221) );
  nand_x1_sg U11663 ( .A(\o_im[7][17] ), .B(n7503), .X(n4223) );
  nand_x1_sg U11664 ( .A(\o_im[2][0] ), .B(n7460), .X(n5056) );
  nand_x1_sg U11665 ( .A(\o_im[2][1] ), .B(n7461), .X(n4543) );
  nand_x1_sg U11666 ( .A(\o_im[2][3] ), .B(n7461), .X(n4402) );
  nand_x1_sg U11667 ( .A(\o_im[2][4] ), .B(n7460), .X(n4459) );
  nand_x1_sg U11668 ( .A(\o_im[2][5] ), .B(n7461), .X(n4667) );
  nand_x1_sg U11669 ( .A(\o_im[2][6] ), .B(n7460), .X(n4709) );
  nand_x1_sg U11670 ( .A(\o_im[2][8] ), .B(n7460), .X(n4581) );
  nand_x1_sg U11671 ( .A(\o_im[2][9] ), .B(n7461), .X(n4919) );
  nand_x1_sg U11672 ( .A(\o_im[2][10] ), .B(n7460), .X(n4965) );
  nand_x1_sg U11673 ( .A(\o_im[2][11] ), .B(n7461), .X(n5054) );
  nand_x1_sg U11674 ( .A(\o_im[2][12] ), .B(n7461), .X(n5060) );
  nand_x1_sg U11675 ( .A(\o_im[2][14] ), .B(n7460), .X(n5062) );
  nand_x1_sg U11676 ( .A(\o_im[2][15] ), .B(n7460), .X(n4835) );
  nand_x1_sg U11677 ( .A(\o_im[2][18] ), .B(n7461), .X(n4793) );
  nand_x1_sg U11678 ( .A(\o_im[3][1] ), .B(n7511), .X(n3996) );
  nand_x1_sg U11679 ( .A(\o_im[3][2] ), .B(n7511), .X(n4014) );
  nand_x1_sg U11680 ( .A(\o_im[3][3] ), .B(n7512), .X(n3988) );
  nand_x1_sg U11681 ( .A(\o_im[3][4] ), .B(n7512), .X(n3975) );
  nand_x1_sg U11682 ( .A(\o_im[3][5] ), .B(n7511), .X(n3990) );
  nand_x1_sg U11683 ( .A(\o_im[3][6] ), .B(n7512), .X(n3982) );
  nand_x1_sg U11684 ( .A(\o_im[3][7] ), .B(n7511), .X(n4008) );
  nand_x1_sg U11685 ( .A(\o_im[3][8] ), .B(n7511), .X(n4002) );
  nand_x1_sg U11686 ( .A(\o_im[3][9] ), .B(n7512), .X(n4012) );
  nand_x1_sg U11687 ( .A(\o_im[3][12] ), .B(n7511), .X(n3978) );
  nand_x1_sg U11688 ( .A(\o_im[3][13] ), .B(n7512), .X(n3994) );
  nand_x1_sg U11689 ( .A(\o_im[3][14] ), .B(n7511), .X(n3984) );
  nand_x1_sg U11690 ( .A(\o_im[3][17] ), .B(n7512), .X(n4006) );
  nand_x1_sg U11691 ( .A(\o_im[3][18] ), .B(n7512), .X(n4000) );
  nand_x1_sg U11692 ( .A(\o_im[6][5] ), .B(n3828), .X(n3850) );
  nand_x1_sg U11693 ( .A(\o_im[6][6] ), .B(n3828), .X(n3841) );
  nand_x1_sg U11694 ( .A(\o_im[6][8] ), .B(n3828), .X(n3859) );
  nand_x1_sg U11695 ( .A(\o_im[6][10] ), .B(n3828), .X(n3832) );
  nand_x1_sg U11696 ( .A(\o_im[6][12] ), .B(n3828), .X(n3868) );
  nand_x1_sg U11697 ( .A(\o_im[6][19] ), .B(n3828), .X(n3877) );
  nand_x2_sg U11698 ( .A(n856), .B(n857), .X(n855) );
  nand_x2_sg U11699 ( .A(n899), .B(n900), .X(n898) );
  nand_x2_sg U11700 ( .A(n1034), .B(n1035), .X(n1033) );
  nand_x2_sg U11701 ( .A(n1067), .B(n1068), .X(n1066) );
  nand_x2_sg U11702 ( .A(n1204), .B(n1205), .X(n1203) );
  nand_x2_sg U11703 ( .A(n1237), .B(n1238), .X(n1236) );
  nand_x2_sg U11704 ( .A(n1372), .B(n1373), .X(n1371) );
  nand_x1_sg U11705 ( .A(\o_im[7][0] ), .B(n4210), .X(n4213) );
  nand_x1_sg U11706 ( .A(\o_im[7][2] ), .B(n4210), .X(n4225) );
  nand_x1_sg U11707 ( .A(\o_im[7][7] ), .B(n4210), .X(n4219) );
  nand_x1_sg U11708 ( .A(\o_im[7][16] ), .B(n4210), .X(n4231) );
  nand_x1_sg U11709 ( .A(\o_im[7][18] ), .B(n4210), .X(n4237) );
  nand_x1_sg U11710 ( .A(\o_im[7][19] ), .B(n4210), .X(n4243) );
  nand_x1_sg U11711 ( .A(\o_im[2][2] ), .B(n4404), .X(n4499) );
  nand_x1_sg U11712 ( .A(\o_im[2][7] ), .B(n4404), .X(n4627) );
  nand_x1_sg U11713 ( .A(\o_im[2][13] ), .B(n4404), .X(n5058) );
  nand_x1_sg U11714 ( .A(\o_im[2][16] ), .B(n4404), .X(n4881) );
  nand_x1_sg U11715 ( .A(\o_im[2][17] ), .B(n4404), .X(n4751) );
  nand_x1_sg U11716 ( .A(\o_im[2][19] ), .B(n4404), .X(n5007) );
  nand_x1_sg U11717 ( .A(\o_im[3][0] ), .B(n3977), .X(n4004) );
  nand_x1_sg U11718 ( .A(\o_im[3][10] ), .B(n3977), .X(n3992) );
  nand_x1_sg U11719 ( .A(\o_im[3][11] ), .B(n3977), .X(n3986) );
  nand_x1_sg U11720 ( .A(\o_im[3][15] ), .B(n3977), .X(n3980) );
  nand_x1_sg U11721 ( .A(\o_im[3][16] ), .B(n3977), .X(n3998) );
  nand_x1_sg U11722 ( .A(\o_im[3][19] ), .B(n3977), .X(n4010) );
  nand_x2_sg U11723 ( .A(n1405), .B(n1406), .X(n1404) );
  nand_x1_sg U11724 ( .A(\o_im[14][0] ), .B(n7515), .X(n3926) );
  nand_x1_sg U11725 ( .A(\o_im[14][2] ), .B(n7516), .X(n3918) );
  nand_x1_sg U11726 ( .A(\o_im[14][3] ), .B(n7515), .X(n3890) );
  nand_x1_sg U11727 ( .A(\o_im[14][4] ), .B(n7516), .X(n3924) );
  nand_x1_sg U11728 ( .A(\o_im[14][5] ), .B(n7515), .X(n3896) );
  nand_x1_sg U11729 ( .A(\o_im[14][6] ), .B(n7515), .X(n3914) );
  nand_x1_sg U11730 ( .A(\o_im[14][7] ), .B(n7515), .X(n3908) );
  nand_x1_sg U11731 ( .A(\o_im[14][8] ), .B(n7516), .X(n3894) );
  nand_x1_sg U11732 ( .A(\o_im[14][9] ), .B(n7515), .X(n3920) );
  nand_x1_sg U11733 ( .A(\o_im[14][12] ), .B(n7516), .X(n3906) );
  nand_x1_sg U11734 ( .A(\o_im[14][13] ), .B(n7516), .X(n3900) );
  nand_x1_sg U11735 ( .A(\o_im[14][14] ), .B(n7515), .X(n3902) );
  nand_x1_sg U11736 ( .A(\o_im[14][16] ), .B(n7516), .X(n3912) );
  nand_x1_sg U11737 ( .A(\o_im[14][18] ), .B(n7516), .X(n3887) );
  nand_x1_sg U11738 ( .A(\o_im[15][0] ), .B(n7501), .X(n4265) );
  nand_x1_sg U11739 ( .A(\o_im[15][2] ), .B(n7501), .X(n4289) );
  nand_x1_sg U11740 ( .A(\o_im[15][3] ), .B(n7501), .X(n4277) );
  nand_x1_sg U11741 ( .A(\o_im[15][4] ), .B(n7502), .X(n4250) );
  nand_x1_sg U11742 ( .A(\o_im[15][6] ), .B(n7502), .X(n4257) );
  nand_x1_sg U11743 ( .A(\o_im[15][7] ), .B(n7501), .X(n4283) );
  nand_x1_sg U11744 ( .A(\o_im[15][9] ), .B(n7502), .X(n4287) );
  nand_x1_sg U11745 ( .A(\o_im[15][10] ), .B(n7502), .X(n4263) );
  nand_x1_sg U11746 ( .A(\o_im[15][12] ), .B(n7501), .X(n4253) );
  nand_x1_sg U11747 ( .A(\o_im[15][13] ), .B(n7501), .X(n4271) );
  nand_x1_sg U11748 ( .A(\o_im[15][14] ), .B(n7501), .X(n4259) );
  nand_x1_sg U11749 ( .A(\o_im[15][16] ), .B(n7502), .X(n4275) );
  nand_x1_sg U11750 ( .A(\o_im[15][17] ), .B(n7502), .X(n4281) );
  nand_x1_sg U11751 ( .A(\o_im[15][18] ), .B(n7502), .X(n4269) );
  nand_x1_sg U11752 ( .A(\o_im[10][0] ), .B(n7458), .X(n5067) );
  nand_x1_sg U11753 ( .A(\o_im[10][1] ), .B(n7459), .X(n4537) );
  nand_x1_sg U11754 ( .A(\o_im[10][3] ), .B(n7459), .X(n4396) );
  nand_x1_sg U11755 ( .A(\o_im[10][4] ), .B(n7458), .X(n4453) );
  nand_x1_sg U11756 ( .A(\o_im[10][5] ), .B(n7459), .X(n4671) );
  nand_x1_sg U11757 ( .A(\o_im[10][6] ), .B(n7458), .X(n4713) );
  nand_x1_sg U11758 ( .A(\o_im[10][8] ), .B(n7458), .X(n4585) );
  nand_x1_sg U11759 ( .A(\o_im[10][9] ), .B(n7459), .X(n4923) );
  nand_x1_sg U11760 ( .A(\o_im[10][10] ), .B(n7458), .X(n4959) );
  nand_x1_sg U11761 ( .A(\o_im[10][11] ), .B(n7458), .X(n5073) );
  nand_x1_sg U11762 ( .A(\o_im[10][12] ), .B(n7459), .X(n5065) );
  nand_x1_sg U11763 ( .A(\o_im[10][14] ), .B(n7459), .X(n5071) );
  nand_x1_sg U11764 ( .A(\o_im[10][15] ), .B(n7458), .X(n4839) );
  nand_x1_sg U11765 ( .A(\o_im[10][18] ), .B(n7459), .X(n4797) );
  nand_x1_sg U11766 ( .A(\o_im[11][0] ), .B(n7514), .X(n3940) );
  nand_x1_sg U11767 ( .A(\o_im[11][1] ), .B(n7513), .X(n3942) );
  nand_x1_sg U11768 ( .A(\o_im[11][2] ), .B(n7513), .X(n3936) );
  nand_x1_sg U11769 ( .A(\o_im[11][4] ), .B(n7514), .X(n3970) );
  nand_x1_sg U11770 ( .A(\o_im[11][5] ), .B(n7513), .X(n3954) );
  nand_x1_sg U11771 ( .A(\o_im[11][6] ), .B(n7514), .X(n3933) );
  nand_x1_sg U11772 ( .A(\o_im[11][7] ), .B(n7513), .X(n3960) );
  nand_x1_sg U11773 ( .A(\o_im[11][8] ), .B(n7514), .X(n3964) );
  nand_x1_sg U11774 ( .A(\o_im[11][9] ), .B(n7513), .X(n3966) );
  nand_x1_sg U11775 ( .A(\o_im[11][10] ), .B(n7514), .X(n3952) );
  nand_x1_sg U11776 ( .A(\o_im[11][12] ), .B(n7514), .X(n3958) );
  nand_x1_sg U11777 ( .A(\o_im[11][13] ), .B(n7513), .X(n3948) );
  nand_x1_sg U11778 ( .A(\o_im[11][14] ), .B(n7513), .X(n3972) );
  nand_x1_sg U11779 ( .A(\o_im[11][18] ), .B(n7514), .X(n3946) );
  nand_x1_sg U11780 ( .A(\o_im[14][1] ), .B(n3889), .X(n3910) );
  nand_x1_sg U11781 ( .A(\o_im[14][10] ), .B(n3889), .X(n3892) );
  nand_x1_sg U11782 ( .A(\o_im[14][11] ), .B(n3889), .X(n3916) );
  nand_x1_sg U11783 ( .A(\o_im[14][15] ), .B(n3889), .X(n3898) );
  nand_x1_sg U11784 ( .A(\o_im[14][17] ), .B(n3889), .X(n3904) );
  nand_x1_sg U11785 ( .A(\o_im[14][19] ), .B(n3889), .X(n3922) );
  nand_x1_sg U11786 ( .A(\o_im[15][1] ), .B(n4252), .X(n4273) );
  nand_x1_sg U11787 ( .A(\o_im[15][5] ), .B(n4252), .X(n4267) );
  nand_x1_sg U11788 ( .A(\o_im[15][8] ), .B(n4252), .X(n4279) );
  nand_x1_sg U11789 ( .A(\o_im[15][11] ), .B(n4252), .X(n4261) );
  nand_x1_sg U11790 ( .A(\o_im[15][15] ), .B(n4252), .X(n4255) );
  nand_x1_sg U11791 ( .A(\o_im[15][19] ), .B(n4252), .X(n4285) );
  nand_x1_sg U11792 ( .A(\o_im[10][2] ), .B(n4398), .X(n4501) );
  nand_x1_sg U11793 ( .A(\o_im[10][7] ), .B(n4398), .X(n4621) );
  nand_x1_sg U11794 ( .A(\o_im[10][13] ), .B(n4398), .X(n5069) );
  nand_x1_sg U11795 ( .A(\o_im[10][16] ), .B(n4398), .X(n4875) );
  nand_x1_sg U11796 ( .A(\o_im[10][17] ), .B(n4398), .X(n4755) );
  nand_x1_sg U11797 ( .A(\o_im[10][19] ), .B(n4398), .X(n5001) );
  nand_x1_sg U11798 ( .A(\o_im[11][3] ), .B(n3935), .X(n3962) );
  nand_x1_sg U11799 ( .A(\o_im[11][11] ), .B(n3935), .X(n3950) );
  nand_x1_sg U11800 ( .A(\o_im[11][15] ), .B(n3935), .X(n3938) );
  nand_x1_sg U11801 ( .A(\o_im[11][16] ), .B(n3935), .X(n3944) );
  nand_x1_sg U11802 ( .A(\o_im[11][17] ), .B(n3935), .X(n3956) );
  nand_x1_sg U11803 ( .A(\o_im[11][19] ), .B(n3935), .X(n3968) );
  nand_x1_sg U11804 ( .A(\o_im[5][6] ), .B(n7404), .X(n4052) );
  nand_x1_sg U11805 ( .A(\o_im[5][8] ), .B(n7446), .X(n4044) );
  nand_x1_sg U11806 ( .A(\o_im[5][9] ), .B(n7446), .X(n4038) );
  nand_x1_sg U11807 ( .A(\o_im[5][18] ), .B(n7446), .X(n4032) );
  nand_x1_sg U11808 ( .A(\o_im[5][1] ), .B(n7446), .X(n4019) );
  nand_x1_sg U11809 ( .A(\o_im[5][2] ), .B(n7404), .X(n4040) );
  nand_x1_sg U11810 ( .A(\o_im[5][4] ), .B(n7404), .X(n4022) );
  nand_x1_sg U11811 ( .A(\o_im[5][0] ), .B(n7404), .X(n4056) );
  nand_x1_sg U11812 ( .A(\o_im[5][10] ), .B(n7446), .X(n4026) );
  nand_x1_sg U11813 ( .A(\o_im[5][11] ), .B(n7404), .X(n4046) );
  nand_x1_sg U11814 ( .A(\o_im[5][12] ), .B(n7404), .X(n5188) );
  nand_x1_sg U11815 ( .A(\o_im[5][13] ), .B(n7404), .X(n4028) );
  nand_x1_sg U11816 ( .A(\o_im[5][14] ), .B(n7404), .X(n4034) );
  nand_x1_sg U11817 ( .A(\o_im[5][19] ), .B(n7446), .X(n4050) );
  nand_x1_sg U11818 ( .A(\o_im[1][5] ), .B(n7405), .X(n4670) );
  nand_x1_sg U11819 ( .A(\o_im[1][6] ), .B(n7455), .X(n4116) );
  nand_x1_sg U11820 ( .A(\o_im[1][7] ), .B(n7455), .X(n4104) );
  nand_x1_sg U11821 ( .A(\o_im[1][16] ), .B(n7455), .X(n4110) );
  nand_x1_sg U11822 ( .A(\o_im[1][18] ), .B(n7405), .X(n4114) );
  nand_x1_sg U11823 ( .A(\o_im[1][1] ), .B(n7405), .X(n4101) );
  nand_x1_sg U11824 ( .A(\o_im[1][2] ), .B(n7455), .X(n4122) );
  nand_x1_sg U11825 ( .A(\o_im[1][3] ), .B(n7455), .X(n4128) );
  nand_x1_sg U11826 ( .A(\o_im[1][0] ), .B(n7405), .X(n4126) );
  nand_x1_sg U11827 ( .A(\o_im[1][10] ), .B(n7405), .X(n4108) );
  nand_x1_sg U11828 ( .A(\o_im[1][11] ), .B(n7405), .X(n4120) );
  nand_x1_sg U11829 ( .A(\o_im[1][12] ), .B(n7405), .X(n4132) );
  nand_x1_sg U11830 ( .A(\o_im[1][14] ), .B(n7455), .X(n5079) );
  nand_x1_sg U11831 ( .A(\o_im[1][19] ), .B(n7455), .X(n4134) );
  nand_x1_sg U11832 ( .A(\o_im[5][3] ), .B(n7404), .X(n4036) );
  nand_x1_sg U11833 ( .A(\o_im[5][5] ), .B(n7404), .X(n4042) );
  nand_x1_sg U11834 ( .A(\o_im[5][7] ), .B(n7446), .X(n4024) );
  nand_x1_sg U11835 ( .A(\o_im[5][15] ), .B(n7404), .X(n4054) );
  nand_x1_sg U11836 ( .A(\o_im[5][16] ), .B(n7446), .X(n4030) );
  nand_x1_sg U11837 ( .A(\o_im[5][17] ), .B(n7404), .X(n4048) );
  nand_x1_sg U11838 ( .A(\o_im[1][4] ), .B(n7405), .X(n4106) );
  nand_x1_sg U11839 ( .A(\o_im[1][8] ), .B(n7455), .X(n4136) );
  nand_x1_sg U11840 ( .A(\o_im[1][9] ), .B(n7405), .X(n4130) );
  nand_x1_sg U11841 ( .A(\o_im[1][13] ), .B(n7405), .X(n4112) );
  nand_x1_sg U11842 ( .A(\o_im[1][15] ), .B(n7405), .X(n4118) );
  nand_x1_sg U11843 ( .A(\o_im[1][17] ), .B(n7405), .X(n4124) );
  nand_x2_sg U11844 ( .A(n992), .B(n993), .X(n971) );
  nand_x2_sg U11845 ( .A(n1025), .B(n1026), .X(n1004) );
  nand_x2_sg U11846 ( .A(n1127), .B(n1128), .X(n1106) );
  nand_x2_sg U11847 ( .A(n1193), .B(n1194), .X(n1172) );
  nand_x2_sg U11848 ( .A(n1297), .B(n1298), .X(n1276) );
  nand_x2_sg U11849 ( .A(n1330), .B(n1331), .X(n1309) );
  nand_x2_sg U11850 ( .A(n1498), .B(n1499), .X(n1477) );
  nand_x2_sg U11851 ( .A(n1534), .B(n1535), .X(n1513) );
  nand_x2_sg U11852 ( .A(n959), .B(n960), .X(n938) );
  nand_x2_sg U11853 ( .A(n1160), .B(n1161), .X(n1139) );
  nand_x2_sg U11854 ( .A(n1363), .B(n1364), .X(n1342) );
  nand_x2_sg U11855 ( .A(n1465), .B(n1466), .X(n1444) );
  nor_x1_sg U11856 ( .A(n1011), .B(n1012), .X(n1010) );
  nand_x2_sg U11857 ( .A(n1013), .B(n1014), .X(n1012) );
  nor_x1_sg U11858 ( .A(n1520), .B(n1521), .X(n1519) );
  nand_x2_sg U11859 ( .A(n1522), .B(n1523), .X(n1521) );
  nor_x1_sg U11860 ( .A(n1349), .B(n1350), .X(n1348) );
  nand_x2_sg U11861 ( .A(n1351), .B(n1352), .X(n1350) );
  nand_x2_sg U11862 ( .A(n1006), .B(n1007), .X(n1005) );
  nand_x1_sg U11863 ( .A(\i_im[11][4] ), .B(n7384), .X(n1007) );
  nand_x2_sg U11864 ( .A(n1174), .B(n1175), .X(n1173) );
  nand_x1_sg U11865 ( .A(\i_im[11][9] ), .B(n7385), .X(n1175) );
  nand_x2_sg U11866 ( .A(n1311), .B(n1312), .X(n1310) );
  nand_x1_sg U11867 ( .A(\i_im[11][13] ), .B(n7384), .X(n1312) );
  nand_x2_sg U11868 ( .A(n1479), .B(n1480), .X(n1478) );
  nand_x1_sg U11869 ( .A(\i_im[11][18] ), .B(n7385), .X(n1480) );
  nand_x2_sg U11870 ( .A(n1515), .B(n1516), .X(n1514) );
  nand_x1_sg U11871 ( .A(\i_im[11][19] ), .B(n7384), .X(n1516) );
  nand_x2_sg U11872 ( .A(n940), .B(n941), .X(n939) );
  nand_x1_sg U11873 ( .A(\i_im[11][2] ), .B(n871), .X(n941) );
  nand_x2_sg U11874 ( .A(n1344), .B(n1345), .X(n1343) );
  nand_x1_sg U11875 ( .A(\i_im[11][14] ), .B(n871), .X(n1345) );
  nand_x2_sg U11876 ( .A(n1000), .B(n1001), .X(n996) );
  nor_x1_sg U11877 ( .A(n1002), .B(n1003), .X(n1000) );
  nand_x2_sg U11878 ( .A(n1168), .B(n1169), .X(n1164) );
  nor_x1_sg U11879 ( .A(n1170), .B(n1171), .X(n1168) );
  nand_x2_sg U11880 ( .A(n1305), .B(n1306), .X(n1301) );
  nor_x1_sg U11881 ( .A(n1307), .B(n1308), .X(n1305) );
  nand_x2_sg U11882 ( .A(n1473), .B(n1474), .X(n1469) );
  nor_x1_sg U11883 ( .A(n1475), .B(n1476), .X(n1473) );
  nand_x2_sg U11884 ( .A(n1506), .B(n1507), .X(n1502) );
  nor_x1_sg U11885 ( .A(n1508), .B(n1509), .X(n1506) );
  nand_x2_sg U11886 ( .A(n934), .B(n935), .X(n930) );
  nor_x1_sg U11887 ( .A(n936), .B(n937), .X(n934) );
  nand_x2_sg U11888 ( .A(n1338), .B(n1339), .X(n1334) );
  nor_x1_sg U11889 ( .A(n1340), .B(n1341), .X(n1338) );
  nand_x2_sg U11890 ( .A(n1181), .B(n1182), .X(n1180) );
  nand_x2_sg U11891 ( .A(n1318), .B(n1319), .X(n1317) );
  nand_x2_sg U11892 ( .A(n1486), .B(n1487), .X(n1485) );
  nand_x2_sg U11893 ( .A(n947), .B(n948), .X(n946) );
  nor_x1_sg U11894 ( .A(n978), .B(n979), .X(n977) );
  nand_x2_sg U11895 ( .A(n980), .B(n981), .X(n979) );
  nor_x1_sg U11896 ( .A(n1113), .B(n1114), .X(n1112) );
  nand_x2_sg U11897 ( .A(n1115), .B(n1116), .X(n1114) );
  nor_x1_sg U11898 ( .A(n1146), .B(n1147), .X(n1145) );
  nand_x2_sg U11899 ( .A(n1148), .B(n1149), .X(n1147) );
  nand_x2_sg U11900 ( .A(n973), .B(n974), .X(n972) );
  nand_x1_sg U11901 ( .A(\i_im[11][3] ), .B(n7385), .X(n974) );
  nand_x2_sg U11902 ( .A(n1108), .B(n1109), .X(n1107) );
  nand_x1_sg U11903 ( .A(\i_im[11][7] ), .B(n7384), .X(n1109) );
  nand_x2_sg U11904 ( .A(n1278), .B(n1279), .X(n1277) );
  nand_x1_sg U11905 ( .A(\i_im[11][12] ), .B(n7385), .X(n1279) );
  nand_x2_sg U11906 ( .A(n1141), .B(n1142), .X(n1140) );
  nand_x1_sg U11907 ( .A(\i_im[11][8] ), .B(n871), .X(n1142) );
  nand_x2_sg U11908 ( .A(n1285), .B(n1286), .X(n1284) );
  nor_x1_sg U11909 ( .A(n1451), .B(n1452), .X(n1450) );
  nand_x2_sg U11910 ( .A(n1453), .B(n1454), .X(n1452) );
  nand_x2_sg U11911 ( .A(n1446), .B(n1447), .X(n1445) );
  nand_x1_sg U11912 ( .A(\i_im[11][17] ), .B(n871), .X(n1447) );
  nand_x2_sg U11913 ( .A(n967), .B(n968), .X(n963) );
  nor_x1_sg U11914 ( .A(n969), .B(n970), .X(n967) );
  nand_x2_sg U11915 ( .A(n1102), .B(n1103), .X(n1098) );
  nor_x1_sg U11916 ( .A(n1104), .B(n1105), .X(n1102) );
  nand_x2_sg U11917 ( .A(n1272), .B(n1273), .X(n1268) );
  nor_x1_sg U11918 ( .A(n1274), .B(n1275), .X(n1272) );
  nand_x2_sg U11919 ( .A(n1135), .B(n1136), .X(n1131) );
  nor_x1_sg U11920 ( .A(n1137), .B(n1138), .X(n1135) );
  nand_x2_sg U11921 ( .A(n1440), .B(n1441), .X(n1436) );
  nor_x1_sg U11922 ( .A(n1442), .B(n1443), .X(n1440) );
  nand_x2_sg U11923 ( .A(n1492), .B(n1493), .X(n1491) );
  nand_x2_sg U11924 ( .A(n932), .B(n933), .X(n931) );
  nand_x2_sg U11925 ( .A(n998), .B(n999), .X(n997) );
  nand_x2_sg U11926 ( .A(n1166), .B(n1167), .X(n1165) );
  nand_x2_sg U11927 ( .A(n1303), .B(n1304), .X(n1302) );
  nand_x2_sg U11928 ( .A(n1336), .B(n1337), .X(n1335) );
  nand_x2_sg U11929 ( .A(n1471), .B(n1472), .X(n1470) );
  nand_x2_sg U11930 ( .A(n1504), .B(n1505), .X(n1503) );
  nand_x2_sg U11931 ( .A(n965), .B(n966), .X(n964) );
  nand_x2_sg U11932 ( .A(n1100), .B(n1101), .X(n1099) );
  nand_x2_sg U11933 ( .A(n1133), .B(n1134), .X(n1132) );
  nand_x2_sg U11934 ( .A(n1270), .B(n1271), .X(n1269) );
  nand_x2_sg U11935 ( .A(n1438), .B(n1439), .X(n1437) );
  nor_x1_sg U11936 ( .A(n1059), .B(n7566), .X(n1058) );
  nor_x1_sg U11937 ( .A(n1092), .B(n7566), .X(n1091) );
  nor_x1_sg U11938 ( .A(n1229), .B(n7564), .X(n1228) );
  nor_x1_sg U11939 ( .A(n1262), .B(n7566), .X(n1261) );
  nor_x1_sg U11940 ( .A(n924), .B(n7566), .X(n923) );
  nor_x1_sg U11941 ( .A(n1397), .B(n7566), .X(n1396) );
  nor_x1_sg U11942 ( .A(n1430), .B(n7566), .X(n1429) );
  nor_x1_sg U11943 ( .A(n890), .B(n7566), .X(n889) );
  nand_x2_sg U11944 ( .A(n5264), .B(n5265), .X(n5243) );
  nand_x2_sg U11945 ( .A(n5245), .B(n5246), .X(n5244) );
  nand_x1_sg U11946 ( .A(n7423), .B(n5537), .X(n5264) );
  nand_x2_sg U11947 ( .A(n4577), .B(n4578), .X(n4556) );
  nand_x2_sg U11948 ( .A(n4558), .B(n4559), .X(n4557) );
  nand_x1_sg U11949 ( .A(n7424), .B(n5526), .X(n4577) );
  nand_x2_sg U11950 ( .A(n4449), .B(n4450), .X(n4424) );
  nand_x2_sg U11951 ( .A(n4426), .B(n4427), .X(n4425) );
  nand_x1_sg U11952 ( .A(n7424), .B(n5504), .X(n4449) );
  nand_x2_sg U11953 ( .A(n4493), .B(n4494), .X(n4472) );
  nand_x2_sg U11954 ( .A(n4474), .B(n4475), .X(n4473) );
  nand_x1_sg U11955 ( .A(n7423), .B(n5493), .X(n4493) );
  nand_x2_sg U11956 ( .A(n4705), .B(n4706), .X(n4684) );
  nand_x2_sg U11957 ( .A(n4686), .B(n4687), .X(n4685) );
  nand_x1_sg U11958 ( .A(n7424), .B(n5482), .X(n4705) );
  nand_x2_sg U11959 ( .A(n4747), .B(n4748), .X(n4726) );
  nand_x2_sg U11960 ( .A(n4728), .B(n4729), .X(n4727) );
  nand_x1_sg U11961 ( .A(n7423), .B(n5471), .X(n4747) );
  nand_x2_sg U11962 ( .A(n4619), .B(n4620), .X(n4598) );
  nand_x2_sg U11963 ( .A(n4600), .B(n4601), .X(n4599) );
  nand_x1_sg U11964 ( .A(n7423), .B(n5449), .X(n4619) );
  nand_x2_sg U11965 ( .A(n4957), .B(n4958), .X(n4936) );
  nand_x2_sg U11966 ( .A(n4938), .B(n4939), .X(n4937) );
  nand_x1_sg U11967 ( .A(n7424), .B(n5438), .X(n4957) );
  nand_x2_sg U11968 ( .A(n4999), .B(n5000), .X(n4978) );
  nand_x2_sg U11969 ( .A(n4980), .B(n4981), .X(n4979) );
  nand_x1_sg U11970 ( .A(n7423), .B(n5427), .X(n4999) );
  nand_x2_sg U11971 ( .A(n5225), .B(n5226), .X(n5204) );
  nand_x2_sg U11972 ( .A(n5206), .B(n5207), .X(n5205) );
  nand_x1_sg U11973 ( .A(n7424), .B(n5405), .X(n5225) );
  nand_x2_sg U11974 ( .A(n5149), .B(n5150), .X(n5128) );
  nand_x2_sg U11975 ( .A(n5130), .B(n5131), .X(n5129) );
  nand_x1_sg U11976 ( .A(n7423), .B(n5394), .X(n5149) );
  nand_x2_sg U11977 ( .A(n5113), .B(n5114), .X(n5092) );
  nand_x2_sg U11978 ( .A(n5094), .B(n5095), .X(n5093) );
  nand_x1_sg U11979 ( .A(n7424), .B(n5383), .X(n5113) );
  nand_x2_sg U11980 ( .A(n4873), .B(n4874), .X(n4852) );
  nand_x2_sg U11981 ( .A(n4854), .B(n4855), .X(n4853) );
  nand_x1_sg U11982 ( .A(n7423), .B(n5372), .X(n4873) );
  nand_x2_sg U11983 ( .A(n4831), .B(n4832), .X(n4810) );
  nand_x2_sg U11984 ( .A(n4812), .B(n4813), .X(n4811) );
  nand_x1_sg U11985 ( .A(n7424), .B(n5339), .X(n4831) );
  nand_x2_sg U11986 ( .A(n4535), .B(n4536), .X(n4514) );
  nand_x2_sg U11987 ( .A(n4516), .B(n4517), .X(n4515) );
  nand_x1_sg U11988 ( .A(n4452), .B(n5515), .X(n4535) );
  nand_x2_sg U11989 ( .A(n4661), .B(n4662), .X(n4640) );
  nand_x2_sg U11990 ( .A(n4642), .B(n4643), .X(n4641) );
  nand_x1_sg U11991 ( .A(n4452), .B(n5460), .X(n4661) );
  nand_x2_sg U11992 ( .A(n5185), .B(n5186), .X(n5164) );
  nand_x2_sg U11993 ( .A(n5166), .B(n5167), .X(n5165) );
  nand_x1_sg U11994 ( .A(n4452), .B(n5416), .X(n5185) );
  nand_x2_sg U11995 ( .A(n4915), .B(n4916), .X(n4894) );
  nand_x2_sg U11996 ( .A(n4896), .B(n4897), .X(n4895) );
  nand_x1_sg U11997 ( .A(n4452), .B(n5361), .X(n4915) );
  nand_x2_sg U11998 ( .A(n4789), .B(n4790), .X(n4768) );
  nand_x2_sg U11999 ( .A(n4770), .B(n4771), .X(n4769) );
  nand_x1_sg U12000 ( .A(n4452), .B(n5350), .X(n4789) );
  nand_x2_sg U12001 ( .A(n5041), .B(n5042), .X(n5020) );
  nand_x2_sg U12002 ( .A(n5022), .B(n5023), .X(n5021) );
  nand_x1_sg U12003 ( .A(n4452), .B(n5328), .X(n5041) );
  nand_x2_sg U12004 ( .A(n4417), .B(n4418), .X(n4411) );
  nand_x2_sg U12005 ( .A(n4413), .B(n4414), .X(n4412) );
  nand_x2_sg U12006 ( .A(n4468), .B(n4469), .X(n4464) );
  nand_x2_sg U12007 ( .A(n4466), .B(n4467), .X(n4465) );
  nand_x2_sg U12008 ( .A(n4680), .B(n4681), .X(n4676) );
  nand_x2_sg U12009 ( .A(n4678), .B(n4679), .X(n4677) );
  nand_x2_sg U12010 ( .A(n4594), .B(n4595), .X(n4590) );
  nand_x2_sg U12011 ( .A(n4592), .B(n4593), .X(n4591) );
  nand_x2_sg U12012 ( .A(n4848), .B(n4849), .X(n4844) );
  nand_x2_sg U12013 ( .A(n4846), .B(n4847), .X(n4845) );
  nand_x2_sg U12014 ( .A(n4806), .B(n4807), .X(n4802) );
  nand_x2_sg U12015 ( .A(n4804), .B(n4805), .X(n4803) );
  nand_x2_sg U12016 ( .A(n4510), .B(n4511), .X(n4506) );
  nand_x2_sg U12017 ( .A(n4508), .B(n4509), .X(n4507) );
  nand_x2_sg U12018 ( .A(n4636), .B(n4637), .X(n4632) );
  nand_x2_sg U12019 ( .A(n4634), .B(n4635), .X(n4633) );
  nand_x2_sg U12020 ( .A(n4890), .B(n4891), .X(n4886) );
  nand_x2_sg U12021 ( .A(n4888), .B(n4889), .X(n4887) );
  nand_x2_sg U12022 ( .A(n5237), .B(n5238), .X(n5232) );
  nand_x2_sg U12023 ( .A(n5234), .B(n5235), .X(n5233) );
  nand_x2_sg U12024 ( .A(n4974), .B(n4975), .X(n4970) );
  nand_x2_sg U12025 ( .A(n4972), .B(n4973), .X(n4971) );
  nand_x2_sg U12026 ( .A(n5200), .B(n5201), .X(n5196) );
  nand_x2_sg U12027 ( .A(n5198), .B(n5199), .X(n5197) );
  nand_x2_sg U12028 ( .A(n5088), .B(n5089), .X(n5084) );
  nand_x2_sg U12029 ( .A(n5086), .B(n5087), .X(n5085) );
  nand_x2_sg U12030 ( .A(n5016), .B(n5017), .X(n5012) );
  nand_x2_sg U12031 ( .A(n5014), .B(n5015), .X(n5013) );
  nor_x1_sg U12032 ( .A(n1023), .B(n7566), .X(n1022) );
  nor_x1_sg U12033 ( .A(n1125), .B(n7566), .X(n1124) );
  nand_x2_sg U12034 ( .A(n4552), .B(n4553), .X(n4548) );
  nand_x2_sg U12035 ( .A(n4550), .B(n4551), .X(n4549) );
  nand_x2_sg U12036 ( .A(n4722), .B(n4723), .X(n4718) );
  nand_x2_sg U12037 ( .A(n4720), .B(n4721), .X(n4719) );
  nand_x2_sg U12038 ( .A(n4932), .B(n4933), .X(n4928) );
  nand_x2_sg U12039 ( .A(n4930), .B(n4931), .X(n4929) );
  nand_x2_sg U12040 ( .A(n5124), .B(n5125), .X(n5120) );
  nand_x2_sg U12041 ( .A(n5122), .B(n5123), .X(n5121) );
  nand_x2_sg U12042 ( .A(n5160), .B(n5161), .X(n5156) );
  nand_x2_sg U12043 ( .A(n5158), .B(n5159), .X(n5157) );
  nand_x2_sg U12044 ( .A(n4764), .B(n4765), .X(n4760) );
  nand_x2_sg U12045 ( .A(n4762), .B(n4763), .X(n4761) );
  nor_x1_sg U12046 ( .A(n957), .B(n7566), .X(n956) );
  nor_x1_sg U12047 ( .A(n990), .B(n7566), .X(n989) );
  nor_x1_sg U12048 ( .A(n1158), .B(n7566), .X(n1157) );
  nor_x1_sg U12049 ( .A(n1191), .B(n7566), .X(n1190) );
  nor_x1_sg U12050 ( .A(n1295), .B(n7566), .X(n1294) );
  nor_x1_sg U12051 ( .A(n1328), .B(n7566), .X(n1327) );
  nor_x1_sg U12052 ( .A(n1361), .B(n7566), .X(n1360) );
  nor_x1_sg U12053 ( .A(n1463), .B(n7564), .X(n1462) );
  nor_x1_sg U12054 ( .A(n1496), .B(n7564), .X(n1495) );
  nand_x2_sg U12055 ( .A(n5252), .B(n5253), .X(n5251) );
  nand_x2_sg U12056 ( .A(n4565), .B(n4566), .X(n4564) );
  nand_x2_sg U12057 ( .A(n4434), .B(n4435), .X(n4433) );
  nand_x2_sg U12058 ( .A(n4481), .B(n4482), .X(n4480) );
  nand_x2_sg U12059 ( .A(n4693), .B(n4694), .X(n4692) );
  nand_x2_sg U12060 ( .A(n4735), .B(n4736), .X(n4734) );
  nand_x2_sg U12061 ( .A(n4607), .B(n4608), .X(n4606) );
  nand_x2_sg U12062 ( .A(n4987), .B(n4988), .X(n4986) );
  nand_x2_sg U12063 ( .A(n4861), .B(n4862), .X(n4860) );
  nand_x2_sg U12064 ( .A(n4819), .B(n4820), .X(n4818) );
  nand_x2_sg U12065 ( .A(n5101), .B(n5102), .X(n5100) );
  nand_x2_sg U12066 ( .A(n4945), .B(n4946), .X(n4944) );
  nand_x2_sg U12067 ( .A(n5213), .B(n5214), .X(n5212) );
  nand_x2_sg U12068 ( .A(n5137), .B(n5138), .X(n5136) );
  nand_x2_sg U12069 ( .A(n4523), .B(n4524), .X(n4522) );
  nand_x2_sg U12070 ( .A(n4649), .B(n4650), .X(n4648) );
  nand_x2_sg U12071 ( .A(n5173), .B(n5174), .X(n5172) );
  nand_x2_sg U12072 ( .A(n4903), .B(n4904), .X(n4902) );
  nand_x2_sg U12073 ( .A(n4777), .B(n4778), .X(n4776) );
  nand_x2_sg U12074 ( .A(n5029), .B(n5030), .X(n5028) );
  nor_x1_sg U12075 ( .A(n1532), .B(n7564), .X(n1531) );
  nand_x2_sg U12076 ( .A(n5269), .B(input_ready), .X(n5268) );
  nor_x1_sg U12077 ( .A(n5990), .B(n5950), .X(n5269) );
  nand_x1_sg U12078 ( .A(n4294), .B(n6381), .X(n4299) );
  nand_x2_sg U12079 ( .A(\update_output_0/n1535 ), .B(n7419), .X(n4307) );
  nand_x2_sg U12080 ( .A(n5263), .B(n7321), .X(n5262) );
  nand_x2_sg U12081 ( .A(n4704), .B(n7321), .X(n4703) );
  nand_x2_sg U12082 ( .A(n4746), .B(n7321), .X(n4745) );
  nand_x2_sg U12083 ( .A(n4660), .B(n7321), .X(n4659) );
  nand_x2_sg U12084 ( .A(n4998), .B(n7321), .X(n4997) );
  nand_x2_sg U12085 ( .A(n5184), .B(n7321), .X(n5183) );
  nand_x2_sg U12086 ( .A(n5112), .B(n7321), .X(n5111) );
  nand_x2_sg U12087 ( .A(n4914), .B(n7321), .X(n4913) );
  nand_x2_sg U12088 ( .A(n4830), .B(n7321), .X(n4829) );
  nand_x2_sg U12089 ( .A(n4576), .B(n7321), .X(n4575) );
  nand_x2_sg U12090 ( .A(n4534), .B(n7321), .X(n4533) );
  nand_x2_sg U12091 ( .A(n4448), .B(n7321), .X(n4447) );
  nand_x2_sg U12092 ( .A(n4492), .B(n7321), .X(n4491) );
  nand_x2_sg U12093 ( .A(n4618), .B(n7321), .X(n4617) );
  nand_x2_sg U12094 ( .A(n5224), .B(n7321), .X(n5223) );
  nand_x2_sg U12095 ( .A(n5148), .B(n7321), .X(n5147) );
  nand_x2_sg U12096 ( .A(n4872), .B(n7321), .X(n4871) );
  nand_x2_sg U12097 ( .A(n4788), .B(n7321), .X(n4787) );
  nand_x2_sg U12098 ( .A(n4956), .B(n7321), .X(n4955) );
  nand_x2_sg U12099 ( .A(n5040), .B(n5991), .X(n5039) );
  nand_x1_sg U12100 ( .A(n9244), .B(n4203), .X(n4198) );
  nand_x1_sg U12101 ( .A(n4200), .B(n5950), .X(n4199) );
  nor_x1_sg U12102 ( .A(n4201), .B(n9196), .X(n4200) );
  nand_x1_sg U12103 ( .A(n4202), .B(n5990), .X(n4205) );
  nand_x1_sg U12104 ( .A(n4203), .B(n4206), .X(n4204) );
  nand_x1_sg U12105 ( .A(n7310), .B(n5926), .X(n5282) );
  nor_x1_sg U12106 ( .A(n9202), .B(n5285), .X(n5281) );
  nand_x1_sg U12107 ( .A(n6254), .B(n7542), .X(n3614) );
  nand_x1_sg U12108 ( .A(n7132), .B(n7542), .X(n3612) );
  nand_x1_sg U12109 ( .A(n6216), .B(n7542), .X(n3610) );
  nand_x1_sg U12110 ( .A(n6100), .B(n7542), .X(n3608) );
  nand_x1_sg U12111 ( .A(n7284), .B(n7542), .X(n3604) );
  nand_x1_sg U12112 ( .A(n6356), .B(n7542), .X(n3602) );
  nand_x1_sg U12113 ( .A(n6130), .B(n7542), .X(n3600) );
  nand_x1_sg U12114 ( .A(n7130), .B(n7552), .X(n3598) );
  nand_x1_sg U12115 ( .A(n7258), .B(n7543), .X(n3596) );
  nand_x1_sg U12116 ( .A(n6330), .B(n7548), .X(n3594) );
  nand_x1_sg U12117 ( .A(n7128), .B(n7552), .X(n3592) );
  nand_x1_sg U12118 ( .A(n6214), .B(n7542), .X(n3590) );
  nand_x1_sg U12119 ( .A(n6098), .B(n7544), .X(n3588) );
  nand_x1_sg U12120 ( .A(n7256), .B(n7550), .X(n3586) );
  nand_x1_sg U12121 ( .A(n6328), .B(n7554), .X(n3584) );
  nand_x1_sg U12122 ( .A(n7126), .B(n7543), .X(n3582) );
  nand_x1_sg U12123 ( .A(n6212), .B(n7548), .X(n3580) );
  nand_x1_sg U12124 ( .A(n6096), .B(n7550), .X(n3578) );
  nand_x1_sg U12125 ( .A(n7254), .B(n7544), .X(n3576) );
  nand_x1_sg U12126 ( .A(n6326), .B(n7543), .X(n3574) );
  nand_x1_sg U12127 ( .A(n7124), .B(n7543), .X(n3572) );
  nand_x1_sg U12128 ( .A(n6210), .B(n7542), .X(n3570) );
  nand_x1_sg U12129 ( .A(n6094), .B(n7554), .X(n3568) );
  nand_x1_sg U12130 ( .A(n7282), .B(n7543), .X(n3564) );
  nand_x1_sg U12131 ( .A(n6354), .B(n7543), .X(n3562) );
  nand_x1_sg U12132 ( .A(n6128), .B(n7543), .X(n3560) );
  nand_x1_sg U12133 ( .A(n7122), .B(n7543), .X(n3558) );
  nand_x1_sg U12134 ( .A(n7178), .B(n7543), .X(n3556) );
  nand_x1_sg U12135 ( .A(n6252), .B(n7543), .X(n3554) );
  nand_x1_sg U12136 ( .A(n7120), .B(n7543), .X(n3552) );
  nand_x1_sg U12137 ( .A(n6208), .B(n7550), .X(n3550) );
  nand_x1_sg U12138 ( .A(n6092), .B(n7554), .X(n3548) );
  nand_x1_sg U12139 ( .A(n7176), .B(n7550), .X(n3546) );
  nand_x1_sg U12140 ( .A(n6250), .B(n7554), .X(n3544) );
  nand_x1_sg U12141 ( .A(n7118), .B(n7550), .X(n3542) );
  nand_x1_sg U12142 ( .A(n6206), .B(n7554), .X(n3540) );
  nand_x1_sg U12143 ( .A(n6090), .B(n7544), .X(n3538) );
  nand_x1_sg U12144 ( .A(n7174), .B(n7542), .X(n3536) );
  nand_x1_sg U12145 ( .A(n6248), .B(n7544), .X(n3534) );
  nand_x1_sg U12146 ( .A(n7116), .B(n7544), .X(n3532) );
  nand_x1_sg U12147 ( .A(n6204), .B(n7544), .X(n3530) );
  nand_x1_sg U12148 ( .A(n6088), .B(n7544), .X(n3528) );
  nand_x1_sg U12149 ( .A(n7280), .B(n7544), .X(n3524) );
  nand_x1_sg U12150 ( .A(n6352), .B(n7544), .X(n3522) );
  nand_x1_sg U12151 ( .A(n6126), .B(n7544), .X(n3520) );
  nand_x1_sg U12152 ( .A(n7114), .B(n7550), .X(n3518) );
  nand_x1_sg U12153 ( .A(n7278), .B(n7554), .X(n3516) );
  nand_x1_sg U12154 ( .A(n6350), .B(n7551), .X(n3514) );
  nand_x1_sg U12155 ( .A(n6124), .B(n7547), .X(n3512) );
  nand_x1_sg U12156 ( .A(n7198), .B(n7544), .X(n3510) );
  nand_x1_sg U12157 ( .A(n6272), .B(n7542), .X(n3508) );
  nand_x1_sg U12158 ( .A(n7276), .B(n7550), .X(n3506) );
  nand_x1_sg U12159 ( .A(n6348), .B(n7554), .X(n3504) );
  nand_x1_sg U12160 ( .A(n6122), .B(n7544), .X(n3502) );
  nand_x1_sg U12161 ( .A(n7196), .B(n7542), .X(n3500) );
  nand_x1_sg U12162 ( .A(n6270), .B(n7554), .X(n3498) );
  nand_x1_sg U12163 ( .A(n7274), .B(n7551), .X(n3496) );
  nand_x1_sg U12164 ( .A(n6346), .B(n7544), .X(n3494) );
  nand_x1_sg U12165 ( .A(n6120), .B(n7550), .X(n3492) );
  nand_x1_sg U12166 ( .A(n7194), .B(n7550), .X(n3490) );
  nand_x1_sg U12167 ( .A(n6268), .B(n7542), .X(n3488) );
  nand_x1_sg U12168 ( .A(n7252), .B(n7554), .X(n3484) );
  nand_x1_sg U12169 ( .A(n6324), .B(n7550), .X(n3482) );
  nand_x1_sg U12170 ( .A(n7112), .B(n7544), .X(n3480) );
  nand_x1_sg U12171 ( .A(n6202), .B(n7543), .X(n3478) );
  nand_x1_sg U12172 ( .A(n7250), .B(n7542), .X(n3476) );
  nand_x1_sg U12173 ( .A(n6322), .B(n7550), .X(n3474) );
  nand_x1_sg U12174 ( .A(n7110), .B(n7542), .X(n3472) );
  nand_x1_sg U12175 ( .A(n6086), .B(n7548), .X(n3470) );
  nand_x1_sg U12176 ( .A(n6040), .B(n7544), .X(n3468) );
  nand_x1_sg U12177 ( .A(n7248), .B(n7545), .X(n3466) );
  nand_x1_sg U12178 ( .A(n6320), .B(n7550), .X(n3464) );
  nand_x1_sg U12179 ( .A(n7108), .B(n7546), .X(n3462) );
  nand_x1_sg U12180 ( .A(n6084), .B(n7552), .X(n3460) );
  nand_x1_sg U12181 ( .A(n6038), .B(n7549), .X(n3458) );
  nand_x1_sg U12182 ( .A(n7246), .B(n7549), .X(n3456) );
  nand_x1_sg U12183 ( .A(n6318), .B(n7550), .X(n3454) );
  nand_x1_sg U12184 ( .A(n7106), .B(n7552), .X(n3452) );
  nand_x1_sg U12185 ( .A(n6082), .B(n7548), .X(n3450) );
  nand_x1_sg U12186 ( .A(n6036), .B(n7554), .X(n3448) );
  nand_x1_sg U12187 ( .A(n7244), .B(n7542), .X(n3444) );
  nand_x1_sg U12188 ( .A(n6316), .B(n7552), .X(n3442) );
  nand_x1_sg U12189 ( .A(n7104), .B(n7549), .X(n3440) );
  nand_x1_sg U12190 ( .A(n7102), .B(n7545), .X(n3438) );
  nand_x1_sg U12191 ( .A(n7242), .B(n7542), .X(n3436) );
  nand_x1_sg U12192 ( .A(n6314), .B(n7545), .X(n3434) );
  nand_x1_sg U12193 ( .A(n7100), .B(n7547), .X(n3432) );
  nand_x1_sg U12194 ( .A(n6200), .B(n7545), .X(n3430) );
  nand_x1_sg U12195 ( .A(n6034), .B(n7551), .X(n3428) );
  nand_x1_sg U12196 ( .A(n7240), .B(n7544), .X(n3426) );
  nand_x1_sg U12197 ( .A(n6312), .B(n7548), .X(n3424) );
  nand_x1_sg U12198 ( .A(n7098), .B(n7554), .X(n3422) );
  nand_x1_sg U12199 ( .A(n6198), .B(n7551), .X(n3420) );
  nand_x1_sg U12200 ( .A(n6032), .B(n7544), .X(n3418) );
  nand_x1_sg U12201 ( .A(n7238), .B(n7554), .X(n3416) );
  nand_x1_sg U12202 ( .A(n6310), .B(n7551), .X(n3414) );
  nand_x1_sg U12203 ( .A(n7096), .B(n7549), .X(n3412) );
  nand_x1_sg U12204 ( .A(n6196), .B(n7550), .X(n3410) );
  nand_x1_sg U12205 ( .A(n6030), .B(n7544), .X(n3408) );
  nand_x1_sg U12206 ( .A(n7094), .B(n7554), .X(n3404) );
  nand_x1_sg U12207 ( .A(n6194), .B(n7542), .X(n3402) );
  nand_x1_sg U12208 ( .A(n7092), .B(n7554), .X(n3398) );
  nand_x1_sg U12209 ( .A(n7172), .B(n7543), .X(n3396) );
  nand_x1_sg U12210 ( .A(n6246), .B(n7554), .X(n3394) );
  nand_x1_sg U12211 ( .A(n7090), .B(n7542), .X(n3392) );
  nand_x1_sg U12212 ( .A(n6192), .B(n7554), .X(n3390) );
  nand_x1_sg U12213 ( .A(n6080), .B(n7544), .X(n3388) );
  nand_x1_sg U12214 ( .A(n7170), .B(n7545), .X(n3386) );
  nand_x1_sg U12215 ( .A(n6244), .B(n7552), .X(n3384) );
  nand_x1_sg U12216 ( .A(n7088), .B(n7542), .X(n3382) );
  nand_x1_sg U12217 ( .A(n6190), .B(n7544), .X(n3380) );
  nand_x1_sg U12218 ( .A(n6078), .B(n7551), .X(n3378) );
  nand_x1_sg U12219 ( .A(n7168), .B(n7542), .X(n3376) );
  nand_x1_sg U12220 ( .A(n6242), .B(n7543), .X(n3374) );
  nand_x1_sg U12221 ( .A(n7086), .B(n7543), .X(n3372) );
  nand_x1_sg U12222 ( .A(n6188), .B(n7543), .X(n3370) );
  nand_x1_sg U12223 ( .A(n6076), .B(n7543), .X(n3368) );
  nand_x1_sg U12224 ( .A(n7084), .B(n7543), .X(n3364) );
  nand_x1_sg U12225 ( .A(n6186), .B(n7543), .X(n3362) );
  nand_x1_sg U12226 ( .A(n7082), .B(n7547), .X(n3358) );
  nand_x1_sg U12227 ( .A(n7166), .B(n7546), .X(n3356) );
  nand_x1_sg U12228 ( .A(n6240), .B(n7545), .X(n3354) );
  nand_x1_sg U12229 ( .A(n7080), .B(n7546), .X(n3352) );
  nand_x1_sg U12230 ( .A(n6184), .B(n7549), .X(n3350) );
  nand_x1_sg U12231 ( .A(n6074), .B(n7546), .X(n3348) );
  nand_x1_sg U12232 ( .A(n7164), .B(n7547), .X(n3346) );
  nand_x1_sg U12233 ( .A(n6238), .B(n7546), .X(n3344) );
  nand_x1_sg U12234 ( .A(n7078), .B(n7546), .X(n3342) );
  nand_x1_sg U12235 ( .A(n6182), .B(n7546), .X(n3340) );
  nand_x1_sg U12236 ( .A(n6072), .B(n7546), .X(n3338) );
  nand_x1_sg U12237 ( .A(n7162), .B(n7546), .X(n3336) );
  nand_x1_sg U12238 ( .A(n6236), .B(n7546), .X(n3334) );
  nand_x1_sg U12239 ( .A(n7076), .B(n7546), .X(n3332) );
  nand_x1_sg U12240 ( .A(n6180), .B(n7546), .X(n3330) );
  nand_x1_sg U12241 ( .A(n6070), .B(n7546), .X(n3328) );
  nand_x1_sg U12242 ( .A(n7074), .B(n7552), .X(n3324) );
  nand_x1_sg U12243 ( .A(n6178), .B(n7551), .X(n3322) );
  nand_x1_sg U12244 ( .A(n7072), .B(n7547), .X(n3318) );
  nand_x1_sg U12245 ( .A(n7236), .B(n7545), .X(n3316) );
  nand_x1_sg U12246 ( .A(n6308), .B(n7549), .X(n3314) );
  nand_x1_sg U12247 ( .A(n6176), .B(n7549), .X(n3312) );
  nand_x1_sg U12248 ( .A(n6068), .B(n7547), .X(n3310) );
  nand_x1_sg U12249 ( .A(n6028), .B(n7545), .X(n3308) );
  nand_x1_sg U12250 ( .A(n7234), .B(n7545), .X(n3306) );
  nand_x1_sg U12251 ( .A(n6306), .B(n7549), .X(n3304) );
  nand_x1_sg U12252 ( .A(n6174), .B(n7542), .X(n3302) );
  nand_x1_sg U12253 ( .A(n6066), .B(n7544), .X(n3300) );
  nand_x1_sg U12254 ( .A(n6026), .B(n7552), .X(n3298) );
  nand_x1_sg U12255 ( .A(n7232), .B(n7543), .X(n3296) );
  nand_x1_sg U12256 ( .A(n6304), .B(n7545), .X(n3294) );
  nand_x1_sg U12257 ( .A(n6172), .B(n7545), .X(n3292) );
  nand_x1_sg U12258 ( .A(n6064), .B(n7545), .X(n3290) );
  nand_x1_sg U12259 ( .A(n6024), .B(n7545), .X(n3288) );
  nand_x1_sg U12260 ( .A(n7070), .B(n7545), .X(n3284) );
  nand_x1_sg U12261 ( .A(n6170), .B(n7545), .X(n3282) );
  nand_x1_sg U12262 ( .A(n7068), .B(n7546), .X(n3278) );
  nand_x1_sg U12263 ( .A(n7230), .B(n7546), .X(n3276) );
  nand_x1_sg U12264 ( .A(n6302), .B(n7546), .X(n3274) );
  nand_x1_sg U12265 ( .A(n7066), .B(n7546), .X(n3272) );
  nand_x1_sg U12266 ( .A(n6168), .B(n7546), .X(n3270) );
  nand_x1_sg U12267 ( .A(n6062), .B(n7546), .X(n3268) );
  nand_x1_sg U12268 ( .A(n7228), .B(n7546), .X(n3266) );
  nand_x1_sg U12269 ( .A(n6300), .B(n7546), .X(n3264) );
  nand_x1_sg U12270 ( .A(n7064), .B(n7547), .X(n3262) );
  nand_x1_sg U12271 ( .A(n6166), .B(n7547), .X(n3260) );
  nand_x1_sg U12272 ( .A(n6060), .B(n7547), .X(n3258) );
  nand_x1_sg U12273 ( .A(n7226), .B(n7547), .X(n3256) );
  nand_x1_sg U12274 ( .A(n6298), .B(n7547), .X(n3254) );
  nand_x1_sg U12275 ( .A(n7062), .B(n7547), .X(n3252) );
  nand_x1_sg U12276 ( .A(n6164), .B(n7547), .X(n3250) );
  nand_x1_sg U12277 ( .A(n6058), .B(n7547), .X(n3248) );
  nand_x1_sg U12278 ( .A(n7192), .B(n7545), .X(n3246) );
  nand_x1_sg U12279 ( .A(n6266), .B(n7547), .X(n3244) );
  nand_x1_sg U12280 ( .A(n7270), .B(n7545), .X(n3240) );
  nand_x1_sg U12281 ( .A(n6118), .B(n7549), .X(n3238) );
  nand_x1_sg U12282 ( .A(n7224), .B(n7551), .X(n3236) );
  nand_x1_sg U12283 ( .A(n6296), .B(n7546), .X(n3234) );
  nand_x1_sg U12284 ( .A(n7060), .B(n7543), .X(n3232) );
  nand_x1_sg U12285 ( .A(n6056), .B(n7552), .X(n3230) );
  nand_x1_sg U12286 ( .A(n6022), .B(n7552), .X(n3228) );
  nand_x1_sg U12287 ( .A(n7222), .B(n7552), .X(n3226) );
  nand_x1_sg U12288 ( .A(n6294), .B(n7552), .X(n3224) );
  nand_x1_sg U12289 ( .A(n7058), .B(n7552), .X(n3222) );
  nand_x1_sg U12290 ( .A(n6054), .B(n7552), .X(n3220) );
  nand_x1_sg U12291 ( .A(n6020), .B(n7549), .X(n3218) );
  nand_x1_sg U12292 ( .A(n7220), .B(n7552), .X(n3216) );
  nand_x1_sg U12293 ( .A(n6292), .B(n7543), .X(n3214) );
  nand_x1_sg U12294 ( .A(n7056), .B(n7548), .X(n3212) );
  nand_x1_sg U12295 ( .A(n6052), .B(n7551), .X(n3210) );
  nand_x1_sg U12296 ( .A(n6018), .B(n7554), .X(n3208) );
  nand_x1_sg U12297 ( .A(n7272), .B(n7554), .X(n3206) );
  nand_x1_sg U12298 ( .A(n6344), .B(n7554), .X(n3204) );
  nand_x1_sg U12299 ( .A(n7268), .B(n7554), .X(n3200) );
  nand_x1_sg U12300 ( .A(n6342), .B(n7547), .X(n3198) );
  nand_x1_sg U12301 ( .A(n7218), .B(n7545), .X(n3196) );
  nand_x1_sg U12302 ( .A(n6290), .B(n7546), .X(n3194) );
  nand_x1_sg U12303 ( .A(n7054), .B(n7543), .X(n3192) );
  nand_x1_sg U12304 ( .A(n6162), .B(n7549), .X(n3190) );
  nand_x1_sg U12305 ( .A(n6016), .B(n7547), .X(n3188) );
  nand_x1_sg U12306 ( .A(n7216), .B(n7548), .X(n3186) );
  nand_x1_sg U12307 ( .A(n6288), .B(n7542), .X(n3184) );
  nand_x1_sg U12308 ( .A(n7052), .B(n7548), .X(n3182) );
  nand_x1_sg U12309 ( .A(n6160), .B(n7547), .X(n3180) );
  nand_x1_sg U12310 ( .A(n6014), .B(n7546), .X(n3178) );
  nand_x1_sg U12311 ( .A(n7214), .B(n7544), .X(n3176) );
  nand_x1_sg U12312 ( .A(n6286), .B(n7542), .X(n3174) );
  nand_x1_sg U12313 ( .A(n7050), .B(n7550), .X(n3172) );
  nand_x1_sg U12314 ( .A(n6158), .B(n7547), .X(n3170) );
  nand_x1_sg U12315 ( .A(n6012), .B(n7549), .X(n3168) );
  nand_x1_sg U12316 ( .A(n7048), .B(n7551), .X(n3110) );
  nand_x1_sg U12317 ( .A(n6340), .B(n7547), .X(n3108) );
  nand_x1_sg U12318 ( .A(n7160), .B(n7545), .X(n3106) );
  nand_x1_sg U12319 ( .A(n6234), .B(n7544), .X(n3103) );
  nand_x1_sg U12320 ( .A(n7542), .B(n5948), .X(n3606) );
  nand_x1_sg U12321 ( .A(n7543), .B(n6006), .X(n3566) );
  nand_x1_sg U12322 ( .A(n7544), .B(n5998), .X(n3526) );
  nand_x1_sg U12323 ( .A(n7550), .B(n6044), .X(n3486) );
  nand_x1_sg U12324 ( .A(n7542), .B(n5986), .X(n3446) );
  nand_x1_sg U12325 ( .A(n7544), .B(n6042), .X(n3406) );
  nand_x1_sg U12326 ( .A(n7543), .B(n7033), .X(n3366) );
  nand_x1_sg U12327 ( .A(n7551), .B(n6004), .X(n3326) );
  nand_x1_sg U12328 ( .A(n7545), .B(n5996), .X(n3286) );
  nand_x1_sg U12329 ( .A(n7548), .B(n7031), .X(n3166) );
  nand_x1_sg U12330 ( .A(n7548), .B(n5984), .X(n3164) );
  nand_x1_sg U12331 ( .A(n7548), .B(n5982), .X(n3162) );
  nand_x1_sg U12332 ( .A(n7548), .B(n5980), .X(n3160) );
  nand_x1_sg U12333 ( .A(n7548), .B(n5946), .X(n3158) );
  nand_x1_sg U12334 ( .A(n7548), .B(n5978), .X(n3156) );
  nand_x1_sg U12335 ( .A(n7548), .B(n5944), .X(n3154) );
  nand_x1_sg U12336 ( .A(n7548), .B(n5942), .X(n3152) );
  nand_x1_sg U12337 ( .A(n7544), .B(n7029), .X(n3150) );
  nand_x1_sg U12338 ( .A(n7552), .B(n5976), .X(n3148) );
  nand_x1_sg U12339 ( .A(n7550), .B(n5974), .X(n3146) );
  nand_x1_sg U12340 ( .A(n7546), .B(n5972), .X(n3144) );
  nand_x1_sg U12341 ( .A(n7547), .B(n5940), .X(n3142) );
  nand_x1_sg U12342 ( .A(n7549), .B(n5970), .X(n3140) );
  nand_x1_sg U12343 ( .A(n7548), .B(n5938), .X(n3138) );
  nand_x1_sg U12344 ( .A(n7549), .B(n5936), .X(n3136) );
  nand_x1_sg U12345 ( .A(n7549), .B(n7027), .X(n3134) );
  nand_x1_sg U12346 ( .A(n7549), .B(n5968), .X(n3132) );
  nand_x1_sg U12347 ( .A(n7549), .B(n5966), .X(n3130) );
  nand_x1_sg U12348 ( .A(n7549), .B(n5964), .X(n3128) );
  nand_x1_sg U12349 ( .A(n7549), .B(n5934), .X(n3126) );
  nand_x1_sg U12350 ( .A(n7549), .B(n5962), .X(n3124) );
  nand_x1_sg U12351 ( .A(n7549), .B(n5932), .X(n3122) );
  nand_x1_sg U12352 ( .A(n7549), .B(n5960), .X(n3120) );
  nand_x1_sg U12353 ( .A(n7549), .B(n7025), .X(n3118) );
  nand_x1_sg U12354 ( .A(n7551), .B(n5958), .X(n3116) );
  nand_x1_sg U12355 ( .A(n7547), .B(n5956), .X(n3114) );
  nand_x1_sg U12356 ( .A(n7550), .B(n5954), .X(n3112) );
  nand_x1_sg U12357 ( .A(n7044), .B(n7547), .X(n3320) );
  nand_x1_sg U12358 ( .A(n7043), .B(n7545), .X(n3280) );
  nand_x1_sg U12359 ( .A(n7042), .B(n7551), .X(n3242) );
  nand_x1_sg U12360 ( .A(n6049), .B(n7554), .X(n3202) );
  nand_x1_sg U12361 ( .A(n7046), .B(n7544), .X(n3400) );
  nand_x1_sg U12362 ( .A(n7045), .B(n7543), .X(n3360) );
  nand_x1_sg U12363 ( .A(n5992), .B(n3092), .X(n3091) );
  nor_x1_sg U12364 ( .A(n3093), .B(n3094), .X(n3090) );
  nand_x1_sg U12365 ( .A(n6146), .B(n7554), .X(n3742) );
  nand_x1_sg U12366 ( .A(n7210), .B(n7552), .X(n3740) );
  nand_x1_sg U12367 ( .A(n6282), .B(n7554), .X(n3738) );
  nand_x1_sg U12368 ( .A(n7298), .B(n7554), .X(n3736) );
  nand_x1_sg U12369 ( .A(n6370), .B(n7543), .X(n3734) );
  nand_x1_sg U12370 ( .A(n6144), .B(n7549), .X(n3732) );
  nand_x1_sg U12371 ( .A(n7208), .B(n7546), .X(n3730) );
  nand_x1_sg U12372 ( .A(n6280), .B(n7549), .X(n3728) );
  nand_x1_sg U12373 ( .A(n7296), .B(n7548), .X(n3724) );
  nand_x1_sg U12374 ( .A(n6368), .B(n7552), .X(n3722) );
  nand_x1_sg U12375 ( .A(n6142), .B(n7548), .X(n3720) );
  nand_x1_sg U12376 ( .A(n7206), .B(n7550), .X(n3718) );
  nand_x1_sg U12377 ( .A(n7294), .B(n7556), .X(n3716) );
  nand_x1_sg U12378 ( .A(n6366), .B(n7551), .X(n3714) );
  nand_x1_sg U12379 ( .A(n6140), .B(n7551), .X(n3712) );
  nand_x1_sg U12380 ( .A(n7204), .B(n7548), .X(n3710) );
  nand_x1_sg U12381 ( .A(n6278), .B(n7551), .X(n3708) );
  nand_x1_sg U12382 ( .A(n7292), .B(n7554), .X(n3706) );
  nand_x1_sg U12383 ( .A(n6364), .B(n7554), .X(n3704) );
  nand_x1_sg U12384 ( .A(n6138), .B(n7554), .X(n3702) );
  nand_x1_sg U12385 ( .A(n7202), .B(n7547), .X(n3700) );
  nand_x1_sg U12386 ( .A(n6276), .B(n7547), .X(n3698) );
  nand_x1_sg U12387 ( .A(n7290), .B(n7554), .X(n3696) );
  nand_x1_sg U12388 ( .A(n6362), .B(n7554), .X(n3694) );
  nand_x1_sg U12389 ( .A(n6136), .B(n7548), .X(n3692) );
  nand_x1_sg U12390 ( .A(n7200), .B(n7552), .X(n3690) );
  nand_x1_sg U12391 ( .A(n6274), .B(n7554), .X(n3688) );
  nand_x1_sg U12392 ( .A(n7288), .B(n7554), .X(n3684) );
  nand_x1_sg U12393 ( .A(n6360), .B(n7552), .X(n3682) );
  nand_x1_sg U12394 ( .A(n6134), .B(n7551), .X(n3680) );
  nand_x1_sg U12395 ( .A(n7146), .B(n7551), .X(n3678) );
  nand_x1_sg U12396 ( .A(n7264), .B(n7554), .X(n3676) );
  nand_x1_sg U12397 ( .A(n6336), .B(n7556), .X(n3674) );
  nand_x1_sg U12398 ( .A(n7144), .B(n7554), .X(n3672) );
  nand_x1_sg U12399 ( .A(n6226), .B(n7554), .X(n3670) );
  nand_x1_sg U12400 ( .A(n6110), .B(n7551), .X(n3668) );
  nand_x1_sg U12401 ( .A(n7262), .B(n7545), .X(n3666) );
  nand_x1_sg U12402 ( .A(n6334), .B(n7554), .X(n3664) );
  nand_x1_sg U12403 ( .A(n7142), .B(n7549), .X(n3662) );
  nand_x1_sg U12404 ( .A(n6224), .B(n7554), .X(n3660) );
  nand_x1_sg U12405 ( .A(n6108), .B(n7550), .X(n3658) );
  nand_x1_sg U12406 ( .A(n7260), .B(n7548), .X(n3656) );
  nand_x1_sg U12407 ( .A(n6332), .B(n7554), .X(n3654) );
  nand_x1_sg U12408 ( .A(n7140), .B(n7550), .X(n3652) );
  nand_x1_sg U12409 ( .A(n6222), .B(n7551), .X(n3650) );
  nand_x1_sg U12410 ( .A(n6106), .B(n7554), .X(n3648) );
  nand_x1_sg U12411 ( .A(n7286), .B(n7552), .X(n3644) );
  nand_x1_sg U12412 ( .A(n6358), .B(n7550), .X(n3642) );
  nand_x1_sg U12413 ( .A(n6132), .B(n7551), .X(n3640) );
  nand_x1_sg U12414 ( .A(n7138), .B(n7547), .X(n3638) );
  nand_x1_sg U12415 ( .A(n7184), .B(n7554), .X(n3636) );
  nand_x1_sg U12416 ( .A(n6258), .B(n7552), .X(n3634) );
  nand_x1_sg U12417 ( .A(n7136), .B(n7554), .X(n3632) );
  nand_x1_sg U12418 ( .A(n6220), .B(n7554), .X(n3630) );
  nand_x1_sg U12419 ( .A(n6104), .B(n7550), .X(n3628) );
  nand_x1_sg U12420 ( .A(n7182), .B(n7554), .X(n3626) );
  nand_x1_sg U12421 ( .A(n6256), .B(n7551), .X(n3624) );
  nand_x1_sg U12422 ( .A(n7134), .B(n7548), .X(n3622) );
  nand_x1_sg U12423 ( .A(n6218), .B(n7545), .X(n3620) );
  nand_x1_sg U12424 ( .A(n6102), .B(n7551), .X(n3618) );
  nand_x1_sg U12425 ( .A(n7180), .B(n7554), .X(n3616) );
  nand_x1_sg U12426 ( .A(n7552), .B(n6046), .X(n3726) );
  nand_x1_sg U12427 ( .A(n7554), .B(n7035), .X(n3686) );
  nand_x1_sg U12428 ( .A(n7554), .B(n6008), .X(n3646) );
  nand_x1_sg U12429 ( .A(n7304), .B(n7552), .X(n3804) );
  nand_x1_sg U12430 ( .A(n6376), .B(n7549), .X(n3802) );
  nand_x1_sg U12431 ( .A(n6150), .B(n7548), .X(n3800) );
  nand_x1_sg U12432 ( .A(n7158), .B(n7547), .X(n3798) );
  nand_x1_sg U12433 ( .A(n7190), .B(n7554), .X(n3796) );
  nand_x1_sg U12434 ( .A(n6264), .B(n7554), .X(n3794) );
  nand_x1_sg U12435 ( .A(n7156), .B(n7550), .X(n3792) );
  nand_x1_sg U12436 ( .A(n6232), .B(n7550), .X(n3790) );
  nand_x1_sg U12437 ( .A(n6116), .B(n7552), .X(n3788) );
  nand_x1_sg U12438 ( .A(n7188), .B(n7554), .X(n3786) );
  nand_x1_sg U12439 ( .A(n6262), .B(n7550), .X(n3784) );
  nand_x1_sg U12440 ( .A(n7154), .B(n7552), .X(n3782) );
  nand_x1_sg U12441 ( .A(n6230), .B(n7545), .X(n3780) );
  nand_x1_sg U12442 ( .A(n6114), .B(n7548), .X(n3778) );
  nand_x1_sg U12443 ( .A(n7186), .B(n7545), .X(n3776) );
  nand_x1_sg U12444 ( .A(n6260), .B(n7554), .X(n3774) );
  nand_x1_sg U12445 ( .A(n7152), .B(n7551), .X(n3772) );
  nand_x1_sg U12446 ( .A(n6228), .B(n7554), .X(n3770) );
  nand_x1_sg U12447 ( .A(n6112), .B(n7545), .X(n3768) );
  nand_x1_sg U12448 ( .A(n7266), .B(n7546), .X(n3764) );
  nand_x1_sg U12449 ( .A(n6338), .B(n7554), .X(n3762) );
  nand_x1_sg U12450 ( .A(n7150), .B(n7550), .X(n3760) );
  nand_x1_sg U12451 ( .A(n7148), .B(n7542), .X(n3758) );
  nand_x1_sg U12452 ( .A(n7302), .B(n7548), .X(n3756) );
  nand_x1_sg U12453 ( .A(n6374), .B(n7552), .X(n3754) );
  nand_x1_sg U12454 ( .A(n6148), .B(n7554), .X(n3752) );
  nand_x1_sg U12455 ( .A(n7212), .B(n7551), .X(n3750) );
  nand_x1_sg U12456 ( .A(n6284), .B(n7549), .X(n3748) );
  nand_x1_sg U12457 ( .A(n7300), .B(n7551), .X(n3746) );
  nand_x1_sg U12458 ( .A(n6372), .B(n7545), .X(n3744) );
  nand_x1_sg U12459 ( .A(n7548), .B(n6010), .X(n3806) );
  nand_x1_sg U12460 ( .A(n7551), .B(n6000), .X(n3766) );
  nand_x1_sg U12461 ( .A(n7312), .B(n3092), .X(n4304) );
  nor_x1_sg U12462 ( .A(n4306), .B(n3092), .X(n4305) );
  nand_x2_sg U12463 ( .A(n7520), .B(n5307), .X(n5310) );
  nand_x2_sg U12464 ( .A(n9214), .B(n7318), .X(n5311) );
  nand_x1_sg U12465 ( .A(n9198), .B(n5988), .X(n5308) );
  nand_x1_sg U12466 ( .A(n5925), .B(n7525), .X(n5309) );
  nand_x1_sg U12467 ( .A(n6152), .B(n4187), .X(n4180) );
  nand_x1_sg U12468 ( .A(n5302), .B(n9203), .X(n5301) );
  nand_x1_sg U12469 ( .A(n6383), .B(n5299), .X(n5300) );
  nand_x1_sg U12470 ( .A(n5305), .B(n9203), .X(n5304) );
  nand_x1_sg U12471 ( .A(n7318), .B(n5277), .X(n5303) );
  nor_x1_sg U12472 ( .A(n7318), .B(n3101), .X(n5305) );
  nand_x1_sg U12473 ( .A(n5927), .B(n3817), .X(n3815) );
  nand_x1_sg U12474 ( .A(n9203), .B(n3818), .X(n3817) );
  nand_x1_sg U12475 ( .A(n7310), .B(n6379), .X(n3818) );
  nand_x1_sg U12476 ( .A(n3812), .B(n3813), .X(n3811) );
  nand_x1_sg U12477 ( .A(n7314), .B(n3815), .X(n3810) );
  nor_x1_sg U12478 ( .A(n7314), .B(n3814), .X(n3812) );
  nand_x1_sg U12479 ( .A(n5280), .B(n3813), .X(n5279) );
  nand_x1_sg U12480 ( .A(n6377), .B(n5926), .X(n5278) );
  nor_x1_sg U12481 ( .A(n6377), .B(n9213), .X(n5280) );
  nand_x1_sg U12482 ( .A(n7308), .B(n5283), .X(n5288) );
  nand_x1_sg U12483 ( .A(n3813), .B(n9213), .X(n5289) );
  nor_x1_sg U12484 ( .A(n5952), .B(n9209), .X(n2070) );
  nor_x1_sg U12485 ( .A(n5326), .B(state[1]), .X(n5325) );
  nor_x1_sg U12486 ( .A(reset), .B(n5322), .X(n19) );
  nand_x2_sg U12487 ( .A(n5320), .B(n9211), .X(n5318) );
  nor_x1_sg U12488 ( .A(n5990), .B(n5952), .X(n5320) );
  nor_x1_sg U12489 ( .A(reset), .B(n5314), .X(n20) );
  nor_x1_sg U12490 ( .A(n9208), .B(n5887), .X(n5315) );
  nor_x1_sg U12491 ( .A(n5317), .B(n9210), .X(n5316) );
  nand_x1_sg U12492 ( .A(n7318), .B(n1998), .X(n1997) );
  nor_x1_sg U12493 ( .A(n2001), .B(n2002), .X(n2000) );
  nor_x1_sg U12494 ( .A(n2007), .B(n2008), .X(n1999) );
  nand_x1_sg U12495 ( .A(n7314), .B(n1854), .X(n1794) );
  nor_x1_sg U12496 ( .A(n1857), .B(n1858), .X(n1856) );
  nor_x1_sg U12497 ( .A(n1877), .B(n1878), .X(n1855) );
  nor_x1_sg U12498 ( .A(n7316), .B(n6234), .X(n2068) );
  nand_x2_sg U12499 ( .A(n1819), .B(n9076), .X(n1818) );
  nor_x1_sg U12500 ( .A(n7270), .B(n6118), .X(n1819) );
  nand_x1_sg U12501 ( .A(n9073), .B(n1665), .X(n1659) );
  nor_x1_sg U12502 ( .A(n6082), .B(n6036), .X(n1666) );
  nor_x1_sg U12503 ( .A(n7106), .B(n9027), .X(n1667) );
  nand_x1_sg U12504 ( .A(n9073), .B(n1729), .X(n1723) );
  nor_x1_sg U12505 ( .A(n6086), .B(n6040), .X(n1730) );
  nor_x1_sg U12506 ( .A(n7110), .B(n9025), .X(n1731) );
  nand_x1_sg U12507 ( .A(n6044), .B(n9073), .X(n1803) );
  nand_x1_sg U12508 ( .A(n9073), .B(n1978), .X(n1972) );
  nor_x1_sg U12509 ( .A(n6084), .B(n6038), .X(n1979) );
  nor_x1_sg U12510 ( .A(n7108), .B(n9026), .X(n1980) );
  nand_x1_sg U12511 ( .A(n9074), .B(n1661), .X(n1660) );
  nor_x1_sg U12512 ( .A(n6196), .B(n6030), .X(n1662) );
  nor_x1_sg U12513 ( .A(n7096), .B(n9031), .X(n1663) );
  nand_x1_sg U12514 ( .A(n9074), .B(n1725), .X(n1724) );
  nor_x1_sg U12515 ( .A(n6200), .B(n6034), .X(n1726) );
  nor_x1_sg U12516 ( .A(n7100), .B(n9029), .X(n1727) );
  nand_x1_sg U12517 ( .A(n5986), .B(n9074), .X(n1804) );
  nand_x1_sg U12518 ( .A(n9074), .B(n1974), .X(n1973) );
  nor_x1_sg U12519 ( .A(n6198), .B(n6032), .X(n1975) );
  nor_x1_sg U12520 ( .A(n7098), .B(n9030), .X(n1976) );
  nand_x1_sg U12521 ( .A(n9076), .B(n1653), .X(n1647) );
  nor_x1_sg U12522 ( .A(n6052), .B(n6018), .X(n1654) );
  nor_x1_sg U12523 ( .A(n7056), .B(n9051), .X(n1655) );
  nand_x1_sg U12524 ( .A(n9076), .B(n1717), .X(n1711) );
  nor_x1_sg U12525 ( .A(n6056), .B(n6022), .X(n1718) );
  nor_x1_sg U12526 ( .A(n7060), .B(n9049), .X(n1719) );
  nand_x1_sg U12527 ( .A(n9076), .B(n1966), .X(n1959) );
  nor_x1_sg U12528 ( .A(n6054), .B(n6020), .X(n1967) );
  nor_x1_sg U12529 ( .A(n7058), .B(n9050), .X(n1968) );
  nand_x2_sg U12530 ( .A(n1823), .B(n9075), .X(n1822) );
  nor_x1_sg U12531 ( .A(n7268), .B(n6342), .X(n1823) );
  nand_x1_sg U12532 ( .A(n9075), .B(n1649), .X(n1648) );
  nor_x1_sg U12533 ( .A(n6158), .B(n6012), .X(n1650) );
  nor_x1_sg U12534 ( .A(n7050), .B(n9055), .X(n1651) );
  nand_x1_sg U12535 ( .A(n9075), .B(n1713), .X(n1712) );
  nor_x1_sg U12536 ( .A(n6162), .B(n6016), .X(n1714) );
  nor_x1_sg U12537 ( .A(n7054), .B(n9053), .X(n1715) );
  nand_x1_sg U12538 ( .A(n9075), .B(n1961), .X(n1960) );
  nor_x1_sg U12539 ( .A(n6160), .B(n6014), .X(n1962) );
  nor_x1_sg U12540 ( .A(n7052), .B(n9054), .X(n1963) );
  nand_x1_sg U12541 ( .A(n9212), .B(n1675), .X(n1669) );
  nor_x1_sg U12542 ( .A(n6064), .B(n6024), .X(n1676) );
  nor_x1_sg U12543 ( .A(n6172), .B(n9043), .X(n1677) );
  nand_x1_sg U12544 ( .A(n9212), .B(n1739), .X(n1733) );
  nor_x1_sg U12545 ( .A(n6068), .B(n6028), .X(n1740) );
  nor_x1_sg U12546 ( .A(n6176), .B(n9041), .X(n1741) );
  nand_x1_sg U12547 ( .A(n9212), .B(n1988), .X(n1982) );
  nor_x1_sg U12548 ( .A(n6066), .B(n6026), .X(n1989) );
  nor_x1_sg U12549 ( .A(n6174), .B(n9042), .X(n1990) );
  nand_x1_sg U12550 ( .A(n5958), .B(n9065), .X(n2053) );
  nand_x1_sg U12551 ( .A(n9057), .B(n5956), .X(n2069) );
  nand_x1_sg U12552 ( .A(n9060), .B(n5954), .X(n2057) );
  nand_x1_sg U12553 ( .A(n5962), .B(n9064), .X(n2036) );
  nand_x1_sg U12554 ( .A(n5960), .B(n9062), .X(n2037) );
  nand_x1_sg U12555 ( .A(n9078), .B(n1590), .X(n1589) );
  nor_x1_sg U12556 ( .A(n6214), .B(n6098), .X(n1591) );
  nor_x1_sg U12557 ( .A(n7128), .B(n9013), .X(n1592) );
  nand_x1_sg U12558 ( .A(n9078), .B(n1639), .X(n1638) );
  nor_x1_sg U12559 ( .A(n6164), .B(n6058), .X(n1640) );
  nor_x1_sg U12560 ( .A(n7062), .B(n9047), .X(n1641) );
  nand_x1_sg U12561 ( .A(n5948), .B(n9078), .X(n1687) );
  nand_x1_sg U12562 ( .A(n9078), .B(n1703), .X(n1702) );
  nor_x1_sg U12563 ( .A(n6168), .B(n6062), .X(n1704) );
  nor_x1_sg U12564 ( .A(n7066), .B(n9045), .X(n1705) );
  nand_x1_sg U12565 ( .A(n9078), .B(n1754), .X(n1753) );
  nor_x1_sg U12566 ( .A(n6212), .B(n6096), .X(n1755) );
  nor_x1_sg U12567 ( .A(n7126), .B(n9014), .X(n1756) );
  nand_x1_sg U12568 ( .A(n9078), .B(n1904), .X(n1903) );
  nor_x1_sg U12569 ( .A(n6210), .B(n6094), .X(n1905) );
  nor_x1_sg U12570 ( .A(n7124), .B(n9015), .X(n1906) );
  nand_x1_sg U12571 ( .A(n9078), .B(n1951), .X(n1950) );
  nor_x1_sg U12572 ( .A(n6166), .B(n6060), .X(n1952) );
  nor_x1_sg U12573 ( .A(n7064), .B(n9046), .X(n1953) );
  inv_x4_sg U12574 ( .A(n1594), .X(n7319) );
  nand_x1_sg U12575 ( .A(n6383), .B(n2063), .X(n2062) );
  nor_x1_sg U12576 ( .A(n2064), .B(n2065), .X(n2063) );
  nor_x1_sg U12577 ( .A(n7158), .B(n3814), .X(n1884) );
  nor_x1_sg U12578 ( .A(n7148), .B(n1845), .X(n1881) );
  nor_x1_sg U12579 ( .A(n7102), .B(n1845), .X(n1842) );
  nand_x2_sg U12580 ( .A(n9056), .B(n9215), .X(n2067) );
  nor_x1_sg U12581 ( .A(n7122), .B(n1876), .X(n1873) );
  nor_x1_sg U12582 ( .A(n7192), .B(n6266), .X(n1820) );
  nor_x1_sg U12583 ( .A(n7074), .B(n6178), .X(n1830) );
  nor_x1_sg U12584 ( .A(n7070), .B(n6170), .X(n1834) );
  nor_x1_sg U12585 ( .A(n7094), .B(n6194), .X(n1850) );
  nor_x1_sg U12586 ( .A(n7084), .B(n6186), .X(n1853) );
  nor_x1_sg U12587 ( .A(n6148), .B(n8997), .X(n1615) );
  nor_x1_sg U12588 ( .A(n6374), .B(n7302), .X(n1616) );
  nor_x1_sg U12589 ( .A(n7212), .B(n6284), .X(n1614) );
  nor_x1_sg U12590 ( .A(n6140), .B(n9001), .X(n1626) );
  nor_x1_sg U12591 ( .A(n6366), .B(n7294), .X(n1627) );
  nor_x1_sg U12592 ( .A(n7204), .B(n6278), .X(n1625) );
  nor_x1_sg U12593 ( .A(n6124), .B(n9021), .X(n1603) );
  nor_x1_sg U12594 ( .A(n6350), .B(n7278), .X(n1604) );
  nor_x1_sg U12595 ( .A(n7198), .B(n6272), .X(n1602) );
  nor_x1_sg U12596 ( .A(n6146), .B(n8998), .X(n1778) );
  nor_x1_sg U12597 ( .A(n6372), .B(n7300), .X(n1779) );
  nor_x1_sg U12598 ( .A(n7210), .B(n6282), .X(n1777) );
  nor_x1_sg U12599 ( .A(n6138), .B(n9002), .X(n1788) );
  nor_x1_sg U12600 ( .A(n6364), .B(n7292), .X(n1789) );
  nor_x1_sg U12601 ( .A(n7202), .B(n6276), .X(n1787) );
  nor_x1_sg U12602 ( .A(n6122), .B(n9022), .X(n1766) );
  nor_x1_sg U12603 ( .A(n6348), .B(n7276), .X(n1767) );
  nor_x1_sg U12604 ( .A(n7196), .B(n6270), .X(n1765) );
  nor_x1_sg U12605 ( .A(n6150), .B(n8992), .X(n1885) );
  nor_x1_sg U12606 ( .A(n6376), .B(n7304), .X(n1886) );
  nor_x1_sg U12607 ( .A(n6142), .B(n9000), .X(n1890) );
  nor_x1_sg U12608 ( .A(n6368), .B(n7296), .X(n1891) );
  nor_x1_sg U12609 ( .A(n7206), .B(n9068), .X(n1889) );
  nor_x1_sg U12610 ( .A(n6132), .B(n9008), .X(n1893) );
  nor_x1_sg U12611 ( .A(n6358), .B(n7286), .X(n1894) );
  nor_x1_sg U12612 ( .A(n6130), .B(n9012), .X(n1862) );
  nor_x1_sg U12613 ( .A(n6356), .B(n7284), .X(n1863) );
  nor_x1_sg U12614 ( .A(n7130), .B(n1833), .X(n1861) );
  nor_x1_sg U12615 ( .A(n6134), .B(n9004), .X(n1865) );
  nor_x1_sg U12616 ( .A(n6360), .B(n7288), .X(n1866) );
  nor_x1_sg U12617 ( .A(n6128), .B(n9016), .X(n1874) );
  nor_x1_sg U12618 ( .A(n6354), .B(n7282), .X(n1875) );
  nor_x1_sg U12619 ( .A(n6126), .B(n9020), .X(n1870) );
  nor_x1_sg U12620 ( .A(n6352), .B(n7280), .X(n1871) );
  nor_x1_sg U12621 ( .A(n6144), .B(n8999), .X(n1928) );
  nor_x1_sg U12622 ( .A(n6370), .B(n7298), .X(n1929) );
  nor_x1_sg U12623 ( .A(n7208), .B(n6280), .X(n1927) );
  nor_x1_sg U12624 ( .A(n6136), .B(n9003), .X(n1938) );
  nor_x1_sg U12625 ( .A(n6362), .B(n7290), .X(n1939) );
  nor_x1_sg U12626 ( .A(n7200), .B(n6274), .X(n1937) );
  nor_x1_sg U12627 ( .A(n6120), .B(n9023), .X(n1916) );
  nor_x1_sg U12628 ( .A(n6346), .B(n7274), .X(n1917) );
  nor_x1_sg U12629 ( .A(n7194), .B(n6268), .X(n1915) );
  nand_x2_sg U12630 ( .A(n1581), .B(n1582), .X(n1580) );
  nand_x1_sg U12631 ( .A(n1632), .B(n9081), .X(n1581) );
  nand_x1_sg U12632 ( .A(n7314), .B(n1583), .X(n1582) );
  nand_x2_sg U12633 ( .A(n1679), .B(n1680), .X(n1579) );
  nand_x1_sg U12634 ( .A(n1696), .B(n9081), .X(n1679) );
  nand_x1_sg U12635 ( .A(n7314), .B(n1681), .X(n1680) );
  nand_x2_sg U12636 ( .A(n1745), .B(n1746), .X(n1744) );
  nand_x1_sg U12637 ( .A(n7314), .B(n1747), .X(n1746) );
  nand_x2_sg U12638 ( .A(n1895), .B(n1896), .X(n1743) );
  nand_x1_sg U12639 ( .A(n1944), .B(n9081), .X(n1895) );
  nand_x1_sg U12640 ( .A(n7314), .B(n1897), .X(n1896) );
  nor_x1_sg U12641 ( .A(n1829), .B(n7072), .X(n1828) );
  nor_x1_sg U12642 ( .A(n1833), .B(n7068), .X(n1832) );
  nor_x1_sg U12643 ( .A(n6264), .B(n7190), .X(n1620) );
  nor_x1_sg U12644 ( .A(n6258), .B(n7184), .X(n1631) );
  nor_x1_sg U12645 ( .A(n6252), .B(n7178), .X(n1608) );
  nor_x1_sg U12646 ( .A(n6242), .B(n7168), .X(n1674) );
  nor_x1_sg U12647 ( .A(n6236), .B(n7162), .X(n1646) );
  nor_x1_sg U12648 ( .A(n6246), .B(n7172), .X(n1738) );
  nor_x1_sg U12649 ( .A(n6240), .B(n7166), .X(n1710) );
  nor_x1_sg U12650 ( .A(n6262), .B(n7188), .X(n1783) );
  nor_x1_sg U12651 ( .A(n6256), .B(n7182), .X(n1793) );
  nor_x1_sg U12652 ( .A(n6250), .B(n7176), .X(n1771) );
  nor_x1_sg U12653 ( .A(n9068), .B(n7092), .X(n1849) );
  nor_x1_sg U12654 ( .A(n9071), .B(n7082), .X(n1852) );
  nor_x1_sg U12655 ( .A(n6324), .B(n7252), .X(n1811) );
  nor_x1_sg U12656 ( .A(n6260), .B(n7186), .X(n1933) );
  nor_x1_sg U12657 ( .A(n6254), .B(n7180), .X(n1943) );
  nor_x1_sg U12658 ( .A(n6248), .B(n7174), .X(n1921) );
  nor_x1_sg U12659 ( .A(n6244), .B(n7170), .X(n1987) );
  nor_x1_sg U12660 ( .A(n6238), .B(n7164), .X(n1958) );
  nand_x1_sg U12661 ( .A(n9217), .B(n2049), .X(n2029) );
  nand_x1_sg U12662 ( .A(n7318), .B(n2031), .X(n2030) );
  nand_x1_sg U12663 ( .A(n7033), .B(n7320), .X(n1799) );
  nand_x2_sg U12664 ( .A(n1799), .B(n9081), .X(n1798) );
  nand_x1_sg U12665 ( .A(n1623), .B(n6042), .X(n1800) );
  nor_x1_sg U12666 ( .A(reset), .B(n9208), .X(n3808) );
  nand_x2_sg U12667 ( .A(n1830), .B(n9040), .X(n1827) );
  nand_x2_sg U12668 ( .A(n1834), .B(n9044), .X(n1831) );
  nand_x2_sg U12669 ( .A(n1850), .B(n9032), .X(n1848) );
  nand_x2_sg U12670 ( .A(n1853), .B(n9036), .X(n1851) );
  nand_x2_sg U12671 ( .A(n2044), .B(n2045), .X(n2043) );
  nand_x1_sg U12672 ( .A(n5966), .B(n9057), .X(n2045) );
  nand_x1_sg U12673 ( .A(n5934), .B(n9216), .X(n2044) );
  nand_x2_sg U12674 ( .A(n2009), .B(n2010), .X(n2008) );
  nand_x1_sg U12675 ( .A(n5982), .B(n9057), .X(n2010) );
  nand_x1_sg U12676 ( .A(n5946), .B(n9216), .X(n2009) );
  nand_x2_sg U12677 ( .A(n2024), .B(n2025), .X(n2023) );
  nand_x1_sg U12678 ( .A(n5974), .B(n9057), .X(n2025) );
  nand_x1_sg U12679 ( .A(n5940), .B(n9216), .X(n2024) );
  nand_x2_sg U12680 ( .A(n1692), .B(n1693), .X(n1691) );
  nand_x1_sg U12681 ( .A(n6000), .B(n9074), .X(n1693) );
  nand_x1_sg U12682 ( .A(n6010), .B(n9073), .X(n1692) );
  nand_x2_sg U12683 ( .A(n1688), .B(n1689), .X(n1684) );
  nand_x1_sg U12684 ( .A(n5998), .B(n9075), .X(n1689) );
  nand_x1_sg U12685 ( .A(n6006), .B(n9076), .X(n1688) );
  nor_x1_sg U12686 ( .A(n6330), .B(n7258), .X(n1593) );
  nor_x1_sg U12687 ( .A(n6336), .B(n7264), .X(n1598) );
  nor_x1_sg U12688 ( .A(n6318), .B(n7246), .X(n1668) );
  nor_x1_sg U12689 ( .A(n6310), .B(n7238), .X(n1664) );
  nor_x1_sg U12690 ( .A(n6304), .B(n7232), .X(n1678) );
  nor_x1_sg U12691 ( .A(n6292), .B(n7220), .X(n1656) );
  nor_x1_sg U12692 ( .A(n6286), .B(n7214), .X(n1652) );
  nor_x1_sg U12693 ( .A(n6298), .B(n7226), .X(n1642) );
  nor_x1_sg U12694 ( .A(n6322), .B(n7250), .X(n1732) );
  nor_x1_sg U12695 ( .A(n6314), .B(n7242), .X(n1728) );
  nor_x1_sg U12696 ( .A(n6308), .B(n7236), .X(n1742) );
  nor_x1_sg U12697 ( .A(n6296), .B(n7224), .X(n1720) );
  nor_x1_sg U12698 ( .A(n6290), .B(n7218), .X(n1716) );
  nor_x1_sg U12699 ( .A(n6302), .B(n7230), .X(n1706) );
  nor_x1_sg U12700 ( .A(n6328), .B(n7256), .X(n1757) );
  nor_x1_sg U12701 ( .A(n6334), .B(n7262), .X(n1761) );
  nor_x1_sg U12702 ( .A(n6338), .B(n7266), .X(n1883) );
  nor_x1_sg U12703 ( .A(n6316), .B(n7244), .X(n1844) );
  nor_x1_sg U12704 ( .A(n6326), .B(n7254), .X(n1907) );
  nor_x1_sg U12705 ( .A(n6332), .B(n7260), .X(n1911) );
  nor_x1_sg U12706 ( .A(n6320), .B(n7248), .X(n1981) );
  nor_x1_sg U12707 ( .A(n6312), .B(n7240), .X(n1977) );
  nor_x1_sg U12708 ( .A(n6306), .B(n7234), .X(n1991) );
  nor_x1_sg U12709 ( .A(n6294), .B(n7222), .X(n1969) );
  nor_x1_sg U12710 ( .A(n6288), .B(n7216), .X(n1964) );
  nor_x1_sg U12711 ( .A(n6300), .B(n7228), .X(n1954) );
  nand_x2_sg U12712 ( .A(n2053), .B(n2054), .X(n2052) );
  nand_x1_sg U12713 ( .A(n7025), .B(n9214), .X(n2054) );
  nand_x2_sg U12714 ( .A(n2047), .B(n2048), .X(n2042) );
  nand_x1_sg U12715 ( .A(n5932), .B(n9063), .X(n2048) );
  nand_x1_sg U12716 ( .A(n5964), .B(n9060), .X(n2047) );
  nand_x2_sg U12717 ( .A(n2011), .B(n2012), .X(n2007) );
  nand_x1_sg U12718 ( .A(n5944), .B(n9063), .X(n2012) );
  nand_x1_sg U12719 ( .A(n5980), .B(n9060), .X(n2011) );
  nand_x2_sg U12720 ( .A(n2026), .B(n2027), .X(n2022) );
  nand_x1_sg U12721 ( .A(n5938), .B(n9063), .X(n2027) );
  nand_x1_sg U12722 ( .A(n5972), .B(n9060), .X(n2026) );
  nand_x2_sg U12723 ( .A(n2040), .B(n2041), .X(n2034) );
  nand_x1_sg U12724 ( .A(n7027), .B(n9214), .X(n2041) );
  nand_x1_sg U12725 ( .A(n5968), .B(n9065), .X(n2040) );
  nand_x2_sg U12726 ( .A(n2005), .B(n2006), .X(n2001) );
  nand_x1_sg U12727 ( .A(n7031), .B(n9214), .X(n2006) );
  nand_x1_sg U12728 ( .A(n5984), .B(n9065), .X(n2005) );
  nand_x2_sg U12729 ( .A(n2020), .B(n2021), .X(n2016) );
  nand_x1_sg U12730 ( .A(n7029), .B(n9214), .X(n2021) );
  nand_x1_sg U12731 ( .A(n5976), .B(n9065), .X(n2020) );
  nand_x2_sg U12732 ( .A(n1694), .B(n1695), .X(n1690) );
  nand_x1_sg U12733 ( .A(n6046), .B(n1623), .X(n1695) );
  nand_x1_sg U12734 ( .A(n6008), .B(n9212), .X(n1694) );
  nand_x2_sg U12735 ( .A(n2003), .B(n2004), .X(n2002) );
  nand_x1_sg U12736 ( .A(n5942), .B(n9062), .X(n2004) );
  nand_x1_sg U12737 ( .A(n5978), .B(n9064), .X(n2003) );
  nand_x2_sg U12738 ( .A(n2018), .B(n2019), .X(n2017) );
  nand_x1_sg U12739 ( .A(n5936), .B(n9062), .X(n2019) );
  nand_x1_sg U12740 ( .A(n5970), .B(n9064), .X(n2018) );
  nor_x1_sg U12741 ( .A(n6226), .B(n6110), .X(n1596) );
  nor_x1_sg U12742 ( .A(n7144), .B(n9005), .X(n1597) );
  nor_x1_sg U12743 ( .A(n6224), .B(n6108), .X(n1759) );
  nor_x1_sg U12744 ( .A(n7142), .B(n9006), .X(n1760) );
  nor_x1_sg U12745 ( .A(n6222), .B(n6106), .X(n1909) );
  nor_x1_sg U12746 ( .A(n7140), .B(n9007), .X(n1910) );
  nor_x1_sg U12747 ( .A(n7112), .B(n9024), .X(n1810) );
  nor_x1_sg U12748 ( .A(n6202), .B(n3814), .X(n1809) );
  nand_x1_sg U12749 ( .A(n1838), .B(n6004), .X(n1837) );
  nand_x1_sg U12750 ( .A(n1839), .B(n5996), .X(n1836) );
  nand_x2_sg U12751 ( .A(n1824), .B(n9052), .X(n1821) );
  nor_x1_sg U12752 ( .A(n7272), .B(n6344), .X(n1824) );
  nor_x1_sg U12753 ( .A(n6232), .B(n6116), .X(n1618) );
  nor_x1_sg U12754 ( .A(n7156), .B(n8993), .X(n1619) );
  nor_x1_sg U12755 ( .A(n6220), .B(n6104), .X(n1629) );
  nor_x1_sg U12756 ( .A(n7136), .B(n9009), .X(n1630) );
  nor_x1_sg U12757 ( .A(n6208), .B(n6092), .X(n1606) );
  nor_x1_sg U12758 ( .A(n7120), .B(n9017), .X(n1607) );
  nor_x1_sg U12759 ( .A(n6188), .B(n6076), .X(n1672) );
  nor_x1_sg U12760 ( .A(n7086), .B(n9035), .X(n1673) );
  nor_x1_sg U12761 ( .A(n6180), .B(n6070), .X(n1644) );
  nor_x1_sg U12762 ( .A(n7076), .B(n9039), .X(n1645) );
  nor_x1_sg U12763 ( .A(n6192), .B(n6080), .X(n1736) );
  nor_x1_sg U12764 ( .A(n7090), .B(n9033), .X(n1737) );
  nor_x1_sg U12765 ( .A(n6184), .B(n6074), .X(n1708) );
  nor_x1_sg U12766 ( .A(n7080), .B(n9037), .X(n1709) );
  nor_x1_sg U12767 ( .A(n6230), .B(n6114), .X(n1781) );
  nor_x1_sg U12768 ( .A(n7154), .B(n8994), .X(n1782) );
  nor_x1_sg U12769 ( .A(n6218), .B(n6102), .X(n1791) );
  nor_x1_sg U12770 ( .A(n7134), .B(n9010), .X(n1792) );
  nor_x1_sg U12771 ( .A(n6206), .B(n6090), .X(n1769) );
  nor_x1_sg U12772 ( .A(n7118), .B(n9018), .X(n1770) );
  nor_x1_sg U12773 ( .A(n6228), .B(n6112), .X(n1931) );
  nor_x1_sg U12774 ( .A(n7152), .B(n8995), .X(n1932) );
  nor_x1_sg U12775 ( .A(n6216), .B(n6100), .X(n1941) );
  nor_x1_sg U12776 ( .A(n7132), .B(n9011), .X(n1942) );
  nor_x1_sg U12777 ( .A(n6204), .B(n6088), .X(n1919) );
  nor_x1_sg U12778 ( .A(n7116), .B(n9019), .X(n1920) );
  nor_x1_sg U12779 ( .A(n6190), .B(n6078), .X(n1985) );
  nor_x1_sg U12780 ( .A(n7088), .B(n9034), .X(n1986) );
  nor_x1_sg U12781 ( .A(n6182), .B(n6072), .X(n1956) );
  nor_x1_sg U12782 ( .A(n7078), .B(n9038), .X(n1957) );
  nand_x2_sg U12783 ( .A(n1840), .B(n1841), .X(n1805) );
  nor_x1_sg U12784 ( .A(n1846), .B(n1847), .X(n1840) );
  nor_x1_sg U12785 ( .A(n7104), .B(n9028), .X(n1843) );
  nand_x2_sg U12786 ( .A(n1879), .B(n1880), .X(n1878) );
  nor_x1_sg U12787 ( .A(n7150), .B(n8996), .X(n1882) );
  nand_x2_sg U12788 ( .A(n1887), .B(n1888), .X(n1877) );
  nor_x1_sg U12789 ( .A(n7138), .B(n1829), .X(n1892) );
  nand_x2_sg U12790 ( .A(n1859), .B(n1860), .X(n1858) );
  nor_x1_sg U12791 ( .A(n7146), .B(n9071), .X(n1864) );
  nand_x2_sg U12792 ( .A(n1867), .B(n1868), .X(n1857) );
  nor_x1_sg U12793 ( .A(n7114), .B(n1872), .X(n1869) );
  inv_x8_sg U12794 ( .A(n7319), .X(n7320) );
  inv_x8_sg U12795 ( .A(n3101), .X(n9214) );
  inv_x8_sg U12796 ( .A(n5992), .X(n7321) );
  inv_x8_sg U12797 ( .A(n7322), .X(n7323) );
  inv_x8_sg U12798 ( .A(n7374), .X(n7324) );
  inv_x8_sg U12799 ( .A(n7372), .X(n7325) );
  inv_x8_sg U12800 ( .A(n7370), .X(n7326) );
  inv_x8_sg U12801 ( .A(n7364), .X(n7327) );
  inv_x8_sg U12802 ( .A(n7362), .X(n7328) );
  inv_x8_sg U12803 ( .A(n7360), .X(n7329) );
  inv_x8_sg U12804 ( .A(n7354), .X(n7330) );
  inv_x8_sg U12805 ( .A(n7352), .X(n7331) );
  inv_x8_sg U12806 ( .A(n7350), .X(n7332) );
  inv_x8_sg U12807 ( .A(n7343), .X(n7333) );
  inv_x8_sg U12808 ( .A(n7341), .X(n7334) );
  inv_x8_sg U12809 ( .A(n7339), .X(n7335) );
  inv_x8_sg U12810 ( .A(n773), .X(n7336) );
  inv_x8_sg U12811 ( .A(n7336), .X(n7337) );
  inv_x8_sg U12812 ( .A(n7338), .X(n7339) );
  inv_x8_sg U12813 ( .A(n7340), .X(n7341) );
  inv_x8_sg U12814 ( .A(n7342), .X(n7343) );
  inv_x8_sg U12815 ( .A(n7344), .X(n7345) );
  inv_x8_sg U12816 ( .A(n7345), .X(n7346) );
  inv_x8_sg U12817 ( .A(n778), .X(n7347) );
  inv_x8_sg U12818 ( .A(n7347), .X(n7348) );
  inv_x8_sg U12819 ( .A(n7349), .X(n7350) );
  inv_x8_sg U12820 ( .A(n7351), .X(n7352) );
  inv_x8_sg U12821 ( .A(n7353), .X(n7354) );
  inv_x8_sg U12822 ( .A(n782), .X(n7355) );
  inv_x8_sg U12823 ( .A(n7355), .X(n7356) );
  inv_x8_sg U12824 ( .A(n783), .X(n7357) );
  inv_x8_sg U12825 ( .A(n7357), .X(n7358) );
  inv_x8_sg U12826 ( .A(n7359), .X(n7360) );
  inv_x8_sg U12827 ( .A(n7361), .X(n7362) );
  inv_x8_sg U12828 ( .A(n7363), .X(n7364) );
  inv_x8_sg U12829 ( .A(n787), .X(n7365) );
  inv_x8_sg U12830 ( .A(n7365), .X(n7366) );
  inv_x8_sg U12831 ( .A(n788), .X(n7367) );
  inv_x8_sg U12832 ( .A(n7367), .X(n7368) );
  inv_x8_sg U12833 ( .A(n7369), .X(n7370) );
  inv_x8_sg U12834 ( .A(n7371), .X(n7372) );
  inv_x8_sg U12835 ( .A(n7373), .X(n7374) );
  inv_x8_sg U12836 ( .A(n6381), .X(n7375) );
  inv_x8_sg U12837 ( .A(n7376), .X(n7377) );
  inv_x8_sg U12838 ( .A(n7378), .X(n7379) );
  nand_x8_sg U12839 ( .A(n1510), .B(n1511), .X(n7380) );
  nand_x8_sg U12840 ( .A(n1510), .B(n1511), .X(n7381) );
  nand_x8_sg U12841 ( .A(n1511), .B(n1512), .X(n7382) );
  nand_x8_sg U12842 ( .A(n1511), .B(n1512), .X(n7383) );
  inv_x8_sg U12843 ( .A(n7386), .X(n7387) );
  inv_x8_sg U12844 ( .A(n7388), .X(n7389) );
  nand_x8_sg U12845 ( .A(n7392), .B(n7568), .X(n7390) );
  nand_x8_sg U12846 ( .A(n7392), .B(n7568), .X(n7391) );
  inv_x8_sg U12847 ( .A(n4196), .X(n7392) );
  inv_x8_sg U12848 ( .A(n4192), .X(n7393) );
  nor_x8_sg U12849 ( .A(n4192), .B(n7569), .X(n7394) );
  nor_x8_sg U12850 ( .A(n4192), .B(n7569), .X(n7395) );
  nor_x8_sg U12851 ( .A(n4192), .B(n7569), .X(n4186) );
  nor_x8_sg U12852 ( .A(n4184), .B(n4196), .X(n7396) );
  nor_x8_sg U12853 ( .A(n4184), .B(n4196), .X(n7397) );
  nor_x8_sg U12854 ( .A(n4184), .B(n4196), .X(n894) );
  inv_x8_sg U12855 ( .A(n6152), .X(n7398) );
  inv_x8_sg U12856 ( .A(n7399), .X(n7400) );
  inv_x8_sg U12857 ( .A(n793), .X(n7401) );
  inv_x8_sg U12858 ( .A(n7401), .X(n7402) );
  inv_x8_sg U12859 ( .A(n7422), .X(n7403) );
  inv_x8_sg U12860 ( .A(n7448), .X(n7404) );
  inv_x8_sg U12861 ( .A(n7457), .X(n7405) );
  inv_x8_sg U12862 ( .A(n7510), .X(n7406) );
  inv_x8_sg U12863 ( .A(n7464), .X(n7407) );
  inv_x8_sg U12864 ( .A(n7497), .X(n7408) );
  inv_x8_sg U12865 ( .A(n7500), .X(n7409) );
  inv_x8_sg U12866 ( .A(n7507), .X(n7410) );
  inv_x8_sg U12867 ( .A(n7459), .X(n7411) );
  inv_x8_sg U12868 ( .A(n7461), .X(n7412) );
  inv_x8_sg U12869 ( .A(n7512), .X(n7413) );
  inv_x8_sg U12870 ( .A(n7514), .X(n7414) );
  inv_x8_sg U12871 ( .A(n7502), .X(n7415) );
  inv_x8_sg U12872 ( .A(n7503), .X(n7416) );
  inv_x8_sg U12873 ( .A(n7516), .X(n7417) );
  inv_x8_sg U12874 ( .A(n7518), .X(n7418) );
  inv_x8_sg U12875 ( .A(n3930), .X(n7419) );
  nor_x8_sg U12876 ( .A(n9245), .B(n3930), .X(n4182) );
  inv_x8_sg U12877 ( .A(n4407), .X(n7420) );
  inv_x8_sg U12878 ( .A(n7420), .X(n7421) );
  inv_x8_sg U12879 ( .A(n7420), .X(n7422) );
  inv_x8_sg U12880 ( .A(n7425), .X(n7426) );
  nand_x8_sg U12881 ( .A(n7570), .B(n7558), .X(n7427) );
  nand_x8_sg U12882 ( .A(n7570), .B(n7558), .X(n7428) );
  nand_x8_sg U12883 ( .A(n7570), .B(n7323), .X(n7429) );
  nor_x8_sg U12884 ( .A(n4297), .B(n7559), .X(n7430) );
  nor_x8_sg U12885 ( .A(n4297), .B(n7559), .X(n7431) );
  nor_x8_sg U12886 ( .A(n4297), .B(n7559), .X(n4428) );
  nand_x8_sg U12887 ( .A(n9240), .B(n5242), .X(n7432) );
  nand_x8_sg U12888 ( .A(n9240), .B(n5242), .X(n7433) );
  nand_x8_sg U12889 ( .A(n9240), .B(n5241), .X(n7434) );
  nand_x8_sg U12890 ( .A(n9240), .B(n5241), .X(n7435) );
  inv_x8_sg U12891 ( .A(n7436), .X(n7437) );
  inv_x8_sg U12892 ( .A(n7438), .X(n7439) );
  inv_x8_sg U12893 ( .A(n7440), .X(n7441) );
  inv_x8_sg U12894 ( .A(n7442), .X(n7443) );
  inv_x8_sg U12895 ( .A(n7444), .X(n7445) );
  inv_x8_sg U12896 ( .A(n4020), .X(n7446) );
  inv_x8_sg U12897 ( .A(n7446), .X(n7447) );
  inv_x8_sg U12898 ( .A(n7446), .X(n7448) );
  inv_x8_sg U12899 ( .A(n7449), .X(n7450) );
  inv_x8_sg U12900 ( .A(n7451), .X(n7452) );
  inv_x8_sg U12901 ( .A(n7453), .X(n7454) );
  inv_x8_sg U12902 ( .A(n4102), .X(n7455) );
  inv_x8_sg U12903 ( .A(n7455), .X(n7456) );
  inv_x8_sg U12904 ( .A(n7455), .X(n7457) );
  nand_x8_sg U12905 ( .A(n5064), .B(n3928), .X(n7458) );
  nand_x8_sg U12906 ( .A(n5064), .B(n3928), .X(n7459) );
  nand_x8_sg U12907 ( .A(n5064), .B(n3886), .X(n7460) );
  nand_x8_sg U12908 ( .A(n5064), .B(n3886), .X(n7461) );
  inv_x8_sg U12909 ( .A(n4401), .X(n7462) );
  inv_x8_sg U12910 ( .A(n7462), .X(n7463) );
  inv_x8_sg U12911 ( .A(n7462), .X(n7464) );
  inv_x8_sg U12912 ( .A(n7465), .X(n7466) );
  inv_x8_sg U12913 ( .A(n7467), .X(n7468) );
  inv_x8_sg U12914 ( .A(n7469), .X(n7470) );
  inv_x8_sg U12915 ( .A(n7471), .X(n7472) );
  inv_x8_sg U12916 ( .A(n7473), .X(n7474) );
  inv_x8_sg U12917 ( .A(n7475), .X(n7476) );
  inv_x8_sg U12918 ( .A(n7477), .X(n7478) );
  inv_x8_sg U12919 ( .A(n7479), .X(n7480) );
  inv_x8_sg U12920 ( .A(n7481), .X(n7482) );
  inv_x8_sg U12921 ( .A(n7483), .X(n7484) );
  inv_x8_sg U12922 ( .A(n7485), .X(n7486) );
  inv_x8_sg U12923 ( .A(n7487), .X(n7488) );
  inv_x8_sg U12924 ( .A(n7489), .X(n7490) );
  inv_x8_sg U12925 ( .A(n7491), .X(n7492) );
  inv_x8_sg U12926 ( .A(n7493), .X(n7494) );
  inv_x8_sg U12927 ( .A(n4352), .X(n7495) );
  inv_x8_sg U12928 ( .A(n7495), .X(n7496) );
  inv_x8_sg U12929 ( .A(n7495), .X(n7497) );
  inv_x8_sg U12930 ( .A(n4310), .X(n7498) );
  inv_x8_sg U12931 ( .A(n7498), .X(n7499) );
  inv_x8_sg U12932 ( .A(n7498), .X(n7500) );
  nand_x8_sg U12933 ( .A(n3928), .B(n4249), .X(n7501) );
  nand_x8_sg U12934 ( .A(n3928), .B(n4249), .X(n7502) );
  nand_x8_sg U12935 ( .A(n3886), .B(n4249), .X(n7503) );
  nand_x8_sg U12936 ( .A(n3886), .B(n4249), .X(n7504) );
  inv_x8_sg U12937 ( .A(n4139), .X(n7505) );
  inv_x8_sg U12938 ( .A(n7505), .X(n7506) );
  inv_x8_sg U12939 ( .A(n7505), .X(n7507) );
  inv_x8_sg U12940 ( .A(n4059), .X(n7508) );
  inv_x8_sg U12941 ( .A(n7508), .X(n7509) );
  inv_x8_sg U12942 ( .A(n7508), .X(n7510) );
  nand_x8_sg U12943 ( .A(n3974), .B(n3886), .X(n7511) );
  nand_x8_sg U12944 ( .A(n3974), .B(n3886), .X(n7512) );
  nand_x8_sg U12945 ( .A(n3974), .B(n3928), .X(n7513) );
  nand_x8_sg U12946 ( .A(n3974), .B(n3928), .X(n7514) );
  nand_x8_sg U12947 ( .A(n9195), .B(n3928), .X(n7515) );
  nand_x8_sg U12948 ( .A(n9195), .B(n3928), .X(n7516) );
  nand_x8_sg U12949 ( .A(n9195), .B(n3886), .X(n7517) );
  nand_x8_sg U12950 ( .A(n9195), .B(n3886), .X(n7518) );
  inv_x8_sg U12951 ( .A(n6154), .X(n7519) );
  inv_x8_sg U12952 ( .A(n7519), .X(n7520) );
  inv_x8_sg U12953 ( .A(n7521), .X(n7522) );
  inv_x8_sg U12954 ( .A(n7524), .X(n7523) );
  inv_x8_sg U12955 ( .A(n4182), .X(n7526) );
  inv_x8_sg U12956 ( .A(n7532), .X(n7527) );
  inv_x8_sg U12957 ( .A(n7532), .X(n7528) );
  inv_x8_sg U12958 ( .A(n7532), .X(n7529) );
  inv_x8_sg U12959 ( .A(n7532), .X(n7530) );
  inv_x8_sg U12960 ( .A(n7532), .X(n7531) );
  inv_x8_sg U12961 ( .A(n7536), .X(n7532) );
  inv_x8_sg U12962 ( .A(n7532), .X(n7533) );
  inv_x8_sg U12963 ( .A(n7532), .X(n7534) );
  inv_x8_sg U12964 ( .A(n7532), .X(n7535) );
  inv_x8_sg U12965 ( .A(n7537), .X(n7536) );
  inv_x8_sg U12966 ( .A(n7553), .X(n7542) );
  inv_x8_sg U12967 ( .A(n7553), .X(n7543) );
  inv_x8_sg U12968 ( .A(n7553), .X(n7544) );
  inv_x8_sg U12969 ( .A(n7553), .X(n7545) );
  inv_x8_sg U12970 ( .A(n7553), .X(n7546) );
  inv_x8_sg U12971 ( .A(n7553), .X(n7547) );
  inv_x8_sg U12972 ( .A(n7553), .X(n7548) );
  inv_x8_sg U12973 ( .A(n7553), .X(n7549) );
  inv_x8_sg U12974 ( .A(n7553), .X(n7550) );
  inv_x8_sg U12975 ( .A(n7553), .X(n7551) );
  inv_x8_sg U12976 ( .A(n7553), .X(n7552) );
  inv_x8_sg U12977 ( .A(n7554), .X(n7553) );
  inv_x8_sg U12978 ( .A(n7555), .X(n7554) );
  inv_x8_sg U12979 ( .A(n7559), .X(n7558) );
  inv_x8_sg U12980 ( .A(n5994), .X(n7559) );
  inv_x8_sg U12981 ( .A(n7562), .X(n7560) );
  inv_x8_sg U12982 ( .A(n7563), .X(n7561) );
  inv_x8_sg U12983 ( .A(n7563), .X(n7562) );
  inv_x8_sg U12984 ( .A(n7039), .X(n7563) );
  inv_x8_sg U12985 ( .A(n7565), .X(n7564) );
  inv_x8_sg U12986 ( .A(n7567), .X(n7566) );
  inv_x4_sg U12987 ( .A(n5895), .X(n7567) );
  inv_x8_sg U12988 ( .A(n7569), .X(n7568) );
  inv_x8_sg U12989 ( .A(n6002), .X(n7569) );
  inv_x8_sg U12990 ( .A(n7571), .X(n7570) );
  inv_x8_sg U12991 ( .A(n6156), .X(n7571) );
  inv_x2_sg U14408 ( .A(n1593), .X(n9013) );
  inv_x2_sg U14409 ( .A(n1598), .X(n9005) );
  inv_x2_sg U14410 ( .A(n1604), .X(n9021) );
  inv_x2_sg U14411 ( .A(n1608), .X(n9017) );
  inv_x2_sg U14412 ( .A(n1616), .X(n8997) );
  inv_x2_sg U14413 ( .A(n1620), .X(n8993) );
  inv_x2_sg U14414 ( .A(n1627), .X(n9001) );
  inv_x2_sg U14415 ( .A(n1631), .X(n9009) );
  inv_x2_sg U14416 ( .A(n1642), .X(n9047) );
  inv_x2_sg U14417 ( .A(n1646), .X(n9039) );
  inv_x2_sg U14418 ( .A(n1652), .X(n9055) );
  inv_x2_sg U14419 ( .A(n1656), .X(n9051) );
  inv_x2_sg U14420 ( .A(n1664), .X(n9031) );
  inv_x2_sg U14421 ( .A(n1668), .X(n9027) );
  inv_x2_sg U14422 ( .A(n1674), .X(n9035) );
  inv_x2_sg U14423 ( .A(n1678), .X(n9043) );
  inv_x2_sg U14424 ( .A(n1706), .X(n9045) );
  inv_x2_sg U14425 ( .A(n1710), .X(n9037) );
  inv_x2_sg U14426 ( .A(n1716), .X(n9053) );
  inv_x2_sg U14427 ( .A(n1720), .X(n9049) );
  inv_x2_sg U14428 ( .A(n1728), .X(n9029) );
  inv_x2_sg U14429 ( .A(n1732), .X(n9025) );
  inv_x2_sg U14430 ( .A(n1738), .X(n9033) );
  inv_x2_sg U14431 ( .A(n1742), .X(n9041) );
  inv_x2_sg U14432 ( .A(n1757), .X(n9014) );
  inv_x2_sg U14433 ( .A(n1761), .X(n9006) );
  inv_x2_sg U14434 ( .A(n1767), .X(n9022) );
  inv_x2_sg U14435 ( .A(n1771), .X(n9018) );
  inv_x2_sg U14436 ( .A(n1779), .X(n8998) );
  inv_x2_sg U14437 ( .A(n1783), .X(n8994) );
  inv_x2_sg U14438 ( .A(n1789), .X(n9002) );
  inv_x2_sg U14439 ( .A(n1793), .X(n9010) );
  inv_x2_sg U14440 ( .A(n1800), .X(n9070) );
  inv_x2_sg U14441 ( .A(n1811), .X(n9024) );
  inv_x2_sg U14442 ( .A(n1828), .X(n9080) );
  inv_x2_sg U14443 ( .A(n1832), .X(n9079) );
  inv_x2_sg U14444 ( .A(n1844), .X(n9028) );
  inv_x2_sg U14445 ( .A(n1849), .X(n9069) );
  inv_x2_sg U14446 ( .A(n1852), .X(n9072) );
  inv_x2_sg U14447 ( .A(n1863), .X(n9012) );
  inv_x2_sg U14448 ( .A(n1866), .X(n9004) );
  inv_x2_sg U14449 ( .A(n1871), .X(n9020) );
  inv_x2_sg U14450 ( .A(n1875), .X(n9016) );
  inv_x2_sg U14451 ( .A(n1883), .X(n8996) );
  inv_x2_sg U14452 ( .A(n1886), .X(n8992) );
  inv_x2_sg U14453 ( .A(n1891), .X(n9000) );
  inv_x2_sg U14454 ( .A(n1894), .X(n9008) );
  inv_x2_sg U14455 ( .A(n1907), .X(n9015) );
  inv_x2_sg U14456 ( .A(n1911), .X(n9007) );
  inv_x2_sg U14457 ( .A(n1917), .X(n9023) );
  inv_x2_sg U14458 ( .A(n1921), .X(n9019) );
  inv_x2_sg U14459 ( .A(n1929), .X(n8999) );
  inv_x2_sg U14460 ( .A(n1933), .X(n8995) );
  inv_x2_sg U14461 ( .A(n1939), .X(n9003) );
  inv_x2_sg U14462 ( .A(n1943), .X(n9011) );
  inv_x2_sg U14463 ( .A(n1954), .X(n9046) );
  inv_x2_sg U14464 ( .A(n1958), .X(n9038) );
  inv_x2_sg U14465 ( .A(n1964), .X(n9054) );
  inv_x2_sg U14466 ( .A(n1969), .X(n9050) );
  inv_x2_sg U14467 ( .A(n1977), .X(n9030) );
  inv_x2_sg U14468 ( .A(n1981), .X(n9026) );
  inv_x2_sg U14469 ( .A(n1987), .X(n9034) );
  inv_x2_sg U14470 ( .A(n1991), .X(n9042) );
  inv_x2_sg U14471 ( .A(n2057), .X(n9061) );
  inv_x2_sg U14472 ( .A(n2062), .X(n9059) );
  inv_x2_sg U14473 ( .A(n2069), .X(n9058) );
  inv_x2_sg U14474 ( .A(n1992), .X(n9185) );
  inv_x2_sg U14475 ( .A(\i_im[13][1] ), .X(n9163) );
  inv_x2_sg U14476 ( .A(\i_im[12][1] ), .X(n9143) );
  inv_x2_sg U14477 ( .A(\i_im[6][1] ), .X(n9103) );
  inv_x2_sg U14478 ( .A(n923), .X(n9083) );
  inv_x2_sg U14479 ( .A(n925), .X(n9123) );
  inv_x2_sg U14480 ( .A(\i_im[13][2] ), .X(n9164) );
  inv_x2_sg U14481 ( .A(\i_im[12][2] ), .X(n9144) );
  inv_x2_sg U14482 ( .A(\i_im[6][2] ), .X(n9104) );
  inv_x2_sg U14483 ( .A(n956), .X(n9084) );
  inv_x2_sg U14484 ( .A(n958), .X(n9124) );
  inv_x2_sg U14485 ( .A(\i_im[13][3] ), .X(n9165) );
  inv_x2_sg U14486 ( .A(\i_im[12][3] ), .X(n9145) );
  inv_x2_sg U14487 ( .A(\i_im[6][3] ), .X(n9105) );
  inv_x2_sg U14488 ( .A(n989), .X(n9085) );
  inv_x2_sg U14489 ( .A(n991), .X(n9125) );
  inv_x2_sg U14490 ( .A(\i_im[13][4] ), .X(n9166) );
  inv_x2_sg U14491 ( .A(\i_im[12][4] ), .X(n9146) );
  inv_x2_sg U14492 ( .A(\i_im[6][4] ), .X(n9106) );
  inv_x2_sg U14493 ( .A(n1022), .X(n9086) );
  inv_x2_sg U14494 ( .A(n1024), .X(n9126) );
  inv_x2_sg U14495 ( .A(\i_im[13][5] ), .X(n9167) );
  inv_x2_sg U14496 ( .A(\i_im[12][5] ), .X(n9147) );
  inv_x2_sg U14497 ( .A(\i_im[6][5] ), .X(n9107) );
  inv_x2_sg U14498 ( .A(n1058), .X(n9087) );
  inv_x2_sg U14499 ( .A(n1060), .X(n9127) );
  inv_x2_sg U14500 ( .A(\i_im[13][6] ), .X(n9168) );
  inv_x2_sg U14501 ( .A(\i_im[12][6] ), .X(n9148) );
  inv_x2_sg U14502 ( .A(\i_im[6][6] ), .X(n9108) );
  inv_x2_sg U14503 ( .A(n1091), .X(n9088) );
  inv_x2_sg U14504 ( .A(n1093), .X(n9128) );
  inv_x2_sg U14505 ( .A(\i_im[13][7] ), .X(n9169) );
  inv_x2_sg U14506 ( .A(\i_im[12][7] ), .X(n9149) );
  inv_x2_sg U14507 ( .A(\i_im[6][7] ), .X(n9109) );
  inv_x2_sg U14508 ( .A(n1124), .X(n9089) );
  inv_x2_sg U14509 ( .A(n1126), .X(n9129) );
  inv_x2_sg U14510 ( .A(\i_im[13][8] ), .X(n9170) );
  inv_x2_sg U14511 ( .A(\i_im[12][8] ), .X(n9150) );
  inv_x2_sg U14512 ( .A(\i_im[6][8] ), .X(n9110) );
  inv_x2_sg U14513 ( .A(n1157), .X(n9090) );
  inv_x2_sg U14514 ( .A(n1159), .X(n9130) );
  inv_x2_sg U14515 ( .A(\i_im[13][9] ), .X(n9171) );
  inv_x2_sg U14516 ( .A(\i_im[12][9] ), .X(n9151) );
  inv_x2_sg U14517 ( .A(\i_im[6][9] ), .X(n9111) );
  inv_x2_sg U14518 ( .A(n1190), .X(n9091) );
  inv_x2_sg U14519 ( .A(n1192), .X(n9131) );
  inv_x2_sg U14520 ( .A(\i_im[13][10] ), .X(n9172) );
  inv_x2_sg U14521 ( .A(\i_im[12][10] ), .X(n9152) );
  inv_x2_sg U14522 ( .A(\i_im[6][10] ), .X(n9112) );
  inv_x2_sg U14523 ( .A(n1228), .X(n9092) );
  inv_x2_sg U14524 ( .A(n1230), .X(n9132) );
  inv_x2_sg U14525 ( .A(\i_im[13][11] ), .X(n9173) );
  inv_x2_sg U14526 ( .A(\i_im[12][11] ), .X(n9153) );
  inv_x2_sg U14527 ( .A(\i_im[6][11] ), .X(n9113) );
  inv_x2_sg U14528 ( .A(n1261), .X(n9093) );
  inv_x2_sg U14529 ( .A(n1263), .X(n9133) );
  inv_x2_sg U14530 ( .A(\i_im[13][12] ), .X(n9174) );
  inv_x2_sg U14531 ( .A(\i_im[12][12] ), .X(n9154) );
  inv_x2_sg U14532 ( .A(\i_im[6][12] ), .X(n9114) );
  inv_x2_sg U14533 ( .A(n1294), .X(n9094) );
  inv_x2_sg U14534 ( .A(n1296), .X(n9134) );
  inv_x2_sg U14535 ( .A(\i_im[13][13] ), .X(n9175) );
  inv_x2_sg U14536 ( .A(\i_im[12][13] ), .X(n9155) );
  inv_x2_sg U14537 ( .A(\i_im[6][13] ), .X(n9115) );
  inv_x2_sg U14538 ( .A(n1327), .X(n9095) );
  inv_x2_sg U14539 ( .A(n1329), .X(n9135) );
  inv_x2_sg U14540 ( .A(\i_im[13][14] ), .X(n9176) );
  inv_x2_sg U14541 ( .A(\i_im[12][14] ), .X(n9156) );
  inv_x2_sg U14542 ( .A(\i_im[6][14] ), .X(n9116) );
  inv_x2_sg U14543 ( .A(n1360), .X(n9096) );
  inv_x2_sg U14544 ( .A(n1362), .X(n9136) );
  inv_x2_sg U14545 ( .A(\i_im[13][15] ), .X(n9177) );
  inv_x2_sg U14546 ( .A(\i_im[12][15] ), .X(n9157) );
  inv_x2_sg U14547 ( .A(\i_im[6][15] ), .X(n9117) );
  inv_x2_sg U14548 ( .A(n1396), .X(n9097) );
  inv_x2_sg U14549 ( .A(n1398), .X(n9137) );
  inv_x2_sg U14550 ( .A(\i_im[13][16] ), .X(n9178) );
  inv_x2_sg U14551 ( .A(\i_im[12][16] ), .X(n9158) );
  inv_x2_sg U14552 ( .A(\i_im[6][16] ), .X(n9118) );
  inv_x2_sg U14553 ( .A(n1429), .X(n9098) );
  inv_x2_sg U14554 ( .A(n1431), .X(n9138) );
  inv_x2_sg U14555 ( .A(\i_im[13][17] ), .X(n9179) );
  inv_x2_sg U14556 ( .A(\i_im[12][17] ), .X(n9159) );
  inv_x2_sg U14557 ( .A(\i_im[6][17] ), .X(n9119) );
  inv_x2_sg U14558 ( .A(n1462), .X(n9099) );
  inv_x2_sg U14559 ( .A(n1464), .X(n9139) );
  inv_x2_sg U14560 ( .A(\i_im[13][18] ), .X(n9180) );
  inv_x2_sg U14561 ( .A(\i_im[12][18] ), .X(n9160) );
  inv_x2_sg U14562 ( .A(\i_im[6][18] ), .X(n9120) );
  inv_x2_sg U14563 ( .A(n1495), .X(n9100) );
  inv_x2_sg U14564 ( .A(n1497), .X(n9140) );
  inv_x2_sg U14565 ( .A(\i_im[13][19] ), .X(n9181) );
  inv_x2_sg U14566 ( .A(\i_im[12][19] ), .X(n9161) );
  inv_x2_sg U14567 ( .A(\i_im[6][19] ), .X(n9121) );
  inv_x2_sg U14568 ( .A(n1531), .X(n9101) );
  inv_x2_sg U14569 ( .A(n1533), .X(n9141) );
  inv_x2_sg U14570 ( .A(\i_im[13][0] ), .X(n9162) );
  inv_x2_sg U14571 ( .A(\i_im[12][0] ), .X(n9142) );
  inv_x2_sg U14572 ( .A(\i_im[6][0] ), .X(n9102) );
  inv_x2_sg U14573 ( .A(n889), .X(n9082) );
  inv_x2_sg U14574 ( .A(n891), .X(n9122) );
  inv_x2_sg U14575 ( .A(n4299), .X(n9190) );
  inv_x2_sg U14576 ( .A(n3092), .X(n9191) );
  inv_x2_sg U14577 ( .A(n5287), .X(n9202) );
endmodule

